module basic_5000_50000_5000_25_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_2428,In_1038);
xnor U1 (N_1,In_3526,In_2700);
nand U2 (N_2,In_108,In_1985);
nand U3 (N_3,In_1336,In_482);
xor U4 (N_4,In_2063,In_966);
nand U5 (N_5,In_3,In_796);
nand U6 (N_6,In_4248,In_3204);
xnor U7 (N_7,In_2711,In_860);
nand U8 (N_8,In_4400,In_1344);
xor U9 (N_9,In_576,In_10);
nor U10 (N_10,In_3080,In_1927);
nor U11 (N_11,In_4022,In_2698);
nor U12 (N_12,In_124,In_4903);
and U13 (N_13,In_76,In_3769);
nor U14 (N_14,In_2313,In_3466);
and U15 (N_15,In_4988,In_1863);
nand U16 (N_16,In_136,In_4801);
or U17 (N_17,In_2572,In_4729);
and U18 (N_18,In_1899,In_1389);
and U19 (N_19,In_2859,In_4666);
and U20 (N_20,In_4263,In_3103);
nor U21 (N_21,In_1052,In_1683);
nor U22 (N_22,In_3013,In_1312);
nand U23 (N_23,In_3282,In_1579);
or U24 (N_24,In_4236,In_2771);
nand U25 (N_25,In_1201,In_998);
and U26 (N_26,In_67,In_3718);
xnor U27 (N_27,In_3191,In_4255);
xor U28 (N_28,In_658,In_4028);
and U29 (N_29,In_997,In_4846);
xnor U30 (N_30,In_4876,In_148);
xor U31 (N_31,In_1841,In_4900);
or U32 (N_32,In_2520,In_4055);
or U33 (N_33,In_984,In_2420);
and U34 (N_34,In_2389,In_4571);
nor U35 (N_35,In_3572,In_4631);
or U36 (N_36,In_918,In_2286);
and U37 (N_37,In_471,In_4741);
nand U38 (N_38,In_4945,In_1861);
xor U39 (N_39,In_1735,In_1252);
nor U40 (N_40,In_2917,In_773);
nand U41 (N_41,In_2619,In_2676);
nand U42 (N_42,In_2151,In_850);
or U43 (N_43,In_3912,In_4805);
or U44 (N_44,In_4182,In_2235);
and U45 (N_45,In_4396,In_1184);
nand U46 (N_46,In_1070,In_2068);
or U47 (N_47,In_1459,In_1028);
nor U48 (N_48,In_2065,In_2720);
and U49 (N_49,In_2758,In_3594);
nand U50 (N_50,In_1705,In_2967);
nand U51 (N_51,In_3982,In_3322);
nor U52 (N_52,In_4598,In_3570);
nand U53 (N_53,In_1465,In_1462);
or U54 (N_54,In_633,In_3837);
nand U55 (N_55,In_2490,In_3200);
xnor U56 (N_56,In_4551,In_3576);
xnor U57 (N_57,In_528,In_3890);
nand U58 (N_58,In_2494,In_762);
nor U59 (N_59,In_1828,In_1265);
and U60 (N_60,In_1891,In_4362);
xor U61 (N_61,In_3375,In_3688);
nor U62 (N_62,In_4897,In_2245);
and U63 (N_63,In_584,In_2540);
xnor U64 (N_64,In_3008,In_2070);
or U65 (N_65,In_2831,In_331);
nand U66 (N_66,In_421,In_3593);
or U67 (N_67,In_4740,In_3365);
nor U68 (N_68,In_3057,In_4195);
or U69 (N_69,In_3207,In_1109);
nor U70 (N_70,In_2322,In_1138);
or U71 (N_71,In_4008,In_1664);
and U72 (N_72,In_3015,In_1729);
xor U73 (N_73,In_1467,In_1875);
or U74 (N_74,In_4485,In_3488);
or U75 (N_75,In_2949,In_2159);
or U76 (N_76,In_3417,In_1178);
xor U77 (N_77,In_3316,In_503);
nor U78 (N_78,In_155,In_2538);
or U79 (N_79,In_3256,In_4386);
nand U80 (N_80,In_1213,In_434);
or U81 (N_81,In_3739,In_4954);
or U82 (N_82,In_1972,In_853);
and U83 (N_83,In_4976,In_4132);
xor U84 (N_84,In_2039,In_1432);
xor U85 (N_85,In_4483,In_546);
and U86 (N_86,In_4151,In_3762);
nor U87 (N_87,In_771,In_3703);
nor U88 (N_88,In_806,In_1088);
or U89 (N_89,In_2597,In_4616);
xor U90 (N_90,In_4721,In_4218);
nand U91 (N_91,In_3574,In_1097);
nand U92 (N_92,In_3535,In_3896);
nor U93 (N_93,In_1965,In_1236);
or U94 (N_94,In_1297,In_1619);
nand U95 (N_95,In_1352,In_458);
and U96 (N_96,In_2689,In_2109);
or U97 (N_97,In_4374,In_290);
and U98 (N_98,In_1077,In_3064);
and U99 (N_99,In_1505,In_2786);
nand U100 (N_100,In_4313,In_4827);
and U101 (N_101,In_4797,In_3969);
xor U102 (N_102,In_3978,In_1200);
xor U103 (N_103,In_1284,In_4981);
and U104 (N_104,In_1530,In_1751);
or U105 (N_105,In_38,In_4607);
or U106 (N_106,In_942,In_2177);
and U107 (N_107,In_1582,In_3782);
and U108 (N_108,In_3989,In_3351);
nand U109 (N_109,In_2115,In_2731);
or U110 (N_110,In_4944,In_1608);
nor U111 (N_111,In_2249,In_3717);
and U112 (N_112,In_3820,In_4747);
nor U113 (N_113,In_1776,In_4057);
nand U114 (N_114,In_359,In_4231);
nand U115 (N_115,In_4475,In_3454);
nor U116 (N_116,In_3612,In_2537);
nand U117 (N_117,In_2452,In_4704);
and U118 (N_118,In_3496,In_666);
or U119 (N_119,In_478,In_2923);
nand U120 (N_120,In_1924,In_944);
xor U121 (N_121,In_307,In_4720);
xnor U122 (N_122,In_4007,In_3074);
and U123 (N_123,In_3771,In_3025);
and U124 (N_124,In_4591,In_72);
nand U125 (N_125,In_3334,In_334);
nor U126 (N_126,In_1492,In_4117);
xor U127 (N_127,In_4638,In_1062);
or U128 (N_128,In_2475,In_1914);
nor U129 (N_129,In_4665,In_3104);
nand U130 (N_130,In_4509,In_1526);
and U131 (N_131,In_429,In_3900);
nor U132 (N_132,In_817,In_3197);
xor U133 (N_133,In_1158,In_864);
nor U134 (N_134,In_1014,In_232);
nand U135 (N_135,In_2964,In_4404);
and U136 (N_136,In_3285,In_2459);
nor U137 (N_137,In_74,In_3350);
and U138 (N_138,In_1149,In_357);
xnor U139 (N_139,In_4952,In_3391);
xnor U140 (N_140,In_198,In_2843);
xnor U141 (N_141,In_1378,In_2193);
and U142 (N_142,In_4697,In_3323);
and U143 (N_143,In_3471,In_3126);
nor U144 (N_144,In_2305,In_862);
and U145 (N_145,In_4641,In_64);
or U146 (N_146,In_789,In_2295);
and U147 (N_147,In_3487,In_4372);
nand U148 (N_148,In_3947,In_2369);
nand U149 (N_149,In_4548,In_2533);
nand U150 (N_150,In_3419,In_4789);
nand U151 (N_151,In_2519,In_2271);
and U152 (N_152,In_624,In_3066);
nand U153 (N_153,In_2956,In_672);
or U154 (N_154,In_704,In_195);
or U155 (N_155,In_725,In_691);
nor U156 (N_156,In_475,In_3672);
and U157 (N_157,In_3687,In_4558);
or U158 (N_158,In_395,In_3084);
and U159 (N_159,In_4545,In_2837);
nand U160 (N_160,In_423,In_2506);
xnor U161 (N_161,In_3175,In_1280);
and U162 (N_162,In_265,In_3675);
nand U163 (N_163,In_35,In_227);
and U164 (N_164,In_4191,In_2349);
nand U165 (N_165,In_2952,In_1534);
nor U166 (N_166,In_693,In_3650);
nor U167 (N_167,In_2411,In_976);
nor U168 (N_168,In_519,In_3482);
or U169 (N_169,In_2820,In_3783);
and U170 (N_170,In_3225,In_3366);
xor U171 (N_171,In_2114,In_443);
or U172 (N_172,In_3331,In_3445);
xnor U173 (N_173,In_3829,In_4133);
xor U174 (N_174,In_881,In_4680);
nand U175 (N_175,In_48,In_581);
nor U176 (N_176,In_23,In_178);
and U177 (N_177,In_466,In_1671);
nand U178 (N_178,In_4220,In_1339);
xor U179 (N_179,In_690,In_4600);
and U180 (N_180,In_3003,In_1399);
nor U181 (N_181,In_4722,In_4877);
nor U182 (N_182,In_2264,In_4724);
nor U183 (N_183,In_480,In_4399);
nand U184 (N_184,In_3630,In_1003);
nand U185 (N_185,In_4727,In_3426);
nand U186 (N_186,In_2968,In_254);
or U187 (N_187,In_3459,In_1880);
nor U188 (N_188,In_4953,In_608);
xor U189 (N_189,In_266,In_2509);
xnor U190 (N_190,In_3186,In_1262);
or U191 (N_191,In_3621,In_613);
nand U192 (N_192,In_511,In_3228);
xor U193 (N_193,In_1528,In_4268);
nor U194 (N_194,In_462,In_2081);
nand U195 (N_195,In_68,In_4001);
xor U196 (N_196,In_2505,In_1890);
nor U197 (N_197,In_711,In_3307);
nand U198 (N_198,In_406,In_1392);
xnor U199 (N_199,In_4002,In_768);
nor U200 (N_200,In_980,In_464);
nand U201 (N_201,In_3063,In_1700);
nor U202 (N_202,In_4705,In_3690);
nor U203 (N_203,In_2189,In_180);
or U204 (N_204,In_728,In_4995);
or U205 (N_205,In_4502,In_3846);
nand U206 (N_206,In_238,In_3081);
or U207 (N_207,In_2621,In_4452);
nor U208 (N_208,In_901,In_3461);
nor U209 (N_209,In_372,In_1132);
nand U210 (N_210,In_601,In_2291);
nand U211 (N_211,In_2395,In_1907);
and U212 (N_212,In_3423,In_3475);
nand U213 (N_213,In_3595,In_420);
and U214 (N_214,In_3995,In_4425);
xnor U215 (N_215,In_299,In_2231);
or U216 (N_216,In_4364,In_4847);
or U217 (N_217,In_4774,In_2629);
xor U218 (N_218,In_4891,In_1440);
xnor U219 (N_219,In_2528,In_4416);
and U220 (N_220,In_1510,In_2052);
nor U221 (N_221,In_748,In_2672);
nand U222 (N_222,In_866,In_4026);
nand U223 (N_223,In_3588,In_2697);
nor U224 (N_224,In_4025,In_3075);
nand U225 (N_225,In_1045,In_4335);
xnor U226 (N_226,In_1259,In_4758);
nor U227 (N_227,In_2806,In_1299);
nor U228 (N_228,In_1728,In_3754);
or U229 (N_229,In_4235,In_1561);
or U230 (N_230,In_1744,In_4515);
nand U231 (N_231,In_1377,In_49);
xnor U232 (N_232,In_2571,In_2257);
or U233 (N_233,In_3509,In_1699);
nor U234 (N_234,In_3881,In_1823);
nor U235 (N_235,In_15,In_755);
or U236 (N_236,In_3528,In_1214);
and U237 (N_237,In_3270,In_2093);
nand U238 (N_238,In_3242,In_803);
nand U239 (N_239,In_4107,In_4890);
nor U240 (N_240,In_1279,In_2724);
nor U241 (N_241,In_4173,In_547);
nor U242 (N_242,In_3255,In_393);
xnor U243 (N_243,In_2995,In_1591);
nor U244 (N_244,In_4264,In_4111);
nand U245 (N_245,In_4510,In_822);
xor U246 (N_246,In_4042,In_1403);
nor U247 (N_247,In_622,In_535);
nand U248 (N_248,In_3811,In_4683);
or U249 (N_249,In_2875,In_3068);
nand U250 (N_250,In_2604,In_29);
nor U251 (N_251,In_1895,In_2921);
nand U252 (N_252,In_602,In_3831);
xor U253 (N_253,In_2350,In_4837);
nor U254 (N_254,In_1866,In_1177);
and U255 (N_255,In_4463,In_2421);
and U256 (N_256,In_3746,In_1657);
nand U257 (N_257,In_1204,In_2550);
or U258 (N_258,In_4148,In_1100);
xor U259 (N_259,In_2282,In_1405);
xnor U260 (N_260,In_1238,In_1532);
xnor U261 (N_261,In_3462,In_206);
nor U262 (N_262,In_558,In_1305);
nor U263 (N_263,In_3664,In_3230);
xor U264 (N_264,In_4760,In_3363);
nand U265 (N_265,In_3768,In_3458);
or U266 (N_266,In_4474,In_447);
or U267 (N_267,In_109,In_2723);
xnor U268 (N_268,In_589,In_318);
or U269 (N_269,In_1298,In_2973);
and U270 (N_270,In_2429,In_2605);
and U271 (N_271,In_2612,In_673);
xnor U272 (N_272,In_3151,In_1707);
xnor U273 (N_273,In_4381,In_2785);
or U274 (N_274,In_4454,In_4032);
or U275 (N_275,In_2582,In_1600);
nor U276 (N_276,In_1709,In_2325);
xor U277 (N_277,In_1370,In_3681);
and U278 (N_278,In_1529,In_1769);
or U279 (N_279,In_4763,In_2853);
xor U280 (N_280,In_4970,In_1949);
nor U281 (N_281,In_3814,In_2154);
xor U282 (N_282,In_3133,In_708);
or U283 (N_283,In_2330,In_738);
xor U284 (N_284,In_1361,In_1642);
xnor U285 (N_285,In_2918,In_1962);
or U286 (N_286,In_2879,In_1746);
nand U287 (N_287,In_1261,In_3100);
nor U288 (N_288,In_929,In_4085);
or U289 (N_289,In_2176,In_2688);
and U290 (N_290,In_1461,In_4690);
or U291 (N_291,In_2076,In_974);
and U292 (N_292,In_3192,In_2372);
nor U293 (N_293,In_947,In_4045);
xor U294 (N_294,In_1845,In_2061);
or U295 (N_295,In_2890,In_3235);
or U296 (N_296,In_4811,In_2543);
xor U297 (N_297,In_3118,In_2882);
and U298 (N_298,In_4013,In_4599);
nor U299 (N_299,In_2760,In_1417);
nor U300 (N_300,In_2686,In_1614);
nand U301 (N_301,In_4130,In_4071);
xnor U302 (N_302,In_1076,In_3745);
nand U303 (N_303,In_1391,In_1822);
or U304 (N_304,In_3825,In_1601);
or U305 (N_305,In_2609,In_4486);
nor U306 (N_306,In_1548,In_2586);
and U307 (N_307,In_2085,In_2324);
and U308 (N_308,In_4385,In_2825);
xor U309 (N_309,In_4802,In_4979);
xor U310 (N_310,In_698,In_1620);
xnor U311 (N_311,In_2376,In_3592);
and U312 (N_312,In_2574,In_382);
nor U313 (N_313,In_2992,In_3658);
and U314 (N_314,In_931,In_4238);
or U315 (N_315,In_3611,In_1205);
nor U316 (N_316,In_1206,In_2774);
xnor U317 (N_317,In_906,In_2266);
nand U318 (N_318,In_3774,In_3977);
and U319 (N_319,In_3360,In_2393);
nor U320 (N_320,In_3985,In_376);
nor U321 (N_321,In_4612,In_1413);
xnor U322 (N_322,In_4658,In_371);
nor U323 (N_323,In_3110,In_1969);
xnor U324 (N_324,In_4768,In_4818);
nand U325 (N_325,In_3042,In_437);
xnor U326 (N_326,In_1476,In_3301);
xor U327 (N_327,In_1419,In_2352);
xnor U328 (N_328,In_717,In_797);
nor U329 (N_329,In_2818,In_4073);
xnor U330 (N_330,In_1933,In_4896);
nor U331 (N_331,In_3937,In_3413);
and U332 (N_332,In_2536,In_3891);
nor U333 (N_333,In_2573,In_1773);
nor U334 (N_334,In_2892,In_2168);
xor U335 (N_335,In_311,In_3813);
nor U336 (N_336,In_4836,In_1785);
or U337 (N_337,In_1429,In_1315);
and U338 (N_338,In_2768,In_2173);
nor U339 (N_339,In_4426,In_1765);
nor U340 (N_340,In_3262,In_2029);
nor U341 (N_341,In_868,In_284);
nor U342 (N_342,In_410,In_98);
xnor U343 (N_343,In_1627,In_472);
or U344 (N_344,In_1568,In_865);
and U345 (N_345,In_3772,In_4996);
and U346 (N_346,In_4792,In_3260);
nand U347 (N_347,In_879,In_4433);
or U348 (N_348,In_3043,In_4329);
and U349 (N_349,In_4547,In_194);
or U350 (N_350,In_3234,In_248);
and U351 (N_351,In_2951,In_4922);
and U352 (N_352,In_278,In_3652);
nor U353 (N_353,In_3590,In_3116);
nand U354 (N_354,In_1692,In_113);
nand U355 (N_355,In_2394,In_894);
and U356 (N_356,In_3828,In_1320);
nand U357 (N_357,In_4645,In_1073);
and U358 (N_358,In_2759,In_832);
and U359 (N_359,In_4712,In_3495);
xnor U360 (N_360,In_4834,In_1025);
nor U361 (N_361,In_2481,In_3897);
nor U362 (N_362,In_4487,In_1793);
xnor U363 (N_363,In_2371,In_1250);
xnor U364 (N_364,In_183,In_2796);
nand U365 (N_365,In_1595,In_418);
and U366 (N_366,In_1334,In_4135);
nand U367 (N_367,In_4788,In_1975);
and U368 (N_368,In_1862,In_3056);
and U369 (N_369,In_94,In_4140);
nand U370 (N_370,In_1628,In_3129);
nor U371 (N_371,In_3016,In_3170);
nor U372 (N_372,In_2991,In_2466);
nand U373 (N_373,In_4549,In_2026);
xnor U374 (N_374,In_1099,In_2464);
and U375 (N_375,In_645,In_4540);
nand U376 (N_376,In_1128,In_6);
nand U377 (N_377,In_1611,In_1103);
xnor U378 (N_378,In_1428,In_620);
and U379 (N_379,In_653,In_4746);
and U380 (N_380,In_4961,In_4241);
xor U381 (N_381,In_3167,In_3399);
nor U382 (N_382,In_3967,In_4201);
xor U383 (N_383,In_1834,In_4735);
nand U384 (N_384,In_1426,In_1263);
and U385 (N_385,In_2740,In_4);
nand U386 (N_386,In_4933,In_3817);
nand U387 (N_387,In_4920,In_422);
xor U388 (N_388,In_1451,In_4556);
nand U389 (N_389,In_2502,In_808);
or U390 (N_390,In_4706,In_2101);
nand U391 (N_391,In_4951,In_3882);
and U392 (N_392,In_4049,In_722);
nand U393 (N_393,In_4284,In_4770);
xor U394 (N_394,In_2966,In_4643);
and U395 (N_395,In_2083,In_3359);
nor U396 (N_396,In_2685,In_534);
nor U397 (N_397,In_4821,In_4608);
xnor U398 (N_398,In_2055,In_2435);
nor U399 (N_399,In_578,In_4141);
or U400 (N_400,In_3000,In_1065);
xor U401 (N_401,In_4059,In_3758);
nor U402 (N_402,In_1143,In_4478);
nor U403 (N_403,In_1267,In_1498);
nor U404 (N_404,In_4505,In_3032);
and U405 (N_405,In_4446,In_476);
nand U406 (N_406,In_1134,In_1680);
nor U407 (N_407,In_3130,In_4767);
and U408 (N_408,In_3784,In_1704);
nand U409 (N_409,In_2750,In_4159);
nand U410 (N_410,In_1021,In_1954);
nor U411 (N_411,In_1418,In_4577);
or U412 (N_412,In_1035,In_1402);
nand U413 (N_413,In_2874,In_917);
and U414 (N_414,In_4113,In_1763);
xnor U415 (N_415,In_150,In_1775);
and U416 (N_416,In_3429,In_982);
and U417 (N_417,In_978,In_3140);
nand U418 (N_418,In_262,In_4652);
nor U419 (N_419,In_1730,In_2816);
or U420 (N_420,In_3226,In_368);
xnor U421 (N_421,In_4533,In_3617);
or U422 (N_422,In_4795,In_3608);
nor U423 (N_423,In_4866,In_1495);
or U424 (N_424,In_2746,In_1698);
xnor U425 (N_425,In_3373,In_3306);
or U426 (N_426,In_2562,In_3227);
nor U427 (N_427,In_241,In_1108);
and U428 (N_428,In_1988,In_197);
nand U429 (N_429,In_2564,In_2832);
and U430 (N_430,In_1078,In_1805);
and U431 (N_431,In_612,In_3099);
nor U432 (N_432,In_3997,In_3984);
nand U433 (N_433,In_617,In_759);
nor U434 (N_434,In_1264,In_742);
and U435 (N_435,In_1142,In_2222);
nand U436 (N_436,In_45,In_3205);
or U437 (N_437,In_1401,In_2942);
nand U438 (N_438,In_370,In_4237);
and U439 (N_439,In_2687,In_3143);
nand U440 (N_440,In_1013,In_1340);
and U441 (N_441,In_871,In_2294);
xnor U442 (N_442,In_1424,In_712);
and U443 (N_443,In_89,In_2644);
xor U444 (N_444,In_785,In_4434);
nand U445 (N_445,In_4947,In_4278);
and U446 (N_446,In_810,In_3097);
nor U447 (N_447,In_235,In_3524);
and U448 (N_448,In_1871,In_2405);
nand U449 (N_449,In_483,In_285);
and U450 (N_450,In_587,In_1585);
nor U451 (N_451,In_292,In_2955);
nor U452 (N_452,In_4293,In_2699);
or U453 (N_453,In_273,In_4376);
or U454 (N_454,In_1547,In_643);
xor U455 (N_455,In_3686,In_330);
and U456 (N_456,In_3878,In_707);
and U457 (N_457,In_3492,In_2870);
or U458 (N_458,In_1521,In_3453);
nand U459 (N_459,In_3856,In_3292);
xnor U460 (N_460,In_1518,In_134);
and U461 (N_461,In_4112,In_814);
and U462 (N_462,In_3736,In_3190);
or U463 (N_463,In_1112,In_3938);
nand U464 (N_464,In_3932,In_3709);
or U465 (N_465,In_402,In_638);
xor U466 (N_466,In_274,In_3950);
nor U467 (N_467,In_1721,In_3615);
or U468 (N_468,In_4047,In_2463);
nand U469 (N_469,In_2167,In_825);
or U470 (N_470,In_17,In_489);
xnor U471 (N_471,In_3059,In_3533);
xnor U472 (N_472,In_1473,In_1710);
nor U473 (N_473,In_342,In_2410);
xnor U474 (N_474,In_4110,In_3113);
nor U475 (N_475,In_1575,In_3378);
xnor U476 (N_476,In_4560,In_3705);
nand U477 (N_477,In_4030,In_4732);
and U478 (N_478,In_2348,In_3580);
or U479 (N_479,In_2377,In_4249);
nor U480 (N_480,In_267,In_2542);
or U481 (N_481,In_1326,In_3922);
xnor U482 (N_482,In_1295,In_4406);
and U483 (N_483,In_2,In_3780);
nand U484 (N_484,In_4621,In_2517);
and U485 (N_485,In_2983,In_1673);
or U486 (N_486,In_448,In_2355);
nor U487 (N_487,In_2179,In_2808);
or U488 (N_488,In_2353,In_4038);
nand U489 (N_489,In_3659,In_676);
nor U490 (N_490,In_1559,In_2359);
and U491 (N_491,In_1323,In_4629);
nand U492 (N_492,In_1039,In_1053);
or U493 (N_493,In_1507,In_1953);
xnor U494 (N_494,In_1641,In_3402);
nand U495 (N_495,In_2467,In_3520);
and U496 (N_496,In_4367,In_3694);
and U497 (N_497,In_3807,In_3834);
or U498 (N_498,In_996,In_1330);
nand U499 (N_499,In_2862,In_2404);
nand U500 (N_500,In_4108,In_2507);
xor U501 (N_501,In_2653,In_839);
nand U502 (N_502,In_3575,In_1854);
or U503 (N_503,In_415,In_4728);
or U504 (N_504,In_1645,In_1524);
nand U505 (N_505,In_31,In_1755);
nor U506 (N_506,In_4627,In_1364);
nand U507 (N_507,In_2777,In_4336);
or U508 (N_508,In_4017,In_360);
xnor U509 (N_509,In_3787,In_1324);
nor U510 (N_510,In_348,In_1269);
nor U511 (N_511,In_2239,In_4080);
and U512 (N_512,In_2113,In_3530);
and U513 (N_513,In_692,In_2782);
xnor U514 (N_514,In_3855,In_4005);
xnor U515 (N_515,In_14,In_1980);
nor U516 (N_516,In_4290,In_3936);
xor U517 (N_517,In_1906,In_3869);
and U518 (N_518,In_3398,In_4227);
xnor U519 (N_519,In_70,In_1555);
or U520 (N_520,In_4941,In_1463);
nand U521 (N_521,In_1190,In_3567);
xor U522 (N_522,In_1054,In_4754);
or U523 (N_523,In_4775,In_3654);
xor U524 (N_524,In_3779,In_510);
xnor U525 (N_525,In_607,In_2584);
nor U526 (N_526,In_3302,In_3765);
xnor U527 (N_527,In_1569,In_4757);
xnor U528 (N_528,In_4084,In_438);
or U529 (N_529,In_615,In_2012);
or U530 (N_530,In_2719,In_3430);
or U531 (N_531,In_473,In_3409);
xnor U532 (N_532,In_276,In_536);
and U533 (N_533,In_4345,In_4437);
and U534 (N_534,In_1359,In_4495);
xnor U535 (N_535,In_1002,In_4966);
and U536 (N_536,In_2171,In_4831);
nand U537 (N_537,In_3436,In_4554);
nor U538 (N_538,In_1126,In_512);
xor U539 (N_539,In_1592,In_219);
or U540 (N_540,In_3879,In_971);
xor U541 (N_541,In_1260,In_1101);
or U542 (N_542,In_3054,In_1797);
nand U543 (N_543,In_2296,In_4192);
and U544 (N_544,In_4880,In_4127);
xnor U545 (N_545,In_3468,In_2362);
or U546 (N_546,In_973,In_3538);
and U547 (N_547,In_2111,In_455);
or U548 (N_548,In_4524,In_399);
nand U549 (N_549,In_4851,In_2197);
xnor U550 (N_550,In_1898,In_205);
and U551 (N_551,In_4442,In_2835);
xor U552 (N_552,In_1543,In_1310);
or U553 (N_553,In_4765,In_3564);
xnor U554 (N_554,In_250,In_3465);
and U555 (N_555,In_3906,In_3741);
nand U556 (N_556,In_353,In_4174);
or U557 (N_557,In_2137,In_247);
or U558 (N_558,In_2157,In_1430);
xor U559 (N_559,In_2329,In_1929);
and U560 (N_560,In_3128,In_2513);
nor U561 (N_561,In_3962,In_2195);
nor U562 (N_562,In_1092,In_3925);
and U563 (N_563,In_577,In_4092);
or U564 (N_564,In_1839,In_4413);
or U565 (N_565,In_2799,In_4019);
nand U566 (N_566,In_3691,In_4178);
and U567 (N_567,In_2664,In_4356);
or U568 (N_568,In_3823,In_3491);
nand U569 (N_569,In_963,In_1852);
or U570 (N_570,In_1123,In_3483);
or U571 (N_571,In_1477,In_3737);
nand U572 (N_572,In_1423,In_363);
nor U573 (N_573,In_2909,In_4303);
nor U574 (N_574,In_3288,In_1990);
nor U575 (N_575,In_4445,In_4275);
and U576 (N_576,In_1516,In_2891);
nor U577 (N_577,In_1395,In_1882);
or U578 (N_578,In_1672,In_701);
or U579 (N_579,In_182,In_338);
and U580 (N_580,In_1131,In_4883);
xnor U581 (N_581,In_4461,In_1064);
and U582 (N_582,In_1122,In_3173);
and U583 (N_583,In_2000,In_4294);
xor U584 (N_584,In_4776,In_3384);
and U585 (N_585,In_3719,In_2846);
nand U586 (N_586,In_3435,In_1621);
xor U587 (N_587,In_675,In_4274);
and U588 (N_588,In_1527,In_3086);
or U589 (N_589,In_3909,In_211);
nor U590 (N_590,In_1009,In_4835);
and U591 (N_591,In_3707,In_2062);
nand U592 (N_592,In_3928,In_110);
or U593 (N_593,In_2960,In_1111);
nand U594 (N_594,In_1512,In_3271);
or U595 (N_595,In_3711,In_4800);
xor U596 (N_596,In_4196,In_2456);
and U597 (N_597,In_391,In_1400);
and U598 (N_598,In_441,In_3805);
and U599 (N_599,In_263,In_3892);
xor U600 (N_600,In_1872,In_4193);
xnor U601 (N_601,In_2181,In_4440);
and U602 (N_602,In_4402,In_4156);
xor U603 (N_603,In_2673,In_1874);
or U604 (N_604,In_2226,In_345);
nand U605 (N_605,In_3497,In_823);
xnor U606 (N_606,In_189,In_3467);
and U607 (N_607,In_1172,In_765);
nor U608 (N_608,In_2031,In_3427);
nand U609 (N_609,In_829,In_4096);
or U610 (N_610,In_1369,In_132);
nor U611 (N_611,In_1993,In_4428);
nor U612 (N_612,In_3631,In_568);
nor U613 (N_613,In_890,In_114);
or U614 (N_614,In_3254,In_1778);
nand U615 (N_615,In_1311,In_1230);
nor U616 (N_616,In_948,In_2416);
and U617 (N_617,In_3558,In_4999);
or U618 (N_618,In_553,In_4341);
xor U619 (N_619,In_4856,In_4992);
nand U620 (N_620,In_2237,In_2522);
or U621 (N_621,In_2267,In_2259);
and U622 (N_622,In_4771,In_4163);
xor U623 (N_623,In_2896,In_401);
nand U624 (N_624,In_2941,In_3845);
nor U625 (N_625,In_428,In_1638);
nor U626 (N_626,In_3806,In_304);
xor U627 (N_627,In_752,In_1435);
nor U628 (N_628,In_1337,In_1317);
xor U629 (N_629,In_2086,In_2826);
or U630 (N_630,In_4798,In_679);
and U631 (N_631,In_4285,In_1162);
or U632 (N_632,In_4686,In_1454);
and U633 (N_633,In_3006,In_4230);
or U634 (N_634,In_1846,In_3797);
nor U635 (N_635,In_264,In_446);
xnor U636 (N_636,In_1282,In_3740);
nand U637 (N_637,In_2493,In_4081);
xnor U638 (N_638,In_1331,In_1702);
and U639 (N_639,In_1174,In_2219);
nand U640 (N_640,In_4414,In_3889);
and U641 (N_641,In_756,In_315);
or U642 (N_642,In_1541,In_2311);
xor U643 (N_643,In_4459,In_2737);
nand U644 (N_644,In_3637,In_326);
or U645 (N_645,In_3087,In_2342);
or U646 (N_646,In_2860,In_4764);
or U647 (N_647,In_2788,In_2281);
nor U648 (N_648,In_3550,In_2095);
and U649 (N_649,In_3863,In_2972);
nand U650 (N_650,In_1163,In_3276);
nand U651 (N_651,In_463,In_3602);
nor U652 (N_652,In_4601,In_4910);
nor U653 (N_653,In_2850,In_1387);
xor U654 (N_654,In_4347,In_706);
and U655 (N_655,In_660,In_2089);
xor U656 (N_656,In_216,In_2308);
xnor U657 (N_657,In_2628,In_930);
nand U658 (N_658,In_4939,In_603);
and U659 (N_659,In_3677,In_3604);
nand U660 (N_660,In_4817,In_3955);
or U661 (N_661,In_4407,In_1093);
and U662 (N_662,In_1464,In_844);
nor U663 (N_663,In_637,In_4338);
xor U664 (N_664,In_4252,In_1644);
nor U665 (N_665,In_2284,In_1074);
nand U666 (N_666,In_2990,In_1791);
nor U667 (N_667,In_4618,In_4708);
nand U668 (N_668,In_3094,In_457);
nand U669 (N_669,In_249,In_4279);
nor U670 (N_670,In_1246,In_3561);
nand U671 (N_671,In_2225,In_187);
nor U672 (N_672,In_2883,In_3424);
xnor U673 (N_673,In_3727,In_3810);
and U674 (N_674,In_1363,In_3603);
nor U675 (N_675,In_3786,In_2255);
and U676 (N_676,In_4094,In_3376);
or U677 (N_677,In_3935,In_2684);
or U678 (N_678,In_1767,In_1919);
xor U679 (N_679,In_4480,In_4879);
or U680 (N_680,In_4403,In_2632);
nor U681 (N_681,In_4990,In_1788);
and U682 (N_682,In_596,In_4626);
nand U683 (N_683,In_2930,In_3924);
nor U684 (N_684,In_1889,In_1982);
nor U685 (N_685,In_3345,In_951);
and U686 (N_686,In_2122,In_2848);
and U687 (N_687,In_1313,In_3903);
or U688 (N_688,In_3265,In_3940);
nor U689 (N_689,In_757,In_1571);
nand U690 (N_690,In_4848,In_8);
or U691 (N_691,In_1651,In_2501);
or U692 (N_692,In_2096,In_449);
and U693 (N_693,In_4962,In_656);
and U694 (N_694,In_1583,In_3387);
and U695 (N_695,In_3809,In_4497);
and U696 (N_696,In_3318,In_1346);
nand U697 (N_697,In_169,In_4370);
nand U698 (N_698,In_2491,In_525);
and U699 (N_699,In_119,In_3648);
and U700 (N_700,In_898,In_1833);
and U701 (N_701,In_644,In_1300);
or U702 (N_702,In_572,In_2828);
nor U703 (N_703,In_2477,In_799);
xnor U704 (N_704,In_3125,In_234);
nor U705 (N_705,In_2561,In_4872);
nand U706 (N_706,In_2567,In_3134);
or U707 (N_707,In_775,In_2473);
or U708 (N_708,In_641,In_3613);
xor U709 (N_709,In_3716,In_1968);
or U710 (N_710,In_3851,In_2006);
and U711 (N_711,In_1383,In_3320);
or U712 (N_712,In_459,In_4000);
xnor U713 (N_713,In_4508,In_935);
or U714 (N_714,In_1987,In_3872);
xnor U715 (N_715,In_3181,In_3330);
nand U716 (N_716,In_2732,In_4889);
or U717 (N_717,In_3770,In_2140);
and U718 (N_718,In_4752,In_1681);
nor U719 (N_719,In_1124,In_3643);
and U720 (N_720,In_1817,In_4301);
and U721 (N_721,In_4761,In_4098);
or U722 (N_722,In_561,In_1589);
and U723 (N_723,In_2110,In_4168);
nor U724 (N_724,In_222,In_377);
nor U725 (N_725,In_229,In_936);
nor U726 (N_726,In_2149,In_2367);
or U727 (N_727,In_914,In_256);
xor U728 (N_728,In_3679,In_1653);
nor U729 (N_729,In_2382,In_3852);
and U730 (N_730,In_635,In_1165);
nor U731 (N_731,In_888,In_579);
xor U732 (N_732,In_492,In_3923);
and U733 (N_733,In_3165,In_3832);
or U734 (N_734,In_4124,In_4965);
xor U735 (N_735,In_2585,In_3039);
nor U736 (N_736,In_3553,In_1256);
nand U737 (N_737,In_2734,In_2422);
xnor U738 (N_738,In_3871,In_3512);
and U739 (N_739,In_2498,In_2439);
xor U740 (N_740,In_3152,In_3542);
nand U741 (N_741,In_3519,In_2557);
or U742 (N_742,In_2797,In_361);
nor U743 (N_743,In_2015,In_4439);
and U744 (N_744,In_3343,In_3115);
xnor U745 (N_745,In_2657,In_2166);
or U746 (N_746,In_3002,In_4075);
or U747 (N_747,In_3362,In_2965);
nor U748 (N_748,In_1740,In_3958);
nand U749 (N_749,In_3875,In_2978);
and U750 (N_750,In_975,In_257);
nand U751 (N_751,In_3021,In_2499);
and U752 (N_752,In_3822,In_2705);
xor U753 (N_753,In_958,In_3842);
and U754 (N_754,In_2958,In_4684);
and U755 (N_755,In_3213,In_3827);
xor U756 (N_756,In_2979,In_782);
nand U757 (N_757,In_3712,In_2046);
nor U758 (N_758,In_50,In_1923);
nor U759 (N_759,In_2642,In_4572);
nor U760 (N_760,In_1581,In_4089);
and U761 (N_761,In_1106,In_875);
nand U762 (N_762,In_4887,In_3112);
xnor U763 (N_763,In_4467,In_995);
or U764 (N_764,In_1042,In_4239);
nor U765 (N_765,In_3193,In_880);
nand U766 (N_766,In_2695,In_517);
nor U767 (N_767,In_833,In_1905);
and U768 (N_768,In_1639,In_1037);
or U769 (N_769,In_2392,In_2982);
and U770 (N_770,In_1234,In_1048);
xnor U771 (N_771,In_2858,In_3551);
and U772 (N_772,In_3437,In_1316);
or U773 (N_773,In_2280,In_4546);
and U774 (N_774,In_4593,In_4873);
or U775 (N_775,In_3026,In_1795);
xnor U776 (N_776,In_1257,In_2224);
or U777 (N_777,In_3494,In_97);
nor U778 (N_778,In_129,In_404);
nand U779 (N_779,In_4544,In_899);
nor U780 (N_780,In_4186,In_987);
and U781 (N_781,In_3513,In_1691);
nand U782 (N_782,In_964,In_2327);
nand U783 (N_783,In_2648,In_3421);
nand U784 (N_784,In_362,In_4035);
and U785 (N_785,In_3224,In_3960);
nor U786 (N_786,In_807,In_920);
nor U787 (N_787,In_4689,In_2943);
and U788 (N_788,In_4520,In_2485);
xor U789 (N_789,In_389,In_674);
nor U790 (N_790,In_2823,In_33);
and U791 (N_791,In_4450,In_2023);
nand U792 (N_792,In_2639,In_1629);
nand U793 (N_793,In_4649,In_1222);
or U794 (N_794,In_2040,In_1441);
xor U795 (N_795,In_3743,In_240);
nor U796 (N_796,In_156,In_417);
nand U797 (N_797,In_1695,In_1393);
nand U798 (N_798,In_498,In_1910);
or U799 (N_799,In_2442,In_4346);
xor U800 (N_800,In_4254,In_4589);
nor U801 (N_801,In_2869,In_1753);
or U802 (N_802,In_495,In_2011);
xnor U803 (N_803,In_1565,In_2091);
nor U804 (N_804,In_4436,In_4020);
xor U805 (N_805,In_2641,In_4304);
nor U806 (N_806,In_2508,In_12);
xor U807 (N_807,In_726,In_4250);
or U808 (N_808,In_2139,In_2622);
nand U809 (N_809,In_3038,In_4432);
and U810 (N_810,In_2233,In_1576);
or U811 (N_811,In_1538,In_1026);
nand U812 (N_812,In_4102,In_85);
or U813 (N_813,In_4575,In_2474);
nand U814 (N_814,In_3324,In_1113);
nand U815 (N_815,In_820,In_2764);
xor U816 (N_816,In_3163,In_3266);
nand U817 (N_817,In_3905,In_4188);
nand U818 (N_818,In_403,In_4916);
or U819 (N_819,In_1915,In_477);
nand U820 (N_820,In_4663,In_977);
xnor U821 (N_821,In_665,In_2492);
or U822 (N_822,In_199,In_2587);
xor U823 (N_823,In_2364,In_764);
xor U824 (N_824,In_1209,In_583);
and U825 (N_825,In_488,In_3154);
nand U826 (N_826,In_4354,In_4868);
xor U827 (N_827,In_1032,In_3372);
xor U828 (N_828,In_2710,In_4871);
nor U829 (N_829,In_723,In_2613);
nor U830 (N_830,In_3798,In_908);
nor U831 (N_831,In_3245,In_1116);
nor U832 (N_832,In_2836,In_3660);
xnor U833 (N_833,In_4060,In_4050);
nor U834 (N_834,In_3916,In_123);
or U835 (N_835,In_1349,In_2135);
nand U836 (N_836,In_461,In_2635);
or U837 (N_837,In_2773,In_1244);
or U838 (N_838,In_3114,In_2565);
nor U839 (N_839,In_804,In_1500);
xor U840 (N_840,In_1155,In_1754);
and U841 (N_841,In_960,In_3329);
nor U842 (N_842,In_2713,In_1741);
nand U843 (N_843,In_2516,In_3532);
nand U844 (N_844,In_151,In_4041);
or U845 (N_845,In_3747,In_1870);
nand U846 (N_846,In_4300,In_2931);
or U847 (N_847,In_3107,In_2008);
nor U848 (N_848,In_3221,In_4937);
nand U849 (N_849,In_2050,In_26);
and U850 (N_850,In_4718,In_3973);
nand U851 (N_851,In_2576,In_4843);
nand U852 (N_852,In_4410,In_1570);
or U853 (N_853,In_3815,In_705);
and U854 (N_854,In_4785,In_2273);
nor U855 (N_855,In_2449,In_1125);
and U856 (N_856,In_1096,In_3579);
and U857 (N_857,In_4408,In_2331);
nand U858 (N_858,In_1615,In_2019);
xor U859 (N_859,In_62,In_78);
nor U860 (N_860,In_3250,In_317);
or U861 (N_861,In_3569,In_1090);
and U862 (N_862,In_3011,In_487);
xnor U863 (N_863,In_1414,In_2326);
nor U864 (N_864,In_2155,In_3247);
nor U865 (N_865,In_3589,In_4647);
or U866 (N_866,In_703,In_3346);
xnor U867 (N_867,In_1715,In_766);
or U868 (N_868,In_2341,In_2560);
or U869 (N_869,In_2887,In_2614);
or U870 (N_870,In_714,In_4234);
nor U871 (N_871,In_694,In_2811);
nor U872 (N_872,In_1545,In_2361);
nand U873 (N_873,In_3433,In_1787);
and U874 (N_874,In_4128,In_2150);
xor U875 (N_875,In_2100,In_835);
xnor U876 (N_876,In_2142,In_1289);
nand U877 (N_877,In_1801,In_514);
nor U878 (N_878,In_3390,In_813);
or U879 (N_879,In_2704,In_1276);
xnor U880 (N_880,In_2589,In_4153);
or U881 (N_881,In_4395,In_2899);
or U882 (N_882,In_545,In_3370);
nand U883 (N_883,In_3258,In_444);
and U884 (N_884,In_1347,In_2174);
or U885 (N_885,In_40,In_4855);
and U886 (N_886,In_128,In_1368);
nand U887 (N_887,In_513,In_3281);
xor U888 (N_888,In_1977,In_4715);
xnor U889 (N_889,In_1777,In_2527);
nand U890 (N_890,In_4913,In_1693);
nand U891 (N_891,In_597,In_3952);
xor U892 (N_892,In_309,In_210);
and U893 (N_893,In_1602,In_4031);
nand U894 (N_894,In_2976,In_2725);
and U895 (N_895,In_1792,In_852);
nand U896 (N_896,In_1437,In_837);
or U897 (N_897,In_4911,In_2380);
nor U898 (N_898,In_700,In_1273);
and U899 (N_899,In_4091,In_2932);
or U900 (N_900,In_4208,In_226);
xor U901 (N_901,In_2360,In_1335);
xor U902 (N_902,In_909,In_3671);
or U903 (N_903,In_3994,In_3439);
nor U904 (N_904,In_1223,In_2601);
nor U905 (N_905,In_1883,In_4762);
nand U906 (N_906,In_486,In_4430);
xor U907 (N_907,In_2742,In_2462);
or U908 (N_908,In_1502,In_1199);
xnor U909 (N_909,In_889,In_1218);
xnor U910 (N_910,In_439,In_1390);
and U911 (N_911,In_2146,In_1770);
and U912 (N_912,In_1407,In_481);
and U913 (N_913,In_4950,In_4247);
and U914 (N_914,In_689,In_3644);
or U915 (N_915,In_2486,In_88);
and U916 (N_916,In_3839,In_2077);
and U917 (N_917,In_1061,In_3357);
nor U918 (N_918,In_0,In_145);
or U919 (N_919,In_1703,In_4882);
nand U920 (N_920,In_1160,In_147);
nor U921 (N_921,In_533,In_3178);
nor U922 (N_922,In_1268,In_3642);
and U923 (N_923,In_1203,In_3527);
nand U924 (N_924,In_2876,In_2004);
nor U925 (N_925,In_2128,In_910);
xnor U926 (N_926,In_3522,In_2242);
or U927 (N_927,In_2524,In_3760);
nor U928 (N_928,In_3641,In_1040);
and U929 (N_929,In_3943,In_560);
nor U930 (N_930,In_4541,In_2530);
nor U931 (N_931,In_2470,In_2407);
xor U932 (N_932,In_2079,In_4125);
xnor U933 (N_933,In_3674,In_303);
nand U934 (N_934,In_751,In_4187);
or U935 (N_935,In_381,In_818);
or U936 (N_936,In_3188,In_4242);
xor U937 (N_937,In_2945,In_3884);
xnor U938 (N_938,In_2221,In_3986);
nand U939 (N_939,In_4157,In_1365);
or U940 (N_940,In_2716,In_4066);
nand U941 (N_941,In_569,In_2243);
nand U942 (N_942,In_527,In_4202);
or U943 (N_943,In_4716,In_4088);
xnor U944 (N_944,In_2677,In_501);
xor U945 (N_945,In_1007,In_4412);
xor U946 (N_946,In_2454,In_1519);
and U947 (N_947,In_3277,In_4368);
or U948 (N_948,In_2388,In_190);
and U949 (N_949,In_2413,In_3199);
nand U950 (N_950,In_2715,In_800);
and U951 (N_951,In_2595,In_1167);
nand U952 (N_952,In_3479,In_2440);
nand U953 (N_953,In_4742,In_3079);
and U954 (N_954,In_1327,In_3452);
nand U955 (N_955,In_1372,In_1921);
nand U956 (N_956,In_538,In_2599);
xor U957 (N_957,In_3085,In_4429);
xnor U958 (N_958,In_3972,In_786);
or U959 (N_959,In_4901,In_4845);
nand U960 (N_960,In_983,In_142);
nor U961 (N_961,In_2339,In_1098);
nor U962 (N_962,In_1503,In_3795);
or U963 (N_963,In_787,In_499);
or U964 (N_964,In_1540,In_1016);
or U965 (N_965,In_2824,In_2333);
nand U966 (N_966,In_4122,In_671);
or U967 (N_967,In_2545,In_61);
nand U968 (N_968,In_286,In_223);
and U969 (N_969,In_1981,In_3578);
or U970 (N_970,In_1609,In_979);
nor U971 (N_971,In_3629,In_4969);
nor U972 (N_972,In_911,In_3730);
or U973 (N_973,In_4244,In_34);
nand U974 (N_974,In_1558,In_1633);
and U975 (N_975,In_2606,In_2541);
nand U976 (N_976,In_2521,In_1553);
and U977 (N_977,In_2415,In_4198);
xnor U978 (N_978,In_1271,In_3560);
nor U979 (N_979,In_2201,In_2911);
and U980 (N_980,In_1853,In_1958);
xor U981 (N_981,In_2489,In_1825);
and U982 (N_982,In_4333,In_3504);
nand U983 (N_983,In_3308,In_2121);
nand U984 (N_984,In_4806,In_3187);
nor U985 (N_985,In_349,In_2772);
nor U986 (N_986,In_319,In_1457);
xnor U987 (N_987,In_1136,In_200);
xor U988 (N_988,In_427,In_4009);
xnor U989 (N_989,In_3867,In_1251);
nor U990 (N_990,In_1747,In_1303);
nand U991 (N_991,In_4317,In_4726);
and U992 (N_992,In_2262,In_614);
or U993 (N_993,In_1759,In_4525);
xor U994 (N_994,In_4259,In_4793);
xor U995 (N_995,In_1974,In_4314);
nand U996 (N_996,In_4422,In_4782);
nor U997 (N_997,In_4339,In_4946);
nand U998 (N_998,In_396,In_2770);
and U999 (N_999,In_4126,In_2336);
xnor U1000 (N_1000,In_91,In_3700);
nand U1001 (N_1001,In_4070,In_3866);
nand U1002 (N_1002,In_3489,In_588);
nand U1003 (N_1003,In_1375,In_699);
nand U1004 (N_1004,In_327,In_1019);
nor U1005 (N_1005,In_2379,In_1536);
nor U1006 (N_1006,In_4309,In_2867);
or U1007 (N_1007,In_3544,In_3833);
xnor U1008 (N_1008,In_4155,In_1436);
or U1009 (N_1009,In_3731,In_369);
xor U1010 (N_1010,In_2981,In_277);
or U1011 (N_1011,In_3177,In_1597);
nor U1012 (N_1012,In_2781,In_4318);
and U1013 (N_1013,In_2626,In_2138);
nor U1014 (N_1014,In_111,In_3744);
xor U1015 (N_1015,In_37,In_3921);
xor U1016 (N_1016,In_3666,In_3121);
nor U1017 (N_1017,In_1858,In_2730);
and U1018 (N_1018,In_2183,In_2714);
or U1019 (N_1019,In_43,In_3680);
xnor U1020 (N_1020,In_4869,In_1318);
xor U1021 (N_1021,In_2256,In_4418);
nand U1022 (N_1022,In_424,In_221);
or U1023 (N_1023,In_3438,In_3953);
nand U1024 (N_1024,In_4606,In_1694);
and U1025 (N_1025,In_4421,In_3470);
nand U1026 (N_1026,In_2417,In_2054);
and U1027 (N_1027,In_4029,In_1830);
and U1028 (N_1028,In_668,In_4907);
or U1029 (N_1029,In_2302,In_312);
xor U1030 (N_1030,In_956,In_177);
or U1031 (N_1031,In_1598,In_4894);
nor U1032 (N_1032,In_333,In_484);
nand U1033 (N_1033,In_55,In_609);
or U1034 (N_1034,In_3348,In_2908);
xnor U1035 (N_1035,In_873,In_4640);
xnor U1036 (N_1036,In_225,In_339);
nor U1037 (N_1037,In_181,In_2679);
and U1038 (N_1038,In_3729,In_32);
nand U1039 (N_1039,In_3088,In_937);
or U1040 (N_1040,In_1187,In_101);
xnor U1041 (N_1041,In_1067,In_4322);
nor U1042 (N_1042,In_4710,In_4003);
or U1043 (N_1043,In_2265,In_968);
or U1044 (N_1044,In_3328,In_2215);
xor U1045 (N_1045,In_4200,In_778);
xor U1046 (N_1046,In_1995,In_2901);
xor U1047 (N_1047,In_3505,In_959);
xor U1048 (N_1048,In_3315,In_1034);
and U1049 (N_1049,In_1147,In_4243);
and U1050 (N_1050,In_2912,In_2568);
xor U1051 (N_1051,In_2652,In_3808);
or U1052 (N_1052,In_280,In_4576);
nor U1053 (N_1053,In_4681,In_2903);
or U1054 (N_1054,In_2810,In_1525);
nand U1055 (N_1055,In_4115,In_3628);
and U1056 (N_1056,In_3127,In_3614);
nor U1057 (N_1057,In_858,In_3093);
xnor U1058 (N_1058,In_1737,In_636);
xor U1059 (N_1059,In_4701,In_2511);
nor U1060 (N_1060,In_2696,In_2726);
nand U1061 (N_1061,In_159,In_4678);
xor U1062 (N_1062,In_2252,In_4468);
and U1063 (N_1063,In_1843,In_2987);
and U1064 (N_1064,In_3785,In_2461);
or U1065 (N_1065,In_1357,In_592);
and U1066 (N_1066,In_1197,In_3061);
or U1067 (N_1067,In_2400,In_604);
or U1068 (N_1068,In_1024,In_4619);
nand U1069 (N_1069,In_41,In_715);
nor U1070 (N_1070,In_688,In_1183);
and U1071 (N_1071,In_4930,In_1900);
nand U1072 (N_1072,In_2757,In_734);
xor U1073 (N_1073,In_1388,In_2335);
and U1074 (N_1074,In_1,In_105);
or U1075 (N_1075,In_2791,In_4532);
nor U1076 (N_1076,In_4331,In_4978);
nor U1077 (N_1077,In_294,In_4943);
or U1078 (N_1078,In_1934,In_1957);
nor U1079 (N_1079,In_2894,In_1665);
nand U1080 (N_1080,In_1838,In_4685);
and U1081 (N_1081,In_1056,In_2934);
xnor U1082 (N_1082,In_571,In_244);
nand U1083 (N_1083,In_2058,In_1782);
and U1084 (N_1084,In_3486,In_3689);
or U1085 (N_1085,In_1104,In_4648);
and U1086 (N_1086,In_2194,In_664);
nor U1087 (N_1087,In_1491,In_485);
or U1088 (N_1088,In_2136,In_903);
and U1089 (N_1089,In_1000,In_1714);
xnor U1090 (N_1090,In_4567,In_293);
or U1091 (N_1091,In_4447,In_1903);
or U1092 (N_1092,In_4858,In_2504);
and U1093 (N_1093,In_4676,In_3102);
or U1094 (N_1094,In_2925,In_2145);
and U1095 (N_1095,In_474,In_1684);
and U1096 (N_1096,In_1573,In_3956);
nand U1097 (N_1097,In_3300,In_1140);
or U1098 (N_1098,In_1046,In_933);
nand U1099 (N_1099,In_2549,In_760);
and U1100 (N_1100,In_1994,In_2794);
or U1101 (N_1101,In_3998,In_3201);
xor U1102 (N_1102,In_2112,In_3232);
xor U1103 (N_1103,In_2650,In_460);
nor U1104 (N_1104,In_3835,In_3485);
nor U1105 (N_1105,In_1637,In_1739);
or U1106 (N_1106,In_2118,In_4632);
nand U1107 (N_1107,In_1724,In_4012);
nor U1108 (N_1108,In_1515,In_4968);
nand U1109 (N_1109,In_4435,In_2938);
or U1110 (N_1110,In_3325,In_3920);
and U1111 (N_1111,In_2753,In_3493);
nor U1112 (N_1112,In_1725,In_1367);
and U1113 (N_1113,In_2532,In_834);
nand U1114 (N_1114,In_1373,In_961);
and U1115 (N_1115,In_3991,In_4702);
nor U1116 (N_1116,In_1355,In_2002);
nor U1117 (N_1117,In_1946,In_2003);
nor U1118 (N_1118,In_3469,In_2778);
nand U1119 (N_1119,In_2847,In_1376);
xnor U1120 (N_1120,In_3076,In_1469);
or U1121 (N_1121,In_2312,In_780);
or U1122 (N_1122,In_2555,In_630);
xnor U1123 (N_1123,In_4330,In_3894);
or U1124 (N_1124,In_1001,In_366);
nand U1125 (N_1125,In_3010,In_4511);
and U1126 (N_1126,In_1291,In_502);
or U1127 (N_1127,In_907,In_4893);
and U1128 (N_1128,In_1416,In_523);
and U1129 (N_1129,In_3510,In_4097);
xor U1130 (N_1130,In_1999,In_4065);
or U1131 (N_1131,In_2132,In_2985);
nor U1132 (N_1132,In_75,In_1050);
or U1133 (N_1133,In_3416,In_4219);
or U1134 (N_1134,In_2354,In_1800);
nor U1135 (N_1135,In_2733,In_122);
nor U1136 (N_1136,In_941,In_1170);
and U1137 (N_1137,In_683,In_4453);
or U1138 (N_1138,In_82,In_4646);
and U1139 (N_1139,In_4984,In_2346);
or U1140 (N_1140,In_4583,In_2678);
or U1141 (N_1141,In_4018,In_3383);
nand U1142 (N_1142,In_3017,In_3649);
and U1143 (N_1143,In_1533,In_1146);
nand U1144 (N_1144,In_2317,In_1186);
nor U1145 (N_1145,In_3927,In_4905);
and U1146 (N_1146,In_3206,In_4784);
or U1147 (N_1147,In_388,In_2946);
and U1148 (N_1148,In_4323,In_2680);
nor U1149 (N_1149,In_3159,In_1850);
nand U1150 (N_1150,In_3028,In_3293);
nor U1151 (N_1151,In_3632,In_237);
xor U1152 (N_1152,In_1066,In_2366);
or U1153 (N_1153,In_130,In_4251);
or U1154 (N_1154,In_1063,In_314);
and U1155 (N_1155,In_876,In_1102);
or U1156 (N_1156,In_2274,In_1697);
nand U1157 (N_1157,In_4384,In_2230);
xnor U1158 (N_1158,In_3065,In_4310);
nor U1159 (N_1159,In_3158,In_2074);
nor U1160 (N_1160,In_4812,In_4458);
and U1161 (N_1161,In_1231,In_1338);
xor U1162 (N_1162,In_3706,In_3053);
or U1163 (N_1163,In_2301,In_158);
nand U1164 (N_1164,In_2199,In_669);
nor U1165 (N_1165,In_3406,In_573);
xor U1166 (N_1166,In_2172,In_4603);
and U1167 (N_1167,In_4865,In_246);
nor U1168 (N_1168,In_3172,In_4733);
or U1169 (N_1169,In_4620,In_4912);
or U1170 (N_1170,In_1410,In_1277);
xnor U1171 (N_1171,In_2546,In_22);
and U1172 (N_1172,In_4743,In_4361);
xor U1173 (N_1173,In_1117,In_1577);
and U1174 (N_1174,In_176,In_4014);
and U1175 (N_1175,In_1151,In_3041);
xnor U1176 (N_1176,In_4053,In_716);
nor U1177 (N_1177,In_4500,In_554);
nor U1178 (N_1178,In_4635,In_4024);
nor U1179 (N_1179,In_1008,In_283);
or U1180 (N_1180,In_3014,In_905);
nor U1181 (N_1181,In_526,In_3150);
and U1182 (N_1182,In_1175,In_2399);
and U1183 (N_1183,In_3939,In_4477);
nand U1184 (N_1184,In_591,In_1425);
and U1185 (N_1185,In_4755,In_4469);
and U1186 (N_1186,In_928,In_3342);
or U1187 (N_1187,In_2953,In_4291);
xor U1188 (N_1188,In_3119,In_1687);
xnor U1189 (N_1189,In_2607,In_3356);
nor U1190 (N_1190,In_153,In_4830);
or U1191 (N_1191,In_3870,In_3915);
xor U1192 (N_1192,In_4653,In_3546);
nand U1193 (N_1193,In_287,In_3304);
nand U1194 (N_1194,In_2103,In_3676);
or U1195 (N_1195,In_2299,In_2084);
or U1196 (N_1196,In_2743,In_470);
and U1197 (N_1197,In_1827,In_3942);
or U1198 (N_1198,In_1790,In_300);
and U1199 (N_1199,In_2974,In_1036);
or U1200 (N_1200,In_3819,In_2658);
nand U1201 (N_1201,In_3537,In_2214);
xnor U1202 (N_1202,In_2547,In_729);
or U1203 (N_1203,In_2258,In_4034);
xor U1204 (N_1204,In_3992,In_4949);
nand U1205 (N_1205,In_2304,In_3153);
nor U1206 (N_1206,In_188,In_3335);
xor U1207 (N_1207,In_1455,In_4292);
and U1208 (N_1208,In_4166,In_2250);
nor U1209 (N_1209,In_4822,In_2106);
or U1210 (N_1210,In_4691,In_24);
nand U1211 (N_1211,In_4857,In_1121);
and U1212 (N_1212,In_912,In_2241);
or U1213 (N_1213,In_4994,In_2670);
nand U1214 (N_1214,In_2210,In_1593);
or U1215 (N_1215,In_1832,In_3412);
xnor U1216 (N_1216,In_1542,In_3450);
nand U1217 (N_1217,In_3431,In_4924);
nor U1218 (N_1218,In_4935,In_4090);
and U1219 (N_1219,In_3895,In_3646);
nand U1220 (N_1220,In_4069,In_4803);
nand U1221 (N_1221,In_3830,In_325);
or U1222 (N_1222,In_4655,In_2306);
and U1223 (N_1223,In_494,In_2588);
xor U1224 (N_1224,In_4960,In_2703);
nand U1225 (N_1225,In_2928,In_1771);
xor U1226 (N_1226,In_1913,In_727);
or U1227 (N_1227,In_2535,In_957);
nand U1228 (N_1228,In_2460,In_3440);
and U1229 (N_1229,In_77,In_2989);
nand U1230 (N_1230,In_4258,In_3386);
xor U1231 (N_1231,In_4711,In_3169);
or U1232 (N_1232,In_4679,In_3752);
nand U1233 (N_1233,In_1967,In_570);
and U1234 (N_1234,In_3394,In_19);
xor U1235 (N_1235,In_3131,In_1133);
nor U1236 (N_1236,In_1481,In_127);
nand U1237 (N_1237,In_4695,In_3844);
or U1238 (N_1238,In_3616,In_819);
and U1239 (N_1239,In_215,In_3369);
and U1240 (N_1240,In_4888,In_2315);
and U1241 (N_1241,In_1879,In_2637);
nand U1242 (N_1242,In_3404,In_2623);
nand U1243 (N_1243,In_4814,In_125);
and U1244 (N_1244,In_373,In_1360);
nand U1245 (N_1245,In_925,In_4820);
nor U1246 (N_1246,In_4494,In_2739);
xnor U1247 (N_1247,In_1483,In_1041);
nand U1248 (N_1248,In_1115,In_4176);
xor U1249 (N_1249,In_3908,In_1584);
nor U1250 (N_1250,In_1325,In_383);
and U1251 (N_1251,In_4388,In_3474);
nand U1252 (N_1252,In_3657,In_685);
xor U1253 (N_1253,In_297,In_4975);
nand U1254 (N_1254,In_1478,In_2598);
nor U1255 (N_1255,In_3354,In_4630);
or U1256 (N_1256,In_2842,In_744);
nor U1257 (N_1257,In_4473,In_3970);
or U1258 (N_1258,In_1071,In_3873);
and U1259 (N_1259,In_4203,In_1936);
xnor U1260 (N_1260,In_2383,In_3702);
nand U1261 (N_1261,In_4215,In_2334);
xor U1262 (N_1262,In_2897,In_1517);
and U1263 (N_1263,In_4074,In_1240);
or U1264 (N_1264,In_3182,In_2701);
xnor U1265 (N_1265,In_1557,In_1966);
nand U1266 (N_1266,In_2228,In_115);
xnor U1267 (N_1267,In_3619,In_761);
nand U1268 (N_1268,In_2169,In_375);
or U1269 (N_1269,In_3755,In_3005);
nand U1270 (N_1270,In_1154,In_2488);
xor U1271 (N_1271,In_2187,In_1343);
xnor U1272 (N_1272,In_4397,In_574);
nand U1273 (N_1273,In_991,In_845);
nand U1274 (N_1274,In_1105,In_3854);
nand U1275 (N_1275,In_4305,In_3557);
xor U1276 (N_1276,In_230,In_3446);
and U1277 (N_1277,In_4867,In_4289);
or U1278 (N_1278,In_599,In_1458);
or U1279 (N_1279,In_3933,In_3341);
nand U1280 (N_1280,In_4566,In_164);
nand U1281 (N_1281,In_3222,In_524);
nand U1282 (N_1282,In_281,In_3949);
nand U1283 (N_1283,In_505,In_4651);
nor U1284 (N_1284,In_4048,In_3311);
or U1285 (N_1285,In_750,In_3361);
nand U1286 (N_1286,In_4725,In_2741);
and U1287 (N_1287,In_92,In_1031);
xnor U1288 (N_1288,In_2358,In_2386);
nand U1289 (N_1289,In_4095,In_1119);
and U1290 (N_1290,In_2053,In_3243);
nand U1291 (N_1291,In_1404,In_1983);
or U1292 (N_1292,In_1472,In_2042);
nand U1293 (N_1293,In_4444,In_3428);
and U1294 (N_1294,In_3216,In_1605);
nor U1295 (N_1295,In_830,In_4523);
nor U1296 (N_1296,In_718,In_3018);
xnor U1297 (N_1297,In_149,In_580);
or U1298 (N_1298,In_563,In_4530);
or U1299 (N_1299,In_4622,In_3638);
or U1300 (N_1300,In_4441,In_3155);
xor U1301 (N_1301,In_2090,In_2185);
or U1302 (N_1302,In_1873,In_1634);
and U1303 (N_1303,In_2620,In_2229);
nand U1304 (N_1304,In_4325,In_1677);
xnor U1305 (N_1305,In_4267,In_3665);
nand U1306 (N_1306,In_4464,In_1678);
or U1307 (N_1307,In_1783,In_1471);
xor U1308 (N_1308,In_4369,In_3775);
nand U1309 (N_1309,In_1768,In_2913);
xnor U1310 (N_1310,In_3961,In_4595);
nand U1311 (N_1311,In_218,In_747);
nor U1312 (N_1312,In_3500,In_4895);
xnor U1313 (N_1313,In_321,In_1631);
nand U1314 (N_1314,In_4224,In_776);
nand U1315 (N_1315,In_1563,In_3476);
or U1316 (N_1316,In_657,In_2433);
nand U1317 (N_1317,In_4134,In_779);
or U1318 (N_1318,In_2693,In_3584);
and U1319 (N_1319,In_1941,In_1130);
xor U1320 (N_1320,In_2915,In_667);
nor U1321 (N_1321,In_1971,In_3861);
xnor U1322 (N_1322,In_2747,In_3781);
and U1323 (N_1323,In_1826,In_2803);
nor U1324 (N_1324,In_3077,In_432);
or U1325 (N_1325,In_166,In_4271);
and U1326 (N_1326,In_364,In_4366);
and U1327 (N_1327,In_4991,In_902);
nand U1328 (N_1328,In_3764,In_1829);
nand U1329 (N_1329,In_3990,In_4717);
or U1330 (N_1330,In_594,In_4116);
and U1331 (N_1331,In_1485,In_1859);
xnor U1332 (N_1332,In_2016,In_2575);
nor U1333 (N_1333,In_3408,In_323);
xnor U1334 (N_1334,In_4183,In_4731);
nor U1335 (N_1335,In_2580,In_3481);
nor U1336 (N_1336,In_2986,In_4861);
xnor U1337 (N_1337,In_4308,In_2127);
and U1338 (N_1338,In_1821,In_1286);
nand U1339 (N_1339,In_529,In_1152);
nor U1340 (N_1340,In_2512,In_938);
and U1341 (N_1341,In_1232,In_4874);
or U1342 (N_1342,In_1942,In_4687);
and U1343 (N_1343,In_1668,In_884);
and U1344 (N_1344,In_1876,In_2751);
xor U1345 (N_1345,In_104,In_1943);
or U1346 (N_1346,In_4958,In_2793);
nor U1347 (N_1347,In_337,In_313);
xnor U1348 (N_1348,In_1341,In_2834);
and U1349 (N_1349,In_924,In_628);
and U1350 (N_1350,In_3444,In_2969);
xor U1351 (N_1351,In_4424,In_3327);
nand U1352 (N_1352,In_1717,In_2032);
and U1353 (N_1353,In_1647,In_677);
nand U1354 (N_1354,In_3788,In_3241);
and U1355 (N_1355,In_4838,In_93);
xor U1356 (N_1356,In_770,In_4340);
xnor U1357 (N_1357,In_3337,In_555);
nor U1358 (N_1358,In_425,In_2087);
and U1359 (N_1359,In_4791,In_1047);
xor U1360 (N_1360,In_567,In_2962);
and U1361 (N_1361,In_440,In_3367);
nor U1362 (N_1362,In_4536,In_4298);
nor U1363 (N_1363,In_2776,In_4398);
xor U1364 (N_1364,In_1433,In_1085);
or U1365 (N_1365,In_4229,In_1157);
and U1366 (N_1366,In_4170,In_4051);
xnor U1367 (N_1367,In_3514,In_772);
and U1368 (N_1368,In_2034,In_1652);
xor U1369 (N_1369,In_351,In_2448);
nor U1370 (N_1370,In_1156,In_4144);
nor U1371 (N_1371,In_2944,In_1191);
nor U1372 (N_1372,In_1885,In_1301);
nand U1373 (N_1373,In_1896,In_3377);
nor U1374 (N_1374,In_1043,In_3555);
nand U1375 (N_1375,In_4010,In_1798);
or U1376 (N_1376,In_355,In_1650);
nor U1377 (N_1377,In_2871,In_4027);
nor U1378 (N_1378,In_3850,In_4438);
or U1379 (N_1379,In_2889,In_3911);
nor U1380 (N_1380,In_1494,In_2066);
or U1381 (N_1381,In_3796,In_3959);
and U1382 (N_1382,In_4114,In_2309);
xnor U1383 (N_1383,In_71,In_2321);
nand U1384 (N_1384,In_654,In_3160);
or U1385 (N_1385,In_3448,In_934);
and U1386 (N_1386,In_2761,In_950);
xnor U1387 (N_1387,In_4934,In_1195);
nor U1388 (N_1388,In_828,In_2005);
xnor U1389 (N_1389,In_826,In_1920);
nor U1390 (N_1390,In_1998,In_897);
nor U1391 (N_1391,In_2927,In_1991);
and U1392 (N_1392,In_2721,In_426);
xor U1393 (N_1393,In_87,In_3023);
nand U1394 (N_1394,In_4054,In_3069);
or U1395 (N_1395,In_3138,In_2865);
xor U1396 (N_1396,In_1764,In_3381);
or U1397 (N_1397,In_1779,In_20);
and U1398 (N_1398,In_3934,In_2099);
and U1399 (N_1399,In_2665,In_2590);
or U1400 (N_1400,In_4449,In_3596);
and U1401 (N_1401,In_2437,In_863);
or U1402 (N_1402,In_2579,In_506);
nand U1403 (N_1403,In_2013,In_3901);
nand U1404 (N_1404,In_4123,In_4870);
and U1405 (N_1405,In_3636,In_1623);
or U1406 (N_1406,In_1171,In_886);
and U1407 (N_1407,In_3599,In_3313);
nor U1408 (N_1408,In_2232,In_220);
xnor U1409 (N_1409,In_4194,In_3536);
or U1410 (N_1410,In_2500,In_626);
nor U1411 (N_1411,In_2484,In_1897);
or U1412 (N_1412,In_2692,In_2343);
and U1413 (N_1413,In_4359,In_1937);
and U1414 (N_1414,In_2445,In_140);
nand U1415 (N_1415,In_4637,In_4272);
or U1416 (N_1416,In_4980,In_1270);
or U1417 (N_1417,In_2984,In_3385);
nand U1418 (N_1418,In_4175,In_2163);
or U1419 (N_1419,In_2398,In_2328);
nor U1420 (N_1420,In_562,In_4016);
or U1421 (N_1421,In_1718,In_3278);
and U1422 (N_1422,In_260,In_1669);
nand U1423 (N_1423,In_2057,In_4859);
nand U1424 (N_1424,In_3219,In_3211);
xor U1425 (N_1425,In_409,In_4276);
and U1426 (N_1426,In_4373,In_3988);
nor U1427 (N_1427,In_3296,In_2939);
xnor U1428 (N_1428,In_2260,In_1173);
nor U1429 (N_1429,In_4535,In_4936);
xnor U1430 (N_1430,In_3996,In_2247);
nand U1431 (N_1431,In_2872,In_1603);
and U1432 (N_1432,In_1406,In_186);
and U1433 (N_1433,In_4561,In_2117);
and U1434 (N_1434,In_1774,In_1084);
and U1435 (N_1435,In_4672,In_4392);
nor U1436 (N_1436,In_4940,In_719);
xor U1437 (N_1437,In_1319,In_3696);
nand U1438 (N_1438,In_1480,In_4470);
nor U1439 (N_1439,In_1743,In_872);
nand U1440 (N_1440,In_302,In_2458);
xnor U1441 (N_1441,In_2234,In_2033);
nor U1442 (N_1442,In_801,In_2316);
xor U1443 (N_1443,In_3007,In_3725);
and U1444 (N_1444,In_2851,In_1732);
xor U1445 (N_1445,In_2631,In_2478);
nand U1446 (N_1446,In_2248,In_2630);
or U1447 (N_1447,In_1030,In_468);
and U1448 (N_1448,In_1068,In_3397);
or U1449 (N_1449,In_1235,In_812);
or U1450 (N_1450,In_1836,In_4415);
or U1451 (N_1451,In_1217,In_1179);
nor U1452 (N_1452,In_1661,In_4169);
nand U1453 (N_1453,In_1916,In_2813);
nor U1454 (N_1454,In_1522,In_162);
nor U1455 (N_1455,In_4154,In_2067);
or U1456 (N_1456,In_4177,In_2998);
or U1457 (N_1457,In_2829,In_3052);
and U1458 (N_1458,In_3174,In_4617);
or U1459 (N_1459,In_1018,In_3132);
nor U1460 (N_1460,In_2021,In_1963);
xor U1461 (N_1461,In_1761,In_2211);
nand U1462 (N_1462,In_3286,In_686);
nor U1463 (N_1463,In_4342,In_4394);
xnor U1464 (N_1464,In_1358,In_1917);
and U1465 (N_1465,In_1752,In_2625);
xnor U1466 (N_1466,In_3778,In_3396);
and U1467 (N_1467,In_1144,In_3698);
nor U1468 (N_1468,In_1816,In_3047);
nor U1469 (N_1469,In_4245,In_4737);
and U1470 (N_1470,In_4036,In_2578);
and U1471 (N_1471,In_1901,In_2356);
nand U1472 (N_1472,In_3275,In_1371);
nor U1473 (N_1473,In_3020,In_2035);
nand U1474 (N_1474,In_2396,In_4581);
nor U1475 (N_1475,In_3684,In_821);
xor U1476 (N_1476,In_2643,In_2651);
nand U1477 (N_1477,In_1766,In_400);
or U1478 (N_1478,In_63,In_4657);
xor U1479 (N_1479,In_4427,In_3971);
xnor U1480 (N_1480,In_4472,In_965);
nor U1481 (N_1481,In_2694,In_1786);
or U1482 (N_1482,In_4693,In_3669);
or U1483 (N_1483,In_926,In_4564);
or U1484 (N_1484,In_2482,In_2165);
xnor U1485 (N_1485,In_2873,In_139);
xnor U1486 (N_1486,In_3968,In_2368);
and U1487 (N_1487,In_2959,In_1226);
or U1488 (N_1488,In_3818,In_3919);
nor U1489 (N_1489,In_3728,In_867);
nor U1490 (N_1490,In_204,In_4993);
and U1491 (N_1491,In_4037,In_4358);
or U1492 (N_1492,In_2048,In_2401);
or U1493 (N_1493,In_1612,In_2345);
nor U1494 (N_1494,In_350,In_1660);
and U1495 (N_1495,In_2244,In_2563);
nor U1496 (N_1496,In_3101,In_2202);
nand U1497 (N_1497,In_537,In_4839);
xor U1498 (N_1498,In_794,In_4222);
nor U1499 (N_1499,In_2514,In_1935);
xnor U1500 (N_1500,In_1869,In_4120);
nor U1501 (N_1501,In_746,In_3203);
or U1502 (N_1502,In_4315,In_2391);
and U1503 (N_1503,In_2844,In_3148);
or U1504 (N_1504,In_3841,In_4389);
nand U1505 (N_1505,In_1237,In_4730);
xor U1506 (N_1506,In_731,In_1196);
nor U1507 (N_1507,In_2801,In_3012);
and U1508 (N_1508,In_564,In_1742);
nor U1509 (N_1509,In_1646,In_2963);
nor U1510 (N_1510,In_42,In_3264);
nand U1511 (N_1511,In_724,In_2904);
nor U1512 (N_1512,In_3701,In_1586);
and U1513 (N_1513,In_365,In_4796);
xnor U1514 (N_1514,In_4448,In_4736);
or U1515 (N_1515,In_1072,In_467);
xor U1516 (N_1516,In_2375,In_3401);
or U1517 (N_1517,In_3004,In_2645);
nor U1518 (N_1518,In_2025,In_4904);
or U1519 (N_1519,In_2162,In_2717);
nor U1520 (N_1520,In_3297,In_4493);
and U1521 (N_1521,In_736,In_1474);
and U1522 (N_1522,In_308,In_831);
and U1523 (N_1523,In_586,In_882);
nand U1524 (N_1524,In_3926,In_999);
nor U1525 (N_1525,In_138,In_2754);
nand U1526 (N_1526,In_1150,In_4101);
nor U1527 (N_1527,In_1847,In_491);
xnor U1528 (N_1528,In_165,In_2496);
or U1529 (N_1529,In_310,In_3753);
nand U1530 (N_1530,In_3231,In_3273);
nand U1531 (N_1531,In_1027,In_518);
nand U1532 (N_1532,In_3902,In_986);
and U1533 (N_1533,In_1394,In_1255);
nor U1534 (N_1534,In_4378,In_1748);
nand U1535 (N_1535,In_3667,In_3049);
or U1536 (N_1536,In_2092,In_1381);
or U1537 (N_1537,In_3715,In_3280);
nor U1538 (N_1538,In_4823,In_3071);
nor U1539 (N_1539,In_4585,In_3251);
and U1540 (N_1540,In_3733,In_4942);
xnor U1541 (N_1541,In_892,In_322);
or U1542 (N_1542,In_2510,In_1438);
xnor U1543 (N_1543,In_623,In_4908);
xnor U1544 (N_1544,In_3120,In_1780);
nor U1545 (N_1545,In_3400,In_4273);
nor U1546 (N_1546,In_141,In_1723);
xor U1547 (N_1547,In_3957,In_921);
or U1548 (N_1548,In_1886,In_552);
nand U1549 (N_1549,In_2954,In_18);
and U1550 (N_1550,In_4150,In_4914);
nor U1551 (N_1551,In_1249,In_1484);
nand U1552 (N_1552,In_2893,In_3531);
or U1553 (N_1553,In_2426,In_4327);
and U1554 (N_1554,In_2143,In_3319);
and U1555 (N_1555,In_2735,In_4083);
and U1556 (N_1556,In_4216,In_3035);
nand U1557 (N_1557,In_3685,In_4262);
nand U1558 (N_1558,In_1479,In_4931);
xnor U1559 (N_1559,In_106,In_1176);
xor U1560 (N_1560,In_255,In_1411);
nor U1561 (N_1561,In_4417,In_4360);
nor U1562 (N_1562,In_2675,In_7);
or U1563 (N_1563,In_2838,In_3040);
and U1564 (N_1564,In_3624,In_981);
nand U1565 (N_1565,In_2798,In_932);
nor U1566 (N_1566,In_2756,In_83);
or U1567 (N_1567,In_3853,In_1091);
nand U1568 (N_1568,In_2766,In_4344);
or U1569 (N_1569,In_1708,In_522);
xor U1570 (N_1570,In_450,In_2412);
nor U1571 (N_1571,In_4623,In_3284);
or U1572 (N_1572,In_3106,In_3742);
and U1573 (N_1573,In_2468,In_3668);
or U1574 (N_1574,In_3661,In_59);
or U1575 (N_1575,In_1020,In_3252);
nor U1576 (N_1576,In_1444,In_107);
xnor U1577 (N_1577,In_1348,In_4923);
and U1578 (N_1578,In_1877,In_3422);
nand U1579 (N_1579,In_4214,In_4636);
nand U1580 (N_1580,In_4067,In_1560);
nand U1581 (N_1581,In_4307,In_1386);
nand U1582 (N_1582,In_1139,In_1544);
and U1583 (N_1583,In_79,In_1546);
and U1584 (N_1584,In_4751,In_922);
nor U1585 (N_1585,In_1328,In_233);
and U1586 (N_1586,In_927,In_4609);
nand U1587 (N_1587,In_25,In_2207);
and U1588 (N_1588,In_4707,In_4781);
nand U1589 (N_1589,In_972,In_2691);
or U1590 (N_1590,In_651,In_453);
or U1591 (N_1591,In_1288,In_2738);
or U1592 (N_1592,In_854,In_891);
or U1593 (N_1593,In_2780,In_3380);
and U1594 (N_1594,In_1023,In_2729);
nor U1595 (N_1595,In_639,In_271);
and U1596 (N_1596,In_4131,In_4602);
and U1597 (N_1597,In_4299,In_2246);
nor U1598 (N_1598,In_1537,In_2805);
nand U1599 (N_1599,In_4892,In_4584);
nor U1600 (N_1600,In_1701,In_4281);
or U1601 (N_1601,In_1610,In_306);
xor U1602 (N_1602,In_3295,In_4056);
nand U1603 (N_1603,In_2158,In_3944);
or U1604 (N_1604,In_2423,In_3776);
or U1605 (N_1605,In_2397,In_1168);
and U1606 (N_1606,In_616,In_3484);
nand U1607 (N_1607,In_288,In_4794);
nand U1608 (N_1608,In_544,In_2839);
or U1609 (N_1609,In_4669,In_1947);
and U1610 (N_1610,In_1574,In_652);
nand U1611 (N_1611,In_2434,In_3713);
nand U1612 (N_1612,In_2661,In_184);
nor U1613 (N_1613,In_4674,In_559);
xor U1614 (N_1614,In_967,In_1513);
nor U1615 (N_1615,In_3734,In_2288);
xnor U1616 (N_1616,In_2344,In_1006);
or U1617 (N_1617,In_231,In_3647);
nand U1618 (N_1618,In_3392,In_1802);
and U1619 (N_1619,In_1844,In_627);
or U1620 (N_1620,In_3478,In_1562);
nor U1621 (N_1621,In_1448,In_4714);
nor U1622 (N_1622,In_3287,In_720);
or U1623 (N_1623,In_2387,In_4982);
or U1624 (N_1624,In_1396,In_1182);
nor U1625 (N_1625,In_824,In_4664);
xor U1626 (N_1626,In_4206,In_2856);
nor U1627 (N_1627,In_3848,In_2708);
nor U1628 (N_1628,In_2914,In_3072);
nor U1629 (N_1629,In_2662,In_595);
and U1630 (N_1630,In_2419,In_4209);
nand U1631 (N_1631,In_4152,In_445);
and U1632 (N_1632,In_1427,In_4488);
or U1633 (N_1633,In_857,In_2037);
nor U1634 (N_1634,In_3124,In_855);
nor U1635 (N_1635,In_1193,In_4749);
or U1636 (N_1636,In_887,In_2634);
nor U1637 (N_1637,In_2338,In_2385);
nand U1638 (N_1638,In_3803,In_1813);
or U1639 (N_1639,In_3460,In_4499);
and U1640 (N_1640,In_56,In_179);
nor U1641 (N_1641,In_3184,In_343);
nand U1642 (N_1642,In_2600,In_1384);
nand U1643 (N_1643,In_3389,In_1884);
xor U1644 (N_1644,In_3480,In_1059);
nor U1645 (N_1645,In_2028,In_354);
or U1646 (N_1646,In_3975,In_4161);
xnor U1647 (N_1647,In_2292,In_2709);
nor U1648 (N_1648,In_1188,In_4312);
xor U1649 (N_1649,In_4925,In_4974);
xor U1650 (N_1650,In_1497,In_2038);
and U1651 (N_1651,In_969,In_4343);
or U1652 (N_1652,In_4185,In_3388);
nand U1653 (N_1653,In_557,In_2209);
nor U1654 (N_1654,In_610,In_743);
nand U1655 (N_1655,In_3582,In_3358);
nor U1656 (N_1656,In_1551,In_2043);
nor U1657 (N_1657,In_3714,In_4334);
xnor U1658 (N_1658,In_4779,In_565);
xnor U1659 (N_1659,In_1501,In_2802);
and U1660 (N_1660,In_753,In_4277);
xor U1661 (N_1661,In_1722,In_4759);
or U1662 (N_1662,In_4539,In_598);
nand U1663 (N_1663,In_253,In_4698);
nor U1664 (N_1664,In_4518,In_4885);
nor U1665 (N_1665,In_1804,In_1486);
or U1666 (N_1666,In_96,In_3983);
and U1667 (N_1667,In_2683,In_3656);
or U1668 (N_1668,In_2378,In_2748);
and U1669 (N_1669,In_4921,In_2718);
nand U1670 (N_1670,In_1580,In_4675);
or U1671 (N_1671,In_4507,In_4682);
nand U1672 (N_1672,In_131,In_663);
and U1673 (N_1673,In_3836,In_1081);
nor U1674 (N_1674,In_4061,In_1986);
xnor U1675 (N_1675,In_3259,In_3763);
and U1676 (N_1676,In_2495,In_1857);
nor U1677 (N_1677,In_2332,In_454);
or U1678 (N_1678,In_3122,In_4884);
xor U1679 (N_1679,In_1762,In_4332);
nor U1680 (N_1680,In_168,In_2436);
or U1681 (N_1681,In_3692,In_2947);
xor U1682 (N_1682,In_4044,In_4058);
and U1683 (N_1683,In_4553,In_4190);
and U1684 (N_1684,In_3790,In_4280);
or U1685 (N_1685,In_4349,In_3290);
xor U1686 (N_1686,In_3030,In_4160);
nor U1687 (N_1687,In_2156,In_117);
and U1688 (N_1688,In_3267,In_1287);
and U1689 (N_1689,In_2340,In_4850);
xor U1690 (N_1690,In_2531,In_3824);
nor U1691 (N_1691,In_39,In_1420);
nor U1692 (N_1692,In_1450,In_3218);
and U1693 (N_1693,In_1241,In_1127);
nor U1694 (N_1694,In_3044,In_702);
nor U1695 (N_1695,In_4597,In_954);
xor U1696 (N_1696,In_3449,In_2276);
or U1697 (N_1697,In_1970,In_1506);
nor U1698 (N_1698,In_1819,In_681);
or U1699 (N_1699,In_3411,In_2518);
nand U1700 (N_1700,In_575,In_1738);
xnor U1701 (N_1701,In_2152,In_1447);
or U1702 (N_1702,In_4078,In_3930);
nand U1703 (N_1703,In_1508,In_4129);
nand U1704 (N_1704,In_4849,In_209);
and U1705 (N_1705,In_2898,In_1379);
and U1706 (N_1706,In_4750,In_2098);
and U1707 (N_1707,In_1840,In_3941);
nand U1708 (N_1708,In_385,In_4955);
nand U1709 (N_1709,In_1345,In_3009);
and U1710 (N_1710,In_3587,In_3179);
or U1711 (N_1711,In_2220,In_4052);
xor U1712 (N_1712,In_4353,In_2551);
or U1713 (N_1713,In_566,In_1756);
nor U1714 (N_1714,In_1682,In_556);
xor U1715 (N_1715,In_2051,In_2270);
nor U1716 (N_1716,In_1434,In_735);
nand U1717 (N_1717,In_2476,In_2868);
xnor U1718 (N_1718,In_4828,In_1590);
or U1719 (N_1719,In_1655,In_4938);
or U1720 (N_1720,In_4555,In_3777);
nor U1721 (N_1721,In_3586,In_3189);
nand U1722 (N_1722,In_332,In_684);
nand U1723 (N_1723,In_2240,In_2977);
or U1724 (N_1724,In_4526,In_172);
nand U1725 (N_1725,In_3598,In_4489);
and U1726 (N_1726,In_2975,In_962);
nand U1727 (N_1727,In_3451,In_4077);
nor U1728 (N_1728,In_1245,In_47);
xor U1729 (N_1729,In_1904,In_1726);
xnor U1730 (N_1730,In_3395,In_2819);
nand U1731 (N_1731,In_4039,In_2206);
nor U1732 (N_1732,In_1616,In_4909);
or U1733 (N_1733,In_2102,In_4023);
or U1734 (N_1734,In_2608,In_2453);
xnor U1735 (N_1735,In_3338,In_3340);
xnor U1736 (N_1736,In_4542,In_2451);
nand U1737 (N_1737,In_4226,In_640);
xor U1738 (N_1738,In_4355,In_2745);
nor U1739 (N_1739,In_3036,In_2300);
nand U1740 (N_1740,In_2556,In_3720);
or U1741 (N_1741,In_4898,In_65);
nand U1742 (N_1742,In_4146,In_2133);
nand U1743 (N_1743,In_3549,In_1453);
nor U1744 (N_1744,In_646,In_955);
nor U1745 (N_1745,In_1960,In_678);
xor U1746 (N_1746,In_2129,In_2441);
and U1747 (N_1747,In_1306,In_1094);
xnor U1748 (N_1748,In_3858,In_4772);
xnor U1749 (N_1749,In_4862,In_1221);
nand U1750 (N_1750,In_4881,In_1488);
and U1751 (N_1751,In_3885,In_3585);
and U1752 (N_1752,In_121,In_2041);
and U1753 (N_1753,In_2365,In_3951);
xnor U1754 (N_1754,In_275,In_802);
xor U1755 (N_1755,In_3149,In_3600);
nand U1756 (N_1756,In_2667,In_1275);
xor U1757 (N_1757,In_754,In_27);
or U1758 (N_1758,In_3229,In_3840);
or U1759 (N_1759,In_749,In_4365);
nor U1760 (N_1760,In_585,In_648);
nor U1761 (N_1761,In_1051,In_3082);
nor U1762 (N_1762,In_1216,In_4211);
and U1763 (N_1763,In_3541,In_2924);
nand U1764 (N_1764,In_3640,In_2027);
or U1765 (N_1765,In_4644,In_3945);
or U1766 (N_1766,In_4465,In_2108);
or U1767 (N_1767,In_2319,In_2007);
nand U1768 (N_1768,In_236,In_2236);
nor U1769 (N_1769,In_1253,In_1153);
and U1770 (N_1770,In_3722,In_4878);
xnor U1771 (N_1771,In_3761,In_4328);
or U1772 (N_1772,In_242,In_2525);
xnor U1773 (N_1773,In_3145,In_3078);
and U1774 (N_1774,In_2948,In_3432);
and U1775 (N_1775,In_2384,In_2852);
and U1776 (N_1776,In_1549,In_1294);
nor U1777 (N_1777,In_2318,In_4324);
nand U1778 (N_1778,In_208,In_1918);
nand U1779 (N_1779,In_2290,In_2895);
nor U1780 (N_1780,In_3859,In_2124);
and U1781 (N_1781,In_4265,In_4816);
nor U1782 (N_1782,In_2749,In_2078);
nand U1783 (N_1783,In_2881,In_2577);
xor U1784 (N_1784,In_2646,In_2855);
nand U1785 (N_1785,In_3490,In_763);
nand U1786 (N_1786,In_3838,In_2654);
xor U1787 (N_1787,In_4181,In_4983);
nor U1788 (N_1788,In_4288,In_1911);
xnor U1789 (N_1789,In_4011,In_2660);
xor U1790 (N_1790,In_4207,In_4082);
and U1791 (N_1791,In_3981,In_4471);
and U1792 (N_1792,In_1005,In_1925);
nor U1793 (N_1793,In_2014,In_3236);
xnor U1794 (N_1794,In_3333,In_1820);
xnor U1795 (N_1795,In_3161,In_1443);
xnor U1796 (N_1796,In_836,In_3954);
or U1797 (N_1797,In_1588,In_4642);
nor U1798 (N_1798,In_2558,In_3456);
and U1799 (N_1799,In_1535,In_590);
nor U1800 (N_1800,In_344,In_3472);
and U1801 (N_1801,In_1865,In_721);
nand U1802 (N_1802,In_4661,In_2886);
nor U1803 (N_1803,In_4956,In_1095);
xor U1804 (N_1804,In_953,In_341);
and U1805 (N_1805,In_4613,In_3108);
nor U1806 (N_1806,In_3750,In_1604);
xor U1807 (N_1807,In_1996,In_3434);
nor U1808 (N_1808,In_3162,In_57);
or U1809 (N_1809,In_798,In_4875);
and U1810 (N_1810,In_3503,In_2190);
nor U1811 (N_1811,In_4139,In_1626);
nand U1812 (N_1812,In_2373,In_4451);
xnor U1813 (N_1813,In_146,In_2712);
xor U1814 (N_1814,In_3208,In_895);
nand U1815 (N_1815,In_600,In_1082);
nor U1816 (N_1816,In_2268,In_4205);
nor U1817 (N_1817,In_4104,In_4232);
xnor U1818 (N_1818,In_2487,In_2861);
nand U1819 (N_1819,In_4927,In_2186);
or U1820 (N_1820,In_4562,In_1842);
nand U1821 (N_1821,In_3518,In_2993);
and U1822 (N_1822,In_3626,In_4986);
or U1823 (N_1823,In_174,In_769);
xnor U1824 (N_1824,In_670,In_3238);
nand U1825 (N_1825,In_2529,In_2196);
xor U1826 (N_1826,In_2656,In_2624);
nand U1827 (N_1827,In_258,In_2088);
or U1828 (N_1828,In_3704,In_3697);
xnor U1829 (N_1829,In_4810,In_2073);
xor U1830 (N_1830,In_4745,In_3135);
nand U1831 (N_1831,In_4587,In_3620);
and U1832 (N_1832,In_3083,In_4068);
nor U1833 (N_1833,In_99,In_4650);
or U1834 (N_1834,In_3164,In_1837);
and U1835 (N_1835,In_2130,In_1322);
nand U1836 (N_1836,In_730,In_1806);
nand U1837 (N_1837,In_1881,In_2594);
nand U1838 (N_1838,In_4167,In_2082);
nor U1839 (N_1839,In_3312,In_2218);
and U1840 (N_1840,In_4604,In_3562);
or U1841 (N_1841,In_2148,In_1181);
nand U1842 (N_1842,In_3511,In_3749);
nand U1843 (N_1843,In_3948,In_4633);
and U1844 (N_1844,In_548,In_4804);
xnor U1845 (N_1845,In_945,In_4668);
nor U1846 (N_1846,In_3732,In_3393);
and U1847 (N_1847,In_3309,In_4513);
xor U1848 (N_1848,In_1366,In_3843);
or U1849 (N_1849,In_2443,In_2097);
and U1850 (N_1850,In_2596,In_713);
nand U1851 (N_1851,In_1979,In_1110);
xnor U1852 (N_1852,In_4766,In_2920);
and U1853 (N_1853,In_848,In_1490);
and U1854 (N_1854,In_2789,In_2961);
or U1855 (N_1855,In_1713,In_4971);
and U1856 (N_1856,In_112,In_877);
or U1857 (N_1857,In_516,In_2591);
and U1858 (N_1858,In_1266,In_3540);
or U1859 (N_1859,In_4199,In_3136);
xnor U1860 (N_1860,In_1749,In_4136);
nand U1861 (N_1861,In_1422,In_5);
or U1862 (N_1862,In_2277,In_4833);
xnor U1863 (N_1863,In_4076,In_3353);
and U1864 (N_1864,In_1587,In_3563);
xor U1865 (N_1865,In_2049,In_885);
and U1866 (N_1866,In_940,In_282);
nor U1867 (N_1867,In_1281,In_2483);
and U1868 (N_1868,In_3523,In_4538);
xnor U1869 (N_1869,In_4302,In_2616);
or U1870 (N_1870,In_3244,In_4719);
and U1871 (N_1871,In_135,In_4756);
nand U1872 (N_1872,In_2427,In_1594);
xnor U1873 (N_1873,In_2627,In_2804);
and U1874 (N_1874,In_3202,In_1956);
or U1875 (N_1875,In_2263,In_3606);
nor U1876 (N_1876,In_861,In_3653);
or U1877 (N_1877,In_2430,In_1902);
or U1878 (N_1878,In_102,In_2849);
nor U1879 (N_1879,In_3240,In_989);
and U1880 (N_1880,In_740,In_4826);
nand U1881 (N_1881,In_3857,In_58);
nand U1882 (N_1882,In_4221,In_2275);
or U1883 (N_1883,In_2682,In_2238);
nand U1884 (N_1884,In_1809,In_2030);
and U1885 (N_1885,In_2182,In_436);
xnor U1886 (N_1886,In_4456,In_4919);
nand U1887 (N_1887,In_1120,In_843);
nor U1888 (N_1888,In_4692,In_4592);
nand U1889 (N_1889,In_532,In_541);
nor U1890 (N_1890,In_4963,In_379);
nand U1891 (N_1891,In_2069,In_387);
or U1892 (N_1892,In_4043,In_4624);
xor U1893 (N_1893,In_2192,In_4228);
and U1894 (N_1894,In_3051,In_1415);
nor U1895 (N_1895,In_2175,In_1952);
nand U1896 (N_1896,In_3477,In_2205);
or U1897 (N_1897,In_3382,In_1470);
or U1898 (N_1898,In_1727,In_2409);
xnor U1899 (N_1899,In_1736,In_2134);
nand U1900 (N_1900,In_1959,In_2602);
or U1901 (N_1901,In_4829,In_3539);
nand U1902 (N_1902,In_1468,In_1258);
xor U1903 (N_1903,In_1812,In_3141);
xor U1904 (N_1904,In_296,In_849);
xor U1905 (N_1905,In_2790,In_4233);
xor U1906 (N_1906,In_4625,In_1912);
or U1907 (N_1907,In_1356,In_3142);
or U1908 (N_1908,In_3073,In_1931);
nand U1909 (N_1909,In_191,In_3583);
nor U1910 (N_1910,In_4671,In_2787);
nor U1911 (N_1911,In_2763,In_4086);
xor U1912 (N_1912,In_2669,In_4256);
nor U1913 (N_1913,In_4948,In_1380);
nand U1914 (N_1914,In_4106,In_2707);
nand U1915 (N_1915,In_4504,In_2814);
and U1916 (N_1916,In_2047,In_185);
nor U1917 (N_1917,In_1202,In_2056);
nand U1918 (N_1918,In_2414,In_1321);
nand U1919 (N_1919,In_2690,In_3913);
and U1920 (N_1920,In_2971,In_3757);
nand U1921 (N_1921,In_4778,In_1015);
nor U1922 (N_1922,In_4093,In_1663);
or U1923 (N_1923,In_217,In_469);
nor U1924 (N_1924,In_2534,In_4534);
nand U1925 (N_1925,In_1350,In_2424);
and U1926 (N_1926,In_1719,In_2216);
and U1927 (N_1927,In_2633,In_3678);
or U1928 (N_1928,In_3263,In_4266);
nor U1929 (N_1929,In_1674,In_73);
and U1930 (N_1930,In_3299,In_1556);
nor U1931 (N_1931,In_1293,In_1848);
nand U1932 (N_1932,In_2278,In_80);
nor U1933 (N_1933,In_904,In_2681);
nand U1934 (N_1934,In_3024,In_4906);
or U1935 (N_1935,In_4306,In_4138);
or U1936 (N_1936,In_4780,In_4709);
or U1937 (N_1937,In_2307,In_2929);
nand U1938 (N_1938,In_1824,In_163);
nand U1939 (N_1939,In_2812,In_1333);
nor U1940 (N_1940,In_4484,In_4295);
xnor U1941 (N_1941,In_2045,In_3194);
nand U1942 (N_1942,In_4351,In_1227);
nand U1943 (N_1943,In_301,In_1940);
nand U1944 (N_1944,In_3239,In_3027);
nor U1945 (N_1945,In_1302,In_2212);
or U1946 (N_1946,In_2457,In_340);
xnor U1947 (N_1947,In_507,In_2200);
and U1948 (N_1948,In_1353,In_1011);
nor U1949 (N_1949,In_1292,In_3517);
or U1950 (N_1950,In_2119,In_3965);
or U1951 (N_1951,In_509,In_4382);
xor U1952 (N_1952,In_4543,In_2310);
nand U1953 (N_1953,In_1864,In_3249);
and U1954 (N_1954,In_3111,In_1198);
and U1955 (N_1955,In_46,In_3473);
and U1956 (N_1956,In_2351,In_2036);
nor U1957 (N_1957,In_3529,In_414);
or U1958 (N_1958,In_3464,In_4522);
nor U1959 (N_1959,In_60,In_4656);
nor U1960 (N_1960,In_4492,In_2539);
or U1961 (N_1961,In_650,In_2298);
and U1962 (N_1962,In_3804,In_3566);
or U1963 (N_1963,In_4860,In_374);
or U1964 (N_1964,In_2120,In_3037);
and U1965 (N_1965,In_2779,In_3499);
and U1966 (N_1966,In_2447,In_4391);
nand U1967 (N_1967,In_4696,In_4062);
and U1968 (N_1968,In_1973,In_900);
xnor U1969 (N_1969,In_2840,In_2293);
and U1970 (N_1970,In_3625,In_2997);
or U1971 (N_1971,In_809,In_3344);
nand U1972 (N_1972,In_2080,In_919);
nand U1973 (N_1973,In_3545,In_4568);
and U1974 (N_1974,In_1169,In_4573);
nand U1975 (N_1975,In_3622,In_84);
nor U1976 (N_1976,In_1180,In_245);
and U1977 (N_1977,In_3168,In_1989);
and U1978 (N_1978,In_4854,In_4744);
and U1979 (N_1979,In_1926,In_2303);
and U1980 (N_1980,In_2888,In_4225);
xnor U1981 (N_1981,In_2064,In_3305);
and U1982 (N_1982,In_1539,In_3682);
and U1983 (N_1983,In_4853,In_710);
or U1984 (N_1984,In_2432,In_3508);
and U1985 (N_1985,In_224,In_4578);
nand U1986 (N_1986,In_239,In_2123);
nand U1987 (N_1987,In_3812,In_3987);
or U1988 (N_1988,In_3633,In_3374);
or U1989 (N_1989,In_212,In_2357);
nand U1990 (N_1990,In_4282,In_1456);
nand U1991 (N_1991,In_2926,In_1799);
and U1992 (N_1992,In_2957,In_593);
and U1993 (N_1993,In_4482,In_4723);
or U1994 (N_1994,In_1814,In_2668);
or U1995 (N_1995,In_793,In_621);
and U1996 (N_1996,In_1079,In_1552);
nor U1997 (N_1997,In_3237,In_2217);
nor U1998 (N_1998,In_3253,In_2105);
nor U1999 (N_1999,In_3067,In_2503);
xor U2000 (N_2000,N_565,In_3257);
nor U2001 (N_2001,N_693,In_2817);
xor U2002 (N_2002,N_1767,In_4072);
nand U2003 (N_2003,N_399,N_29);
xnor U2004 (N_2004,N_130,In_4886);
and U2005 (N_2005,N_1013,N_36);
and U2006 (N_2006,N_1176,N_615);
and U2007 (N_2007,In_397,N_1991);
nand U2008 (N_2008,N_449,In_69);
xnor U2009 (N_2009,In_846,N_1916);
nor U2010 (N_2010,N_1247,N_1713);
nor U2011 (N_2011,N_1367,N_1688);
or U2012 (N_2012,N_1964,N_1698);
xnor U2013 (N_2013,In_3261,In_3847);
nand U2014 (N_2014,N_730,N_1124);
nor U2015 (N_2015,N_1224,In_3195);
nor U2016 (N_2016,N_1941,In_4119);
xor U2017 (N_2017,In_874,N_393);
and U2018 (N_2018,In_2884,In_4204);
nor U2019 (N_2019,In_1696,In_2125);
xnor U2020 (N_2020,N_310,In_1409);
and U2021 (N_2021,N_109,In_4667);
and U2022 (N_2022,N_1527,In_3321);
nor U2023 (N_2023,N_616,In_4476);
xnor U2024 (N_2024,N_311,In_992);
xnor U2025 (N_2025,N_715,In_3899);
nor U2026 (N_2026,N_1596,N_1403);
xnor U2027 (N_2027,In_1137,In_392);
and U2028 (N_2028,In_291,N_1297);
and U2029 (N_2029,N_544,N_423);
xnor U2030 (N_2030,N_1405,N_1167);
and U2031 (N_2031,N_738,In_358);
or U2032 (N_2032,N_573,N_1834);
and U2033 (N_2033,N_1590,N_1120);
xnor U2034 (N_2034,N_1915,N_721);
and U2035 (N_2035,N_1877,In_416);
and U2036 (N_2036,N_1707,N_280);
and U2037 (N_2037,In_2279,In_1004);
nor U2038 (N_2038,N_1463,N_245);
and U2039 (N_2039,N_614,N_270);
and U2040 (N_2040,N_30,N_1032);
nand U2041 (N_2041,N_1576,N_605);
and U2042 (N_2042,N_1676,N_1191);
and U2043 (N_2043,N_479,N_1036);
xor U2044 (N_2044,In_192,N_1432);
nand U2045 (N_2045,N_725,N_476);
and U2046 (N_2046,N_1634,N_118);
and U2047 (N_2047,N_1479,N_1739);
nor U2048 (N_2048,In_659,In_4363);
and U2049 (N_2049,In_2289,N_1101);
nor U2050 (N_2050,N_1069,N_666);
nand U2051 (N_2051,In_3597,N_390);
or U2052 (N_2052,N_463,N_980);
xor U2053 (N_2053,N_765,N_690);
and U2054 (N_2054,N_1773,In_2213);
xor U2055 (N_2055,In_543,N_697);
xnor U2056 (N_2056,N_1113,In_1296);
or U2057 (N_2057,In_1676,N_1374);
nand U2058 (N_2058,N_665,In_3693);
nor U2059 (N_2059,In_347,In_1835);
nor U2060 (N_2060,In_3368,N_1090);
xor U2061 (N_2061,N_890,In_201);
xor U2062 (N_2062,In_1398,N_1960);
nand U2063 (N_2063,In_4261,N_1437);
or U2064 (N_2064,N_481,In_2347);
nand U2065 (N_2065,N_1709,N_1165);
and U2066 (N_2066,N_1125,In_4844);
or U2067 (N_2067,N_967,In_540);
nand U2068 (N_2068,N_1440,N_453);
xor U2069 (N_2069,N_1265,N_985);
nor U2070 (N_2070,N_660,In_390);
nor U2071 (N_2071,N_1984,In_2170);
nor U2072 (N_2072,N_1901,N_1768);
nand U2073 (N_2073,N_1725,In_783);
nor U2074 (N_2074,N_862,N_363);
and U2075 (N_2075,N_1734,In_272);
and U2076 (N_2076,N_952,N_1205);
xnor U2077 (N_2077,In_1908,N_120);
xnor U2078 (N_2078,N_112,In_3868);
nor U2079 (N_2079,In_3314,In_243);
nor U2080 (N_2080,In_915,N_684);
nor U2081 (N_2081,In_1815,N_1539);
and U2082 (N_2082,N_255,In_3272);
and U2083 (N_2083,In_4586,N_912);
or U2084 (N_2084,N_1956,N_526);
or U2085 (N_2085,N_1343,In_4352);
xor U2086 (N_2086,N_1587,In_1831);
nor U2087 (N_2087,N_809,N_101);
and U2088 (N_2088,N_55,In_412);
nor U2089 (N_2089,N_142,N_602);
nand U2090 (N_2090,In_4713,In_4998);
and U2091 (N_2091,N_1782,In_2208);
nor U2092 (N_2092,N_1801,N_762);
and U2093 (N_2093,In_1716,In_2297);
nor U2094 (N_2094,N_1225,N_1067);
xor U2095 (N_2095,N_1600,N_838);
nand U2096 (N_2096,N_1800,N_1366);
nand U2097 (N_2097,In_2910,N_1959);
nand U2098 (N_2098,N_1663,N_1997);
nand U2099 (N_2099,N_842,In_36);
xor U2100 (N_2100,N_777,N_205);
nor U2101 (N_2101,In_4703,In_1617);
nor U2102 (N_2102,In_3070,In_3966);
xnor U2103 (N_2103,In_496,N_1859);
xor U2104 (N_2104,In_3062,N_571);
nand U2105 (N_2105,N_870,N_1728);
nand U2106 (N_2106,N_1717,In_3723);
nand U2107 (N_2107,In_4118,N_563);
and U2108 (N_2108,N_400,In_3534);
or U2109 (N_2109,N_591,N_577);
nand U2110 (N_2110,In_1044,N_16);
xnor U2111 (N_2111,In_2863,N_1481);
and U2112 (N_2112,In_1711,N_408);
nor U2113 (N_2113,In_816,In_1274);
and U2114 (N_2114,N_1502,In_1757);
xor U2115 (N_2115,In_2022,In_2390);
or U2116 (N_2116,In_1950,N_859);
nand U2117 (N_2117,N_794,In_1332);
nor U2118 (N_2118,N_982,N_1529);
and U2119 (N_2119,In_3849,N_1427);
nor U2120 (N_2120,N_1078,In_4321);
nor U2121 (N_2121,N_394,N_358);
or U2122 (N_2122,N_1239,N_1687);
and U2123 (N_2123,In_3347,N_185);
nor U2124 (N_2124,In_3098,N_1862);
nand U2125 (N_2125,N_1434,N_268);
or U2126 (N_2126,N_1455,N_1616);
nor U2127 (N_2127,N_1757,N_1885);
nand U2128 (N_2128,N_317,In_1141);
or U2129 (N_2129,In_2902,In_521);
nand U2130 (N_2130,N_1344,In_4688);
nor U2131 (N_2131,In_1944,N_1809);
or U2132 (N_2132,In_3048,N_1290);
and U2133 (N_2133,N_798,N_628);
nor U2134 (N_2134,N_552,N_1549);
xnor U2135 (N_2135,N_286,N_769);
xor U2136 (N_2136,In_2744,In_791);
nor U2137 (N_2137,N_195,N_953);
nand U2138 (N_2138,N_1094,In_2996);
nor U2139 (N_2139,In_739,N_718);
and U2140 (N_2140,N_915,N_1003);
nand U2141 (N_2141,N_1945,N_1640);
or U2142 (N_2142,In_1622,N_578);
nand U2143 (N_2143,N_419,N_1417);
or U2144 (N_2144,N_241,N_1790);
xnor U2145 (N_2145,In_4379,N_81);
nand U2146 (N_2146,In_1189,In_2722);
xnor U2147 (N_2147,N_1515,N_1064);
or U2148 (N_2148,In_3317,In_994);
and U2149 (N_2149,In_1978,N_1321);
and U2150 (N_2150,N_1411,N_780);
and U2151 (N_2151,N_1714,N_1431);
nand U2152 (N_2152,In_3876,N_1339);
nor U2153 (N_2153,N_1678,N_389);
nand U2154 (N_2154,N_743,In_167);
nand U2155 (N_2155,N_1471,N_719);
and U2156 (N_2156,N_1001,N_349);
and U2157 (N_2157,In_993,N_708);
nor U2158 (N_2158,N_1871,N_728);
xor U2159 (N_2159,N_1820,In_1493);
and U2160 (N_2160,N_787,N_168);
and U2161 (N_2161,N_844,N_1169);
nand U2162 (N_2162,In_2553,In_2075);
xor U2163 (N_2163,N_1690,N_231);
nand U2164 (N_2164,In_1278,N_958);
nand U2165 (N_2165,N_1751,N_652);
xnor U2166 (N_2166,N_1581,N_1115);
nor U2167 (N_2167,N_222,N_1319);
or U2168 (N_2168,N_314,N_627);
nor U2169 (N_2169,N_1720,In_430);
nand U2170 (N_2170,N_1159,N_478);
nand U2171 (N_2171,In_4411,In_2994);
and U2172 (N_2172,N_1781,N_1618);
nand U2173 (N_2173,N_990,N_546);
xnor U2174 (N_2174,N_681,N_116);
xor U2175 (N_2175,In_2727,N_82);
or U2176 (N_2176,N_397,In_2752);
nor U2177 (N_2177,N_486,N_1489);
and U2178 (N_2178,In_1554,N_1804);
nand U2179 (N_2179,In_2649,N_1095);
xor U2180 (N_2180,In_2269,N_307);
and U2181 (N_2181,In_790,N_603);
nor U2182 (N_2182,In_497,N_1512);
nor U2183 (N_2183,N_1715,N_1844);
and U2184 (N_2184,In_4405,N_1729);
and U2185 (N_2185,N_209,In_4596);
nor U2186 (N_2186,N_1301,N_341);
or U2187 (N_2187,N_1891,In_4006);
and U2188 (N_2188,In_1194,N_43);
nand U2189 (N_2189,N_1708,N_1175);
nor U2190 (N_2190,N_1458,N_773);
xnor U2191 (N_2191,N_144,N_403);
nor U2192 (N_2192,In_3568,N_941);
and U2193 (N_2193,N_10,N_644);
and U2194 (N_2194,N_1314,In_4004);
and U2195 (N_2195,N_867,In_3605);
and U2196 (N_2196,N_568,N_1164);
nand U2197 (N_2197,N_20,N_1174);
and U2198 (N_2198,N_531,N_1599);
xnor U2199 (N_2199,In_2374,N_562);
xnor U2200 (N_2200,N_800,N_702);
nand U2201 (N_2201,N_1197,In_1868);
xor U2202 (N_2202,In_203,In_3726);
and U2203 (N_2203,In_2116,N_1626);
or U2204 (N_2204,In_3559,In_1939);
nor U2205 (N_2205,N_1075,In_1810);
or U2206 (N_2206,N_827,In_3171);
nand U2207 (N_2207,In_270,N_1752);
nand U2208 (N_2208,N_342,In_2581);
nand U2209 (N_2209,N_1380,N_372);
and U2210 (N_2210,N_1921,In_3651);
and U2211 (N_2211,N_1705,In_4466);
nand U2212 (N_2212,In_3821,N_1149);
or U2213 (N_2213,N_1128,In_4455);
nor U2214 (N_2214,In_3212,N_1361);
and U2215 (N_2215,In_3581,N_1689);
xnor U2216 (N_2216,N_832,In_1107);
xnor U2217 (N_2217,N_1419,N_1209);
nand U2218 (N_2218,In_1685,In_508);
nand U2219 (N_2219,N_1105,N_1242);
nand U2220 (N_2220,In_154,In_515);
nand U2221 (N_2221,N_1841,In_490);
xor U2222 (N_2222,N_1724,N_1934);
and U2223 (N_2223,In_1564,N_805);
xnor U2224 (N_2224,N_1811,N_1016);
xor U2225 (N_2225,In_3274,N_249);
xnor U2226 (N_2226,N_1249,N_613);
nand U2227 (N_2227,N_736,In_1520);
or U2228 (N_2228,N_1755,N_1202);
nand U2229 (N_2229,In_946,N_1156);
nor U2230 (N_2230,N_276,In_4928);
xor U2231 (N_2231,N_1478,N_95);
xnor U2232 (N_2232,N_1513,N_1495);
or U2233 (N_2233,In_4137,N_237);
xor U2234 (N_2234,In_1225,N_700);
xor U2235 (N_2235,N_1723,In_2919);
nor U2236 (N_2236,In_1161,N_57);
and U2237 (N_2237,N_696,In_2094);
nand U2238 (N_2238,N_1368,N_891);
xor U2239 (N_2239,In_869,N_1233);
nand U2240 (N_2240,In_2337,N_1312);
and U2241 (N_2241,N_1805,N_617);
xnor U2242 (N_2242,N_402,N_1280);
xnor U2243 (N_2243,N_495,N_0);
nand U2244 (N_2244,In_214,N_983);
nor U2245 (N_2245,In_1606,N_1140);
or U2246 (N_2246,N_373,N_764);
xnor U2247 (N_2247,N_1111,N_1644);
nand U2248 (N_2248,N_496,N_648);
nor U2249 (N_2249,N_117,In_137);
nor U2250 (N_2250,In_1636,N_904);
nand U2251 (N_2251,N_242,N_290);
nor U2252 (N_2252,N_1462,N_566);
xnor U2253 (N_2253,N_1822,N_98);
and U2254 (N_2254,In_3655,In_4105);
nor U2255 (N_2255,In_2178,N_789);
nand U2256 (N_2256,N_1065,N_907);
or U2257 (N_2257,N_735,In_1860);
nand U2258 (N_2258,N_1056,N_1665);
nand U2259 (N_2259,In_2526,In_431);
nor U2260 (N_2260,N_444,In_4809);
nor U2261 (N_2261,N_1993,N_1584);
nand U2262 (N_2262,N_1027,N_1578);
nor U2263 (N_2263,N_384,In_949);
nand U2264 (N_2264,In_827,N_585);
or U2265 (N_2265,N_1173,N_1252);
nor U2266 (N_2266,In_1385,In_3610);
or U2267 (N_2267,N_998,In_386);
nor U2268 (N_2268,N_623,N_63);
or U2269 (N_2269,In_4401,N_815);
and U2270 (N_2270,N_1237,N_923);
and U2271 (N_2271,N_1015,N_763);
and U2272 (N_2272,N_1737,In_3695);
xnor U2273 (N_2273,N_8,N_159);
nand U2274 (N_2274,In_2807,In_1445);
xnor U2275 (N_2275,N_380,In_697);
and U2276 (N_2276,N_491,In_3826);
nand U2277 (N_2277,N_1979,N_406);
or U2278 (N_2278,In_2795,N_643);
xor U2279 (N_2279,N_72,N_1031);
and U2280 (N_2280,In_1618,N_1438);
nor U2281 (N_2281,N_320,N_19);
or U2282 (N_2282,In_970,N_1410);
and U2283 (N_2283,In_1304,In_3976);
nor U2284 (N_2284,In_4501,N_733);
and U2285 (N_2285,N_23,N_1499);
nor U2286 (N_2286,In_1909,N_1926);
and U2287 (N_2287,In_1012,N_843);
xnor U2288 (N_2288,N_1170,N_1098);
nor U2289 (N_2289,In_2444,In_465);
and U2290 (N_2290,N_1295,In_3418);
or U2291 (N_2291,In_2203,In_2164);
xor U2292 (N_2292,N_885,N_1682);
nand U2293 (N_2293,N_92,N_1882);
and U2294 (N_2294,N_121,N_271);
xor U2295 (N_2295,In_696,N_278);
and U2296 (N_2296,In_1397,In_3166);
and U2297 (N_2297,N_1735,N_178);
and U2298 (N_2298,N_1396,In_4316);
or U2299 (N_2299,N_1068,N_1992);
xor U2300 (N_2300,N_1691,N_283);
nor U2301 (N_2301,N_1546,N_163);
nor U2302 (N_2302,N_490,In_4799);
or U2303 (N_2303,N_662,In_4902);
xnor U2304 (N_2304,N_1789,N_1622);
or U2305 (N_2305,In_126,N_1185);
or U2306 (N_2306,N_6,N_969);
nand U2307 (N_2307,N_1198,N_974);
nand U2308 (N_2308,In_4662,N_336);
nand U2309 (N_2309,N_1172,N_143);
nand U2310 (N_2310,In_3865,N_1565);
and U2311 (N_2311,N_1765,N_175);
or U2312 (N_2312,N_180,N_1254);
and U2313 (N_2313,N_1081,In_2403);
or U2314 (N_2314,In_3670,N_981);
or U2315 (N_2315,In_1166,N_1995);
xor U2316 (N_2316,N_1588,In_4569);
nor U2317 (N_2317,In_3410,N_381);
or U2318 (N_2318,N_1107,In_1239);
or U2319 (N_2319,In_1248,In_4734);
xor U2320 (N_2320,N_1726,In_4899);
and U2321 (N_2321,N_1122,N_308);
xor U2322 (N_2322,N_1399,N_897);
nor U2323 (N_2323,N_1074,In_913);
nand U2324 (N_2324,N_108,In_335);
nand U2325 (N_2325,In_3893,N_846);
or U2326 (N_2326,N_1594,N_47);
or U2327 (N_2327,N_1694,In_2402);
nor U2328 (N_2328,N_1292,In_4350);
or U2329 (N_2329,In_2618,N_169);
or U2330 (N_2330,N_487,N_1968);
nand U2331 (N_2331,N_529,N_1129);
and U2332 (N_2332,In_1351,In_4832);
nor U2333 (N_2333,N_1392,N_401);
or U2334 (N_2334,In_157,In_4739);
xor U2335 (N_2335,In_4164,In_4286);
or U2336 (N_2336,N_774,N_303);
and U2337 (N_2337,N_1575,In_4197);
nand U2338 (N_2338,N_1365,N_1195);
nand U2339 (N_2339,N_716,N_1668);
xnor U2340 (N_2340,N_385,N_756);
or U2341 (N_2341,N_900,N_61);
xnor U2342 (N_2342,In_3223,In_4699);
and U2343 (N_2343,N_1730,N_368);
or U2344 (N_2344,N_1573,In_1878);
nor U2345 (N_2345,In_745,N_1922);
xor U2346 (N_2346,In_1932,N_821);
nor U2347 (N_2347,In_2455,In_840);
nand U2348 (N_2348,N_1266,In_1362);
nand U2349 (N_2349,N_1073,N_824);
or U2350 (N_2350,In_1720,N_947);
and U2351 (N_2351,N_1039,In_883);
and U2352 (N_2352,In_3198,N_1219);
nand U2353 (N_2353,N_877,N_987);
nand U2354 (N_2354,N_517,In_2980);
or U2355 (N_2355,N_942,In_228);
nand U2356 (N_2356,In_1022,In_442);
and U2357 (N_2357,In_4337,N_1385);
and U2358 (N_2358,In_3999,N_976);
and U2359 (N_2359,In_1578,In_1784);
and U2360 (N_2360,N_1300,N_726);
xnor U2361 (N_2361,In_2765,N_946);
nor U2362 (N_2362,In_2363,In_3095);
and U2363 (N_2363,In_4807,N_1500);
xor U2364 (N_2364,N_706,N_1748);
and U2365 (N_2365,N_1311,N_598);
nand U2366 (N_2366,In_4529,N_522);
xor U2367 (N_2367,N_1452,N_1157);
and U2368 (N_2368,N_1116,In_2800);
nor U2369 (N_2369,N_1313,N_851);
or U2370 (N_2370,In_4773,In_1285);
nor U2371 (N_2371,In_985,N_96);
nor U2372 (N_2372,N_682,In_520);
nor U2373 (N_2373,N_1398,In_1374);
nor U2374 (N_2374,In_3498,In_1922);
nor U2375 (N_2375,N_1099,In_4852);
and U2376 (N_2376,N_1126,In_1159);
nand U2377 (N_2377,N_1060,N_1658);
nor U2378 (N_2378,In_4957,In_1803);
nor U2379 (N_2379,In_4842,N_1066);
or U2380 (N_2380,In_1219,In_2161);
nand U2381 (N_2381,In_1961,In_2592);
nand U2382 (N_2382,In_1475,In_2144);
xor U2383 (N_2383,N_633,In_3910);
nor U2384 (N_2384,N_1041,N_1672);
nor U2385 (N_2385,In_1382,N_1675);
nand U2386 (N_2386,N_329,N_1555);
nor U2387 (N_2387,N_714,In_3880);
nor U2388 (N_2388,In_4393,N_812);
and U2389 (N_2389,In_2762,N_14);
xor U2390 (N_2390,N_273,N_31);
and U2391 (N_2391,N_836,N_1449);
xor U2392 (N_2392,N_1829,N_115);
nand U2393 (N_2393,In_4240,N_1670);
xnor U2394 (N_2394,N_1702,N_212);
and U2395 (N_2395,N_1302,In_2569);
and U2396 (N_2396,N_197,N_191);
nor U2397 (N_2397,N_604,N_1942);
nand U2398 (N_2398,In_3441,N_1950);
or U2399 (N_2399,N_1780,N_1271);
and U2400 (N_2400,N_1453,N_1044);
nand U2401 (N_2401,N_454,In_2552);
xnor U2402 (N_2402,In_4973,N_1425);
or U2403 (N_2403,N_421,In_2017);
nand U2404 (N_2404,N_1619,In_2755);
nor U2405 (N_2405,N_1653,In_4063);
nor U2406 (N_2406,N_335,In_4918);
or U2407 (N_2407,N_398,N_289);
xnor U2408 (N_2408,N_410,N_474);
xor U2409 (N_2409,N_768,N_1308);
or U2410 (N_2410,In_2044,N_1467);
or U2411 (N_2411,N_1217,N_284);
nand U2412 (N_2412,N_1643,N_1152);
and U2413 (N_2413,In_3974,In_1446);
xnor U2414 (N_2414,N_671,N_1181);
xor U2415 (N_2415,N_1335,N_438);
xnor U2416 (N_2416,N_431,N_1999);
xnor U2417 (N_2417,In_939,In_2900);
and U2418 (N_2418,N_1954,N_1029);
nand U2419 (N_2419,N_866,N_704);
or U2420 (N_2420,In_252,N_140);
and U2421 (N_2421,N_819,N_1774);
and U2422 (N_2422,N_1583,In_4142);
or U2423 (N_2423,In_1089,In_305);
xnor U2424 (N_2424,N_1040,N_1610);
nand U2425 (N_2425,N_731,In_4769);
and U2426 (N_2426,N_1320,In_815);
nand U2427 (N_2427,In_3352,N_675);
and U2428 (N_2428,N_1764,N_1420);
or U2429 (N_2429,N_227,N_1349);
nand U2430 (N_2430,In_2841,N_129);
nand U2431 (N_2431,N_260,N_1418);
nand U2432 (N_2432,N_636,N_182);
nor U2433 (N_2433,N_968,N_688);
nor U2434 (N_2434,N_93,In_2830);
or U2435 (N_2435,N_1637,In_3443);
and U2436 (N_2436,N_767,In_1760);
or U2437 (N_2437,N_1283,N_1540);
xnor U2438 (N_2438,In_3710,In_1856);
nand U2439 (N_2439,N_975,In_1523);
nor U2440 (N_2440,N_931,In_2603);
and U2441 (N_2441,N_1645,N_493);
nor U2442 (N_2442,N_1315,In_2285);
xnor U2443 (N_2443,In_328,In_1807);
nand U2444 (N_2444,N_1598,N_484);
nor U2445 (N_2445,N_305,In_3507);
and U2446 (N_2446,In_647,N_1893);
xnor U2447 (N_2447,N_219,N_107);
nand U2448 (N_2448,In_4959,N_411);
and U2449 (N_2449,N_147,In_4503);
and U2450 (N_2450,N_841,N_814);
nand U2451 (N_2451,N_1356,N_1293);
nor U2452 (N_2452,In_100,N_988);
nand U2453 (N_2453,In_3918,N_1632);
nor U2454 (N_2454,N_1072,N_855);
or U2455 (N_2455,N_1097,N_1784);
nand U2456 (N_2456,N_1797,N_464);
or U2457 (N_2457,N_1255,N_808);
or U2458 (N_2458,N_261,N_513);
nand U2459 (N_2459,N_1771,In_251);
nor U2460 (N_2460,In_3556,N_1566);
nand U2461 (N_2461,In_413,N_631);
xnor U2462 (N_2462,N_739,N_1900);
or U2463 (N_2463,In_3874,N_301);
or U2464 (N_2464,N_823,N_1490);
nand U2465 (N_2465,In_1049,N_224);
xnor U2466 (N_2466,In_2857,N_938);
nand U2467 (N_2467,N_46,N_1135);
xnor U2468 (N_2468,In_1060,In_289);
nand U2469 (N_2469,In_1057,N_637);
nand U2470 (N_2470,In_3721,In_4517);
nand U2471 (N_2471,N_629,N_1704);
xnor U2472 (N_2472,N_871,N_527);
xnor U2473 (N_2473,N_1206,N_1613);
and U2474 (N_2474,N_1203,In_1550);
xor U2475 (N_2475,N_1162,In_3050);
xnor U2476 (N_2476,N_433,N_354);
xor U2477 (N_2477,N_1407,N_1150);
or U2478 (N_2478,N_376,In_3904);
or U2479 (N_2479,In_1781,N_1370);
nand U2480 (N_2480,N_171,In_4519);
and U2481 (N_2481,N_1369,In_2018);
or U2482 (N_2482,N_122,In_261);
and U2483 (N_2483,N_392,N_1477);
nor U2484 (N_2484,N_1669,N_1087);
and U2485 (N_2485,N_1919,N_443);
xnor U2486 (N_2486,In_175,N_1360);
nand U2487 (N_2487,N_321,N_295);
nor U2488 (N_2488,N_1416,N_1278);
nor U2489 (N_2489,N_737,N_7);
nor U2490 (N_2490,N_1674,In_4287);
xor U2491 (N_2491,N_165,N_337);
nand U2492 (N_2492,N_960,N_569);
and U2493 (N_2493,N_687,N_1953);
xnor U2494 (N_2494,N_1615,N_414);
nand U2495 (N_2495,N_970,In_419);
xnor U2496 (N_2496,N_297,N_11);
and U2497 (N_2497,N_1808,N_1794);
nand U2498 (N_2498,N_1747,In_661);
and U2499 (N_2499,In_3289,N_1325);
nor U2500 (N_2500,N_1299,In_2446);
nand U2501 (N_2501,N_1910,N_325);
xor U2502 (N_2502,In_3816,N_1806);
and U2503 (N_2503,In_1938,N_570);
and U2504 (N_2504,N_620,In_3886);
or U2505 (N_2505,N_468,In_733);
nand U2506 (N_2506,In_2880,In_1228);
xnor U2507 (N_2507,N_1194,N_1006);
and U2508 (N_2508,N_471,N_345);
nand U2509 (N_2509,N_788,N_943);
xor U2510 (N_2510,N_741,In_4915);
xnor U2511 (N_2511,In_4565,N_1978);
nand U2512 (N_2512,N_170,N_1210);
xnor U2513 (N_2513,In_3096,N_556);
or U2514 (N_2514,N_1372,N_1685);
nor U2515 (N_2515,In_1145,N_1232);
or U2516 (N_2516,In_777,N_825);
or U2517 (N_2517,N_547,In_2866);
or U2518 (N_2518,In_1796,N_752);
nand U2519 (N_2519,N_1881,N_1306);
xor U2520 (N_2520,In_1955,N_1838);
and U2521 (N_2521,N_1756,N_1840);
nor U2522 (N_2522,N_1522,In_767);
xnor U2523 (N_2523,In_479,N_1980);
or U2524 (N_2524,In_2253,N_811);
nor U2525 (N_2525,N_3,N_1857);
and U2526 (N_2526,N_1058,N_1281);
nand U2527 (N_2527,N_1955,In_4297);
nor U2528 (N_2528,N_1819,N_1719);
and U2529 (N_2529,N_1519,N_79);
xnor U2530 (N_2530,N_1826,N_469);
xnor U2531 (N_2531,N_161,N_458);
nor U2532 (N_2532,N_750,N_1604);
nor U2533 (N_2533,N_1683,N_150);
or U2534 (N_2534,In_851,N_748);
and U2535 (N_2535,N_246,In_504);
xnor U2536 (N_2536,N_1851,N_148);
xnor U2537 (N_2537,N_371,N_432);
and U2538 (N_2538,N_1018,N_456);
nor U2539 (N_2539,N_1208,In_3183);
nor U2540 (N_2540,N_35,N_1330);
nor U2541 (N_2541,N_816,In_4380);
xor U2542 (N_2542,N_608,In_1945);
and U2543 (N_2543,In_28,In_4165);
or U2544 (N_2544,N_1516,In_1888);
xnor U2545 (N_2545,N_677,N_646);
and U2546 (N_2546,N_428,N_676);
nor U2547 (N_2547,N_1641,N_1245);
nand U2548 (N_2548,N_1045,In_2153);
xnor U2549 (N_2549,In_2821,N_1951);
and U2550 (N_2550,N_1484,In_631);
nor U2551 (N_2551,In_3415,In_1460);
nand U2552 (N_2552,N_939,N_1507);
nand U2553 (N_2553,In_805,N_581);
or U2554 (N_2554,N_378,N_1384);
nand U2555 (N_2555,N_1913,N_876);
xor U2556 (N_2556,In_3310,N_1938);
nor U2557 (N_2557,N_886,N_53);
nor U2558 (N_2558,N_860,N_587);
xor U2559 (N_2559,In_3092,N_437);
and U2560 (N_2560,In_3210,N_695);
or U2561 (N_2561,N_482,N_187);
nand U2562 (N_2562,N_1580,In_1511);
and U2563 (N_2563,N_796,In_1712);
nor U2564 (N_2564,N_1629,N_184);
nand U2565 (N_2565,In_4841,N_1070);
nor U2566 (N_2566,N_839,N_1592);
and U2567 (N_2567,N_864,N_795);
or U2568 (N_2568,N_1258,In_118);
nand U2569 (N_2569,In_4253,In_784);
or U2570 (N_2570,N_818,N_48);
xnor U2571 (N_2571,N_312,N_62);
nand U2572 (N_2572,In_4559,N_1608);
and U2573 (N_2573,N_1914,N_1807);
nand U2574 (N_2574,In_2593,N_1563);
nand U2575 (N_2575,In_2497,N_1218);
nand U2576 (N_2576,In_4283,N_954);
nor U2577 (N_2577,In_3326,N_90);
nand U2578 (N_2578,N_1250,N_1422);
and U2579 (N_2579,N_52,N_534);
xor U2580 (N_2580,N_1024,In_1867);
or U2581 (N_2581,N_964,N_56);
nor U2582 (N_2582,In_2272,In_4512);
and U2583 (N_2583,N_903,N_1746);
xnor U2584 (N_2584,In_1314,N_1119);
and U2585 (N_2585,N_680,N_1874);
nand U2586 (N_2586,N_1815,In_4223);
xnor U2587 (N_2587,N_322,N_1007);
nand U2588 (N_2588,In_3298,N_1446);
and U2589 (N_2589,N_1470,In_2548);
or U2590 (N_2590,N_155,In_4787);
nor U2591 (N_2591,N_1611,In_2784);
nand U2592 (N_2592,N_535,In_3364);
nand U2593 (N_2593,N_799,N_1760);
nand U2594 (N_2594,In_269,In_3156);
or U2595 (N_2595,In_1635,N_430);
nand U2596 (N_2596,In_3185,In_3888);
and U2597 (N_2597,N_1358,N_97);
nor U2598 (N_2598,In_2059,In_792);
and U2599 (N_2599,N_54,In_1408);
and U2600 (N_2600,In_3979,N_1505);
nor U2601 (N_2601,N_1082,N_1322);
or U2602 (N_2602,N_1294,In_1656);
xnor U2603 (N_2603,N_1286,N_1718);
nor U2604 (N_2604,N_1442,In_3802);
xor U2605 (N_2605,N_73,N_1667);
nand U2606 (N_2606,In_2736,N_1700);
nand U2607 (N_2607,N_705,In_4753);
xor U2608 (N_2608,In_542,In_741);
and U2609 (N_2609,N_1837,N_810);
and U2610 (N_2610,N_1429,In_1851);
and U2611 (N_2611,In_3883,N_70);
xnor U2612 (N_2612,In_4677,N_898);
or U2613 (N_2613,N_618,In_923);
and U2614 (N_2614,N_207,N_259);
nor U2615 (N_2615,N_502,N_760);
and U2616 (N_2616,In_3463,N_651);
xor U2617 (N_2617,In_2188,N_668);
or U2618 (N_2618,N_1770,N_1414);
nor U2619 (N_2619,N_318,N_514);
nor U2620 (N_2620,N_131,N_1376);
nand U2621 (N_2621,In_4270,N_1002);
nor U2622 (N_2622,N_1977,N_1277);
and U2623 (N_2623,N_51,N_1423);
and U2624 (N_2624,In_3055,N_1614);
nand U2625 (N_2625,In_3801,N_216);
xor U2626 (N_2626,In_4462,N_1550);
and U2627 (N_2627,N_882,N_1166);
and U2628 (N_2628,In_4460,In_3548);
nand U2629 (N_2629,N_835,N_1270);
or U2630 (N_2630,N_217,N_1889);
xnor U2631 (N_2631,N_1989,N_497);
and U2632 (N_2632,N_254,In_2431);
nand U2633 (N_2633,In_4162,N_1853);
and U2634 (N_2634,In_3405,N_1927);
nor U2635 (N_2635,In_408,N_560);
and U2636 (N_2636,N_1091,N_1201);
nand U2637 (N_2637,In_2610,N_1973);
or U2638 (N_2638,N_383,N_609);
or U2639 (N_2639,In_3371,N_447);
or U2640 (N_2640,N_868,N_639);
nand U2641 (N_2641,N_1092,N_1537);
and U2642 (N_2642,In_3748,N_837);
nor U2643 (N_2643,N_1758,In_3279);
and U2644 (N_2644,N_1856,N_1231);
and U2645 (N_2645,N_908,N_906);
or U2646 (N_2646,N_1867,N_1061);
nand U2647 (N_2647,N_1759,In_1658);
nor U2648 (N_2648,N_1686,In_4109);
nand U2649 (N_2649,In_655,N_584);
xnor U2650 (N_2650,N_356,N_1404);
and U2651 (N_2651,In_3898,N_1288);
or U2652 (N_2652,N_1260,N_657);
nand U2653 (N_2653,N_833,N_1076);
nand U2654 (N_2654,In_4605,In_2907);
nand U2655 (N_2655,N_75,N_1110);
nand U2656 (N_2656,N_1444,In_3176);
and U2657 (N_2657,In_3248,N_1930);
nand U2658 (N_2658,N_364,N_1823);
nand U2659 (N_2659,In_4383,N_896);
and U2660 (N_2660,N_1287,N_1732);
and U2661 (N_2661,In_1412,N_1982);
nor U2662 (N_2662,N_553,N_1184);
and U2663 (N_2663,In_781,In_3907);
or U2664 (N_2664,N_515,N_937);
or U2665 (N_2665,N_510,N_930);
xor U2666 (N_2666,In_4189,N_1079);
nor U2667 (N_2667,N_1524,In_4180);
or U2668 (N_2668,In_680,N_1188);
and U2669 (N_2669,N_1476,N_462);
or U2670 (N_2670,N_306,N_905);
nand U2671 (N_2671,N_111,N_516);
xnor U2672 (N_2672,N_369,In_398);
xor U2673 (N_2673,In_1706,N_386);
and U2674 (N_2674,In_3862,In_2854);
nand U2675 (N_2675,In_1607,N_1243);
xor U2676 (N_2676,N_1981,In_3738);
and U2677 (N_2677,N_1778,N_382);
nand U2678 (N_2678,N_1328,In_11);
xor U2679 (N_2679,In_2320,N_567);
and U2680 (N_2680,In_1220,N_854);
nand U2681 (N_2681,N_1154,N_901);
nand U2682 (N_2682,N_1114,In_1745);
nor U2683 (N_2683,In_3455,N_265);
nand U2684 (N_2684,N_722,N_1680);
xor U2685 (N_2685,N_1464,In_2160);
nor U2686 (N_2686,N_1869,In_2010);
nand U2687 (N_2687,N_642,In_1613);
xor U2688 (N_2688,In_3860,N_1733);
nor U2689 (N_2689,In_896,N_102);
or U2690 (N_2690,N_655,N_1742);
and U2691 (N_2691,N_879,In_3623);
and U2692 (N_2692,In_2180,N_802);
nor U2693 (N_2693,N_753,N_649);
nor U2694 (N_2694,N_1080,N_1063);
nand U2695 (N_2695,N_1296,N_783);
nor U2696 (N_2696,N_592,N_200);
nand U2697 (N_2697,N_1638,In_2815);
nor U2698 (N_2698,In_394,N_1532);
and U2699 (N_2699,N_1899,N_1391);
nor U2700 (N_2700,N_523,N_694);
and U2701 (N_2701,In_611,In_3379);
xnor U2702 (N_2702,N_746,N_405);
nor U2703 (N_2703,N_994,N_895);
nand U2704 (N_2704,In_1080,N_1741);
xnor U2705 (N_2705,N_720,In_3502);
or U2706 (N_2706,In_3147,In_1254);
nand U2707 (N_2707,In_1247,In_1794);
and U2708 (N_2708,In_1772,N_554);
nor U2709 (N_2709,In_143,N_579);
or U2710 (N_2710,In_3091,N_404);
nor U2711 (N_2711,N_1049,N_1509);
nor U2712 (N_2712,N_747,N_1654);
nand U2713 (N_2713,N_1738,N_1944);
and U2714 (N_2714,In_1630,N_1636);
or U2715 (N_2715,N_1931,In_788);
nor U2716 (N_2716,N_1264,N_1473);
nor U2717 (N_2717,N_1214,N_559);
xnor U2718 (N_2718,In_2767,N_650);
xnor U2719 (N_2719,N_4,N_266);
and U2720 (N_2720,In_2864,N_1351);
and U2721 (N_2721,In_4825,N_638);
and U2722 (N_2722,N_1633,N_5);
nand U2723 (N_2723,N_1259,N_713);
or U2724 (N_2724,In_4580,In_2465);
nor U2725 (N_2725,N_1394,In_352);
nand U2726 (N_2726,N_1345,N_1200);
or U2727 (N_2727,N_858,In_4443);
and U2728 (N_2728,In_2107,In_2287);
or U2729 (N_2729,In_3554,In_2659);
nor U2730 (N_2730,In_116,N_225);
nand U2731 (N_2731,N_89,N_1331);
or U2732 (N_2732,N_723,N_1753);
nor U2733 (N_2733,In_3046,N_277);
or U2734 (N_2734,N_1386,N_1253);
nand U2735 (N_2735,N_1817,In_2655);
nor U2736 (N_2736,N_834,N_894);
or U2737 (N_2737,N_489,N_669);
nor U2738 (N_2738,In_4171,In_3877);
or U2739 (N_2739,N_228,N_173);
and U2740 (N_2740,N_294,N_1603);
nor U2741 (N_2741,N_119,N_1496);
and U2742 (N_2742,N_924,N_106);
or U2743 (N_2743,N_267,N_1799);
and U2744 (N_2744,N_583,In_4260);
nor U2745 (N_2745,N_202,In_2611);
nor U2746 (N_2746,In_4972,In_2663);
nand U2747 (N_2747,In_1482,In_1964);
or U2748 (N_2748,N_1560,N_87);
nor U2749 (N_2749,N_483,N_1355);
and U2750 (N_2750,In_4269,N_293);
and U2751 (N_2751,In_4748,In_2617);
or U2752 (N_2752,In_4552,In_618);
xnor U2753 (N_2753,N_370,N_755);
or U2754 (N_2754,N_208,N_1946);
or U2755 (N_2755,In_2922,N_1178);
or U2756 (N_2756,N_1333,In_2009);
xnor U2757 (N_2757,In_4582,N_1364);
nand U2758 (N_2758,N_391,N_1268);
and U2759 (N_2759,In_2469,N_1917);
and U2760 (N_2760,In_2515,N_1047);
nand U2761 (N_2761,In_2936,N_1706);
xnor U2762 (N_2762,N_512,N_1035);
xor U2763 (N_2763,N_27,N_1121);
nor U2764 (N_2764,In_4079,N_1928);
and U2765 (N_2765,In_3663,N_331);
nor U2766 (N_2766,N_211,N_1936);
xnor U2767 (N_2767,N_1052,In_4967);
or U2768 (N_2768,N_925,N_1377);
or U2769 (N_2769,N_999,In_916);
xor U2770 (N_2770,N_422,N_965);
or U2771 (N_2771,In_2198,N_1701);
and U2772 (N_2772,In_320,N_425);
and U2773 (N_2773,N_679,In_44);
xnor U2774 (N_2774,In_3573,In_4147);
or U2775 (N_2775,N_580,In_4550);
or U2776 (N_2776,N_611,N_1138);
xor U2777 (N_2777,N_1744,N_1791);
or U2778 (N_2778,N_873,N_1852);
nand U2779 (N_2779,N_1492,N_1551);
nand U2780 (N_2780,In_2406,N_533);
and U2781 (N_2781,N_1605,N_83);
nand U2782 (N_2782,In_3609,In_619);
or U2783 (N_2783,N_683,In_3708);
nor U2784 (N_2784,N_1474,N_304);
nor U2785 (N_2785,N_359,N_1085);
or U2786 (N_2786,N_727,In_2418);
and U2787 (N_2787,N_1557,N_1042);
nand U2788 (N_2788,N_1627,In_1951);
or U2789 (N_2789,N_439,N_1180);
nor U2790 (N_2790,N_28,N_1990);
xor U2791 (N_2791,In_2523,N_139);
xor U2792 (N_2792,N_1642,N_911);
xnor U2793 (N_2793,N_299,N_1722);
xnor U2794 (N_2794,N_1480,N_919);
nand U2795 (N_2795,N_786,In_1283);
or U2796 (N_2796,In_2950,In_4926);
or U2797 (N_2797,N_1038,In_1599);
or U2798 (N_2798,In_346,In_120);
and U2799 (N_2799,N_1582,N_330);
or U2800 (N_2800,N_316,N_1133);
or U2801 (N_2801,N_1612,N_1601);
and U2802 (N_2802,N_807,N_1193);
nand U2803 (N_2803,N_506,In_4431);
xor U2804 (N_2804,N_588,N_689);
nor U2805 (N_2805,In_3294,N_653);
and U2806 (N_2806,N_113,In_4790);
and U2807 (N_2807,N_125,N_1435);
and U2808 (N_2808,N_1602,N_543);
nor U2809 (N_2809,N_1307,In_4700);
nand U2810 (N_2810,N_1284,N_857);
or U2811 (N_2811,N_1846,N_1925);
nand U2812 (N_2812,N_257,N_1939);
xnor U2813 (N_2813,N_840,N_1639);
nand U2814 (N_2814,N_902,In_1224);
nand U2815 (N_2815,N_1679,N_1591);
nor U2816 (N_2816,In_86,In_893);
xnor U2817 (N_2817,N_539,N_1362);
xor U2818 (N_2818,N_1059,N_1567);
nor U2819 (N_2819,In_4099,N_355);
nand U2820 (N_2820,In_3355,In_2254);
xor U2821 (N_2821,In_380,N_630);
nand U2822 (N_2822,N_883,N_215);
nand U2823 (N_2823,N_1625,N_85);
and U2824 (N_2824,N_918,In_1215);
and U2825 (N_2825,N_1163,N_550);
nand U2826 (N_2826,In_1997,N_327);
xor U2827 (N_2827,N_1896,N_1469);
or U2828 (N_2828,N_775,In_758);
xnor U2829 (N_2829,N_1215,N_1402);
or U2830 (N_2830,In_3214,N_1317);
nand U2831 (N_2831,In_4813,N_1848);
xnor U2832 (N_2832,N_1228,N_1506);
nand U2833 (N_2833,N_1332,N_25);
or U2834 (N_2834,In_30,In_405);
or U2835 (N_2835,In_4496,In_3033);
and U2836 (N_2836,N_672,In_3146);
and U2837 (N_2837,In_1466,N_190);
and U2838 (N_2838,N_888,N_830);
nor U2839 (N_2839,N_183,N_1711);
and U2840 (N_2840,N_262,In_4964);
or U2841 (N_2841,N_1818,In_4390);
nand U2842 (N_2842,N_1545,N_521);
nor U2843 (N_2843,N_749,N_1421);
and U2844 (N_2844,In_1689,In_4615);
nor U2845 (N_2845,N_1593,In_4046);
nor U2846 (N_2846,N_1112,N_1657);
nand U2847 (N_2847,N_1009,In_2615);
nand U2848 (N_2848,In_990,N_238);
or U2849 (N_2849,In_3591,N_149);
and U2850 (N_2850,N_334,N_1631);
nor U2851 (N_2851,N_1441,In_1632);
xnor U2852 (N_2852,N_1878,N_1792);
or U2853 (N_2853,In_3627,N_1491);
and U2854 (N_2854,N_1227,In_3217);
or U2855 (N_2855,N_829,N_110);
or U2856 (N_2856,N_426,N_132);
nand U2857 (N_2857,N_1662,N_1244);
or U2858 (N_2858,N_201,N_576);
or U2859 (N_2859,In_1572,In_3864);
and U2860 (N_2860,N_1544,N_1528);
nor U2861 (N_2861,N_772,N_1501);
nand U2862 (N_2862,N_17,In_2438);
or U2863 (N_2863,In_682,In_384);
or U2864 (N_2864,N_692,In_2184);
nand U2865 (N_2865,In_213,In_1984);
xnor U2866 (N_2866,N_1975,N_1017);
nor U2867 (N_2867,N_1207,N_792);
xnor U2868 (N_2868,In_3209,N_88);
nor U2869 (N_2869,In_173,In_4824);
xor U2870 (N_2870,N_1409,N_193);
nand U2871 (N_2871,In_2071,N_460);
and U2872 (N_2872,N_971,N_248);
nor U2873 (N_2873,In_2227,In_207);
nor U2874 (N_2874,N_1493,N_49);
nor U2875 (N_2875,In_3525,N_784);
and U2876 (N_2876,N_166,N_1648);
nor U2877 (N_2877,N_1498,N_759);
or U2878 (N_2878,N_899,N_498);
or U2879 (N_2879,N_440,N_659);
nor U2880 (N_2880,In_988,N_828);
and U2881 (N_2881,N_1727,In_1309);
or U2882 (N_2882,N_1160,N_1461);
xor U2883 (N_2883,In_1229,In_2988);
xnor U2884 (N_2884,N_635,N_1443);
xor U2885 (N_2885,In_1148,In_1992);
xor U2886 (N_2886,In_1010,N_177);
nor U2887 (N_2887,N_377,N_1677);
and U2888 (N_2888,N_67,N_1466);
and U2889 (N_2889,N_1827,N_436);
nand U2890 (N_2890,In_838,N_174);
nor U2891 (N_2891,N_388,N_1761);
nand U2892 (N_2892,N_564,N_1972);
and U2893 (N_2893,In_4064,N_1721);
nor U2894 (N_2894,N_18,N_32);
nand U2895 (N_2895,N_658,N_275);
and U2896 (N_2896,In_2544,N_1710);
and U2897 (N_2897,N_1998,N_1022);
and U2898 (N_2898,N_1855,N_1161);
xnor U2899 (N_2899,N_928,In_2471);
or U2900 (N_2900,N_984,N_1189);
xnor U2901 (N_2901,N_1316,N_1230);
and U2902 (N_2902,N_607,In_133);
xor U2903 (N_2903,N_123,N_1357);
nor U2904 (N_2904,N_24,N_661);
nor U2905 (N_2905,N_934,N_1586);
and U2906 (N_2906,N_1865,N_1892);
and U2907 (N_2907,N_1887,N_707);
nor U2908 (N_2908,N_1650,In_847);
nor U2909 (N_2909,N_1875,N_236);
or U2910 (N_2910,In_3645,In_582);
nand U2911 (N_2911,N_1262,N_1326);
or U2912 (N_2912,N_1348,N_1693);
and U2913 (N_2913,N_909,N_285);
nor U2914 (N_2914,N_847,N_1439);
xnor U2915 (N_2915,N_1510,N_1952);
or U2916 (N_2916,In_2251,N_929);
and U2917 (N_2917,In_549,In_3571);
nor U2918 (N_2918,N_1511,N_137);
nor U2919 (N_2919,N_253,In_1808);
nor U2920 (N_2920,N_230,In_2408);
xor U2921 (N_2921,In_3794,In_3269);
nor U2922 (N_2922,N_1987,N_1447);
or U2923 (N_2923,In_1894,In_1504);
and U2924 (N_2924,In_1192,In_1625);
or U2925 (N_2925,N_451,N_251);
or U2926 (N_2926,In_4654,N_188);
xor U2927 (N_2927,In_4213,N_779);
and U2928 (N_2928,In_3521,N_1833);
xor U2929 (N_2929,N_1158,N_1263);
nor U2930 (N_2930,N_1933,N_582);
xnor U2931 (N_2931,N_339,N_272);
nand U2932 (N_2932,N_1963,N_1962);
or U2933 (N_2933,N_1323,N_622);
nor U2934 (N_2934,N_1935,N_1554);
nor U2935 (N_2935,N_761,N_1514);
nor U2936 (N_2936,In_1208,In_4783);
xor U2937 (N_2937,N_126,N_1957);
xnor U2938 (N_2938,In_3552,N_548);
xnor U2939 (N_2939,N_41,In_4660);
or U2940 (N_2940,In_1308,In_539);
nor U2941 (N_2941,N_26,In_695);
xnor U2942 (N_2942,N_360,N_991);
or U2943 (N_2943,N_1274,N_1026);
and U2944 (N_2944,In_2638,N_324);
and U2945 (N_2945,N_1766,In_1129);
and U2946 (N_2946,In_4670,N_40);
nor U2947 (N_2947,N_435,N_1415);
and U2948 (N_2948,In_4103,In_3029);
nand U2949 (N_2949,N_1890,N_298);
nor U2950 (N_2950,N_1966,N_199);
and U2951 (N_2951,N_258,In_1509);
or U2952 (N_2952,N_724,N_1585);
and U2953 (N_2953,In_4087,In_2636);
or U2954 (N_2954,In_452,N_1559);
xnor U2955 (N_2955,N_348,In_4409);
xnor U2956 (N_2956,N_962,N_541);
nand U2957 (N_2957,In_2833,In_3058);
nor U2958 (N_2958,In_642,In_4527);
or U2959 (N_2959,N_1754,N_420);
and U2960 (N_2960,In_1596,N_1353);
or U2961 (N_2961,In_367,N_624);
or U2962 (N_2962,N_872,In_2769);
and U2963 (N_2963,N_1883,In_1667);
or U2964 (N_2964,N_1318,In_4172);
nand U2965 (N_2965,N_1552,In_4864);
and U2966 (N_2966,In_4777,N_461);
nor U2967 (N_2967,N_452,In_4614);
xnor U2968 (N_2968,N_632,In_1893);
or U2969 (N_2969,N_1216,N_1338);
and U2970 (N_2970,N_1030,In_2640);
and U2971 (N_2971,N_1276,N_1408);
and U2972 (N_2972,In_4659,N_670);
xor U2973 (N_2973,N_555,N_1903);
nand U2974 (N_2974,N_1054,N_1775);
xor U2975 (N_2975,N_863,In_1734);
xor U2976 (N_2976,N_1155,In_1083);
xnor U2977 (N_2977,N_1812,N_1285);
or U2978 (N_2978,In_316,N_42);
nor U2979 (N_2979,N_875,N_831);
nand U2980 (N_2980,N_1961,In_4481);
nor U2981 (N_2981,N_1518,N_1898);
nand U2982 (N_2982,N_619,N_1847);
nor U2983 (N_2983,N_1787,N_344);
or U2984 (N_2984,N_203,In_3724);
and U2985 (N_2985,N_179,N_1530);
nor U2986 (N_2986,N_1740,In_1449);
xnor U2987 (N_2987,N_350,In_709);
nor U2988 (N_2988,In_324,In_2223);
nor U2989 (N_2989,N_1517,In_3980);
nor U2990 (N_2990,In_2937,N_1199);
xnor U2991 (N_2991,N_757,N_1996);
and U2992 (N_2992,N_1712,N_949);
xor U2993 (N_2993,In_1272,N_1269);
or U2994 (N_2994,N_561,N_597);
xnor U2995 (N_2995,In_259,N_1589);
and U2996 (N_2996,In_3963,N_1858);
or U2997 (N_2997,N_507,N_1354);
or U2998 (N_2998,N_1543,In_3914);
nand U2999 (N_2999,N_204,N_1192);
xnor U3000 (N_3000,N_1569,N_1538);
and U3001 (N_3001,N_656,N_699);
or U3002 (N_3002,N_1671,N_1267);
nor U3003 (N_3003,In_268,In_531);
xnor U3004 (N_3004,N_1430,N_80);
xnor U3005 (N_3005,In_4557,N_849);
nand U3006 (N_3006,In_4387,In_2261);
and U3007 (N_3007,N_367,In_3793);
xnor U3008 (N_3008,N_536,N_549);
and U3009 (N_3009,In_3117,N_1118);
or U3010 (N_3010,N_1897,In_81);
or U3011 (N_3011,N_782,N_957);
nand U3012 (N_3012,N_1151,N_485);
xnor U3013 (N_3013,In_3766,N_1986);
nand U3014 (N_3014,In_4531,N_1117);
or U3015 (N_3015,In_1789,N_820);
nor U3016 (N_3016,N_375,N_1236);
nand U3017 (N_3017,N_387,In_1211);
xnor U3018 (N_3018,N_922,In_1733);
xor U3019 (N_3019,In_103,N_1666);
nand U3020 (N_3020,N_1123,In_2935);
nor U3021 (N_3021,N_771,In_3683);
xnor U3022 (N_3022,In_4375,In_3634);
and U3023 (N_3023,In_1452,N_845);
or U3024 (N_3024,N_1863,In_1679);
xnor U3025 (N_3025,N_508,N_678);
nand U3026 (N_3026,N_1104,In_4033);
and U3027 (N_3027,N_395,N_1579);
xnor U3028 (N_3028,N_1413,N_424);
xor U3029 (N_3029,In_13,In_295);
or U3030 (N_3030,N_221,N_247);
nor U3031 (N_3031,N_1387,N_162);
nor U3032 (N_3032,In_3501,N_1745);
and U3033 (N_3033,N_1659,N_1139);
nand U3034 (N_3034,N_634,In_1242);
or U3035 (N_3035,N_1656,N_1831);
nor U3036 (N_3036,N_263,N_1508);
or U3037 (N_3037,In_3034,N_1168);
or U3038 (N_3038,N_1574,In_3220);
and U3039 (N_3039,N_153,N_1617);
nand U3040 (N_3040,N_351,In_1649);
xor U3041 (N_3041,In_4212,N_1895);
nor U3042 (N_3042,In_3800,In_3403);
xor U3043 (N_3043,N_1086,In_4611);
nor U3044 (N_3044,N_887,N_1750);
and U3045 (N_3045,N_1279,In_4158);
xnor U3046 (N_3046,N_1736,N_1572);
xnor U3047 (N_3047,N_1483,N_1854);
nand U3048 (N_3048,N_1187,In_1624);
or U3049 (N_3049,N_1472,N_1796);
or U3050 (N_3050,In_1855,In_2283);
and U3051 (N_3051,N_673,N_505);
and U3052 (N_3052,N_45,N_326);
nand U3053 (N_3053,N_250,N_1607);
nand U3054 (N_3054,N_357,N_1136);
nand U3055 (N_3055,N_156,In_737);
nand U3056 (N_3056,N_574,N_333);
and U3057 (N_3057,In_144,N_1424);
or U3058 (N_3058,In_4326,N_935);
or U3059 (N_3059,N_134,N_966);
and U3060 (N_3060,N_141,N_599);
xnor U3061 (N_3061,In_1017,In_1818);
and U3062 (N_3062,N_1147,N_315);
and U3063 (N_3063,N_1226,In_4371);
and U3064 (N_3064,N_530,N_1132);
xor U3065 (N_3065,N_1071,In_2666);
nand U3066 (N_3066,In_3283,N_806);
nand U3067 (N_3067,In_2141,N_450);
nor U3068 (N_3068,N_1920,N_1832);
nor U3069 (N_3069,N_917,N_674);
nand U3070 (N_3070,N_243,N_595);
or U3071 (N_3071,In_2827,N_1562);
or U3072 (N_3072,N_1949,In_3105);
nand U3073 (N_3073,N_1876,N_302);
nand U3074 (N_3074,N_235,N_856);
or U3075 (N_3075,In_1058,In_3303);
and U3076 (N_3076,In_811,N_1673);
or U3077 (N_3077,In_4100,N_932);
nor U3078 (N_3078,N_50,N_287);
or U3079 (N_3079,N_1062,N_1525);
and U3080 (N_3080,N_1145,N_1488);
nand U3081 (N_3081,In_1207,N_446);
nor U3082 (N_3082,In_1342,N_164);
and U3083 (N_3083,N_1347,N_1204);
and U3084 (N_3084,N_1021,N_1089);
nor U3085 (N_3085,N_711,N_1000);
nand U3086 (N_3086,N_710,N_1034);
nand U3087 (N_3087,In_1210,In_4490);
xor U3088 (N_3088,N_1521,N_1523);
nand U3089 (N_3089,N_365,N_1137);
nor U3090 (N_3090,N_1235,In_329);
xnor U3091 (N_3091,N_916,N_323);
xnor U3092 (N_3092,N_189,In_732);
nand U3093 (N_3093,In_3547,In_3662);
nand U3094 (N_3094,In_634,In_4514);
or U3095 (N_3095,N_1352,N_1456);
xnor U3096 (N_3096,In_1849,N_1635);
or U3097 (N_3097,In_2906,N_542);
and U3098 (N_3098,In_2933,In_1118);
and U3099 (N_3099,N_742,N_1912);
or U3100 (N_3100,N_12,In_1948);
or U3101 (N_3101,In_4021,N_44);
or U3102 (N_3102,N_1451,N_1393);
and U3103 (N_3103,N_133,In_1887);
or U3104 (N_3104,N_138,N_226);
nand U3105 (N_3105,In_3090,N_1486);
nand U3106 (N_3106,N_978,N_1023);
nor U3107 (N_3107,In_3339,N_1661);
or U3108 (N_3108,N_74,N_1621);
or U3109 (N_3109,N_551,In_3792);
or U3110 (N_3110,N_160,In_1758);
or U3111 (N_3111,In_1496,In_3332);
and U3112 (N_3112,N_1948,N_1005);
and U3113 (N_3113,In_4521,N_1872);
nor U3114 (N_3114,N_1976,In_1290);
nand U3115 (N_3115,N_1487,N_1220);
nand U3116 (N_3116,N_995,N_770);
xor U3117 (N_3117,N_252,N_959);
nor U3118 (N_3118,N_803,N_229);
nor U3119 (N_3119,In_3414,In_629);
nor U3120 (N_3120,N_448,In_2583);
nor U3121 (N_3121,In_493,N_1025);
xnor U3122 (N_3122,N_993,N_1699);
nand U3123 (N_3123,N_22,In_9);
or U3124 (N_3124,N_1821,N_1212);
or U3125 (N_3125,N_418,N_1556);
and U3126 (N_3126,In_3001,N_1577);
nor U3127 (N_3127,N_1541,N_804);
or U3128 (N_3128,N_1273,N_1788);
nor U3129 (N_3129,N_429,N_920);
and U3130 (N_3130,N_1609,N_1088);
xnor U3131 (N_3131,In_2970,In_4537);
nor U3132 (N_3132,In_4694,N_501);
nor U3133 (N_3133,In_2728,N_1905);
xor U3134 (N_3134,In_3447,N_1141);
nor U3135 (N_3135,N_1520,N_151);
nor U3136 (N_3136,In_1114,N_135);
and U3137 (N_3137,N_1906,N_1043);
nor U3138 (N_3138,N_292,In_3506);
and U3139 (N_3139,N_1902,N_220);
nor U3140 (N_3140,N_740,N_1448);
and U3141 (N_3141,N_927,N_1433);
nor U3142 (N_3142,In_841,In_1690);
or U3143 (N_3143,N_1329,N_1873);
or U3144 (N_3144,In_4929,In_1648);
nor U3145 (N_3145,N_1494,N_1229);
or U3146 (N_3146,In_2020,N_1649);
xnor U3147 (N_3147,N_538,In_1566);
xor U3148 (N_3148,N_1697,N_955);
and U3149 (N_3149,N_492,In_4121);
nand U3150 (N_3150,In_4320,In_435);
nor U3151 (N_3151,N_124,N_86);
and U3152 (N_3152,N_1342,In_1675);
xor U3153 (N_3153,N_1824,In_4040);
nor U3154 (N_3154,N_1504,In_3022);
xor U3155 (N_3155,N_309,N_206);
and U3156 (N_3156,In_551,In_1811);
and U3157 (N_3157,N_128,In_3123);
and U3158 (N_3158,In_3515,In_1135);
or U3159 (N_3159,N_663,N_956);
nor U3160 (N_3160,N_413,N_69);
and U3161 (N_3161,N_256,In_1531);
nor U3162 (N_3162,N_1010,In_3425);
nand U3163 (N_3163,In_3031,N_1535);
or U3164 (N_3164,N_475,N_781);
and U3165 (N_3165,N_914,N_1646);
and U3166 (N_3166,N_223,N_477);
and U3167 (N_3167,N_1304,N_1310);
or U3168 (N_3168,N_778,N_1412);
xnor U3169 (N_3169,In_4257,N_972);
xor U3170 (N_3170,N_65,N_1864);
and U3171 (N_3171,N_518,N_1703);
and U3172 (N_3172,N_1390,N_466);
and U3173 (N_3173,In_550,In_2792);
or U3174 (N_3174,N_1533,N_313);
nand U3175 (N_3175,N_850,N_861);
or U3176 (N_3176,N_524,N_1373);
nand U3177 (N_3177,N_647,N_996);
or U3178 (N_3178,In_4457,In_4563);
nand U3179 (N_3179,In_625,In_4570);
or U3180 (N_3180,In_3246,In_2647);
and U3181 (N_3181,N_427,N_480);
nor U3182 (N_3182,N_104,N_15);
xnor U3183 (N_3183,N_1497,N_944);
nand U3184 (N_3184,In_3767,N_1436);
nand U3185 (N_3185,In_1439,N_754);
nand U3186 (N_3186,In_1750,N_813);
nand U3187 (N_3187,N_853,N_232);
and U3188 (N_3188,In_3137,N_1911);
or U3189 (N_3189,N_654,N_751);
and U3190 (N_3190,In_3917,N_214);
or U3191 (N_3191,In_161,In_356);
and U3192 (N_3192,In_1069,N_1144);
nand U3193 (N_3193,N_557,In_378);
nor U3194 (N_3194,N_1012,In_649);
or U3195 (N_3195,N_1561,N_1346);
and U3196 (N_3196,In_4863,N_114);
nand U3197 (N_3197,N_1083,N_1795);
nand U3198 (N_3198,In_4419,In_52);
and U3199 (N_3199,N_1460,N_1014);
nand U3200 (N_3200,In_1212,N_1179);
nand U3201 (N_3201,N_1190,N_612);
and U3202 (N_3202,N_167,N_105);
and U3203 (N_3203,N_1106,N_1248);
and U3204 (N_3204,N_1937,N_1547);
or U3205 (N_3205,N_279,In_3019);
xnor U3206 (N_3206,N_1994,N_1655);
nor U3207 (N_3207,N_1186,N_1275);
and U3208 (N_3208,N_1772,In_1670);
or U3209 (N_3209,N_78,In_4145);
nand U3210 (N_3210,In_2916,In_4628);
xor U3211 (N_3211,N_703,In_4786);
or U3212 (N_3212,In_2314,N_785);
and U3213 (N_3213,In_2809,N_1327);
and U3214 (N_3214,In_3601,N_691);
and U3215 (N_3215,In_2559,N_218);
or U3216 (N_3216,N_500,N_1860);
xnor U3217 (N_3217,In_4506,N_2);
xor U3218 (N_3218,N_94,N_1143);
and U3219 (N_3219,In_1185,N_1130);
xor U3220 (N_3220,In_1662,N_545);
or U3221 (N_3221,N_1033,N_878);
nor U3222 (N_3222,N_1240,In_2131);
and U3223 (N_3223,In_4296,In_16);
xor U3224 (N_3224,N_1093,N_319);
or U3225 (N_3225,N_76,In_943);
nand U3226 (N_3226,N_1813,N_152);
and U3227 (N_3227,N_1623,In_1976);
xor U3228 (N_3228,N_1019,N_1880);
and U3229 (N_3229,In_2671,In_1354);
nand U3230 (N_3230,In_2204,N_1965);
and U3231 (N_3231,N_1558,N_625);
and U3232 (N_3232,In_1087,N_511);
xor U3233 (N_3233,N_1324,In_3887);
nand U3234 (N_3234,In_3635,N_1211);
nor U3235 (N_3235,In_4377,N_1309);
or U3236 (N_3236,N_1046,N_338);
and U3237 (N_3237,N_1802,N_1395);
xnor U3238 (N_3238,N_441,N_417);
nand U3239 (N_3239,N_601,N_940);
nor U3240 (N_3240,N_38,N_1148);
nor U3241 (N_3241,In_878,N_186);
and U3242 (N_3242,N_176,N_1454);
nor U3243 (N_3243,N_1100,N_346);
nand U3244 (N_3244,N_240,N_1050);
xor U3245 (N_3245,N_709,N_817);
or U3246 (N_3246,N_455,In_411);
xnor U3247 (N_3247,N_9,N_396);
nor U3248 (N_3248,N_961,N_869);
nand U3249 (N_3249,N_1630,In_500);
or U3250 (N_3250,N_239,N_744);
and U3251 (N_3251,In_2450,In_3791);
nand U3252 (N_3252,N_951,In_21);
and U3253 (N_3253,In_4989,N_328);
or U3254 (N_3254,N_366,N_1884);
or U3255 (N_3255,N_1241,N_589);
nand U3256 (N_3256,N_1692,N_1298);
xnor U3257 (N_3257,In_1055,N_1861);
nor U3258 (N_3258,N_1234,N_1108);
or U3259 (N_3259,N_1743,In_606);
nand U3260 (N_3260,N_973,N_1553);
nor U3261 (N_3261,In_2999,N_963);
nand U3262 (N_3262,In_1567,In_859);
nand U3263 (N_3263,N_494,N_685);
nor U3264 (N_3264,N_1651,N_596);
or U3265 (N_3265,In_4819,In_3929);
or U3266 (N_3266,N_1053,In_3180);
nand U3267 (N_3267,N_361,In_196);
or U3268 (N_3268,N_488,N_1213);
nand U3269 (N_3269,In_1487,N_1568);
nor U3270 (N_3270,N_921,N_558);
nor U3271 (N_3271,In_1431,N_992);
nor U3272 (N_3272,In_3789,N_1828);
or U3273 (N_3273,In_3756,N_1223);
or U3274 (N_3274,N_37,N_989);
or U3275 (N_3275,N_1918,In_1233);
xnor U3276 (N_3276,In_2845,In_4579);
xor U3277 (N_3277,In_4590,N_997);
nand U3278 (N_3278,In_90,In_2674);
and U3279 (N_3279,In_870,N_1843);
nor U3280 (N_3280,N_913,N_1388);
xnor U3281 (N_3281,N_745,N_1459);
nand U3282 (N_3282,N_1971,N_68);
or U3283 (N_3283,In_1033,N_39);
or U3284 (N_3284,In_3233,N_352);
xor U3285 (N_3285,In_4574,N_409);
and U3286 (N_3286,N_1531,In_3577);
xor U3287 (N_3287,In_3268,N_1967);
nor U3288 (N_3288,In_4808,In_2566);
xnor U3289 (N_3289,In_4610,In_1307);
and U3290 (N_3290,In_1659,In_407);
nand U3291 (N_3291,N_1842,In_160);
or U3292 (N_3292,N_977,In_3457);
or U3293 (N_3293,In_2472,In_3060);
and U3294 (N_3294,N_1810,N_1008);
xor U3295 (N_3295,In_4987,N_892);
or U3296 (N_3296,N_146,N_801);
nor U3297 (N_3297,In_1654,N_300);
nand U3298 (N_3298,N_1786,N_1681);
and U3299 (N_3299,N_282,In_3931);
nor U3300 (N_3300,In_2060,N_1020);
nor U3301 (N_3301,In_632,In_4932);
nor U3302 (N_3302,N_100,N_537);
nand U3303 (N_3303,N_58,In_1892);
nor U3304 (N_3304,N_822,N_1816);
and U3305 (N_3305,In_3699,N_1845);
or U3306 (N_3306,N_1221,N_374);
nand U3307 (N_3307,N_233,In_1643);
xor U3308 (N_3308,N_884,N_1196);
xor U3309 (N_3309,In_2940,N_1785);
nand U3310 (N_3310,N_154,In_3618);
xnor U3311 (N_3311,N_1103,In_3751);
nand U3312 (N_3312,N_1055,In_2702);
xnor U3313 (N_3313,N_797,N_504);
xnor U3314 (N_3314,N_1830,N_610);
nor U3315 (N_3315,N_1146,In_952);
xor U3316 (N_3316,In_3407,In_856);
xnor U3317 (N_3317,N_1303,N_281);
xor U3318 (N_3318,N_1849,N_600);
xor U3319 (N_3319,N_1970,N_641);
xor U3320 (N_3320,N_936,In_2126);
nand U3321 (N_3321,N_60,N_1798);
nor U3322 (N_3322,N_667,N_1879);
nand U3323 (N_3323,In_170,N_758);
and U3324 (N_3324,In_4634,N_826);
xnor U3325 (N_3325,In_3215,In_4420);
xnor U3326 (N_3326,In_4184,N_645);
nor U3327 (N_3327,N_33,N_244);
xnor U3328 (N_3328,N_269,N_1051);
nand U3329 (N_3329,N_1974,N_1246);
or U3330 (N_3330,In_3964,N_1943);
and U3331 (N_3331,In_2479,N_1426);
or U3332 (N_3332,N_1886,N_1251);
nand U3333 (N_3333,N_766,N_84);
nand U3334 (N_3334,In_662,N_1923);
nor U3335 (N_3335,N_1037,N_1988);
xor U3336 (N_3336,In_687,N_412);
nor U3337 (N_3337,In_3442,N_1793);
or U3338 (N_3338,N_1363,In_2877);
xnor U3339 (N_3339,N_926,In_4673);
nor U3340 (N_3340,N_1660,N_1109);
and U3341 (N_3341,N_621,In_3673);
nor U3342 (N_3342,N_979,N_210);
or U3343 (N_3343,N_1762,N_1769);
and U3344 (N_3344,N_1749,N_353);
xnor U3345 (N_3345,N_1291,N_1177);
and U3346 (N_3346,N_1929,In_3516);
nand U3347 (N_3347,In_1686,N_1028);
xnor U3348 (N_3348,In_3565,N_1503);
and U3349 (N_3349,N_1382,In_4917);
and U3350 (N_3350,In_298,N_1468);
xnor U3351 (N_3351,N_194,In_1421);
and U3352 (N_3352,In_451,N_1803);
xnor U3353 (N_3353,In_2554,N_1011);
or U3354 (N_3354,N_509,In_4217);
nand U3355 (N_3355,N_1261,In_53);
and U3356 (N_3356,N_407,In_4985);
xor U3357 (N_3357,N_1475,N_172);
xor U3358 (N_3358,N_445,In_433);
nor U3359 (N_3359,In_2885,In_4594);
and U3360 (N_3360,N_520,N_1664);
nand U3361 (N_3361,N_790,N_340);
xor U3362 (N_3362,In_3139,N_848);
nor U3363 (N_3363,In_95,N_874);
nor U3364 (N_3364,N_34,In_4423);
nand U3365 (N_3365,N_1378,In_1640);
nand U3366 (N_3366,N_264,N_1428);
nor U3367 (N_3367,In_1329,In_456);
or U3368 (N_3368,N_1985,N_893);
xor U3369 (N_3369,N_712,In_3144);
xnor U3370 (N_3370,In_4639,In_3993);
nand U3371 (N_3371,N_1375,In_1164);
and U3372 (N_3372,In_4179,N_196);
nor U3373 (N_3373,In_2147,N_701);
xor U3374 (N_3374,N_865,N_776);
xnor U3375 (N_3375,N_77,N_1825);
and U3376 (N_3376,N_540,N_1932);
or U3377 (N_3377,In_795,N_362);
and U3378 (N_3378,N_586,N_1445);
or U3379 (N_3379,N_1379,N_145);
nand U3380 (N_3380,N_1222,N_950);
xnor U3381 (N_3381,N_1381,N_1401);
and U3382 (N_3382,In_2072,N_572);
nor U3383 (N_3383,N_157,N_519);
nor U3384 (N_3384,N_933,N_594);
nor U3385 (N_3385,In_3639,N_1776);
and U3386 (N_3386,N_1628,In_4143);
or U3387 (N_3387,N_525,N_470);
nor U3388 (N_3388,In_1489,In_4815);
xnor U3389 (N_3389,In_66,N_1127);
xnor U3390 (N_3390,In_3759,N_881);
and U3391 (N_3391,N_1542,N_948);
xnor U3392 (N_3392,N_234,N_434);
or U3393 (N_3393,N_640,N_213);
nor U3394 (N_3394,N_532,N_1624);
xor U3395 (N_3395,In_2783,N_1256);
and U3396 (N_3396,In_4210,In_2104);
and U3397 (N_3397,N_1526,N_1866);
xor U3398 (N_3398,In_1930,In_1075);
and U3399 (N_3399,N_1457,N_1131);
xnor U3400 (N_3400,In_1928,N_347);
or U3401 (N_3401,N_1983,N_127);
and U3402 (N_3402,In_4479,In_4149);
nor U3403 (N_3403,In_3543,In_4840);
and U3404 (N_3404,N_1684,N_473);
xor U3405 (N_3405,N_1057,N_1397);
nor U3406 (N_3406,N_1341,N_1272);
or U3407 (N_3407,N_1868,N_1958);
or U3408 (N_3408,N_21,In_336);
xnor U3409 (N_3409,N_1777,N_880);
nand U3410 (N_3410,N_1814,In_2706);
xor U3411 (N_3411,N_343,N_1564);
and U3412 (N_3412,N_852,In_51);
nor U3413 (N_3413,In_2480,In_605);
nor U3414 (N_3414,N_1238,N_606);
nand U3415 (N_3415,N_590,N_729);
and U3416 (N_3416,N_575,N_791);
or U3417 (N_3417,In_2775,N_91);
xor U3418 (N_3418,N_698,N_1548);
xnor U3419 (N_3419,In_279,In_193);
xor U3420 (N_3420,In_2381,N_99);
and U3421 (N_3421,N_415,In_1442);
nor U3422 (N_3422,N_889,In_4977);
nand U3423 (N_3423,In_3157,N_198);
xnor U3424 (N_3424,In_1666,N_1400);
nor U3425 (N_3425,In_1243,N_442);
nor U3426 (N_3426,N_1763,N_1096);
nor U3427 (N_3427,In_1499,In_1086);
nor U3428 (N_3428,N_379,N_291);
nor U3429 (N_3429,N_288,N_1595);
xnor U3430 (N_3430,N_1171,N_1305);
and U3431 (N_3431,N_1406,N_1606);
nor U3432 (N_3432,N_1839,N_686);
nand U3433 (N_3433,N_64,N_1909);
nand U3434 (N_3434,N_1947,In_4528);
nor U3435 (N_3435,N_332,N_528);
or U3436 (N_3436,In_2001,In_4246);
and U3437 (N_3437,N_1371,In_3607);
and U3438 (N_3438,N_1570,N_1597);
and U3439 (N_3439,In_3336,N_1620);
xnor U3440 (N_3440,N_465,In_4491);
nor U3441 (N_3441,In_3946,N_1924);
or U3442 (N_3442,N_1908,N_1696);
xor U3443 (N_3443,N_1102,N_13);
xnor U3444 (N_3444,In_1688,N_1334);
nor U3445 (N_3445,N_136,In_2024);
nand U3446 (N_3446,In_3196,N_1359);
and U3447 (N_3447,N_1716,N_1850);
or U3448 (N_3448,N_274,N_593);
and U3449 (N_3449,In_3773,N_1835);
or U3450 (N_3450,In_2905,N_1182);
and U3451 (N_3451,N_181,N_1904);
xnor U3452 (N_3452,In_4319,In_3420);
nand U3453 (N_3453,N_1134,In_4498);
xnor U3454 (N_3454,N_1907,In_1029);
or U3455 (N_3455,In_3799,N_1336);
xor U3456 (N_3456,In_3349,N_66);
nand U3457 (N_3457,N_1482,In_202);
or U3458 (N_3458,N_1731,N_945);
and U3459 (N_3459,N_296,In_4015);
nand U3460 (N_3460,N_1894,N_457);
xor U3461 (N_3461,N_416,N_664);
or U3462 (N_3462,N_1153,N_793);
and U3463 (N_3463,N_1077,N_1350);
nand U3464 (N_3464,In_3109,In_4738);
xnor U3465 (N_3465,N_467,N_1870);
nor U3466 (N_3466,N_1450,N_59);
xor U3467 (N_3467,N_1534,N_1465);
and U3468 (N_3468,In_1514,In_3291);
nand U3469 (N_3469,In_4588,In_2425);
or U3470 (N_3470,N_717,N_1779);
and U3471 (N_3471,In_2323,N_1536);
or U3472 (N_3472,N_103,N_1389);
nand U3473 (N_3473,In_4997,N_1571);
and U3474 (N_3474,In_2878,N_503);
xor U3475 (N_3475,N_1836,N_1485);
nor U3476 (N_3476,N_459,N_1783);
or U3477 (N_3477,N_986,N_472);
or U3478 (N_3478,N_1257,N_1048);
and U3479 (N_3479,N_734,In_3045);
xor U3480 (N_3480,In_4357,N_1383);
xor U3481 (N_3481,N_1183,N_1969);
nand U3482 (N_3482,N_158,In_3089);
and U3483 (N_3483,In_2570,N_1940);
nor U3484 (N_3484,In_4516,In_2822);
nand U3485 (N_3485,In_4348,N_1084);
or U3486 (N_3486,N_732,N_192);
and U3487 (N_3487,N_1340,N_1695);
xor U3488 (N_3488,N_1004,In_1731);
nand U3489 (N_3489,In_54,N_1888);
xor U3490 (N_3490,N_1647,In_3735);
nor U3491 (N_3491,N_1282,In_774);
or U3492 (N_3492,N_1142,In_2191);
nor U3493 (N_3493,In_152,In_2370);
xnor U3494 (N_3494,N_499,N_1337);
nor U3495 (N_3495,N_1652,N_71);
xnor U3496 (N_3496,In_4311,N_910);
nor U3497 (N_3497,In_171,N_626);
nand U3498 (N_3498,N_1,N_1289);
or U3499 (N_3499,In_530,In_842);
and U3500 (N_3500,N_1803,In_3655);
nor U3501 (N_3501,In_2775,N_1832);
xnor U3502 (N_3502,In_3233,In_3045);
nor U3503 (N_3503,N_1660,N_1689);
or U3504 (N_3504,N_603,In_1696);
and U3505 (N_3505,N_430,In_2593);
nor U3506 (N_3506,In_3724,In_4033);
nand U3507 (N_3507,N_1535,N_827);
xnor U3508 (N_3508,In_3098,N_1619);
xnor U3509 (N_3509,In_90,N_1843);
or U3510 (N_3510,N_1876,In_1445);
nor U3511 (N_3511,N_1522,N_511);
xnor U3512 (N_3512,N_939,In_697);
and U3513 (N_3513,N_573,N_138);
or U3514 (N_3514,N_1562,In_682);
nand U3515 (N_3515,N_1912,N_427);
or U3516 (N_3516,In_118,N_1542);
xor U3517 (N_3517,In_4928,N_136);
nand U3518 (N_3518,N_1297,In_1675);
or U3519 (N_3519,N_402,N_1090);
nand U3520 (N_3520,N_1675,N_1696);
and U3521 (N_3521,N_181,N_1902);
nor U3522 (N_3522,N_478,N_168);
and U3523 (N_3523,In_2906,N_1946);
and U3524 (N_3524,N_346,In_2775);
nor U3525 (N_3525,N_375,In_1892);
and U3526 (N_3526,N_323,In_990);
and U3527 (N_3527,In_1630,In_4287);
or U3528 (N_3528,N_1709,In_1666);
nor U3529 (N_3529,N_1260,N_502);
nor U3530 (N_3530,N_216,In_4660);
and U3531 (N_3531,N_1323,In_3964);
nor U3532 (N_3532,N_408,N_1607);
xor U3533 (N_3533,N_420,N_1436);
xor U3534 (N_3534,N_1259,N_1780);
and U3535 (N_3535,N_1827,N_1466);
nand U3536 (N_3536,N_804,In_3898);
nand U3537 (N_3537,N_1012,In_4586);
nor U3538 (N_3538,In_4257,N_1649);
xor U3539 (N_3539,N_427,In_2706);
and U3540 (N_3540,In_21,In_4033);
nand U3541 (N_3541,In_2347,N_1455);
or U3542 (N_3542,N_1355,In_4989);
nor U3543 (N_3543,N_930,N_822);
xor U3544 (N_3544,In_2223,N_926);
nand U3545 (N_3545,N_1230,In_741);
nor U3546 (N_3546,In_380,In_137);
nand U3547 (N_3547,N_1921,In_2857);
xor U3548 (N_3548,N_246,In_90);
and U3549 (N_3549,N_1568,N_455);
nor U3550 (N_3550,In_1784,N_238);
and U3551 (N_3551,In_1408,In_1930);
nor U3552 (N_3552,In_1855,In_213);
and U3553 (N_3553,N_356,N_1158);
and U3554 (N_3554,N_417,N_206);
nand U3555 (N_3555,N_871,N_1810);
nor U3556 (N_3556,N_967,N_410);
and U3557 (N_3557,N_1323,In_356);
xnor U3558 (N_3558,In_1688,In_4787);
nor U3559 (N_3559,N_1584,N_664);
nand U3560 (N_3560,In_2647,N_1173);
nand U3561 (N_3561,N_694,In_1080);
nor U3562 (N_3562,N_1774,N_1898);
xnor U3563 (N_3563,N_1815,N_1687);
nor U3564 (N_3564,In_1711,N_1483);
xor U3565 (N_3565,N_910,N_569);
nor U3566 (N_3566,In_3019,N_705);
or U3567 (N_3567,N_447,N_1638);
nor U3568 (N_3568,In_1308,N_725);
xnor U3569 (N_3569,In_2144,N_1063);
nand U3570 (N_3570,In_3534,N_256);
xor U3571 (N_3571,N_1754,In_2204);
and U3572 (N_3572,In_1564,In_1760);
nor U3573 (N_3573,In_442,In_1636);
or U3574 (N_3574,In_4662,N_1916);
xor U3575 (N_3575,N_1142,N_1256);
nand U3576 (N_3576,N_397,In_659);
and U3577 (N_3577,N_558,N_829);
and U3578 (N_3578,N_994,N_1186);
nor U3579 (N_3579,N_266,In_2916);
nor U3580 (N_3580,In_419,N_1403);
or U3581 (N_3581,N_1758,N_246);
or U3582 (N_3582,N_1291,N_353);
nor U3583 (N_3583,N_762,N_1724);
nand U3584 (N_3584,In_4531,N_1318);
nor U3585 (N_3585,In_4825,In_869);
or U3586 (N_3586,N_968,N_1396);
nand U3587 (N_3587,N_70,N_1255);
nor U3588 (N_3588,N_1036,In_508);
xnor U3589 (N_3589,N_151,In_625);
xnor U3590 (N_3590,In_2907,N_80);
nand U3591 (N_3591,N_219,N_826);
or U3592 (N_3592,N_1460,N_1483);
and U3593 (N_3593,N_259,N_1681);
or U3594 (N_3594,N_902,N_944);
and U3595 (N_3595,In_4840,In_1033);
xor U3596 (N_3596,N_209,N_1501);
nor U3597 (N_3597,N_283,In_346);
nand U3598 (N_3598,In_1086,N_432);
nor U3599 (N_3599,N_805,N_123);
nand U3600 (N_3600,N_1490,N_1334);
nand U3601 (N_3601,N_1707,N_260);
nor U3602 (N_3602,In_2444,N_1174);
nand U3603 (N_3603,N_784,N_1474);
nand U3604 (N_3604,N_357,N_909);
or U3605 (N_3605,N_1922,N_1039);
and U3606 (N_3606,N_401,In_3791);
and U3607 (N_3607,In_251,In_3091);
and U3608 (N_3608,In_1523,N_1933);
or U3609 (N_3609,N_343,In_856);
nor U3610 (N_3610,In_4172,N_1289);
and U3611 (N_3611,N_4,In_4296);
nand U3612 (N_3612,N_1349,In_170);
or U3613 (N_3613,N_1456,N_858);
or U3614 (N_3614,N_498,N_218);
nor U3615 (N_3615,In_1496,In_3157);
nand U3616 (N_3616,N_1595,N_1857);
xnor U3617 (N_3617,N_195,N_1553);
or U3618 (N_3618,N_1648,In_4807);
nor U3619 (N_3619,In_3792,N_1955);
and U3620 (N_3620,N_1487,In_3457);
nor U3621 (N_3621,N_1163,In_3789);
xor U3622 (N_3622,In_2438,N_279);
xor U3623 (N_3623,N_630,In_69);
xnor U3624 (N_3624,N_1811,N_897);
and U3625 (N_3625,In_550,N_1810);
nor U3626 (N_3626,N_1299,In_550);
nor U3627 (N_3627,In_795,In_1908);
nor U3628 (N_3628,In_1012,N_1324);
xor U3629 (N_3629,N_1272,N_1474);
nand U3630 (N_3630,In_21,In_4119);
nand U3631 (N_3631,N_1951,N_246);
nand U3632 (N_3632,N_1981,N_1666);
nor U3633 (N_3633,N_660,In_11);
nor U3634 (N_3634,In_1567,In_2905);
nor U3635 (N_3635,N_863,In_618);
nand U3636 (N_3636,N_1286,In_2736);
or U3637 (N_3637,In_3379,N_1044);
and U3638 (N_3638,N_1324,N_1202);
nand U3639 (N_3639,In_4605,In_1439);
nor U3640 (N_3640,N_136,N_118);
or U3641 (N_3641,In_625,N_1941);
xnor U3642 (N_3642,N_14,In_625);
or U3643 (N_3643,N_730,N_1048);
and U3644 (N_3644,N_557,In_3695);
xor U3645 (N_3645,N_703,N_1500);
xor U3646 (N_3646,N_1288,N_469);
or U3647 (N_3647,N_880,N_713);
and U3648 (N_3648,In_4223,N_834);
xor U3649 (N_3649,In_3521,N_1070);
and U3650 (N_3650,N_1359,N_1691);
nor U3651 (N_3651,N_1986,N_918);
xnor U3652 (N_3652,N_197,In_167);
and U3653 (N_3653,N_1085,N_445);
nor U3654 (N_3654,In_659,In_1622);
nor U3655 (N_3655,N_1053,N_690);
and U3656 (N_3656,N_714,N_675);
xnor U3657 (N_3657,N_949,N_989);
and U3658 (N_3658,In_4103,N_1508);
xnor U3659 (N_3659,In_3651,In_3355);
and U3660 (N_3660,N_203,N_931);
nand U3661 (N_3661,N_1776,N_1428);
xor U3662 (N_3662,N_1046,N_686);
or U3663 (N_3663,In_4783,N_1866);
nor U3664 (N_3664,N_471,In_1572);
and U3665 (N_3665,N_444,In_3166);
nor U3666 (N_3666,N_126,N_268);
and U3667 (N_3667,N_1284,N_729);
or U3668 (N_3668,N_337,In_4985);
or U3669 (N_3669,In_4503,N_860);
xor U3670 (N_3670,N_1491,N_808);
nor U3671 (N_3671,N_47,N_518);
nand U3672 (N_3672,In_3502,N_122);
nand U3673 (N_3673,In_3248,N_625);
xnor U3674 (N_3674,N_347,In_2845);
and U3675 (N_3675,In_2164,N_606);
nand U3676 (N_3676,N_1430,In_4985);
xor U3677 (N_3677,N_1843,In_4409);
xnor U3678 (N_3678,In_3212,In_3759);
and U3679 (N_3679,N_351,In_324);
and U3680 (N_3680,N_820,N_664);
or U3681 (N_3681,N_342,N_428);
nor U3682 (N_3682,N_1313,N_1560);
xnor U3683 (N_3683,In_1219,N_1247);
and U3684 (N_3684,N_341,N_546);
and U3685 (N_3685,In_3534,N_1569);
and U3686 (N_3686,N_678,In_435);
xnor U3687 (N_3687,In_2935,In_4703);
and U3688 (N_3688,N_1838,In_1229);
nand U3689 (N_3689,In_1398,N_1401);
and U3690 (N_3690,N_1720,N_1270);
nand U3691 (N_3691,N_1270,N_1575);
xnor U3692 (N_3692,N_896,N_1844);
nor U3693 (N_3693,N_595,N_1149);
and U3694 (N_3694,In_3220,N_1855);
and U3695 (N_3695,N_611,N_1454);
nand U3696 (N_3696,N_817,N_117);
and U3697 (N_3697,In_2603,In_3183);
and U3698 (N_3698,N_774,N_1655);
nor U3699 (N_3699,N_1934,N_1997);
nand U3700 (N_3700,N_681,N_879);
or U3701 (N_3701,N_1211,In_2438);
or U3702 (N_3702,N_1704,N_1148);
nor U3703 (N_3703,N_175,N_819);
nor U3704 (N_3704,N_1986,N_1189);
nor U3705 (N_3705,N_1622,N_1771);
nand U3706 (N_3706,N_1255,N_1978);
and U3707 (N_3707,N_129,N_1447);
or U3708 (N_3708,In_1922,In_1164);
nor U3709 (N_3709,In_4841,N_986);
or U3710 (N_3710,N_657,N_1024);
and U3711 (N_3711,In_767,N_1959);
and U3712 (N_3712,N_1354,N_205);
and U3713 (N_3713,N_1446,N_386);
nor U3714 (N_3714,In_985,N_1559);
and U3715 (N_3715,N_1973,In_3693);
xnor U3716 (N_3716,N_1047,N_1195);
nand U3717 (N_3717,N_1355,In_745);
and U3718 (N_3718,In_2213,N_357);
and U3719 (N_3719,N_205,N_1133);
nor U3720 (N_3720,N_1369,N_1460);
nor U3721 (N_3721,In_994,N_517);
or U3722 (N_3722,N_506,N_425);
nand U3723 (N_3723,N_1693,N_549);
nor U3724 (N_3724,N_840,N_1902);
or U3725 (N_3725,N_692,N_1408);
or U3726 (N_3726,In_4479,N_212);
nor U3727 (N_3727,In_3904,In_1248);
nand U3728 (N_3728,In_2728,In_2970);
and U3729 (N_3729,N_1649,N_1791);
nor U3730 (N_3730,N_189,N_1912);
and U3731 (N_3731,N_1079,In_4197);
and U3732 (N_3732,In_4521,N_656);
nor U3733 (N_3733,N_1048,N_662);
nor U3734 (N_3734,N_518,N_1985);
xnor U3735 (N_3735,N_1808,N_352);
xnor U3736 (N_3736,In_3233,N_1781);
xor U3737 (N_3737,In_2431,N_630);
nor U3738 (N_3738,In_3946,In_4673);
and U3739 (N_3739,N_1095,In_36);
or U3740 (N_3740,In_3425,N_858);
xor U3741 (N_3741,In_1446,N_1216);
or U3742 (N_3742,In_496,N_593);
xor U3743 (N_3743,N_668,N_356);
or U3744 (N_3744,N_1484,N_933);
nor U3745 (N_3745,N_148,In_3146);
xor U3746 (N_3746,N_894,N_830);
or U3747 (N_3747,In_2935,N_1410);
xnor U3748 (N_3748,N_671,N_1592);
and U3749 (N_3749,In_1243,In_2970);
and U3750 (N_3750,N_764,N_630);
or U3751 (N_3751,In_2728,N_512);
nor U3752 (N_3752,In_336,N_871);
nor U3753 (N_3753,N_588,N_1409);
nor U3754 (N_3754,N_830,N_1465);
and U3755 (N_3755,N_1523,N_1163);
and U3756 (N_3756,N_908,N_36);
nand U3757 (N_3757,N_159,N_1342);
xnor U3758 (N_3758,In_2178,N_1401);
and U3759 (N_3759,N_316,N_1945);
and U3760 (N_3760,N_208,N_1692);
and U3761 (N_3761,N_1452,N_752);
xnor U3762 (N_3762,N_1348,N_486);
xnor U3763 (N_3763,N_1224,N_698);
or U3764 (N_3764,N_434,N_1469);
xor U3765 (N_3765,N_1085,N_592);
and U3766 (N_3766,In_4673,N_540);
xor U3767 (N_3767,N_1179,N_418);
and U3768 (N_3768,N_837,N_1314);
and U3769 (N_3769,In_3176,N_1900);
or U3770 (N_3770,In_632,N_757);
nand U3771 (N_3771,In_3645,In_3979);
nand U3772 (N_3772,N_218,N_2);
nor U3773 (N_3773,N_1995,N_1349);
nor U3774 (N_3774,N_1162,N_1266);
xnor U3775 (N_3775,N_703,N_377);
nor U3776 (N_3776,N_1417,In_1686);
nand U3777 (N_3777,In_2617,N_1582);
xor U3778 (N_3778,In_2638,In_3272);
xor U3779 (N_3779,In_1382,N_389);
xnor U3780 (N_3780,In_739,In_3974);
nand U3781 (N_3781,N_1920,In_3048);
and U3782 (N_3782,N_284,N_1435);
and U3783 (N_3783,In_2666,In_2523);
xnor U3784 (N_3784,In_1654,In_3929);
nand U3785 (N_3785,In_3708,N_1607);
nand U3786 (N_3786,In_4926,In_3055);
nor U3787 (N_3787,N_1328,N_794);
or U3788 (N_3788,N_511,N_1584);
and U3789 (N_3789,N_906,N_513);
nand U3790 (N_3790,N_164,N_1798);
nor U3791 (N_3791,In_631,In_4634);
nor U3792 (N_3792,In_3157,N_1910);
xor U3793 (N_3793,N_1149,N_1091);
or U3794 (N_3794,N_560,N_1343);
and U3795 (N_3795,N_1684,N_178);
and U3796 (N_3796,N_951,N_885);
xnor U3797 (N_3797,N_1736,N_1791);
nor U3798 (N_3798,N_1814,In_2022);
and U3799 (N_3799,In_3261,N_1879);
and U3800 (N_3800,N_290,In_1228);
nand U3801 (N_3801,N_1751,N_1811);
nand U3802 (N_3802,N_127,N_1177);
nor U3803 (N_3803,N_1214,N_1129);
nor U3804 (N_3804,N_388,N_682);
and U3805 (N_3805,N_514,N_194);
nor U3806 (N_3806,In_465,N_1992);
and U3807 (N_3807,N_1006,N_169);
nor U3808 (N_3808,N_1914,In_4490);
nor U3809 (N_3809,N_468,N_392);
or U3810 (N_3810,N_908,N_595);
xor U3811 (N_3811,N_929,N_287);
or U3812 (N_3812,In_497,N_1014);
nand U3813 (N_3813,In_4985,In_2905);
and U3814 (N_3814,N_430,In_4119);
nor U3815 (N_3815,N_1291,N_878);
nor U3816 (N_3816,In_3198,N_971);
xor U3817 (N_3817,N_201,N_774);
or U3818 (N_3818,In_777,In_1649);
nor U3819 (N_3819,N_1954,N_1666);
xnor U3820 (N_3820,N_553,In_51);
xor U3821 (N_3821,In_3123,N_1479);
or U3822 (N_3822,N_1998,N_1297);
and U3823 (N_3823,In_431,N_50);
nand U3824 (N_3824,N_205,N_721);
xnor U3825 (N_3825,N_1927,N_893);
and U3826 (N_3826,In_531,N_287);
nor U3827 (N_3827,In_411,In_2559);
or U3828 (N_3828,In_133,In_3279);
xnor U3829 (N_3829,N_1048,In_1566);
xor U3830 (N_3830,N_1142,N_56);
xnor U3831 (N_3831,N_148,N_1575);
or U3832 (N_3832,N_1085,N_1748);
or U3833 (N_3833,N_1064,N_110);
and U3834 (N_3834,N_1761,In_2559);
xnor U3835 (N_3835,N_1828,In_2018);
nand U3836 (N_3836,In_4457,N_389);
or U3837 (N_3837,N_209,In_4213);
and U3838 (N_3838,N_925,N_453);
nor U3839 (N_3839,In_3886,N_745);
and U3840 (N_3840,In_1596,In_1148);
nand U3841 (N_3841,N_994,N_197);
or U3842 (N_3842,In_175,In_1159);
nand U3843 (N_3843,N_1421,N_743);
and U3844 (N_3844,In_1309,In_2104);
nor U3845 (N_3845,In_4145,N_1348);
or U3846 (N_3846,N_383,In_3415);
and U3847 (N_3847,In_3726,N_1460);
nor U3848 (N_3848,N_1174,N_692);
or U3849 (N_3849,N_909,In_4457);
xor U3850 (N_3850,N_833,In_1211);
nand U3851 (N_3851,In_1689,N_1767);
xor U3852 (N_3852,N_147,N_1517);
nor U3853 (N_3853,N_1500,In_2390);
and U3854 (N_3854,N_813,N_181);
or U3855 (N_3855,In_3269,N_1523);
and U3856 (N_3856,N_1890,In_1452);
nand U3857 (N_3857,N_1545,N_1243);
or U3858 (N_3858,N_1187,N_866);
xnor U3859 (N_3859,N_854,In_582);
nand U3860 (N_3860,N_1001,N_269);
xnor U3861 (N_3861,N_1123,N_1646);
xor U3862 (N_3862,In_2736,N_256);
or U3863 (N_3863,N_1535,In_1220);
nor U3864 (N_3864,In_3210,N_1291);
xor U3865 (N_3865,N_37,N_1797);
nand U3866 (N_3866,N_1935,N_1617);
xnor U3867 (N_3867,N_1183,N_397);
nor U3868 (N_3868,In_4040,N_931);
xnor U3869 (N_3869,N_57,In_2297);
and U3870 (N_3870,N_1202,N_1471);
and U3871 (N_3871,N_1703,N_627);
and U3872 (N_3872,N_941,In_192);
nor U3873 (N_3873,In_3914,N_851);
nor U3874 (N_3874,N_1009,In_2830);
and U3875 (N_3875,N_1566,N_613);
nor U3876 (N_3876,N_894,In_1690);
nor U3877 (N_3877,N_1911,In_4594);
xnor U3878 (N_3878,N_389,N_1108);
nor U3879 (N_3879,N_524,In_3195);
and U3880 (N_3880,N_1194,N_824);
and U3881 (N_3881,N_1175,In_3751);
or U3882 (N_3882,N_1856,N_1939);
and U3883 (N_3883,In_4840,N_496);
nand U3884 (N_3884,N_298,N_24);
nand U3885 (N_3885,In_4162,N_1364);
nor U3886 (N_3886,In_2636,In_2775);
xnor U3887 (N_3887,N_1772,N_1096);
nor U3888 (N_3888,N_632,N_1354);
or U3889 (N_3889,N_1511,In_405);
nor U3890 (N_3890,In_3929,In_4462);
nor U3891 (N_3891,N_837,N_1006);
and U3892 (N_3892,N_1481,N_1703);
and U3893 (N_3893,In_28,N_658);
and U3894 (N_3894,N_53,N_294);
and U3895 (N_3895,In_4240,In_3463);
and U3896 (N_3896,N_1268,N_137);
or U3897 (N_3897,In_1750,N_1063);
nor U3898 (N_3898,N_923,In_1856);
or U3899 (N_3899,N_104,N_1672);
or U3900 (N_3900,N_1459,N_933);
and U3901 (N_3901,N_283,N_1162);
or U3902 (N_3902,N_1442,In_4813);
or U3903 (N_3903,N_1325,N_1371);
nor U3904 (N_3904,N_286,In_4137);
and U3905 (N_3905,N_1130,N_360);
and U3906 (N_3906,In_120,N_1594);
xor U3907 (N_3907,N_1225,N_1200);
or U3908 (N_3908,N_309,In_4917);
and U3909 (N_3909,N_1947,N_1748);
and U3910 (N_3910,In_4105,N_73);
or U3911 (N_3911,N_446,In_1617);
xor U3912 (N_3912,In_3048,N_257);
nand U3913 (N_3913,N_1143,In_3974);
nand U3914 (N_3914,N_2,N_732);
nor U3915 (N_3915,In_1667,N_964);
and U3916 (N_3916,N_1671,N_135);
xnor U3917 (N_3917,N_1311,N_872);
nand U3918 (N_3918,N_440,N_1210);
xor U3919 (N_3919,N_589,In_3767);
or U3920 (N_3920,N_1658,N_1285);
xnor U3921 (N_3921,N_1009,N_1277);
or U3922 (N_3922,N_1027,N_1845);
nor U3923 (N_3923,In_4431,N_210);
xnor U3924 (N_3924,N_1964,N_847);
and U3925 (N_3925,N_1892,N_1124);
and U3926 (N_3926,N_735,N_352);
nor U3927 (N_3927,In_2822,N_1662);
nand U3928 (N_3928,N_70,N_722);
xor U3929 (N_3929,In_508,N_57);
nand U3930 (N_3930,In_3272,N_627);
or U3931 (N_3931,In_3096,N_1963);
nand U3932 (N_3932,In_3060,N_1044);
and U3933 (N_3933,N_1388,N_1076);
or U3934 (N_3934,N_312,In_4419);
nand U3935 (N_3935,N_51,In_1012);
nor U3936 (N_3936,N_379,N_1331);
and U3937 (N_3937,N_1743,N_776);
nor U3938 (N_3938,In_4253,N_1679);
or U3939 (N_3939,N_675,N_1279);
or U3940 (N_3940,In_95,In_4844);
nor U3941 (N_3941,N_963,In_4582);
nor U3942 (N_3942,N_951,In_2655);
or U3943 (N_3943,N_1004,In_1055);
nor U3944 (N_3944,In_3198,N_471);
or U3945 (N_3945,N_457,N_175);
xnor U3946 (N_3946,N_769,N_1862);
xor U3947 (N_3947,N_766,In_741);
nand U3948 (N_3948,N_1611,N_1962);
nand U3949 (N_3949,N_1148,N_1172);
and U3950 (N_3950,N_1079,In_1636);
xnor U3951 (N_3951,N_727,N_1757);
xnor U3952 (N_3952,In_4180,In_3918);
or U3953 (N_3953,N_1552,N_732);
and U3954 (N_3954,In_2936,In_1475);
nor U3955 (N_3955,N_1527,In_3332);
nand U3956 (N_3956,N_809,N_1330);
or U3957 (N_3957,In_4660,In_2191);
xor U3958 (N_3958,N_1196,In_4786);
nand U3959 (N_3959,N_1447,In_4964);
and U3960 (N_3960,N_1162,N_1184);
nor U3961 (N_3961,In_4813,In_1087);
nand U3962 (N_3962,N_98,N_125);
nor U3963 (N_3963,N_1739,N_785);
and U3964 (N_3964,N_297,In_1166);
or U3965 (N_3965,N_1816,N_1616);
and U3966 (N_3966,N_1561,N_444);
and U3967 (N_3967,In_1080,N_899);
or U3968 (N_3968,N_774,N_250);
nand U3969 (N_3969,N_1705,N_712);
nand U3970 (N_3970,In_1489,N_29);
nor U3971 (N_3971,N_1461,N_1088);
and U3972 (N_3972,N_1359,In_4734);
nand U3973 (N_3973,N_184,N_73);
nor U3974 (N_3974,In_4537,In_3019);
and U3975 (N_3975,N_1905,In_827);
xor U3976 (N_3976,N_591,N_1028);
nand U3977 (N_3977,In_51,N_1195);
or U3978 (N_3978,N_29,N_7);
nand U3979 (N_3979,In_1649,N_137);
or U3980 (N_3980,N_1438,N_920);
nand U3981 (N_3981,N_901,N_909);
xor U3982 (N_3982,N_1220,N_1219);
nor U3983 (N_3983,N_61,N_1872);
and U3984 (N_3984,In_3979,N_1264);
or U3985 (N_3985,N_666,N_1334);
nor U3986 (N_3986,In_1135,N_1985);
xor U3987 (N_3987,N_922,In_465);
or U3988 (N_3988,N_839,N_1768);
xnor U3989 (N_3989,N_1458,In_3751);
nand U3990 (N_3990,N_157,N_197);
and U3991 (N_3991,N_1714,In_2755);
nor U3992 (N_3992,N_889,N_1217);
and U3993 (N_3993,N_1627,N_284);
and U3994 (N_3994,N_1777,In_838);
or U3995 (N_3995,N_1413,N_1985);
nand U3996 (N_3996,N_305,N_347);
or U3997 (N_3997,In_3635,N_1541);
and U3998 (N_3998,In_3355,In_1596);
nor U3999 (N_3999,N_369,N_1278);
xnor U4000 (N_4000,N_3841,N_2802);
nor U4001 (N_4001,N_3799,N_2095);
xor U4002 (N_4002,N_3739,N_3989);
nand U4003 (N_4003,N_3816,N_3161);
nand U4004 (N_4004,N_3391,N_2386);
xnor U4005 (N_4005,N_3591,N_3599);
nor U4006 (N_4006,N_2151,N_2799);
or U4007 (N_4007,N_3221,N_3865);
xnor U4008 (N_4008,N_3588,N_2755);
xnor U4009 (N_4009,N_2690,N_3966);
nand U4010 (N_4010,N_2679,N_3534);
and U4011 (N_4011,N_3371,N_3993);
or U4012 (N_4012,N_3255,N_2632);
and U4013 (N_4013,N_2722,N_2869);
or U4014 (N_4014,N_2963,N_2599);
xor U4015 (N_4015,N_2486,N_2245);
and U4016 (N_4016,N_2258,N_3230);
nor U4017 (N_4017,N_3565,N_2495);
nand U4018 (N_4018,N_2224,N_2041);
or U4019 (N_4019,N_2945,N_2510);
nand U4020 (N_4020,N_2838,N_2100);
nor U4021 (N_4021,N_2540,N_3846);
nand U4022 (N_4022,N_2545,N_3504);
nand U4023 (N_4023,N_2767,N_2373);
nand U4024 (N_4024,N_3090,N_3603);
nand U4025 (N_4025,N_2840,N_2173);
or U4026 (N_4026,N_3491,N_2193);
nor U4027 (N_4027,N_2729,N_3992);
nand U4028 (N_4028,N_3858,N_3696);
nand U4029 (N_4029,N_3542,N_2648);
nand U4030 (N_4030,N_3853,N_2324);
xor U4031 (N_4031,N_3044,N_2715);
and U4032 (N_4032,N_2481,N_3855);
xor U4033 (N_4033,N_3906,N_2942);
xor U4034 (N_4034,N_3208,N_3220);
xnor U4035 (N_4035,N_3765,N_3422);
nor U4036 (N_4036,N_2321,N_3000);
nor U4037 (N_4037,N_3583,N_3913);
nor U4038 (N_4038,N_2288,N_2307);
nand U4039 (N_4039,N_3875,N_3554);
and U4040 (N_4040,N_2754,N_2081);
nand U4041 (N_4041,N_3782,N_2940);
nand U4042 (N_4042,N_3613,N_2693);
and U4043 (N_4043,N_3470,N_3424);
xor U4044 (N_4044,N_2121,N_2624);
or U4045 (N_4045,N_2088,N_3452);
nand U4046 (N_4046,N_3411,N_2422);
nand U4047 (N_4047,N_2985,N_2670);
or U4048 (N_4048,N_2226,N_3012);
xor U4049 (N_4049,N_2549,N_2944);
and U4050 (N_4050,N_3407,N_3789);
and U4051 (N_4051,N_2885,N_2805);
nand U4052 (N_4052,N_3793,N_2663);
nand U4053 (N_4053,N_3496,N_3253);
nand U4054 (N_4054,N_2357,N_2308);
or U4055 (N_4055,N_2494,N_2439);
xor U4056 (N_4056,N_2039,N_3773);
nand U4057 (N_4057,N_2829,N_3500);
xor U4058 (N_4058,N_2106,N_3118);
nand U4059 (N_4059,N_2820,N_2008);
xor U4060 (N_4060,N_2668,N_3248);
nor U4061 (N_4061,N_2231,N_2279);
and U4062 (N_4062,N_3974,N_2711);
nor U4063 (N_4063,N_3414,N_3301);
xnor U4064 (N_4064,N_2118,N_2076);
nand U4065 (N_4065,N_3363,N_2793);
xnor U4066 (N_4066,N_2168,N_3561);
xor U4067 (N_4067,N_2534,N_3081);
or U4068 (N_4068,N_2927,N_3082);
or U4069 (N_4069,N_3651,N_3333);
and U4070 (N_4070,N_2678,N_3174);
xor U4071 (N_4071,N_3949,N_3585);
nor U4072 (N_4072,N_2917,N_2742);
nor U4073 (N_4073,N_3204,N_2841);
xor U4074 (N_4074,N_3990,N_3733);
nand U4075 (N_4075,N_3014,N_2908);
xor U4076 (N_4076,N_3056,N_3652);
nor U4077 (N_4077,N_2227,N_3962);
or U4078 (N_4078,N_3266,N_2865);
nand U4079 (N_4079,N_3813,N_3912);
nand U4080 (N_4080,N_3274,N_3537);
xor U4081 (N_4081,N_2978,N_2241);
and U4082 (N_4082,N_3375,N_3843);
nor U4083 (N_4083,N_3305,N_2748);
xor U4084 (N_4084,N_3807,N_2541);
nor U4085 (N_4085,N_2646,N_3478);
nor U4086 (N_4086,N_2370,N_2752);
xor U4087 (N_4087,N_3590,N_2075);
or U4088 (N_4088,N_3804,N_2220);
nor U4089 (N_4089,N_3063,N_2511);
xor U4090 (N_4090,N_2776,N_2239);
nand U4091 (N_4091,N_2016,N_2395);
nor U4092 (N_4092,N_3918,N_3594);
nand U4093 (N_4093,N_2828,N_2294);
nor U4094 (N_4094,N_3265,N_3051);
xor U4095 (N_4095,N_3776,N_2257);
and U4096 (N_4096,N_2033,N_3271);
or U4097 (N_4097,N_2929,N_3954);
nor U4098 (N_4098,N_2751,N_3436);
and U4099 (N_4099,N_3764,N_2249);
or U4100 (N_4100,N_2098,N_2652);
and U4101 (N_4101,N_3278,N_3034);
nor U4102 (N_4102,N_2529,N_3038);
and U4103 (N_4103,N_3575,N_2247);
nor U4104 (N_4104,N_3730,N_3545);
nand U4105 (N_4105,N_2737,N_3008);
or U4106 (N_4106,N_2961,N_2795);
nand U4107 (N_4107,N_2096,N_2590);
nor U4108 (N_4108,N_2285,N_3142);
nand U4109 (N_4109,N_3931,N_3708);
or U4110 (N_4110,N_2103,N_3828);
nand U4111 (N_4111,N_2413,N_3472);
or U4112 (N_4112,N_3516,N_3896);
nand U4113 (N_4113,N_2287,N_2237);
nor U4114 (N_4114,N_3936,N_2275);
and U4115 (N_4115,N_3379,N_3717);
nor U4116 (N_4116,N_2804,N_3748);
xnor U4117 (N_4117,N_3810,N_3935);
nor U4118 (N_4118,N_2566,N_2146);
xor U4119 (N_4119,N_2252,N_2688);
nand U4120 (N_4120,N_3718,N_3223);
and U4121 (N_4121,N_3699,N_3953);
and U4122 (N_4122,N_2801,N_2968);
nand U4123 (N_4123,N_2049,N_2570);
and U4124 (N_4124,N_2438,N_2617);
and U4125 (N_4125,N_3499,N_3326);
xnor U4126 (N_4126,N_3626,N_2926);
nand U4127 (N_4127,N_3300,N_3049);
and U4128 (N_4128,N_3335,N_2139);
xnor U4129 (N_4129,N_3394,N_2880);
and U4130 (N_4130,N_3131,N_3299);
xnor U4131 (N_4131,N_3930,N_2922);
and U4132 (N_4132,N_2325,N_3361);
xor U4133 (N_4133,N_2901,N_3829);
nand U4134 (N_4134,N_3842,N_2791);
and U4135 (N_4135,N_2107,N_3506);
and U4136 (N_4136,N_2085,N_2971);
nand U4137 (N_4137,N_3308,N_3721);
and U4138 (N_4138,N_3997,N_2983);
nand U4139 (N_4139,N_3083,N_2519);
xnor U4140 (N_4140,N_2293,N_3244);
nand U4141 (N_4141,N_2994,N_3973);
nand U4142 (N_4142,N_2572,N_2444);
nor U4143 (N_4143,N_3454,N_2728);
nand U4144 (N_4144,N_3323,N_3830);
nand U4145 (N_4145,N_3701,N_3844);
nand U4146 (N_4146,N_2031,N_2695);
nand U4147 (N_4147,N_3285,N_3911);
nor U4148 (N_4148,N_3073,N_2027);
nor U4149 (N_4149,N_3756,N_2195);
xor U4150 (N_4150,N_2595,N_3181);
nor U4151 (N_4151,N_3010,N_2986);
and U4152 (N_4152,N_3279,N_3895);
nand U4153 (N_4153,N_2750,N_3729);
nor U4154 (N_4154,N_3381,N_2565);
xnor U4155 (N_4155,N_3768,N_3901);
or U4156 (N_4156,N_2777,N_2077);
nand U4157 (N_4157,N_3130,N_3840);
nand U4158 (N_4158,N_3540,N_3463);
nor U4159 (N_4159,N_3283,N_3607);
nand U4160 (N_4160,N_3571,N_3137);
xor U4161 (N_4161,N_3801,N_3218);
nand U4162 (N_4162,N_2764,N_2980);
or U4163 (N_4163,N_3369,N_3107);
and U4164 (N_4164,N_2347,N_3523);
nor U4165 (N_4165,N_3526,N_2503);
or U4166 (N_4166,N_3883,N_2655);
or U4167 (N_4167,N_2127,N_3176);
or U4168 (N_4168,N_2708,N_3473);
or U4169 (N_4169,N_3580,N_3129);
xnor U4170 (N_4170,N_2666,N_2061);
or U4171 (N_4171,N_2558,N_2500);
xor U4172 (N_4172,N_2618,N_3178);
and U4173 (N_4173,N_3249,N_3400);
nor U4174 (N_4174,N_2399,N_3502);
xnor U4175 (N_4175,N_2587,N_2768);
nand U4176 (N_4176,N_2485,N_2034);
xor U4177 (N_4177,N_3541,N_3268);
or U4178 (N_4178,N_3643,N_3483);
xnor U4179 (N_4179,N_2640,N_2406);
and U4180 (N_4180,N_2866,N_3630);
nand U4181 (N_4181,N_2067,N_3031);
xnor U4182 (N_4182,N_3444,N_2235);
xnor U4183 (N_4183,N_3214,N_3548);
or U4184 (N_4184,N_3040,N_2845);
and U4185 (N_4185,N_3766,N_2142);
or U4186 (N_4186,N_2643,N_2291);
and U4187 (N_4187,N_2456,N_2167);
or U4188 (N_4188,N_2197,N_2114);
xor U4189 (N_4189,N_3557,N_2082);
nand U4190 (N_4190,N_3486,N_2011);
xnor U4191 (N_4191,N_3309,N_2527);
nand U4192 (N_4192,N_2327,N_3201);
and U4193 (N_4193,N_3886,N_3149);
nand U4194 (N_4194,N_3426,N_2786);
xor U4195 (N_4195,N_2478,N_2302);
nand U4196 (N_4196,N_3354,N_3552);
or U4197 (N_4197,N_2977,N_3744);
or U4198 (N_4198,N_2248,N_2369);
nor U4199 (N_4199,N_3724,N_2615);
xor U4200 (N_4200,N_2610,N_3209);
nor U4201 (N_4201,N_2789,N_2255);
or U4202 (N_4202,N_3295,N_3888);
and U4203 (N_4203,N_2178,N_3314);
nor U4204 (N_4204,N_3634,N_2130);
nand U4205 (N_4205,N_2554,N_2072);
or U4206 (N_4206,N_3374,N_3487);
nand U4207 (N_4207,N_3934,N_3995);
and U4208 (N_4208,N_3264,N_2959);
and U4209 (N_4209,N_3958,N_2600);
nor U4210 (N_4210,N_2625,N_3240);
and U4211 (N_4211,N_2488,N_2660);
and U4212 (N_4212,N_3179,N_2411);
nand U4213 (N_4213,N_2561,N_2743);
nor U4214 (N_4214,N_2872,N_3796);
or U4215 (N_4215,N_3458,N_3380);
nor U4216 (N_4216,N_3382,N_2837);
nor U4217 (N_4217,N_3774,N_2057);
xor U4218 (N_4218,N_3342,N_3141);
xnor U4219 (N_4219,N_2188,N_2713);
xnor U4220 (N_4220,N_3908,N_3693);
and U4221 (N_4221,N_2148,N_3133);
or U4222 (N_4222,N_2576,N_3654);
nor U4223 (N_4223,N_3680,N_2622);
or U4224 (N_4224,N_2087,N_3648);
or U4225 (N_4225,N_2437,N_3398);
xor U4226 (N_4226,N_2110,N_2425);
and U4227 (N_4227,N_3315,N_3926);
nor U4228 (N_4228,N_3100,N_2333);
or U4229 (N_4229,N_3370,N_3755);
nor U4230 (N_4230,N_3408,N_2256);
nand U4231 (N_4231,N_3015,N_2338);
xnor U4232 (N_4232,N_2296,N_2734);
nor U4233 (N_4233,N_3011,N_2273);
or U4234 (N_4234,N_3869,N_2380);
nand U4235 (N_4235,N_3199,N_3356);
and U4236 (N_4236,N_3719,N_2318);
or U4237 (N_4237,N_3505,N_3597);
and U4238 (N_4238,N_3263,N_2292);
nand U4239 (N_4239,N_3684,N_2430);
and U4240 (N_4240,N_3642,N_2807);
and U4241 (N_4241,N_2521,N_2765);
nand U4242 (N_4242,N_3509,N_2138);
xor U4243 (N_4243,N_2557,N_2390);
nor U4244 (N_4244,N_3318,N_2991);
nor U4245 (N_4245,N_3903,N_2211);
nor U4246 (N_4246,N_3212,N_3441);
xor U4247 (N_4247,N_3944,N_3569);
or U4248 (N_4248,N_3294,N_2040);
xor U4249 (N_4249,N_3405,N_2973);
or U4250 (N_4250,N_3564,N_3861);
and U4251 (N_4251,N_2209,N_2900);
nor U4252 (N_4252,N_3809,N_2161);
nand U4253 (N_4253,N_2493,N_3749);
or U4254 (N_4254,N_2140,N_2054);
and U4255 (N_4255,N_3258,N_3093);
nand U4256 (N_4256,N_3827,N_2024);
or U4257 (N_4257,N_2830,N_3215);
or U4258 (N_4258,N_3211,N_2542);
or U4259 (N_4259,N_2143,N_2998);
or U4260 (N_4260,N_3728,N_3153);
nor U4261 (N_4261,N_2391,N_2176);
or U4262 (N_4262,N_2170,N_3267);
or U4263 (N_4263,N_2310,N_2923);
or U4264 (N_4264,N_2070,N_3501);
xor U4265 (N_4265,N_3753,N_2996);
nor U4266 (N_4266,N_3399,N_3546);
or U4267 (N_4267,N_3567,N_2361);
and U4268 (N_4268,N_3225,N_3256);
or U4269 (N_4269,N_3835,N_2069);
or U4270 (N_4270,N_3115,N_3951);
and U4271 (N_4271,N_2891,N_3175);
or U4272 (N_4272,N_2320,N_3821);
nor U4273 (N_4273,N_2903,N_3233);
nand U4274 (N_4274,N_3982,N_3635);
and U4275 (N_4275,N_2536,N_2946);
and U4276 (N_4276,N_2912,N_2634);
nor U4277 (N_4277,N_2126,N_2638);
and U4278 (N_4278,N_2233,N_2145);
or U4279 (N_4279,N_2407,N_2890);
and U4280 (N_4280,N_3905,N_2611);
nand U4281 (N_4281,N_2440,N_2303);
nand U4282 (N_4282,N_2585,N_2109);
or U4283 (N_4283,N_3515,N_3018);
xnor U4284 (N_4284,N_3046,N_2770);
and U4285 (N_4285,N_3289,N_3525);
nor U4286 (N_4286,N_3581,N_3879);
or U4287 (N_4287,N_2219,N_3146);
and U4288 (N_4288,N_2272,N_3067);
xnor U4289 (N_4289,N_2642,N_2524);
and U4290 (N_4290,N_3519,N_3372);
nor U4291 (N_4291,N_3938,N_3324);
or U4292 (N_4292,N_2414,N_2965);
and U4293 (N_4293,N_3440,N_3064);
nand U4294 (N_4294,N_3328,N_3579);
nor U4295 (N_4295,N_3893,N_2271);
nor U4296 (N_4296,N_2925,N_2286);
and U4297 (N_4297,N_3102,N_3672);
nand U4298 (N_4298,N_2892,N_3980);
nand U4299 (N_4299,N_2852,N_3638);
nor U4300 (N_4300,N_2990,N_2471);
or U4301 (N_4301,N_2396,N_2836);
and U4302 (N_4302,N_3885,N_2919);
nand U4303 (N_4303,N_2862,N_2215);
xor U4304 (N_4304,N_2939,N_2179);
nand U4305 (N_4305,N_3725,N_3060);
xnor U4306 (N_4306,N_2367,N_2060);
nor U4307 (N_4307,N_3057,N_2479);
and U4308 (N_4308,N_3661,N_2026);
and U4309 (N_4309,N_2492,N_2019);
xnor U4310 (N_4310,N_3246,N_3600);
and U4311 (N_4311,N_3815,N_3033);
xnor U4312 (N_4312,N_2433,N_2342);
xnor U4313 (N_4313,N_2629,N_2556);
or U4314 (N_4314,N_2879,N_3132);
xor U4315 (N_4315,N_3737,N_3117);
nor U4316 (N_4316,N_3147,N_3606);
nor U4317 (N_4317,N_2465,N_3723);
nor U4318 (N_4318,N_2544,N_3593);
or U4319 (N_4319,N_3862,N_3197);
nor U4320 (N_4320,N_3646,N_3629);
nor U4321 (N_4321,N_2006,N_3494);
and U4322 (N_4322,N_3670,N_2874);
nand U4323 (N_4323,N_3679,N_3668);
nor U4324 (N_4324,N_2048,N_2654);
or U4325 (N_4325,N_2208,N_3800);
and U4326 (N_4326,N_2066,N_2575);
nor U4327 (N_4327,N_3514,N_2135);
and U4328 (N_4328,N_3711,N_2468);
or U4329 (N_4329,N_3450,N_3775);
nand U4330 (N_4330,N_2482,N_3251);
nand U4331 (N_4331,N_2893,N_2210);
nor U4332 (N_4332,N_2661,N_2045);
and U4333 (N_4333,N_3608,N_2354);
or U4334 (N_4334,N_3448,N_3669);
or U4335 (N_4335,N_2009,N_3415);
nor U4336 (N_4336,N_3019,N_2833);
xnor U4337 (N_4337,N_2111,N_2372);
xnor U4338 (N_4338,N_3162,N_3769);
or U4339 (N_4339,N_3662,N_2888);
xor U4340 (N_4340,N_2032,N_2094);
and U4341 (N_4341,N_2234,N_2763);
nand U4342 (N_4342,N_3657,N_3316);
or U4343 (N_4343,N_3229,N_3006);
and U4344 (N_4344,N_3462,N_3104);
or U4345 (N_4345,N_2749,N_3849);
xnor U4346 (N_4346,N_3868,N_2059);
nor U4347 (N_4347,N_2201,N_3059);
and U4348 (N_4348,N_2603,N_2964);
nand U4349 (N_4349,N_2924,N_3103);
and U4350 (N_4350,N_2086,N_3467);
nand U4351 (N_4351,N_2309,N_2577);
or U4352 (N_4352,N_3280,N_2207);
or U4353 (N_4353,N_3836,N_2199);
nor U4354 (N_4354,N_3427,N_3975);
nor U4355 (N_4355,N_2403,N_2689);
and U4356 (N_4356,N_2868,N_2680);
and U4357 (N_4357,N_2571,N_3021);
nand U4358 (N_4358,N_2604,N_2909);
or U4359 (N_4359,N_2475,N_2899);
nor U4360 (N_4360,N_3517,N_3979);
nor U4361 (N_4361,N_2499,N_2254);
or U4362 (N_4362,N_3741,N_3872);
or U4363 (N_4363,N_2867,N_3080);
and U4364 (N_4364,N_3282,N_2636);
xor U4365 (N_4365,N_3108,N_3653);
xnor U4366 (N_4366,N_2317,N_2474);
and U4367 (N_4367,N_3751,N_2366);
xnor U4368 (N_4368,N_2788,N_2123);
or U4369 (N_4369,N_3095,N_3678);
nor U4370 (N_4370,N_3584,N_3094);
nor U4371 (N_4371,N_3947,N_2739);
nor U4372 (N_4372,N_3464,N_3009);
xnor U4373 (N_4373,N_2261,N_3601);
nand U4374 (N_4374,N_2567,N_3121);
nor U4375 (N_4375,N_3705,N_2731);
and U4376 (N_4376,N_2476,N_3859);
and U4377 (N_4377,N_3417,N_3919);
and U4378 (N_4378,N_3633,N_3035);
or U4379 (N_4379,N_3819,N_3941);
or U4380 (N_4380,N_3479,N_3984);
or U4381 (N_4381,N_3216,N_3163);
or U4382 (N_4382,N_3961,N_3948);
xnor U4383 (N_4383,N_2163,N_3043);
nor U4384 (N_4384,N_2483,N_2811);
and U4385 (N_4385,N_3784,N_2677);
xor U4386 (N_4386,N_2269,N_3402);
and U4387 (N_4387,N_2972,N_3732);
or U4388 (N_4388,N_3053,N_3498);
nor U4389 (N_4389,N_3845,N_2259);
or U4390 (N_4390,N_3965,N_2953);
or U4391 (N_4391,N_3419,N_2270);
and U4392 (N_4392,N_3114,N_3239);
nand U4393 (N_4393,N_2284,N_2472);
or U4394 (N_4394,N_3978,N_3671);
or U4395 (N_4395,N_3425,N_2598);
nor U4396 (N_4396,N_2954,N_3898);
or U4397 (N_4397,N_3574,N_2800);
xor U4398 (N_4398,N_2581,N_2131);
and U4399 (N_4399,N_3549,N_3072);
xnor U4400 (N_4400,N_3917,N_3771);
and U4401 (N_4401,N_2671,N_3418);
nand U4402 (N_4402,N_3281,N_3207);
or U4403 (N_4403,N_3122,N_2504);
or U4404 (N_4404,N_2623,N_2274);
nand U4405 (N_4405,N_2683,N_2280);
xor U4406 (N_4406,N_3303,N_3939);
nand U4407 (N_4407,N_2522,N_3431);
and U4408 (N_4408,N_3320,N_2855);
xnor U4409 (N_4409,N_2993,N_3459);
and U4410 (N_4410,N_3481,N_3442);
xnor U4411 (N_4411,N_3412,N_2563);
and U4412 (N_4412,N_2970,N_3946);
and U4413 (N_4413,N_3077,N_3359);
or U4414 (N_4414,N_2267,N_2778);
xor U4415 (N_4415,N_3192,N_2952);
nand U4416 (N_4416,N_3030,N_3928);
nand U4417 (N_4417,N_3779,N_3173);
xnor U4418 (N_4418,N_2134,N_2229);
nand U4419 (N_4419,N_3864,N_2477);
xor U4420 (N_4420,N_2716,N_3937);
nor U4421 (N_4421,N_2136,N_2621);
and U4422 (N_4422,N_2796,N_2160);
and U4423 (N_4423,N_3378,N_3269);
nand U4424 (N_4424,N_2336,N_3409);
or U4425 (N_4425,N_2079,N_3139);
nor U4426 (N_4426,N_2526,N_3558);
nor U4427 (N_4427,N_2808,N_3511);
or U4428 (N_4428,N_2348,N_3276);
and U4429 (N_4429,N_2817,N_3145);
xor U4430 (N_4430,N_3169,N_2873);
xor U4431 (N_4431,N_3120,N_2289);
xnor U4432 (N_4432,N_2304,N_3039);
or U4433 (N_4433,N_3362,N_2305);
and U4434 (N_4434,N_2794,N_3631);
or U4435 (N_4435,N_3609,N_3856);
nand U4436 (N_4436,N_3522,N_3002);
nor U4437 (N_4437,N_3164,N_3451);
nor U4438 (N_4438,N_3636,N_2513);
and U4439 (N_4439,N_2108,N_2378);
and U4440 (N_4440,N_3924,N_2810);
nor U4441 (N_4441,N_2191,N_3736);
or U4442 (N_4442,N_2446,N_3570);
nand U4443 (N_4443,N_3433,N_3143);
xor U4444 (N_4444,N_2605,N_2218);
and U4445 (N_4445,N_3313,N_2155);
xnor U4446 (N_4446,N_2735,N_2958);
or U4447 (N_4447,N_2686,N_2343);
or U4448 (N_4448,N_3017,N_2803);
and U4449 (N_4449,N_2637,N_3337);
xnor U4450 (N_4450,N_2185,N_3183);
xor U4451 (N_4451,N_3406,N_3687);
xor U4452 (N_4452,N_3507,N_3388);
or U4453 (N_4453,N_2449,N_2417);
xor U4454 (N_4454,N_2460,N_3620);
nor U4455 (N_4455,N_3759,N_3111);
or U4456 (N_4456,N_2911,N_2601);
or U4457 (N_4457,N_2962,N_3389);
nand U4458 (N_4458,N_3468,N_3837);
nor U4459 (N_4459,N_2064,N_2698);
and U4460 (N_4460,N_2594,N_2806);
nor U4461 (N_4461,N_2129,N_2074);
or U4462 (N_4462,N_2265,N_2694);
nor U4463 (N_4463,N_3113,N_2532);
and U4464 (N_4464,N_2498,N_2659);
or U4465 (N_4465,N_2651,N_2989);
xor U4466 (N_4466,N_3834,N_2117);
nand U4467 (N_4467,N_3848,N_2895);
and U4468 (N_4468,N_3887,N_2539);
nor U4469 (N_4469,N_2152,N_2453);
or U4470 (N_4470,N_3177,N_2635);
xnor U4471 (N_4471,N_2051,N_2010);
or U4472 (N_4472,N_2382,N_3101);
nor U4473 (N_4473,N_3760,N_2533);
and U4474 (N_4474,N_3128,N_3761);
and U4475 (N_4475,N_3092,N_2782);
and U4476 (N_4476,N_2746,N_3559);
or U4477 (N_4477,N_3503,N_2757);
or U4478 (N_4478,N_2166,N_3539);
nor U4479 (N_4479,N_3762,N_3054);
nor U4480 (N_4480,N_2685,N_3871);
and U4481 (N_4481,N_3079,N_2337);
nand U4482 (N_4482,N_2180,N_2781);
nand U4483 (N_4483,N_3803,N_2171);
or U4484 (N_4484,N_2712,N_3219);
or U4485 (N_4485,N_2720,N_2022);
and U4486 (N_4486,N_2353,N_2740);
nand U4487 (N_4487,N_2362,N_3692);
and U4488 (N_4488,N_2835,N_2555);
nand U4489 (N_4489,N_2863,N_3640);
nand U4490 (N_4490,N_2298,N_2410);
nand U4491 (N_4491,N_3618,N_2282);
xor U4492 (N_4492,N_2150,N_2232);
and U4493 (N_4493,N_3573,N_2169);
or U4494 (N_4494,N_3825,N_2931);
and U4495 (N_4495,N_3242,N_3656);
and U4496 (N_4496,N_3791,N_3780);
or U4497 (N_4497,N_3685,N_2470);
or U4498 (N_4498,N_2091,N_3622);
nand U4499 (N_4499,N_2394,N_3619);
nor U4500 (N_4500,N_2859,N_2156);
nand U4501 (N_4501,N_2930,N_2606);
nand U4502 (N_4502,N_3206,N_3710);
and U4503 (N_4503,N_2672,N_3644);
nor U4504 (N_4504,N_3048,N_3460);
nand U4505 (N_4505,N_2976,N_3469);
nor U4506 (N_4506,N_3932,N_3790);
or U4507 (N_4507,N_2200,N_2662);
nor U4508 (N_4508,N_3332,N_3513);
and U4509 (N_4509,N_3832,N_3550);
nand U4510 (N_4510,N_3186,N_3476);
and U4511 (N_4511,N_3495,N_3614);
or U4512 (N_4512,N_2774,N_3838);
nand U4513 (N_4513,N_3602,N_2316);
xnor U4514 (N_4514,N_3658,N_3555);
or U4515 (N_4515,N_2339,N_3783);
or U4516 (N_4516,N_2723,N_3527);
xor U4517 (N_4517,N_2627,N_2424);
and U4518 (N_4518,N_3287,N_3061);
and U4519 (N_4519,N_2507,N_3125);
nor U4520 (N_4520,N_2432,N_2276);
nor U4521 (N_4521,N_2246,N_2824);
or U4522 (N_4522,N_2260,N_2352);
xnor U4523 (N_4523,N_2915,N_3387);
or U4524 (N_4524,N_3488,N_2484);
nand U4525 (N_4525,N_2047,N_2564);
and U4526 (N_4526,N_3284,N_3676);
and U4527 (N_4527,N_3312,N_2984);
nor U4528 (N_4528,N_2351,N_2408);
or U4529 (N_4529,N_2614,N_2137);
or U4530 (N_4530,N_3493,N_3528);
nor U4531 (N_4531,N_3976,N_2080);
and U4532 (N_4532,N_3876,N_2910);
xor U4533 (N_4533,N_2725,N_2738);
xnor U4534 (N_4534,N_3675,N_3490);
nor U4535 (N_4535,N_3410,N_2692);
nor U4536 (N_4536,N_2398,N_2950);
nor U4537 (N_4537,N_2999,N_2847);
nor U4538 (N_4538,N_2423,N_2882);
and U4539 (N_4539,N_2790,N_2431);
nand U4540 (N_4540,N_3532,N_2724);
nand U4541 (N_4541,N_2797,N_3329);
xor U4542 (N_4542,N_3920,N_3972);
or U4543 (N_4543,N_3860,N_3377);
and U4544 (N_4544,N_2462,N_3797);
xor U4545 (N_4545,N_2773,N_2102);
xnor U4546 (N_4546,N_2848,N_2987);
nor U4547 (N_4547,N_3632,N_3826);
or U4548 (N_4548,N_2875,N_3623);
and U4549 (N_4549,N_3074,N_2042);
nor U4550 (N_4550,N_2938,N_2175);
or U4551 (N_4551,N_3392,N_3345);
nand U4552 (N_4552,N_3822,N_2898);
xor U4553 (N_4553,N_2568,N_2251);
xor U4554 (N_4554,N_3850,N_3076);
nand U4555 (N_4555,N_3649,N_3727);
and U4556 (N_4556,N_3738,N_2012);
xor U4557 (N_4557,N_3105,N_3004);
or U4558 (N_4558,N_3851,N_2125);
xor U4559 (N_4559,N_3228,N_3187);
or U4560 (N_4560,N_3945,N_2906);
nor U4561 (N_4561,N_3191,N_3706);
or U4562 (N_4562,N_2681,N_2747);
or U4563 (N_4563,N_3655,N_3884);
xnor U4564 (N_4564,N_3322,N_3307);
nor U4565 (N_4565,N_3624,N_3817);
xor U4566 (N_4566,N_3551,N_2023);
nand U4567 (N_4567,N_2839,N_3794);
or U4568 (N_4568,N_2083,N_3891);
nand U4569 (N_4569,N_2537,N_3743);
or U4570 (N_4570,N_2459,N_3112);
xor U4571 (N_4571,N_3690,N_3712);
nand U4572 (N_4572,N_2913,N_2376);
nor U4573 (N_4573,N_3866,N_3275);
or U4574 (N_4574,N_3942,N_2955);
and U4575 (N_4575,N_2402,N_2543);
nor U4576 (N_4576,N_2512,N_3716);
or U4577 (N_4577,N_3290,N_2182);
nor U4578 (N_4578,N_3172,N_3365);
nand U4579 (N_4579,N_3272,N_3533);
nor U4580 (N_4580,N_2214,N_3005);
and U4581 (N_4581,N_3025,N_2467);
nor U4582 (N_4582,N_2093,N_3754);
and U4583 (N_4583,N_2328,N_3098);
nand U4584 (N_4584,N_3792,N_3330);
and U4585 (N_4585,N_3196,N_3273);
nand U4586 (N_4586,N_2957,N_3109);
and U4587 (N_4587,N_2877,N_3231);
xor U4588 (N_4588,N_3259,N_3957);
nor U4589 (N_4589,N_2818,N_2050);
xnor U4590 (N_4590,N_3445,N_2326);
nand U4591 (N_4591,N_3075,N_3024);
xor U4592 (N_4592,N_2078,N_3171);
xor U4593 (N_4593,N_2497,N_2489);
xnor U4594 (N_4594,N_2871,N_3547);
nor U4595 (N_4595,N_2089,N_3434);
and U4596 (N_4596,N_3022,N_3262);
and U4597 (N_4597,N_2823,N_2569);
xnor U4598 (N_4598,N_2014,N_2969);
and U4599 (N_4599,N_2916,N_3304);
nand U4600 (N_4600,N_3795,N_2616);
xor U4601 (N_4601,N_3820,N_2612);
xnor U4602 (N_4602,N_2853,N_3852);
xnor U4603 (N_4603,N_3786,N_3346);
or U4604 (N_4604,N_3050,N_2619);
and U4605 (N_4605,N_3742,N_2473);
xor U4606 (N_4606,N_3438,N_3689);
and U4607 (N_4607,N_2266,N_3894);
xnor U4608 (N_4608,N_2223,N_3007);
nand U4609 (N_4609,N_3616,N_3461);
nand U4610 (N_4610,N_2018,N_2858);
nor U4611 (N_4611,N_2189,N_3747);
nand U4612 (N_4612,N_2592,N_2918);
and U4613 (N_4613,N_3047,N_3235);
xor U4614 (N_4614,N_3683,N_3252);
or U4615 (N_4615,N_3420,N_2429);
or U4616 (N_4616,N_3787,N_2884);
nand U4617 (N_4617,N_2345,N_2461);
and U4618 (N_4618,N_3612,N_3116);
nor U4619 (N_4619,N_3099,N_3151);
and U4620 (N_4620,N_2517,N_3874);
xnor U4621 (N_4621,N_2198,N_3126);
xnor U4622 (N_4622,N_3155,N_3432);
nand U4623 (N_4623,N_3562,N_2330);
xor U4624 (N_4624,N_2092,N_3510);
or U4625 (N_4625,N_3715,N_3956);
xor U4626 (N_4626,N_3368,N_2787);
xnor U4627 (N_4627,N_2037,N_3664);
nand U4628 (N_4628,N_2158,N_2626);
nor U4629 (N_4629,N_2052,N_2596);
nand U4630 (N_4630,N_2584,N_3097);
nand U4631 (N_4631,N_2658,N_3396);
nor U4632 (N_4632,N_2508,N_2933);
or U4633 (N_4633,N_3996,N_3847);
nor U4634 (N_4634,N_2613,N_2084);
xnor U4635 (N_4635,N_2936,N_3971);
or U4636 (N_4636,N_2350,N_2726);
xor U4637 (N_4637,N_3933,N_2727);
and U4638 (N_4638,N_2535,N_3878);
and U4639 (N_4639,N_2277,N_2332);
nand U4640 (N_4640,N_2821,N_2502);
or U4641 (N_4641,N_2186,N_3811);
or U4642 (N_4642,N_2664,N_2881);
or U4643 (N_4643,N_3088,N_3041);
or U4644 (N_4644,N_3222,N_3697);
nor U4645 (N_4645,N_2719,N_3350);
or U4646 (N_4646,N_2988,N_3189);
or U4647 (N_4647,N_2520,N_2547);
nand U4648 (N_4648,N_3217,N_2981);
and U4649 (N_4649,N_3645,N_3677);
nand U4650 (N_4650,N_3205,N_2409);
or U4651 (N_4651,N_3416,N_2886);
nor U4652 (N_4652,N_3232,N_3798);
xor U4653 (N_4653,N_3288,N_3480);
and U4654 (N_4654,N_2013,N_3037);
and U4655 (N_4655,N_3226,N_3682);
xnor U4656 (N_4656,N_2812,N_3310);
nand U4657 (N_4657,N_3203,N_2714);
or U4658 (N_4658,N_2974,N_3777);
nand U4659 (N_4659,N_3812,N_3731);
or U4660 (N_4660,N_2870,N_2753);
or U4661 (N_4661,N_2177,N_3306);
nor U4662 (N_4662,N_2721,N_3302);
nand U4663 (N_4663,N_2044,N_2697);
or U4664 (N_4664,N_2609,N_3681);
and U4665 (N_4665,N_3563,N_3625);
nor U4666 (N_4666,N_2744,N_3297);
nand U4667 (N_4667,N_3123,N_2063);
and U4668 (N_4668,N_2458,N_3909);
xnor U4669 (N_4669,N_2344,N_2043);
nand U4670 (N_4670,N_3621,N_3720);
or U4671 (N_4671,N_2673,N_3700);
and U4672 (N_4672,N_2300,N_3998);
nand U4673 (N_4673,N_2928,N_3556);
and U4674 (N_4674,N_2992,N_3032);
or U4675 (N_4675,N_2667,N_3960);
nor U4676 (N_4676,N_3386,N_3344);
and U4677 (N_4677,N_2216,N_2639);
xor U4678 (N_4678,N_2466,N_2115);
and U4679 (N_4679,N_2358,N_3160);
nand U4680 (N_4680,N_3802,N_2665);
nor U4681 (N_4681,N_3453,N_3355);
nand U4682 (N_4682,N_2213,N_2384);
nor U4683 (N_4683,N_3213,N_2515);
or U4684 (N_4684,N_3358,N_2703);
or U4685 (N_4685,N_2894,N_2937);
nor U4686 (N_4686,N_2450,N_3292);
or U4687 (N_4687,N_2240,N_3003);
or U4688 (N_4688,N_3311,N_3071);
nand U4689 (N_4689,N_2691,N_2181);
nand U4690 (N_4690,N_2704,N_2202);
and U4691 (N_4691,N_2844,N_3397);
or U4692 (N_4692,N_3923,N_2035);
nor U4693 (N_4693,N_3227,N_2878);
nand U4694 (N_4694,N_3767,N_2580);
nor U4695 (N_4695,N_3376,N_3224);
xor U4696 (N_4696,N_3028,N_3535);
xor U4697 (N_4697,N_2419,N_3695);
and U4698 (N_4698,N_2128,N_3013);
nor U4699 (N_4699,N_3950,N_2000);
and U4700 (N_4700,N_2206,N_2448);
xor U4701 (N_4701,N_2586,N_3757);
nand U4702 (N_4702,N_2434,N_2331);
or U4703 (N_4703,N_3135,N_3892);
nor U4704 (N_4704,N_2834,N_2525);
nor U4705 (N_4705,N_2184,N_3994);
nor U4706 (N_4706,N_3156,N_2015);
xnor U4707 (N_4707,N_2154,N_2588);
nand U4708 (N_4708,N_3058,N_2701);
or U4709 (N_4709,N_2124,N_3910);
xor U4710 (N_4710,N_3647,N_2745);
or U4711 (N_4711,N_3138,N_2196);
or U4712 (N_4712,N_2732,N_3465);
nand U4713 (N_4713,N_3566,N_2225);
xor U4714 (N_4714,N_2187,N_2920);
xor U4715 (N_4715,N_2113,N_2644);
or U4716 (N_4716,N_2204,N_2030);
and U4717 (N_4717,N_3395,N_3598);
or U4718 (N_4718,N_3423,N_3045);
or U4719 (N_4719,N_2967,N_2203);
nor U4720 (N_4720,N_2392,N_2975);
xnor U4721 (N_4721,N_2290,N_3384);
or U4722 (N_4722,N_3351,N_2283);
nand U4723 (N_4723,N_3691,N_2707);
nor U4724 (N_4724,N_2949,N_2190);
or U4725 (N_4725,N_3870,N_2278);
and U4726 (N_4726,N_2335,N_2851);
or U4727 (N_4727,N_2645,N_2491);
or U4728 (N_4728,N_2506,N_3578);
or U4729 (N_4729,N_2120,N_3474);
or U4730 (N_4730,N_2730,N_2205);
or U4731 (N_4731,N_3257,N_2675);
nor U4732 (N_4732,N_2029,N_2228);
xnor U4733 (N_4733,N_3703,N_2766);
xor U4734 (N_4734,N_2244,N_3091);
or U4735 (N_4735,N_2383,N_2579);
nor U4736 (N_4736,N_2427,N_2001);
or U4737 (N_4737,N_2454,N_2560);
or U4738 (N_4738,N_2020,N_3746);
nand U4739 (N_4739,N_2597,N_2887);
xor U4740 (N_4740,N_2705,N_3512);
nor U4741 (N_4741,N_2153,N_2551);
nor U4742 (N_4742,N_3148,N_3673);
xnor U4743 (N_4743,N_3319,N_2375);
nor U4744 (N_4744,N_2116,N_3968);
xor U4745 (N_4745,N_3674,N_2412);
xor U4746 (N_4746,N_2736,N_2105);
nand U4747 (N_4747,N_2090,N_3611);
nand U4748 (N_4748,N_2144,N_3357);
xnor U4749 (N_4749,N_3881,N_2349);
nor U4750 (N_4750,N_2772,N_2490);
xnor U4751 (N_4751,N_2299,N_3202);
and U4752 (N_4752,N_3986,N_2784);
xnor U4753 (N_4753,N_3688,N_3430);
or U4754 (N_4754,N_2897,N_3814);
and U4755 (N_4755,N_3615,N_2162);
and U4756 (N_4756,N_2559,N_2819);
and U4757 (N_4757,N_3068,N_2388);
xor U4758 (N_4758,N_2825,N_3752);
or U4759 (N_4759,N_3666,N_3985);
or U4760 (N_4760,N_2792,N_2798);
or U4761 (N_4761,N_2548,N_2827);
and U4762 (N_4762,N_3194,N_2849);
or U4763 (N_4763,N_3435,N_2602);
xnor U4764 (N_4764,N_3750,N_2119);
xor U4765 (N_4765,N_3334,N_3234);
nor U4766 (N_4766,N_3052,N_2650);
or U4767 (N_4767,N_2172,N_2761);
xnor U4768 (N_4768,N_3340,N_2573);
nand U4769 (N_4769,N_3027,N_3144);
xnor U4770 (N_4770,N_3497,N_2416);
nand U4771 (N_4771,N_2436,N_3925);
nand U4772 (N_4772,N_3617,N_2487);
nor U4773 (N_4773,N_3106,N_2856);
or U4774 (N_4774,N_3243,N_2531);
nor U4775 (N_4775,N_2387,N_3066);
nand U4776 (N_4776,N_3952,N_3023);
nor U4777 (N_4777,N_3124,N_2706);
nor U4778 (N_4778,N_2400,N_2036);
nor U4779 (N_4779,N_3713,N_2389);
xnor U4780 (N_4780,N_2702,N_3321);
nor U4781 (N_4781,N_2649,N_3735);
and U4782 (N_4782,N_2003,N_2656);
nor U4783 (N_4783,N_2004,N_2062);
nand U4784 (N_4784,N_3413,N_2501);
xnor U4785 (N_4785,N_2876,N_2311);
and U4786 (N_4786,N_3134,N_3296);
nor U4787 (N_4787,N_2363,N_3200);
xnor U4788 (N_4788,N_3833,N_3195);
nand U4789 (N_4789,N_3900,N_2371);
nand U4790 (N_4790,N_2314,N_2771);
xor U4791 (N_4791,N_3250,N_2966);
nor U4792 (N_4792,N_2301,N_2591);
xnor U4793 (N_4793,N_2381,N_3360);
and U4794 (N_4794,N_2709,N_3854);
and U4795 (N_4795,N_2578,N_2262);
nand U4796 (N_4796,N_2359,N_2469);
and U4797 (N_4797,N_3922,N_2951);
and U4798 (N_4798,N_2435,N_3627);
xor U4799 (N_4799,N_2046,N_3531);
and U4800 (N_4800,N_3999,N_3650);
or U4801 (N_4801,N_2312,N_3663);
nand U4802 (N_4802,N_3457,N_2831);
and U4803 (N_4803,N_3036,N_3245);
and U4804 (N_4804,N_2905,N_3824);
xnor U4805 (N_4805,N_3343,N_3353);
xor U4806 (N_4806,N_3325,N_3484);
nor U4807 (N_4807,N_2099,N_2212);
and U4808 (N_4808,N_2242,N_2684);
and U4809 (N_4809,N_3001,N_2306);
and U4810 (N_4810,N_2864,N_2364);
nor U4811 (N_4811,N_2758,N_3443);
or U4812 (N_4812,N_3277,N_2322);
xor U4813 (N_4813,N_3403,N_3367);
or U4814 (N_4814,N_2250,N_2038);
xor U4815 (N_4815,N_3704,N_2368);
nor U4816 (N_4816,N_2514,N_2574);
nor U4817 (N_4817,N_2762,N_2315);
xor U4818 (N_4818,N_2682,N_3065);
nand U4819 (N_4819,N_2846,N_3714);
or U4820 (N_4820,N_3987,N_3210);
and U4821 (N_4821,N_2687,N_2329);
nor U4822 (N_4822,N_2159,N_3969);
or U4823 (N_4823,N_3818,N_2593);
nand U4824 (N_4824,N_2718,N_3349);
xor U4825 (N_4825,N_2676,N_2769);
xnor U4826 (N_4826,N_3763,N_3026);
and U4827 (N_4827,N_2323,N_2264);
nor U4828 (N_4828,N_3449,N_3270);
and U4829 (N_4829,N_3839,N_2053);
or U4830 (N_4830,N_3429,N_2814);
xnor U4831 (N_4831,N_3639,N_3286);
or U4832 (N_4832,N_2842,N_2297);
or U4833 (N_4833,N_3694,N_2149);
nand U4834 (N_4834,N_3456,N_3152);
nand U4835 (N_4835,N_3929,N_3029);
and U4836 (N_4836,N_2860,N_2374);
or U4837 (N_4837,N_3536,N_3785);
nand U4838 (N_4838,N_3238,N_2943);
nor U4839 (N_4839,N_3062,N_3963);
xor U4840 (N_4840,N_3475,N_2700);
nand U4841 (N_4841,N_3863,N_3867);
or U4842 (N_4842,N_2377,N_2854);
or U4843 (N_4843,N_2157,N_3991);
nor U4844 (N_4844,N_2982,N_3988);
and U4845 (N_4845,N_2222,N_2295);
and U4846 (N_4846,N_3902,N_3823);
nor U4847 (N_4847,N_2710,N_3589);
and U4848 (N_4848,N_2445,N_2889);
or U4849 (N_4849,N_2447,N_3977);
xnor U4850 (N_4850,N_2941,N_3364);
nor U4851 (N_4851,N_2002,N_3069);
nor U4852 (N_4852,N_3582,N_3568);
and U4853 (N_4853,N_2165,N_3157);
xnor U4854 (N_4854,N_2068,N_3915);
xor U4855 (N_4855,N_2997,N_3291);
xnor U4856 (N_4856,N_3543,N_3492);
nor U4857 (N_4857,N_2243,N_2073);
and U4858 (N_4858,N_3390,N_3981);
or U4859 (N_4859,N_3338,N_3158);
xor U4860 (N_4860,N_2365,N_3331);
nor U4861 (N_4861,N_3236,N_2192);
and U4862 (N_4862,N_2025,N_3182);
nor U4863 (N_4863,N_2021,N_2562);
and U4864 (N_4864,N_2775,N_2132);
nand U4865 (N_4865,N_3529,N_2313);
or U4866 (N_4866,N_3168,N_3758);
or U4867 (N_4867,N_3166,N_2346);
xor U4868 (N_4868,N_2826,N_3439);
and U4869 (N_4869,N_2385,N_3707);
nor U4870 (N_4870,N_2509,N_2058);
or U4871 (N_4871,N_2921,N_2779);
nand U4872 (N_4872,N_2907,N_3772);
xnor U4873 (N_4873,N_3298,N_3089);
nand U4874 (N_4874,N_3605,N_3907);
nand U4875 (N_4875,N_3165,N_3185);
nor U4876 (N_4876,N_2759,N_3890);
or U4877 (N_4877,N_2760,N_2420);
or U4878 (N_4878,N_2194,N_3560);
nand U4879 (N_4879,N_2904,N_2451);
nor U4880 (N_4880,N_3482,N_3421);
nand U4881 (N_4881,N_2334,N_3336);
and U4882 (N_4882,N_2641,N_2340);
xor U4883 (N_4883,N_3637,N_3604);
xnor U4884 (N_4884,N_3959,N_3641);
nand U4885 (N_4885,N_2948,N_2523);
or U4886 (N_4886,N_3159,N_3595);
or U4887 (N_4887,N_2816,N_2813);
xor U4888 (N_4888,N_2133,N_3348);
nand U4889 (N_4889,N_2028,N_3184);
or U4890 (N_4890,N_3347,N_3446);
xnor U4891 (N_4891,N_2426,N_2418);
xnor U4892 (N_4892,N_2530,N_3317);
and U4893 (N_4893,N_3521,N_2696);
nor U4894 (N_4894,N_2657,N_3889);
nand U4895 (N_4895,N_3086,N_2979);
nor U4896 (N_4896,N_3726,N_2442);
xnor U4897 (N_4897,N_2947,N_3857);
nand U4898 (N_4898,N_2902,N_3383);
nand U4899 (N_4899,N_2463,N_3084);
nand U4900 (N_4900,N_3261,N_2017);
nor U4901 (N_4901,N_2379,N_3899);
or U4902 (N_4902,N_3055,N_3587);
nand U4903 (N_4903,N_2582,N_2401);
nor U4904 (N_4904,N_2785,N_2056);
xor U4905 (N_4905,N_3659,N_2393);
xor U4906 (N_4906,N_3808,N_3916);
nand U4907 (N_4907,N_3341,N_3964);
and U4908 (N_4908,N_3489,N_2850);
nor U4909 (N_4909,N_2174,N_3880);
xnor U4910 (N_4910,N_2263,N_3198);
or U4911 (N_4911,N_2452,N_3553);
nand U4912 (N_4912,N_2097,N_3921);
and U4913 (N_4913,N_3610,N_3241);
xor U4914 (N_4914,N_2464,N_3477);
nand U4915 (N_4915,N_3393,N_3665);
nor U4916 (N_4916,N_2717,N_2783);
nor U4917 (N_4917,N_2230,N_2608);
nor U4918 (N_4918,N_3327,N_2647);
nand U4919 (N_4919,N_3085,N_2883);
nand U4920 (N_4920,N_3524,N_3293);
nand U4921 (N_4921,N_3592,N_3660);
nor U4922 (N_4922,N_2236,N_2455);
nand U4923 (N_4923,N_3110,N_3538);
and U4924 (N_4924,N_3190,N_2065);
or U4925 (N_4925,N_3167,N_2809);
or U4926 (N_4926,N_3260,N_2415);
nor U4927 (N_4927,N_2589,N_2355);
xor U4928 (N_4928,N_3940,N_3873);
nor U4929 (N_4929,N_2756,N_2319);
nor U4930 (N_4930,N_2607,N_3970);
xor U4931 (N_4931,N_3897,N_2221);
or U4932 (N_4932,N_2620,N_2935);
or U4933 (N_4933,N_3577,N_2550);
nand U4934 (N_4934,N_3428,N_2546);
and U4935 (N_4935,N_3466,N_3385);
xnor U4936 (N_4936,N_3373,N_2281);
nand U4937 (N_4937,N_3967,N_3254);
nand U4938 (N_4938,N_3404,N_3070);
nor U4939 (N_4939,N_2628,N_3572);
nand U4940 (N_4940,N_3366,N_3628);
nand U4941 (N_4941,N_3042,N_3455);
xnor U4942 (N_4942,N_3020,N_2843);
nor U4943 (N_4943,N_3722,N_2356);
nor U4944 (N_4944,N_2141,N_3983);
and U4945 (N_4945,N_2104,N_3805);
nor U4946 (N_4946,N_3136,N_3518);
nand U4947 (N_4947,N_3778,N_2630);
nor U4948 (N_4948,N_2071,N_3831);
xnor U4949 (N_4949,N_2914,N_2268);
and U4950 (N_4950,N_2428,N_3914);
nor U4951 (N_4951,N_3667,N_3882);
xor U4952 (N_4952,N_3788,N_3877);
nor U4953 (N_4953,N_3170,N_3734);
and U4954 (N_4954,N_3447,N_3096);
or U4955 (N_4955,N_2934,N_2583);
xor U4956 (N_4956,N_2780,N_2932);
nand U4957 (N_4957,N_2669,N_2122);
or U4958 (N_4958,N_2457,N_2995);
and U4959 (N_4959,N_2518,N_3520);
or U4960 (N_4960,N_3339,N_3437);
nand U4961 (N_4961,N_2147,N_3596);
nor U4962 (N_4962,N_2360,N_3686);
and U4963 (N_4963,N_2699,N_2443);
or U4964 (N_4964,N_2404,N_3781);
xor U4965 (N_4965,N_3078,N_3127);
and U4966 (N_4966,N_2253,N_2341);
nand U4967 (N_4967,N_2674,N_3806);
or U4968 (N_4968,N_2538,N_3576);
or U4969 (N_4969,N_2007,N_3401);
and U4970 (N_4970,N_2896,N_2741);
or U4971 (N_4971,N_3943,N_2421);
and U4972 (N_4972,N_3180,N_2822);
or U4973 (N_4973,N_2441,N_3016);
nor U4974 (N_4974,N_3955,N_3544);
and U4975 (N_4975,N_3586,N_3485);
nand U4976 (N_4976,N_3770,N_3471);
and U4977 (N_4977,N_3740,N_2217);
nand U4978 (N_4978,N_2733,N_3698);
or U4979 (N_4979,N_3709,N_2238);
nor U4980 (N_4980,N_3237,N_2528);
xnor U4981 (N_4981,N_2960,N_3352);
nand U4982 (N_4982,N_2183,N_3508);
or U4983 (N_4983,N_2101,N_2480);
nand U4984 (N_4984,N_3140,N_2552);
nor U4985 (N_4985,N_2553,N_2633);
xnor U4986 (N_4986,N_2956,N_2653);
and U4987 (N_4987,N_3154,N_2815);
nand U4988 (N_4988,N_2505,N_2405);
or U4989 (N_4989,N_3904,N_3193);
or U4990 (N_4990,N_3119,N_2112);
and U4991 (N_4991,N_3150,N_2861);
xor U4992 (N_4992,N_2005,N_2397);
nor U4993 (N_4993,N_3927,N_2516);
or U4994 (N_4994,N_2631,N_3188);
and U4995 (N_4995,N_3745,N_3087);
nand U4996 (N_4996,N_2164,N_3247);
nor U4997 (N_4997,N_2857,N_3530);
or U4998 (N_4998,N_3702,N_2832);
nor U4999 (N_4999,N_2055,N_2496);
nor U5000 (N_5000,N_3765,N_2419);
nor U5001 (N_5001,N_2263,N_3707);
nand U5002 (N_5002,N_2156,N_2373);
xnor U5003 (N_5003,N_2106,N_2847);
or U5004 (N_5004,N_2130,N_2642);
xnor U5005 (N_5005,N_2054,N_3498);
nor U5006 (N_5006,N_3904,N_3643);
or U5007 (N_5007,N_2556,N_3318);
nor U5008 (N_5008,N_3974,N_3992);
and U5009 (N_5009,N_2356,N_2883);
xor U5010 (N_5010,N_3101,N_2408);
nor U5011 (N_5011,N_2681,N_3853);
and U5012 (N_5012,N_2674,N_3662);
xor U5013 (N_5013,N_2368,N_2068);
nand U5014 (N_5014,N_3043,N_3065);
nand U5015 (N_5015,N_3271,N_2331);
and U5016 (N_5016,N_2454,N_2680);
nor U5017 (N_5017,N_2145,N_3751);
nor U5018 (N_5018,N_3866,N_2711);
or U5019 (N_5019,N_2817,N_2323);
or U5020 (N_5020,N_2319,N_3237);
nand U5021 (N_5021,N_2111,N_2609);
or U5022 (N_5022,N_2323,N_3018);
nand U5023 (N_5023,N_3033,N_3578);
nor U5024 (N_5024,N_2645,N_3262);
nand U5025 (N_5025,N_3646,N_3634);
nand U5026 (N_5026,N_3261,N_3185);
or U5027 (N_5027,N_3372,N_3870);
nor U5028 (N_5028,N_2407,N_3496);
xor U5029 (N_5029,N_3902,N_3334);
nor U5030 (N_5030,N_2456,N_3276);
nand U5031 (N_5031,N_3326,N_2125);
xor U5032 (N_5032,N_3931,N_2675);
xor U5033 (N_5033,N_2168,N_3094);
nand U5034 (N_5034,N_2178,N_3050);
nand U5035 (N_5035,N_3495,N_2210);
or U5036 (N_5036,N_3180,N_3826);
xor U5037 (N_5037,N_3183,N_3624);
and U5038 (N_5038,N_3405,N_3875);
or U5039 (N_5039,N_2264,N_3597);
nor U5040 (N_5040,N_2502,N_2472);
and U5041 (N_5041,N_2777,N_3044);
xor U5042 (N_5042,N_2506,N_3981);
or U5043 (N_5043,N_3239,N_3461);
and U5044 (N_5044,N_2432,N_2873);
or U5045 (N_5045,N_2500,N_3262);
xor U5046 (N_5046,N_2203,N_3063);
nand U5047 (N_5047,N_3877,N_3553);
nand U5048 (N_5048,N_2910,N_2585);
nand U5049 (N_5049,N_3572,N_2908);
and U5050 (N_5050,N_2675,N_2223);
nand U5051 (N_5051,N_3890,N_3994);
and U5052 (N_5052,N_2797,N_3920);
nand U5053 (N_5053,N_2523,N_2385);
nor U5054 (N_5054,N_2812,N_3131);
nand U5055 (N_5055,N_3946,N_3303);
or U5056 (N_5056,N_3450,N_3314);
nand U5057 (N_5057,N_3991,N_2345);
nor U5058 (N_5058,N_2239,N_3855);
xor U5059 (N_5059,N_2679,N_3046);
and U5060 (N_5060,N_2218,N_2174);
nor U5061 (N_5061,N_3297,N_2218);
nand U5062 (N_5062,N_3973,N_3807);
or U5063 (N_5063,N_2204,N_2437);
xor U5064 (N_5064,N_2253,N_2926);
xor U5065 (N_5065,N_3490,N_2528);
xor U5066 (N_5066,N_3538,N_2680);
nand U5067 (N_5067,N_2594,N_3388);
nand U5068 (N_5068,N_2178,N_2224);
nor U5069 (N_5069,N_3738,N_3816);
xnor U5070 (N_5070,N_3780,N_2909);
and U5071 (N_5071,N_2764,N_2830);
nor U5072 (N_5072,N_2743,N_2475);
or U5073 (N_5073,N_2940,N_2663);
or U5074 (N_5074,N_2900,N_3542);
nand U5075 (N_5075,N_2335,N_2761);
nor U5076 (N_5076,N_3635,N_3024);
nor U5077 (N_5077,N_3135,N_3949);
and U5078 (N_5078,N_2009,N_3152);
xor U5079 (N_5079,N_2668,N_3778);
or U5080 (N_5080,N_2037,N_2152);
nor U5081 (N_5081,N_3013,N_2159);
nand U5082 (N_5082,N_2489,N_3447);
xor U5083 (N_5083,N_3473,N_2842);
nand U5084 (N_5084,N_3846,N_3282);
and U5085 (N_5085,N_2947,N_2710);
nand U5086 (N_5086,N_2236,N_3030);
nand U5087 (N_5087,N_2518,N_2670);
and U5088 (N_5088,N_3512,N_2428);
nor U5089 (N_5089,N_3636,N_2100);
or U5090 (N_5090,N_2838,N_3112);
or U5091 (N_5091,N_2120,N_2803);
nor U5092 (N_5092,N_3776,N_3523);
and U5093 (N_5093,N_3623,N_3545);
or U5094 (N_5094,N_3582,N_2647);
and U5095 (N_5095,N_3475,N_3224);
nor U5096 (N_5096,N_3494,N_2266);
nor U5097 (N_5097,N_2710,N_3352);
nor U5098 (N_5098,N_3024,N_2529);
and U5099 (N_5099,N_3712,N_3329);
nor U5100 (N_5100,N_2612,N_3169);
or U5101 (N_5101,N_3279,N_3319);
nand U5102 (N_5102,N_2280,N_2981);
or U5103 (N_5103,N_3483,N_2743);
or U5104 (N_5104,N_3975,N_2126);
nor U5105 (N_5105,N_2478,N_2830);
or U5106 (N_5106,N_3769,N_3152);
and U5107 (N_5107,N_3173,N_2900);
and U5108 (N_5108,N_3555,N_3676);
nand U5109 (N_5109,N_2547,N_3113);
and U5110 (N_5110,N_2386,N_2450);
nand U5111 (N_5111,N_3996,N_3594);
xor U5112 (N_5112,N_2865,N_3527);
or U5113 (N_5113,N_2343,N_3310);
nor U5114 (N_5114,N_3808,N_3216);
nand U5115 (N_5115,N_3636,N_3274);
nand U5116 (N_5116,N_2987,N_2762);
or U5117 (N_5117,N_2828,N_3305);
or U5118 (N_5118,N_3421,N_2110);
xor U5119 (N_5119,N_3768,N_2804);
xnor U5120 (N_5120,N_3128,N_3694);
or U5121 (N_5121,N_2142,N_2764);
or U5122 (N_5122,N_2486,N_3843);
nor U5123 (N_5123,N_2373,N_3612);
nor U5124 (N_5124,N_3983,N_2154);
nor U5125 (N_5125,N_2300,N_3545);
xnor U5126 (N_5126,N_3606,N_2766);
nand U5127 (N_5127,N_2060,N_2390);
nor U5128 (N_5128,N_2213,N_3684);
or U5129 (N_5129,N_2817,N_3856);
nor U5130 (N_5130,N_2626,N_2131);
nand U5131 (N_5131,N_3119,N_2654);
nor U5132 (N_5132,N_2966,N_3478);
nand U5133 (N_5133,N_3273,N_3938);
nor U5134 (N_5134,N_2813,N_3492);
nor U5135 (N_5135,N_3579,N_2627);
nand U5136 (N_5136,N_3175,N_2682);
or U5137 (N_5137,N_2733,N_2197);
nor U5138 (N_5138,N_3893,N_3708);
nand U5139 (N_5139,N_3930,N_2861);
nand U5140 (N_5140,N_3929,N_2013);
nand U5141 (N_5141,N_2885,N_3201);
nor U5142 (N_5142,N_3716,N_2080);
xor U5143 (N_5143,N_2082,N_3036);
nand U5144 (N_5144,N_2823,N_3801);
or U5145 (N_5145,N_3444,N_3048);
nor U5146 (N_5146,N_2677,N_2913);
and U5147 (N_5147,N_2834,N_3678);
or U5148 (N_5148,N_2060,N_3753);
or U5149 (N_5149,N_3641,N_2577);
or U5150 (N_5150,N_3249,N_3512);
or U5151 (N_5151,N_2342,N_2102);
xnor U5152 (N_5152,N_2310,N_2369);
nor U5153 (N_5153,N_3036,N_3606);
nor U5154 (N_5154,N_3903,N_2901);
and U5155 (N_5155,N_3433,N_3755);
and U5156 (N_5156,N_3737,N_2722);
xnor U5157 (N_5157,N_2569,N_3432);
xor U5158 (N_5158,N_3526,N_2484);
nor U5159 (N_5159,N_3862,N_2217);
and U5160 (N_5160,N_2227,N_3008);
nand U5161 (N_5161,N_3377,N_2827);
and U5162 (N_5162,N_2423,N_2392);
nand U5163 (N_5163,N_2961,N_3514);
or U5164 (N_5164,N_2915,N_3706);
xor U5165 (N_5165,N_2388,N_2115);
xor U5166 (N_5166,N_2172,N_2303);
or U5167 (N_5167,N_2433,N_3943);
or U5168 (N_5168,N_2251,N_2747);
nand U5169 (N_5169,N_2058,N_3240);
and U5170 (N_5170,N_2252,N_3506);
and U5171 (N_5171,N_2671,N_2519);
nor U5172 (N_5172,N_3840,N_2292);
nand U5173 (N_5173,N_3075,N_3834);
or U5174 (N_5174,N_2912,N_3306);
nand U5175 (N_5175,N_2284,N_3105);
xnor U5176 (N_5176,N_3611,N_3347);
nor U5177 (N_5177,N_3085,N_3580);
nor U5178 (N_5178,N_2794,N_2233);
xnor U5179 (N_5179,N_2596,N_2168);
nand U5180 (N_5180,N_3365,N_3798);
and U5181 (N_5181,N_3584,N_2973);
or U5182 (N_5182,N_3827,N_3921);
nor U5183 (N_5183,N_2268,N_2570);
nor U5184 (N_5184,N_2306,N_3049);
nand U5185 (N_5185,N_3924,N_2952);
nand U5186 (N_5186,N_3762,N_2325);
and U5187 (N_5187,N_3283,N_3770);
nor U5188 (N_5188,N_2396,N_3387);
xor U5189 (N_5189,N_3595,N_2488);
nand U5190 (N_5190,N_3191,N_3537);
and U5191 (N_5191,N_2979,N_3860);
or U5192 (N_5192,N_3899,N_3435);
xor U5193 (N_5193,N_3762,N_2634);
or U5194 (N_5194,N_2796,N_3297);
and U5195 (N_5195,N_3569,N_2982);
xnor U5196 (N_5196,N_3089,N_3763);
or U5197 (N_5197,N_3059,N_3766);
xor U5198 (N_5198,N_2618,N_2426);
nand U5199 (N_5199,N_2723,N_2055);
or U5200 (N_5200,N_2543,N_3483);
or U5201 (N_5201,N_3315,N_2741);
or U5202 (N_5202,N_2325,N_2858);
and U5203 (N_5203,N_2788,N_2200);
xor U5204 (N_5204,N_3675,N_2535);
nor U5205 (N_5205,N_2717,N_3775);
nor U5206 (N_5206,N_3446,N_2828);
nor U5207 (N_5207,N_3004,N_2965);
nor U5208 (N_5208,N_2425,N_3924);
and U5209 (N_5209,N_3161,N_3205);
nor U5210 (N_5210,N_3335,N_2221);
xor U5211 (N_5211,N_3598,N_2406);
and U5212 (N_5212,N_3119,N_3665);
and U5213 (N_5213,N_3948,N_3565);
and U5214 (N_5214,N_2885,N_2315);
nor U5215 (N_5215,N_3305,N_3950);
nor U5216 (N_5216,N_3286,N_2693);
or U5217 (N_5217,N_3100,N_3007);
nor U5218 (N_5218,N_3656,N_3798);
xor U5219 (N_5219,N_2999,N_2667);
nor U5220 (N_5220,N_3723,N_2334);
nand U5221 (N_5221,N_2607,N_3285);
and U5222 (N_5222,N_3958,N_3671);
or U5223 (N_5223,N_3344,N_2045);
nor U5224 (N_5224,N_2654,N_3853);
and U5225 (N_5225,N_2219,N_2866);
or U5226 (N_5226,N_2740,N_3827);
nand U5227 (N_5227,N_3949,N_3737);
xnor U5228 (N_5228,N_2178,N_3516);
nor U5229 (N_5229,N_3065,N_2927);
xor U5230 (N_5230,N_3076,N_3936);
nor U5231 (N_5231,N_3528,N_2236);
xnor U5232 (N_5232,N_3651,N_2371);
or U5233 (N_5233,N_2648,N_3116);
and U5234 (N_5234,N_3269,N_3302);
or U5235 (N_5235,N_2055,N_2215);
and U5236 (N_5236,N_3569,N_2841);
nor U5237 (N_5237,N_3229,N_3968);
or U5238 (N_5238,N_3178,N_3842);
nand U5239 (N_5239,N_2666,N_3118);
and U5240 (N_5240,N_3388,N_3188);
and U5241 (N_5241,N_2211,N_2954);
or U5242 (N_5242,N_2023,N_2540);
or U5243 (N_5243,N_3432,N_3299);
or U5244 (N_5244,N_2927,N_2594);
nand U5245 (N_5245,N_2771,N_2910);
and U5246 (N_5246,N_2523,N_2329);
nor U5247 (N_5247,N_2537,N_3986);
or U5248 (N_5248,N_3184,N_3031);
nand U5249 (N_5249,N_3919,N_2827);
nand U5250 (N_5250,N_3550,N_2481);
and U5251 (N_5251,N_2096,N_2808);
xor U5252 (N_5252,N_2864,N_3282);
nor U5253 (N_5253,N_3071,N_3355);
nor U5254 (N_5254,N_3128,N_2836);
and U5255 (N_5255,N_2588,N_3245);
xor U5256 (N_5256,N_3667,N_2307);
nor U5257 (N_5257,N_3156,N_3410);
nor U5258 (N_5258,N_2130,N_2224);
xnor U5259 (N_5259,N_3877,N_3878);
or U5260 (N_5260,N_2356,N_3850);
nor U5261 (N_5261,N_3066,N_3652);
and U5262 (N_5262,N_2701,N_3854);
or U5263 (N_5263,N_3414,N_2541);
or U5264 (N_5264,N_3478,N_3480);
nor U5265 (N_5265,N_2347,N_3109);
and U5266 (N_5266,N_3548,N_2659);
xnor U5267 (N_5267,N_3932,N_2849);
and U5268 (N_5268,N_2899,N_3077);
nand U5269 (N_5269,N_3913,N_2709);
xor U5270 (N_5270,N_2563,N_2073);
xnor U5271 (N_5271,N_2964,N_3098);
and U5272 (N_5272,N_2479,N_2921);
and U5273 (N_5273,N_3818,N_3179);
or U5274 (N_5274,N_3005,N_3708);
or U5275 (N_5275,N_3082,N_3514);
and U5276 (N_5276,N_2158,N_2320);
or U5277 (N_5277,N_2833,N_3398);
and U5278 (N_5278,N_2804,N_2171);
xnor U5279 (N_5279,N_3529,N_3661);
xor U5280 (N_5280,N_3593,N_2425);
nand U5281 (N_5281,N_3067,N_2003);
nand U5282 (N_5282,N_2530,N_3419);
and U5283 (N_5283,N_3190,N_2969);
nand U5284 (N_5284,N_3523,N_3548);
or U5285 (N_5285,N_3819,N_2507);
and U5286 (N_5286,N_2530,N_2338);
nor U5287 (N_5287,N_3782,N_3374);
xnor U5288 (N_5288,N_3822,N_3633);
xnor U5289 (N_5289,N_2464,N_2247);
xor U5290 (N_5290,N_2112,N_2843);
nand U5291 (N_5291,N_2772,N_3463);
nand U5292 (N_5292,N_2153,N_3814);
or U5293 (N_5293,N_2843,N_3421);
xor U5294 (N_5294,N_3428,N_3734);
xnor U5295 (N_5295,N_3130,N_3050);
nand U5296 (N_5296,N_3541,N_2171);
and U5297 (N_5297,N_3737,N_3982);
and U5298 (N_5298,N_2860,N_2318);
and U5299 (N_5299,N_3405,N_3433);
nor U5300 (N_5300,N_3074,N_3815);
nand U5301 (N_5301,N_2441,N_3040);
nor U5302 (N_5302,N_3835,N_3704);
nor U5303 (N_5303,N_3600,N_2543);
nor U5304 (N_5304,N_2328,N_2273);
nor U5305 (N_5305,N_3319,N_2146);
nor U5306 (N_5306,N_2816,N_2822);
nor U5307 (N_5307,N_3193,N_2398);
xnor U5308 (N_5308,N_2925,N_3960);
xor U5309 (N_5309,N_2046,N_3512);
nand U5310 (N_5310,N_2686,N_2747);
and U5311 (N_5311,N_3887,N_3905);
xnor U5312 (N_5312,N_2381,N_3850);
xor U5313 (N_5313,N_2750,N_3063);
or U5314 (N_5314,N_2843,N_2241);
nor U5315 (N_5315,N_2899,N_2998);
nor U5316 (N_5316,N_3674,N_3951);
nand U5317 (N_5317,N_3804,N_3624);
xnor U5318 (N_5318,N_2765,N_2295);
nor U5319 (N_5319,N_3195,N_2970);
and U5320 (N_5320,N_2416,N_2720);
nor U5321 (N_5321,N_3224,N_2842);
xor U5322 (N_5322,N_2164,N_3475);
or U5323 (N_5323,N_2454,N_2552);
nor U5324 (N_5324,N_3100,N_2153);
or U5325 (N_5325,N_3733,N_3847);
xnor U5326 (N_5326,N_2489,N_2374);
nand U5327 (N_5327,N_3794,N_3140);
xor U5328 (N_5328,N_3099,N_2961);
or U5329 (N_5329,N_2524,N_3182);
or U5330 (N_5330,N_2702,N_2930);
nor U5331 (N_5331,N_3584,N_2832);
xor U5332 (N_5332,N_2768,N_2919);
xor U5333 (N_5333,N_3432,N_3641);
nand U5334 (N_5334,N_2397,N_2622);
or U5335 (N_5335,N_2100,N_3564);
or U5336 (N_5336,N_2830,N_2788);
nand U5337 (N_5337,N_3639,N_2727);
or U5338 (N_5338,N_2647,N_2575);
xor U5339 (N_5339,N_2518,N_2588);
nand U5340 (N_5340,N_3259,N_2358);
nor U5341 (N_5341,N_2770,N_2536);
and U5342 (N_5342,N_3464,N_2011);
nand U5343 (N_5343,N_3545,N_3294);
and U5344 (N_5344,N_3599,N_3613);
nor U5345 (N_5345,N_3966,N_3960);
and U5346 (N_5346,N_2994,N_3847);
and U5347 (N_5347,N_2918,N_3134);
nand U5348 (N_5348,N_2915,N_3600);
and U5349 (N_5349,N_3512,N_2546);
nor U5350 (N_5350,N_2459,N_3054);
nand U5351 (N_5351,N_3234,N_3045);
or U5352 (N_5352,N_2089,N_2093);
xnor U5353 (N_5353,N_3184,N_3934);
or U5354 (N_5354,N_2218,N_2023);
or U5355 (N_5355,N_3951,N_2354);
xor U5356 (N_5356,N_2774,N_3522);
xor U5357 (N_5357,N_3562,N_3584);
and U5358 (N_5358,N_3625,N_2785);
xor U5359 (N_5359,N_3844,N_2420);
nand U5360 (N_5360,N_2520,N_3051);
and U5361 (N_5361,N_3542,N_2277);
nor U5362 (N_5362,N_2426,N_3635);
xor U5363 (N_5363,N_3628,N_2932);
nand U5364 (N_5364,N_3725,N_3111);
xor U5365 (N_5365,N_3980,N_2711);
or U5366 (N_5366,N_2101,N_2868);
or U5367 (N_5367,N_2472,N_2087);
or U5368 (N_5368,N_3209,N_2225);
nand U5369 (N_5369,N_2000,N_3653);
nand U5370 (N_5370,N_2077,N_2966);
or U5371 (N_5371,N_3380,N_3276);
nor U5372 (N_5372,N_3559,N_3486);
nor U5373 (N_5373,N_3666,N_2491);
nor U5374 (N_5374,N_2780,N_3692);
xnor U5375 (N_5375,N_3409,N_3255);
xor U5376 (N_5376,N_3187,N_2046);
nor U5377 (N_5377,N_3871,N_2604);
and U5378 (N_5378,N_2556,N_3672);
xnor U5379 (N_5379,N_2040,N_2600);
nor U5380 (N_5380,N_3485,N_3258);
xor U5381 (N_5381,N_2914,N_3382);
nand U5382 (N_5382,N_3545,N_3926);
nand U5383 (N_5383,N_3336,N_2367);
nand U5384 (N_5384,N_3122,N_2751);
or U5385 (N_5385,N_2450,N_3979);
or U5386 (N_5386,N_2552,N_2939);
nand U5387 (N_5387,N_2478,N_3397);
or U5388 (N_5388,N_3034,N_2724);
xor U5389 (N_5389,N_3508,N_3881);
and U5390 (N_5390,N_2546,N_3901);
nor U5391 (N_5391,N_3676,N_2222);
xor U5392 (N_5392,N_2641,N_2093);
nand U5393 (N_5393,N_3849,N_3266);
nand U5394 (N_5394,N_3938,N_2073);
nand U5395 (N_5395,N_2054,N_3181);
and U5396 (N_5396,N_2781,N_2760);
xnor U5397 (N_5397,N_3482,N_2455);
and U5398 (N_5398,N_3844,N_3003);
nand U5399 (N_5399,N_3175,N_3825);
and U5400 (N_5400,N_2169,N_2209);
nand U5401 (N_5401,N_2933,N_3983);
or U5402 (N_5402,N_2123,N_3868);
and U5403 (N_5403,N_3627,N_2205);
or U5404 (N_5404,N_2257,N_3975);
nor U5405 (N_5405,N_3295,N_3894);
nand U5406 (N_5406,N_3795,N_3277);
nor U5407 (N_5407,N_3753,N_2279);
nand U5408 (N_5408,N_3955,N_2110);
xnor U5409 (N_5409,N_2178,N_2283);
xor U5410 (N_5410,N_2099,N_2748);
and U5411 (N_5411,N_3134,N_3249);
or U5412 (N_5412,N_3021,N_2578);
nand U5413 (N_5413,N_2990,N_2695);
or U5414 (N_5414,N_2274,N_2154);
or U5415 (N_5415,N_3295,N_2267);
nor U5416 (N_5416,N_2828,N_3136);
and U5417 (N_5417,N_2488,N_2544);
nand U5418 (N_5418,N_3134,N_2422);
xor U5419 (N_5419,N_2887,N_2344);
and U5420 (N_5420,N_2533,N_3984);
and U5421 (N_5421,N_2483,N_3433);
and U5422 (N_5422,N_2139,N_3315);
nand U5423 (N_5423,N_2626,N_3238);
nor U5424 (N_5424,N_3230,N_3280);
nor U5425 (N_5425,N_2475,N_2109);
and U5426 (N_5426,N_3313,N_3739);
nand U5427 (N_5427,N_3642,N_2233);
nor U5428 (N_5428,N_3675,N_3674);
and U5429 (N_5429,N_2980,N_3688);
or U5430 (N_5430,N_3888,N_3293);
xor U5431 (N_5431,N_3877,N_3259);
or U5432 (N_5432,N_2495,N_2958);
or U5433 (N_5433,N_2574,N_2927);
or U5434 (N_5434,N_3779,N_2640);
and U5435 (N_5435,N_3440,N_2153);
xnor U5436 (N_5436,N_3306,N_2427);
and U5437 (N_5437,N_2716,N_3522);
or U5438 (N_5438,N_2620,N_2239);
nand U5439 (N_5439,N_3913,N_2144);
and U5440 (N_5440,N_3443,N_2615);
and U5441 (N_5441,N_2447,N_2768);
xor U5442 (N_5442,N_2534,N_3047);
and U5443 (N_5443,N_2202,N_3844);
and U5444 (N_5444,N_2859,N_2506);
and U5445 (N_5445,N_3054,N_3808);
and U5446 (N_5446,N_2956,N_2394);
nor U5447 (N_5447,N_2085,N_3410);
or U5448 (N_5448,N_3779,N_2626);
nor U5449 (N_5449,N_2739,N_2920);
or U5450 (N_5450,N_3532,N_3947);
nand U5451 (N_5451,N_3120,N_3194);
nand U5452 (N_5452,N_3030,N_3098);
nand U5453 (N_5453,N_2013,N_2773);
nor U5454 (N_5454,N_3888,N_2267);
xnor U5455 (N_5455,N_3471,N_3029);
nor U5456 (N_5456,N_3176,N_2447);
nand U5457 (N_5457,N_2909,N_2740);
nand U5458 (N_5458,N_3752,N_3490);
nand U5459 (N_5459,N_2544,N_3446);
nand U5460 (N_5460,N_3746,N_2487);
or U5461 (N_5461,N_3623,N_2945);
nor U5462 (N_5462,N_3383,N_2319);
xor U5463 (N_5463,N_3106,N_3039);
or U5464 (N_5464,N_3185,N_3472);
xor U5465 (N_5465,N_2397,N_2781);
or U5466 (N_5466,N_3520,N_2084);
nand U5467 (N_5467,N_2261,N_3845);
and U5468 (N_5468,N_3176,N_2383);
and U5469 (N_5469,N_2164,N_3524);
or U5470 (N_5470,N_3307,N_3959);
nor U5471 (N_5471,N_3023,N_3352);
nor U5472 (N_5472,N_3316,N_2386);
nand U5473 (N_5473,N_2849,N_2157);
xnor U5474 (N_5474,N_3626,N_2705);
and U5475 (N_5475,N_2216,N_3628);
nand U5476 (N_5476,N_3704,N_3574);
nand U5477 (N_5477,N_2708,N_2922);
xor U5478 (N_5478,N_2806,N_2531);
or U5479 (N_5479,N_3259,N_2703);
and U5480 (N_5480,N_3547,N_3481);
nand U5481 (N_5481,N_2783,N_2385);
or U5482 (N_5482,N_2945,N_3491);
nand U5483 (N_5483,N_3642,N_3960);
or U5484 (N_5484,N_2317,N_3270);
xnor U5485 (N_5485,N_2710,N_3225);
nand U5486 (N_5486,N_3010,N_3132);
or U5487 (N_5487,N_3043,N_3615);
xor U5488 (N_5488,N_2835,N_3138);
or U5489 (N_5489,N_3872,N_2153);
and U5490 (N_5490,N_2765,N_3101);
nor U5491 (N_5491,N_2061,N_3446);
xnor U5492 (N_5492,N_2033,N_3549);
nand U5493 (N_5493,N_3205,N_3519);
nor U5494 (N_5494,N_2286,N_3039);
xnor U5495 (N_5495,N_3080,N_3135);
nand U5496 (N_5496,N_3245,N_3846);
nor U5497 (N_5497,N_3518,N_3905);
nor U5498 (N_5498,N_3346,N_3300);
and U5499 (N_5499,N_3002,N_2581);
and U5500 (N_5500,N_2143,N_3587);
and U5501 (N_5501,N_2192,N_2761);
nand U5502 (N_5502,N_2671,N_3465);
nand U5503 (N_5503,N_2999,N_3278);
xnor U5504 (N_5504,N_3065,N_2026);
nand U5505 (N_5505,N_3936,N_3901);
nor U5506 (N_5506,N_2120,N_3224);
nor U5507 (N_5507,N_3129,N_2120);
or U5508 (N_5508,N_3519,N_3001);
and U5509 (N_5509,N_2333,N_2006);
and U5510 (N_5510,N_2730,N_3125);
and U5511 (N_5511,N_2977,N_3641);
xor U5512 (N_5512,N_2027,N_3909);
nand U5513 (N_5513,N_3948,N_3411);
or U5514 (N_5514,N_3115,N_2500);
nand U5515 (N_5515,N_3870,N_2724);
nor U5516 (N_5516,N_2086,N_2864);
xor U5517 (N_5517,N_3625,N_2847);
or U5518 (N_5518,N_3843,N_2757);
xnor U5519 (N_5519,N_3855,N_3424);
xnor U5520 (N_5520,N_2163,N_3661);
and U5521 (N_5521,N_2138,N_2387);
nor U5522 (N_5522,N_2443,N_2748);
and U5523 (N_5523,N_3137,N_2715);
nand U5524 (N_5524,N_2049,N_3560);
and U5525 (N_5525,N_3752,N_2863);
and U5526 (N_5526,N_3200,N_3612);
nand U5527 (N_5527,N_2019,N_2667);
nor U5528 (N_5528,N_3632,N_2729);
xnor U5529 (N_5529,N_2826,N_3761);
nand U5530 (N_5530,N_3173,N_2705);
nand U5531 (N_5531,N_2631,N_3429);
nor U5532 (N_5532,N_2866,N_3477);
nor U5533 (N_5533,N_2710,N_2072);
and U5534 (N_5534,N_3391,N_3076);
and U5535 (N_5535,N_2809,N_3443);
nor U5536 (N_5536,N_2086,N_3860);
nor U5537 (N_5537,N_3568,N_3543);
or U5538 (N_5538,N_2632,N_2363);
nor U5539 (N_5539,N_2043,N_2132);
and U5540 (N_5540,N_3327,N_3616);
or U5541 (N_5541,N_3282,N_3302);
nand U5542 (N_5542,N_3401,N_2548);
nor U5543 (N_5543,N_2442,N_2350);
and U5544 (N_5544,N_2263,N_3802);
nor U5545 (N_5545,N_2165,N_3341);
and U5546 (N_5546,N_2729,N_3517);
nand U5547 (N_5547,N_3236,N_2433);
nor U5548 (N_5548,N_3135,N_3327);
nor U5549 (N_5549,N_2342,N_3478);
nor U5550 (N_5550,N_2311,N_3650);
nor U5551 (N_5551,N_2807,N_3236);
and U5552 (N_5552,N_2417,N_3539);
nor U5553 (N_5553,N_3920,N_2531);
or U5554 (N_5554,N_3634,N_2880);
or U5555 (N_5555,N_3324,N_2201);
nand U5556 (N_5556,N_2824,N_3331);
and U5557 (N_5557,N_3182,N_3341);
and U5558 (N_5558,N_3254,N_2723);
or U5559 (N_5559,N_2647,N_3398);
xnor U5560 (N_5560,N_2483,N_3657);
and U5561 (N_5561,N_3554,N_3427);
or U5562 (N_5562,N_2035,N_3272);
nand U5563 (N_5563,N_2523,N_2204);
nand U5564 (N_5564,N_2235,N_3738);
or U5565 (N_5565,N_3760,N_2621);
xnor U5566 (N_5566,N_3212,N_3975);
nor U5567 (N_5567,N_2128,N_2763);
and U5568 (N_5568,N_2081,N_3853);
nor U5569 (N_5569,N_3143,N_3501);
and U5570 (N_5570,N_3600,N_2656);
nor U5571 (N_5571,N_3954,N_2071);
or U5572 (N_5572,N_2991,N_2170);
xnor U5573 (N_5573,N_2614,N_3468);
and U5574 (N_5574,N_2684,N_3620);
nand U5575 (N_5575,N_2516,N_3117);
and U5576 (N_5576,N_2046,N_3997);
or U5577 (N_5577,N_2479,N_2293);
and U5578 (N_5578,N_2890,N_3880);
or U5579 (N_5579,N_3733,N_3038);
and U5580 (N_5580,N_3967,N_2043);
nor U5581 (N_5581,N_2240,N_2637);
xor U5582 (N_5582,N_3399,N_3473);
nor U5583 (N_5583,N_2741,N_3717);
xnor U5584 (N_5584,N_3594,N_2399);
xnor U5585 (N_5585,N_2206,N_2109);
nor U5586 (N_5586,N_3769,N_3258);
or U5587 (N_5587,N_2001,N_3476);
nand U5588 (N_5588,N_3879,N_3614);
nor U5589 (N_5589,N_2051,N_3213);
nor U5590 (N_5590,N_3405,N_3046);
or U5591 (N_5591,N_2254,N_2233);
or U5592 (N_5592,N_3541,N_3712);
and U5593 (N_5593,N_3059,N_3078);
xnor U5594 (N_5594,N_2440,N_2716);
xor U5595 (N_5595,N_2334,N_3481);
or U5596 (N_5596,N_3639,N_3163);
nand U5597 (N_5597,N_2928,N_3539);
nor U5598 (N_5598,N_3070,N_3639);
or U5599 (N_5599,N_2932,N_2077);
or U5600 (N_5600,N_3359,N_3831);
nand U5601 (N_5601,N_2756,N_3549);
xor U5602 (N_5602,N_3774,N_3473);
or U5603 (N_5603,N_2308,N_3363);
nand U5604 (N_5604,N_2930,N_2035);
and U5605 (N_5605,N_3616,N_3353);
nand U5606 (N_5606,N_2566,N_3058);
or U5607 (N_5607,N_2208,N_2799);
nor U5608 (N_5608,N_2965,N_2595);
xor U5609 (N_5609,N_3001,N_2873);
nor U5610 (N_5610,N_3191,N_2459);
and U5611 (N_5611,N_3476,N_3713);
and U5612 (N_5612,N_2010,N_3221);
nand U5613 (N_5613,N_3832,N_3193);
nand U5614 (N_5614,N_3707,N_3632);
xor U5615 (N_5615,N_3729,N_2018);
or U5616 (N_5616,N_2491,N_2567);
and U5617 (N_5617,N_3831,N_2644);
xor U5618 (N_5618,N_2029,N_2336);
and U5619 (N_5619,N_2131,N_2780);
xor U5620 (N_5620,N_2588,N_2212);
and U5621 (N_5621,N_2517,N_2005);
xor U5622 (N_5622,N_2331,N_2291);
xnor U5623 (N_5623,N_2886,N_3037);
or U5624 (N_5624,N_2742,N_3853);
or U5625 (N_5625,N_3232,N_3792);
nand U5626 (N_5626,N_3372,N_2205);
and U5627 (N_5627,N_2786,N_3271);
xor U5628 (N_5628,N_3063,N_2194);
and U5629 (N_5629,N_3030,N_3443);
xnor U5630 (N_5630,N_2215,N_3808);
xor U5631 (N_5631,N_2507,N_2319);
nand U5632 (N_5632,N_2095,N_2381);
and U5633 (N_5633,N_3024,N_2642);
xor U5634 (N_5634,N_3569,N_3389);
xnor U5635 (N_5635,N_3485,N_3721);
xnor U5636 (N_5636,N_2085,N_3467);
nand U5637 (N_5637,N_3687,N_2977);
xor U5638 (N_5638,N_3767,N_3293);
xnor U5639 (N_5639,N_2362,N_3007);
xor U5640 (N_5640,N_3106,N_2950);
or U5641 (N_5641,N_2936,N_2695);
xor U5642 (N_5642,N_2298,N_2270);
nand U5643 (N_5643,N_3642,N_3873);
nor U5644 (N_5644,N_3483,N_3552);
and U5645 (N_5645,N_3870,N_2797);
and U5646 (N_5646,N_2502,N_2386);
and U5647 (N_5647,N_3791,N_3213);
or U5648 (N_5648,N_3179,N_2191);
nand U5649 (N_5649,N_2410,N_3745);
nor U5650 (N_5650,N_3508,N_3238);
xnor U5651 (N_5651,N_3294,N_2602);
nor U5652 (N_5652,N_3659,N_3286);
nand U5653 (N_5653,N_2675,N_2663);
and U5654 (N_5654,N_2273,N_2353);
nand U5655 (N_5655,N_3374,N_2274);
nor U5656 (N_5656,N_2988,N_2750);
nor U5657 (N_5657,N_3289,N_2053);
nand U5658 (N_5658,N_3898,N_2919);
and U5659 (N_5659,N_3805,N_2772);
nor U5660 (N_5660,N_2708,N_2645);
xnor U5661 (N_5661,N_2954,N_2963);
and U5662 (N_5662,N_2763,N_2915);
xnor U5663 (N_5663,N_2853,N_3226);
nand U5664 (N_5664,N_2464,N_2916);
and U5665 (N_5665,N_2568,N_2483);
xor U5666 (N_5666,N_3129,N_2705);
xor U5667 (N_5667,N_2839,N_3907);
xor U5668 (N_5668,N_3470,N_3777);
nor U5669 (N_5669,N_2863,N_3194);
and U5670 (N_5670,N_3279,N_2577);
nand U5671 (N_5671,N_3707,N_2878);
xor U5672 (N_5672,N_3263,N_2156);
or U5673 (N_5673,N_2498,N_3535);
xor U5674 (N_5674,N_3623,N_3025);
nor U5675 (N_5675,N_3260,N_3219);
nor U5676 (N_5676,N_2288,N_2016);
xor U5677 (N_5677,N_3288,N_2559);
or U5678 (N_5678,N_2382,N_3434);
xnor U5679 (N_5679,N_3325,N_3192);
nor U5680 (N_5680,N_3923,N_2224);
nor U5681 (N_5681,N_2519,N_2437);
nor U5682 (N_5682,N_3952,N_2067);
xor U5683 (N_5683,N_3380,N_2619);
nand U5684 (N_5684,N_3239,N_3943);
nand U5685 (N_5685,N_3065,N_3502);
xor U5686 (N_5686,N_3227,N_3874);
nor U5687 (N_5687,N_2011,N_2890);
nand U5688 (N_5688,N_2900,N_2447);
nor U5689 (N_5689,N_3796,N_3524);
and U5690 (N_5690,N_3813,N_3606);
nand U5691 (N_5691,N_3724,N_2524);
and U5692 (N_5692,N_2734,N_2977);
or U5693 (N_5693,N_3818,N_3595);
and U5694 (N_5694,N_3955,N_3163);
xnor U5695 (N_5695,N_2796,N_3209);
and U5696 (N_5696,N_3765,N_2058);
or U5697 (N_5697,N_2695,N_2295);
xnor U5698 (N_5698,N_2298,N_2174);
and U5699 (N_5699,N_2241,N_2580);
or U5700 (N_5700,N_3564,N_2973);
or U5701 (N_5701,N_2144,N_2462);
xor U5702 (N_5702,N_3470,N_2734);
nand U5703 (N_5703,N_2469,N_2764);
xnor U5704 (N_5704,N_3623,N_3097);
and U5705 (N_5705,N_3909,N_3846);
nand U5706 (N_5706,N_2782,N_2841);
or U5707 (N_5707,N_2155,N_2411);
xnor U5708 (N_5708,N_3054,N_2866);
nor U5709 (N_5709,N_3221,N_2358);
xor U5710 (N_5710,N_3161,N_3327);
xor U5711 (N_5711,N_2921,N_3713);
xor U5712 (N_5712,N_2194,N_3101);
and U5713 (N_5713,N_2340,N_3824);
xnor U5714 (N_5714,N_3152,N_2586);
nand U5715 (N_5715,N_3946,N_2822);
or U5716 (N_5716,N_3258,N_3477);
and U5717 (N_5717,N_3359,N_2240);
xor U5718 (N_5718,N_3037,N_3180);
xor U5719 (N_5719,N_2800,N_2263);
or U5720 (N_5720,N_2153,N_2010);
nand U5721 (N_5721,N_3842,N_3612);
and U5722 (N_5722,N_3226,N_3315);
or U5723 (N_5723,N_3800,N_3765);
nand U5724 (N_5724,N_2394,N_3299);
nor U5725 (N_5725,N_3140,N_2556);
nand U5726 (N_5726,N_3917,N_2346);
nor U5727 (N_5727,N_3346,N_3565);
xnor U5728 (N_5728,N_3787,N_2747);
nand U5729 (N_5729,N_3562,N_3889);
xor U5730 (N_5730,N_3129,N_2110);
nor U5731 (N_5731,N_2879,N_2436);
and U5732 (N_5732,N_3319,N_3187);
nand U5733 (N_5733,N_2664,N_3135);
nand U5734 (N_5734,N_2802,N_3439);
nand U5735 (N_5735,N_2339,N_2979);
nor U5736 (N_5736,N_2383,N_3934);
nand U5737 (N_5737,N_2746,N_2623);
and U5738 (N_5738,N_2610,N_2115);
xor U5739 (N_5739,N_3611,N_2494);
nand U5740 (N_5740,N_2389,N_3020);
or U5741 (N_5741,N_2651,N_3800);
xor U5742 (N_5742,N_3290,N_2210);
and U5743 (N_5743,N_3999,N_3147);
or U5744 (N_5744,N_3370,N_2153);
xor U5745 (N_5745,N_3292,N_2072);
nand U5746 (N_5746,N_2429,N_3161);
and U5747 (N_5747,N_2919,N_3964);
nor U5748 (N_5748,N_3307,N_2251);
nor U5749 (N_5749,N_3314,N_2619);
or U5750 (N_5750,N_3304,N_2590);
nand U5751 (N_5751,N_2546,N_2289);
and U5752 (N_5752,N_3897,N_2052);
or U5753 (N_5753,N_2134,N_3930);
nand U5754 (N_5754,N_2394,N_2000);
or U5755 (N_5755,N_3815,N_2280);
xnor U5756 (N_5756,N_3462,N_3293);
and U5757 (N_5757,N_3177,N_2761);
xor U5758 (N_5758,N_2040,N_2553);
and U5759 (N_5759,N_3955,N_3349);
or U5760 (N_5760,N_2662,N_3348);
nand U5761 (N_5761,N_2065,N_2145);
or U5762 (N_5762,N_2642,N_2845);
and U5763 (N_5763,N_3490,N_3170);
nand U5764 (N_5764,N_2485,N_2145);
nor U5765 (N_5765,N_2930,N_2250);
or U5766 (N_5766,N_2285,N_2880);
nor U5767 (N_5767,N_3707,N_2088);
and U5768 (N_5768,N_3426,N_3066);
or U5769 (N_5769,N_3203,N_2174);
xnor U5770 (N_5770,N_2795,N_2448);
xnor U5771 (N_5771,N_3401,N_3587);
nor U5772 (N_5772,N_2562,N_2503);
nand U5773 (N_5773,N_3841,N_2769);
nor U5774 (N_5774,N_2785,N_2709);
or U5775 (N_5775,N_3368,N_2599);
or U5776 (N_5776,N_3837,N_2605);
or U5777 (N_5777,N_3043,N_2951);
nand U5778 (N_5778,N_3675,N_3898);
nand U5779 (N_5779,N_2878,N_2451);
or U5780 (N_5780,N_2715,N_2269);
nand U5781 (N_5781,N_3113,N_3667);
and U5782 (N_5782,N_3599,N_2505);
nand U5783 (N_5783,N_3771,N_3389);
nand U5784 (N_5784,N_2216,N_2157);
nand U5785 (N_5785,N_3964,N_2606);
and U5786 (N_5786,N_2282,N_2684);
xnor U5787 (N_5787,N_3126,N_3775);
xor U5788 (N_5788,N_3080,N_2528);
nor U5789 (N_5789,N_2249,N_2290);
nor U5790 (N_5790,N_2806,N_2192);
or U5791 (N_5791,N_2586,N_3312);
and U5792 (N_5792,N_2008,N_3079);
and U5793 (N_5793,N_2117,N_2241);
xor U5794 (N_5794,N_2878,N_2655);
nor U5795 (N_5795,N_2730,N_2201);
nor U5796 (N_5796,N_3274,N_3334);
and U5797 (N_5797,N_2467,N_3884);
or U5798 (N_5798,N_3846,N_3815);
xnor U5799 (N_5799,N_3863,N_2554);
nand U5800 (N_5800,N_3568,N_3912);
xor U5801 (N_5801,N_3309,N_3418);
and U5802 (N_5802,N_2712,N_3968);
nor U5803 (N_5803,N_3348,N_3774);
and U5804 (N_5804,N_3198,N_2090);
or U5805 (N_5805,N_2190,N_3645);
and U5806 (N_5806,N_3208,N_2027);
or U5807 (N_5807,N_3090,N_3251);
nor U5808 (N_5808,N_3416,N_2665);
nor U5809 (N_5809,N_2295,N_2867);
and U5810 (N_5810,N_3877,N_3532);
and U5811 (N_5811,N_3198,N_3805);
xor U5812 (N_5812,N_2644,N_2256);
and U5813 (N_5813,N_3933,N_2856);
nand U5814 (N_5814,N_2180,N_3654);
or U5815 (N_5815,N_3333,N_3192);
nor U5816 (N_5816,N_2463,N_3354);
nor U5817 (N_5817,N_3438,N_3984);
xor U5818 (N_5818,N_2139,N_2007);
xor U5819 (N_5819,N_3694,N_3125);
or U5820 (N_5820,N_3621,N_2987);
xnor U5821 (N_5821,N_3783,N_2231);
and U5822 (N_5822,N_3166,N_2573);
nor U5823 (N_5823,N_2623,N_2462);
and U5824 (N_5824,N_3512,N_3761);
xnor U5825 (N_5825,N_2035,N_2349);
xnor U5826 (N_5826,N_2823,N_3325);
nand U5827 (N_5827,N_3482,N_2341);
xor U5828 (N_5828,N_3659,N_3971);
xor U5829 (N_5829,N_3010,N_3098);
and U5830 (N_5830,N_3371,N_3829);
nor U5831 (N_5831,N_2578,N_2855);
or U5832 (N_5832,N_2898,N_3384);
nand U5833 (N_5833,N_2003,N_3187);
and U5834 (N_5834,N_3272,N_2975);
xor U5835 (N_5835,N_3396,N_2654);
nor U5836 (N_5836,N_3440,N_2415);
xor U5837 (N_5837,N_3388,N_3146);
and U5838 (N_5838,N_3135,N_3624);
xor U5839 (N_5839,N_2164,N_2740);
nor U5840 (N_5840,N_2632,N_2522);
xnor U5841 (N_5841,N_3369,N_2043);
nand U5842 (N_5842,N_2420,N_2538);
xor U5843 (N_5843,N_2788,N_3309);
nand U5844 (N_5844,N_2001,N_3077);
xnor U5845 (N_5845,N_3991,N_3157);
nor U5846 (N_5846,N_2358,N_2623);
or U5847 (N_5847,N_3647,N_2278);
nand U5848 (N_5848,N_3664,N_3393);
xnor U5849 (N_5849,N_2863,N_2992);
and U5850 (N_5850,N_2627,N_2397);
nand U5851 (N_5851,N_3864,N_3416);
or U5852 (N_5852,N_2789,N_3802);
or U5853 (N_5853,N_3988,N_2414);
and U5854 (N_5854,N_2324,N_2751);
xor U5855 (N_5855,N_2179,N_3367);
or U5856 (N_5856,N_3365,N_3436);
nor U5857 (N_5857,N_2429,N_2813);
and U5858 (N_5858,N_2182,N_2352);
nor U5859 (N_5859,N_3810,N_2025);
and U5860 (N_5860,N_2356,N_3974);
or U5861 (N_5861,N_3185,N_2546);
xor U5862 (N_5862,N_3030,N_3692);
xor U5863 (N_5863,N_3605,N_2903);
nor U5864 (N_5864,N_2827,N_2131);
or U5865 (N_5865,N_2030,N_2164);
nor U5866 (N_5866,N_3374,N_2086);
xor U5867 (N_5867,N_2439,N_3802);
nand U5868 (N_5868,N_2299,N_3861);
or U5869 (N_5869,N_3215,N_2143);
nand U5870 (N_5870,N_3727,N_2154);
xor U5871 (N_5871,N_2711,N_3013);
nand U5872 (N_5872,N_3800,N_3605);
nand U5873 (N_5873,N_2836,N_2854);
nand U5874 (N_5874,N_2333,N_3597);
xor U5875 (N_5875,N_3706,N_3011);
and U5876 (N_5876,N_2064,N_2108);
and U5877 (N_5877,N_2402,N_2281);
or U5878 (N_5878,N_2038,N_3590);
nand U5879 (N_5879,N_2881,N_2197);
nand U5880 (N_5880,N_3510,N_3206);
nand U5881 (N_5881,N_2475,N_3768);
xnor U5882 (N_5882,N_3527,N_3247);
or U5883 (N_5883,N_3439,N_3356);
or U5884 (N_5884,N_2729,N_2759);
or U5885 (N_5885,N_2775,N_3093);
and U5886 (N_5886,N_3378,N_2673);
and U5887 (N_5887,N_2968,N_2551);
xor U5888 (N_5888,N_3621,N_3077);
and U5889 (N_5889,N_2459,N_2491);
and U5890 (N_5890,N_2324,N_2042);
and U5891 (N_5891,N_2182,N_3643);
nand U5892 (N_5892,N_2159,N_2285);
nand U5893 (N_5893,N_3174,N_2902);
nor U5894 (N_5894,N_3420,N_3350);
nand U5895 (N_5895,N_3280,N_2689);
nand U5896 (N_5896,N_2251,N_2064);
xor U5897 (N_5897,N_3111,N_3449);
and U5898 (N_5898,N_2801,N_3003);
and U5899 (N_5899,N_2168,N_3572);
nand U5900 (N_5900,N_3267,N_3372);
or U5901 (N_5901,N_3477,N_2626);
nor U5902 (N_5902,N_2586,N_3469);
or U5903 (N_5903,N_3994,N_3922);
or U5904 (N_5904,N_2901,N_2767);
nand U5905 (N_5905,N_2181,N_3827);
nand U5906 (N_5906,N_2196,N_2393);
xor U5907 (N_5907,N_3393,N_3614);
nand U5908 (N_5908,N_2580,N_2254);
and U5909 (N_5909,N_3655,N_2100);
or U5910 (N_5910,N_2743,N_2401);
nand U5911 (N_5911,N_3024,N_3550);
nand U5912 (N_5912,N_3344,N_2229);
nand U5913 (N_5913,N_3095,N_3275);
nor U5914 (N_5914,N_2907,N_2952);
xor U5915 (N_5915,N_2523,N_2660);
nor U5916 (N_5916,N_2472,N_2036);
nand U5917 (N_5917,N_2044,N_2986);
and U5918 (N_5918,N_3824,N_2401);
xor U5919 (N_5919,N_3342,N_2498);
xor U5920 (N_5920,N_3720,N_2968);
or U5921 (N_5921,N_3435,N_3451);
xor U5922 (N_5922,N_2999,N_3724);
nand U5923 (N_5923,N_3243,N_2625);
or U5924 (N_5924,N_2321,N_2076);
nand U5925 (N_5925,N_3443,N_3689);
or U5926 (N_5926,N_2358,N_2853);
and U5927 (N_5927,N_3450,N_3321);
nor U5928 (N_5928,N_3720,N_3137);
xnor U5929 (N_5929,N_2352,N_2193);
nand U5930 (N_5930,N_3871,N_3982);
nor U5931 (N_5931,N_3905,N_2399);
and U5932 (N_5932,N_2630,N_2593);
or U5933 (N_5933,N_2439,N_3564);
nand U5934 (N_5934,N_3044,N_3809);
nand U5935 (N_5935,N_2108,N_3230);
or U5936 (N_5936,N_2405,N_3833);
xor U5937 (N_5937,N_2653,N_3409);
xor U5938 (N_5938,N_2897,N_2310);
nor U5939 (N_5939,N_2566,N_2601);
or U5940 (N_5940,N_3655,N_2720);
or U5941 (N_5941,N_3516,N_2977);
or U5942 (N_5942,N_3220,N_3847);
xnor U5943 (N_5943,N_2543,N_3184);
nor U5944 (N_5944,N_2375,N_2002);
xor U5945 (N_5945,N_3043,N_3652);
or U5946 (N_5946,N_3348,N_2438);
xnor U5947 (N_5947,N_2666,N_3507);
or U5948 (N_5948,N_2356,N_2390);
xor U5949 (N_5949,N_3928,N_3938);
nand U5950 (N_5950,N_2776,N_3587);
and U5951 (N_5951,N_2723,N_2742);
xnor U5952 (N_5952,N_2822,N_2328);
or U5953 (N_5953,N_3255,N_2326);
nor U5954 (N_5954,N_3154,N_2136);
nand U5955 (N_5955,N_3035,N_2389);
or U5956 (N_5956,N_2000,N_2696);
nand U5957 (N_5957,N_2037,N_2576);
or U5958 (N_5958,N_2202,N_2695);
or U5959 (N_5959,N_2708,N_2514);
nor U5960 (N_5960,N_3453,N_2695);
nand U5961 (N_5961,N_2455,N_2074);
nand U5962 (N_5962,N_3636,N_3942);
nand U5963 (N_5963,N_3739,N_2062);
nand U5964 (N_5964,N_3145,N_2594);
or U5965 (N_5965,N_2116,N_2510);
and U5966 (N_5966,N_3917,N_2640);
or U5967 (N_5967,N_2972,N_2491);
xnor U5968 (N_5968,N_3232,N_2122);
and U5969 (N_5969,N_3462,N_2268);
nor U5970 (N_5970,N_2933,N_2944);
or U5971 (N_5971,N_2929,N_2861);
nand U5972 (N_5972,N_3066,N_3710);
and U5973 (N_5973,N_3036,N_2548);
or U5974 (N_5974,N_3103,N_2492);
and U5975 (N_5975,N_2403,N_3389);
nor U5976 (N_5976,N_3978,N_3086);
or U5977 (N_5977,N_3574,N_3456);
xnor U5978 (N_5978,N_2621,N_3746);
xor U5979 (N_5979,N_3290,N_3382);
nand U5980 (N_5980,N_2925,N_2691);
or U5981 (N_5981,N_3462,N_3612);
nor U5982 (N_5982,N_3722,N_2251);
nor U5983 (N_5983,N_2530,N_2575);
or U5984 (N_5984,N_2502,N_3081);
nand U5985 (N_5985,N_3871,N_2155);
and U5986 (N_5986,N_2092,N_3077);
nor U5987 (N_5987,N_3220,N_2293);
and U5988 (N_5988,N_3375,N_2740);
and U5989 (N_5989,N_3264,N_2616);
xnor U5990 (N_5990,N_3163,N_2811);
xor U5991 (N_5991,N_3925,N_3864);
or U5992 (N_5992,N_2315,N_2816);
and U5993 (N_5993,N_2819,N_3443);
and U5994 (N_5994,N_3852,N_3139);
and U5995 (N_5995,N_3078,N_3208);
nor U5996 (N_5996,N_3273,N_3185);
nor U5997 (N_5997,N_2401,N_2626);
or U5998 (N_5998,N_2359,N_2587);
and U5999 (N_5999,N_3127,N_2249);
nor U6000 (N_6000,N_5658,N_4380);
or U6001 (N_6001,N_4591,N_5387);
nand U6002 (N_6002,N_4204,N_4556);
and U6003 (N_6003,N_4953,N_5632);
or U6004 (N_6004,N_5721,N_4702);
or U6005 (N_6005,N_4580,N_4922);
nor U6006 (N_6006,N_4816,N_4798);
nand U6007 (N_6007,N_5202,N_4385);
nand U6008 (N_6008,N_4202,N_5532);
xnor U6009 (N_6009,N_5492,N_4085);
nor U6010 (N_6010,N_5230,N_5946);
and U6011 (N_6011,N_4485,N_4075);
and U6012 (N_6012,N_4447,N_5138);
and U6013 (N_6013,N_4043,N_4864);
nor U6014 (N_6014,N_4635,N_4583);
and U6015 (N_6015,N_5649,N_4826);
and U6016 (N_6016,N_5941,N_5173);
or U6017 (N_6017,N_5035,N_4523);
nor U6018 (N_6018,N_4434,N_4531);
or U6019 (N_6019,N_4018,N_4374);
nor U6020 (N_6020,N_5166,N_5309);
or U6021 (N_6021,N_5994,N_5159);
or U6022 (N_6022,N_5084,N_5473);
nand U6023 (N_6023,N_4569,N_5811);
and U6024 (N_6024,N_5080,N_5477);
and U6025 (N_6025,N_5681,N_5813);
and U6026 (N_6026,N_4463,N_5752);
nand U6027 (N_6027,N_4770,N_4733);
nand U6028 (N_6028,N_4909,N_4608);
and U6029 (N_6029,N_4779,N_4517);
and U6030 (N_6030,N_5419,N_5585);
and U6031 (N_6031,N_5075,N_4561);
or U6032 (N_6032,N_5863,N_4326);
or U6033 (N_6033,N_4653,N_4068);
and U6034 (N_6034,N_4592,N_5076);
xnor U6035 (N_6035,N_5133,N_4707);
nor U6036 (N_6036,N_4032,N_4114);
nand U6037 (N_6037,N_4044,N_4851);
and U6038 (N_6038,N_4400,N_5805);
and U6039 (N_6039,N_4247,N_4107);
nor U6040 (N_6040,N_4530,N_4721);
nor U6041 (N_6041,N_4926,N_5100);
nor U6042 (N_6042,N_4141,N_5695);
nand U6043 (N_6043,N_5364,N_4727);
and U6044 (N_6044,N_5136,N_5406);
nand U6045 (N_6045,N_5883,N_4841);
or U6046 (N_6046,N_5229,N_5810);
and U6047 (N_6047,N_5359,N_5090);
and U6048 (N_6048,N_4180,N_4519);
xnor U6049 (N_6049,N_4259,N_4318);
nor U6050 (N_6050,N_4302,N_5693);
xnor U6051 (N_6051,N_4128,N_5451);
and U6052 (N_6052,N_4056,N_5105);
or U6053 (N_6053,N_4263,N_5439);
nand U6054 (N_6054,N_5969,N_4045);
or U6055 (N_6055,N_5302,N_4507);
nor U6056 (N_6056,N_5809,N_5489);
nor U6057 (N_6057,N_4634,N_4740);
xor U6058 (N_6058,N_5029,N_5791);
or U6059 (N_6059,N_5264,N_4737);
nand U6060 (N_6060,N_5245,N_4091);
xor U6061 (N_6061,N_4810,N_5518);
xor U6062 (N_6062,N_5192,N_4459);
xor U6063 (N_6063,N_4039,N_4799);
xnor U6064 (N_6064,N_4551,N_5835);
nand U6065 (N_6065,N_5277,N_5279);
or U6066 (N_6066,N_5360,N_4143);
xnor U6067 (N_6067,N_4852,N_5787);
or U6068 (N_6068,N_5899,N_4418);
and U6069 (N_6069,N_5161,N_4994);
and U6070 (N_6070,N_4613,N_4245);
nand U6071 (N_6071,N_4225,N_5862);
and U6072 (N_6072,N_4422,N_5502);
nor U6073 (N_6073,N_4911,N_5789);
nor U6074 (N_6074,N_5861,N_4682);
xor U6075 (N_6075,N_5276,N_5108);
xor U6076 (N_6076,N_5307,N_5725);
xor U6077 (N_6077,N_4274,N_5400);
or U6078 (N_6078,N_4815,N_5234);
or U6079 (N_6079,N_4771,N_4515);
nand U6080 (N_6080,N_5221,N_5933);
nor U6081 (N_6081,N_4450,N_5280);
xnor U6082 (N_6082,N_5524,N_4562);
or U6083 (N_6083,N_4933,N_5853);
nor U6084 (N_6084,N_4321,N_4865);
and U6085 (N_6085,N_4490,N_4335);
nand U6086 (N_6086,N_5298,N_4837);
nor U6087 (N_6087,N_4488,N_5538);
or U6088 (N_6088,N_5717,N_5475);
nor U6089 (N_6089,N_4630,N_5187);
nand U6090 (N_6090,N_5978,N_5959);
nand U6091 (N_6091,N_4260,N_4236);
and U6092 (N_6092,N_5023,N_4929);
nor U6093 (N_6093,N_4339,N_5579);
and U6094 (N_6094,N_4035,N_5212);
and U6095 (N_6095,N_5513,N_4549);
nand U6096 (N_6096,N_4688,N_4381);
nor U6097 (N_6097,N_4176,N_5416);
nor U6098 (N_6098,N_5860,N_5103);
or U6099 (N_6099,N_5637,N_5461);
or U6100 (N_6100,N_4221,N_5713);
nand U6101 (N_6101,N_5190,N_5252);
or U6102 (N_6102,N_4062,N_5610);
xor U6103 (N_6103,N_4969,N_4522);
nor U6104 (N_6104,N_4252,N_5420);
xor U6105 (N_6105,N_5909,N_5737);
and U6106 (N_6106,N_4642,N_5139);
or U6107 (N_6107,N_4121,N_5736);
and U6108 (N_6108,N_5673,N_5446);
nand U6109 (N_6109,N_5501,N_4391);
nor U6110 (N_6110,N_5609,N_4654);
nand U6111 (N_6111,N_4670,N_4655);
nand U6112 (N_6112,N_5481,N_4430);
or U6113 (N_6113,N_5655,N_4208);
xnor U6114 (N_6114,N_5115,N_4359);
or U6115 (N_6115,N_5907,N_4570);
and U6116 (N_6116,N_5799,N_5879);
or U6117 (N_6117,N_5278,N_5121);
xnor U6118 (N_6118,N_5843,N_4355);
xor U6119 (N_6119,N_4178,N_5095);
and U6120 (N_6120,N_5082,N_4352);
and U6121 (N_6121,N_4006,N_5766);
xor U6122 (N_6122,N_4306,N_5089);
xnor U6123 (N_6123,N_5028,N_4061);
and U6124 (N_6124,N_5623,N_5614);
xnor U6125 (N_6125,N_5816,N_5603);
xnor U6126 (N_6126,N_5218,N_4219);
xnor U6127 (N_6127,N_4340,N_5059);
nand U6128 (N_6128,N_4750,N_5832);
or U6129 (N_6129,N_4965,N_4899);
xnor U6130 (N_6130,N_5025,N_5804);
nand U6131 (N_6131,N_4948,N_5402);
nor U6132 (N_6132,N_4404,N_5060);
xnor U6133 (N_6133,N_5581,N_4500);
xor U6134 (N_6134,N_4917,N_4802);
nand U6135 (N_6135,N_5165,N_5778);
nand U6136 (N_6136,N_4298,N_5346);
xnor U6137 (N_6137,N_5859,N_4297);
and U6138 (N_6138,N_5846,N_4597);
nand U6139 (N_6139,N_4330,N_5898);
or U6140 (N_6140,N_5668,N_4262);
xor U6141 (N_6141,N_4593,N_4610);
xnor U6142 (N_6142,N_5543,N_4902);
nand U6143 (N_6143,N_5185,N_5742);
xor U6144 (N_6144,N_4257,N_5085);
or U6145 (N_6145,N_4809,N_5203);
or U6146 (N_6146,N_4543,N_5345);
or U6147 (N_6147,N_5018,N_5246);
nor U6148 (N_6148,N_4441,N_5908);
xor U6149 (N_6149,N_4557,N_5504);
or U6150 (N_6150,N_5304,N_4784);
xor U6151 (N_6151,N_5901,N_5850);
and U6152 (N_6152,N_5453,N_4310);
and U6153 (N_6153,N_4130,N_5892);
or U6154 (N_6154,N_4416,N_4405);
nor U6155 (N_6155,N_4331,N_5236);
nor U6156 (N_6156,N_5485,N_4712);
nor U6157 (N_6157,N_4907,N_5378);
nand U6158 (N_6158,N_5064,N_5775);
nor U6159 (N_6159,N_4442,N_4454);
and U6160 (N_6160,N_4206,N_5339);
and U6161 (N_6161,N_5282,N_4234);
xor U6162 (N_6162,N_4883,N_4836);
and U6163 (N_6163,N_4590,N_4753);
or U6164 (N_6164,N_4898,N_4487);
or U6165 (N_6165,N_4726,N_4859);
xnor U6166 (N_6166,N_4893,N_5071);
or U6167 (N_6167,N_4240,N_4084);
and U6168 (N_6168,N_4144,N_4065);
nand U6169 (N_6169,N_4042,N_5594);
and U6170 (N_6170,N_5716,N_5956);
and U6171 (N_6171,N_5865,N_5993);
nand U6172 (N_6172,N_4586,N_4066);
nand U6173 (N_6173,N_5448,N_5338);
nand U6174 (N_6174,N_4364,N_5949);
nand U6175 (N_6175,N_5318,N_5176);
nor U6176 (N_6176,N_4333,N_4376);
nor U6177 (N_6177,N_5315,N_4518);
or U6178 (N_6178,N_5327,N_4276);
or U6179 (N_6179,N_5821,N_5251);
or U6180 (N_6180,N_5456,N_5152);
and U6181 (N_6181,N_4256,N_4289);
or U6182 (N_6182,N_5967,N_5938);
or U6183 (N_6183,N_5174,N_4021);
or U6184 (N_6184,N_4429,N_4460);
and U6185 (N_6185,N_4271,N_4249);
and U6186 (N_6186,N_4956,N_5091);
nand U6187 (N_6187,N_5881,N_5828);
xor U6188 (N_6188,N_5094,N_4356);
nand U6189 (N_6189,N_5217,N_4278);
or U6190 (N_6190,N_5694,N_5773);
xnor U6191 (N_6191,N_5321,N_4217);
xor U6192 (N_6192,N_5690,N_5559);
xnor U6193 (N_6193,N_4981,N_5914);
or U6194 (N_6194,N_4897,N_4366);
nor U6195 (N_6195,N_4226,N_5033);
or U6196 (N_6196,N_4976,N_4351);
nand U6197 (N_6197,N_5684,N_5534);
and U6198 (N_6198,N_4623,N_5476);
or U6199 (N_6199,N_4197,N_5873);
nor U6200 (N_6200,N_5560,N_4011);
nand U6201 (N_6201,N_5745,N_4272);
xor U6202 (N_6202,N_4511,N_5348);
and U6203 (N_6203,N_5397,N_5488);
and U6204 (N_6204,N_5388,N_4057);
nor U6205 (N_6205,N_4343,N_5718);
nand U6206 (N_6206,N_5535,N_5353);
xnor U6207 (N_6207,N_4076,N_5126);
nand U6208 (N_6208,N_5039,N_5744);
xor U6209 (N_6209,N_4058,N_4193);
nor U6210 (N_6210,N_4906,N_5047);
or U6211 (N_6211,N_4679,N_5659);
and U6212 (N_6212,N_5548,N_4329);
nor U6213 (N_6213,N_5068,N_4819);
and U6214 (N_6214,N_5206,N_4509);
nor U6215 (N_6215,N_4703,N_5827);
or U6216 (N_6216,N_4891,N_5552);
and U6217 (N_6217,N_5641,N_5983);
or U6218 (N_6218,N_5057,N_4394);
nand U6219 (N_6219,N_4473,N_4269);
or U6220 (N_6220,N_5072,N_5630);
nand U6221 (N_6221,N_5757,N_5436);
nor U6222 (N_6222,N_5177,N_4150);
nand U6223 (N_6223,N_5750,N_5463);
and U6224 (N_6224,N_5670,N_4233);
xnor U6225 (N_6225,N_4002,N_5242);
and U6226 (N_6226,N_5045,N_5031);
xnor U6227 (N_6227,N_5925,N_4393);
xnor U6228 (N_6228,N_4083,N_4827);
nor U6229 (N_6229,N_5553,N_5010);
xor U6230 (N_6230,N_5733,N_4480);
xnor U6231 (N_6231,N_4714,N_4413);
and U6232 (N_6232,N_5458,N_5297);
or U6233 (N_6233,N_4110,N_4535);
and U6234 (N_6234,N_4573,N_5927);
and U6235 (N_6235,N_5871,N_4311);
or U6236 (N_6236,N_4942,N_5970);
or U6237 (N_6237,N_4617,N_5478);
xnor U6238 (N_6238,N_4506,N_5947);
xnor U6239 (N_6239,N_4415,N_5022);
and U6240 (N_6240,N_5760,N_5329);
nand U6241 (N_6241,N_4754,N_5558);
nand U6242 (N_6242,N_5429,N_5496);
nand U6243 (N_6243,N_5920,N_5261);
xor U6244 (N_6244,N_4175,N_5564);
xor U6245 (N_6245,N_4315,N_4761);
or U6246 (N_6246,N_5196,N_4451);
and U6247 (N_6247,N_5851,N_4345);
or U6248 (N_6248,N_4533,N_5688);
and U6249 (N_6249,N_5584,N_4123);
nand U6250 (N_6250,N_5888,N_4813);
nand U6251 (N_6251,N_5830,N_5870);
or U6252 (N_6252,N_4466,N_5512);
xor U6253 (N_6253,N_4763,N_4181);
or U6254 (N_6254,N_5132,N_5770);
nor U6255 (N_6255,N_4805,N_4191);
xor U6256 (N_6256,N_5957,N_5923);
and U6257 (N_6257,N_5296,N_5714);
nor U6258 (N_6258,N_4769,N_4677);
nor U6259 (N_6259,N_4882,N_4694);
nand U6260 (N_6260,N_5749,N_4401);
nand U6261 (N_6261,N_4860,N_5195);
or U6262 (N_6262,N_5286,N_5563);
and U6263 (N_6263,N_5320,N_4885);
xnor U6264 (N_6264,N_4894,N_5437);
nor U6265 (N_6265,N_5454,N_5991);
nor U6266 (N_6266,N_4713,N_5213);
or U6267 (N_6267,N_5066,N_5743);
nor U6268 (N_6268,N_5118,N_5131);
nor U6269 (N_6269,N_4382,N_5178);
and U6270 (N_6270,N_5671,N_4800);
and U6271 (N_6271,N_5772,N_4698);
and U6272 (N_6272,N_5274,N_4649);
xor U6273 (N_6273,N_5367,N_4986);
and U6274 (N_6274,N_5113,N_5288);
and U6275 (N_6275,N_4720,N_5792);
and U6276 (N_6276,N_4681,N_4879);
or U6277 (N_6277,N_5249,N_4973);
nor U6278 (N_6278,N_5875,N_4495);
and U6279 (N_6279,N_4532,N_5571);
and U6280 (N_6280,N_5876,N_4288);
and U6281 (N_6281,N_5989,N_4790);
nand U6282 (N_6282,N_5506,N_5998);
nor U6283 (N_6283,N_5435,N_5273);
nand U6284 (N_6284,N_4555,N_5644);
nor U6285 (N_6285,N_4453,N_5308);
and U6286 (N_6286,N_5423,N_5052);
or U6287 (N_6287,N_5299,N_5682);
and U6288 (N_6288,N_5974,N_4088);
and U6289 (N_6289,N_4216,N_4829);
xor U6290 (N_6290,N_4054,N_4692);
nor U6291 (N_6291,N_5697,N_5602);
nor U6292 (N_6292,N_5394,N_5629);
or U6293 (N_6293,N_5497,N_5699);
nor U6294 (N_6294,N_5017,N_4468);
nand U6295 (N_6295,N_4748,N_5490);
nand U6296 (N_6296,N_4873,N_5884);
nand U6297 (N_6297,N_5472,N_4647);
or U6298 (N_6298,N_5040,N_5164);
nor U6299 (N_6299,N_4470,N_5233);
and U6300 (N_6300,N_4818,N_4398);
and U6301 (N_6301,N_4735,N_5369);
xor U6302 (N_6302,N_5767,N_4215);
nand U6303 (N_6303,N_5326,N_4988);
xor U6304 (N_6304,N_5676,N_5445);
xnor U6305 (N_6305,N_4605,N_4938);
xor U6306 (N_6306,N_4200,N_4205);
and U6307 (N_6307,N_4270,N_4987);
nand U6308 (N_6308,N_4697,N_5328);
or U6309 (N_6309,N_4086,N_5114);
and U6310 (N_6310,N_4063,N_5723);
xnor U6311 (N_6311,N_4001,N_5536);
xnor U6312 (N_6312,N_5844,N_4772);
and U6313 (N_6313,N_5486,N_5070);
nand U6314 (N_6314,N_5911,N_4918);
nor U6315 (N_6315,N_5250,N_4105);
and U6316 (N_6316,N_5146,N_4547);
and U6317 (N_6317,N_4845,N_4833);
nand U6318 (N_6318,N_4629,N_4164);
or U6319 (N_6319,N_4069,N_5526);
or U6320 (N_6320,N_5036,N_4149);
nand U6321 (N_6321,N_4627,N_5205);
nand U6322 (N_6322,N_4683,N_5839);
or U6323 (N_6323,N_5209,N_5452);
nand U6324 (N_6324,N_5396,N_5573);
nand U6325 (N_6325,N_4253,N_5626);
nor U6326 (N_6326,N_4999,N_5223);
nor U6327 (N_6327,N_4529,N_5739);
nor U6328 (N_6328,N_4636,N_4241);
nand U6329 (N_6329,N_4528,N_4040);
xnor U6330 (N_6330,N_5984,N_5729);
or U6331 (N_6331,N_5724,N_5365);
and U6332 (N_6332,N_4187,N_5568);
nor U6333 (N_6333,N_4975,N_5459);
nor U6334 (N_6334,N_4758,N_4477);
xnor U6335 (N_6335,N_5395,N_5952);
nand U6336 (N_6336,N_5426,N_5499);
nor U6337 (N_6337,N_4546,N_4541);
or U6338 (N_6338,N_4407,N_4751);
nand U6339 (N_6339,N_5924,N_5399);
nand U6340 (N_6340,N_5283,N_5539);
xnor U6341 (N_6341,N_4525,N_4337);
xor U6342 (N_6342,N_4675,N_4194);
and U6343 (N_6343,N_4534,N_5981);
xor U6344 (N_6344,N_4765,N_4138);
or U6345 (N_6345,N_5352,N_4777);
and U6346 (N_6346,N_4478,N_5702);
nor U6347 (N_6347,N_4139,N_5913);
xnor U6348 (N_6348,N_5817,N_5508);
nor U6349 (N_6349,N_5030,N_4632);
xnor U6350 (N_6350,N_4266,N_4725);
or U6351 (N_6351,N_5631,N_5333);
xor U6352 (N_6352,N_5265,N_5134);
and U6353 (N_6353,N_5323,N_5712);
and U6354 (N_6354,N_5520,N_4250);
nand U6355 (N_6355,N_5374,N_4280);
nor U6356 (N_6356,N_4710,N_4255);
and U6357 (N_6357,N_5407,N_5516);
or U6358 (N_6358,N_5301,N_4379);
nand U6359 (N_6359,N_5878,N_5701);
nand U6360 (N_6360,N_5886,N_5119);
nand U6361 (N_6361,N_4700,N_4465);
nor U6362 (N_6362,N_5825,N_5386);
nand U6363 (N_6363,N_5596,N_5601);
nand U6364 (N_6364,N_5608,N_4844);
nand U6365 (N_6365,N_5042,N_5484);
or U6366 (N_6366,N_5565,N_5800);
nor U6367 (N_6367,N_5410,N_5300);
or U6368 (N_6368,N_4157,N_5127);
or U6369 (N_6369,N_4027,N_4611);
xor U6370 (N_6370,N_5027,N_5618);
xnor U6371 (N_6371,N_4439,N_4475);
or U6372 (N_6372,N_5592,N_5376);
and U6373 (N_6373,N_4974,N_4734);
and U6374 (N_6374,N_5430,N_4552);
and U6375 (N_6375,N_5709,N_4984);
and U6376 (N_6376,N_5877,N_4145);
and U6377 (N_6377,N_4730,N_4585);
nor U6378 (N_6378,N_5487,N_5021);
or U6379 (N_6379,N_5026,N_4009);
nand U6380 (N_6380,N_4195,N_5557);
or U6381 (N_6381,N_5549,N_5403);
nor U6382 (N_6382,N_5305,N_4186);
xnor U6383 (N_6383,N_4888,N_4448);
nor U6384 (N_6384,N_4743,N_5551);
and U6385 (N_6385,N_4034,N_4210);
xor U6386 (N_6386,N_5193,N_5428);
nand U6387 (N_6387,N_5505,N_4952);
and U6388 (N_6388,N_5793,N_5211);
and U6389 (N_6389,N_4689,N_5143);
or U6390 (N_6390,N_4967,N_4571);
or U6391 (N_6391,N_5855,N_4936);
nor U6392 (N_6392,N_4866,N_5689);
nor U6393 (N_6393,N_5015,N_5016);
and U6394 (N_6394,N_5857,N_5613);
and U6395 (N_6395,N_5527,N_4457);
nand U6396 (N_6396,N_4308,N_5104);
nor U6397 (N_6397,N_5838,N_4626);
and U6398 (N_6398,N_4174,N_4410);
or U6399 (N_6399,N_4196,N_4395);
nand U6400 (N_6400,N_5053,N_5183);
or U6401 (N_6401,N_4294,N_4370);
xor U6402 (N_6402,N_5275,N_4954);
nor U6403 (N_6403,N_4317,N_5916);
nor U6404 (N_6404,N_5995,N_5652);
or U6405 (N_6405,N_4872,N_5208);
nand U6406 (N_6406,N_5657,N_4991);
or U6407 (N_6407,N_4417,N_4334);
nor U6408 (N_6408,N_5096,N_4505);
and U6409 (N_6409,N_5986,N_5814);
and U6410 (N_6410,N_5591,N_4628);
or U6411 (N_6411,N_5093,N_5281);
and U6412 (N_6412,N_5703,N_4461);
nor U6413 (N_6413,N_5337,N_4959);
xnor U6414 (N_6414,N_4868,N_5331);
or U6415 (N_6415,N_4875,N_4792);
or U6416 (N_6416,N_5482,N_5184);
nand U6417 (N_6417,N_4773,N_4222);
or U6418 (N_6418,N_4961,N_5172);
nor U6419 (N_6419,N_5316,N_5541);
nand U6420 (N_6420,N_4133,N_4668);
nor U6421 (N_6421,N_4612,N_4237);
nor U6422 (N_6422,N_5985,N_5171);
nand U6423 (N_6423,N_4576,N_5124);
or U6424 (N_6424,N_5322,N_4619);
and U6425 (N_6425,N_4855,N_5795);
nand U6426 (N_6426,N_4674,N_5580);
xnor U6427 (N_6427,N_4966,N_5444);
nor U6428 (N_6428,N_4427,N_4440);
xor U6429 (N_6429,N_4172,N_4097);
and U6430 (N_6430,N_5141,N_4299);
and U6431 (N_6431,N_4614,N_4838);
and U6432 (N_6432,N_5401,N_4745);
and U6433 (N_6433,N_5806,N_4137);
and U6434 (N_6434,N_4971,N_4687);
nand U6435 (N_6435,N_5756,N_5902);
xor U6436 (N_6436,N_4680,N_4168);
nand U6437 (N_6437,N_5291,N_4804);
nor U6438 (N_6438,N_5140,N_4502);
xnor U6439 (N_6439,N_5041,N_4695);
xnor U6440 (N_6440,N_4747,N_5646);
xnor U6441 (N_6441,N_4760,N_4645);
or U6442 (N_6442,N_4584,N_5829);
nor U6443 (N_6443,N_4484,N_4286);
nand U6444 (N_6444,N_4831,N_5882);
and U6445 (N_6445,N_4048,N_4052);
nand U6446 (N_6446,N_4101,N_4708);
nand U6447 (N_6447,N_4169,N_4323);
and U6448 (N_6448,N_5120,N_5932);
xnor U6449 (N_6449,N_4793,N_5145);
nand U6450 (N_6450,N_5762,N_4412);
xor U6451 (N_6451,N_5255,N_4915);
xor U6452 (N_6452,N_5332,N_5162);
and U6453 (N_6453,N_5889,N_4029);
nor U6454 (N_6454,N_5024,N_4977);
xnor U6455 (N_6455,N_5706,N_4079);
or U6456 (N_6456,N_5988,N_4111);
xor U6457 (N_6457,N_4741,N_4017);
nand U6458 (N_6458,N_5272,N_4671);
xnor U6459 (N_6459,N_5929,N_5928);
nand U6460 (N_6460,N_4661,N_4055);
nor U6461 (N_6461,N_5607,N_4498);
nor U6462 (N_6462,N_4100,N_4738);
xnor U6463 (N_6463,N_4408,N_5460);
nand U6464 (N_6464,N_5639,N_4167);
nor U6465 (N_6465,N_4213,N_5577);
nor U6466 (N_6466,N_4947,N_5599);
or U6467 (N_6467,N_5008,N_4098);
and U6468 (N_6468,N_4823,N_5605);
xor U6469 (N_6469,N_4824,N_5392);
nor U6470 (N_6470,N_4663,N_4696);
and U6471 (N_6471,N_4438,N_5554);
and U6472 (N_6472,N_5013,N_5434);
nand U6473 (N_6473,N_4122,N_4349);
nand U6474 (N_6474,N_5540,N_4968);
xnor U6475 (N_6475,N_5294,N_4154);
nor U6476 (N_6476,N_4676,N_5960);
nand U6477 (N_6477,N_5874,N_4115);
nand U6478 (N_6478,N_4458,N_5848);
xnor U6479 (N_6479,N_4625,N_4047);
nor U6480 (N_6480,N_5635,N_4578);
nor U6481 (N_6481,N_5958,N_5412);
nand U6482 (N_6482,N_4667,N_4113);
nor U6483 (N_6483,N_4419,N_4443);
nand U6484 (N_6484,N_4600,N_4296);
or U6485 (N_6485,N_4732,N_5720);
nor U6486 (N_6486,N_5836,N_5731);
xor U6487 (N_6487,N_5285,N_5771);
or U6488 (N_6488,N_5917,N_4828);
nor U6489 (N_6489,N_4426,N_5621);
xnor U6490 (N_6490,N_4397,N_4548);
and U6491 (N_6491,N_4637,N_4080);
xnor U6492 (N_6492,N_4820,N_5740);
xor U6493 (N_6493,N_5842,N_5390);
and U6494 (N_6494,N_5764,N_4471);
xor U6495 (N_6495,N_5144,N_4151);
nor U6496 (N_6496,N_4706,N_4716);
nand U6497 (N_6497,N_5674,N_5169);
nand U6498 (N_6498,N_5111,N_4096);
xnor U6499 (N_6499,N_5200,N_5783);
or U6500 (N_6500,N_4267,N_5625);
nand U6501 (N_6501,N_4540,N_4010);
nand U6502 (N_6502,N_5616,N_5663);
or U6503 (N_6503,N_4136,N_5081);
nor U6504 (N_6504,N_4003,N_4643);
xnor U6505 (N_6505,N_5046,N_4633);
or U6506 (N_6506,N_5759,N_5732);
or U6507 (N_6507,N_4449,N_5313);
or U6508 (N_6508,N_4783,N_4327);
or U6509 (N_6509,N_5334,N_5191);
and U6510 (N_6510,N_4863,N_5887);
or U6511 (N_6511,N_5785,N_4701);
and U6512 (N_6512,N_5826,N_4007);
nand U6513 (N_6513,N_4858,N_4558);
xor U6514 (N_6514,N_4300,N_4207);
xnor U6515 (N_6515,N_4261,N_4658);
and U6516 (N_6516,N_4705,N_5224);
xor U6517 (N_6517,N_5550,N_4962);
nor U6518 (N_6518,N_5263,N_5244);
and U6519 (N_6519,N_4589,N_4344);
nand U6520 (N_6520,N_4067,N_5248);
xor U6521 (N_6521,N_4749,N_5831);
or U6522 (N_6522,N_5225,N_4126);
and U6523 (N_6523,N_4389,N_4757);
nand U6524 (N_6524,N_5897,N_4423);
nand U6525 (N_6525,N_5798,N_5455);
or U6526 (N_6526,N_5465,N_4078);
or U6527 (N_6527,N_5530,N_4943);
nand U6528 (N_6528,N_5683,N_4527);
nand U6529 (N_6529,N_4112,N_5471);
or U6530 (N_6530,N_5295,N_4941);
and U6531 (N_6531,N_4014,N_4153);
and U6532 (N_6532,N_5253,N_4104);
xnor U6533 (N_6533,N_4744,N_5201);
xnor U6534 (N_6534,N_4989,N_4539);
or U6535 (N_6535,N_4163,N_5382);
and U6536 (N_6536,N_5112,N_5562);
xnor U6537 (N_6537,N_5915,N_4847);
nor U6538 (N_6538,N_4566,N_5758);
and U6539 (N_6539,N_5698,N_4762);
nor U6540 (N_6540,N_4092,N_4788);
or U6541 (N_6541,N_4303,N_5566);
nor U6542 (N_6542,N_4232,N_5306);
xnor U6543 (N_6543,N_4949,N_4012);
nor U6544 (N_6544,N_5715,N_4718);
xnor U6545 (N_6545,N_4903,N_5678);
nand U6546 (N_6546,N_4189,N_4103);
nor U6547 (N_6547,N_5355,N_5470);
xnor U6548 (N_6548,N_4910,N_4806);
or U6549 (N_6549,N_5587,N_5801);
and U6550 (N_6550,N_4409,N_5198);
or U6551 (N_6551,N_5950,N_4158);
xnor U6552 (N_6552,N_5239,N_4752);
xor U6553 (N_6553,N_4684,N_4579);
nor U6554 (N_6554,N_5968,N_5340);
and U6555 (N_6555,N_5727,N_5619);
or U6556 (N_6556,N_5377,N_5935);
xor U6557 (N_6557,N_5393,N_4399);
nor U6558 (N_6558,N_5708,N_5074);
and U6559 (N_6559,N_5357,N_4287);
nand U6560 (N_6560,N_5647,N_5002);
nand U6561 (N_6561,N_5680,N_4870);
nor U6562 (N_6562,N_4901,N_4588);
or U6563 (N_6563,N_5356,N_4406);
or U6564 (N_6564,N_4281,N_5219);
nand U6565 (N_6565,N_4774,N_5312);
or U6566 (N_6566,N_5617,N_4446);
nor U6567 (N_6567,N_4550,N_5819);
nor U6568 (N_6568,N_5310,N_5834);
xor U6569 (N_6569,N_5354,N_5414);
xor U6570 (N_6570,N_4129,N_4537);
xnor U6571 (N_6571,N_5181,N_5411);
xor U6572 (N_6572,N_4433,N_5254);
nor U6573 (N_6573,N_5362,N_5058);
and U6574 (N_6574,N_4188,N_4147);
xnor U6575 (N_6575,N_5123,N_4292);
and U6576 (N_6576,N_4324,N_4731);
or U6577 (N_6577,N_5292,N_4336);
nand U6578 (N_6578,N_5624,N_5578);
xnor U6579 (N_6579,N_5197,N_5687);
nand U6580 (N_6580,N_4884,N_5421);
and U6581 (N_6581,N_4814,N_5235);
and U6582 (N_6582,N_5438,N_4979);
nand U6583 (N_6583,N_5077,N_4646);
nand U6584 (N_6584,N_5383,N_4290);
xnor U6585 (N_6585,N_5593,N_5073);
or U6586 (N_6586,N_5856,N_5086);
nor U6587 (N_6587,N_5228,N_5044);
and U6588 (N_6588,N_5556,N_4026);
and U6589 (N_6589,N_4031,N_4019);
nor U6590 (N_6590,N_5336,N_5262);
nor U6591 (N_6591,N_5510,N_4691);
xor U6592 (N_6592,N_5885,N_5427);
xnor U6593 (N_6593,N_5479,N_4265);
or U6594 (N_6594,N_4890,N_5906);
nand U6595 (N_6595,N_4786,N_5433);
nand U6596 (N_6596,N_5943,N_5271);
and U6597 (N_6597,N_5638,N_5665);
nand U6598 (N_6598,N_4644,N_4620);
and U6599 (N_6599,N_5269,N_5586);
xnor U6600 (N_6600,N_5468,N_5738);
or U6601 (N_6601,N_5576,N_5953);
nor U6602 (N_6602,N_4669,N_4998);
xnor U6603 (N_6603,N_4504,N_5361);
xor U6604 (N_6604,N_4889,N_5858);
and U6605 (N_6605,N_5589,N_5645);
nor U6606 (N_6606,N_4483,N_5975);
nand U6607 (N_6607,N_5944,N_4420);
xnor U6608 (N_6608,N_4024,N_5845);
nor U6609 (N_6609,N_5755,N_4319);
and U6610 (N_6610,N_5006,N_4095);
nor U6611 (N_6611,N_4955,N_4652);
xor U6612 (N_6612,N_4223,N_5777);
nand U6613 (N_6613,N_4717,N_5818);
xor U6614 (N_6614,N_5570,N_4782);
and U6615 (N_6615,N_5011,N_4880);
nor U6616 (N_6616,N_5188,N_5964);
nor U6617 (N_6617,N_4709,N_5866);
nand U6618 (N_6618,N_5852,N_4070);
nand U6619 (N_6619,N_5371,N_5754);
xnor U6620 (N_6620,N_5005,N_4332);
nor U6621 (N_6621,N_4607,N_5544);
xnor U6622 (N_6622,N_5168,N_5867);
and U6623 (N_6623,N_5664,N_4120);
nor U6624 (N_6624,N_4134,N_5824);
nand U6625 (N_6625,N_4008,N_4462);
xor U6626 (N_6626,N_5175,N_5432);
or U6627 (N_6627,N_4514,N_5519);
nor U6628 (N_6628,N_4742,N_5149);
xnor U6629 (N_6629,N_5786,N_4985);
nor U6630 (N_6630,N_5317,N_4609);
nand U6631 (N_6631,N_5065,N_5533);
or U6632 (N_6632,N_5156,N_5598);
nor U6633 (N_6633,N_4375,N_4131);
nor U6634 (N_6634,N_4524,N_5768);
xnor U6635 (N_6635,N_4028,N_4492);
nand U6636 (N_6636,N_4900,N_5779);
xor U6637 (N_6637,N_5335,N_5686);
nor U6638 (N_6638,N_4924,N_5803);
nand U6639 (N_6639,N_4821,N_5097);
nor U6640 (N_6640,N_5375,N_4854);
nor U6641 (N_6641,N_5128,N_5256);
or U6642 (N_6642,N_4445,N_4560);
nor U6643 (N_6643,N_4074,N_5270);
nand U6644 (N_6644,N_4361,N_5934);
nor U6645 (N_6645,N_4279,N_4768);
xnor U6646 (N_6646,N_5521,N_5366);
xnor U6647 (N_6647,N_5972,N_5194);
and U6648 (N_6648,N_4246,N_4925);
nor U6649 (N_6649,N_4251,N_4273);
nand U6650 (N_6650,N_4574,N_5424);
and U6651 (N_6651,N_5525,N_5158);
nor U6652 (N_6652,N_5973,N_5350);
nand U6653 (N_6653,N_5088,N_5186);
xor U6654 (N_6654,N_5034,N_5636);
and U6655 (N_6655,N_4624,N_4963);
nor U6656 (N_6656,N_4230,N_5214);
xnor U6657 (N_6657,N_5822,N_4049);
and U6658 (N_6658,N_4102,N_5293);
and U6659 (N_6659,N_5961,N_5268);
xor U6660 (N_6660,N_4931,N_5780);
or U6661 (N_6661,N_4722,N_4358);
and U6662 (N_6662,N_5373,N_5627);
or U6663 (N_6663,N_5849,N_4639);
xor U6664 (N_6664,N_4807,N_4803);
or U6665 (N_6665,N_4199,N_4595);
and U6666 (N_6666,N_4723,N_4467);
xor U6667 (N_6667,N_5125,N_5815);
nand U6668 (N_6668,N_4958,N_5951);
nand U6669 (N_6669,N_4384,N_5153);
nand U6670 (N_6670,N_4372,N_4161);
xor U6671 (N_6671,N_4797,N_4817);
nor U6672 (N_6672,N_4565,N_4939);
and U6673 (N_6673,N_4444,N_5370);
or U6674 (N_6674,N_4914,N_4436);
nand U6675 (N_6675,N_4293,N_4839);
and U6676 (N_6676,N_4037,N_5155);
xor U6677 (N_6677,N_4602,N_4160);
xnor U6678 (N_6678,N_4563,N_5467);
nor U6679 (N_6679,N_5669,N_5311);
xor U6680 (N_6680,N_4497,N_5893);
xnor U6681 (N_6681,N_4089,N_4390);
nor U6682 (N_6682,N_5147,N_5936);
nor U6683 (N_6683,N_4673,N_4437);
and U6684 (N_6684,N_4386,N_5287);
or U6685 (N_6685,N_5231,N_4020);
xnor U6686 (N_6686,N_5660,N_4756);
or U6687 (N_6687,N_4455,N_5531);
and U6688 (N_6688,N_4598,N_4935);
nor U6689 (N_6689,N_4135,N_5963);
and U6690 (N_6690,N_5150,N_5794);
xnor U6691 (N_6691,N_4767,N_4489);
nor U6692 (N_6692,N_4140,N_5199);
nand U6693 (N_6693,N_5137,N_5606);
nor U6694 (N_6694,N_5784,N_5880);
or U6695 (N_6695,N_4544,N_4657);
or U6696 (N_6696,N_5157,N_5368);
nand U6697 (N_6697,N_4496,N_5457);
nand U6698 (N_6698,N_5494,N_5257);
nand U6699 (N_6699,N_5009,N_4360);
nand U6700 (N_6700,N_4229,N_5389);
xor U6701 (N_6701,N_4621,N_4951);
and U6702 (N_6702,N_5284,N_5869);
xnor U6703 (N_6703,N_5384,N_5163);
and U6704 (N_6704,N_4313,N_5450);
xor U6705 (N_6705,N_4690,N_4932);
and U6706 (N_6706,N_4403,N_4218);
or U6707 (N_6707,N_5349,N_5449);
nor U6708 (N_6708,N_4736,N_4728);
xor U6709 (N_6709,N_5003,N_5904);
xor U6710 (N_6710,N_4764,N_4822);
nand U6711 (N_6711,N_5769,N_5634);
nor U6712 (N_6712,N_4980,N_4004);
or U6713 (N_6713,N_5447,N_4796);
or U6714 (N_6714,N_4108,N_5788);
xnor U6715 (N_6715,N_5344,N_4481);
nand U6716 (N_6716,N_5215,N_4377);
or U6717 (N_6717,N_5700,N_5987);
and U6718 (N_6718,N_5722,N_5507);
or U6719 (N_6719,N_5921,N_5474);
nand U6720 (N_6720,N_4913,N_5528);
nand U6721 (N_6721,N_5314,N_4493);
xnor U6722 (N_6722,N_4997,N_4542);
or U6723 (N_6723,N_4388,N_5980);
nand U6724 (N_6724,N_5661,N_5032);
nand U6725 (N_6725,N_4789,N_4755);
nand U6726 (N_6726,N_5640,N_4046);
or U6727 (N_6727,N_4059,N_4957);
and U6728 (N_6728,N_4711,N_4378);
nand U6729 (N_6729,N_5122,N_4051);
and U6730 (N_6730,N_5847,N_4982);
nand U6731 (N_6731,N_5555,N_5833);
and U6732 (N_6732,N_4348,N_5222);
xor U6733 (N_6733,N_5441,N_4201);
and U6734 (N_6734,N_4411,N_4486);
and U6735 (N_6735,N_5405,N_4970);
nor U6736 (N_6736,N_5398,N_4934);
and U6737 (N_6737,N_4013,N_4582);
nand U6738 (N_6738,N_4699,N_4309);
nor U6739 (N_6739,N_4577,N_4775);
xor U6740 (N_6740,N_5226,N_4357);
or U6741 (N_6741,N_5588,N_4342);
or U6742 (N_6742,N_5747,N_5583);
and U6743 (N_6743,N_5751,N_4867);
or U6744 (N_6744,N_4812,N_5500);
xnor U6745 (N_6745,N_4887,N_5135);
and U6746 (N_6746,N_4142,N_4235);
and U6747 (N_6747,N_5996,N_5653);
xnor U6748 (N_6748,N_4030,N_4148);
nor U6749 (N_6749,N_5408,N_5067);
nor U6750 (N_6750,N_4082,N_4604);
nor U6751 (N_6751,N_4650,N_4877);
and U6752 (N_6752,N_4554,N_5945);
nor U6753 (N_6753,N_5823,N_4526);
or U6754 (N_6754,N_5079,N_5628);
and U6755 (N_6755,N_5054,N_5001);
or U6756 (N_6756,N_4920,N_5910);
and U6757 (N_6757,N_4156,N_5259);
nand U6758 (N_6758,N_4165,N_5545);
nand U6759 (N_6759,N_5948,N_5087);
xor U6760 (N_6760,N_4119,N_5692);
and U6761 (N_6761,N_4601,N_5651);
nor U6762 (N_6762,N_4192,N_4036);
nor U6763 (N_6763,N_5069,N_4362);
or U6764 (N_6764,N_5890,N_4050);
nor U6765 (N_6765,N_4258,N_5351);
and U6766 (N_6766,N_5012,N_5704);
nand U6767 (N_6767,N_5004,N_5726);
or U6768 (N_6768,N_4015,N_4363);
or U6769 (N_6769,N_5600,N_5117);
nor U6770 (N_6770,N_5992,N_4795);
or U6771 (N_6771,N_5043,N_4322);
nor U6772 (N_6772,N_4184,N_5710);
xor U6773 (N_6773,N_5918,N_4435);
xor U6774 (N_6774,N_4996,N_4152);
nor U6775 (N_6775,N_4428,N_5480);
and U6776 (N_6776,N_4664,N_5891);
xor U6777 (N_6777,N_5962,N_4678);
nand U6778 (N_6778,N_4759,N_4277);
or U6779 (N_6779,N_5170,N_4944);
nand U6780 (N_6780,N_4648,N_5049);
xor U6781 (N_6781,N_4990,N_5303);
or U6782 (N_6782,N_4660,N_5207);
nor U6783 (N_6783,N_4567,N_5656);
nor U6784 (N_6784,N_5633,N_4995);
or U6785 (N_6785,N_5498,N_5782);
xnor U6786 (N_6786,N_4392,N_5517);
nand U6787 (N_6787,N_4693,N_4282);
and U6788 (N_6788,N_4268,N_4077);
and U6789 (N_6789,N_5106,N_5379);
or U6790 (N_6790,N_4469,N_5347);
xnor U6791 (N_6791,N_5160,N_4572);
nand U6792 (N_6792,N_4159,N_4846);
and U6793 (N_6793,N_4640,N_5063);
xnor U6794 (N_6794,N_4094,N_5761);
and U6795 (N_6795,N_4368,N_5189);
and U6796 (N_6796,N_5864,N_4886);
xor U6797 (N_6797,N_4116,N_4000);
nand U6798 (N_6798,N_4396,N_5142);
nor U6799 (N_6799,N_4365,N_4005);
nand U6800 (N_6800,N_4238,N_4564);
nand U6801 (N_6801,N_5574,N_5107);
and U6802 (N_6802,N_5999,N_5572);
xnor U6803 (N_6803,N_4243,N_5922);
and U6804 (N_6804,N_5051,N_5466);
nor U6805 (N_6805,N_4568,N_4704);
and U6806 (N_6806,N_4127,N_5919);
nand U6807 (N_6807,N_5895,N_5820);
nor U6808 (N_6808,N_5763,N_5154);
nor U6809 (N_6809,N_4862,N_5931);
nand U6810 (N_6810,N_5083,N_5464);
xor U6811 (N_6811,N_5976,N_5385);
nor U6812 (N_6812,N_4651,N_4724);
and U6813 (N_6813,N_5179,N_4124);
and U6814 (N_6814,N_5654,N_4383);
xnor U6815 (N_6815,N_4559,N_4264);
or U6816 (N_6816,N_4946,N_5007);
and U6817 (N_6817,N_5728,N_4672);
and U6818 (N_6818,N_4641,N_5575);
xnor U6819 (N_6819,N_4993,N_5522);
or U6820 (N_6820,N_4285,N_5442);
nor U6821 (N_6821,N_4616,N_5705);
xor U6822 (N_6822,N_4402,N_4041);
or U6823 (N_6823,N_4190,N_4842);
and U6824 (N_6824,N_4203,N_5325);
or U6825 (N_6825,N_4840,N_4662);
and U6826 (N_6826,N_4248,N_5675);
nand U6827 (N_6827,N_4871,N_4835);
xor U6828 (N_6828,N_4923,N_4811);
nand U6829 (N_6829,N_5116,N_4848);
or U6830 (N_6830,N_4414,N_4876);
nor U6831 (N_6831,N_4295,N_4109);
and U6832 (N_6832,N_4666,N_4594);
and U6833 (N_6833,N_4781,N_5056);
nand U6834 (N_6834,N_4254,N_4878);
xor U6835 (N_6835,N_5971,N_4861);
or U6836 (N_6836,N_4581,N_5413);
nand U6837 (N_6837,N_4746,N_5099);
nor U6838 (N_6838,N_4794,N_5078);
xor U6839 (N_6839,N_4341,N_5781);
xor U6840 (N_6840,N_5038,N_5391);
nand U6841 (N_6841,N_5404,N_5243);
or U6842 (N_6842,N_5290,N_5514);
nand U6843 (N_6843,N_5240,N_4212);
and U6844 (N_6844,N_5267,N_5650);
nor U6845 (N_6845,N_4983,N_5942);
or U6846 (N_6846,N_4503,N_5900);
nor U6847 (N_6847,N_4501,N_5363);
and U6848 (N_6848,N_4715,N_4338);
xnor U6849 (N_6849,N_5493,N_4464);
nand U6850 (N_6850,N_4387,N_4347);
xor U6851 (N_6851,N_5940,N_5216);
or U6852 (N_6852,N_4896,N_5515);
nand U6853 (N_6853,N_4927,N_4869);
nand U6854 (N_6854,N_4791,N_4132);
nor U6855 (N_6855,N_4171,N_4787);
nand U6856 (N_6856,N_5417,N_4346);
nand U6857 (N_6857,N_5696,N_4118);
nand U6858 (N_6858,N_5582,N_5774);
xnor U6859 (N_6859,N_4320,N_4472);
nor U6860 (N_6860,N_4231,N_5912);
or U6861 (N_6861,N_4284,N_4304);
xnor U6862 (N_6862,N_4538,N_5227);
xnor U6863 (N_6863,N_4291,N_5247);
or U6864 (N_6864,N_4023,N_5258);
or U6865 (N_6865,N_5443,N_4978);
and U6866 (N_6866,N_4183,N_5807);
nand U6867 (N_6867,N_5569,N_5102);
nor U6868 (N_6868,N_4830,N_4686);
nor U6869 (N_6869,N_5491,N_4060);
or U6870 (N_6870,N_5685,N_4937);
nor U6871 (N_6871,N_5204,N_5796);
nor U6872 (N_6872,N_5110,N_4665);
nor U6873 (N_6873,N_4227,N_4596);
xnor U6874 (N_6874,N_5055,N_5547);
xnor U6875 (N_6875,N_4022,N_5241);
nand U6876 (N_6876,N_4892,N_5939);
or U6877 (N_6877,N_5101,N_5431);
nand U6878 (N_6878,N_5180,N_4214);
or U6879 (N_6879,N_4520,N_4476);
nand U6880 (N_6880,N_4545,N_4073);
or U6881 (N_6881,N_4513,N_4510);
nand U6882 (N_6882,N_5812,N_5469);
and U6883 (N_6883,N_4432,N_5741);
xnor U6884 (N_6884,N_4170,N_4587);
or U6885 (N_6885,N_5691,N_4606);
and U6886 (N_6886,N_4211,N_4038);
and U6887 (N_6887,N_4283,N_5148);
or U6888 (N_6888,N_5503,N_5977);
or U6889 (N_6889,N_5595,N_4479);
nand U6890 (N_6890,N_4090,N_5020);
and U6891 (N_6891,N_4328,N_5372);
or U6892 (N_6892,N_4832,N_4603);
and U6893 (N_6893,N_4224,N_5380);
xnor U6894 (N_6894,N_4857,N_5648);
and U6895 (N_6895,N_4553,N_5167);
xnor U6896 (N_6896,N_5615,N_5260);
or U6897 (N_6897,N_4316,N_5422);
and U6898 (N_6898,N_4307,N_4033);
and U6899 (N_6899,N_5612,N_5730);
or U6900 (N_6900,N_4916,N_4908);
and U6901 (N_6901,N_4239,N_5341);
and U6902 (N_6902,N_4173,N_5289);
nor U6903 (N_6903,N_4354,N_4244);
xor U6904 (N_6904,N_4305,N_5000);
or U6905 (N_6905,N_4198,N_5381);
or U6906 (N_6906,N_5776,N_5997);
nor U6907 (N_6907,N_4638,N_5342);
or U6908 (N_6908,N_5092,N_4081);
and U6909 (N_6909,N_4369,N_4125);
and U6910 (N_6910,N_4785,N_4964);
and U6911 (N_6911,N_4575,N_5037);
xor U6912 (N_6912,N_4599,N_4739);
and U6913 (N_6913,N_5098,N_5872);
xnor U6914 (N_6914,N_5130,N_5537);
nor U6915 (N_6915,N_4881,N_5542);
or U6916 (N_6916,N_5735,N_5418);
nand U6917 (N_6917,N_5266,N_4071);
or U6918 (N_6918,N_5319,N_5937);
and U6919 (N_6919,N_4512,N_5604);
nor U6920 (N_6920,N_5062,N_4622);
xnor U6921 (N_6921,N_5955,N_4353);
xnor U6922 (N_6922,N_5220,N_4972);
nand U6923 (N_6923,N_5666,N_4945);
nand U6924 (N_6924,N_4659,N_4106);
xor U6925 (N_6925,N_4940,N_4424);
nand U6926 (N_6926,N_4155,N_5930);
and U6927 (N_6927,N_5896,N_5894);
nand U6928 (N_6928,N_5905,N_4521);
or U6929 (N_6929,N_4780,N_4499);
nand U6930 (N_6930,N_5048,N_5868);
nand U6931 (N_6931,N_4228,N_5982);
nand U6932 (N_6932,N_4950,N_4631);
nor U6933 (N_6933,N_4685,N_4849);
nand U6934 (N_6934,N_4474,N_5990);
nand U6935 (N_6935,N_4919,N_4162);
nand U6936 (N_6936,N_5840,N_4850);
nand U6937 (N_6937,N_4314,N_5966);
or U6938 (N_6938,N_5903,N_4117);
nand U6939 (N_6939,N_5061,N_4053);
and U6940 (N_6940,N_5546,N_4729);
xnor U6941 (N_6941,N_4242,N_5677);
or U6942 (N_6942,N_5129,N_5965);
or U6943 (N_6943,N_5237,N_4834);
nor U6944 (N_6944,N_5238,N_4874);
nor U6945 (N_6945,N_5425,N_5511);
nor U6946 (N_6946,N_5642,N_5019);
or U6947 (N_6947,N_5109,N_5210);
or U6948 (N_6948,N_4766,N_4808);
and U6949 (N_6949,N_5802,N_4904);
and U6950 (N_6950,N_4456,N_5808);
xnor U6951 (N_6951,N_4367,N_4825);
nor U6952 (N_6952,N_4482,N_5797);
nor U6953 (N_6953,N_4025,N_4921);
and U6954 (N_6954,N_5483,N_4431);
nor U6955 (N_6955,N_4146,N_4656);
nor U6956 (N_6956,N_4618,N_5719);
or U6957 (N_6957,N_4992,N_4312);
and U6958 (N_6958,N_4853,N_5462);
and U6959 (N_6959,N_4325,N_5954);
nand U6960 (N_6960,N_5409,N_5662);
or U6961 (N_6961,N_5926,N_5765);
nor U6962 (N_6962,N_4072,N_4301);
and U6963 (N_6963,N_4928,N_5672);
or U6964 (N_6964,N_4350,N_4179);
nand U6965 (N_6965,N_4895,N_5590);
and U6966 (N_6966,N_5620,N_5358);
and U6967 (N_6967,N_4776,N_5707);
and U6968 (N_6968,N_4778,N_5529);
xor U6969 (N_6969,N_5014,N_5841);
nand U6970 (N_6970,N_5330,N_5182);
and U6971 (N_6971,N_4177,N_4905);
xor U6972 (N_6972,N_4843,N_5495);
xor U6973 (N_6973,N_5748,N_5561);
nand U6974 (N_6974,N_4064,N_5050);
nand U6975 (N_6975,N_4209,N_5597);
nor U6976 (N_6976,N_4182,N_5151);
nand U6977 (N_6977,N_4220,N_5790);
xor U6978 (N_6978,N_4099,N_5753);
nand U6979 (N_6979,N_5667,N_4373);
xnor U6980 (N_6980,N_5711,N_5232);
nand U6981 (N_6981,N_5854,N_5611);
and U6982 (N_6982,N_4421,N_5415);
nand U6983 (N_6983,N_4093,N_4615);
xor U6984 (N_6984,N_5523,N_4491);
xor U6985 (N_6985,N_4508,N_4960);
and U6986 (N_6986,N_4371,N_5734);
nor U6987 (N_6987,N_5837,N_5567);
nor U6988 (N_6988,N_4425,N_5440);
or U6989 (N_6989,N_5679,N_5643);
or U6990 (N_6990,N_4930,N_4856);
xor U6991 (N_6991,N_4166,N_4452);
xor U6992 (N_6992,N_4912,N_5979);
nand U6993 (N_6993,N_4536,N_5509);
nand U6994 (N_6994,N_4801,N_4719);
nand U6995 (N_6995,N_5343,N_4087);
xnor U6996 (N_6996,N_5746,N_5324);
or U6997 (N_6997,N_5622,N_4516);
nand U6998 (N_6998,N_4185,N_4016);
or U6999 (N_6999,N_4494,N_4275);
and U7000 (N_7000,N_5636,N_5432);
or U7001 (N_7001,N_4227,N_4500);
nand U7002 (N_7002,N_4480,N_5832);
or U7003 (N_7003,N_5230,N_4957);
or U7004 (N_7004,N_4469,N_5123);
nand U7005 (N_7005,N_5581,N_5875);
or U7006 (N_7006,N_5181,N_5202);
or U7007 (N_7007,N_5730,N_4105);
xnor U7008 (N_7008,N_4419,N_4853);
or U7009 (N_7009,N_5669,N_4200);
nand U7010 (N_7010,N_5411,N_5719);
nor U7011 (N_7011,N_4588,N_5569);
and U7012 (N_7012,N_4012,N_4039);
nor U7013 (N_7013,N_4059,N_5641);
or U7014 (N_7014,N_4276,N_4917);
and U7015 (N_7015,N_4039,N_5428);
xnor U7016 (N_7016,N_5500,N_4132);
or U7017 (N_7017,N_4386,N_4269);
and U7018 (N_7018,N_5664,N_4909);
and U7019 (N_7019,N_5756,N_5130);
nand U7020 (N_7020,N_5759,N_4180);
xor U7021 (N_7021,N_4070,N_4871);
xor U7022 (N_7022,N_4139,N_4903);
or U7023 (N_7023,N_4117,N_5446);
nor U7024 (N_7024,N_5843,N_4288);
or U7025 (N_7025,N_5270,N_5211);
nor U7026 (N_7026,N_4393,N_4450);
nand U7027 (N_7027,N_4988,N_5609);
and U7028 (N_7028,N_5505,N_5742);
nand U7029 (N_7029,N_4208,N_4496);
nand U7030 (N_7030,N_4799,N_5445);
nand U7031 (N_7031,N_4612,N_4226);
nand U7032 (N_7032,N_4815,N_5766);
nand U7033 (N_7033,N_4145,N_5372);
xnor U7034 (N_7034,N_5565,N_5692);
nand U7035 (N_7035,N_4611,N_4637);
nor U7036 (N_7036,N_5165,N_5585);
xnor U7037 (N_7037,N_5968,N_4682);
nand U7038 (N_7038,N_4216,N_4112);
xor U7039 (N_7039,N_4839,N_4429);
or U7040 (N_7040,N_5613,N_4687);
or U7041 (N_7041,N_4446,N_4349);
nor U7042 (N_7042,N_5298,N_5972);
nor U7043 (N_7043,N_4209,N_5664);
and U7044 (N_7044,N_4754,N_5546);
or U7045 (N_7045,N_4468,N_5848);
xnor U7046 (N_7046,N_5477,N_4134);
or U7047 (N_7047,N_5155,N_5088);
or U7048 (N_7048,N_4052,N_5848);
and U7049 (N_7049,N_5685,N_4779);
xor U7050 (N_7050,N_5031,N_5702);
nor U7051 (N_7051,N_5677,N_4521);
nor U7052 (N_7052,N_4067,N_5163);
nand U7053 (N_7053,N_5123,N_4882);
xor U7054 (N_7054,N_5215,N_4974);
xnor U7055 (N_7055,N_5716,N_5088);
nor U7056 (N_7056,N_4793,N_4947);
and U7057 (N_7057,N_4791,N_4802);
and U7058 (N_7058,N_4825,N_5220);
nand U7059 (N_7059,N_4432,N_5918);
or U7060 (N_7060,N_4318,N_5172);
or U7061 (N_7061,N_4456,N_4243);
xor U7062 (N_7062,N_4142,N_4237);
and U7063 (N_7063,N_4509,N_4946);
nand U7064 (N_7064,N_5963,N_4571);
or U7065 (N_7065,N_4033,N_4481);
or U7066 (N_7066,N_5189,N_4788);
and U7067 (N_7067,N_4242,N_4009);
nor U7068 (N_7068,N_4320,N_4377);
or U7069 (N_7069,N_5106,N_5204);
nand U7070 (N_7070,N_5528,N_5411);
or U7071 (N_7071,N_5456,N_5854);
and U7072 (N_7072,N_4037,N_5335);
nand U7073 (N_7073,N_5320,N_4379);
or U7074 (N_7074,N_5503,N_5428);
or U7075 (N_7075,N_5805,N_5284);
and U7076 (N_7076,N_5545,N_4079);
nand U7077 (N_7077,N_4856,N_4073);
nand U7078 (N_7078,N_5798,N_4544);
and U7079 (N_7079,N_4845,N_4820);
and U7080 (N_7080,N_4835,N_5305);
nand U7081 (N_7081,N_5898,N_4928);
or U7082 (N_7082,N_4857,N_5396);
or U7083 (N_7083,N_5595,N_5413);
and U7084 (N_7084,N_5627,N_4420);
xnor U7085 (N_7085,N_4415,N_4842);
xor U7086 (N_7086,N_4255,N_5090);
or U7087 (N_7087,N_4138,N_4245);
xor U7088 (N_7088,N_5043,N_4986);
and U7089 (N_7089,N_4887,N_4723);
or U7090 (N_7090,N_5694,N_4700);
and U7091 (N_7091,N_5539,N_5186);
nor U7092 (N_7092,N_4053,N_5267);
nand U7093 (N_7093,N_5799,N_5222);
nor U7094 (N_7094,N_4470,N_4979);
nor U7095 (N_7095,N_5378,N_5720);
nor U7096 (N_7096,N_4202,N_5207);
nand U7097 (N_7097,N_5966,N_5960);
nand U7098 (N_7098,N_4253,N_5269);
or U7099 (N_7099,N_4165,N_4667);
or U7100 (N_7100,N_4618,N_4474);
xnor U7101 (N_7101,N_4928,N_5412);
nor U7102 (N_7102,N_5016,N_4603);
or U7103 (N_7103,N_4657,N_5526);
xor U7104 (N_7104,N_5132,N_5883);
xor U7105 (N_7105,N_5945,N_4399);
and U7106 (N_7106,N_4088,N_5594);
and U7107 (N_7107,N_4873,N_5201);
nand U7108 (N_7108,N_4728,N_5888);
xor U7109 (N_7109,N_5014,N_4445);
and U7110 (N_7110,N_4197,N_5331);
nand U7111 (N_7111,N_4515,N_4236);
or U7112 (N_7112,N_5020,N_4520);
nand U7113 (N_7113,N_4659,N_4545);
nand U7114 (N_7114,N_4440,N_4698);
and U7115 (N_7115,N_4184,N_4595);
nand U7116 (N_7116,N_5066,N_4075);
and U7117 (N_7117,N_4785,N_5292);
nand U7118 (N_7118,N_5379,N_5452);
nor U7119 (N_7119,N_5995,N_5384);
nor U7120 (N_7120,N_5835,N_5285);
and U7121 (N_7121,N_4707,N_5380);
and U7122 (N_7122,N_5235,N_5975);
and U7123 (N_7123,N_4641,N_4136);
nand U7124 (N_7124,N_5995,N_5610);
nand U7125 (N_7125,N_4239,N_5864);
nand U7126 (N_7126,N_5323,N_4013);
and U7127 (N_7127,N_5923,N_4611);
nand U7128 (N_7128,N_4659,N_5693);
xor U7129 (N_7129,N_5595,N_4381);
nor U7130 (N_7130,N_4672,N_5043);
and U7131 (N_7131,N_5876,N_4687);
or U7132 (N_7132,N_5652,N_4078);
or U7133 (N_7133,N_5776,N_4421);
nor U7134 (N_7134,N_4635,N_4028);
nor U7135 (N_7135,N_4828,N_4084);
or U7136 (N_7136,N_5919,N_5670);
xnor U7137 (N_7137,N_5192,N_5868);
nand U7138 (N_7138,N_5235,N_5399);
and U7139 (N_7139,N_5397,N_4341);
or U7140 (N_7140,N_5569,N_5807);
nor U7141 (N_7141,N_4440,N_5515);
nand U7142 (N_7142,N_4474,N_4290);
and U7143 (N_7143,N_4300,N_5645);
and U7144 (N_7144,N_5994,N_4390);
nand U7145 (N_7145,N_4392,N_4921);
xor U7146 (N_7146,N_5497,N_4323);
nand U7147 (N_7147,N_5548,N_5193);
xor U7148 (N_7148,N_4515,N_5193);
or U7149 (N_7149,N_4230,N_5912);
and U7150 (N_7150,N_5317,N_5177);
or U7151 (N_7151,N_5261,N_5824);
and U7152 (N_7152,N_5548,N_5380);
xnor U7153 (N_7153,N_5822,N_5173);
or U7154 (N_7154,N_4970,N_4764);
or U7155 (N_7155,N_4054,N_5220);
nor U7156 (N_7156,N_5295,N_4684);
nor U7157 (N_7157,N_5266,N_4229);
xor U7158 (N_7158,N_4912,N_4621);
nor U7159 (N_7159,N_4259,N_4087);
and U7160 (N_7160,N_5905,N_5680);
xor U7161 (N_7161,N_4650,N_5349);
nor U7162 (N_7162,N_5062,N_5850);
and U7163 (N_7163,N_5171,N_5172);
nand U7164 (N_7164,N_5019,N_5571);
xnor U7165 (N_7165,N_5288,N_4027);
and U7166 (N_7166,N_5962,N_4367);
and U7167 (N_7167,N_5328,N_5106);
nor U7168 (N_7168,N_5285,N_5813);
or U7169 (N_7169,N_4523,N_5541);
nor U7170 (N_7170,N_4442,N_4817);
nor U7171 (N_7171,N_5684,N_4882);
xnor U7172 (N_7172,N_5175,N_5387);
xor U7173 (N_7173,N_5364,N_5068);
or U7174 (N_7174,N_5560,N_4464);
and U7175 (N_7175,N_4376,N_4304);
xor U7176 (N_7176,N_5756,N_5322);
xnor U7177 (N_7177,N_4103,N_5498);
nand U7178 (N_7178,N_5092,N_4939);
and U7179 (N_7179,N_5697,N_5577);
nand U7180 (N_7180,N_4877,N_5945);
nand U7181 (N_7181,N_4710,N_5502);
nand U7182 (N_7182,N_4067,N_4042);
nor U7183 (N_7183,N_5342,N_4251);
xnor U7184 (N_7184,N_5716,N_5386);
and U7185 (N_7185,N_5149,N_4217);
or U7186 (N_7186,N_4240,N_5860);
nand U7187 (N_7187,N_5032,N_5789);
or U7188 (N_7188,N_5519,N_4139);
or U7189 (N_7189,N_4057,N_4082);
and U7190 (N_7190,N_4557,N_5597);
and U7191 (N_7191,N_4317,N_5990);
xnor U7192 (N_7192,N_4279,N_4340);
nand U7193 (N_7193,N_5129,N_5357);
and U7194 (N_7194,N_5219,N_5010);
nor U7195 (N_7195,N_4422,N_5073);
nand U7196 (N_7196,N_4301,N_4538);
xnor U7197 (N_7197,N_5252,N_4753);
or U7198 (N_7198,N_4978,N_4319);
or U7199 (N_7199,N_5636,N_4150);
xnor U7200 (N_7200,N_5595,N_4263);
and U7201 (N_7201,N_5107,N_5327);
or U7202 (N_7202,N_4335,N_4214);
or U7203 (N_7203,N_5318,N_5024);
and U7204 (N_7204,N_4151,N_4708);
nor U7205 (N_7205,N_4566,N_4615);
and U7206 (N_7206,N_4148,N_5578);
xnor U7207 (N_7207,N_4545,N_4611);
and U7208 (N_7208,N_5133,N_4423);
nor U7209 (N_7209,N_4726,N_4444);
and U7210 (N_7210,N_4049,N_4177);
nor U7211 (N_7211,N_4905,N_4748);
xor U7212 (N_7212,N_4494,N_4711);
or U7213 (N_7213,N_5004,N_5927);
xor U7214 (N_7214,N_4274,N_5817);
xor U7215 (N_7215,N_4722,N_4878);
or U7216 (N_7216,N_5266,N_4114);
nor U7217 (N_7217,N_5572,N_5940);
and U7218 (N_7218,N_5337,N_4939);
nor U7219 (N_7219,N_5852,N_4362);
or U7220 (N_7220,N_5593,N_4455);
nor U7221 (N_7221,N_4627,N_5491);
or U7222 (N_7222,N_5231,N_5026);
nor U7223 (N_7223,N_4485,N_4193);
nand U7224 (N_7224,N_4921,N_4991);
nand U7225 (N_7225,N_4211,N_5023);
or U7226 (N_7226,N_5074,N_4085);
xnor U7227 (N_7227,N_4724,N_4110);
nand U7228 (N_7228,N_4472,N_5284);
xor U7229 (N_7229,N_5915,N_5529);
nand U7230 (N_7230,N_4971,N_5238);
nor U7231 (N_7231,N_5800,N_5617);
nand U7232 (N_7232,N_4869,N_5139);
nand U7233 (N_7233,N_4504,N_5732);
nor U7234 (N_7234,N_5189,N_4080);
xnor U7235 (N_7235,N_4466,N_5544);
or U7236 (N_7236,N_4202,N_4648);
nand U7237 (N_7237,N_4590,N_5217);
nand U7238 (N_7238,N_5200,N_5831);
and U7239 (N_7239,N_5652,N_4990);
nor U7240 (N_7240,N_4088,N_4090);
and U7241 (N_7241,N_5958,N_5039);
nor U7242 (N_7242,N_5900,N_5141);
or U7243 (N_7243,N_5619,N_4147);
xor U7244 (N_7244,N_5210,N_5613);
nand U7245 (N_7245,N_5958,N_5541);
and U7246 (N_7246,N_5486,N_5192);
and U7247 (N_7247,N_4806,N_5137);
or U7248 (N_7248,N_5454,N_5997);
nor U7249 (N_7249,N_5197,N_5209);
xor U7250 (N_7250,N_5358,N_4692);
and U7251 (N_7251,N_4115,N_5299);
and U7252 (N_7252,N_4646,N_4630);
xor U7253 (N_7253,N_5046,N_5420);
nand U7254 (N_7254,N_4085,N_4015);
and U7255 (N_7255,N_5210,N_5228);
nor U7256 (N_7256,N_5852,N_5207);
or U7257 (N_7257,N_5033,N_4560);
and U7258 (N_7258,N_4264,N_5017);
or U7259 (N_7259,N_4160,N_4008);
or U7260 (N_7260,N_5413,N_5409);
xor U7261 (N_7261,N_5203,N_5125);
and U7262 (N_7262,N_4581,N_4035);
nor U7263 (N_7263,N_5050,N_5875);
xor U7264 (N_7264,N_4060,N_5211);
nor U7265 (N_7265,N_5400,N_4361);
or U7266 (N_7266,N_5491,N_4182);
or U7267 (N_7267,N_5432,N_5882);
and U7268 (N_7268,N_5402,N_4708);
nor U7269 (N_7269,N_5667,N_4378);
nand U7270 (N_7270,N_4398,N_5353);
and U7271 (N_7271,N_4114,N_4547);
nand U7272 (N_7272,N_5380,N_5104);
nand U7273 (N_7273,N_5386,N_5481);
or U7274 (N_7274,N_4027,N_4044);
nand U7275 (N_7275,N_4783,N_5027);
nor U7276 (N_7276,N_5940,N_5029);
nand U7277 (N_7277,N_4610,N_5723);
nor U7278 (N_7278,N_5431,N_5509);
xor U7279 (N_7279,N_5816,N_5468);
and U7280 (N_7280,N_5565,N_5635);
nand U7281 (N_7281,N_4070,N_4718);
or U7282 (N_7282,N_5153,N_5994);
or U7283 (N_7283,N_4062,N_5178);
and U7284 (N_7284,N_4584,N_4810);
nand U7285 (N_7285,N_4610,N_5460);
or U7286 (N_7286,N_5569,N_5215);
xnor U7287 (N_7287,N_5033,N_5520);
or U7288 (N_7288,N_4732,N_5166);
and U7289 (N_7289,N_5842,N_4480);
nand U7290 (N_7290,N_4949,N_5409);
xnor U7291 (N_7291,N_4059,N_5458);
or U7292 (N_7292,N_4420,N_4793);
nand U7293 (N_7293,N_5613,N_4819);
xor U7294 (N_7294,N_5771,N_4932);
xnor U7295 (N_7295,N_4005,N_5667);
and U7296 (N_7296,N_5326,N_4084);
or U7297 (N_7297,N_5216,N_4747);
nor U7298 (N_7298,N_4200,N_5229);
xnor U7299 (N_7299,N_5795,N_5558);
nor U7300 (N_7300,N_4653,N_5627);
or U7301 (N_7301,N_5061,N_5695);
nor U7302 (N_7302,N_5710,N_5052);
and U7303 (N_7303,N_4049,N_5320);
or U7304 (N_7304,N_4363,N_4813);
and U7305 (N_7305,N_4311,N_5495);
and U7306 (N_7306,N_4107,N_5746);
and U7307 (N_7307,N_4409,N_4581);
xnor U7308 (N_7308,N_4272,N_4776);
nor U7309 (N_7309,N_4220,N_5412);
nand U7310 (N_7310,N_5635,N_4120);
nand U7311 (N_7311,N_4519,N_5060);
nor U7312 (N_7312,N_5085,N_4777);
xnor U7313 (N_7313,N_4566,N_5134);
or U7314 (N_7314,N_5056,N_5003);
or U7315 (N_7315,N_5857,N_5642);
and U7316 (N_7316,N_5428,N_4143);
and U7317 (N_7317,N_5454,N_4969);
and U7318 (N_7318,N_5413,N_5322);
xnor U7319 (N_7319,N_5443,N_5807);
nand U7320 (N_7320,N_5172,N_5984);
or U7321 (N_7321,N_4526,N_5836);
nor U7322 (N_7322,N_5439,N_4619);
nor U7323 (N_7323,N_5380,N_4714);
xor U7324 (N_7324,N_4722,N_5537);
xor U7325 (N_7325,N_4737,N_4431);
nand U7326 (N_7326,N_5782,N_5739);
or U7327 (N_7327,N_4998,N_4294);
nor U7328 (N_7328,N_5880,N_4747);
or U7329 (N_7329,N_4602,N_4442);
nor U7330 (N_7330,N_4071,N_4790);
xor U7331 (N_7331,N_4496,N_4292);
and U7332 (N_7332,N_5340,N_4148);
or U7333 (N_7333,N_4816,N_5713);
and U7334 (N_7334,N_5554,N_5567);
nor U7335 (N_7335,N_5803,N_4652);
nor U7336 (N_7336,N_4014,N_4313);
and U7337 (N_7337,N_4415,N_5786);
and U7338 (N_7338,N_4851,N_4676);
nor U7339 (N_7339,N_5099,N_5460);
xnor U7340 (N_7340,N_5845,N_4612);
nand U7341 (N_7341,N_4789,N_5657);
nor U7342 (N_7342,N_4296,N_4417);
xor U7343 (N_7343,N_4487,N_5357);
nor U7344 (N_7344,N_4696,N_4398);
nand U7345 (N_7345,N_4329,N_5466);
and U7346 (N_7346,N_5074,N_4170);
and U7347 (N_7347,N_5346,N_4422);
xor U7348 (N_7348,N_4498,N_5790);
nor U7349 (N_7349,N_5459,N_5269);
xor U7350 (N_7350,N_4311,N_4499);
nand U7351 (N_7351,N_5492,N_4943);
or U7352 (N_7352,N_4176,N_5686);
nand U7353 (N_7353,N_4112,N_5263);
nor U7354 (N_7354,N_4036,N_4374);
nand U7355 (N_7355,N_5156,N_5451);
and U7356 (N_7356,N_4422,N_5439);
nor U7357 (N_7357,N_4556,N_5218);
or U7358 (N_7358,N_4146,N_4269);
nor U7359 (N_7359,N_4429,N_5981);
nor U7360 (N_7360,N_5244,N_5932);
nand U7361 (N_7361,N_5490,N_5665);
nand U7362 (N_7362,N_4228,N_4667);
and U7363 (N_7363,N_5913,N_4936);
or U7364 (N_7364,N_4901,N_4647);
nand U7365 (N_7365,N_5737,N_4283);
and U7366 (N_7366,N_4301,N_5522);
and U7367 (N_7367,N_5494,N_5787);
nor U7368 (N_7368,N_5018,N_4618);
and U7369 (N_7369,N_4989,N_4942);
nand U7370 (N_7370,N_4704,N_4622);
nand U7371 (N_7371,N_5374,N_5688);
or U7372 (N_7372,N_4164,N_4923);
nand U7373 (N_7373,N_4706,N_5426);
nand U7374 (N_7374,N_5969,N_5953);
and U7375 (N_7375,N_4852,N_5137);
or U7376 (N_7376,N_5862,N_5000);
xnor U7377 (N_7377,N_4030,N_4933);
xnor U7378 (N_7378,N_5354,N_4130);
or U7379 (N_7379,N_4247,N_5199);
or U7380 (N_7380,N_4144,N_4923);
or U7381 (N_7381,N_4134,N_5056);
nor U7382 (N_7382,N_5424,N_4832);
nor U7383 (N_7383,N_4003,N_4184);
or U7384 (N_7384,N_4298,N_4522);
xor U7385 (N_7385,N_4723,N_4280);
nand U7386 (N_7386,N_5837,N_4239);
nor U7387 (N_7387,N_4399,N_5105);
nor U7388 (N_7388,N_4663,N_5950);
nand U7389 (N_7389,N_4225,N_4128);
nor U7390 (N_7390,N_4555,N_5668);
nor U7391 (N_7391,N_4288,N_5744);
or U7392 (N_7392,N_4038,N_5324);
nand U7393 (N_7393,N_5337,N_4967);
and U7394 (N_7394,N_5438,N_5234);
nand U7395 (N_7395,N_5975,N_5344);
nand U7396 (N_7396,N_4027,N_5604);
or U7397 (N_7397,N_4633,N_4355);
or U7398 (N_7398,N_5972,N_5920);
xor U7399 (N_7399,N_5684,N_5809);
xnor U7400 (N_7400,N_5529,N_4797);
nand U7401 (N_7401,N_4011,N_4225);
nor U7402 (N_7402,N_4621,N_5201);
and U7403 (N_7403,N_4130,N_5896);
nand U7404 (N_7404,N_5826,N_5750);
and U7405 (N_7405,N_5669,N_5262);
and U7406 (N_7406,N_4782,N_5234);
or U7407 (N_7407,N_5179,N_4033);
nand U7408 (N_7408,N_4961,N_4222);
or U7409 (N_7409,N_5706,N_5499);
and U7410 (N_7410,N_5013,N_4497);
and U7411 (N_7411,N_5486,N_4467);
xnor U7412 (N_7412,N_4262,N_5360);
xor U7413 (N_7413,N_4897,N_4966);
nand U7414 (N_7414,N_4533,N_4363);
and U7415 (N_7415,N_4554,N_4052);
xor U7416 (N_7416,N_5389,N_5725);
xnor U7417 (N_7417,N_5743,N_5037);
nand U7418 (N_7418,N_4965,N_5721);
or U7419 (N_7419,N_5974,N_4915);
xnor U7420 (N_7420,N_5963,N_4294);
and U7421 (N_7421,N_4297,N_5566);
and U7422 (N_7422,N_4184,N_4611);
nand U7423 (N_7423,N_5516,N_4221);
nor U7424 (N_7424,N_4888,N_4970);
and U7425 (N_7425,N_5906,N_4648);
nand U7426 (N_7426,N_5128,N_4707);
nand U7427 (N_7427,N_4872,N_4934);
nand U7428 (N_7428,N_4600,N_5702);
nor U7429 (N_7429,N_5291,N_5161);
nor U7430 (N_7430,N_5721,N_4438);
nand U7431 (N_7431,N_4896,N_4077);
and U7432 (N_7432,N_5378,N_4100);
or U7433 (N_7433,N_4838,N_5963);
nor U7434 (N_7434,N_4635,N_4845);
xor U7435 (N_7435,N_5094,N_5363);
and U7436 (N_7436,N_5625,N_4665);
or U7437 (N_7437,N_4302,N_5608);
and U7438 (N_7438,N_4953,N_4153);
nor U7439 (N_7439,N_5699,N_5966);
nand U7440 (N_7440,N_5351,N_4643);
xor U7441 (N_7441,N_4416,N_4252);
and U7442 (N_7442,N_5025,N_4200);
nand U7443 (N_7443,N_5101,N_4246);
nand U7444 (N_7444,N_5074,N_5040);
or U7445 (N_7445,N_5457,N_5320);
nand U7446 (N_7446,N_4639,N_4911);
and U7447 (N_7447,N_5778,N_5674);
or U7448 (N_7448,N_5735,N_4786);
nor U7449 (N_7449,N_4518,N_5474);
nand U7450 (N_7450,N_5149,N_5303);
or U7451 (N_7451,N_5659,N_4256);
nand U7452 (N_7452,N_4546,N_4432);
xnor U7453 (N_7453,N_5785,N_5035);
nand U7454 (N_7454,N_5390,N_5702);
or U7455 (N_7455,N_4517,N_5536);
nor U7456 (N_7456,N_5011,N_4022);
and U7457 (N_7457,N_5715,N_4401);
or U7458 (N_7458,N_4509,N_5409);
or U7459 (N_7459,N_5708,N_5444);
nor U7460 (N_7460,N_5666,N_5607);
or U7461 (N_7461,N_5142,N_5042);
xnor U7462 (N_7462,N_4303,N_5907);
and U7463 (N_7463,N_4517,N_4590);
xor U7464 (N_7464,N_4271,N_4815);
or U7465 (N_7465,N_5843,N_4028);
xor U7466 (N_7466,N_5188,N_5575);
nor U7467 (N_7467,N_4057,N_5280);
nand U7468 (N_7468,N_4943,N_4811);
or U7469 (N_7469,N_4417,N_5912);
nor U7470 (N_7470,N_5651,N_5902);
xnor U7471 (N_7471,N_4634,N_4838);
xnor U7472 (N_7472,N_5795,N_4909);
nand U7473 (N_7473,N_5104,N_5491);
nor U7474 (N_7474,N_4502,N_5878);
xor U7475 (N_7475,N_5855,N_5574);
or U7476 (N_7476,N_5027,N_4429);
nor U7477 (N_7477,N_4473,N_5296);
and U7478 (N_7478,N_4581,N_5464);
nand U7479 (N_7479,N_4025,N_5880);
nand U7480 (N_7480,N_4320,N_5306);
xor U7481 (N_7481,N_5625,N_5059);
or U7482 (N_7482,N_4219,N_4480);
or U7483 (N_7483,N_5285,N_4999);
nand U7484 (N_7484,N_4206,N_5003);
or U7485 (N_7485,N_5181,N_4049);
xor U7486 (N_7486,N_5118,N_4017);
and U7487 (N_7487,N_4532,N_5262);
and U7488 (N_7488,N_4326,N_5149);
nand U7489 (N_7489,N_5480,N_5942);
and U7490 (N_7490,N_5398,N_4040);
or U7491 (N_7491,N_5870,N_5239);
or U7492 (N_7492,N_5313,N_4344);
or U7493 (N_7493,N_4710,N_5614);
nand U7494 (N_7494,N_5404,N_4804);
nand U7495 (N_7495,N_5527,N_4021);
and U7496 (N_7496,N_5198,N_4887);
nor U7497 (N_7497,N_5937,N_5882);
and U7498 (N_7498,N_5368,N_4695);
xor U7499 (N_7499,N_4936,N_4089);
or U7500 (N_7500,N_5214,N_5697);
and U7501 (N_7501,N_4640,N_4071);
nand U7502 (N_7502,N_5340,N_5108);
or U7503 (N_7503,N_5026,N_4678);
and U7504 (N_7504,N_5913,N_5757);
xnor U7505 (N_7505,N_5109,N_5660);
nor U7506 (N_7506,N_4026,N_4274);
nand U7507 (N_7507,N_4517,N_4626);
nor U7508 (N_7508,N_4629,N_4721);
or U7509 (N_7509,N_4047,N_5969);
nand U7510 (N_7510,N_5953,N_4485);
xnor U7511 (N_7511,N_5640,N_4871);
or U7512 (N_7512,N_4874,N_5228);
or U7513 (N_7513,N_5164,N_5179);
or U7514 (N_7514,N_5333,N_5651);
and U7515 (N_7515,N_4879,N_5030);
or U7516 (N_7516,N_4524,N_5233);
and U7517 (N_7517,N_5044,N_5409);
or U7518 (N_7518,N_5841,N_4626);
nand U7519 (N_7519,N_5491,N_4948);
and U7520 (N_7520,N_5406,N_5972);
xnor U7521 (N_7521,N_5107,N_5603);
or U7522 (N_7522,N_5477,N_4889);
xnor U7523 (N_7523,N_4795,N_5850);
nand U7524 (N_7524,N_5434,N_5022);
nand U7525 (N_7525,N_5312,N_4402);
and U7526 (N_7526,N_4595,N_5548);
and U7527 (N_7527,N_4740,N_5013);
nor U7528 (N_7528,N_4036,N_5183);
nand U7529 (N_7529,N_4093,N_4401);
and U7530 (N_7530,N_5502,N_4962);
nor U7531 (N_7531,N_4355,N_4976);
and U7532 (N_7532,N_5394,N_5716);
nand U7533 (N_7533,N_4875,N_4368);
xor U7534 (N_7534,N_4864,N_4623);
nor U7535 (N_7535,N_5101,N_5646);
and U7536 (N_7536,N_4085,N_4428);
or U7537 (N_7537,N_4793,N_4499);
or U7538 (N_7538,N_5024,N_4691);
or U7539 (N_7539,N_5295,N_4443);
xor U7540 (N_7540,N_5009,N_5335);
nand U7541 (N_7541,N_5047,N_5556);
nand U7542 (N_7542,N_5398,N_5762);
nand U7543 (N_7543,N_5837,N_4743);
nand U7544 (N_7544,N_4333,N_5092);
nand U7545 (N_7545,N_4981,N_5663);
nor U7546 (N_7546,N_5044,N_4095);
and U7547 (N_7547,N_5930,N_4393);
nand U7548 (N_7548,N_5108,N_5168);
or U7549 (N_7549,N_4388,N_5521);
and U7550 (N_7550,N_5038,N_5431);
nand U7551 (N_7551,N_4769,N_5858);
or U7552 (N_7552,N_5783,N_5771);
and U7553 (N_7553,N_4616,N_4555);
and U7554 (N_7554,N_5467,N_4831);
and U7555 (N_7555,N_4116,N_5050);
and U7556 (N_7556,N_5661,N_4828);
nor U7557 (N_7557,N_5164,N_5287);
nand U7558 (N_7558,N_5950,N_5185);
nor U7559 (N_7559,N_4849,N_4750);
and U7560 (N_7560,N_4453,N_5447);
nand U7561 (N_7561,N_4732,N_5910);
nand U7562 (N_7562,N_5703,N_5002);
and U7563 (N_7563,N_5843,N_5248);
and U7564 (N_7564,N_4398,N_5780);
nand U7565 (N_7565,N_4047,N_5681);
or U7566 (N_7566,N_4394,N_5134);
xnor U7567 (N_7567,N_4845,N_5711);
nand U7568 (N_7568,N_5200,N_5404);
and U7569 (N_7569,N_5145,N_4911);
or U7570 (N_7570,N_5054,N_4132);
or U7571 (N_7571,N_5642,N_4153);
or U7572 (N_7572,N_5988,N_5269);
and U7573 (N_7573,N_4469,N_4572);
and U7574 (N_7574,N_5640,N_4052);
and U7575 (N_7575,N_4184,N_5920);
nand U7576 (N_7576,N_5504,N_4928);
or U7577 (N_7577,N_5208,N_4207);
and U7578 (N_7578,N_4062,N_4111);
nor U7579 (N_7579,N_5112,N_4635);
or U7580 (N_7580,N_4541,N_5000);
nand U7581 (N_7581,N_4991,N_4830);
xor U7582 (N_7582,N_4783,N_5929);
xnor U7583 (N_7583,N_5358,N_4760);
or U7584 (N_7584,N_4295,N_4363);
nand U7585 (N_7585,N_5285,N_5927);
or U7586 (N_7586,N_5287,N_5787);
nand U7587 (N_7587,N_5514,N_5225);
xor U7588 (N_7588,N_4994,N_5150);
nand U7589 (N_7589,N_5961,N_4464);
nor U7590 (N_7590,N_5931,N_5461);
and U7591 (N_7591,N_5277,N_4532);
nor U7592 (N_7592,N_4556,N_5980);
and U7593 (N_7593,N_5326,N_5044);
nand U7594 (N_7594,N_5072,N_5396);
or U7595 (N_7595,N_4832,N_4540);
or U7596 (N_7596,N_4438,N_4642);
xnor U7597 (N_7597,N_4187,N_4853);
or U7598 (N_7598,N_4247,N_5813);
nor U7599 (N_7599,N_5158,N_4957);
nor U7600 (N_7600,N_4173,N_5941);
nand U7601 (N_7601,N_5099,N_5253);
nor U7602 (N_7602,N_5875,N_4524);
nand U7603 (N_7603,N_4712,N_5402);
nand U7604 (N_7604,N_5103,N_5770);
and U7605 (N_7605,N_4872,N_5175);
nor U7606 (N_7606,N_5610,N_4713);
or U7607 (N_7607,N_4177,N_5546);
or U7608 (N_7608,N_4099,N_4585);
or U7609 (N_7609,N_5388,N_5736);
and U7610 (N_7610,N_5524,N_5221);
nor U7611 (N_7611,N_4777,N_5612);
nor U7612 (N_7612,N_5917,N_5682);
and U7613 (N_7613,N_5837,N_5506);
and U7614 (N_7614,N_4612,N_5004);
or U7615 (N_7615,N_4257,N_4185);
nor U7616 (N_7616,N_5610,N_4270);
nand U7617 (N_7617,N_4745,N_4650);
or U7618 (N_7618,N_4139,N_4046);
nand U7619 (N_7619,N_4768,N_5896);
xor U7620 (N_7620,N_4744,N_5780);
or U7621 (N_7621,N_4866,N_5601);
and U7622 (N_7622,N_4448,N_5382);
xor U7623 (N_7623,N_5503,N_5526);
or U7624 (N_7624,N_4022,N_5318);
nor U7625 (N_7625,N_5275,N_5081);
xor U7626 (N_7626,N_5124,N_4811);
nor U7627 (N_7627,N_4595,N_5338);
nand U7628 (N_7628,N_4282,N_5530);
xnor U7629 (N_7629,N_4833,N_5173);
nand U7630 (N_7630,N_5275,N_4427);
nor U7631 (N_7631,N_5155,N_5459);
nor U7632 (N_7632,N_4165,N_4715);
xnor U7633 (N_7633,N_5791,N_5201);
nand U7634 (N_7634,N_5205,N_4303);
or U7635 (N_7635,N_4889,N_5451);
nand U7636 (N_7636,N_5128,N_4867);
and U7637 (N_7637,N_4964,N_5890);
xnor U7638 (N_7638,N_5026,N_5778);
xor U7639 (N_7639,N_4571,N_5106);
or U7640 (N_7640,N_5252,N_4939);
nor U7641 (N_7641,N_4032,N_4326);
and U7642 (N_7642,N_5334,N_5452);
or U7643 (N_7643,N_5930,N_4947);
nand U7644 (N_7644,N_5015,N_5997);
or U7645 (N_7645,N_4056,N_5072);
nor U7646 (N_7646,N_4046,N_4013);
xor U7647 (N_7647,N_5482,N_5658);
nor U7648 (N_7648,N_4103,N_5970);
and U7649 (N_7649,N_4101,N_4555);
xor U7650 (N_7650,N_4218,N_5485);
nor U7651 (N_7651,N_5945,N_5585);
nand U7652 (N_7652,N_5359,N_4342);
nor U7653 (N_7653,N_4223,N_5956);
xor U7654 (N_7654,N_4492,N_5596);
xor U7655 (N_7655,N_4677,N_4133);
or U7656 (N_7656,N_5037,N_5283);
or U7657 (N_7657,N_4191,N_4413);
or U7658 (N_7658,N_4017,N_4877);
xor U7659 (N_7659,N_4691,N_5749);
or U7660 (N_7660,N_4556,N_4198);
and U7661 (N_7661,N_5470,N_4610);
or U7662 (N_7662,N_5290,N_5079);
nand U7663 (N_7663,N_5192,N_5034);
nand U7664 (N_7664,N_5774,N_4694);
and U7665 (N_7665,N_5630,N_5155);
nor U7666 (N_7666,N_5187,N_5654);
and U7667 (N_7667,N_5232,N_4952);
nand U7668 (N_7668,N_5547,N_4656);
and U7669 (N_7669,N_5318,N_4403);
and U7670 (N_7670,N_5448,N_4316);
xnor U7671 (N_7671,N_5647,N_5271);
nand U7672 (N_7672,N_5996,N_4919);
nand U7673 (N_7673,N_5915,N_4806);
nor U7674 (N_7674,N_5288,N_5660);
or U7675 (N_7675,N_5821,N_4969);
or U7676 (N_7676,N_5069,N_5957);
nor U7677 (N_7677,N_5054,N_5431);
nand U7678 (N_7678,N_5138,N_5066);
or U7679 (N_7679,N_4498,N_5859);
nor U7680 (N_7680,N_4334,N_5694);
xnor U7681 (N_7681,N_5879,N_4340);
xnor U7682 (N_7682,N_5503,N_4055);
or U7683 (N_7683,N_5742,N_5607);
and U7684 (N_7684,N_4739,N_4419);
and U7685 (N_7685,N_4431,N_5457);
nand U7686 (N_7686,N_5390,N_5157);
and U7687 (N_7687,N_4706,N_5531);
xor U7688 (N_7688,N_5073,N_4602);
and U7689 (N_7689,N_5130,N_4500);
and U7690 (N_7690,N_5545,N_4966);
xnor U7691 (N_7691,N_5074,N_5856);
nand U7692 (N_7692,N_5787,N_5194);
nand U7693 (N_7693,N_5856,N_4592);
or U7694 (N_7694,N_5212,N_4511);
and U7695 (N_7695,N_5120,N_5585);
and U7696 (N_7696,N_4063,N_4166);
nor U7697 (N_7697,N_4331,N_4853);
and U7698 (N_7698,N_4033,N_4437);
nor U7699 (N_7699,N_5969,N_5127);
xor U7700 (N_7700,N_5469,N_5704);
or U7701 (N_7701,N_4131,N_4399);
or U7702 (N_7702,N_5677,N_5540);
nor U7703 (N_7703,N_5078,N_4169);
xnor U7704 (N_7704,N_5352,N_4288);
nor U7705 (N_7705,N_5875,N_4870);
and U7706 (N_7706,N_5788,N_4950);
nor U7707 (N_7707,N_4930,N_4202);
or U7708 (N_7708,N_4558,N_5247);
nand U7709 (N_7709,N_4570,N_4072);
nor U7710 (N_7710,N_5967,N_5191);
and U7711 (N_7711,N_5503,N_5316);
xor U7712 (N_7712,N_5318,N_4759);
xor U7713 (N_7713,N_5948,N_5013);
xnor U7714 (N_7714,N_4142,N_4380);
or U7715 (N_7715,N_4018,N_5023);
nand U7716 (N_7716,N_5238,N_4652);
or U7717 (N_7717,N_4981,N_5678);
nand U7718 (N_7718,N_5351,N_4983);
or U7719 (N_7719,N_5817,N_4378);
and U7720 (N_7720,N_5902,N_5562);
nor U7721 (N_7721,N_5864,N_5396);
nor U7722 (N_7722,N_4770,N_4467);
nor U7723 (N_7723,N_4643,N_4607);
nor U7724 (N_7724,N_4515,N_4319);
nand U7725 (N_7725,N_4388,N_4041);
nor U7726 (N_7726,N_5104,N_5252);
nor U7727 (N_7727,N_5467,N_5779);
or U7728 (N_7728,N_5850,N_4426);
xnor U7729 (N_7729,N_5503,N_4699);
or U7730 (N_7730,N_5966,N_5292);
or U7731 (N_7731,N_4733,N_5625);
nand U7732 (N_7732,N_4469,N_4352);
or U7733 (N_7733,N_5849,N_4879);
nand U7734 (N_7734,N_4344,N_5721);
xor U7735 (N_7735,N_5174,N_4351);
or U7736 (N_7736,N_5550,N_4427);
nand U7737 (N_7737,N_5578,N_4107);
nand U7738 (N_7738,N_5652,N_5181);
nand U7739 (N_7739,N_5394,N_4590);
nor U7740 (N_7740,N_5336,N_5833);
nor U7741 (N_7741,N_5916,N_4468);
or U7742 (N_7742,N_5928,N_5963);
xor U7743 (N_7743,N_4363,N_4935);
nor U7744 (N_7744,N_5660,N_5377);
nand U7745 (N_7745,N_5764,N_4915);
or U7746 (N_7746,N_5209,N_5169);
nor U7747 (N_7747,N_4379,N_4089);
and U7748 (N_7748,N_5750,N_4549);
nor U7749 (N_7749,N_5719,N_4049);
nor U7750 (N_7750,N_4099,N_5140);
nand U7751 (N_7751,N_5198,N_4992);
xor U7752 (N_7752,N_5027,N_4983);
and U7753 (N_7753,N_4965,N_5248);
nor U7754 (N_7754,N_4700,N_4895);
nand U7755 (N_7755,N_5098,N_5751);
xor U7756 (N_7756,N_5462,N_4026);
and U7757 (N_7757,N_4617,N_5193);
and U7758 (N_7758,N_4073,N_4387);
nor U7759 (N_7759,N_5488,N_4953);
nor U7760 (N_7760,N_4875,N_4879);
or U7761 (N_7761,N_4711,N_5862);
or U7762 (N_7762,N_4222,N_4653);
and U7763 (N_7763,N_5581,N_5874);
and U7764 (N_7764,N_4663,N_5638);
or U7765 (N_7765,N_5368,N_4312);
nor U7766 (N_7766,N_5585,N_5604);
or U7767 (N_7767,N_5085,N_4157);
xor U7768 (N_7768,N_5010,N_4996);
nor U7769 (N_7769,N_5277,N_5271);
xor U7770 (N_7770,N_5332,N_5898);
xor U7771 (N_7771,N_5659,N_4146);
xnor U7772 (N_7772,N_5242,N_5447);
or U7773 (N_7773,N_4985,N_5244);
or U7774 (N_7774,N_4342,N_4724);
nor U7775 (N_7775,N_4775,N_4796);
or U7776 (N_7776,N_5793,N_4935);
nor U7777 (N_7777,N_4865,N_4179);
nand U7778 (N_7778,N_4424,N_4441);
nor U7779 (N_7779,N_5609,N_4856);
and U7780 (N_7780,N_4143,N_4916);
nor U7781 (N_7781,N_5452,N_4332);
nand U7782 (N_7782,N_5406,N_5019);
nand U7783 (N_7783,N_4210,N_4441);
or U7784 (N_7784,N_5147,N_5019);
nand U7785 (N_7785,N_4869,N_5916);
xor U7786 (N_7786,N_4704,N_5969);
nand U7787 (N_7787,N_4393,N_4328);
and U7788 (N_7788,N_5522,N_4701);
nand U7789 (N_7789,N_5676,N_4581);
xnor U7790 (N_7790,N_4788,N_5105);
or U7791 (N_7791,N_4276,N_5510);
or U7792 (N_7792,N_5161,N_5948);
nor U7793 (N_7793,N_5380,N_4610);
and U7794 (N_7794,N_5759,N_5315);
and U7795 (N_7795,N_4538,N_5138);
xnor U7796 (N_7796,N_4564,N_5970);
or U7797 (N_7797,N_5161,N_5541);
nor U7798 (N_7798,N_4697,N_4290);
and U7799 (N_7799,N_5254,N_4820);
and U7800 (N_7800,N_5555,N_4450);
xnor U7801 (N_7801,N_4513,N_5331);
or U7802 (N_7802,N_4421,N_5020);
and U7803 (N_7803,N_4378,N_4140);
or U7804 (N_7804,N_4965,N_5530);
xnor U7805 (N_7805,N_4287,N_5455);
nor U7806 (N_7806,N_5689,N_5907);
nand U7807 (N_7807,N_5980,N_5864);
nor U7808 (N_7808,N_5426,N_4119);
or U7809 (N_7809,N_5998,N_5123);
nand U7810 (N_7810,N_5574,N_4813);
xnor U7811 (N_7811,N_4849,N_5597);
nor U7812 (N_7812,N_4519,N_5626);
nand U7813 (N_7813,N_4283,N_5989);
and U7814 (N_7814,N_5456,N_4333);
xor U7815 (N_7815,N_5601,N_5419);
xor U7816 (N_7816,N_4852,N_4376);
or U7817 (N_7817,N_5463,N_5460);
nor U7818 (N_7818,N_4867,N_4279);
or U7819 (N_7819,N_5587,N_5435);
xnor U7820 (N_7820,N_4498,N_5906);
xnor U7821 (N_7821,N_4564,N_5447);
and U7822 (N_7822,N_4043,N_4731);
nand U7823 (N_7823,N_4153,N_5008);
or U7824 (N_7824,N_4366,N_4044);
nor U7825 (N_7825,N_4089,N_4913);
nand U7826 (N_7826,N_4211,N_4212);
and U7827 (N_7827,N_4108,N_4756);
xnor U7828 (N_7828,N_5325,N_5096);
and U7829 (N_7829,N_5984,N_4852);
xor U7830 (N_7830,N_4718,N_4813);
and U7831 (N_7831,N_4055,N_4563);
xnor U7832 (N_7832,N_4081,N_4840);
xnor U7833 (N_7833,N_4978,N_5442);
nor U7834 (N_7834,N_4322,N_5545);
or U7835 (N_7835,N_4243,N_4593);
or U7836 (N_7836,N_5567,N_5899);
nand U7837 (N_7837,N_4978,N_5046);
xnor U7838 (N_7838,N_4324,N_5407);
or U7839 (N_7839,N_4628,N_5636);
nand U7840 (N_7840,N_4683,N_5375);
nand U7841 (N_7841,N_5718,N_4394);
or U7842 (N_7842,N_5272,N_4412);
nor U7843 (N_7843,N_5078,N_5092);
or U7844 (N_7844,N_5041,N_4349);
nor U7845 (N_7845,N_4499,N_5676);
and U7846 (N_7846,N_4619,N_5796);
nor U7847 (N_7847,N_4904,N_5702);
nand U7848 (N_7848,N_4570,N_5200);
xnor U7849 (N_7849,N_5463,N_4159);
nor U7850 (N_7850,N_4894,N_5174);
or U7851 (N_7851,N_4178,N_5609);
or U7852 (N_7852,N_5632,N_4071);
or U7853 (N_7853,N_5427,N_4971);
xnor U7854 (N_7854,N_5756,N_4130);
or U7855 (N_7855,N_5071,N_5538);
xor U7856 (N_7856,N_5892,N_4396);
and U7857 (N_7857,N_5520,N_5078);
xor U7858 (N_7858,N_4744,N_4374);
and U7859 (N_7859,N_4727,N_4415);
nand U7860 (N_7860,N_4340,N_5089);
nor U7861 (N_7861,N_5637,N_5082);
nor U7862 (N_7862,N_5936,N_4766);
or U7863 (N_7863,N_4841,N_4181);
nor U7864 (N_7864,N_5902,N_5086);
xnor U7865 (N_7865,N_4329,N_5235);
xnor U7866 (N_7866,N_5885,N_5123);
nor U7867 (N_7867,N_4314,N_5905);
nor U7868 (N_7868,N_4418,N_5783);
nor U7869 (N_7869,N_5128,N_4745);
nand U7870 (N_7870,N_5941,N_4106);
nor U7871 (N_7871,N_5049,N_4279);
and U7872 (N_7872,N_4499,N_4554);
xor U7873 (N_7873,N_4674,N_4858);
nor U7874 (N_7874,N_4334,N_5159);
and U7875 (N_7875,N_5691,N_4017);
nand U7876 (N_7876,N_5152,N_4307);
or U7877 (N_7877,N_4042,N_5618);
nand U7878 (N_7878,N_4928,N_5029);
nor U7879 (N_7879,N_5765,N_4434);
or U7880 (N_7880,N_4208,N_4819);
or U7881 (N_7881,N_5445,N_5123);
xor U7882 (N_7882,N_4659,N_5650);
or U7883 (N_7883,N_5385,N_5000);
xnor U7884 (N_7884,N_4953,N_5688);
xnor U7885 (N_7885,N_5747,N_5858);
xor U7886 (N_7886,N_5386,N_4851);
xnor U7887 (N_7887,N_5607,N_5851);
nand U7888 (N_7888,N_5811,N_5807);
nand U7889 (N_7889,N_5084,N_4099);
nand U7890 (N_7890,N_4791,N_4900);
nand U7891 (N_7891,N_5465,N_4743);
and U7892 (N_7892,N_4171,N_5785);
and U7893 (N_7893,N_4061,N_4990);
xnor U7894 (N_7894,N_5052,N_5337);
xor U7895 (N_7895,N_4692,N_4377);
xnor U7896 (N_7896,N_4988,N_5316);
and U7897 (N_7897,N_4046,N_5131);
and U7898 (N_7898,N_5539,N_4298);
nand U7899 (N_7899,N_5330,N_5026);
xor U7900 (N_7900,N_5449,N_5142);
or U7901 (N_7901,N_4846,N_4214);
nand U7902 (N_7902,N_5105,N_5727);
xor U7903 (N_7903,N_4842,N_4582);
nand U7904 (N_7904,N_4202,N_5412);
nor U7905 (N_7905,N_4109,N_4282);
xnor U7906 (N_7906,N_5281,N_4673);
xor U7907 (N_7907,N_4724,N_4626);
or U7908 (N_7908,N_4363,N_5475);
nand U7909 (N_7909,N_5472,N_5989);
or U7910 (N_7910,N_4227,N_4789);
nor U7911 (N_7911,N_5018,N_5672);
and U7912 (N_7912,N_5842,N_4681);
or U7913 (N_7913,N_4279,N_5035);
or U7914 (N_7914,N_4989,N_5778);
and U7915 (N_7915,N_5146,N_5695);
nor U7916 (N_7916,N_5292,N_4791);
or U7917 (N_7917,N_4845,N_5671);
or U7918 (N_7918,N_5378,N_4850);
nand U7919 (N_7919,N_4035,N_5049);
and U7920 (N_7920,N_4577,N_4642);
xnor U7921 (N_7921,N_5557,N_4451);
nor U7922 (N_7922,N_5841,N_5200);
or U7923 (N_7923,N_5925,N_4519);
nor U7924 (N_7924,N_4251,N_4587);
and U7925 (N_7925,N_5943,N_5397);
xnor U7926 (N_7926,N_5217,N_5330);
and U7927 (N_7927,N_4895,N_5508);
nand U7928 (N_7928,N_5545,N_4213);
and U7929 (N_7929,N_4912,N_4811);
nand U7930 (N_7930,N_4198,N_4919);
xor U7931 (N_7931,N_4118,N_4394);
or U7932 (N_7932,N_4411,N_4061);
nor U7933 (N_7933,N_5457,N_4555);
xnor U7934 (N_7934,N_4590,N_4397);
nand U7935 (N_7935,N_5378,N_5069);
nor U7936 (N_7936,N_5776,N_5162);
nand U7937 (N_7937,N_5485,N_5719);
and U7938 (N_7938,N_5518,N_4291);
xnor U7939 (N_7939,N_4487,N_4325);
nor U7940 (N_7940,N_5128,N_5010);
nor U7941 (N_7941,N_5317,N_4613);
xnor U7942 (N_7942,N_5662,N_5283);
nand U7943 (N_7943,N_5809,N_5410);
nor U7944 (N_7944,N_4271,N_5254);
or U7945 (N_7945,N_5181,N_5085);
and U7946 (N_7946,N_5063,N_5915);
xor U7947 (N_7947,N_4496,N_4300);
xor U7948 (N_7948,N_4690,N_4777);
and U7949 (N_7949,N_4613,N_5760);
nand U7950 (N_7950,N_4542,N_5891);
xnor U7951 (N_7951,N_4286,N_5487);
xor U7952 (N_7952,N_4200,N_4851);
nor U7953 (N_7953,N_4838,N_5772);
xor U7954 (N_7954,N_5312,N_5375);
or U7955 (N_7955,N_4383,N_4791);
and U7956 (N_7956,N_5655,N_4205);
nor U7957 (N_7957,N_5072,N_5764);
xor U7958 (N_7958,N_5167,N_5638);
nor U7959 (N_7959,N_4450,N_4812);
xor U7960 (N_7960,N_4304,N_4094);
or U7961 (N_7961,N_4588,N_4634);
xor U7962 (N_7962,N_5015,N_4336);
and U7963 (N_7963,N_4579,N_5088);
nand U7964 (N_7964,N_5834,N_5385);
nor U7965 (N_7965,N_5332,N_5758);
nor U7966 (N_7966,N_5879,N_5907);
nor U7967 (N_7967,N_5473,N_4809);
or U7968 (N_7968,N_4403,N_4282);
or U7969 (N_7969,N_5254,N_5920);
xnor U7970 (N_7970,N_5917,N_4088);
nor U7971 (N_7971,N_5470,N_4915);
and U7972 (N_7972,N_4912,N_5403);
nor U7973 (N_7973,N_5756,N_5753);
xor U7974 (N_7974,N_5591,N_5042);
nand U7975 (N_7975,N_4505,N_4040);
nor U7976 (N_7976,N_4839,N_5618);
nor U7977 (N_7977,N_4862,N_4939);
or U7978 (N_7978,N_4538,N_4763);
nand U7979 (N_7979,N_5156,N_4669);
xnor U7980 (N_7980,N_4273,N_4211);
nand U7981 (N_7981,N_4622,N_5127);
or U7982 (N_7982,N_5471,N_4068);
nor U7983 (N_7983,N_5957,N_4582);
and U7984 (N_7984,N_5649,N_4504);
nor U7985 (N_7985,N_4232,N_4366);
or U7986 (N_7986,N_4005,N_4097);
or U7987 (N_7987,N_4481,N_5821);
and U7988 (N_7988,N_5764,N_4538);
and U7989 (N_7989,N_4987,N_4018);
xnor U7990 (N_7990,N_4332,N_4735);
nor U7991 (N_7991,N_5411,N_5094);
xor U7992 (N_7992,N_4789,N_4403);
and U7993 (N_7993,N_5087,N_5873);
and U7994 (N_7994,N_5494,N_4398);
nand U7995 (N_7995,N_4357,N_5925);
nand U7996 (N_7996,N_4392,N_4334);
nand U7997 (N_7997,N_4328,N_5650);
nor U7998 (N_7998,N_5632,N_4175);
or U7999 (N_7999,N_4449,N_5600);
or U8000 (N_8000,N_7012,N_7099);
nor U8001 (N_8001,N_6342,N_6164);
or U8002 (N_8002,N_6626,N_6753);
xor U8003 (N_8003,N_7866,N_7686);
or U8004 (N_8004,N_6155,N_6898);
nand U8005 (N_8005,N_6369,N_7248);
nand U8006 (N_8006,N_7245,N_7307);
and U8007 (N_8007,N_7218,N_7938);
nor U8008 (N_8008,N_7534,N_7903);
nand U8009 (N_8009,N_6226,N_7716);
or U8010 (N_8010,N_7732,N_6008);
nand U8011 (N_8011,N_6782,N_7035);
or U8012 (N_8012,N_6133,N_7522);
xor U8013 (N_8013,N_7382,N_6525);
xnor U8014 (N_8014,N_6653,N_7525);
and U8015 (N_8015,N_7396,N_7523);
nand U8016 (N_8016,N_6070,N_7741);
xnor U8017 (N_8017,N_6655,N_6946);
nor U8018 (N_8018,N_7119,N_7558);
nor U8019 (N_8019,N_7477,N_6681);
xnor U8020 (N_8020,N_6746,N_7833);
xor U8021 (N_8021,N_6974,N_7220);
and U8022 (N_8022,N_6509,N_6494);
or U8023 (N_8023,N_7536,N_6751);
or U8024 (N_8024,N_7424,N_7851);
nor U8025 (N_8025,N_6693,N_7830);
xnor U8026 (N_8026,N_6086,N_7438);
and U8027 (N_8027,N_6855,N_6214);
or U8028 (N_8028,N_6059,N_6588);
nor U8029 (N_8029,N_7472,N_7392);
or U8030 (N_8030,N_7189,N_6606);
or U8031 (N_8031,N_7963,N_6137);
or U8032 (N_8032,N_6835,N_6194);
or U8033 (N_8033,N_7107,N_6540);
or U8034 (N_8034,N_7004,N_7764);
and U8035 (N_8035,N_7071,N_6654);
and U8036 (N_8036,N_6221,N_7208);
or U8037 (N_8037,N_6850,N_7855);
nor U8038 (N_8038,N_7212,N_7291);
and U8039 (N_8039,N_6297,N_7226);
nand U8040 (N_8040,N_6901,N_6429);
or U8041 (N_8041,N_7805,N_6403);
and U8042 (N_8042,N_6911,N_6439);
nand U8043 (N_8043,N_6293,N_6852);
xor U8044 (N_8044,N_7254,N_7919);
and U8045 (N_8045,N_7677,N_7806);
nor U8046 (N_8046,N_6413,N_7784);
xnor U8047 (N_8047,N_7801,N_6251);
nor U8048 (N_8048,N_6119,N_6033);
xor U8049 (N_8049,N_7809,N_7352);
or U8050 (N_8050,N_6092,N_7211);
and U8051 (N_8051,N_7090,N_7600);
or U8052 (N_8052,N_6093,N_7386);
nand U8053 (N_8053,N_7023,N_6388);
and U8054 (N_8054,N_7264,N_7846);
or U8055 (N_8055,N_7783,N_7008);
and U8056 (N_8056,N_7973,N_6064);
nand U8057 (N_8057,N_6382,N_7769);
xnor U8058 (N_8058,N_6202,N_6205);
and U8059 (N_8059,N_7387,N_6153);
nand U8060 (N_8060,N_6181,N_7638);
xor U8061 (N_8061,N_7876,N_6673);
and U8062 (N_8062,N_7708,N_7966);
xor U8063 (N_8063,N_6377,N_7130);
nor U8064 (N_8064,N_6818,N_6283);
nand U8065 (N_8065,N_6604,N_7055);
or U8066 (N_8066,N_7104,N_7391);
and U8067 (N_8067,N_7077,N_6068);
xnor U8068 (N_8068,N_7648,N_6727);
and U8069 (N_8069,N_6415,N_7798);
or U8070 (N_8070,N_7453,N_7166);
and U8071 (N_8071,N_7637,N_7429);
or U8072 (N_8072,N_7026,N_6146);
nor U8073 (N_8073,N_6278,N_6858);
and U8074 (N_8074,N_7021,N_7549);
nand U8075 (N_8075,N_6501,N_6065);
and U8076 (N_8076,N_7383,N_7969);
nand U8077 (N_8077,N_7298,N_6284);
or U8078 (N_8078,N_6275,N_6612);
and U8079 (N_8079,N_7405,N_6390);
or U8080 (N_8080,N_7266,N_6322);
and U8081 (N_8081,N_6058,N_6291);
xnor U8082 (N_8082,N_6255,N_7149);
and U8083 (N_8083,N_6699,N_7188);
or U8084 (N_8084,N_6476,N_7230);
and U8085 (N_8085,N_6748,N_6618);
and U8086 (N_8086,N_7002,N_6016);
xor U8087 (N_8087,N_6042,N_7222);
nand U8088 (N_8088,N_7605,N_7569);
or U8089 (N_8089,N_6201,N_6270);
xnor U8090 (N_8090,N_6338,N_7874);
and U8091 (N_8091,N_7738,N_6096);
xor U8092 (N_8092,N_7714,N_7645);
and U8093 (N_8093,N_6491,N_6661);
or U8094 (N_8094,N_7904,N_6250);
or U8095 (N_8095,N_6922,N_6504);
nand U8096 (N_8096,N_7895,N_6453);
xnor U8097 (N_8097,N_6641,N_7807);
nand U8098 (N_8098,N_6507,N_6132);
xnor U8099 (N_8099,N_7095,N_6109);
and U8100 (N_8100,N_6582,N_6812);
and U8101 (N_8101,N_6515,N_7554);
nand U8102 (N_8102,N_7029,N_7682);
nand U8103 (N_8103,N_7467,N_6943);
nand U8104 (N_8104,N_7186,N_6502);
or U8105 (N_8105,N_7848,N_6028);
and U8106 (N_8106,N_7864,N_7819);
nor U8107 (N_8107,N_7878,N_7482);
xnor U8108 (N_8108,N_7260,N_6517);
xor U8109 (N_8109,N_6066,N_6303);
nand U8110 (N_8110,N_7345,N_7237);
or U8111 (N_8111,N_6667,N_6021);
and U8112 (N_8112,N_7681,N_6671);
or U8113 (N_8113,N_6258,N_7193);
nor U8114 (N_8114,N_6268,N_7883);
xnor U8115 (N_8115,N_6956,N_6315);
nor U8116 (N_8116,N_6822,N_6728);
nor U8117 (N_8117,N_6643,N_6682);
nor U8118 (N_8118,N_7421,N_7794);
xor U8119 (N_8119,N_7695,N_6634);
xor U8120 (N_8120,N_6873,N_7700);
nand U8121 (N_8121,N_6983,N_6075);
nor U8122 (N_8122,N_7852,N_6454);
nand U8123 (N_8123,N_6773,N_7824);
nand U8124 (N_8124,N_7688,N_7750);
and U8125 (N_8125,N_7793,N_7684);
or U8126 (N_8126,N_6804,N_6039);
nand U8127 (N_8127,N_6496,N_6934);
and U8128 (N_8128,N_6617,N_6740);
and U8129 (N_8129,N_6077,N_6690);
xor U8130 (N_8130,N_6849,N_6761);
nand U8131 (N_8131,N_6677,N_7669);
nor U8132 (N_8132,N_7013,N_7484);
nor U8133 (N_8133,N_6100,N_6289);
or U8134 (N_8134,N_7827,N_7584);
nand U8135 (N_8135,N_7845,N_7885);
xnor U8136 (N_8136,N_7358,N_6900);
and U8137 (N_8137,N_6586,N_6170);
nor U8138 (N_8138,N_7890,N_7555);
and U8139 (N_8139,N_6490,N_7325);
and U8140 (N_8140,N_6431,N_7713);
or U8141 (N_8141,N_6723,N_7849);
and U8142 (N_8142,N_7236,N_6295);
and U8143 (N_8143,N_6862,N_7834);
or U8144 (N_8144,N_6895,N_7347);
nand U8145 (N_8145,N_7642,N_7504);
nand U8146 (N_8146,N_6487,N_6354);
nand U8147 (N_8147,N_6788,N_6584);
and U8148 (N_8148,N_7984,N_6676);
xnor U8149 (N_8149,N_6393,N_7458);
and U8150 (N_8150,N_7986,N_7277);
and U8151 (N_8151,N_6962,N_7777);
xor U8152 (N_8152,N_7877,N_7436);
or U8153 (N_8153,N_7418,N_7944);
nor U8154 (N_8154,N_6704,N_7346);
nor U8155 (N_8155,N_6921,N_6763);
nand U8156 (N_8156,N_6513,N_7658);
or U8157 (N_8157,N_7698,N_7153);
or U8158 (N_8158,N_6929,N_6874);
xor U8159 (N_8159,N_6449,N_6142);
or U8160 (N_8160,N_7094,N_6144);
xnor U8161 (N_8161,N_6152,N_6233);
nand U8162 (N_8162,N_7295,N_6422);
or U8163 (N_8163,N_6022,N_7072);
or U8164 (N_8164,N_6433,N_7152);
nand U8165 (N_8165,N_7056,N_6477);
nor U8166 (N_8166,N_6769,N_7991);
nor U8167 (N_8167,N_6854,N_7974);
or U8168 (N_8168,N_6495,N_7279);
nor U8169 (N_8169,N_6814,N_6915);
and U8170 (N_8170,N_7620,N_6813);
nor U8171 (N_8171,N_7593,N_6566);
or U8172 (N_8172,N_7164,N_6972);
nor U8173 (N_8173,N_6599,N_7433);
xnor U8174 (N_8174,N_6656,N_6380);
xnor U8175 (N_8175,N_7838,N_6242);
or U8176 (N_8176,N_7893,N_6640);
nand U8177 (N_8177,N_7694,N_6691);
or U8178 (N_8178,N_6460,N_7616);
and U8179 (N_8179,N_6330,N_6914);
and U8180 (N_8180,N_6309,N_6452);
xor U8181 (N_8181,N_6172,N_6466);
nor U8182 (N_8182,N_7921,N_7626);
nand U8183 (N_8183,N_7790,N_7262);
and U8184 (N_8184,N_6939,N_6731);
or U8185 (N_8185,N_7803,N_7203);
nor U8186 (N_8186,N_7887,N_6421);
or U8187 (N_8187,N_6179,N_6623);
nand U8188 (N_8188,N_6680,N_7144);
and U8189 (N_8189,N_6547,N_7630);
nand U8190 (N_8190,N_6907,N_6944);
xnor U8191 (N_8191,N_7967,N_6969);
nand U8192 (N_8192,N_7689,N_6530);
xnor U8193 (N_8193,N_7712,N_7194);
xor U8194 (N_8194,N_6206,N_7321);
xnor U8195 (N_8195,N_6948,N_6591);
or U8196 (N_8196,N_6356,N_6197);
xnor U8197 (N_8197,N_7551,N_7242);
or U8198 (N_8198,N_6572,N_6475);
or U8199 (N_8199,N_6575,N_7303);
and U8200 (N_8200,N_7380,N_7081);
nor U8201 (N_8201,N_7489,N_6381);
nor U8202 (N_8202,N_6000,N_7430);
xor U8203 (N_8203,N_7531,N_7859);
nand U8204 (N_8204,N_7267,N_7441);
nand U8205 (N_8205,N_7509,N_6050);
nand U8206 (N_8206,N_7412,N_7755);
or U8207 (N_8207,N_6244,N_6310);
and U8208 (N_8208,N_7579,N_6138);
nand U8209 (N_8209,N_7044,N_6364);
or U8210 (N_8210,N_7749,N_7332);
and U8211 (N_8211,N_7093,N_6407);
or U8212 (N_8212,N_7080,N_6658);
nand U8213 (N_8213,N_6965,N_6002);
nand U8214 (N_8214,N_7941,N_7711);
nand U8215 (N_8215,N_6807,N_7381);
xor U8216 (N_8216,N_7572,N_7324);
xor U8217 (N_8217,N_6510,N_7238);
nand U8218 (N_8218,N_7117,N_7936);
or U8219 (N_8219,N_7273,N_7180);
nand U8220 (N_8220,N_7082,N_6684);
and U8221 (N_8221,N_6889,N_6130);
nand U8222 (N_8222,N_7888,N_7257);
xor U8223 (N_8223,N_6084,N_6327);
xnor U8224 (N_8224,N_7223,N_6955);
and U8225 (N_8225,N_7280,N_7213);
and U8226 (N_8226,N_7914,N_7653);
and U8227 (N_8227,N_6714,N_7719);
and U8228 (N_8228,N_6760,N_7519);
or U8229 (N_8229,N_7483,N_6314);
nand U8230 (N_8230,N_7891,N_6389);
xnor U8231 (N_8231,N_6605,N_7882);
nor U8232 (N_8232,N_7995,N_7444);
nand U8233 (N_8233,N_7802,N_7401);
nor U8234 (N_8234,N_6775,N_6443);
and U8235 (N_8235,N_7249,N_6892);
or U8236 (N_8236,N_6593,N_6902);
nor U8237 (N_8237,N_6425,N_6537);
nor U8238 (N_8238,N_6869,N_6712);
xnor U8239 (N_8239,N_7825,N_7502);
and U8240 (N_8240,N_7108,N_6912);
or U8241 (N_8241,N_6536,N_6811);
or U8242 (N_8242,N_6660,N_7114);
nand U8243 (N_8243,N_6230,N_6808);
and U8244 (N_8244,N_7058,N_6702);
or U8245 (N_8245,N_7410,N_7420);
nand U8246 (N_8246,N_6675,N_6235);
or U8247 (N_8247,N_6007,N_7491);
and U8248 (N_8248,N_7946,N_7678);
xnor U8249 (N_8249,N_7590,N_6896);
nor U8250 (N_8250,N_7167,N_6821);
xor U8251 (N_8251,N_7020,N_7028);
nand U8252 (N_8252,N_7661,N_6737);
nand U8253 (N_8253,N_7751,N_7469);
and U8254 (N_8254,N_7473,N_6734);
xor U8255 (N_8255,N_7479,N_7190);
and U8256 (N_8256,N_6228,N_7317);
xor U8257 (N_8257,N_7357,N_6282);
nand U8258 (N_8258,N_7539,N_6175);
xor U8259 (N_8259,N_7870,N_6952);
xor U8260 (N_8260,N_6920,N_7553);
or U8261 (N_8261,N_7364,N_6074);
nor U8262 (N_8262,N_7770,N_7564);
nand U8263 (N_8263,N_6925,N_6827);
nand U8264 (N_8264,N_6333,N_7290);
or U8265 (N_8265,N_7550,N_6880);
nor U8266 (N_8266,N_7591,N_6707);
nor U8267 (N_8267,N_7319,N_6145);
nand U8268 (N_8268,N_6512,N_7097);
and U8269 (N_8269,N_7624,N_7414);
xor U8270 (N_8270,N_6608,N_6385);
nor U8271 (N_8271,N_7641,N_7463);
nand U8272 (N_8272,N_6110,N_7943);
nand U8273 (N_8273,N_6999,N_7475);
and U8274 (N_8274,N_7202,N_7465);
nand U8275 (N_8275,N_7087,N_7360);
nor U8276 (N_8276,N_7983,N_6287);
nand U8277 (N_8277,N_6456,N_7792);
nor U8278 (N_8278,N_6447,N_7393);
and U8279 (N_8279,N_7089,N_7693);
xor U8280 (N_8280,N_6882,N_6531);
or U8281 (N_8281,N_6072,N_7231);
nor U8282 (N_8282,N_6474,N_6908);
nand U8283 (N_8283,N_7384,N_6799);
xnor U8284 (N_8284,N_7690,N_7448);
xnor U8285 (N_8285,N_6106,N_6638);
or U8286 (N_8286,N_6844,N_6749);
xor U8287 (N_8287,N_6919,N_6082);
or U8288 (N_8288,N_7659,N_7839);
xnor U8289 (N_8289,N_6200,N_7623);
and U8290 (N_8290,N_7906,N_7379);
nand U8291 (N_8291,N_6135,N_6624);
or U8292 (N_8292,N_7990,N_7141);
nand U8293 (N_8293,N_7631,N_7156);
or U8294 (N_8294,N_7667,N_6906);
nand U8295 (N_8295,N_7437,N_7568);
xor U8296 (N_8296,N_6781,N_7910);
nand U8297 (N_8297,N_7820,N_7111);
or U8298 (N_8298,N_7768,N_6426);
nor U8299 (N_8299,N_6971,N_7588);
or U8300 (N_8300,N_7432,N_7251);
and U8301 (N_8301,N_6635,N_6321);
xnor U8302 (N_8302,N_6355,N_6428);
xor U8303 (N_8303,N_6863,N_7622);
and U8304 (N_8304,N_6055,N_6716);
nor U8305 (N_8305,N_7204,N_7070);
or U8306 (N_8306,N_6815,N_7704);
xnor U8307 (N_8307,N_6669,N_7278);
or U8308 (N_8308,N_7778,N_6750);
or U8309 (N_8309,N_6089,N_7235);
nand U8310 (N_8310,N_7710,N_6967);
nor U8311 (N_8311,N_6448,N_6442);
and U8312 (N_8312,N_6613,N_6402);
or U8313 (N_8313,N_7901,N_6725);
xor U8314 (N_8314,N_7284,N_6348);
xor U8315 (N_8315,N_7499,N_6825);
nor U8316 (N_8316,N_7581,N_7275);
nor U8317 (N_8317,N_6549,N_7655);
nor U8318 (N_8318,N_6829,N_6410);
or U8319 (N_8319,N_7179,N_6427);
and U8320 (N_8320,N_6409,N_6195);
nand U8321 (N_8321,N_6719,N_6933);
nor U8322 (N_8322,N_7999,N_7935);
nor U8323 (N_8323,N_7971,N_7181);
xor U8324 (N_8324,N_7857,N_6806);
nor U8325 (N_8325,N_7942,N_6583);
nand U8326 (N_8326,N_7385,N_6423);
or U8327 (N_8327,N_7316,N_6163);
and U8328 (N_8328,N_6573,N_7786);
nor U8329 (N_8329,N_7757,N_7478);
nor U8330 (N_8330,N_6718,N_7310);
xnor U8331 (N_8331,N_7195,N_6891);
or U8332 (N_8332,N_7959,N_7449);
nand U8333 (N_8333,N_7045,N_6336);
xor U8334 (N_8334,N_6325,N_7061);
nand U8335 (N_8335,N_7454,N_7606);
or U8336 (N_8336,N_6396,N_7402);
nor U8337 (N_8337,N_7322,N_7718);
nor U8338 (N_8338,N_6736,N_6938);
xnor U8339 (N_8339,N_7486,N_6023);
or U8340 (N_8340,N_6498,N_6918);
nor U8341 (N_8341,N_7060,N_6772);
nor U8342 (N_8342,N_6899,N_7185);
nand U8343 (N_8343,N_6541,N_6665);
xor U8344 (N_8344,N_6768,N_7940);
or U8345 (N_8345,N_6991,N_6024);
or U8346 (N_8346,N_7541,N_7889);
nor U8347 (N_8347,N_6243,N_7243);
nand U8348 (N_8348,N_6574,N_7823);
nor U8349 (N_8349,N_6265,N_7355);
nand U8350 (N_8350,N_6455,N_6697);
and U8351 (N_8351,N_6954,N_7840);
and U8352 (N_8352,N_6105,N_7907);
xnor U8353 (N_8353,N_7348,N_7398);
nor U8354 (N_8354,N_7397,N_7431);
or U8355 (N_8355,N_7426,N_7344);
xor U8356 (N_8356,N_6183,N_6668);
xor U8357 (N_8357,N_7327,N_6417);
or U8358 (N_8358,N_6151,N_6099);
xnor U8359 (N_8359,N_7892,N_7916);
and U8360 (N_8360,N_7762,N_7372);
nor U8361 (N_8361,N_7696,N_6692);
nor U8362 (N_8362,N_6212,N_6196);
or U8363 (N_8363,N_6752,N_6071);
nand U8364 (N_8364,N_6198,N_6418);
and U8365 (N_8365,N_7530,N_7950);
xor U8366 (N_8366,N_6279,N_7488);
nand U8367 (N_8367,N_7511,N_7116);
xnor U8368 (N_8368,N_6091,N_6516);
and U8369 (N_8369,N_6276,N_6136);
and U8370 (N_8370,N_6457,N_7404);
nand U8371 (N_8371,N_7528,N_6597);
and U8372 (N_8372,N_6580,N_7607);
and U8373 (N_8373,N_6328,N_6615);
or U8374 (N_8374,N_6116,N_6069);
or U8375 (N_8375,N_6534,N_6579);
xnor U8376 (N_8376,N_7542,N_7014);
or U8377 (N_8377,N_6674,N_6114);
nor U8378 (N_8378,N_6386,N_7610);
and U8379 (N_8379,N_6705,N_7516);
xor U8380 (N_8380,N_6533,N_7746);
and U8381 (N_8381,N_6993,N_7731);
xnor U8382 (N_8382,N_6182,N_6405);
and U8383 (N_8383,N_6506,N_6011);
xor U8384 (N_8384,N_6203,N_7214);
and U8385 (N_8385,N_6786,N_6785);
or U8386 (N_8386,N_6395,N_6611);
nand U8387 (N_8387,N_7773,N_7334);
xor U8388 (N_8388,N_6802,N_6770);
nor U8389 (N_8389,N_7977,N_6963);
or U8390 (N_8390,N_6787,N_7356);
nor U8391 (N_8391,N_7505,N_7027);
nand U8392 (N_8392,N_6581,N_6756);
nor U8393 (N_8393,N_6412,N_7343);
nand U8394 (N_8394,N_6294,N_7970);
and U8395 (N_8395,N_7651,N_7952);
nor U8396 (N_8396,N_6543,N_6240);
and U8397 (N_8397,N_7933,N_7615);
nand U8398 (N_8398,N_6539,N_7250);
or U8399 (N_8399,N_7987,N_6659);
nor U8400 (N_8400,N_6738,N_7754);
or U8401 (N_8401,N_7672,N_7873);
and U8402 (N_8402,N_7856,N_7617);
nand U8403 (N_8403,N_7515,N_6741);
nand U8404 (N_8404,N_7366,N_7931);
nand U8405 (N_8405,N_6492,N_6332);
xor U8406 (N_8406,N_6758,N_7320);
nand U8407 (N_8407,N_6966,N_7602);
xor U8408 (N_8408,N_6609,N_7676);
xor U8409 (N_8409,N_7302,N_6222);
xnor U8410 (N_8410,N_6298,N_7406);
nand U8411 (N_8411,N_7359,N_7122);
and U8412 (N_8412,N_7139,N_7526);
nand U8413 (N_8413,N_7197,N_7015);
or U8414 (N_8414,N_7705,N_6984);
or U8415 (N_8415,N_6358,N_6465);
xor U8416 (N_8416,N_7604,N_7299);
nor U8417 (N_8417,N_6627,N_6292);
xnor U8418 (N_8418,N_6006,N_6865);
nor U8419 (N_8419,N_6592,N_7633);
xor U8420 (N_8420,N_7073,N_6757);
or U8421 (N_8421,N_6027,N_7103);
and U8422 (N_8422,N_6990,N_7474);
xor U8423 (N_8423,N_6497,N_6419);
and U8424 (N_8424,N_7373,N_7837);
nand U8425 (N_8425,N_6797,N_7246);
nand U8426 (N_8426,N_6924,N_7143);
or U8427 (N_8427,N_6823,N_6809);
and U8428 (N_8428,N_6249,N_6038);
and U8429 (N_8429,N_7543,N_7649);
or U8430 (N_8430,N_7326,N_7261);
or U8431 (N_8431,N_7416,N_7092);
and U8432 (N_8432,N_6125,N_7340);
xor U8433 (N_8433,N_7628,N_6040);
and U8434 (N_8434,N_7304,N_7062);
or U8435 (N_8435,N_7662,N_7679);
or U8436 (N_8436,N_7374,N_7905);
and U8437 (N_8437,N_6432,N_7774);
nand U8438 (N_8438,N_6557,N_7796);
xor U8439 (N_8439,N_7314,N_6124);
xnor U8440 (N_8440,N_7595,N_7154);
nand U8441 (N_8441,N_6141,N_6032);
nor U8442 (N_8442,N_7621,N_7232);
nor U8443 (N_8443,N_6185,N_7200);
or U8444 (N_8444,N_6398,N_6715);
nor U8445 (N_8445,N_7086,N_6562);
xnor U8446 (N_8446,N_7187,N_7759);
nor U8447 (N_8447,N_6199,N_6817);
xnor U8448 (N_8448,N_7168,N_6029);
nor U8449 (N_8449,N_7618,N_7003);
and U8450 (N_8450,N_6774,N_6538);
nor U8451 (N_8451,N_7134,N_6805);
nand U8452 (N_8452,N_7052,N_6140);
or U8453 (N_8453,N_7652,N_7634);
and U8454 (N_8454,N_7102,N_7567);
and U8455 (N_8455,N_6870,N_7730);
nand U8456 (N_8456,N_6798,N_6462);
nand U8457 (N_8457,N_7041,N_7727);
and U8458 (N_8458,N_6037,N_6678);
nand U8459 (N_8459,N_6632,N_6098);
xor U8460 (N_8460,N_7367,N_6411);
nand U8461 (N_8461,N_7274,N_7255);
nand U8462 (N_8462,N_7858,N_7442);
xnor U8463 (N_8463,N_6437,N_6980);
xnor U8464 (N_8464,N_6383,N_7050);
xor U8465 (N_8465,N_6630,N_6049);
and U8466 (N_8466,N_6568,N_6834);
xnor U8467 (N_8467,N_7763,N_7654);
or U8468 (N_8468,N_7172,N_7018);
nand U8469 (N_8469,N_6633,N_6646);
xor U8470 (N_8470,N_6111,N_6441);
and U8471 (N_8471,N_7100,N_6994);
nand U8472 (N_8472,N_7766,N_6489);
and U8473 (N_8473,N_6372,N_6832);
and U8474 (N_8474,N_7996,N_7583);
nor U8475 (N_8475,N_7934,N_7191);
nand U8476 (N_8476,N_6794,N_6430);
xor U8477 (N_8477,N_7835,N_7884);
xnor U8478 (N_8478,N_6169,N_6192);
nand U8479 (N_8479,N_6215,N_7377);
xor U8480 (N_8480,N_7640,N_7150);
nand U8481 (N_8481,N_6729,N_7924);
and U8482 (N_8482,N_6464,N_6435);
and U8483 (N_8483,N_7368,N_7112);
and U8484 (N_8484,N_6610,N_6471);
xor U8485 (N_8485,N_7059,N_6998);
nand U8486 (N_8486,N_7199,N_6227);
and U8487 (N_8487,N_6436,N_7140);
nor U8488 (N_8488,N_6054,N_6434);
or U8489 (N_8489,N_7601,N_6184);
nor U8490 (N_8490,N_6601,N_7354);
xnor U8491 (N_8491,N_7956,N_7850);
nor U8492 (N_8492,N_7594,N_7462);
or U8493 (N_8493,N_6733,N_7863);
xor U8494 (N_8494,N_7580,N_6840);
nand U8495 (N_8495,N_7138,N_7105);
and U8496 (N_8496,N_7228,N_6500);
or U8497 (N_8497,N_6387,N_7341);
xnor U8498 (N_8498,N_6220,N_7955);
and U8499 (N_8499,N_6178,N_6936);
xor U8500 (N_8500,N_7297,N_7501);
or U8501 (N_8501,N_7918,N_6073);
nand U8502 (N_8502,N_6177,N_6468);
nand U8503 (N_8503,N_6828,N_7720);
xor U8504 (N_8504,N_6997,N_7953);
nor U8505 (N_8505,N_6080,N_6743);
xnor U8506 (N_8506,N_6062,N_7980);
or U8507 (N_8507,N_7577,N_6337);
and U8508 (N_8508,N_6014,N_6686);
and U8509 (N_8509,N_7725,N_7571);
and U8510 (N_8510,N_7810,N_6404);
nand U8511 (N_8511,N_7075,N_6585);
nor U8512 (N_8512,N_6253,N_7209);
nor U8513 (N_8513,N_7234,N_6945);
xnor U8514 (N_8514,N_7038,N_6139);
xor U8515 (N_8515,N_7147,N_6937);
and U8516 (N_8516,N_6267,N_6783);
nand U8517 (N_8517,N_6960,N_7434);
and U8518 (N_8518,N_6979,N_6546);
or U8519 (N_8519,N_6162,N_6663);
nand U8520 (N_8520,N_6217,N_6313);
or U8521 (N_8521,N_6713,N_6903);
nor U8522 (N_8522,N_7960,N_6883);
or U8523 (N_8523,N_6264,N_7016);
nor U8524 (N_8524,N_6005,N_6406);
xnor U8525 (N_8525,N_7155,N_6045);
xnor U8526 (N_8526,N_7271,N_7411);
or U8527 (N_8527,N_7445,N_6154);
or U8528 (N_8528,N_7958,N_6717);
nand U8529 (N_8529,N_7084,N_6120);
or U8530 (N_8530,N_7464,N_7123);
nand U8531 (N_8531,N_7459,N_7521);
nand U8532 (N_8532,N_6553,N_7721);
nor U8533 (N_8533,N_6085,N_7947);
and U8534 (N_8534,N_6157,N_7548);
or U8535 (N_8535,N_7125,N_6857);
and U8536 (N_8536,N_6843,N_6569);
and U8537 (N_8537,N_7954,N_7733);
nor U8538 (N_8538,N_7636,N_6652);
or U8539 (N_8539,N_6044,N_6376);
nand U8540 (N_8540,N_7201,N_6360);
nor U8541 (N_8541,N_6416,N_7451);
xor U8542 (N_8542,N_6020,N_6013);
xnor U8543 (N_8543,N_7664,N_7282);
nand U8544 (N_8544,N_7709,N_6709);
and U8545 (N_8545,N_7268,N_7407);
nand U8546 (N_8546,N_7363,N_7818);
and U8547 (N_8547,N_7470,N_7496);
nor U8548 (N_8548,N_7917,N_6176);
xor U8549 (N_8549,N_7962,N_7808);
nor U8550 (N_8550,N_6363,N_6622);
xor U8551 (N_8551,N_7207,N_6101);
and U8552 (N_8552,N_6987,N_6619);
xnor U8553 (N_8553,N_6424,N_7930);
xor U8554 (N_8554,N_7293,N_7176);
and U8555 (N_8555,N_7128,N_7113);
nand U8556 (N_8556,N_6650,N_7843);
xnor U8557 (N_8557,N_7663,N_6819);
or U8558 (N_8558,N_7000,N_6689);
and U8559 (N_8559,N_7177,N_7342);
or U8560 (N_8560,N_6570,N_6532);
or U8561 (N_8561,N_6842,N_7133);
xor U8562 (N_8562,N_7395,N_7512);
or U8563 (N_8563,N_6340,N_7163);
or U8564 (N_8564,N_6263,N_6446);
nand U8565 (N_8565,N_7896,N_7068);
nor U8566 (N_8566,N_6160,N_7854);
and U8567 (N_8567,N_6810,N_6368);
xor U8568 (N_8568,N_7428,N_6942);
nor U8569 (N_8569,N_7258,N_6866);
nor U8570 (N_8570,N_7455,N_7899);
and U8571 (N_8571,N_6958,N_7547);
or U8572 (N_8572,N_6795,N_7365);
and U8573 (N_8573,N_6732,N_7836);
and U8574 (N_8574,N_7665,N_7025);
xnor U8575 (N_8575,N_6951,N_7224);
nor U8576 (N_8576,N_7817,N_7545);
and U8577 (N_8577,N_7544,N_7625);
and U8578 (N_8578,N_6296,N_6479);
nand U8579 (N_8579,N_6596,N_7323);
xnor U8580 (N_8580,N_6559,N_7171);
xnor U8581 (N_8581,N_7717,N_6651);
nor U8582 (N_8582,N_7239,N_7780);
and U8583 (N_8583,N_6246,N_6259);
nand U8584 (N_8584,N_6127,N_6090);
xnor U8585 (N_8585,N_7233,N_6511);
nor U8586 (N_8586,N_6526,N_7135);
xor U8587 (N_8587,N_7842,N_7205);
xor U8588 (N_8588,N_6522,N_6587);
xor U8589 (N_8589,N_7513,N_6041);
or U8590 (N_8590,N_6548,N_7985);
nand U8591 (N_8591,N_6129,N_6837);
nor U8592 (N_8592,N_6694,N_7120);
nor U8593 (N_8593,N_6603,N_7540);
or U8594 (N_8594,N_6087,N_7722);
and U8595 (N_8595,N_7378,N_7972);
and U8596 (N_8596,N_7573,N_6839);
or U8597 (N_8597,N_6989,N_7847);
or U8598 (N_8598,N_7256,N_6706);
nand U8599 (N_8599,N_6366,N_6231);
nand U8600 (N_8600,N_7085,N_7495);
nor U8601 (N_8601,N_6662,N_7409);
nor U8602 (N_8602,N_7487,N_7032);
xnor U8603 (N_8603,N_7869,N_7399);
nand U8604 (N_8604,N_6107,N_7328);
xor U8605 (N_8605,N_6156,N_7419);
xnor U8606 (N_8606,N_6950,N_7939);
nor U8607 (N_8607,N_7098,N_6560);
nor U8608 (N_8608,N_6949,N_7643);
xor U8609 (N_8609,N_7048,N_6521);
nor U8610 (N_8610,N_6996,N_7745);
xor U8611 (N_8611,N_6118,N_6057);
nor U8612 (N_8612,N_7083,N_6365);
and U8613 (N_8613,N_6930,N_7375);
xor U8614 (N_8614,N_7797,N_6459);
xor U8615 (N_8615,N_6273,N_6371);
nor U8616 (N_8616,N_7037,N_6563);
nand U8617 (N_8617,N_7670,N_7216);
and U8618 (N_8618,N_7219,N_6234);
and U8619 (N_8619,N_6097,N_6735);
nor U8620 (N_8620,N_6916,N_6347);
nand U8621 (N_8621,N_7639,N_7456);
or U8622 (N_8622,N_7269,N_6685);
nand U8623 (N_8623,N_7656,N_7657);
nor U8624 (N_8624,N_7311,N_6349);
or U8625 (N_8625,N_6458,N_7868);
or U8626 (N_8626,N_6595,N_6326);
nor U8627 (N_8627,N_7076,N_6344);
nand U8628 (N_8628,N_7017,N_7440);
and U8629 (N_8629,N_6306,N_7761);
xor U8630 (N_8630,N_6629,N_6056);
nor U8631 (N_8631,N_6343,N_6362);
or U8632 (N_8632,N_6274,N_6308);
and U8633 (N_8633,N_7285,N_6645);
and U8634 (N_8634,N_7508,N_7198);
or U8635 (N_8635,N_7598,N_7063);
xnor U8636 (N_8636,N_7608,N_7007);
nand U8637 (N_8637,N_6288,N_7853);
nand U8638 (N_8638,N_6790,N_7518);
and U8639 (N_8639,N_6018,N_7031);
nand U8640 (N_8640,N_7978,N_6271);
or U8641 (N_8641,N_6373,N_7740);
or U8642 (N_8642,N_6171,N_7900);
xor U8643 (N_8643,N_6147,N_7353);
or U8644 (N_8644,N_6143,N_6803);
and U8645 (N_8645,N_7747,N_7335);
and U8646 (N_8646,N_7728,N_7992);
nand U8647 (N_8647,N_6043,N_6520);
nand U8648 (N_8648,N_6260,N_6975);
xor U8649 (N_8649,N_7101,N_7546);
nand U8650 (N_8650,N_7920,N_7989);
nand U8651 (N_8651,N_7131,N_7447);
nand U8652 (N_8652,N_7370,N_6616);
xor U8653 (N_8653,N_7912,N_6917);
and U8654 (N_8654,N_6224,N_7151);
and U8655 (N_8655,N_6300,N_7829);
or U8656 (N_8656,N_6905,N_7309);
nor U8657 (N_8657,N_7812,N_7351);
nand U8658 (N_8658,N_6571,N_7159);
nand U8659 (N_8659,N_6856,N_6467);
nor U8660 (N_8660,N_7337,N_7051);
nor U8661 (N_8661,N_7789,N_7795);
nor U8662 (N_8662,N_7815,N_6564);
nand U8663 (N_8663,N_6598,N_6542);
or U8664 (N_8664,N_6126,N_6518);
nor U8665 (N_8665,N_7066,N_7841);
and U8666 (N_8666,N_6158,N_6614);
xnor U8667 (N_8667,N_7263,N_6524);
nor U8668 (N_8668,N_7865,N_6888);
or U8669 (N_8669,N_7306,N_6625);
and U8670 (N_8670,N_6012,N_7259);
nand U8671 (N_8671,N_6252,N_7668);
xnor U8672 (N_8672,N_6193,N_6600);
xnor U8673 (N_8673,N_6982,N_6875);
or U8674 (N_8674,N_6478,N_7288);
or U8675 (N_8675,N_6556,N_6115);
xnor U8676 (N_8676,N_7091,N_6010);
nor U8677 (N_8677,N_6302,N_6961);
nand U8678 (N_8678,N_7192,N_7715);
nand U8679 (N_8679,N_7592,N_6724);
and U8680 (N_8680,N_6864,N_7908);
nor U8681 (N_8681,N_7915,N_7527);
nand U8682 (N_8682,N_7964,N_7788);
nand U8683 (N_8683,N_6695,N_7862);
nor U8684 (N_8684,N_6816,N_7333);
or U8685 (N_8685,N_7799,N_7183);
nor U8686 (N_8686,N_7109,N_7276);
or U8687 (N_8687,N_7286,N_7734);
or U8688 (N_8688,N_6721,N_6004);
and U8689 (N_8689,N_7034,N_7574);
nand U8690 (N_8690,N_7979,N_6469);
and U8691 (N_8691,N_6451,N_6237);
xor U8692 (N_8692,N_6637,N_6166);
and U8693 (N_8693,N_6281,N_6112);
xor U8694 (N_8694,N_7422,N_7030);
or U8695 (N_8695,N_7039,N_7556);
xor U8696 (N_8696,N_6095,N_6762);
or U8697 (N_8697,N_6826,N_7452);
nand U8698 (N_8698,N_7132,N_7313);
nor U8699 (N_8699,N_6320,N_7800);
and U8700 (N_8700,N_6767,N_7570);
xor U8701 (N_8701,N_6216,N_7775);
nand U8702 (N_8702,N_7779,N_7737);
and U8703 (N_8703,N_6047,N_6764);
or U8704 (N_8704,N_7443,N_6861);
xor U8705 (N_8705,N_6351,N_7371);
xor U8706 (N_8706,N_7106,N_6361);
nand U8707 (N_8707,N_6527,N_7010);
nor U8708 (N_8708,N_6508,N_7493);
nor U8709 (N_8709,N_6341,N_7088);
and U8710 (N_8710,N_6977,N_6988);
or U8711 (N_8711,N_6545,N_7064);
or U8712 (N_8712,N_6893,N_6493);
nand U8713 (N_8713,N_6311,N_7948);
nand U8714 (N_8714,N_6256,N_6223);
nor U8715 (N_8715,N_6438,N_7461);
or U8716 (N_8716,N_6359,N_6887);
or U8717 (N_8717,N_7227,N_6104);
nor U8718 (N_8718,N_7880,N_6890);
xor U8719 (N_8719,N_7881,N_6932);
or U8720 (N_8720,N_7951,N_7148);
nor U8721 (N_8721,N_6859,N_6319);
or U8722 (N_8722,N_6391,N_7736);
or U8723 (N_8723,N_7042,N_6710);
nand U8724 (N_8724,N_6913,N_6312);
nor U8725 (N_8725,N_6853,N_6470);
or U8726 (N_8726,N_6053,N_7145);
xnor U8727 (N_8727,N_6463,N_6210);
or U8728 (N_8728,N_6346,N_6036);
xor U8729 (N_8729,N_7949,N_7514);
nand U8730 (N_8730,N_6976,N_7578);
xnor U8731 (N_8731,N_6408,N_7599);
or U8732 (N_8732,N_6048,N_6910);
and U8733 (N_8733,N_6204,N_7160);
xor U8734 (N_8734,N_6035,N_6824);
nor U8735 (N_8735,N_7561,N_6280);
or U8736 (N_8736,N_6026,N_7126);
nand U8737 (N_8737,N_7127,N_7388);
and U8738 (N_8738,N_7494,N_7687);
nand U8739 (N_8739,N_6081,N_7362);
xnor U8740 (N_8740,N_7826,N_7965);
xor U8741 (N_8741,N_7609,N_6830);
and U8742 (N_8742,N_6959,N_7247);
nor U8743 (N_8743,N_6061,N_6079);
or U8744 (N_8744,N_6232,N_7968);
xor U8745 (N_8745,N_7596,N_7047);
and U8746 (N_8746,N_6208,N_6149);
nand U8747 (N_8747,N_7586,N_7206);
or U8748 (N_8748,N_7680,N_7040);
xnor U8749 (N_8749,N_7339,N_7925);
and U8750 (N_8750,N_7520,N_6698);
xnor U8751 (N_8751,N_7415,N_6700);
xor U8752 (N_8752,N_6286,N_7926);
and U8753 (N_8753,N_7785,N_7997);
xnor U8754 (N_8754,N_6789,N_7929);
or U8755 (N_8755,N_6552,N_6254);
and U8756 (N_8756,N_6894,N_6379);
and U8757 (N_8757,N_7982,N_7053);
or U8758 (N_8758,N_6307,N_6666);
or U8759 (N_8759,N_6778,N_6188);
xnor U8760 (N_8760,N_7945,N_7614);
or U8761 (N_8761,N_6088,N_7221);
or U8762 (N_8762,N_7635,N_6046);
nand U8763 (N_8763,N_7559,N_6186);
xnor U8764 (N_8764,N_7330,N_6352);
nor U8765 (N_8765,N_7315,N_6482);
nand U8766 (N_8766,N_6881,N_7036);
nor U8767 (N_8767,N_7724,N_7225);
nor U8768 (N_8768,N_7660,N_6577);
and U8769 (N_8769,N_6884,N_7142);
or U8770 (N_8770,N_6631,N_6696);
or U8771 (N_8771,N_7821,N_7065);
xor U8772 (N_8772,N_7619,N_7726);
nand U8773 (N_8773,N_7457,N_7162);
xor U8774 (N_8774,N_7510,N_7707);
and U8775 (N_8775,N_7692,N_6397);
nor U8776 (N_8776,N_7024,N_7993);
or U8777 (N_8777,N_7006,N_7196);
xor U8778 (N_8778,N_6218,N_7612);
nand U8779 (N_8779,N_7173,N_6879);
and U8780 (N_8780,N_6121,N_7079);
nor U8781 (N_8781,N_6174,N_6730);
nor U8782 (N_8782,N_7533,N_7408);
or U8783 (N_8783,N_6897,N_7423);
nor U8784 (N_8784,N_7471,N_6277);
and U8785 (N_8785,N_7781,N_6503);
nor U8786 (N_8786,N_6290,N_7476);
or U8787 (N_8787,N_7957,N_6978);
nor U8788 (N_8788,N_7932,N_7361);
nand U8789 (N_8789,N_6711,N_7175);
or U8790 (N_8790,N_6399,N_7532);
nand U8791 (N_8791,N_7137,N_6094);
nor U8792 (N_8792,N_6019,N_7331);
or U8793 (N_8793,N_7691,N_6868);
xor U8794 (N_8794,N_7703,N_7739);
xor U8795 (N_8795,N_6067,N_7158);
xnor U8796 (N_8796,N_6957,N_7772);
nand U8797 (N_8797,N_6590,N_6122);
xnor U8798 (N_8798,N_7913,N_7281);
xnor U8799 (N_8799,N_7435,N_6285);
or U8800 (N_8800,N_7110,N_6484);
nor U8801 (N_8801,N_6030,N_6187);
nor U8802 (N_8802,N_6034,N_7450);
and U8803 (N_8803,N_6331,N_7816);
or U8804 (N_8804,N_7129,N_6687);
or U8805 (N_8805,N_7729,N_6384);
nor U8806 (N_8806,N_6241,N_7701);
xnor U8807 (N_8807,N_7240,N_6670);
xnor U8808 (N_8808,N_6947,N_7697);
xnor U8809 (N_8809,N_6535,N_6009);
nor U8810 (N_8810,N_7485,N_7814);
or U8811 (N_8811,N_6219,N_7500);
nor U8812 (N_8812,N_6485,N_7170);
and U8813 (N_8813,N_7270,N_6339);
or U8814 (N_8814,N_7922,N_7832);
and U8815 (N_8815,N_7603,N_7861);
xnor U8816 (N_8816,N_7871,N_6392);
or U8817 (N_8817,N_6357,N_7894);
or U8818 (N_8818,N_7706,N_6551);
and U8819 (N_8819,N_6940,N_6777);
and U8820 (N_8820,N_7389,N_7182);
nand U8821 (N_8821,N_6304,N_6134);
nand U8822 (N_8822,N_6639,N_7121);
nor U8823 (N_8823,N_6180,N_7683);
nor U8824 (N_8824,N_7161,N_6473);
xor U8825 (N_8825,N_6867,N_6148);
nor U8826 (N_8826,N_7498,N_7300);
nor U8827 (N_8827,N_6031,N_6846);
nor U8828 (N_8828,N_6836,N_7735);
xor U8829 (N_8829,N_7552,N_6878);
nand U8830 (N_8830,N_6793,N_7647);
xor U8831 (N_8831,N_6450,N_7184);
and U8832 (N_8832,N_6657,N_7480);
nor U8833 (N_8833,N_6519,N_6607);
or U8834 (N_8834,N_6329,N_6964);
and U8835 (N_8835,N_7283,N_6877);
and U8836 (N_8836,N_6262,N_7998);
nor U8837 (N_8837,N_6636,N_7394);
or U8838 (N_8838,N_7096,N_7427);
and U8839 (N_8839,N_7287,N_7879);
or U8840 (N_8840,N_6003,N_7831);
nand U8841 (N_8841,N_6872,N_7400);
and U8842 (N_8842,N_6647,N_7787);
nor U8843 (N_8843,N_6791,N_7524);
nor U8844 (N_8844,N_7597,N_7666);
or U8845 (N_8845,N_7229,N_7067);
nand U8846 (N_8846,N_7481,N_7376);
nor U8847 (N_8847,N_7844,N_6644);
and U8848 (N_8848,N_7582,N_6189);
nand U8849 (N_8849,N_7902,N_6350);
and U8850 (N_8850,N_7791,N_6766);
and U8851 (N_8851,N_6578,N_6480);
nor U8852 (N_8852,N_6420,N_6375);
and U8853 (N_8853,N_7898,N_7529);
and U8854 (N_8854,N_7174,N_6554);
and U8855 (N_8855,N_7671,N_6051);
or U8856 (N_8856,N_7217,N_7403);
or U8857 (N_8857,N_6995,N_7022);
or U8858 (N_8858,N_7756,N_6845);
or U8859 (N_8859,N_7043,N_6567);
or U8860 (N_8860,N_7460,N_6848);
nand U8861 (N_8861,N_6239,N_6621);
and U8862 (N_8862,N_6168,N_7244);
nor U8863 (N_8863,N_6904,N_6213);
or U8864 (N_8864,N_6558,N_7294);
or U8865 (N_8865,N_6973,N_6926);
and U8866 (N_8866,N_6440,N_6173);
xnor U8867 (N_8867,N_6514,N_6565);
or U8868 (N_8868,N_7760,N_6602);
nand U8869 (N_8869,N_6649,N_6472);
or U8870 (N_8870,N_6078,N_6353);
nand U8871 (N_8871,N_7054,N_7535);
and U8872 (N_8872,N_6860,N_6461);
nand U8873 (N_8873,N_7976,N_7178);
or U8874 (N_8874,N_7329,N_7937);
nor U8875 (N_8875,N_6935,N_7776);
nor U8876 (N_8876,N_7417,N_7702);
or U8877 (N_8877,N_6269,N_6229);
nand U8878 (N_8878,N_7981,N_7507);
nand U8879 (N_8879,N_7822,N_6672);
nor U8880 (N_8880,N_6780,N_6744);
xor U8881 (N_8881,N_7210,N_7742);
xnor U8882 (N_8882,N_7253,N_6544);
or U8883 (N_8883,N_6150,N_7562);
nand U8884 (N_8884,N_7492,N_6576);
nor U8885 (N_8885,N_6483,N_7685);
xor U8886 (N_8886,N_6801,N_6796);
or U8887 (N_8887,N_6334,N_6701);
and U8888 (N_8888,N_6499,N_6060);
xor U8889 (N_8889,N_7804,N_7743);
nor U8890 (N_8890,N_7627,N_6941);
nand U8891 (N_8891,N_6261,N_6015);
and U8892 (N_8892,N_7165,N_6820);
nand U8893 (N_8893,N_7563,N_7439);
nor U8894 (N_8894,N_6236,N_6683);
nand U8895 (N_8895,N_7566,N_6209);
or U8896 (N_8896,N_6191,N_6968);
xnor U8897 (N_8897,N_7644,N_6063);
nor U8898 (N_8898,N_6771,N_6953);
xnor U8899 (N_8899,N_6776,N_6370);
nand U8900 (N_8900,N_7753,N_7009);
nand U8901 (N_8901,N_7961,N_7369);
and U8902 (N_8902,N_6841,N_7771);
and U8903 (N_8903,N_7272,N_7265);
or U8904 (N_8904,N_6345,N_6102);
and U8905 (N_8905,N_7124,N_7557);
xor U8906 (N_8906,N_6394,N_6703);
and U8907 (N_8907,N_7975,N_6765);
nor U8908 (N_8908,N_7585,N_6400);
and U8909 (N_8909,N_7468,N_7646);
nor U8910 (N_8910,N_6103,N_6335);
nor U8911 (N_8911,N_6318,N_6628);
nor U8912 (N_8912,N_6754,N_6981);
or U8913 (N_8913,N_7252,N_6708);
nor U8914 (N_8914,N_7466,N_7860);
or U8915 (N_8915,N_6257,N_6555);
xor U8916 (N_8916,N_7506,N_7312);
or U8917 (N_8917,N_6128,N_7744);
or U8918 (N_8918,N_7517,N_7503);
and U8919 (N_8919,N_7390,N_7994);
or U8920 (N_8920,N_6838,N_6159);
xor U8921 (N_8921,N_6167,N_6117);
and U8922 (N_8922,N_6272,N_7767);
and U8923 (N_8923,N_6792,N_7425);
and U8924 (N_8924,N_7675,N_6550);
nor U8925 (N_8925,N_7723,N_6985);
nor U8926 (N_8926,N_6986,N_7813);
nor U8927 (N_8927,N_7537,N_7349);
and U8928 (N_8928,N_7118,N_7576);
nor U8929 (N_8929,N_6871,N_6927);
or U8930 (N_8930,N_7629,N_6742);
nand U8931 (N_8931,N_6779,N_6305);
xor U8932 (N_8932,N_6726,N_6211);
nor U8933 (N_8933,N_6248,N_6113);
nor U8934 (N_8934,N_7897,N_7074);
nor U8935 (N_8935,N_7587,N_7650);
and U8936 (N_8936,N_7872,N_6266);
xnor U8937 (N_8937,N_6620,N_7560);
or U8938 (N_8938,N_6992,N_6784);
nor U8939 (N_8939,N_7928,N_6800);
nand U8940 (N_8940,N_6909,N_7988);
and U8941 (N_8941,N_6970,N_7292);
nand U8942 (N_8942,N_6444,N_6324);
nand U8943 (N_8943,N_7305,N_6642);
or U8944 (N_8944,N_6589,N_6123);
nand U8945 (N_8945,N_6445,N_6414);
nor U8946 (N_8946,N_7875,N_6247);
nand U8947 (N_8947,N_6720,N_7611);
nand U8948 (N_8948,N_6025,N_7575);
xnor U8949 (N_8949,N_6759,N_6886);
nand U8950 (N_8950,N_6876,N_6374);
nand U8951 (N_8951,N_6679,N_6594);
xor U8952 (N_8952,N_6528,N_6317);
nor U8953 (N_8953,N_7613,N_7699);
and U8954 (N_8954,N_7336,N_6923);
and U8955 (N_8955,N_7069,N_6648);
and U8956 (N_8956,N_6316,N_7674);
or U8957 (N_8957,N_6225,N_7115);
and U8958 (N_8958,N_6745,N_6207);
or U8959 (N_8959,N_7308,N_7765);
xor U8960 (N_8960,N_6323,N_6481);
nand U8961 (N_8961,N_7782,N_6928);
or U8962 (N_8962,N_6931,N_6747);
xor U8963 (N_8963,N_6664,N_7169);
nor U8964 (N_8964,N_6108,N_7019);
xor U8965 (N_8965,N_6885,N_6833);
or U8966 (N_8966,N_7909,N_6052);
nand U8967 (N_8967,N_6561,N_6238);
xnor U8968 (N_8968,N_6367,N_7338);
xor U8969 (N_8969,N_7632,N_7446);
nand U8970 (N_8970,N_6847,N_6523);
or U8971 (N_8971,N_7911,N_7490);
nand U8972 (N_8972,N_7923,N_7673);
nor U8973 (N_8973,N_7001,N_7057);
nor U8974 (N_8974,N_7748,N_7828);
or U8975 (N_8975,N_6161,N_7146);
nand U8976 (N_8976,N_7011,N_7296);
nand U8977 (N_8977,N_6165,N_6739);
nor U8978 (N_8978,N_7538,N_7758);
nor U8979 (N_8979,N_7497,N_7752);
xnor U8980 (N_8980,N_6245,N_7413);
xnor U8981 (N_8981,N_6755,N_7136);
nand U8982 (N_8982,N_7301,N_6505);
xnor U8983 (N_8983,N_6017,N_7241);
nand U8984 (N_8984,N_6190,N_7033);
nor U8985 (N_8985,N_6083,N_6851);
nor U8986 (N_8986,N_7049,N_7046);
nor U8987 (N_8987,N_7078,N_7811);
xor U8988 (N_8988,N_6301,N_6722);
nand U8989 (N_8989,N_7927,N_6131);
and U8990 (N_8990,N_7867,N_7565);
xor U8991 (N_8991,N_7157,N_6378);
or U8992 (N_8992,N_6299,N_7289);
nor U8993 (N_8993,N_6076,N_6688);
nand U8994 (N_8994,N_6001,N_7005);
nor U8995 (N_8995,N_6488,N_7350);
xnor U8996 (N_8996,N_7318,N_6529);
nor U8997 (N_8997,N_6486,N_6831);
or U8998 (N_8998,N_7589,N_7886);
and U8999 (N_8999,N_7215,N_6401);
and U9000 (N_9000,N_7404,N_7369);
or U9001 (N_9001,N_7441,N_6735);
or U9002 (N_9002,N_7247,N_7677);
xor U9003 (N_9003,N_7532,N_6981);
xnor U9004 (N_9004,N_7777,N_7624);
and U9005 (N_9005,N_6728,N_6465);
xnor U9006 (N_9006,N_6587,N_7163);
xnor U9007 (N_9007,N_6149,N_7453);
nor U9008 (N_9008,N_6867,N_6060);
or U9009 (N_9009,N_7381,N_7936);
and U9010 (N_9010,N_7799,N_7662);
nor U9011 (N_9011,N_6600,N_7446);
xor U9012 (N_9012,N_7219,N_6620);
or U9013 (N_9013,N_7699,N_6554);
nand U9014 (N_9014,N_7227,N_6597);
or U9015 (N_9015,N_7175,N_6762);
xnor U9016 (N_9016,N_6606,N_6996);
xor U9017 (N_9017,N_7283,N_7220);
or U9018 (N_9018,N_7078,N_6394);
or U9019 (N_9019,N_6543,N_7491);
or U9020 (N_9020,N_6002,N_7359);
or U9021 (N_9021,N_7969,N_7633);
nand U9022 (N_9022,N_6426,N_6342);
nor U9023 (N_9023,N_7486,N_6162);
and U9024 (N_9024,N_6423,N_7550);
and U9025 (N_9025,N_6447,N_7523);
or U9026 (N_9026,N_6453,N_6819);
and U9027 (N_9027,N_7368,N_7232);
xnor U9028 (N_9028,N_7378,N_6108);
and U9029 (N_9029,N_7635,N_7174);
and U9030 (N_9030,N_7177,N_6206);
nor U9031 (N_9031,N_7154,N_6078);
and U9032 (N_9032,N_6498,N_7916);
or U9033 (N_9033,N_7854,N_7413);
and U9034 (N_9034,N_7272,N_7873);
or U9035 (N_9035,N_7364,N_7826);
xor U9036 (N_9036,N_7395,N_6276);
nand U9037 (N_9037,N_6899,N_7748);
or U9038 (N_9038,N_7596,N_7070);
and U9039 (N_9039,N_6009,N_6436);
nand U9040 (N_9040,N_6989,N_6730);
or U9041 (N_9041,N_7607,N_6319);
or U9042 (N_9042,N_7914,N_6069);
nand U9043 (N_9043,N_7788,N_7960);
nor U9044 (N_9044,N_6058,N_6758);
or U9045 (N_9045,N_6616,N_7672);
nand U9046 (N_9046,N_6266,N_6317);
nor U9047 (N_9047,N_6396,N_6661);
or U9048 (N_9048,N_6987,N_7795);
or U9049 (N_9049,N_6201,N_6305);
or U9050 (N_9050,N_7604,N_6824);
nor U9051 (N_9051,N_7981,N_7653);
xor U9052 (N_9052,N_6913,N_6639);
xnor U9053 (N_9053,N_7753,N_6611);
nand U9054 (N_9054,N_6413,N_7766);
nand U9055 (N_9055,N_6025,N_6873);
xnor U9056 (N_9056,N_7325,N_7890);
or U9057 (N_9057,N_6599,N_7898);
or U9058 (N_9058,N_7803,N_7194);
nand U9059 (N_9059,N_6395,N_7652);
nor U9060 (N_9060,N_6300,N_6317);
nor U9061 (N_9061,N_6699,N_6478);
or U9062 (N_9062,N_6993,N_7966);
nand U9063 (N_9063,N_7694,N_6555);
xnor U9064 (N_9064,N_6996,N_6793);
xor U9065 (N_9065,N_7515,N_6349);
nand U9066 (N_9066,N_7633,N_6266);
nand U9067 (N_9067,N_7900,N_7920);
nand U9068 (N_9068,N_7869,N_6801);
nor U9069 (N_9069,N_7357,N_6592);
xnor U9070 (N_9070,N_6698,N_6022);
xnor U9071 (N_9071,N_7746,N_6207);
nand U9072 (N_9072,N_7951,N_6414);
or U9073 (N_9073,N_6936,N_7654);
and U9074 (N_9074,N_7915,N_7323);
and U9075 (N_9075,N_7293,N_7402);
xor U9076 (N_9076,N_7045,N_6716);
or U9077 (N_9077,N_7867,N_7208);
and U9078 (N_9078,N_7641,N_6061);
nor U9079 (N_9079,N_6001,N_7011);
nand U9080 (N_9080,N_6651,N_6700);
xnor U9081 (N_9081,N_7086,N_7545);
nor U9082 (N_9082,N_6512,N_7454);
or U9083 (N_9083,N_6429,N_6683);
nor U9084 (N_9084,N_7974,N_7539);
nor U9085 (N_9085,N_7361,N_6419);
and U9086 (N_9086,N_7150,N_6873);
nand U9087 (N_9087,N_7427,N_6352);
nor U9088 (N_9088,N_6561,N_7484);
or U9089 (N_9089,N_6426,N_7491);
xnor U9090 (N_9090,N_6372,N_6341);
or U9091 (N_9091,N_7158,N_7892);
nor U9092 (N_9092,N_6465,N_7977);
nor U9093 (N_9093,N_6549,N_7287);
or U9094 (N_9094,N_7105,N_6042);
xnor U9095 (N_9095,N_7059,N_6753);
nor U9096 (N_9096,N_7537,N_7485);
nand U9097 (N_9097,N_6705,N_7766);
nor U9098 (N_9098,N_7754,N_6478);
and U9099 (N_9099,N_6858,N_6182);
nand U9100 (N_9100,N_6299,N_7366);
nand U9101 (N_9101,N_7307,N_6416);
and U9102 (N_9102,N_7272,N_7793);
xor U9103 (N_9103,N_7482,N_6059);
nand U9104 (N_9104,N_7972,N_6545);
nor U9105 (N_9105,N_7427,N_7236);
nor U9106 (N_9106,N_7855,N_7158);
or U9107 (N_9107,N_7858,N_6673);
and U9108 (N_9108,N_7458,N_6164);
or U9109 (N_9109,N_7258,N_7558);
nand U9110 (N_9110,N_7093,N_7159);
nor U9111 (N_9111,N_7411,N_7942);
nor U9112 (N_9112,N_7554,N_6647);
and U9113 (N_9113,N_7408,N_6099);
xor U9114 (N_9114,N_6378,N_7717);
nand U9115 (N_9115,N_6151,N_7076);
xnor U9116 (N_9116,N_7960,N_7364);
xor U9117 (N_9117,N_6674,N_7924);
nor U9118 (N_9118,N_6140,N_6528);
nor U9119 (N_9119,N_6708,N_6180);
or U9120 (N_9120,N_7984,N_7533);
xor U9121 (N_9121,N_7329,N_6866);
xnor U9122 (N_9122,N_6750,N_6625);
nor U9123 (N_9123,N_6289,N_7748);
nand U9124 (N_9124,N_6919,N_7416);
and U9125 (N_9125,N_7566,N_6287);
xnor U9126 (N_9126,N_6292,N_6154);
and U9127 (N_9127,N_6168,N_6174);
xnor U9128 (N_9128,N_7267,N_6907);
and U9129 (N_9129,N_6256,N_6033);
xnor U9130 (N_9130,N_6568,N_6014);
xnor U9131 (N_9131,N_7251,N_6623);
xnor U9132 (N_9132,N_7313,N_6613);
xor U9133 (N_9133,N_7474,N_7165);
xor U9134 (N_9134,N_7899,N_7402);
and U9135 (N_9135,N_6514,N_7902);
or U9136 (N_9136,N_6374,N_6584);
xor U9137 (N_9137,N_6059,N_7869);
or U9138 (N_9138,N_7615,N_7519);
xnor U9139 (N_9139,N_6204,N_6899);
nor U9140 (N_9140,N_7929,N_6964);
nor U9141 (N_9141,N_6686,N_6870);
xnor U9142 (N_9142,N_6883,N_6630);
nand U9143 (N_9143,N_6674,N_7581);
and U9144 (N_9144,N_7975,N_6496);
nor U9145 (N_9145,N_6136,N_6368);
nor U9146 (N_9146,N_6000,N_6298);
and U9147 (N_9147,N_6327,N_6172);
or U9148 (N_9148,N_7236,N_6294);
nand U9149 (N_9149,N_7197,N_7334);
nand U9150 (N_9150,N_6410,N_7973);
xnor U9151 (N_9151,N_7281,N_7661);
nor U9152 (N_9152,N_7552,N_7698);
xor U9153 (N_9153,N_7457,N_7754);
and U9154 (N_9154,N_7893,N_6413);
or U9155 (N_9155,N_7452,N_7952);
nor U9156 (N_9156,N_6207,N_7266);
nor U9157 (N_9157,N_6966,N_6117);
nand U9158 (N_9158,N_6719,N_7119);
nor U9159 (N_9159,N_7439,N_6380);
or U9160 (N_9160,N_7129,N_7928);
or U9161 (N_9161,N_6170,N_7969);
xor U9162 (N_9162,N_6083,N_6442);
xor U9163 (N_9163,N_7239,N_6885);
and U9164 (N_9164,N_7637,N_7865);
or U9165 (N_9165,N_7850,N_6654);
or U9166 (N_9166,N_6904,N_7469);
nor U9167 (N_9167,N_7542,N_6187);
nor U9168 (N_9168,N_7288,N_7350);
and U9169 (N_9169,N_7593,N_6201);
and U9170 (N_9170,N_6132,N_6117);
xnor U9171 (N_9171,N_6675,N_6358);
nor U9172 (N_9172,N_7150,N_6489);
or U9173 (N_9173,N_7371,N_6922);
or U9174 (N_9174,N_6398,N_6245);
nand U9175 (N_9175,N_7613,N_7342);
nand U9176 (N_9176,N_6712,N_6542);
and U9177 (N_9177,N_7298,N_6884);
or U9178 (N_9178,N_7302,N_6269);
and U9179 (N_9179,N_6691,N_7321);
or U9180 (N_9180,N_6096,N_6666);
nand U9181 (N_9181,N_7580,N_6425);
or U9182 (N_9182,N_6685,N_7521);
xnor U9183 (N_9183,N_6230,N_7512);
nor U9184 (N_9184,N_7467,N_7441);
nor U9185 (N_9185,N_7968,N_7500);
nor U9186 (N_9186,N_7342,N_6946);
nand U9187 (N_9187,N_6783,N_7218);
nor U9188 (N_9188,N_7647,N_7936);
nor U9189 (N_9189,N_7090,N_6638);
xor U9190 (N_9190,N_7375,N_6645);
and U9191 (N_9191,N_6107,N_7607);
and U9192 (N_9192,N_6802,N_6886);
nor U9193 (N_9193,N_6798,N_7971);
xor U9194 (N_9194,N_6925,N_6051);
or U9195 (N_9195,N_6812,N_6505);
xor U9196 (N_9196,N_7498,N_6568);
nand U9197 (N_9197,N_6939,N_6027);
xnor U9198 (N_9198,N_6399,N_6103);
xor U9199 (N_9199,N_7296,N_6933);
nand U9200 (N_9200,N_7798,N_7918);
and U9201 (N_9201,N_6146,N_7323);
xor U9202 (N_9202,N_7047,N_6251);
and U9203 (N_9203,N_6650,N_7133);
or U9204 (N_9204,N_6313,N_6979);
xor U9205 (N_9205,N_7730,N_7275);
and U9206 (N_9206,N_7040,N_6353);
or U9207 (N_9207,N_7802,N_6456);
xor U9208 (N_9208,N_6880,N_7796);
or U9209 (N_9209,N_6557,N_6576);
xor U9210 (N_9210,N_6399,N_6681);
xnor U9211 (N_9211,N_6797,N_6012);
or U9212 (N_9212,N_7205,N_7194);
nor U9213 (N_9213,N_7811,N_7558);
and U9214 (N_9214,N_6624,N_7224);
or U9215 (N_9215,N_6827,N_6803);
xor U9216 (N_9216,N_6105,N_6119);
or U9217 (N_9217,N_6060,N_6805);
xor U9218 (N_9218,N_6539,N_7370);
or U9219 (N_9219,N_7076,N_6770);
and U9220 (N_9220,N_6852,N_6270);
xor U9221 (N_9221,N_6121,N_7628);
and U9222 (N_9222,N_7930,N_6902);
nor U9223 (N_9223,N_7200,N_7315);
or U9224 (N_9224,N_7988,N_6888);
and U9225 (N_9225,N_7592,N_7211);
nor U9226 (N_9226,N_6128,N_7202);
nand U9227 (N_9227,N_6563,N_6502);
or U9228 (N_9228,N_6890,N_6663);
nand U9229 (N_9229,N_6033,N_6159);
nor U9230 (N_9230,N_7406,N_6946);
and U9231 (N_9231,N_6062,N_6536);
and U9232 (N_9232,N_7563,N_7758);
nand U9233 (N_9233,N_6952,N_6793);
nand U9234 (N_9234,N_7242,N_6523);
or U9235 (N_9235,N_6481,N_6478);
and U9236 (N_9236,N_6749,N_7647);
nand U9237 (N_9237,N_7469,N_6999);
or U9238 (N_9238,N_7941,N_7918);
nor U9239 (N_9239,N_7848,N_7129);
nand U9240 (N_9240,N_6910,N_7768);
nand U9241 (N_9241,N_7522,N_7608);
or U9242 (N_9242,N_6035,N_7086);
and U9243 (N_9243,N_7345,N_6962);
nor U9244 (N_9244,N_7655,N_6135);
nor U9245 (N_9245,N_6931,N_6054);
and U9246 (N_9246,N_7424,N_7169);
nor U9247 (N_9247,N_6363,N_7375);
nand U9248 (N_9248,N_6651,N_7643);
or U9249 (N_9249,N_6474,N_6661);
or U9250 (N_9250,N_6680,N_6389);
and U9251 (N_9251,N_6207,N_7306);
xnor U9252 (N_9252,N_7274,N_6551);
and U9253 (N_9253,N_6629,N_7126);
nand U9254 (N_9254,N_6223,N_7881);
or U9255 (N_9255,N_7623,N_7265);
or U9256 (N_9256,N_7757,N_7509);
nand U9257 (N_9257,N_7286,N_7865);
nor U9258 (N_9258,N_7869,N_6096);
xor U9259 (N_9259,N_6245,N_7770);
nor U9260 (N_9260,N_6389,N_7886);
or U9261 (N_9261,N_7651,N_6684);
and U9262 (N_9262,N_7355,N_7477);
or U9263 (N_9263,N_7874,N_7931);
nor U9264 (N_9264,N_6366,N_7532);
nor U9265 (N_9265,N_7060,N_6222);
xor U9266 (N_9266,N_7226,N_7472);
nand U9267 (N_9267,N_6897,N_6178);
and U9268 (N_9268,N_6848,N_6683);
nand U9269 (N_9269,N_7312,N_6917);
or U9270 (N_9270,N_7184,N_6299);
and U9271 (N_9271,N_6955,N_6362);
and U9272 (N_9272,N_6371,N_7547);
nand U9273 (N_9273,N_7749,N_7326);
or U9274 (N_9274,N_7556,N_7074);
xnor U9275 (N_9275,N_6815,N_7086);
nor U9276 (N_9276,N_7139,N_6634);
or U9277 (N_9277,N_7201,N_7628);
and U9278 (N_9278,N_6085,N_6228);
nand U9279 (N_9279,N_6134,N_7991);
xor U9280 (N_9280,N_7375,N_6958);
nand U9281 (N_9281,N_6549,N_7929);
and U9282 (N_9282,N_7496,N_7512);
or U9283 (N_9283,N_6502,N_7250);
xnor U9284 (N_9284,N_6944,N_7017);
nor U9285 (N_9285,N_7055,N_7585);
nand U9286 (N_9286,N_6427,N_6733);
and U9287 (N_9287,N_6717,N_6788);
nand U9288 (N_9288,N_6222,N_6096);
xor U9289 (N_9289,N_7074,N_7767);
and U9290 (N_9290,N_6940,N_6918);
or U9291 (N_9291,N_7774,N_7380);
nor U9292 (N_9292,N_7404,N_6234);
or U9293 (N_9293,N_6233,N_6586);
nand U9294 (N_9294,N_6508,N_6444);
nand U9295 (N_9295,N_6950,N_7501);
or U9296 (N_9296,N_7916,N_7909);
nor U9297 (N_9297,N_7427,N_6372);
and U9298 (N_9298,N_7151,N_6445);
nor U9299 (N_9299,N_7074,N_7085);
xor U9300 (N_9300,N_6726,N_7900);
nand U9301 (N_9301,N_7648,N_6711);
xnor U9302 (N_9302,N_6668,N_6866);
nand U9303 (N_9303,N_6354,N_7624);
and U9304 (N_9304,N_7945,N_6182);
xor U9305 (N_9305,N_7323,N_7161);
nand U9306 (N_9306,N_6455,N_6849);
xor U9307 (N_9307,N_7870,N_6704);
nor U9308 (N_9308,N_7309,N_6390);
xor U9309 (N_9309,N_6770,N_6210);
nand U9310 (N_9310,N_6724,N_6395);
and U9311 (N_9311,N_7206,N_7868);
and U9312 (N_9312,N_7575,N_7364);
xnor U9313 (N_9313,N_7576,N_7638);
and U9314 (N_9314,N_6308,N_7357);
xor U9315 (N_9315,N_6767,N_6228);
or U9316 (N_9316,N_6045,N_7449);
nand U9317 (N_9317,N_6114,N_6659);
and U9318 (N_9318,N_7824,N_6315);
nor U9319 (N_9319,N_7037,N_6511);
or U9320 (N_9320,N_7439,N_7074);
xor U9321 (N_9321,N_6078,N_6349);
and U9322 (N_9322,N_6728,N_6055);
and U9323 (N_9323,N_7121,N_7374);
nor U9324 (N_9324,N_6078,N_6766);
nand U9325 (N_9325,N_6527,N_6670);
or U9326 (N_9326,N_6424,N_7850);
and U9327 (N_9327,N_6460,N_7585);
or U9328 (N_9328,N_6416,N_7655);
nand U9329 (N_9329,N_6444,N_7930);
or U9330 (N_9330,N_6692,N_7481);
nand U9331 (N_9331,N_6994,N_7249);
nor U9332 (N_9332,N_7502,N_7145);
and U9333 (N_9333,N_7072,N_6729);
nand U9334 (N_9334,N_6647,N_6382);
nor U9335 (N_9335,N_7466,N_6643);
xnor U9336 (N_9336,N_6010,N_6752);
nor U9337 (N_9337,N_7887,N_6564);
and U9338 (N_9338,N_7896,N_7902);
nand U9339 (N_9339,N_6549,N_6506);
nand U9340 (N_9340,N_6145,N_6712);
nand U9341 (N_9341,N_6451,N_7164);
nor U9342 (N_9342,N_6861,N_7112);
nand U9343 (N_9343,N_7184,N_7373);
or U9344 (N_9344,N_6399,N_6333);
xnor U9345 (N_9345,N_7533,N_7321);
xor U9346 (N_9346,N_7295,N_7575);
nand U9347 (N_9347,N_6350,N_7915);
nand U9348 (N_9348,N_7510,N_6069);
nor U9349 (N_9349,N_6541,N_7397);
nor U9350 (N_9350,N_7131,N_7730);
nor U9351 (N_9351,N_6626,N_7621);
and U9352 (N_9352,N_7460,N_6457);
nor U9353 (N_9353,N_6039,N_7442);
nand U9354 (N_9354,N_7620,N_7802);
or U9355 (N_9355,N_6733,N_7083);
xor U9356 (N_9356,N_7875,N_6896);
nor U9357 (N_9357,N_7234,N_6467);
and U9358 (N_9358,N_7500,N_7348);
xor U9359 (N_9359,N_6241,N_7909);
and U9360 (N_9360,N_7057,N_7820);
xnor U9361 (N_9361,N_7286,N_7233);
nor U9362 (N_9362,N_7098,N_6293);
and U9363 (N_9363,N_7226,N_7534);
nor U9364 (N_9364,N_7755,N_6232);
nor U9365 (N_9365,N_6887,N_7665);
xnor U9366 (N_9366,N_7903,N_6776);
xnor U9367 (N_9367,N_7149,N_7333);
or U9368 (N_9368,N_6772,N_6220);
nand U9369 (N_9369,N_6611,N_7472);
xnor U9370 (N_9370,N_7780,N_6092);
and U9371 (N_9371,N_7895,N_7095);
or U9372 (N_9372,N_6898,N_7768);
and U9373 (N_9373,N_6791,N_6904);
or U9374 (N_9374,N_7492,N_6327);
and U9375 (N_9375,N_6991,N_6862);
nor U9376 (N_9376,N_7686,N_7733);
nand U9377 (N_9377,N_7047,N_6234);
and U9378 (N_9378,N_7959,N_6240);
or U9379 (N_9379,N_6985,N_6137);
nand U9380 (N_9380,N_7206,N_6698);
nor U9381 (N_9381,N_6331,N_7963);
and U9382 (N_9382,N_7757,N_7181);
nand U9383 (N_9383,N_6661,N_7760);
nand U9384 (N_9384,N_7210,N_6832);
nor U9385 (N_9385,N_7393,N_7755);
and U9386 (N_9386,N_6066,N_6669);
xor U9387 (N_9387,N_6914,N_7907);
or U9388 (N_9388,N_6998,N_7156);
nand U9389 (N_9389,N_7724,N_7959);
or U9390 (N_9390,N_6186,N_7800);
or U9391 (N_9391,N_6272,N_7944);
xor U9392 (N_9392,N_6455,N_7131);
nor U9393 (N_9393,N_6299,N_7198);
nor U9394 (N_9394,N_7595,N_7354);
and U9395 (N_9395,N_7467,N_6057);
and U9396 (N_9396,N_7550,N_6781);
xor U9397 (N_9397,N_6010,N_7909);
or U9398 (N_9398,N_6931,N_6596);
nor U9399 (N_9399,N_6664,N_6755);
nand U9400 (N_9400,N_7825,N_7094);
and U9401 (N_9401,N_6185,N_7830);
and U9402 (N_9402,N_6630,N_6298);
and U9403 (N_9403,N_6798,N_6048);
or U9404 (N_9404,N_7849,N_7636);
and U9405 (N_9405,N_7338,N_7232);
xnor U9406 (N_9406,N_7528,N_6794);
nand U9407 (N_9407,N_6344,N_6773);
xnor U9408 (N_9408,N_7558,N_6185);
xor U9409 (N_9409,N_7108,N_7001);
nand U9410 (N_9410,N_7889,N_6498);
nor U9411 (N_9411,N_6915,N_7366);
and U9412 (N_9412,N_6453,N_7847);
and U9413 (N_9413,N_6869,N_6607);
or U9414 (N_9414,N_7727,N_6781);
nor U9415 (N_9415,N_7034,N_7520);
nor U9416 (N_9416,N_6333,N_7552);
nor U9417 (N_9417,N_6691,N_7603);
xor U9418 (N_9418,N_6585,N_6260);
xor U9419 (N_9419,N_6360,N_6916);
nor U9420 (N_9420,N_7009,N_7851);
nand U9421 (N_9421,N_7940,N_7256);
nand U9422 (N_9422,N_6036,N_6681);
or U9423 (N_9423,N_6745,N_7767);
or U9424 (N_9424,N_7031,N_7190);
nor U9425 (N_9425,N_6466,N_6075);
and U9426 (N_9426,N_7797,N_6060);
or U9427 (N_9427,N_6931,N_6004);
xor U9428 (N_9428,N_6572,N_7925);
or U9429 (N_9429,N_7918,N_7219);
nor U9430 (N_9430,N_7758,N_6912);
and U9431 (N_9431,N_7147,N_6103);
nor U9432 (N_9432,N_6343,N_6984);
or U9433 (N_9433,N_7641,N_7559);
or U9434 (N_9434,N_7905,N_6210);
nand U9435 (N_9435,N_7590,N_7647);
nand U9436 (N_9436,N_7012,N_6507);
xor U9437 (N_9437,N_7534,N_7565);
nand U9438 (N_9438,N_7585,N_7076);
nand U9439 (N_9439,N_7343,N_7856);
nand U9440 (N_9440,N_7473,N_7384);
xor U9441 (N_9441,N_7641,N_7464);
or U9442 (N_9442,N_6066,N_6477);
nor U9443 (N_9443,N_7498,N_6043);
nand U9444 (N_9444,N_6863,N_6720);
or U9445 (N_9445,N_6882,N_6618);
or U9446 (N_9446,N_6295,N_7639);
xor U9447 (N_9447,N_6311,N_7088);
nor U9448 (N_9448,N_6246,N_7425);
nand U9449 (N_9449,N_7193,N_7101);
and U9450 (N_9450,N_7512,N_6001);
or U9451 (N_9451,N_7590,N_6987);
nand U9452 (N_9452,N_6656,N_6307);
and U9453 (N_9453,N_7183,N_6059);
nand U9454 (N_9454,N_6469,N_6986);
xnor U9455 (N_9455,N_7822,N_7889);
xor U9456 (N_9456,N_7997,N_7299);
or U9457 (N_9457,N_6526,N_7468);
nand U9458 (N_9458,N_6603,N_6212);
and U9459 (N_9459,N_6971,N_6477);
nor U9460 (N_9460,N_7442,N_6758);
and U9461 (N_9461,N_6879,N_7509);
and U9462 (N_9462,N_7949,N_6703);
or U9463 (N_9463,N_7051,N_7572);
and U9464 (N_9464,N_7786,N_6393);
or U9465 (N_9465,N_7340,N_6107);
nand U9466 (N_9466,N_7578,N_7404);
and U9467 (N_9467,N_6187,N_6717);
and U9468 (N_9468,N_6573,N_7669);
and U9469 (N_9469,N_7903,N_7765);
nor U9470 (N_9470,N_7302,N_6346);
nor U9471 (N_9471,N_6818,N_6708);
and U9472 (N_9472,N_7892,N_6421);
nor U9473 (N_9473,N_7453,N_7288);
or U9474 (N_9474,N_6615,N_7063);
and U9475 (N_9475,N_6960,N_7101);
nor U9476 (N_9476,N_6260,N_7344);
or U9477 (N_9477,N_6887,N_6567);
and U9478 (N_9478,N_7526,N_6686);
xor U9479 (N_9479,N_6408,N_7956);
nor U9480 (N_9480,N_6350,N_7143);
xor U9481 (N_9481,N_7892,N_7439);
nor U9482 (N_9482,N_6881,N_7770);
nand U9483 (N_9483,N_7549,N_6812);
nor U9484 (N_9484,N_7103,N_7463);
nor U9485 (N_9485,N_6525,N_6890);
xnor U9486 (N_9486,N_7818,N_6313);
nand U9487 (N_9487,N_7237,N_7133);
or U9488 (N_9488,N_7534,N_6865);
xnor U9489 (N_9489,N_7495,N_7607);
nand U9490 (N_9490,N_6847,N_7863);
or U9491 (N_9491,N_6590,N_7686);
or U9492 (N_9492,N_6273,N_6120);
nand U9493 (N_9493,N_7403,N_6757);
and U9494 (N_9494,N_7878,N_7981);
nand U9495 (N_9495,N_6800,N_6794);
xor U9496 (N_9496,N_6091,N_6149);
xor U9497 (N_9497,N_6718,N_6736);
or U9498 (N_9498,N_7712,N_6028);
nand U9499 (N_9499,N_7300,N_7428);
nand U9500 (N_9500,N_6178,N_6778);
and U9501 (N_9501,N_6618,N_7162);
and U9502 (N_9502,N_6829,N_7994);
xor U9503 (N_9503,N_6264,N_7395);
and U9504 (N_9504,N_7492,N_7997);
xor U9505 (N_9505,N_7890,N_6877);
or U9506 (N_9506,N_7684,N_6663);
nor U9507 (N_9507,N_6590,N_6065);
nand U9508 (N_9508,N_7341,N_6323);
nor U9509 (N_9509,N_6460,N_7146);
xor U9510 (N_9510,N_6325,N_6301);
and U9511 (N_9511,N_6664,N_6978);
and U9512 (N_9512,N_7625,N_7663);
xnor U9513 (N_9513,N_7427,N_6108);
nor U9514 (N_9514,N_6876,N_7902);
and U9515 (N_9515,N_7091,N_7243);
nand U9516 (N_9516,N_6466,N_7048);
nand U9517 (N_9517,N_6944,N_7976);
and U9518 (N_9518,N_6055,N_7615);
nor U9519 (N_9519,N_7571,N_6709);
nor U9520 (N_9520,N_7382,N_7723);
and U9521 (N_9521,N_6699,N_6697);
xnor U9522 (N_9522,N_6843,N_7561);
and U9523 (N_9523,N_7244,N_6190);
xnor U9524 (N_9524,N_6752,N_7305);
nand U9525 (N_9525,N_6202,N_7884);
and U9526 (N_9526,N_6623,N_7167);
and U9527 (N_9527,N_7289,N_7743);
nand U9528 (N_9528,N_7472,N_6023);
nor U9529 (N_9529,N_6015,N_6611);
or U9530 (N_9530,N_7471,N_6596);
and U9531 (N_9531,N_7670,N_7077);
nor U9532 (N_9532,N_7049,N_6794);
or U9533 (N_9533,N_6573,N_7134);
xnor U9534 (N_9534,N_7446,N_7651);
and U9535 (N_9535,N_6459,N_6120);
nand U9536 (N_9536,N_7952,N_7404);
xnor U9537 (N_9537,N_6623,N_7948);
nor U9538 (N_9538,N_7697,N_7797);
and U9539 (N_9539,N_7390,N_6127);
nor U9540 (N_9540,N_6789,N_7976);
xnor U9541 (N_9541,N_6378,N_7380);
or U9542 (N_9542,N_6802,N_6362);
nor U9543 (N_9543,N_7873,N_6995);
or U9544 (N_9544,N_7704,N_6862);
and U9545 (N_9545,N_7541,N_7448);
nand U9546 (N_9546,N_7131,N_7317);
xnor U9547 (N_9547,N_6113,N_6525);
or U9548 (N_9548,N_6547,N_7592);
nor U9549 (N_9549,N_6135,N_6693);
and U9550 (N_9550,N_7864,N_7101);
or U9551 (N_9551,N_6500,N_7419);
nand U9552 (N_9552,N_7133,N_6567);
or U9553 (N_9553,N_7319,N_7418);
xnor U9554 (N_9554,N_6656,N_6402);
nor U9555 (N_9555,N_7801,N_7348);
or U9556 (N_9556,N_7629,N_6507);
and U9557 (N_9557,N_6467,N_6627);
nand U9558 (N_9558,N_7420,N_6777);
xnor U9559 (N_9559,N_6177,N_6657);
or U9560 (N_9560,N_7978,N_6017);
and U9561 (N_9561,N_7671,N_6618);
nand U9562 (N_9562,N_6902,N_6283);
or U9563 (N_9563,N_7205,N_6668);
nor U9564 (N_9564,N_7429,N_7546);
nor U9565 (N_9565,N_7586,N_7944);
nand U9566 (N_9566,N_7339,N_6785);
and U9567 (N_9567,N_7850,N_6855);
nor U9568 (N_9568,N_7011,N_7650);
or U9569 (N_9569,N_6459,N_7418);
and U9570 (N_9570,N_7625,N_7955);
nor U9571 (N_9571,N_6749,N_7068);
and U9572 (N_9572,N_6934,N_6442);
nor U9573 (N_9573,N_7037,N_7792);
xnor U9574 (N_9574,N_7448,N_6968);
nand U9575 (N_9575,N_6641,N_6843);
xor U9576 (N_9576,N_7476,N_6377);
nand U9577 (N_9577,N_7275,N_6958);
nand U9578 (N_9578,N_7773,N_6453);
and U9579 (N_9579,N_6027,N_6854);
nor U9580 (N_9580,N_6740,N_7403);
nor U9581 (N_9581,N_6631,N_7167);
xnor U9582 (N_9582,N_7837,N_6320);
nand U9583 (N_9583,N_6167,N_6559);
or U9584 (N_9584,N_6423,N_7733);
nand U9585 (N_9585,N_6300,N_6121);
nand U9586 (N_9586,N_7142,N_6952);
nand U9587 (N_9587,N_6450,N_6045);
xnor U9588 (N_9588,N_7409,N_7913);
and U9589 (N_9589,N_7311,N_6695);
xnor U9590 (N_9590,N_6056,N_7259);
nor U9591 (N_9591,N_6077,N_7095);
nor U9592 (N_9592,N_7453,N_6415);
xor U9593 (N_9593,N_6094,N_7700);
xor U9594 (N_9594,N_7827,N_6193);
nor U9595 (N_9595,N_6060,N_6906);
and U9596 (N_9596,N_7042,N_6736);
or U9597 (N_9597,N_6341,N_7536);
and U9598 (N_9598,N_7618,N_6042);
xnor U9599 (N_9599,N_7191,N_6215);
nand U9600 (N_9600,N_6872,N_7989);
or U9601 (N_9601,N_6628,N_7649);
nor U9602 (N_9602,N_6614,N_6226);
nor U9603 (N_9603,N_7111,N_7161);
and U9604 (N_9604,N_7835,N_7788);
nor U9605 (N_9605,N_7395,N_7641);
nor U9606 (N_9606,N_6501,N_7524);
nand U9607 (N_9607,N_6452,N_6342);
and U9608 (N_9608,N_6936,N_7268);
nor U9609 (N_9609,N_7727,N_6494);
and U9610 (N_9610,N_7651,N_6798);
xnor U9611 (N_9611,N_7300,N_6228);
or U9612 (N_9612,N_6659,N_7509);
nor U9613 (N_9613,N_6537,N_7125);
nor U9614 (N_9614,N_7453,N_7501);
nor U9615 (N_9615,N_6779,N_7718);
or U9616 (N_9616,N_6461,N_6058);
and U9617 (N_9617,N_6354,N_7517);
nand U9618 (N_9618,N_7359,N_7601);
and U9619 (N_9619,N_6258,N_7586);
nand U9620 (N_9620,N_6301,N_7038);
and U9621 (N_9621,N_7864,N_7144);
or U9622 (N_9622,N_6376,N_6568);
nand U9623 (N_9623,N_6073,N_6362);
nor U9624 (N_9624,N_7619,N_7413);
or U9625 (N_9625,N_7879,N_7431);
nor U9626 (N_9626,N_7310,N_7714);
nand U9627 (N_9627,N_7447,N_7217);
nor U9628 (N_9628,N_7215,N_7412);
and U9629 (N_9629,N_6876,N_7027);
and U9630 (N_9630,N_6956,N_7697);
nor U9631 (N_9631,N_7803,N_7675);
and U9632 (N_9632,N_7589,N_6454);
or U9633 (N_9633,N_7469,N_6765);
nand U9634 (N_9634,N_6282,N_7881);
and U9635 (N_9635,N_7634,N_6624);
or U9636 (N_9636,N_7511,N_7391);
xnor U9637 (N_9637,N_6690,N_6997);
and U9638 (N_9638,N_7877,N_7997);
nand U9639 (N_9639,N_7752,N_6709);
and U9640 (N_9640,N_6329,N_6393);
or U9641 (N_9641,N_6904,N_7913);
nor U9642 (N_9642,N_6691,N_7841);
or U9643 (N_9643,N_7949,N_7287);
nand U9644 (N_9644,N_6247,N_7472);
xor U9645 (N_9645,N_6554,N_7568);
and U9646 (N_9646,N_7278,N_7157);
nor U9647 (N_9647,N_6247,N_6246);
nand U9648 (N_9648,N_6358,N_7377);
or U9649 (N_9649,N_6458,N_6860);
or U9650 (N_9650,N_6131,N_6893);
nand U9651 (N_9651,N_6664,N_7814);
nand U9652 (N_9652,N_6923,N_7175);
xor U9653 (N_9653,N_6519,N_7489);
and U9654 (N_9654,N_7775,N_6621);
nand U9655 (N_9655,N_6528,N_6922);
nor U9656 (N_9656,N_6704,N_6966);
or U9657 (N_9657,N_7056,N_7168);
nor U9658 (N_9658,N_7667,N_7661);
xnor U9659 (N_9659,N_7979,N_6124);
and U9660 (N_9660,N_7490,N_7021);
nand U9661 (N_9661,N_7969,N_7947);
nor U9662 (N_9662,N_7853,N_7230);
and U9663 (N_9663,N_6360,N_7923);
xor U9664 (N_9664,N_7680,N_6577);
xor U9665 (N_9665,N_6838,N_7734);
xnor U9666 (N_9666,N_7087,N_7978);
nand U9667 (N_9667,N_7174,N_7037);
nor U9668 (N_9668,N_6387,N_6151);
and U9669 (N_9669,N_6843,N_6017);
or U9670 (N_9670,N_6389,N_7320);
or U9671 (N_9671,N_7393,N_7161);
or U9672 (N_9672,N_6049,N_7626);
or U9673 (N_9673,N_6767,N_7042);
nand U9674 (N_9674,N_6493,N_6450);
or U9675 (N_9675,N_7381,N_6719);
nand U9676 (N_9676,N_6351,N_7869);
and U9677 (N_9677,N_7017,N_6689);
xor U9678 (N_9678,N_6183,N_7940);
and U9679 (N_9679,N_7185,N_7911);
or U9680 (N_9680,N_6089,N_7944);
nand U9681 (N_9681,N_6707,N_7399);
xor U9682 (N_9682,N_7292,N_6420);
nand U9683 (N_9683,N_6554,N_7939);
or U9684 (N_9684,N_6060,N_6717);
nor U9685 (N_9685,N_6017,N_6006);
nor U9686 (N_9686,N_7028,N_7928);
nor U9687 (N_9687,N_6706,N_6257);
nand U9688 (N_9688,N_6505,N_6906);
nand U9689 (N_9689,N_6433,N_6134);
or U9690 (N_9690,N_7321,N_6612);
nand U9691 (N_9691,N_7090,N_7144);
nand U9692 (N_9692,N_6269,N_7488);
nand U9693 (N_9693,N_7489,N_6911);
or U9694 (N_9694,N_6106,N_6102);
and U9695 (N_9695,N_7473,N_6872);
nand U9696 (N_9696,N_6449,N_7354);
xnor U9697 (N_9697,N_6215,N_7667);
and U9698 (N_9698,N_7189,N_7659);
and U9699 (N_9699,N_7174,N_6656);
xor U9700 (N_9700,N_6666,N_7032);
xor U9701 (N_9701,N_7974,N_6802);
nor U9702 (N_9702,N_7742,N_7581);
xor U9703 (N_9703,N_6583,N_7128);
xnor U9704 (N_9704,N_6898,N_7100);
nand U9705 (N_9705,N_7916,N_6312);
nor U9706 (N_9706,N_6886,N_6831);
and U9707 (N_9707,N_6994,N_6273);
nand U9708 (N_9708,N_6060,N_7742);
nor U9709 (N_9709,N_6675,N_7771);
nand U9710 (N_9710,N_6518,N_7335);
xor U9711 (N_9711,N_7293,N_6963);
nand U9712 (N_9712,N_6035,N_6705);
xor U9713 (N_9713,N_6713,N_7918);
nand U9714 (N_9714,N_7605,N_6721);
nor U9715 (N_9715,N_7041,N_6082);
or U9716 (N_9716,N_7032,N_6472);
and U9717 (N_9717,N_7458,N_7536);
nand U9718 (N_9718,N_7635,N_6459);
xor U9719 (N_9719,N_6260,N_6928);
nand U9720 (N_9720,N_7039,N_6475);
or U9721 (N_9721,N_7446,N_7765);
nor U9722 (N_9722,N_7848,N_7705);
xnor U9723 (N_9723,N_7699,N_7570);
and U9724 (N_9724,N_6920,N_6202);
xor U9725 (N_9725,N_6733,N_6553);
or U9726 (N_9726,N_6492,N_6513);
or U9727 (N_9727,N_6932,N_6515);
or U9728 (N_9728,N_7184,N_6496);
nor U9729 (N_9729,N_7488,N_7252);
or U9730 (N_9730,N_6875,N_6185);
nand U9731 (N_9731,N_7315,N_6913);
and U9732 (N_9732,N_7193,N_6404);
and U9733 (N_9733,N_7585,N_7881);
nand U9734 (N_9734,N_7986,N_6246);
and U9735 (N_9735,N_6883,N_7243);
or U9736 (N_9736,N_6577,N_6575);
nand U9737 (N_9737,N_7741,N_6296);
or U9738 (N_9738,N_6085,N_6188);
and U9739 (N_9739,N_6801,N_6943);
or U9740 (N_9740,N_7995,N_6346);
xor U9741 (N_9741,N_7036,N_6363);
and U9742 (N_9742,N_7349,N_6686);
nor U9743 (N_9743,N_7988,N_6917);
nor U9744 (N_9744,N_6571,N_7805);
nand U9745 (N_9745,N_7551,N_7004);
and U9746 (N_9746,N_6718,N_7886);
nor U9747 (N_9747,N_6761,N_7061);
or U9748 (N_9748,N_7555,N_6155);
xor U9749 (N_9749,N_7880,N_6563);
xnor U9750 (N_9750,N_7029,N_7777);
nor U9751 (N_9751,N_7677,N_6950);
and U9752 (N_9752,N_7642,N_7150);
nor U9753 (N_9753,N_6096,N_7436);
nand U9754 (N_9754,N_7856,N_6374);
xor U9755 (N_9755,N_6933,N_7665);
xnor U9756 (N_9756,N_6446,N_6979);
or U9757 (N_9757,N_7199,N_7323);
or U9758 (N_9758,N_6862,N_6847);
xor U9759 (N_9759,N_7502,N_6920);
nor U9760 (N_9760,N_7025,N_6628);
and U9761 (N_9761,N_6459,N_7701);
xnor U9762 (N_9762,N_7767,N_7153);
nand U9763 (N_9763,N_6083,N_7708);
or U9764 (N_9764,N_7828,N_6702);
nor U9765 (N_9765,N_6458,N_6985);
xnor U9766 (N_9766,N_7600,N_7627);
or U9767 (N_9767,N_7188,N_6185);
xnor U9768 (N_9768,N_7160,N_6435);
nand U9769 (N_9769,N_7719,N_6773);
xor U9770 (N_9770,N_6031,N_6602);
or U9771 (N_9771,N_6400,N_6972);
and U9772 (N_9772,N_6530,N_7764);
nor U9773 (N_9773,N_7168,N_6363);
nand U9774 (N_9774,N_6597,N_6881);
xor U9775 (N_9775,N_7124,N_6514);
or U9776 (N_9776,N_6537,N_6033);
nand U9777 (N_9777,N_7877,N_6436);
xnor U9778 (N_9778,N_7874,N_7163);
or U9779 (N_9779,N_6288,N_7232);
xnor U9780 (N_9780,N_6293,N_6883);
or U9781 (N_9781,N_7736,N_6577);
xor U9782 (N_9782,N_6341,N_6764);
nand U9783 (N_9783,N_7393,N_7635);
nor U9784 (N_9784,N_6054,N_7368);
nand U9785 (N_9785,N_6911,N_7130);
nand U9786 (N_9786,N_7051,N_7936);
nor U9787 (N_9787,N_7801,N_7048);
or U9788 (N_9788,N_7199,N_6763);
nand U9789 (N_9789,N_6147,N_7711);
nand U9790 (N_9790,N_7666,N_6571);
xnor U9791 (N_9791,N_7715,N_6220);
nand U9792 (N_9792,N_7063,N_7303);
nand U9793 (N_9793,N_7813,N_6510);
or U9794 (N_9794,N_6174,N_6741);
nor U9795 (N_9795,N_6887,N_6688);
nand U9796 (N_9796,N_7224,N_6102);
nand U9797 (N_9797,N_7842,N_6160);
nand U9798 (N_9798,N_7150,N_6432);
and U9799 (N_9799,N_7647,N_6599);
nand U9800 (N_9800,N_7131,N_7874);
nor U9801 (N_9801,N_7499,N_6002);
nor U9802 (N_9802,N_7789,N_7199);
xnor U9803 (N_9803,N_7542,N_7213);
and U9804 (N_9804,N_6714,N_6658);
or U9805 (N_9805,N_6097,N_7103);
xnor U9806 (N_9806,N_6640,N_6720);
nor U9807 (N_9807,N_6075,N_7743);
or U9808 (N_9808,N_6794,N_6873);
and U9809 (N_9809,N_6305,N_7410);
and U9810 (N_9810,N_6948,N_6613);
and U9811 (N_9811,N_6920,N_7443);
and U9812 (N_9812,N_7399,N_7375);
nand U9813 (N_9813,N_6847,N_6842);
nor U9814 (N_9814,N_6875,N_7646);
nor U9815 (N_9815,N_7096,N_6942);
nor U9816 (N_9816,N_6939,N_6832);
nand U9817 (N_9817,N_6328,N_6595);
and U9818 (N_9818,N_6598,N_7581);
or U9819 (N_9819,N_7024,N_6688);
xor U9820 (N_9820,N_6503,N_6312);
nor U9821 (N_9821,N_7722,N_6384);
and U9822 (N_9822,N_6050,N_7661);
nor U9823 (N_9823,N_7182,N_6739);
or U9824 (N_9824,N_7082,N_6293);
nand U9825 (N_9825,N_6369,N_7395);
nor U9826 (N_9826,N_6313,N_7653);
nor U9827 (N_9827,N_7071,N_6813);
and U9828 (N_9828,N_7088,N_7270);
and U9829 (N_9829,N_7868,N_6983);
nor U9830 (N_9830,N_6381,N_6157);
nand U9831 (N_9831,N_6036,N_7216);
and U9832 (N_9832,N_7712,N_7236);
nand U9833 (N_9833,N_6676,N_6603);
xor U9834 (N_9834,N_7047,N_6133);
or U9835 (N_9835,N_6937,N_6529);
nor U9836 (N_9836,N_6453,N_7150);
nor U9837 (N_9837,N_6624,N_6269);
nand U9838 (N_9838,N_6673,N_6930);
nor U9839 (N_9839,N_7887,N_7855);
xor U9840 (N_9840,N_7168,N_7647);
or U9841 (N_9841,N_7987,N_7975);
xnor U9842 (N_9842,N_6341,N_7626);
and U9843 (N_9843,N_7394,N_6267);
or U9844 (N_9844,N_7338,N_6079);
nor U9845 (N_9845,N_7640,N_7921);
or U9846 (N_9846,N_6728,N_6432);
nand U9847 (N_9847,N_7752,N_7867);
nor U9848 (N_9848,N_7118,N_6259);
xor U9849 (N_9849,N_7522,N_6764);
nand U9850 (N_9850,N_7244,N_6114);
nand U9851 (N_9851,N_6565,N_6717);
nor U9852 (N_9852,N_7935,N_6345);
xnor U9853 (N_9853,N_7216,N_7472);
nand U9854 (N_9854,N_7435,N_7544);
or U9855 (N_9855,N_6635,N_6002);
and U9856 (N_9856,N_6710,N_7836);
nor U9857 (N_9857,N_6428,N_6729);
xor U9858 (N_9858,N_7584,N_6423);
and U9859 (N_9859,N_6621,N_7818);
nor U9860 (N_9860,N_6617,N_6890);
or U9861 (N_9861,N_6753,N_6310);
and U9862 (N_9862,N_7442,N_7245);
nand U9863 (N_9863,N_7184,N_7634);
or U9864 (N_9864,N_6802,N_6891);
nand U9865 (N_9865,N_7661,N_6745);
nor U9866 (N_9866,N_6514,N_7331);
xnor U9867 (N_9867,N_7163,N_7483);
nor U9868 (N_9868,N_7782,N_7259);
xor U9869 (N_9869,N_6520,N_7960);
nor U9870 (N_9870,N_6083,N_7936);
or U9871 (N_9871,N_6956,N_7409);
nand U9872 (N_9872,N_7635,N_7155);
xnor U9873 (N_9873,N_7694,N_6013);
or U9874 (N_9874,N_6481,N_6738);
nor U9875 (N_9875,N_6320,N_6722);
and U9876 (N_9876,N_7222,N_6197);
or U9877 (N_9877,N_6857,N_6895);
or U9878 (N_9878,N_6124,N_7829);
nor U9879 (N_9879,N_7705,N_6496);
or U9880 (N_9880,N_6473,N_6297);
and U9881 (N_9881,N_7810,N_6547);
xnor U9882 (N_9882,N_6685,N_6373);
xor U9883 (N_9883,N_6685,N_6302);
nand U9884 (N_9884,N_6509,N_7188);
nand U9885 (N_9885,N_6515,N_6434);
xnor U9886 (N_9886,N_6192,N_6763);
and U9887 (N_9887,N_7782,N_7931);
nor U9888 (N_9888,N_7569,N_7884);
xor U9889 (N_9889,N_6757,N_6285);
xnor U9890 (N_9890,N_6223,N_6069);
xor U9891 (N_9891,N_6036,N_6937);
and U9892 (N_9892,N_6829,N_7406);
nor U9893 (N_9893,N_6122,N_6815);
nand U9894 (N_9894,N_7929,N_7345);
and U9895 (N_9895,N_6078,N_7272);
nand U9896 (N_9896,N_7901,N_7525);
nand U9897 (N_9897,N_7235,N_6117);
or U9898 (N_9898,N_7888,N_7948);
nor U9899 (N_9899,N_7170,N_6553);
and U9900 (N_9900,N_6023,N_7730);
nor U9901 (N_9901,N_6892,N_6357);
and U9902 (N_9902,N_6365,N_6865);
nor U9903 (N_9903,N_6774,N_6009);
and U9904 (N_9904,N_6772,N_6372);
nand U9905 (N_9905,N_6302,N_7207);
nand U9906 (N_9906,N_7198,N_7693);
and U9907 (N_9907,N_7419,N_7046);
or U9908 (N_9908,N_7761,N_6414);
nor U9909 (N_9909,N_7707,N_7176);
xnor U9910 (N_9910,N_6457,N_7796);
and U9911 (N_9911,N_7603,N_7539);
and U9912 (N_9912,N_6477,N_6139);
or U9913 (N_9913,N_7329,N_7420);
or U9914 (N_9914,N_7883,N_7674);
xnor U9915 (N_9915,N_7978,N_7830);
or U9916 (N_9916,N_6546,N_6847);
nor U9917 (N_9917,N_7413,N_6052);
nand U9918 (N_9918,N_7819,N_7573);
and U9919 (N_9919,N_6478,N_6684);
xor U9920 (N_9920,N_7592,N_7044);
nor U9921 (N_9921,N_7578,N_6784);
nor U9922 (N_9922,N_7975,N_7679);
nand U9923 (N_9923,N_7346,N_6608);
and U9924 (N_9924,N_6310,N_7401);
xnor U9925 (N_9925,N_7647,N_7923);
nor U9926 (N_9926,N_6069,N_6490);
xnor U9927 (N_9927,N_6567,N_6246);
xor U9928 (N_9928,N_6825,N_6046);
and U9929 (N_9929,N_6700,N_6009);
xor U9930 (N_9930,N_7406,N_6397);
and U9931 (N_9931,N_7233,N_7191);
nand U9932 (N_9932,N_7853,N_7963);
and U9933 (N_9933,N_6285,N_6722);
xnor U9934 (N_9934,N_6223,N_7654);
xnor U9935 (N_9935,N_7798,N_6165);
and U9936 (N_9936,N_7862,N_7627);
xnor U9937 (N_9937,N_7438,N_6695);
and U9938 (N_9938,N_6056,N_7497);
and U9939 (N_9939,N_7310,N_6085);
or U9940 (N_9940,N_7959,N_6453);
nand U9941 (N_9941,N_7751,N_7664);
and U9942 (N_9942,N_6151,N_6064);
nor U9943 (N_9943,N_6025,N_7958);
or U9944 (N_9944,N_6924,N_6773);
or U9945 (N_9945,N_7914,N_6873);
xor U9946 (N_9946,N_6064,N_7766);
and U9947 (N_9947,N_7134,N_7401);
and U9948 (N_9948,N_7320,N_6746);
nand U9949 (N_9949,N_6342,N_7653);
and U9950 (N_9950,N_6295,N_7969);
nor U9951 (N_9951,N_6667,N_7969);
nor U9952 (N_9952,N_6821,N_6935);
and U9953 (N_9953,N_6380,N_6888);
xor U9954 (N_9954,N_6576,N_6648);
and U9955 (N_9955,N_6372,N_7841);
nand U9956 (N_9956,N_7488,N_7671);
and U9957 (N_9957,N_6834,N_6711);
nand U9958 (N_9958,N_7705,N_6664);
and U9959 (N_9959,N_7855,N_6531);
or U9960 (N_9960,N_6941,N_7588);
or U9961 (N_9961,N_6953,N_7960);
nor U9962 (N_9962,N_6826,N_6386);
and U9963 (N_9963,N_7189,N_7069);
and U9964 (N_9964,N_6345,N_7680);
or U9965 (N_9965,N_6108,N_6929);
nand U9966 (N_9966,N_6524,N_7586);
and U9967 (N_9967,N_7227,N_7220);
nor U9968 (N_9968,N_6250,N_7013);
or U9969 (N_9969,N_7119,N_7232);
nand U9970 (N_9970,N_7130,N_7115);
xnor U9971 (N_9971,N_6648,N_6663);
and U9972 (N_9972,N_7207,N_7454);
or U9973 (N_9973,N_6946,N_6516);
and U9974 (N_9974,N_6954,N_6181);
and U9975 (N_9975,N_7876,N_6286);
or U9976 (N_9976,N_6175,N_6307);
and U9977 (N_9977,N_7975,N_6405);
nand U9978 (N_9978,N_7970,N_6273);
xor U9979 (N_9979,N_6229,N_7687);
and U9980 (N_9980,N_6804,N_7266);
nor U9981 (N_9981,N_7160,N_6007);
xor U9982 (N_9982,N_7501,N_7871);
xor U9983 (N_9983,N_6998,N_6582);
and U9984 (N_9984,N_7977,N_7361);
xnor U9985 (N_9985,N_7409,N_7662);
and U9986 (N_9986,N_6637,N_6246);
and U9987 (N_9987,N_6733,N_6792);
nand U9988 (N_9988,N_6201,N_6203);
and U9989 (N_9989,N_7011,N_6664);
nand U9990 (N_9990,N_7480,N_7903);
nor U9991 (N_9991,N_7297,N_7969);
or U9992 (N_9992,N_7535,N_6034);
or U9993 (N_9993,N_6645,N_7395);
xnor U9994 (N_9994,N_6376,N_6326);
nand U9995 (N_9995,N_6841,N_7409);
and U9996 (N_9996,N_6327,N_7178);
and U9997 (N_9997,N_6702,N_6671);
and U9998 (N_9998,N_7202,N_6140);
or U9999 (N_9999,N_7971,N_6358);
or U10000 (N_10000,N_8619,N_9603);
xnor U10001 (N_10001,N_9222,N_9392);
nor U10002 (N_10002,N_8717,N_9031);
and U10003 (N_10003,N_8061,N_9868);
xnor U10004 (N_10004,N_9946,N_8279);
and U10005 (N_10005,N_9561,N_9905);
xor U10006 (N_10006,N_9146,N_9303);
and U10007 (N_10007,N_8082,N_9852);
and U10008 (N_10008,N_8382,N_8875);
or U10009 (N_10009,N_9756,N_9958);
nor U10010 (N_10010,N_9359,N_9520);
and U10011 (N_10011,N_8750,N_8495);
and U10012 (N_10012,N_8353,N_9036);
or U10013 (N_10013,N_9932,N_8240);
and U10014 (N_10014,N_9763,N_9995);
xor U10015 (N_10015,N_8987,N_8460);
and U10016 (N_10016,N_9509,N_8904);
or U10017 (N_10017,N_9039,N_8538);
nor U10018 (N_10018,N_8981,N_8907);
or U10019 (N_10019,N_9267,N_8975);
nand U10020 (N_10020,N_9655,N_9634);
or U10021 (N_10021,N_8653,N_9348);
or U10022 (N_10022,N_8193,N_8811);
nand U10023 (N_10023,N_8142,N_8326);
or U10024 (N_10024,N_8604,N_8462);
xnor U10025 (N_10025,N_9123,N_8349);
or U10026 (N_10026,N_8077,N_8576);
nand U10027 (N_10027,N_8288,N_9815);
or U10028 (N_10028,N_8978,N_9882);
nand U10029 (N_10029,N_9542,N_9687);
xor U10030 (N_10030,N_9027,N_8095);
nand U10031 (N_10031,N_8085,N_8650);
nand U10032 (N_10032,N_8493,N_9975);
and U10033 (N_10033,N_9326,N_8407);
and U10034 (N_10034,N_8552,N_8694);
nand U10035 (N_10035,N_9840,N_8524);
or U10036 (N_10036,N_9909,N_8503);
nand U10037 (N_10037,N_9902,N_8320);
nand U10038 (N_10038,N_8639,N_9989);
or U10039 (N_10039,N_9481,N_8476);
nor U10040 (N_10040,N_8344,N_8005);
nor U10041 (N_10041,N_8010,N_8885);
and U10042 (N_10042,N_8754,N_8469);
and U10043 (N_10043,N_9839,N_8678);
xor U10044 (N_10044,N_8009,N_9884);
or U10045 (N_10045,N_8986,N_8846);
xnor U10046 (N_10046,N_8672,N_9974);
xnor U10047 (N_10047,N_9112,N_8209);
and U10048 (N_10048,N_9014,N_9981);
nor U10049 (N_10049,N_8671,N_8249);
nor U10050 (N_10050,N_9492,N_9104);
and U10051 (N_10051,N_8970,N_9085);
xnor U10052 (N_10052,N_9211,N_9578);
and U10053 (N_10053,N_8393,N_9693);
nand U10054 (N_10054,N_9056,N_9565);
nand U10055 (N_10055,N_8951,N_8898);
nor U10056 (N_10056,N_9444,N_9695);
xnor U10057 (N_10057,N_8843,N_9585);
nor U10058 (N_10058,N_9507,N_9860);
or U10059 (N_10059,N_8993,N_9851);
nand U10060 (N_10060,N_9414,N_9790);
nand U10061 (N_10061,N_9455,N_8497);
or U10062 (N_10062,N_9526,N_9635);
nor U10063 (N_10063,N_9762,N_8835);
nand U10064 (N_10064,N_8395,N_8807);
xnor U10065 (N_10065,N_9018,N_8120);
nor U10066 (N_10066,N_9160,N_9499);
nand U10067 (N_10067,N_9233,N_9559);
xor U10068 (N_10068,N_9803,N_8518);
nand U10069 (N_10069,N_9052,N_9793);
nand U10070 (N_10070,N_9020,N_9646);
xnor U10071 (N_10071,N_9013,N_8565);
nor U10072 (N_10072,N_9470,N_9371);
or U10073 (N_10073,N_8832,N_9741);
xnor U10074 (N_10074,N_9290,N_8684);
xnor U10075 (N_10075,N_8610,N_8205);
or U10076 (N_10076,N_9870,N_8931);
and U10077 (N_10077,N_9777,N_9621);
nor U10078 (N_10078,N_9260,N_9453);
nand U10079 (N_10079,N_8555,N_9562);
nor U10080 (N_10080,N_8372,N_9147);
xor U10081 (N_10081,N_9678,N_9019);
nand U10082 (N_10082,N_8453,N_9990);
nor U10083 (N_10083,N_8556,N_9458);
xnor U10084 (N_10084,N_8314,N_9699);
xnor U10085 (N_10085,N_9308,N_9084);
xor U10086 (N_10086,N_9152,N_9843);
and U10087 (N_10087,N_8974,N_8581);
xnor U10088 (N_10088,N_8631,N_8792);
nand U10089 (N_10089,N_8128,N_8673);
nor U10090 (N_10090,N_9487,N_8138);
or U10091 (N_10091,N_8785,N_8066);
nor U10092 (N_10092,N_9814,N_9548);
and U10093 (N_10093,N_9445,N_8794);
or U10094 (N_10094,N_8165,N_8661);
xnor U10095 (N_10095,N_9657,N_8872);
nand U10096 (N_10096,N_9755,N_9854);
nand U10097 (N_10097,N_9199,N_9407);
or U10098 (N_10098,N_9970,N_8068);
or U10099 (N_10099,N_9093,N_8571);
or U10100 (N_10100,N_9006,N_9313);
xor U10101 (N_10101,N_8432,N_9328);
xor U10102 (N_10102,N_8458,N_8282);
xnor U10103 (N_10103,N_9581,N_8482);
nand U10104 (N_10104,N_9978,N_9866);
nand U10105 (N_10105,N_8607,N_9571);
and U10106 (N_10106,N_8481,N_9365);
nand U10107 (N_10107,N_9450,N_9574);
or U10108 (N_10108,N_8763,N_9523);
nor U10109 (N_10109,N_9602,N_8541);
or U10110 (N_10110,N_8884,N_9711);
or U10111 (N_10111,N_8246,N_8426);
and U10112 (N_10112,N_8122,N_8459);
xor U10113 (N_10113,N_9441,N_8755);
and U10114 (N_10114,N_9545,N_9721);
nor U10115 (N_10115,N_8420,N_9652);
nand U10116 (N_10116,N_9368,N_9694);
and U10117 (N_10117,N_8615,N_9753);
nor U10118 (N_10118,N_9676,N_8505);
and U10119 (N_10119,N_9286,N_8150);
nand U10120 (N_10120,N_9688,N_8402);
nand U10121 (N_10121,N_9667,N_8212);
xor U10122 (N_10122,N_9847,N_8062);
and U10123 (N_10123,N_8035,N_9181);
xnor U10124 (N_10124,N_8688,N_9088);
nand U10125 (N_10125,N_8526,N_9894);
and U10126 (N_10126,N_9564,N_8919);
nor U10127 (N_10127,N_9383,N_8419);
nor U10128 (N_10128,N_8707,N_9399);
nor U10129 (N_10129,N_9483,N_9660);
xor U10130 (N_10130,N_9729,N_8943);
and U10131 (N_10131,N_8852,N_8112);
nor U10132 (N_10132,N_8236,N_9580);
nor U10133 (N_10133,N_9416,N_8733);
nor U10134 (N_10134,N_9338,N_9618);
xor U10135 (N_10135,N_9924,N_9102);
and U10136 (N_10136,N_9789,N_9823);
nor U10137 (N_10137,N_9236,N_8247);
and U10138 (N_10138,N_9288,N_8043);
and U10139 (N_10139,N_9411,N_9091);
and U10140 (N_10140,N_8848,N_8297);
and U10141 (N_10141,N_9496,N_8421);
nor U10142 (N_10142,N_9828,N_9433);
xor U10143 (N_10143,N_9883,N_9751);
nor U10144 (N_10144,N_9108,N_9479);
nand U10145 (N_10145,N_8098,N_8337);
xor U10146 (N_10146,N_8296,N_8765);
xnor U10147 (N_10147,N_8913,N_9872);
and U10148 (N_10148,N_8443,N_8753);
nand U10149 (N_10149,N_9931,N_8548);
nor U10150 (N_10150,N_9037,N_8024);
nand U10151 (N_10151,N_9822,N_9612);
nor U10152 (N_10152,N_8135,N_9702);
and U10153 (N_10153,N_9493,N_8273);
or U10154 (N_10154,N_9586,N_9448);
xor U10155 (N_10155,N_9669,N_8598);
and U10156 (N_10156,N_8194,N_8131);
xnor U10157 (N_10157,N_9438,N_9215);
or U10158 (N_10158,N_9206,N_9528);
or U10159 (N_10159,N_8034,N_9896);
xnor U10160 (N_10160,N_9053,N_8562);
nand U10161 (N_10161,N_8351,N_9798);
nand U10162 (N_10162,N_8429,N_9259);
nor U10163 (N_10163,N_9796,N_9550);
or U10164 (N_10164,N_8487,N_9302);
or U10165 (N_10165,N_9754,N_8080);
and U10166 (N_10166,N_8692,N_9757);
or U10167 (N_10167,N_8090,N_9390);
or U10168 (N_10168,N_9935,N_8032);
nand U10169 (N_10169,N_8257,N_9269);
nand U10170 (N_10170,N_9519,N_9849);
and U10171 (N_10171,N_8015,N_9381);
and U10172 (N_10172,N_8990,N_9633);
nand U10173 (N_10173,N_8761,N_8837);
or U10174 (N_10174,N_8801,N_9068);
or U10175 (N_10175,N_9820,N_9340);
xor U10176 (N_10176,N_8243,N_8530);
xor U10177 (N_10177,N_9224,N_9255);
and U10178 (N_10178,N_8532,N_8815);
nor U10179 (N_10179,N_9128,N_8767);
and U10180 (N_10180,N_8472,N_8804);
or U10181 (N_10181,N_8543,N_9250);
or U10182 (N_10182,N_8840,N_9080);
xor U10183 (N_10183,N_8011,N_9058);
nor U10184 (N_10184,N_9012,N_8861);
nor U10185 (N_10185,N_8014,N_8119);
nand U10186 (N_10186,N_8307,N_8991);
nand U10187 (N_10187,N_8293,N_8225);
nand U10188 (N_10188,N_8322,N_8271);
or U10189 (N_10189,N_8527,N_8570);
and U10190 (N_10190,N_9280,N_9029);
xor U10191 (N_10191,N_9874,N_9945);
and U10192 (N_10192,N_8736,N_9715);
and U10193 (N_10193,N_8188,N_8957);
nand U10194 (N_10194,N_8850,N_8721);
nor U10195 (N_10195,N_8594,N_9773);
nor U10196 (N_10196,N_8523,N_8956);
xor U10197 (N_10197,N_9588,N_9464);
and U10198 (N_10198,N_8298,N_8466);
or U10199 (N_10199,N_8500,N_8782);
or U10200 (N_10200,N_8896,N_9189);
xnor U10201 (N_10201,N_9480,N_8741);
nor U10202 (N_10202,N_8364,N_9157);
nand U10203 (N_10203,N_9327,N_9130);
xnor U10204 (N_10204,N_9765,N_9343);
and U10205 (N_10205,N_9266,N_8501);
xnor U10206 (N_10206,N_9619,N_9997);
and U10207 (N_10207,N_8882,N_9195);
and U10208 (N_10208,N_9363,N_9922);
xor U10209 (N_10209,N_9462,N_9783);
nor U10210 (N_10210,N_9065,N_9625);
and U10211 (N_10211,N_9473,N_8666);
nand U10212 (N_10212,N_8702,N_8033);
or U10213 (N_10213,N_8647,N_9366);
nand U10214 (N_10214,N_9126,N_8625);
nand U10215 (N_10215,N_9097,N_8632);
nand U10216 (N_10216,N_8396,N_8371);
nor U10217 (N_10217,N_9747,N_8922);
and U10218 (N_10218,N_9074,N_8595);
xor U10219 (N_10219,N_8324,N_9400);
xnor U10220 (N_10220,N_8863,N_8667);
nor U10221 (N_10221,N_8827,N_8682);
nand U10222 (N_10222,N_9976,N_9651);
and U10223 (N_10223,N_8210,N_9082);
nor U10224 (N_10224,N_8108,N_8474);
xor U10225 (N_10225,N_8067,N_9424);
nand U10226 (N_10226,N_9560,N_8113);
nand U10227 (N_10227,N_8367,N_8468);
and U10228 (N_10228,N_9077,N_8308);
xnor U10229 (N_10229,N_9961,N_9740);
nor U10230 (N_10230,N_9437,N_9021);
xor U10231 (N_10231,N_8952,N_9934);
and U10232 (N_10232,N_8747,N_9731);
xor U10233 (N_10233,N_9686,N_9109);
nand U10234 (N_10234,N_9972,N_8380);
nor U10235 (N_10235,N_8039,N_9467);
nor U10236 (N_10236,N_8637,N_9792);
nand U10237 (N_10237,N_8788,N_8584);
xor U10238 (N_10238,N_8044,N_9570);
xor U10239 (N_10239,N_9265,N_9514);
nand U10240 (N_10240,N_9275,N_9857);
or U10241 (N_10241,N_9436,N_9712);
or U10242 (N_10242,N_9639,N_9833);
or U10243 (N_10243,N_9370,N_8040);
nor U10244 (N_10244,N_8966,N_8877);
nor U10245 (N_10245,N_8596,N_8916);
and U10246 (N_10246,N_8302,N_9826);
nor U10247 (N_10247,N_8285,N_9393);
nand U10248 (N_10248,N_8398,N_9957);
nor U10249 (N_10249,N_9501,N_8305);
xor U10250 (N_10250,N_9384,N_8700);
nand U10251 (N_10251,N_9221,N_9690);
and U10252 (N_10252,N_8146,N_9720);
nor U10253 (N_10253,N_9807,N_9168);
nor U10254 (N_10254,N_9906,N_9994);
xnor U10255 (N_10255,N_9697,N_9780);
or U10256 (N_10256,N_9203,N_8434);
nor U10257 (N_10257,N_8016,N_8265);
and U10258 (N_10258,N_8448,N_8748);
xor U10259 (N_10259,N_9670,N_9626);
xor U10260 (N_10260,N_9888,N_8758);
xor U10261 (N_10261,N_9644,N_9497);
or U10262 (N_10262,N_9853,N_8480);
nand U10263 (N_10263,N_8655,N_9532);
and U10264 (N_10264,N_8464,N_9611);
and U10265 (N_10265,N_9703,N_8105);
nand U10266 (N_10266,N_8699,N_8333);
and U10267 (N_10267,N_9179,N_8502);
nand U10268 (N_10268,N_8687,N_8259);
and U10269 (N_10269,N_8433,N_8190);
nor U10270 (N_10270,N_8086,N_9643);
nand U10271 (N_10271,N_9461,N_8202);
or U10272 (N_10272,N_9427,N_9816);
nor U10273 (N_10273,N_9622,N_8787);
nor U10274 (N_10274,N_8118,N_9926);
nand U10275 (N_10275,N_8348,N_9795);
xnor U10276 (N_10276,N_9916,N_8979);
nand U10277 (N_10277,N_8718,N_8473);
nand U10278 (N_10278,N_8756,N_8779);
xnor U10279 (N_10279,N_9017,N_8231);
or U10280 (N_10280,N_9447,N_9836);
and U10281 (N_10281,N_8477,N_9598);
or U10282 (N_10282,N_8719,N_8720);
xor U10283 (N_10283,N_9724,N_8329);
nor U10284 (N_10284,N_9537,N_8002);
xor U10285 (N_10285,N_9351,N_8134);
or U10286 (N_10286,N_9806,N_9330);
xor U10287 (N_10287,N_9398,N_8640);
nor U10288 (N_10288,N_8844,N_8816);
and U10289 (N_10289,N_8154,N_8689);
and U10290 (N_10290,N_9797,N_8441);
and U10291 (N_10291,N_9805,N_8902);
nor U10292 (N_10292,N_8341,N_9425);
or U10293 (N_10293,N_8544,N_8310);
xor U10294 (N_10294,N_9463,N_9318);
xor U10295 (N_10295,N_9775,N_8802);
nor U10296 (N_10296,N_9918,N_9204);
xnor U10297 (N_10297,N_9738,N_8964);
nand U10298 (N_10298,N_8643,N_9417);
nor U10299 (N_10299,N_8511,N_9558);
or U10300 (N_10300,N_9604,N_8186);
or U10301 (N_10301,N_9245,N_8597);
xnor U10302 (N_10302,N_8173,N_8892);
nor U10303 (N_10303,N_8006,N_8217);
nand U10304 (N_10304,N_8281,N_9979);
and U10305 (N_10305,N_8102,N_8819);
nand U10306 (N_10306,N_8440,N_9165);
xnor U10307 (N_10307,N_8343,N_8680);
and U10308 (N_10308,N_9734,N_9406);
nor U10309 (N_10309,N_9120,N_9389);
or U10310 (N_10310,N_8796,N_8063);
nor U10311 (N_10311,N_9886,N_8050);
or U10312 (N_10312,N_9048,N_8908);
nand U10313 (N_10313,N_8143,N_9388);
or U10314 (N_10314,N_9525,N_8430);
xnor U10315 (N_10315,N_8409,N_9664);
xor U10316 (N_10316,N_9372,N_9426);
or U10317 (N_10317,N_8490,N_9422);
or U10318 (N_10318,N_8554,N_9730);
xor U10319 (N_10319,N_8886,N_8470);
xnor U10320 (N_10320,N_9547,N_9282);
nand U10321 (N_10321,N_8946,N_8375);
nor U10322 (N_10322,N_8723,N_9614);
or U10323 (N_10323,N_9767,N_8764);
nor U10324 (N_10324,N_8439,N_9605);
xor U10325 (N_10325,N_9881,N_9156);
or U10326 (N_10326,N_9878,N_8897);
or U10327 (N_10327,N_8879,N_9268);
nor U10328 (N_10328,N_9040,N_9373);
or U10329 (N_10329,N_9219,N_9837);
and U10330 (N_10330,N_9107,N_8578);
and U10331 (N_10331,N_9804,N_8603);
xnor U10332 (N_10332,N_8001,N_9539);
and U10333 (N_10333,N_8740,N_8325);
and U10334 (N_10334,N_8726,N_8809);
or U10335 (N_10335,N_8638,N_8945);
or U10336 (N_10336,N_8444,N_9025);
nor U10337 (N_10337,N_9759,N_8561);
and U10338 (N_10338,N_9358,N_8838);
xnor U10339 (N_10339,N_8590,N_8608);
or U10340 (N_10340,N_8483,N_8323);
xnor U10341 (N_10341,N_8905,N_9124);
or U10342 (N_10342,N_9440,N_8864);
nand U10343 (N_10343,N_9022,N_9246);
nand U10344 (N_10344,N_9354,N_9861);
and U10345 (N_10345,N_9682,N_8114);
nand U10346 (N_10346,N_8315,N_9799);
nor U10347 (N_10347,N_8769,N_8036);
nor U10348 (N_10348,N_8287,N_9319);
nor U10349 (N_10349,N_9379,N_8642);
xnor U10350 (N_10350,N_9394,N_9498);
xor U10351 (N_10351,N_9166,N_8139);
or U10352 (N_10352,N_8378,N_8716);
or U10353 (N_10353,N_9555,N_9835);
nand U10354 (N_10354,N_9593,N_8727);
and U10355 (N_10355,N_9725,N_8703);
and U10356 (N_10356,N_9845,N_8573);
or U10357 (N_10357,N_9346,N_8049);
or U10358 (N_10358,N_9484,N_8064);
xnor U10359 (N_10359,N_8575,N_8903);
nand U10360 (N_10360,N_8232,N_9158);
xor U10361 (N_10361,N_8182,N_8600);
xnor U10362 (N_10362,N_8037,N_8332);
or U10363 (N_10363,N_8317,N_8950);
nand U10364 (N_10364,N_9198,N_8158);
and U10365 (N_10365,N_8256,N_9940);
or U10366 (N_10366,N_8424,N_9364);
xnor U10367 (N_10367,N_8599,N_8374);
and U10368 (N_10368,N_9210,N_9901);
nand U10369 (N_10369,N_9985,N_8346);
nor U10370 (N_10370,N_9925,N_9802);
xor U10371 (N_10371,N_9701,N_9412);
and U10372 (N_10372,N_8521,N_8651);
nand U10373 (N_10373,N_9929,N_9276);
nand U10374 (N_10374,N_8883,N_9552);
nand U10375 (N_10375,N_8629,N_8274);
nand U10376 (N_10376,N_8797,N_8551);
and U10377 (N_10377,N_9530,N_8592);
nor U10378 (N_10378,N_9468,N_9681);
xnor U10379 (N_10379,N_9505,N_8550);
or U10380 (N_10380,N_8825,N_9596);
nand U10381 (N_10381,N_9449,N_9794);
nor U10382 (N_10382,N_8805,N_8289);
and U10383 (N_10383,N_9671,N_9067);
and U10384 (N_10384,N_9167,N_8888);
nand U10385 (N_10385,N_8226,N_8609);
and U10386 (N_10386,N_8025,N_8878);
xor U10387 (N_10387,N_8253,N_9549);
nor U10388 (N_10388,N_9451,N_8160);
or U10389 (N_10389,N_9457,N_8789);
nor U10390 (N_10390,N_9324,N_9674);
nand U10391 (N_10391,N_8413,N_8645);
and U10392 (N_10392,N_8177,N_9594);
nor U10393 (N_10393,N_9534,N_9201);
nand U10394 (N_10394,N_8512,N_8620);
xnor U10395 (N_10395,N_9111,N_9270);
or U10396 (N_10396,N_9685,N_9531);
or U10397 (N_10397,N_9766,N_8277);
or U10398 (N_10398,N_8577,N_8152);
nand U10399 (N_10399,N_9274,N_9791);
or U10400 (N_10400,N_9758,N_8774);
xor U10401 (N_10401,N_9778,N_8073);
and U10402 (N_10402,N_8762,N_9915);
or U10403 (N_10403,N_9010,N_8627);
or U10404 (N_10404,N_8547,N_8397);
and U10405 (N_10405,N_9421,N_8646);
nor U10406 (N_10406,N_9933,N_9876);
nor U10407 (N_10407,N_9912,N_8557);
xor U10408 (N_10408,N_9454,N_9873);
nand U10409 (N_10409,N_9846,N_8821);
nor U10410 (N_10410,N_9941,N_9174);
xor U10411 (N_10411,N_8242,N_8633);
nor U10412 (N_10412,N_9408,N_9774);
nand U10413 (N_10413,N_9164,N_8893);
nor U10414 (N_10414,N_9956,N_9714);
and U10415 (N_10415,N_9554,N_9927);
nand U10416 (N_10416,N_8553,N_8824);
or U10417 (N_10417,N_9887,N_9046);
xor U10418 (N_10418,N_9698,N_9051);
xnor U10419 (N_10419,N_8621,N_8301);
nand U10420 (N_10420,N_8130,N_8766);
and U10421 (N_10421,N_9446,N_8405);
and U10422 (N_10422,N_8545,N_9435);
nor U10423 (N_10423,N_8982,N_8685);
xor U10424 (N_10424,N_8569,N_8461);
xor U10425 (N_10425,N_9810,N_8187);
xor U10426 (N_10426,N_8536,N_8652);
xnor U10427 (N_10427,N_8962,N_9648);
xor U10428 (N_10428,N_9175,N_9289);
nand U10429 (N_10429,N_9551,N_9154);
and U10430 (N_10430,N_9576,N_8076);
nand U10431 (N_10431,N_8808,N_8911);
and U10432 (N_10432,N_9101,N_9035);
xnor U10433 (N_10433,N_8047,N_9728);
xor U10434 (N_10434,N_9817,N_8665);
nand U10435 (N_10435,N_9063,N_9813);
xor U10436 (N_10436,N_9098,N_9103);
and U10437 (N_10437,N_9196,N_9726);
xnor U10438 (N_10438,N_8294,N_8427);
nor U10439 (N_10439,N_9137,N_9538);
or U10440 (N_10440,N_9248,N_9298);
and U10441 (N_10441,N_8742,N_8959);
nor U10442 (N_10442,N_8997,N_9066);
and U10443 (N_10443,N_9362,N_8038);
or U10444 (N_10444,N_8944,N_8504);
and U10445 (N_10445,N_8963,N_9138);
or U10446 (N_10446,N_9824,N_8948);
or U10447 (N_10447,N_9613,N_9234);
or U10448 (N_10448,N_8084,N_8304);
nor U10449 (N_10449,N_8980,N_8901);
and U10450 (N_10450,N_8677,N_9903);
nand U10451 (N_10451,N_9277,N_9044);
nor U10452 (N_10452,N_8972,N_8436);
or U10453 (N_10453,N_9966,N_9984);
nor U10454 (N_10454,N_9291,N_8075);
nand U10455 (N_10455,N_8938,N_8059);
nor U10456 (N_10456,N_9704,N_9415);
nand U10457 (N_10457,N_8841,N_8412);
xnor U10458 (N_10458,N_8830,N_8617);
and U10459 (N_10459,N_9899,N_9991);
xor U10460 (N_10460,N_8255,N_8089);
xnor U10461 (N_10461,N_9038,N_9629);
nand U10462 (N_10462,N_9008,N_8862);
nor U10463 (N_10463,N_9808,N_9423);
and U10464 (N_10464,N_8391,N_9785);
and U10465 (N_10465,N_8347,N_9919);
and U10466 (N_10466,N_9344,N_8601);
nor U10467 (N_10467,N_8664,N_9567);
and U10468 (N_10468,N_8517,N_8201);
and U10469 (N_10469,N_9404,N_9471);
xnor U10470 (N_10470,N_9689,N_9591);
nor U10471 (N_10471,N_8096,N_9663);
or U10472 (N_10472,N_9092,N_9659);
and U10473 (N_10473,N_9079,N_8379);
nand U10474 (N_10474,N_9508,N_9015);
and U10475 (N_10475,N_9375,N_8213);
nor U10476 (N_10476,N_9769,N_8939);
and U10477 (N_10477,N_8008,N_8491);
nor U10478 (N_10478,N_8737,N_9786);
xor U10479 (N_10479,N_9069,N_9396);
nand U10480 (N_10480,N_9113,N_9485);
nor U10481 (N_10481,N_9736,N_8934);
nor U10482 (N_10482,N_9263,N_8318);
xnor U10483 (N_10483,N_9475,N_9335);
xnor U10484 (N_10484,N_8280,N_8313);
nand U10485 (N_10485,N_8184,N_9942);
or U10486 (N_10486,N_9770,N_8568);
or U10487 (N_10487,N_8052,N_9750);
or U10488 (N_10488,N_9776,N_9026);
and U10489 (N_10489,N_9176,N_8299);
xor U10490 (N_10490,N_9477,N_8269);
or U10491 (N_10491,N_8151,N_8350);
nand U10492 (N_10492,N_8057,N_8670);
xor U10493 (N_10493,N_8091,N_8106);
and U10494 (N_10494,N_8780,N_9227);
nand U10495 (N_10495,N_8546,N_8284);
nand U10496 (N_10496,N_8218,N_9656);
nand U10497 (N_10497,N_9439,N_8923);
nor U10498 (N_10498,N_9996,N_8083);
nor U10499 (N_10499,N_9739,N_9054);
xnor U10500 (N_10500,N_8199,N_9830);
and U10501 (N_10501,N_8869,N_8989);
and U10502 (N_10502,N_9281,N_8705);
nand U10503 (N_10503,N_9161,N_8206);
nor U10504 (N_10504,N_8880,N_9615);
nor U10505 (N_10505,N_9705,N_9336);
and U10506 (N_10506,N_8960,N_9380);
xnor U10507 (N_10507,N_8278,N_8836);
or U10508 (N_10508,N_8856,N_8549);
and U10509 (N_10509,N_9768,N_8924);
nor U10510 (N_10510,N_9000,N_9959);
and U10511 (N_10511,N_8339,N_9331);
nor U10512 (N_10512,N_8826,N_9139);
and U10513 (N_10513,N_9541,N_9601);
and U10514 (N_10514,N_9304,N_8626);
or U10515 (N_10515,N_8053,N_8858);
or U10516 (N_10516,N_8810,N_9980);
nand U10517 (N_10517,N_9858,N_9148);
xnor U10518 (N_10518,N_8484,N_8567);
and U10519 (N_10519,N_8370,N_9679);
xor U10520 (N_10520,N_8196,N_8401);
nand U10521 (N_10521,N_9301,N_8634);
and U10522 (N_10522,N_9235,N_8799);
and U10523 (N_10523,N_9350,N_8749);
or U10524 (N_10524,N_8657,N_8947);
or U10525 (N_10525,N_8069,N_8498);
or U10526 (N_10526,N_9131,N_9913);
nor U10527 (N_10527,N_8812,N_8178);
or U10528 (N_10528,N_9049,N_9320);
and U10529 (N_10529,N_8855,N_9251);
xnor U10530 (N_10530,N_8697,N_9993);
and U10531 (N_10531,N_9733,N_8051);
nor U10532 (N_10532,N_8630,N_9095);
xor U10533 (N_10533,N_8912,N_9352);
nor U10534 (N_10534,N_8081,N_8522);
nand U10535 (N_10535,N_8528,N_8996);
xor U10536 (N_10536,N_8909,N_9465);
nor U10537 (N_10537,N_9050,N_9502);
or U10538 (N_10538,N_8784,N_9361);
nor U10539 (N_10539,N_9583,N_8928);
nor U10540 (N_10540,N_8715,N_8475);
and U10541 (N_10541,N_8360,N_8334);
nor U10542 (N_10542,N_8696,N_8262);
or U10543 (N_10543,N_8701,N_9937);
or U10544 (N_10544,N_9977,N_8712);
and U10545 (N_10545,N_8790,N_8157);
and U10546 (N_10546,N_8589,N_9231);
nor U10547 (N_10547,N_9610,N_8890);
and U10548 (N_10548,N_9118,N_8820);
or U10549 (N_10549,N_9764,N_8985);
xnor U10550 (N_10550,N_8239,N_8013);
or U10551 (N_10551,N_8478,N_8669);
nand U10552 (N_10552,N_8926,N_8676);
and U10553 (N_10553,N_9030,N_8456);
or U10554 (N_10554,N_8492,N_8170);
and U10555 (N_10555,N_8215,N_9413);
nand U10556 (N_10556,N_8731,N_9781);
nand U10557 (N_10557,N_9105,N_8839);
nor U10558 (N_10558,N_9722,N_9316);
nor U10559 (N_10559,N_9033,N_8183);
xnor U10560 (N_10560,N_9954,N_9880);
nor U10561 (N_10561,N_8261,N_9761);
nand U10562 (N_10562,N_9047,N_9673);
and U10563 (N_10563,N_9829,N_8539);
and U10564 (N_10564,N_9294,N_8219);
and U10565 (N_10565,N_9595,N_9947);
xnor U10566 (N_10566,N_9078,N_9043);
or U10567 (N_10567,N_8300,N_8961);
xor U10568 (N_10568,N_9510,N_9297);
nand U10569 (N_10569,N_8849,N_8254);
nor U10570 (N_10570,N_9258,N_8734);
and U10571 (N_10571,N_9513,N_8115);
and U10572 (N_10572,N_8874,N_9184);
nor U10573 (N_10573,N_8531,N_8778);
xor U10574 (N_10574,N_9240,N_8935);
and U10575 (N_10575,N_9228,N_9329);
or U10576 (N_10576,N_8203,N_9938);
or U10577 (N_10577,N_8007,N_8342);
nor U10578 (N_10578,N_8887,N_9662);
xnor U10579 (N_10579,N_8866,N_8463);
nor U10580 (N_10580,N_9936,N_8221);
nor U10581 (N_10581,N_9784,N_8148);
or U10582 (N_10582,N_9237,N_8168);
or U10583 (N_10583,N_9200,N_9299);
and U10584 (N_10584,N_9072,N_9710);
nand U10585 (N_10585,N_8127,N_9232);
or U10586 (N_10586,N_9332,N_9821);
nor U10587 (N_10587,N_8854,N_8927);
nor U10588 (N_10588,N_8408,N_8829);
nand U10589 (N_10589,N_8316,N_8361);
and U10590 (N_10590,N_9623,N_8070);
nor U10591 (N_10591,N_8161,N_9382);
xor U10592 (N_10592,N_9600,N_8983);
or U10593 (N_10593,N_8616,N_8410);
xnor U10594 (N_10594,N_8169,N_9864);
and U10595 (N_10595,N_8965,N_9127);
or U10596 (N_10596,N_9135,N_8691);
nor U10597 (N_10597,N_8662,N_9986);
nor U10598 (N_10598,N_8713,N_8582);
nand U10599 (N_10599,N_9296,N_8233);
nand U10600 (N_10600,N_8976,N_9489);
nand U10601 (N_10601,N_9386,N_9708);
xnor U10602 (N_10602,N_9914,N_8823);
xnor U10603 (N_10603,N_8452,N_8932);
nand U10604 (N_10604,N_9748,N_8681);
xor U10605 (N_10605,N_9125,N_8937);
nor U10606 (N_10606,N_8977,N_9247);
xnor U10607 (N_10607,N_8454,N_8605);
xor U10608 (N_10608,N_9832,N_8675);
nor U10609 (N_10609,N_8865,N_9322);
xor U10610 (N_10610,N_8704,N_9194);
xnor U10611 (N_10611,N_8435,N_8414);
xor U10612 (N_10612,N_9252,N_8759);
and U10613 (N_10613,N_8847,N_8229);
xnor U10614 (N_10614,N_8358,N_9772);
xnor U10615 (N_10615,N_9202,N_9007);
xor U10616 (N_10616,N_8588,N_9818);
xnor U10617 (N_10617,N_8654,N_8906);
nor U10618 (N_10618,N_8074,N_8079);
and U10619 (N_10619,N_8772,N_8563);
or U10620 (N_10620,N_8881,N_8026);
nor U10621 (N_10621,N_8376,N_8097);
nand U10622 (N_10622,N_8735,N_9410);
nor U10623 (N_10623,N_8660,N_8003);
xor U10624 (N_10624,N_8450,N_9587);
xnor U10625 (N_10625,N_8999,N_9630);
nor U10626 (N_10626,N_8828,N_9185);
nand U10627 (N_10627,N_8529,N_8399);
and U10628 (N_10628,N_8775,N_9811);
or U10629 (N_10629,N_9208,N_9420);
and U10630 (N_10630,N_8593,N_9192);
xnor U10631 (N_10631,N_9086,N_9556);
or U10632 (N_10632,N_9142,N_9609);
nand U10633 (N_10633,N_8258,N_8058);
nand U10634 (N_10634,N_9838,N_9672);
or U10635 (N_10635,N_9005,N_9675);
nor U10636 (N_10636,N_8163,N_8635);
nand U10637 (N_10637,N_8352,N_9136);
xor U10638 (N_10638,N_8579,N_9094);
or U10639 (N_10639,N_8228,N_9190);
and U10640 (N_10640,N_9223,N_9355);
xor U10641 (N_10641,N_9443,N_8771);
and U10642 (N_10642,N_9511,N_8770);
nand U10643 (N_10643,N_9023,N_8175);
or U10644 (N_10644,N_8123,N_8994);
xnor U10645 (N_10645,N_9073,N_9254);
and U10646 (N_10646,N_8611,N_9921);
nand U10647 (N_10647,N_8695,N_9998);
and U10648 (N_10648,N_9300,N_8428);
xor U10649 (N_10649,N_8394,N_9582);
nor U10650 (N_10650,N_8649,N_8817);
or U10651 (N_10651,N_9284,N_8969);
and U10652 (N_10652,N_9920,N_9771);
and U10653 (N_10653,N_9314,N_9209);
and U10654 (N_10654,N_8319,N_9917);
nor U10655 (N_10655,N_9746,N_8252);
nand U10656 (N_10656,N_9879,N_9645);
nand U10657 (N_10657,N_8383,N_9885);
nor U10658 (N_10658,N_8690,N_8622);
nor U10659 (N_10659,N_9272,N_8519);
nand U10660 (N_10660,N_8744,N_8743);
nand U10661 (N_10661,N_9628,N_8018);
or U10662 (N_10662,N_9939,N_9982);
nor U10663 (N_10663,N_9287,N_8418);
and U10664 (N_10664,N_8822,N_9983);
and U10665 (N_10665,N_8133,N_8560);
and U10666 (N_10666,N_9692,N_9647);
and U10667 (N_10667,N_8377,N_9661);
nor U10668 (N_10668,N_8683,N_8729);
nor U10669 (N_10669,N_9034,N_9306);
or U10670 (N_10670,N_8499,N_8048);
nor U10671 (N_10671,N_8768,N_8533);
or U10672 (N_10672,N_8191,N_8189);
nand U10673 (N_10673,N_8968,N_9649);
or U10674 (N_10674,N_9869,N_8384);
or U10675 (N_10675,N_9114,N_8998);
and U10676 (N_10676,N_8208,N_9032);
and U10677 (N_10677,N_9512,N_8783);
and U10678 (N_10678,N_8386,N_8251);
or U10679 (N_10679,N_8023,N_9476);
nand U10680 (N_10680,N_8354,N_9096);
and U10681 (N_10681,N_9875,N_9121);
and U10682 (N_10682,N_9169,N_8535);
or U10683 (N_10683,N_8515,N_9460);
xor U10684 (N_10684,N_8751,N_9141);
xor U10685 (N_10685,N_9178,N_9521);
and U10686 (N_10686,N_8818,N_9402);
or U10687 (N_10687,N_9787,N_9491);
nor U10688 (N_10688,N_9907,N_9391);
xnor U10689 (N_10689,N_8200,N_8117);
or U10690 (N_10690,N_9419,N_8942);
xnor U10691 (N_10691,N_9191,N_8659);
xor U10692 (N_10692,N_9244,N_8489);
xor U10693 (N_10693,N_9650,N_8357);
or U10694 (N_10694,N_8275,N_8292);
nand U10695 (N_10695,N_8859,N_9723);
and U10696 (N_10696,N_8663,N_9533);
or U10697 (N_10697,N_8895,N_9323);
and U10698 (N_10698,N_9638,N_8853);
xor U10699 (N_10699,N_8129,N_8156);
nor U10700 (N_10700,N_8752,N_9469);
xnor U10701 (N_10701,N_9242,N_9897);
nor U10702 (N_10702,N_9944,N_9271);
xor U10703 (N_10703,N_8416,N_9599);
xor U10704 (N_10704,N_8776,N_9517);
xnor U10705 (N_10705,N_8510,N_9950);
nor U10706 (N_10706,N_9405,N_9825);
nand U10707 (N_10707,N_8078,N_8107);
xor U10708 (N_10708,N_8583,N_8915);
or U10709 (N_10709,N_9948,N_8936);
nor U10710 (N_10710,N_9295,N_9841);
nand U10711 (N_10711,N_9225,N_9606);
and U10712 (N_10712,N_8425,N_8363);
or U10713 (N_10713,N_8728,N_8447);
or U10714 (N_10714,N_8648,N_9357);
nor U10715 (N_10715,N_9642,N_8141);
or U10716 (N_10716,N_8263,N_8693);
or U10717 (N_10717,N_8929,N_9910);
or U10718 (N_10718,N_9238,N_8111);
nor U10719 (N_10719,N_9334,N_9713);
nand U10720 (N_10720,N_9064,N_8155);
or U10721 (N_10721,N_9495,N_9001);
and U10722 (N_10722,N_9877,N_9760);
and U10723 (N_10723,N_8870,N_9430);
nor U10724 (N_10724,N_9486,N_9133);
and U10725 (N_10725,N_8270,N_9700);
and U10726 (N_10726,N_9684,N_9253);
xnor U10727 (N_10727,N_9083,N_9653);
xnor U10728 (N_10728,N_9011,N_9812);
and U10729 (N_10729,N_9749,N_8041);
nor U10730 (N_10730,N_9557,N_8000);
or U10731 (N_10731,N_8746,N_8021);
xnor U10732 (N_10732,N_8054,N_9418);
nor U10733 (N_10733,N_9273,N_8368);
nor U10734 (N_10734,N_9856,N_9953);
xnor U10735 (N_10735,N_8359,N_9898);
nand U10736 (N_10736,N_8658,N_8973);
and U10737 (N_10737,N_9212,N_8224);
and U10738 (N_10738,N_9627,N_9009);
or U10739 (N_10739,N_8004,N_9187);
xor U10740 (N_10740,N_9145,N_9665);
xor U10741 (N_10741,N_9339,N_8028);
xor U10742 (N_10742,N_9801,N_8910);
and U10743 (N_10743,N_8223,N_9041);
and U10744 (N_10744,N_8591,N_8803);
xnor U10745 (N_10745,N_8471,N_9850);
nand U10746 (N_10746,N_9395,N_8438);
nor U10747 (N_10747,N_9143,N_9683);
or U10748 (N_10748,N_9385,N_9960);
or U10749 (N_10749,N_9170,N_8558);
xnor U10750 (N_10750,N_8967,N_8136);
xnor U10751 (N_10751,N_8668,N_9967);
nand U10752 (N_10752,N_8507,N_8921);
nand U10753 (N_10753,N_9374,N_9516);
nor U10754 (N_10754,N_8109,N_9230);
nor U10755 (N_10755,N_8030,N_8101);
xnor U10756 (N_10756,N_8791,N_9640);
or U10757 (N_10757,N_8406,N_8404);
xnor U10758 (N_10758,N_9590,N_9999);
nand U10759 (N_10759,N_9800,N_9264);
and U10760 (N_10760,N_9891,N_8508);
nor U10761 (N_10761,N_8525,N_8800);
nor U10762 (N_10762,N_8708,N_9459);
xnor U10763 (N_10763,N_9973,N_9862);
nand U10764 (N_10764,N_9620,N_8509);
xnor U10765 (N_10765,N_8092,N_9317);
and U10766 (N_10766,N_9149,N_8268);
nor U10767 (N_10767,N_8137,N_8389);
nor U10768 (N_10768,N_8814,N_9024);
nand U10769 (N_10769,N_8722,N_8385);
or U10770 (N_10770,N_8714,N_8045);
nand U10771 (N_10771,N_8520,N_9589);
and U10772 (N_10772,N_9522,N_8873);
xnor U10773 (N_10773,N_8777,N_9536);
nand U10774 (N_10774,N_9285,N_8295);
nor U10775 (N_10775,N_8710,N_8309);
nor U10776 (N_10776,N_9397,N_9220);
nor U10777 (N_10777,N_9930,N_8834);
nand U10778 (N_10778,N_8506,N_9356);
nand U10779 (N_10779,N_9177,N_9709);
nand U10780 (N_10780,N_9293,N_8781);
xor U10781 (N_10781,N_9305,N_9428);
and U10782 (N_10782,N_9827,N_8871);
xor U10783 (N_10783,N_8250,N_9333);
xor U10784 (N_10784,N_8730,N_9923);
nand U10785 (N_10785,N_8586,N_9378);
nor U10786 (N_10786,N_8618,N_9106);
and U10787 (N_10787,N_9257,N_9871);
and U10788 (N_10788,N_9431,N_8711);
nand U10789 (N_10789,N_9745,N_9188);
nor U10790 (N_10790,N_9955,N_9535);
nor U10791 (N_10791,N_8335,N_9243);
xor U10792 (N_10792,N_9442,N_8925);
nor U10793 (N_10793,N_8366,N_8988);
nor U10794 (N_10794,N_8954,N_8159);
nor U10795 (N_10795,N_9969,N_8709);
or U10796 (N_10796,N_8496,N_8486);
nor U10797 (N_10797,N_8798,N_9071);
and U10798 (N_10798,N_9341,N_9844);
xor U10799 (N_10799,N_8345,N_8857);
xor U10800 (N_10800,N_8833,N_8423);
xor U10801 (N_10801,N_9159,N_8636);
or U10802 (N_10802,N_8216,N_9719);
xor U10803 (N_10803,N_8914,N_9680);
xnor U10804 (N_10804,N_8185,N_9577);
or U10805 (N_10805,N_8773,N_9387);
nor U10806 (N_10806,N_9952,N_9151);
or U10807 (N_10807,N_9345,N_8894);
nand U10808 (N_10808,N_8328,N_8312);
nand U10809 (N_10809,N_9500,N_9003);
and U10810 (N_10810,N_8147,N_9403);
nor U10811 (N_10811,N_9732,N_9488);
and U10812 (N_10812,N_8920,N_8172);
xor U10813 (N_10813,N_8264,N_9456);
xor U10814 (N_10814,N_8171,N_9060);
nand U10815 (N_10815,N_9089,N_9893);
xnor U10816 (N_10816,N_8167,N_8940);
or U10817 (N_10817,N_8116,N_8267);
xnor U10818 (N_10818,N_8235,N_9226);
nand U10819 (N_10819,N_9075,N_8060);
and U10820 (N_10820,N_9434,N_8411);
and U10821 (N_10821,N_8534,N_8286);
nand U10822 (N_10822,N_9213,N_8140);
and U10823 (N_10823,N_8056,N_9090);
xnor U10824 (N_10824,N_9472,N_8564);
nand U10825 (N_10825,N_8104,N_8455);
or U10826 (N_10826,N_8451,N_8362);
or U10827 (N_10827,N_9908,N_9057);
and U10828 (N_10828,N_8181,N_9658);
xnor U10829 (N_10829,N_9217,N_8124);
xor U10830 (N_10830,N_9788,N_8027);
or U10831 (N_10831,N_9988,N_8306);
xnor U10832 (N_10832,N_9173,N_8479);
nor U10833 (N_10833,N_9241,N_9218);
nor U10834 (N_10834,N_9597,N_8400);
or U10835 (N_10835,N_9307,N_8022);
or U10836 (N_10836,N_8153,N_9115);
nor U10837 (N_10837,N_9632,N_9119);
nor U10838 (N_10838,N_9518,N_9490);
and U10839 (N_10839,N_8392,N_8738);
and U10840 (N_10840,N_8889,N_9150);
nand U10841 (N_10841,N_9311,N_9949);
nand U10842 (N_10842,N_8485,N_8851);
or U10843 (N_10843,N_8516,N_8340);
or U10844 (N_10844,N_9968,N_9309);
or U10845 (N_10845,N_9855,N_9377);
nor U10846 (N_10846,N_9342,N_9707);
xor U10847 (N_10847,N_8046,N_9409);
xor U10848 (N_10848,N_8237,N_8204);
nand U10849 (N_10849,N_8706,N_8180);
nand U10850 (N_10850,N_9087,N_9900);
xnor U10851 (N_10851,N_8446,N_9834);
or U10852 (N_10852,N_8984,N_8248);
or U10853 (N_10853,N_9964,N_9546);
or U10854 (N_10854,N_8559,N_8587);
or U10855 (N_10855,N_9249,N_8327);
or U10856 (N_10856,N_9863,N_9134);
nand U10857 (N_10857,N_8786,N_8930);
nand U10858 (N_10858,N_8900,N_9608);
or U10859 (N_10859,N_8031,N_9677);
nor U10860 (N_10860,N_9216,N_8793);
xor U10861 (N_10861,N_9055,N_9261);
or U10862 (N_10862,N_8422,N_9592);
nand U10863 (N_10863,N_9140,N_8065);
nor U10864 (N_10864,N_8126,N_8388);
xnor U10865 (N_10865,N_9506,N_9256);
and U10866 (N_10866,N_9325,N_8806);
and U10867 (N_10867,N_8145,N_9744);
xor U10868 (N_10868,N_9347,N_8012);
or U10869 (N_10869,N_8941,N_9666);
xnor U10870 (N_10870,N_9717,N_8121);
and U10871 (N_10871,N_9572,N_9752);
nand U10872 (N_10872,N_9737,N_9239);
xnor U10873 (N_10873,N_9278,N_8876);
xnor U10874 (N_10874,N_9016,N_9004);
nor U10875 (N_10875,N_8745,N_8971);
and U10876 (N_10876,N_8390,N_8088);
nor U10877 (N_10877,N_9292,N_8207);
xnor U10878 (N_10878,N_8757,N_9193);
or U10879 (N_10879,N_8195,N_8211);
nor U10880 (N_10880,N_9116,N_9691);
and U10881 (N_10881,N_8260,N_8029);
and U10882 (N_10882,N_9515,N_9895);
or U10883 (N_10883,N_8132,N_8099);
nor U10884 (N_10884,N_8628,N_9965);
nor U10885 (N_10885,N_8760,N_9819);
nand U10886 (N_10886,N_8387,N_9070);
xnor U10887 (N_10887,N_9831,N_9452);
nor U10888 (N_10888,N_8356,N_9214);
nand U10889 (N_10889,N_8087,N_9735);
and U10890 (N_10890,N_9474,N_9617);
or U10891 (N_10891,N_8336,N_9859);
or U10892 (N_10892,N_8679,N_8241);
nand U10893 (N_10893,N_9129,N_8860);
or U10894 (N_10894,N_8019,N_8641);
or U10895 (N_10895,N_8891,N_8071);
or U10896 (N_10896,N_8656,N_9262);
and U10897 (N_10897,N_9099,N_9573);
nor U10898 (N_10898,N_9279,N_8513);
or U10899 (N_10899,N_8125,N_8276);
nand U10900 (N_10900,N_9637,N_9987);
nor U10901 (N_10901,N_9197,N_8110);
nand U10902 (N_10902,N_8093,N_8415);
xor U10903 (N_10903,N_8020,N_9172);
nand U10904 (N_10904,N_9706,N_8238);
or U10905 (N_10905,N_8574,N_9062);
and U10906 (N_10906,N_8540,N_9575);
or U10907 (N_10907,N_8542,N_9943);
nand U10908 (N_10908,N_8623,N_8192);
and U10909 (N_10909,N_8613,N_9229);
nand U10910 (N_10910,N_8732,N_8698);
or U10911 (N_10911,N_8234,N_8899);
nor U10912 (N_10912,N_9045,N_9478);
and U10913 (N_10913,N_9321,N_8179);
or U10914 (N_10914,N_8953,N_8955);
or U10915 (N_10915,N_9892,N_8842);
nand U10916 (N_10916,N_8725,N_8813);
and U10917 (N_10917,N_9059,N_9186);
and U10918 (N_10918,N_9002,N_9081);
xor U10919 (N_10919,N_9527,N_9636);
nand U10920 (N_10920,N_9616,N_9171);
and U10921 (N_10921,N_9503,N_8149);
nand U10922 (N_10922,N_8949,N_8227);
nor U10923 (N_10923,N_8330,N_9809);
nor U10924 (N_10924,N_8369,N_9122);
and U10925 (N_10925,N_9100,N_8176);
xnor U10926 (N_10926,N_8686,N_9042);
and U10927 (N_10927,N_8331,N_8724);
xor U10928 (N_10928,N_8457,N_9207);
nor U10929 (N_10929,N_9992,N_9727);
xnor U10930 (N_10930,N_9742,N_8612);
or U10931 (N_10931,N_9962,N_8995);
and U10932 (N_10932,N_8321,N_8290);
nor U10933 (N_10933,N_9544,N_9696);
and U10934 (N_10934,N_8585,N_9155);
xnor U10935 (N_10935,N_8266,N_9779);
nand U10936 (N_10936,N_9432,N_9654);
or U10937 (N_10937,N_9641,N_8933);
nor U10938 (N_10938,N_9494,N_9718);
and U10939 (N_10939,N_9568,N_9716);
and U10940 (N_10940,N_8867,N_8245);
nand U10941 (N_10941,N_8214,N_9117);
nand U10942 (N_10942,N_8222,N_9028);
xnor U10943 (N_10943,N_9504,N_9668);
or U10944 (N_10944,N_9529,N_9367);
nand U10945 (N_10945,N_8144,N_8220);
nor U10946 (N_10946,N_8614,N_8417);
or U10947 (N_10947,N_9890,N_8100);
nand U10948 (N_10948,N_9624,N_8230);
xor U10949 (N_10949,N_9429,N_9553);
nand U10950 (N_10950,N_9144,N_9963);
and U10951 (N_10951,N_9337,N_8055);
or U10952 (N_10952,N_9482,N_9182);
and U10953 (N_10953,N_9563,N_8442);
or U10954 (N_10954,N_8845,N_8373);
or U10955 (N_10955,N_9743,N_8272);
nor U10956 (N_10956,N_9904,N_9163);
xor U10957 (N_10957,N_9283,N_8283);
and U10958 (N_10958,N_8918,N_8403);
nand U10959 (N_10959,N_9061,N_8958);
and U10960 (N_10960,N_9867,N_8338);
nor U10961 (N_10961,N_8488,N_8602);
xnor U10962 (N_10962,N_9566,N_8166);
or U10963 (N_10963,N_8103,N_9153);
nor U10964 (N_10964,N_8795,N_9911);
nor U10965 (N_10965,N_9353,N_8465);
xor U10966 (N_10966,N_9180,N_9569);
nand U10967 (N_10967,N_8992,N_9360);
and U10968 (N_10968,N_9132,N_8624);
or U10969 (N_10969,N_8674,N_8437);
nor U10970 (N_10970,N_8303,N_9205);
xnor U10971 (N_10971,N_8494,N_9928);
and U10972 (N_10972,N_9466,N_8162);
and U10973 (N_10973,N_8197,N_8094);
nor U10974 (N_10974,N_8572,N_8244);
xor U10975 (N_10975,N_8355,N_8445);
nand U10976 (N_10976,N_9369,N_9865);
or U10977 (N_10977,N_8644,N_9543);
xor U10978 (N_10978,N_9631,N_9889);
xor U10979 (N_10979,N_8739,N_8537);
nand U10980 (N_10980,N_8174,N_9349);
and U10981 (N_10981,N_8467,N_8514);
and U10982 (N_10982,N_8431,N_9607);
xnor U10983 (N_10983,N_8365,N_8164);
and U10984 (N_10984,N_8198,N_9076);
xnor U10985 (N_10985,N_8917,N_8449);
nand U10986 (N_10986,N_9310,N_9524);
xor U10987 (N_10987,N_8580,N_8072);
and U10988 (N_10988,N_9782,N_9376);
nor U10989 (N_10989,N_9848,N_9842);
or U10990 (N_10990,N_9540,N_9110);
nor U10991 (N_10991,N_8868,N_9315);
nor U10992 (N_10992,N_9579,N_8291);
or U10993 (N_10993,N_9951,N_8606);
nand U10994 (N_10994,N_8042,N_9312);
and U10995 (N_10995,N_9584,N_9183);
and U10996 (N_10996,N_8831,N_9401);
and U10997 (N_10997,N_8017,N_8381);
nor U10998 (N_10998,N_9971,N_8311);
or U10999 (N_10999,N_8566,N_9162);
nand U11000 (N_11000,N_9565,N_9397);
xnor U11001 (N_11001,N_9379,N_8761);
nand U11002 (N_11002,N_8299,N_8345);
nand U11003 (N_11003,N_9115,N_9884);
xnor U11004 (N_11004,N_8795,N_9460);
nand U11005 (N_11005,N_9072,N_8374);
xnor U11006 (N_11006,N_9077,N_8815);
or U11007 (N_11007,N_9706,N_9658);
nand U11008 (N_11008,N_8710,N_9302);
or U11009 (N_11009,N_9170,N_9781);
or U11010 (N_11010,N_8845,N_9674);
and U11011 (N_11011,N_8015,N_9617);
nand U11012 (N_11012,N_8031,N_9915);
nor U11013 (N_11013,N_8081,N_9414);
nand U11014 (N_11014,N_9029,N_8079);
xnor U11015 (N_11015,N_9979,N_8541);
xnor U11016 (N_11016,N_8226,N_8312);
and U11017 (N_11017,N_9259,N_8759);
or U11018 (N_11018,N_9854,N_9113);
xor U11019 (N_11019,N_8363,N_9520);
xor U11020 (N_11020,N_9309,N_9146);
or U11021 (N_11021,N_9193,N_9816);
and U11022 (N_11022,N_8719,N_8942);
xnor U11023 (N_11023,N_9280,N_9304);
xnor U11024 (N_11024,N_9755,N_9916);
or U11025 (N_11025,N_9489,N_9922);
xor U11026 (N_11026,N_8392,N_9700);
and U11027 (N_11027,N_9707,N_9818);
and U11028 (N_11028,N_8572,N_8474);
nand U11029 (N_11029,N_8064,N_8995);
nor U11030 (N_11030,N_8914,N_8488);
nand U11031 (N_11031,N_8634,N_9263);
xnor U11032 (N_11032,N_9908,N_8228);
or U11033 (N_11033,N_9351,N_8835);
or U11034 (N_11034,N_8753,N_8269);
or U11035 (N_11035,N_9904,N_8268);
nand U11036 (N_11036,N_8217,N_8127);
nand U11037 (N_11037,N_8595,N_8849);
nand U11038 (N_11038,N_9899,N_9318);
nor U11039 (N_11039,N_9780,N_9614);
or U11040 (N_11040,N_9067,N_8877);
or U11041 (N_11041,N_9678,N_8847);
nand U11042 (N_11042,N_9232,N_9949);
nor U11043 (N_11043,N_9327,N_8317);
xnor U11044 (N_11044,N_8698,N_8119);
xor U11045 (N_11045,N_8612,N_8115);
or U11046 (N_11046,N_9839,N_8589);
nand U11047 (N_11047,N_8642,N_9795);
or U11048 (N_11048,N_8766,N_8206);
or U11049 (N_11049,N_9226,N_9018);
xor U11050 (N_11050,N_9767,N_8746);
or U11051 (N_11051,N_9873,N_9624);
xnor U11052 (N_11052,N_8889,N_8549);
and U11053 (N_11053,N_8314,N_9336);
nand U11054 (N_11054,N_9508,N_8423);
nor U11055 (N_11055,N_9637,N_8988);
xor U11056 (N_11056,N_9414,N_9306);
nand U11057 (N_11057,N_9124,N_9493);
or U11058 (N_11058,N_8091,N_8609);
or U11059 (N_11059,N_9160,N_9009);
and U11060 (N_11060,N_9307,N_9823);
nor U11061 (N_11061,N_8289,N_8167);
nand U11062 (N_11062,N_8428,N_9808);
or U11063 (N_11063,N_8479,N_9601);
nor U11064 (N_11064,N_8976,N_9195);
and U11065 (N_11065,N_8984,N_8127);
nand U11066 (N_11066,N_8135,N_8239);
nor U11067 (N_11067,N_9914,N_8410);
nor U11068 (N_11068,N_9582,N_9678);
nand U11069 (N_11069,N_9216,N_8259);
nor U11070 (N_11070,N_9626,N_9028);
nor U11071 (N_11071,N_8197,N_9608);
and U11072 (N_11072,N_8655,N_8979);
nor U11073 (N_11073,N_9737,N_9780);
nand U11074 (N_11074,N_8493,N_9581);
and U11075 (N_11075,N_8458,N_9012);
nor U11076 (N_11076,N_9603,N_9067);
nor U11077 (N_11077,N_9366,N_9422);
or U11078 (N_11078,N_9480,N_9321);
nor U11079 (N_11079,N_9908,N_8026);
xor U11080 (N_11080,N_8442,N_9072);
and U11081 (N_11081,N_8244,N_8923);
xor U11082 (N_11082,N_8199,N_8177);
or U11083 (N_11083,N_9096,N_9800);
and U11084 (N_11084,N_9934,N_8174);
and U11085 (N_11085,N_8355,N_9205);
nor U11086 (N_11086,N_9794,N_9353);
or U11087 (N_11087,N_9803,N_8860);
xnor U11088 (N_11088,N_9153,N_9238);
nor U11089 (N_11089,N_8741,N_9113);
or U11090 (N_11090,N_9963,N_8682);
and U11091 (N_11091,N_8623,N_9514);
nor U11092 (N_11092,N_8102,N_9926);
or U11093 (N_11093,N_9311,N_8425);
and U11094 (N_11094,N_8765,N_9087);
or U11095 (N_11095,N_8799,N_9786);
or U11096 (N_11096,N_8460,N_8119);
or U11097 (N_11097,N_8701,N_8035);
nor U11098 (N_11098,N_9629,N_8816);
and U11099 (N_11099,N_8167,N_8407);
xor U11100 (N_11100,N_9266,N_8654);
or U11101 (N_11101,N_8386,N_8249);
nor U11102 (N_11102,N_8888,N_8966);
or U11103 (N_11103,N_8333,N_9682);
xnor U11104 (N_11104,N_9368,N_8212);
or U11105 (N_11105,N_8416,N_9842);
xor U11106 (N_11106,N_9514,N_9828);
xor U11107 (N_11107,N_8217,N_8112);
nand U11108 (N_11108,N_8570,N_9728);
or U11109 (N_11109,N_8641,N_9290);
nand U11110 (N_11110,N_9990,N_9118);
xnor U11111 (N_11111,N_9190,N_8937);
or U11112 (N_11112,N_8903,N_8227);
and U11113 (N_11113,N_8944,N_8454);
and U11114 (N_11114,N_9008,N_9477);
and U11115 (N_11115,N_9867,N_8974);
xnor U11116 (N_11116,N_8268,N_9068);
nand U11117 (N_11117,N_8108,N_9818);
or U11118 (N_11118,N_9612,N_9993);
nor U11119 (N_11119,N_9082,N_8658);
xor U11120 (N_11120,N_9984,N_9000);
nand U11121 (N_11121,N_8685,N_8173);
nor U11122 (N_11122,N_9200,N_8236);
xnor U11123 (N_11123,N_8285,N_8756);
nor U11124 (N_11124,N_8774,N_8029);
and U11125 (N_11125,N_9828,N_9922);
nor U11126 (N_11126,N_8566,N_9104);
or U11127 (N_11127,N_8696,N_8381);
nor U11128 (N_11128,N_8445,N_8325);
and U11129 (N_11129,N_8361,N_9357);
and U11130 (N_11130,N_9636,N_8002);
nand U11131 (N_11131,N_8305,N_8901);
xnor U11132 (N_11132,N_8692,N_8422);
nand U11133 (N_11133,N_8055,N_9028);
nand U11134 (N_11134,N_8090,N_9433);
or U11135 (N_11135,N_9453,N_9083);
xor U11136 (N_11136,N_9828,N_9626);
nand U11137 (N_11137,N_9678,N_8792);
xor U11138 (N_11138,N_8493,N_9722);
and U11139 (N_11139,N_9612,N_8565);
nand U11140 (N_11140,N_9058,N_9233);
and U11141 (N_11141,N_9351,N_8152);
nand U11142 (N_11142,N_8510,N_9314);
or U11143 (N_11143,N_8456,N_8682);
xor U11144 (N_11144,N_8528,N_8878);
or U11145 (N_11145,N_8230,N_9457);
nand U11146 (N_11146,N_8648,N_9740);
nand U11147 (N_11147,N_9148,N_9927);
nor U11148 (N_11148,N_9024,N_9638);
nor U11149 (N_11149,N_9904,N_9362);
nor U11150 (N_11150,N_8384,N_8947);
or U11151 (N_11151,N_8548,N_9890);
nor U11152 (N_11152,N_8630,N_9176);
and U11153 (N_11153,N_8265,N_8257);
or U11154 (N_11154,N_8920,N_9112);
nor U11155 (N_11155,N_8948,N_8914);
or U11156 (N_11156,N_9281,N_9333);
nand U11157 (N_11157,N_9128,N_9207);
nand U11158 (N_11158,N_9010,N_9018);
nor U11159 (N_11159,N_9716,N_8134);
nand U11160 (N_11160,N_9751,N_9169);
nor U11161 (N_11161,N_9136,N_8244);
nor U11162 (N_11162,N_8591,N_8306);
and U11163 (N_11163,N_9174,N_8828);
nor U11164 (N_11164,N_9902,N_9705);
nor U11165 (N_11165,N_8086,N_8146);
nand U11166 (N_11166,N_8646,N_9854);
or U11167 (N_11167,N_9802,N_8694);
xnor U11168 (N_11168,N_9420,N_9031);
or U11169 (N_11169,N_8716,N_9295);
xnor U11170 (N_11170,N_8855,N_8000);
nor U11171 (N_11171,N_9580,N_9812);
and U11172 (N_11172,N_9037,N_9674);
and U11173 (N_11173,N_9644,N_8164);
and U11174 (N_11174,N_8183,N_8634);
or U11175 (N_11175,N_8162,N_9875);
and U11176 (N_11176,N_8330,N_9688);
nand U11177 (N_11177,N_8736,N_9066);
nor U11178 (N_11178,N_9732,N_9207);
and U11179 (N_11179,N_8844,N_9326);
xor U11180 (N_11180,N_8860,N_8279);
or U11181 (N_11181,N_8100,N_9532);
nand U11182 (N_11182,N_9592,N_9629);
nand U11183 (N_11183,N_8307,N_8287);
nand U11184 (N_11184,N_8544,N_8479);
and U11185 (N_11185,N_8821,N_9946);
or U11186 (N_11186,N_9973,N_8345);
nor U11187 (N_11187,N_9421,N_8293);
nand U11188 (N_11188,N_8245,N_9824);
xor U11189 (N_11189,N_8441,N_9845);
nand U11190 (N_11190,N_9283,N_8454);
or U11191 (N_11191,N_8281,N_8162);
and U11192 (N_11192,N_9193,N_9391);
nand U11193 (N_11193,N_9100,N_9910);
and U11194 (N_11194,N_8877,N_8047);
nand U11195 (N_11195,N_9768,N_8539);
nor U11196 (N_11196,N_9869,N_9380);
and U11197 (N_11197,N_8865,N_8875);
and U11198 (N_11198,N_8374,N_8722);
nor U11199 (N_11199,N_8624,N_9214);
nor U11200 (N_11200,N_8803,N_8733);
xnor U11201 (N_11201,N_8306,N_9110);
nand U11202 (N_11202,N_8522,N_8507);
nand U11203 (N_11203,N_9781,N_8811);
nor U11204 (N_11204,N_8640,N_8024);
or U11205 (N_11205,N_9063,N_8761);
nand U11206 (N_11206,N_9269,N_9866);
and U11207 (N_11207,N_8740,N_9164);
nand U11208 (N_11208,N_8634,N_9214);
and U11209 (N_11209,N_9103,N_8303);
xnor U11210 (N_11210,N_8170,N_8633);
or U11211 (N_11211,N_8241,N_9917);
xnor U11212 (N_11212,N_8893,N_9293);
nor U11213 (N_11213,N_8417,N_9071);
xnor U11214 (N_11214,N_9708,N_9757);
and U11215 (N_11215,N_8628,N_9840);
or U11216 (N_11216,N_8498,N_8222);
nand U11217 (N_11217,N_8758,N_8511);
nand U11218 (N_11218,N_9081,N_9057);
or U11219 (N_11219,N_9125,N_8973);
xnor U11220 (N_11220,N_9416,N_8178);
xnor U11221 (N_11221,N_9625,N_8391);
and U11222 (N_11222,N_8543,N_9434);
xnor U11223 (N_11223,N_9342,N_9194);
and U11224 (N_11224,N_8542,N_9158);
nor U11225 (N_11225,N_9433,N_8884);
xnor U11226 (N_11226,N_9656,N_9858);
nor U11227 (N_11227,N_8068,N_8033);
and U11228 (N_11228,N_8271,N_8704);
xor U11229 (N_11229,N_8537,N_9110);
nor U11230 (N_11230,N_9481,N_8240);
nand U11231 (N_11231,N_8641,N_8872);
or U11232 (N_11232,N_9705,N_9386);
nor U11233 (N_11233,N_8193,N_9949);
and U11234 (N_11234,N_8294,N_8475);
nand U11235 (N_11235,N_8490,N_9033);
and U11236 (N_11236,N_9973,N_8774);
xor U11237 (N_11237,N_8720,N_8297);
nand U11238 (N_11238,N_8521,N_9130);
or U11239 (N_11239,N_9802,N_8422);
xor U11240 (N_11240,N_8145,N_8728);
and U11241 (N_11241,N_9374,N_8513);
nor U11242 (N_11242,N_8151,N_8464);
or U11243 (N_11243,N_8833,N_8210);
nor U11244 (N_11244,N_8521,N_8868);
or U11245 (N_11245,N_9979,N_8178);
xnor U11246 (N_11246,N_9355,N_9793);
nor U11247 (N_11247,N_8685,N_9789);
and U11248 (N_11248,N_8391,N_8519);
nor U11249 (N_11249,N_8458,N_8799);
nor U11250 (N_11250,N_9197,N_8126);
nor U11251 (N_11251,N_9894,N_9862);
nor U11252 (N_11252,N_9751,N_8731);
nor U11253 (N_11253,N_9574,N_9565);
nor U11254 (N_11254,N_8733,N_9676);
and U11255 (N_11255,N_9460,N_9428);
nor U11256 (N_11256,N_8978,N_8195);
nand U11257 (N_11257,N_8544,N_8929);
nand U11258 (N_11258,N_9543,N_9672);
nor U11259 (N_11259,N_9622,N_9692);
nor U11260 (N_11260,N_9234,N_9338);
nor U11261 (N_11261,N_8537,N_8226);
and U11262 (N_11262,N_9060,N_9904);
xnor U11263 (N_11263,N_9806,N_9234);
or U11264 (N_11264,N_8795,N_8065);
and U11265 (N_11265,N_9726,N_8606);
nand U11266 (N_11266,N_8802,N_9219);
and U11267 (N_11267,N_8523,N_9206);
xnor U11268 (N_11268,N_9418,N_9446);
nand U11269 (N_11269,N_8347,N_8668);
xor U11270 (N_11270,N_9620,N_9294);
and U11271 (N_11271,N_8129,N_9574);
xnor U11272 (N_11272,N_8477,N_8562);
nand U11273 (N_11273,N_9903,N_9606);
nand U11274 (N_11274,N_9255,N_8550);
xnor U11275 (N_11275,N_8531,N_8896);
or U11276 (N_11276,N_8208,N_8833);
nor U11277 (N_11277,N_8972,N_8301);
nor U11278 (N_11278,N_9087,N_8895);
nor U11279 (N_11279,N_8028,N_9769);
xnor U11280 (N_11280,N_9160,N_8768);
nor U11281 (N_11281,N_8470,N_8560);
and U11282 (N_11282,N_8608,N_9747);
or U11283 (N_11283,N_9597,N_9943);
and U11284 (N_11284,N_8790,N_9594);
or U11285 (N_11285,N_9330,N_9465);
nand U11286 (N_11286,N_9747,N_9148);
nor U11287 (N_11287,N_9037,N_9582);
and U11288 (N_11288,N_8493,N_9417);
or U11289 (N_11289,N_8536,N_9006);
nor U11290 (N_11290,N_8188,N_8843);
nand U11291 (N_11291,N_9399,N_9847);
and U11292 (N_11292,N_9703,N_9082);
xnor U11293 (N_11293,N_9004,N_8889);
xor U11294 (N_11294,N_8306,N_8654);
or U11295 (N_11295,N_9365,N_8914);
or U11296 (N_11296,N_8700,N_9902);
nor U11297 (N_11297,N_8677,N_8183);
and U11298 (N_11298,N_9605,N_9481);
nor U11299 (N_11299,N_9534,N_8402);
xor U11300 (N_11300,N_9760,N_9346);
nand U11301 (N_11301,N_9748,N_8039);
and U11302 (N_11302,N_8533,N_8520);
nor U11303 (N_11303,N_8295,N_8778);
nand U11304 (N_11304,N_9941,N_8989);
and U11305 (N_11305,N_8498,N_9363);
and U11306 (N_11306,N_9198,N_8284);
and U11307 (N_11307,N_9666,N_8803);
or U11308 (N_11308,N_9998,N_8749);
or U11309 (N_11309,N_8583,N_9879);
and U11310 (N_11310,N_8675,N_8338);
nor U11311 (N_11311,N_9338,N_8412);
nand U11312 (N_11312,N_9115,N_9970);
or U11313 (N_11313,N_9078,N_8507);
and U11314 (N_11314,N_9877,N_9719);
nor U11315 (N_11315,N_9184,N_8656);
xor U11316 (N_11316,N_8928,N_9502);
nor U11317 (N_11317,N_9509,N_9677);
and U11318 (N_11318,N_9461,N_9113);
or U11319 (N_11319,N_8728,N_9752);
nor U11320 (N_11320,N_8478,N_9024);
or U11321 (N_11321,N_8057,N_9143);
nand U11322 (N_11322,N_9800,N_8918);
xor U11323 (N_11323,N_8452,N_9581);
and U11324 (N_11324,N_8935,N_8033);
nand U11325 (N_11325,N_9193,N_9732);
xor U11326 (N_11326,N_8773,N_8989);
nand U11327 (N_11327,N_8834,N_9826);
and U11328 (N_11328,N_8043,N_8280);
or U11329 (N_11329,N_9253,N_9126);
nor U11330 (N_11330,N_8335,N_9684);
or U11331 (N_11331,N_9749,N_8136);
xor U11332 (N_11332,N_8472,N_9516);
or U11333 (N_11333,N_8822,N_9865);
nand U11334 (N_11334,N_9711,N_9229);
or U11335 (N_11335,N_8171,N_9161);
nor U11336 (N_11336,N_8949,N_8443);
nand U11337 (N_11337,N_9383,N_8559);
nand U11338 (N_11338,N_8893,N_9356);
xnor U11339 (N_11339,N_9775,N_8594);
xor U11340 (N_11340,N_9667,N_8657);
and U11341 (N_11341,N_9074,N_8534);
and U11342 (N_11342,N_9233,N_9882);
nand U11343 (N_11343,N_8047,N_9422);
xnor U11344 (N_11344,N_9198,N_8456);
and U11345 (N_11345,N_9203,N_9128);
and U11346 (N_11346,N_9801,N_8621);
xnor U11347 (N_11347,N_9465,N_9289);
nand U11348 (N_11348,N_9480,N_8103);
nand U11349 (N_11349,N_8130,N_8600);
nand U11350 (N_11350,N_9465,N_9883);
nor U11351 (N_11351,N_9658,N_9476);
nor U11352 (N_11352,N_9263,N_9026);
and U11353 (N_11353,N_8730,N_9350);
nor U11354 (N_11354,N_8436,N_8777);
and U11355 (N_11355,N_8273,N_8786);
or U11356 (N_11356,N_8444,N_9335);
and U11357 (N_11357,N_9953,N_9874);
nand U11358 (N_11358,N_8919,N_9430);
nor U11359 (N_11359,N_8903,N_9335);
or U11360 (N_11360,N_9167,N_8524);
or U11361 (N_11361,N_8715,N_8985);
nand U11362 (N_11362,N_9445,N_8357);
xnor U11363 (N_11363,N_8125,N_9714);
and U11364 (N_11364,N_9708,N_9694);
or U11365 (N_11365,N_9675,N_9734);
and U11366 (N_11366,N_8272,N_9110);
nand U11367 (N_11367,N_9183,N_9786);
xor U11368 (N_11368,N_9789,N_8041);
nand U11369 (N_11369,N_9296,N_9979);
and U11370 (N_11370,N_9254,N_9601);
xnor U11371 (N_11371,N_9069,N_8931);
xnor U11372 (N_11372,N_9673,N_8042);
nor U11373 (N_11373,N_9432,N_9770);
and U11374 (N_11374,N_9338,N_9911);
or U11375 (N_11375,N_9351,N_8310);
nand U11376 (N_11376,N_9161,N_9096);
nor U11377 (N_11377,N_9108,N_9453);
or U11378 (N_11378,N_8133,N_8856);
and U11379 (N_11379,N_9394,N_8168);
nor U11380 (N_11380,N_8040,N_8187);
or U11381 (N_11381,N_8881,N_8465);
nand U11382 (N_11382,N_8375,N_9589);
and U11383 (N_11383,N_8202,N_8441);
and U11384 (N_11384,N_8004,N_9888);
nor U11385 (N_11385,N_9631,N_9977);
and U11386 (N_11386,N_9455,N_9805);
and U11387 (N_11387,N_8512,N_8054);
nor U11388 (N_11388,N_9887,N_9659);
nor U11389 (N_11389,N_9512,N_8593);
xnor U11390 (N_11390,N_8133,N_9763);
xor U11391 (N_11391,N_9113,N_9257);
or U11392 (N_11392,N_9004,N_9897);
xor U11393 (N_11393,N_9265,N_8658);
and U11394 (N_11394,N_9724,N_8876);
and U11395 (N_11395,N_8457,N_8933);
nand U11396 (N_11396,N_8835,N_8863);
nand U11397 (N_11397,N_9829,N_9618);
nor U11398 (N_11398,N_8885,N_8359);
and U11399 (N_11399,N_9071,N_8398);
or U11400 (N_11400,N_8203,N_8639);
nand U11401 (N_11401,N_9017,N_8985);
and U11402 (N_11402,N_9977,N_9529);
or U11403 (N_11403,N_8659,N_8675);
and U11404 (N_11404,N_9676,N_8523);
and U11405 (N_11405,N_9941,N_9123);
and U11406 (N_11406,N_8026,N_8425);
nand U11407 (N_11407,N_8688,N_9689);
or U11408 (N_11408,N_9333,N_9713);
nor U11409 (N_11409,N_9570,N_9182);
and U11410 (N_11410,N_8977,N_9283);
or U11411 (N_11411,N_8817,N_9274);
nor U11412 (N_11412,N_8352,N_9547);
or U11413 (N_11413,N_9213,N_9425);
nor U11414 (N_11414,N_8869,N_9575);
or U11415 (N_11415,N_8379,N_9986);
and U11416 (N_11416,N_8988,N_8771);
nand U11417 (N_11417,N_9065,N_9988);
nor U11418 (N_11418,N_9536,N_9044);
nand U11419 (N_11419,N_8347,N_8880);
nand U11420 (N_11420,N_8118,N_9742);
and U11421 (N_11421,N_9495,N_9318);
nor U11422 (N_11422,N_9127,N_9987);
or U11423 (N_11423,N_8431,N_9259);
nor U11424 (N_11424,N_8054,N_9759);
or U11425 (N_11425,N_8549,N_8886);
nor U11426 (N_11426,N_9934,N_9864);
or U11427 (N_11427,N_8367,N_8061);
or U11428 (N_11428,N_8888,N_9599);
nand U11429 (N_11429,N_8547,N_9348);
or U11430 (N_11430,N_8251,N_8227);
nor U11431 (N_11431,N_9624,N_9963);
nor U11432 (N_11432,N_8390,N_9094);
nand U11433 (N_11433,N_9892,N_8906);
and U11434 (N_11434,N_9777,N_8386);
xor U11435 (N_11435,N_8118,N_8147);
xnor U11436 (N_11436,N_9476,N_9657);
and U11437 (N_11437,N_9296,N_9387);
and U11438 (N_11438,N_8240,N_8759);
nor U11439 (N_11439,N_9391,N_8890);
and U11440 (N_11440,N_9061,N_8672);
and U11441 (N_11441,N_8451,N_9014);
nor U11442 (N_11442,N_8753,N_9357);
nor U11443 (N_11443,N_9925,N_9743);
and U11444 (N_11444,N_9753,N_8389);
nor U11445 (N_11445,N_8027,N_8735);
nor U11446 (N_11446,N_9218,N_8358);
xnor U11447 (N_11447,N_9679,N_9487);
nor U11448 (N_11448,N_9803,N_9708);
nand U11449 (N_11449,N_8762,N_8650);
nand U11450 (N_11450,N_9450,N_8235);
xnor U11451 (N_11451,N_9053,N_9389);
nor U11452 (N_11452,N_9518,N_9927);
and U11453 (N_11453,N_9192,N_8578);
xor U11454 (N_11454,N_9476,N_8535);
nand U11455 (N_11455,N_9958,N_8797);
xor U11456 (N_11456,N_9465,N_8043);
or U11457 (N_11457,N_9275,N_8610);
nor U11458 (N_11458,N_9962,N_8792);
and U11459 (N_11459,N_9004,N_9249);
nand U11460 (N_11460,N_8424,N_9994);
or U11461 (N_11461,N_9390,N_9602);
nand U11462 (N_11462,N_8651,N_8768);
xnor U11463 (N_11463,N_8491,N_9038);
and U11464 (N_11464,N_8671,N_8779);
and U11465 (N_11465,N_9457,N_9423);
xor U11466 (N_11466,N_9541,N_8161);
nand U11467 (N_11467,N_8112,N_9335);
or U11468 (N_11468,N_9154,N_8956);
nand U11469 (N_11469,N_8152,N_8645);
nand U11470 (N_11470,N_9201,N_9797);
and U11471 (N_11471,N_8094,N_9363);
nand U11472 (N_11472,N_8716,N_9322);
and U11473 (N_11473,N_8692,N_8671);
and U11474 (N_11474,N_8585,N_8594);
or U11475 (N_11475,N_8848,N_9974);
and U11476 (N_11476,N_8777,N_9881);
nand U11477 (N_11477,N_9833,N_9887);
or U11478 (N_11478,N_8969,N_8515);
and U11479 (N_11479,N_9689,N_9283);
xor U11480 (N_11480,N_8408,N_8646);
and U11481 (N_11481,N_9971,N_8040);
or U11482 (N_11482,N_9939,N_8887);
and U11483 (N_11483,N_9121,N_8343);
nand U11484 (N_11484,N_8940,N_9323);
and U11485 (N_11485,N_9894,N_9879);
or U11486 (N_11486,N_9864,N_9625);
nor U11487 (N_11487,N_9667,N_8327);
nand U11488 (N_11488,N_8551,N_9554);
nand U11489 (N_11489,N_9841,N_9306);
nor U11490 (N_11490,N_9984,N_8283);
nor U11491 (N_11491,N_8057,N_8716);
or U11492 (N_11492,N_8469,N_8185);
xnor U11493 (N_11493,N_8880,N_8881);
or U11494 (N_11494,N_8848,N_9208);
nor U11495 (N_11495,N_8126,N_8887);
nand U11496 (N_11496,N_9223,N_8440);
nand U11497 (N_11497,N_8840,N_9556);
nand U11498 (N_11498,N_8330,N_9675);
or U11499 (N_11499,N_8681,N_9447);
nand U11500 (N_11500,N_9935,N_8230);
nor U11501 (N_11501,N_9355,N_8017);
or U11502 (N_11502,N_9997,N_9485);
xor U11503 (N_11503,N_8430,N_9916);
xor U11504 (N_11504,N_8497,N_8451);
or U11505 (N_11505,N_8887,N_8155);
and U11506 (N_11506,N_8663,N_8843);
nor U11507 (N_11507,N_8083,N_8150);
xnor U11508 (N_11508,N_8959,N_8163);
or U11509 (N_11509,N_9400,N_8422);
nor U11510 (N_11510,N_8199,N_9375);
nand U11511 (N_11511,N_8891,N_8241);
nor U11512 (N_11512,N_9230,N_9091);
xnor U11513 (N_11513,N_8583,N_8248);
and U11514 (N_11514,N_9743,N_8465);
or U11515 (N_11515,N_8957,N_9704);
nor U11516 (N_11516,N_9904,N_9300);
xnor U11517 (N_11517,N_8798,N_8251);
xor U11518 (N_11518,N_9128,N_8971);
or U11519 (N_11519,N_8317,N_9773);
and U11520 (N_11520,N_9463,N_9460);
xor U11521 (N_11521,N_9414,N_9274);
or U11522 (N_11522,N_9999,N_8184);
or U11523 (N_11523,N_8005,N_9795);
nand U11524 (N_11524,N_9368,N_8712);
nor U11525 (N_11525,N_8670,N_9105);
nand U11526 (N_11526,N_9116,N_9030);
or U11527 (N_11527,N_8200,N_9130);
or U11528 (N_11528,N_9119,N_8930);
nor U11529 (N_11529,N_9583,N_8174);
and U11530 (N_11530,N_9037,N_8902);
and U11531 (N_11531,N_8557,N_9069);
or U11532 (N_11532,N_8060,N_9741);
nor U11533 (N_11533,N_8024,N_8381);
nand U11534 (N_11534,N_9663,N_8944);
nand U11535 (N_11535,N_8610,N_8726);
nor U11536 (N_11536,N_9480,N_9482);
xnor U11537 (N_11537,N_8952,N_9712);
and U11538 (N_11538,N_8804,N_8891);
nand U11539 (N_11539,N_9433,N_8626);
and U11540 (N_11540,N_8425,N_9549);
nor U11541 (N_11541,N_9601,N_9932);
or U11542 (N_11542,N_8602,N_9819);
and U11543 (N_11543,N_8276,N_9600);
nor U11544 (N_11544,N_8950,N_9426);
and U11545 (N_11545,N_8988,N_9765);
nor U11546 (N_11546,N_8305,N_8248);
nand U11547 (N_11547,N_8301,N_8162);
nor U11548 (N_11548,N_9860,N_9231);
nor U11549 (N_11549,N_8959,N_9851);
and U11550 (N_11550,N_8664,N_9245);
and U11551 (N_11551,N_9054,N_8628);
nand U11552 (N_11552,N_9342,N_9053);
nor U11553 (N_11553,N_9099,N_8317);
and U11554 (N_11554,N_9806,N_9827);
or U11555 (N_11555,N_9231,N_9426);
and U11556 (N_11556,N_8026,N_9740);
xor U11557 (N_11557,N_9644,N_8870);
or U11558 (N_11558,N_8358,N_8980);
and U11559 (N_11559,N_8252,N_9235);
xnor U11560 (N_11560,N_8163,N_8228);
nor U11561 (N_11561,N_8561,N_8213);
or U11562 (N_11562,N_9500,N_8711);
or U11563 (N_11563,N_9659,N_9861);
nor U11564 (N_11564,N_9105,N_9517);
xor U11565 (N_11565,N_9076,N_9019);
and U11566 (N_11566,N_8260,N_9531);
xor U11567 (N_11567,N_9775,N_9920);
xor U11568 (N_11568,N_8864,N_9572);
nor U11569 (N_11569,N_9103,N_8737);
and U11570 (N_11570,N_9926,N_9346);
nor U11571 (N_11571,N_9023,N_9389);
xnor U11572 (N_11572,N_8385,N_8180);
nand U11573 (N_11573,N_8076,N_8642);
xor U11574 (N_11574,N_8605,N_9254);
xor U11575 (N_11575,N_8340,N_8107);
xor U11576 (N_11576,N_9412,N_8397);
and U11577 (N_11577,N_8440,N_9462);
nand U11578 (N_11578,N_8830,N_8857);
or U11579 (N_11579,N_8956,N_8665);
nor U11580 (N_11580,N_9728,N_9666);
or U11581 (N_11581,N_8560,N_8504);
nand U11582 (N_11582,N_8408,N_9340);
nand U11583 (N_11583,N_9468,N_8542);
or U11584 (N_11584,N_9986,N_8317);
or U11585 (N_11585,N_9442,N_8304);
nand U11586 (N_11586,N_9702,N_8822);
and U11587 (N_11587,N_9887,N_8116);
nor U11588 (N_11588,N_9306,N_9257);
nand U11589 (N_11589,N_9856,N_8252);
or U11590 (N_11590,N_9866,N_8015);
nor U11591 (N_11591,N_8095,N_8986);
nor U11592 (N_11592,N_8619,N_8173);
or U11593 (N_11593,N_8760,N_8293);
and U11594 (N_11594,N_9092,N_8548);
or U11595 (N_11595,N_9473,N_9540);
xnor U11596 (N_11596,N_8445,N_9693);
or U11597 (N_11597,N_9495,N_8833);
xnor U11598 (N_11598,N_9568,N_8672);
or U11599 (N_11599,N_8291,N_9886);
nor U11600 (N_11600,N_9727,N_9215);
nor U11601 (N_11601,N_8085,N_9081);
nand U11602 (N_11602,N_8029,N_8376);
nor U11603 (N_11603,N_8745,N_8703);
and U11604 (N_11604,N_9867,N_8598);
xor U11605 (N_11605,N_9768,N_8423);
or U11606 (N_11606,N_8642,N_8100);
nand U11607 (N_11607,N_9826,N_9878);
xor U11608 (N_11608,N_9978,N_9415);
and U11609 (N_11609,N_8318,N_8742);
or U11610 (N_11610,N_9854,N_8168);
nand U11611 (N_11611,N_8207,N_8202);
nand U11612 (N_11612,N_8685,N_8674);
and U11613 (N_11613,N_8172,N_9636);
xnor U11614 (N_11614,N_9897,N_8232);
xor U11615 (N_11615,N_8929,N_9382);
xor U11616 (N_11616,N_8300,N_8097);
nand U11617 (N_11617,N_9121,N_8161);
or U11618 (N_11618,N_8699,N_9439);
nor U11619 (N_11619,N_9466,N_9953);
nor U11620 (N_11620,N_9008,N_8393);
nand U11621 (N_11621,N_9763,N_9978);
nand U11622 (N_11622,N_9825,N_8011);
and U11623 (N_11623,N_9550,N_9477);
xnor U11624 (N_11624,N_8968,N_9025);
and U11625 (N_11625,N_9806,N_8377);
nand U11626 (N_11626,N_9976,N_9539);
nor U11627 (N_11627,N_8502,N_8554);
and U11628 (N_11628,N_9514,N_8170);
or U11629 (N_11629,N_9490,N_9347);
and U11630 (N_11630,N_9712,N_9640);
xnor U11631 (N_11631,N_8525,N_9325);
nor U11632 (N_11632,N_9570,N_9175);
nand U11633 (N_11633,N_9337,N_9626);
nor U11634 (N_11634,N_8940,N_8918);
nor U11635 (N_11635,N_9195,N_9055);
nor U11636 (N_11636,N_8175,N_8708);
nor U11637 (N_11637,N_8210,N_8641);
and U11638 (N_11638,N_9275,N_8285);
nand U11639 (N_11639,N_9653,N_8263);
xor U11640 (N_11640,N_9164,N_9323);
or U11641 (N_11641,N_8996,N_8971);
and U11642 (N_11642,N_8833,N_9480);
or U11643 (N_11643,N_9797,N_8996);
xor U11644 (N_11644,N_8696,N_9068);
or U11645 (N_11645,N_9103,N_8740);
or U11646 (N_11646,N_9310,N_8190);
and U11647 (N_11647,N_8550,N_9895);
xor U11648 (N_11648,N_8959,N_8084);
xor U11649 (N_11649,N_8303,N_8571);
nor U11650 (N_11650,N_9679,N_8255);
or U11651 (N_11651,N_9061,N_8410);
or U11652 (N_11652,N_8548,N_8657);
and U11653 (N_11653,N_9094,N_8166);
and U11654 (N_11654,N_8665,N_8077);
nand U11655 (N_11655,N_9390,N_9802);
or U11656 (N_11656,N_9556,N_9333);
and U11657 (N_11657,N_9936,N_8222);
xnor U11658 (N_11658,N_8229,N_8092);
xor U11659 (N_11659,N_9768,N_8441);
and U11660 (N_11660,N_8508,N_9699);
and U11661 (N_11661,N_9882,N_9787);
nand U11662 (N_11662,N_9480,N_8469);
or U11663 (N_11663,N_9441,N_9947);
or U11664 (N_11664,N_9400,N_9294);
xor U11665 (N_11665,N_8549,N_8312);
and U11666 (N_11666,N_8383,N_9928);
xnor U11667 (N_11667,N_8853,N_8692);
or U11668 (N_11668,N_9649,N_9507);
nor U11669 (N_11669,N_9992,N_9820);
or U11670 (N_11670,N_8103,N_9985);
nor U11671 (N_11671,N_9888,N_9087);
or U11672 (N_11672,N_9833,N_8584);
and U11673 (N_11673,N_8315,N_8352);
or U11674 (N_11674,N_8039,N_8654);
nand U11675 (N_11675,N_9929,N_9905);
nor U11676 (N_11676,N_9341,N_9316);
and U11677 (N_11677,N_9748,N_8990);
xnor U11678 (N_11678,N_9651,N_8947);
nand U11679 (N_11679,N_9874,N_8715);
or U11680 (N_11680,N_9776,N_9365);
nand U11681 (N_11681,N_8366,N_9304);
and U11682 (N_11682,N_9273,N_9042);
or U11683 (N_11683,N_9469,N_8249);
nand U11684 (N_11684,N_9054,N_8446);
or U11685 (N_11685,N_8213,N_9792);
xor U11686 (N_11686,N_9355,N_9494);
nand U11687 (N_11687,N_9707,N_9973);
nor U11688 (N_11688,N_9664,N_8271);
nor U11689 (N_11689,N_8160,N_9903);
xor U11690 (N_11690,N_9565,N_9442);
and U11691 (N_11691,N_9732,N_9806);
or U11692 (N_11692,N_8409,N_9781);
nand U11693 (N_11693,N_8099,N_8855);
nand U11694 (N_11694,N_9368,N_8709);
xnor U11695 (N_11695,N_9166,N_9485);
or U11696 (N_11696,N_8126,N_8832);
nor U11697 (N_11697,N_8233,N_8305);
and U11698 (N_11698,N_8638,N_8026);
nand U11699 (N_11699,N_8580,N_8065);
and U11700 (N_11700,N_9020,N_9921);
and U11701 (N_11701,N_8042,N_8376);
nor U11702 (N_11702,N_9493,N_8212);
xor U11703 (N_11703,N_8999,N_8780);
or U11704 (N_11704,N_9996,N_8294);
and U11705 (N_11705,N_8952,N_9913);
and U11706 (N_11706,N_8677,N_8975);
and U11707 (N_11707,N_8689,N_9457);
or U11708 (N_11708,N_8731,N_9917);
and U11709 (N_11709,N_9704,N_9661);
xor U11710 (N_11710,N_9574,N_9816);
or U11711 (N_11711,N_9139,N_9933);
nand U11712 (N_11712,N_8989,N_8091);
xnor U11713 (N_11713,N_8604,N_8626);
and U11714 (N_11714,N_9275,N_8062);
xor U11715 (N_11715,N_9921,N_9038);
or U11716 (N_11716,N_9350,N_8148);
or U11717 (N_11717,N_8761,N_8989);
or U11718 (N_11718,N_8972,N_8908);
nor U11719 (N_11719,N_8531,N_9762);
nor U11720 (N_11720,N_8384,N_8050);
nand U11721 (N_11721,N_8995,N_9977);
or U11722 (N_11722,N_8367,N_9535);
xor U11723 (N_11723,N_9889,N_9211);
or U11724 (N_11724,N_8323,N_8525);
xor U11725 (N_11725,N_9882,N_8907);
nand U11726 (N_11726,N_8356,N_8492);
nand U11727 (N_11727,N_8408,N_9452);
nor U11728 (N_11728,N_9321,N_8701);
nand U11729 (N_11729,N_8990,N_8743);
xnor U11730 (N_11730,N_9744,N_8593);
and U11731 (N_11731,N_8760,N_8415);
and U11732 (N_11732,N_9613,N_9538);
or U11733 (N_11733,N_8698,N_9541);
xnor U11734 (N_11734,N_9966,N_8211);
or U11735 (N_11735,N_8346,N_9526);
xor U11736 (N_11736,N_8907,N_8283);
nand U11737 (N_11737,N_9873,N_9921);
nor U11738 (N_11738,N_9795,N_9780);
nand U11739 (N_11739,N_8173,N_9003);
nand U11740 (N_11740,N_9530,N_8741);
and U11741 (N_11741,N_9207,N_8323);
nor U11742 (N_11742,N_9128,N_9746);
nor U11743 (N_11743,N_9100,N_8929);
and U11744 (N_11744,N_8565,N_8710);
and U11745 (N_11745,N_9556,N_9875);
xor U11746 (N_11746,N_8228,N_9748);
xnor U11747 (N_11747,N_8979,N_9457);
or U11748 (N_11748,N_8043,N_9747);
nor U11749 (N_11749,N_8517,N_9271);
xnor U11750 (N_11750,N_9979,N_9965);
nand U11751 (N_11751,N_9463,N_9805);
nand U11752 (N_11752,N_8847,N_9657);
or U11753 (N_11753,N_8736,N_9999);
xnor U11754 (N_11754,N_8318,N_8703);
xor U11755 (N_11755,N_9995,N_8833);
and U11756 (N_11756,N_8214,N_9976);
or U11757 (N_11757,N_9705,N_8840);
and U11758 (N_11758,N_8549,N_8275);
xnor U11759 (N_11759,N_8136,N_9072);
nor U11760 (N_11760,N_9994,N_9147);
nor U11761 (N_11761,N_9951,N_9621);
and U11762 (N_11762,N_9182,N_9063);
and U11763 (N_11763,N_8694,N_8264);
nor U11764 (N_11764,N_8562,N_9533);
or U11765 (N_11765,N_9830,N_8129);
nand U11766 (N_11766,N_8218,N_8486);
and U11767 (N_11767,N_9079,N_8890);
nand U11768 (N_11768,N_8361,N_9440);
nand U11769 (N_11769,N_9138,N_9488);
and U11770 (N_11770,N_9181,N_8378);
nor U11771 (N_11771,N_8160,N_8896);
or U11772 (N_11772,N_8381,N_8430);
xor U11773 (N_11773,N_8755,N_9328);
nand U11774 (N_11774,N_9356,N_9913);
and U11775 (N_11775,N_8582,N_8333);
nor U11776 (N_11776,N_9850,N_9241);
xnor U11777 (N_11777,N_8591,N_9475);
xnor U11778 (N_11778,N_9392,N_9369);
xnor U11779 (N_11779,N_8545,N_8613);
or U11780 (N_11780,N_9294,N_8855);
xnor U11781 (N_11781,N_8227,N_9141);
xnor U11782 (N_11782,N_9985,N_8389);
or U11783 (N_11783,N_8169,N_9061);
nor U11784 (N_11784,N_9443,N_8306);
nand U11785 (N_11785,N_8278,N_9565);
nor U11786 (N_11786,N_9087,N_8744);
and U11787 (N_11787,N_8996,N_9020);
or U11788 (N_11788,N_9184,N_9669);
nor U11789 (N_11789,N_9234,N_9933);
and U11790 (N_11790,N_9433,N_9213);
and U11791 (N_11791,N_8767,N_8139);
nand U11792 (N_11792,N_8697,N_8480);
or U11793 (N_11793,N_9978,N_9473);
nor U11794 (N_11794,N_9232,N_8870);
nand U11795 (N_11795,N_8675,N_9343);
nor U11796 (N_11796,N_8237,N_9591);
or U11797 (N_11797,N_8560,N_8605);
nand U11798 (N_11798,N_8050,N_8105);
xor U11799 (N_11799,N_9968,N_9272);
and U11800 (N_11800,N_9655,N_8765);
xnor U11801 (N_11801,N_9779,N_9745);
or U11802 (N_11802,N_9621,N_8713);
xor U11803 (N_11803,N_9001,N_8519);
xnor U11804 (N_11804,N_8570,N_8403);
or U11805 (N_11805,N_9092,N_8913);
nand U11806 (N_11806,N_8737,N_8885);
and U11807 (N_11807,N_8033,N_8732);
and U11808 (N_11808,N_9657,N_9406);
and U11809 (N_11809,N_9455,N_9430);
or U11810 (N_11810,N_8259,N_9653);
and U11811 (N_11811,N_8626,N_8671);
and U11812 (N_11812,N_9912,N_9863);
and U11813 (N_11813,N_8457,N_9592);
nor U11814 (N_11814,N_9030,N_9303);
and U11815 (N_11815,N_9549,N_8656);
nand U11816 (N_11816,N_8050,N_8984);
and U11817 (N_11817,N_8094,N_9349);
or U11818 (N_11818,N_8605,N_9287);
nor U11819 (N_11819,N_9219,N_8857);
xnor U11820 (N_11820,N_8980,N_8501);
xnor U11821 (N_11821,N_9279,N_9322);
nand U11822 (N_11822,N_8938,N_8906);
xnor U11823 (N_11823,N_8779,N_8538);
and U11824 (N_11824,N_9849,N_8588);
nand U11825 (N_11825,N_9621,N_8654);
and U11826 (N_11826,N_9025,N_9328);
xor U11827 (N_11827,N_8926,N_8826);
nand U11828 (N_11828,N_9519,N_8408);
nand U11829 (N_11829,N_9163,N_9717);
and U11830 (N_11830,N_9263,N_9752);
nor U11831 (N_11831,N_8103,N_9177);
and U11832 (N_11832,N_9117,N_9854);
nand U11833 (N_11833,N_9142,N_9793);
nor U11834 (N_11834,N_8696,N_9915);
xor U11835 (N_11835,N_9440,N_9725);
nor U11836 (N_11836,N_9644,N_8906);
nor U11837 (N_11837,N_9477,N_9213);
nand U11838 (N_11838,N_9194,N_8504);
nor U11839 (N_11839,N_9744,N_9108);
nor U11840 (N_11840,N_8302,N_9311);
or U11841 (N_11841,N_9291,N_8209);
and U11842 (N_11842,N_8455,N_8498);
or U11843 (N_11843,N_9574,N_8004);
xnor U11844 (N_11844,N_9818,N_8853);
xor U11845 (N_11845,N_9417,N_9995);
or U11846 (N_11846,N_8268,N_9681);
or U11847 (N_11847,N_8817,N_9976);
nand U11848 (N_11848,N_9657,N_9786);
or U11849 (N_11849,N_9207,N_8135);
xor U11850 (N_11850,N_8578,N_9152);
nand U11851 (N_11851,N_8975,N_8273);
nand U11852 (N_11852,N_8527,N_9882);
xor U11853 (N_11853,N_8608,N_8915);
nor U11854 (N_11854,N_9447,N_8918);
nor U11855 (N_11855,N_9923,N_9683);
xnor U11856 (N_11856,N_9178,N_9631);
or U11857 (N_11857,N_9997,N_8081);
xor U11858 (N_11858,N_8989,N_9630);
xor U11859 (N_11859,N_8602,N_8228);
xor U11860 (N_11860,N_9606,N_8600);
xnor U11861 (N_11861,N_8801,N_9897);
xnor U11862 (N_11862,N_9096,N_8463);
nand U11863 (N_11863,N_8650,N_8591);
nand U11864 (N_11864,N_8194,N_9124);
nor U11865 (N_11865,N_9004,N_9595);
and U11866 (N_11866,N_9296,N_9348);
xnor U11867 (N_11867,N_9566,N_8402);
nand U11868 (N_11868,N_8617,N_8871);
nor U11869 (N_11869,N_8802,N_8484);
or U11870 (N_11870,N_9500,N_8782);
and U11871 (N_11871,N_9738,N_8761);
or U11872 (N_11872,N_8580,N_8492);
or U11873 (N_11873,N_9375,N_8525);
xor U11874 (N_11874,N_9881,N_9309);
and U11875 (N_11875,N_9727,N_8516);
nor U11876 (N_11876,N_8848,N_9851);
xor U11877 (N_11877,N_8454,N_8967);
nand U11878 (N_11878,N_9197,N_9928);
xnor U11879 (N_11879,N_8651,N_9760);
or U11880 (N_11880,N_8546,N_8395);
or U11881 (N_11881,N_8877,N_8408);
and U11882 (N_11882,N_9989,N_9612);
or U11883 (N_11883,N_8849,N_8006);
or U11884 (N_11884,N_9342,N_8123);
nor U11885 (N_11885,N_8625,N_9607);
and U11886 (N_11886,N_9400,N_9851);
nand U11887 (N_11887,N_9401,N_8860);
or U11888 (N_11888,N_8179,N_9334);
nor U11889 (N_11889,N_8594,N_8226);
nand U11890 (N_11890,N_9942,N_9554);
and U11891 (N_11891,N_8017,N_9606);
and U11892 (N_11892,N_8962,N_9642);
xnor U11893 (N_11893,N_8731,N_9605);
nand U11894 (N_11894,N_9823,N_9831);
or U11895 (N_11895,N_8958,N_9057);
and U11896 (N_11896,N_8484,N_8934);
or U11897 (N_11897,N_9329,N_9104);
nand U11898 (N_11898,N_8776,N_8861);
nor U11899 (N_11899,N_9839,N_8613);
xor U11900 (N_11900,N_9903,N_8191);
xor U11901 (N_11901,N_9919,N_9543);
and U11902 (N_11902,N_9646,N_9991);
nor U11903 (N_11903,N_9876,N_8331);
or U11904 (N_11904,N_8396,N_8739);
nor U11905 (N_11905,N_8061,N_9211);
and U11906 (N_11906,N_9409,N_9636);
nand U11907 (N_11907,N_8562,N_9193);
and U11908 (N_11908,N_8760,N_8563);
nand U11909 (N_11909,N_8715,N_8962);
or U11910 (N_11910,N_9306,N_8512);
nand U11911 (N_11911,N_8494,N_9979);
and U11912 (N_11912,N_9900,N_8732);
xor U11913 (N_11913,N_8100,N_9027);
nand U11914 (N_11914,N_8357,N_9863);
or U11915 (N_11915,N_9837,N_9081);
and U11916 (N_11916,N_9840,N_8118);
xor U11917 (N_11917,N_9655,N_9331);
xor U11918 (N_11918,N_8387,N_8233);
and U11919 (N_11919,N_8852,N_9941);
or U11920 (N_11920,N_8681,N_8372);
nand U11921 (N_11921,N_8824,N_9163);
and U11922 (N_11922,N_9332,N_8398);
nor U11923 (N_11923,N_8213,N_9744);
nand U11924 (N_11924,N_8570,N_9225);
or U11925 (N_11925,N_8733,N_9920);
and U11926 (N_11926,N_8923,N_8700);
or U11927 (N_11927,N_8790,N_8429);
or U11928 (N_11928,N_9787,N_9804);
and U11929 (N_11929,N_9114,N_9908);
xor U11930 (N_11930,N_9654,N_9528);
or U11931 (N_11931,N_9365,N_8910);
nand U11932 (N_11932,N_8474,N_8886);
nand U11933 (N_11933,N_9448,N_8485);
nand U11934 (N_11934,N_8354,N_9771);
nand U11935 (N_11935,N_9962,N_8726);
and U11936 (N_11936,N_8358,N_9621);
nand U11937 (N_11937,N_9723,N_9480);
nand U11938 (N_11938,N_8878,N_9024);
or U11939 (N_11939,N_8402,N_9350);
and U11940 (N_11940,N_8884,N_8393);
nand U11941 (N_11941,N_9397,N_8488);
nand U11942 (N_11942,N_9774,N_9059);
nor U11943 (N_11943,N_9551,N_8652);
nor U11944 (N_11944,N_8282,N_9919);
and U11945 (N_11945,N_8422,N_9077);
nor U11946 (N_11946,N_9980,N_9808);
and U11947 (N_11947,N_9465,N_9522);
nand U11948 (N_11948,N_9068,N_9354);
or U11949 (N_11949,N_8179,N_9819);
xor U11950 (N_11950,N_9111,N_9510);
and U11951 (N_11951,N_9978,N_9496);
or U11952 (N_11952,N_9441,N_9882);
or U11953 (N_11953,N_8851,N_9068);
or U11954 (N_11954,N_8194,N_9260);
and U11955 (N_11955,N_9658,N_9948);
nand U11956 (N_11956,N_8616,N_9337);
nor U11957 (N_11957,N_9885,N_8033);
nand U11958 (N_11958,N_9946,N_8305);
nor U11959 (N_11959,N_8670,N_8916);
and U11960 (N_11960,N_8549,N_9734);
xnor U11961 (N_11961,N_8707,N_8668);
nand U11962 (N_11962,N_9276,N_8561);
and U11963 (N_11963,N_8761,N_9579);
nand U11964 (N_11964,N_8681,N_9991);
or U11965 (N_11965,N_8402,N_9429);
nand U11966 (N_11966,N_9944,N_8417);
xnor U11967 (N_11967,N_9553,N_9816);
xor U11968 (N_11968,N_9516,N_9437);
xnor U11969 (N_11969,N_9049,N_8252);
nor U11970 (N_11970,N_8393,N_9428);
and U11971 (N_11971,N_8730,N_8452);
nor U11972 (N_11972,N_9281,N_8680);
nor U11973 (N_11973,N_9313,N_9409);
nand U11974 (N_11974,N_9445,N_9771);
xor U11975 (N_11975,N_8898,N_8686);
or U11976 (N_11976,N_9505,N_9788);
nor U11977 (N_11977,N_8543,N_8370);
and U11978 (N_11978,N_9993,N_8832);
or U11979 (N_11979,N_8365,N_9562);
and U11980 (N_11980,N_8105,N_9672);
nor U11981 (N_11981,N_9750,N_9030);
xnor U11982 (N_11982,N_8535,N_8770);
nand U11983 (N_11983,N_8916,N_8441);
nand U11984 (N_11984,N_8511,N_9868);
nor U11985 (N_11985,N_9611,N_8385);
nand U11986 (N_11986,N_8887,N_8130);
nand U11987 (N_11987,N_9323,N_9500);
nor U11988 (N_11988,N_9214,N_8242);
nor U11989 (N_11989,N_8398,N_9645);
and U11990 (N_11990,N_9253,N_9674);
xor U11991 (N_11991,N_9965,N_8297);
xnor U11992 (N_11992,N_8908,N_9808);
or U11993 (N_11993,N_8640,N_8074);
nor U11994 (N_11994,N_9846,N_9647);
or U11995 (N_11995,N_8283,N_8340);
nor U11996 (N_11996,N_9615,N_8397);
nor U11997 (N_11997,N_8220,N_8763);
or U11998 (N_11998,N_8656,N_9473);
and U11999 (N_11999,N_9793,N_9346);
nor U12000 (N_12000,N_10392,N_10058);
xnor U12001 (N_12001,N_11283,N_10326);
or U12002 (N_12002,N_11812,N_10386);
xnor U12003 (N_12003,N_11734,N_10404);
nor U12004 (N_12004,N_11501,N_10249);
xnor U12005 (N_12005,N_10912,N_11519);
nor U12006 (N_12006,N_11621,N_11492);
and U12007 (N_12007,N_10821,N_10554);
nand U12008 (N_12008,N_10409,N_11825);
or U12009 (N_12009,N_10188,N_11919);
and U12010 (N_12010,N_11399,N_11182);
and U12011 (N_12011,N_10028,N_11290);
xnor U12012 (N_12012,N_11297,N_10921);
nor U12013 (N_12013,N_11231,N_10811);
or U12014 (N_12014,N_10783,N_10178);
and U12015 (N_12015,N_11292,N_10238);
xor U12016 (N_12016,N_11334,N_10705);
or U12017 (N_12017,N_11991,N_10573);
and U12018 (N_12018,N_10172,N_10299);
nand U12019 (N_12019,N_11324,N_11217);
or U12020 (N_12020,N_10544,N_11916);
xor U12021 (N_12021,N_10570,N_10946);
nor U12022 (N_12022,N_11474,N_10785);
and U12023 (N_12023,N_10070,N_10711);
and U12024 (N_12024,N_10190,N_11874);
and U12025 (N_12025,N_10723,N_10839);
and U12026 (N_12026,N_10750,N_11814);
and U12027 (N_12027,N_10248,N_11136);
nor U12028 (N_12028,N_11248,N_10482);
nor U12029 (N_12029,N_11244,N_10470);
xor U12030 (N_12030,N_11102,N_11711);
nand U12031 (N_12031,N_11934,N_11583);
or U12032 (N_12032,N_10904,N_10709);
or U12033 (N_12033,N_10804,N_10187);
nand U12034 (N_12034,N_11398,N_11932);
nand U12035 (N_12035,N_11296,N_11428);
nor U12036 (N_12036,N_11479,N_11571);
or U12037 (N_12037,N_10346,N_10211);
nand U12038 (N_12038,N_11420,N_11444);
and U12039 (N_12039,N_10976,N_11116);
xor U12040 (N_12040,N_11109,N_10356);
nand U12041 (N_12041,N_11277,N_10111);
xnor U12042 (N_12042,N_10651,N_10538);
xor U12043 (N_12043,N_11707,N_10893);
xnor U12044 (N_12044,N_10018,N_11467);
or U12045 (N_12045,N_11702,N_11122);
nor U12046 (N_12046,N_11772,N_11154);
nor U12047 (N_12047,N_10202,N_10982);
nor U12048 (N_12048,N_10144,N_11347);
nor U12049 (N_12049,N_11215,N_10714);
and U12050 (N_12050,N_10305,N_11715);
and U12051 (N_12051,N_10297,N_11352);
nor U12052 (N_12052,N_11885,N_10378);
and U12053 (N_12053,N_11038,N_10966);
and U12054 (N_12054,N_11658,N_10360);
nor U12055 (N_12055,N_10184,N_10294);
and U12056 (N_12056,N_10557,N_10933);
nand U12057 (N_12057,N_10826,N_10990);
and U12058 (N_12058,N_10043,N_11505);
nand U12059 (N_12059,N_11235,N_10510);
or U12060 (N_12060,N_11357,N_11859);
xor U12061 (N_12061,N_11729,N_11705);
nand U12062 (N_12062,N_10082,N_10108);
nor U12063 (N_12063,N_10436,N_10756);
nand U12064 (N_12064,N_10331,N_11411);
and U12065 (N_12065,N_11550,N_11644);
xnor U12066 (N_12066,N_10149,N_11521);
nand U12067 (N_12067,N_11737,N_10931);
nand U12068 (N_12068,N_11977,N_10948);
or U12069 (N_12069,N_10846,N_10063);
and U12070 (N_12070,N_11405,N_10799);
nand U12071 (N_12071,N_10423,N_10822);
and U12072 (N_12072,N_10340,N_11273);
or U12073 (N_12073,N_10408,N_11433);
nor U12074 (N_12074,N_10022,N_11745);
nand U12075 (N_12075,N_11738,N_11897);
or U12076 (N_12076,N_10730,N_11019);
or U12077 (N_12077,N_11686,N_11335);
and U12078 (N_12078,N_10926,N_10576);
and U12079 (N_12079,N_11969,N_10774);
nand U12080 (N_12080,N_11671,N_10000);
nor U12081 (N_12081,N_11599,N_11927);
and U12082 (N_12082,N_11093,N_11301);
and U12083 (N_12083,N_10629,N_10984);
nand U12084 (N_12084,N_11082,N_11889);
xor U12085 (N_12085,N_10319,N_10041);
or U12086 (N_12086,N_10498,N_10875);
xnor U12087 (N_12087,N_10377,N_10133);
xnor U12088 (N_12088,N_10692,N_11643);
xnor U12089 (N_12089,N_10825,N_11802);
and U12090 (N_12090,N_11875,N_11533);
nand U12091 (N_12091,N_11662,N_11960);
nand U12092 (N_12092,N_10306,N_10492);
or U12093 (N_12093,N_10139,N_11890);
or U12094 (N_12094,N_11508,N_10191);
xor U12095 (N_12095,N_11120,N_11060);
nand U12096 (N_12096,N_10488,N_11475);
nor U12097 (N_12097,N_11843,N_10770);
xnor U12098 (N_12098,N_10957,N_10769);
and U12099 (N_12099,N_11480,N_10527);
nand U12100 (N_12100,N_11194,N_11504);
nor U12101 (N_12101,N_10645,N_11684);
nand U12102 (N_12102,N_10707,N_11453);
nor U12103 (N_12103,N_11949,N_11080);
nand U12104 (N_12104,N_11333,N_11162);
or U12105 (N_12105,N_10517,N_11717);
nand U12106 (N_12106,N_11641,N_11003);
nand U12107 (N_12107,N_10633,N_11421);
nor U12108 (N_12108,N_11650,N_10228);
xor U12109 (N_12109,N_11085,N_11022);
xor U12110 (N_12110,N_10788,N_11225);
nand U12111 (N_12111,N_11213,N_10892);
nand U12112 (N_12112,N_11633,N_10585);
xnor U12113 (N_12113,N_10442,N_10214);
nor U12114 (N_12114,N_11664,N_11354);
and U12115 (N_12115,N_11037,N_10158);
nor U12116 (N_12116,N_10568,N_11951);
xor U12117 (N_12117,N_11337,N_11219);
and U12118 (N_12118,N_10480,N_11071);
nor U12119 (N_12119,N_11667,N_11973);
xnor U12120 (N_12120,N_11168,N_11013);
or U12121 (N_12121,N_10174,N_11941);
or U12122 (N_12122,N_11576,N_10417);
or U12123 (N_12123,N_11692,N_10981);
nand U12124 (N_12124,N_10474,N_11079);
xor U12125 (N_12125,N_11310,N_10900);
or U12126 (N_12126,N_10073,N_11557);
nor U12127 (N_12127,N_10422,N_11672);
nor U12128 (N_12128,N_11754,N_11130);
nor U12129 (N_12129,N_10901,N_10757);
xnor U12130 (N_12130,N_11285,N_10563);
and U12131 (N_12131,N_11952,N_10837);
nand U12132 (N_12132,N_11512,N_10192);
nor U12133 (N_12133,N_10885,N_11903);
xnor U12134 (N_12134,N_10850,N_10878);
xor U12135 (N_12135,N_10452,N_10704);
and U12136 (N_12136,N_10123,N_10213);
xnor U12137 (N_12137,N_10764,N_10273);
xor U12138 (N_12138,N_10592,N_11258);
or U12139 (N_12139,N_10676,N_10514);
or U12140 (N_12140,N_10153,N_11904);
xor U12141 (N_12141,N_10109,N_10464);
or U12142 (N_12142,N_10366,N_11156);
nor U12143 (N_12143,N_11778,N_11094);
and U12144 (N_12144,N_10141,N_10486);
nor U12145 (N_12145,N_11348,N_10848);
and U12146 (N_12146,N_10828,N_11000);
and U12147 (N_12147,N_10119,N_10795);
xnor U12148 (N_12148,N_11107,N_11493);
xor U12149 (N_12149,N_10674,N_10542);
nand U12150 (N_12150,N_11375,N_10503);
and U12151 (N_12151,N_10967,N_10530);
and U12152 (N_12152,N_10965,N_11978);
xor U12153 (N_12153,N_11514,N_10852);
xor U12154 (N_12154,N_10759,N_10155);
or U12155 (N_12155,N_11647,N_10565);
or U12156 (N_12156,N_10716,N_10260);
or U12157 (N_12157,N_10905,N_10719);
and U12158 (N_12158,N_11926,N_11098);
nand U12159 (N_12159,N_10708,N_10425);
or U12160 (N_12160,N_10148,N_11852);
and U12161 (N_12161,N_10620,N_10625);
nand U12162 (N_12162,N_10091,N_11468);
or U12163 (N_12163,N_10463,N_10194);
nand U12164 (N_12164,N_11770,N_11328);
xor U12165 (N_12165,N_11992,N_11575);
nand U12166 (N_12166,N_11842,N_10993);
nor U12167 (N_12167,N_11946,N_10044);
nand U12168 (N_12168,N_10333,N_10817);
nor U12169 (N_12169,N_11742,N_11645);
and U12170 (N_12170,N_11840,N_10964);
nand U12171 (N_12171,N_10956,N_10626);
nor U12172 (N_12172,N_10315,N_10135);
xnor U12173 (N_12173,N_10084,N_10874);
xnor U12174 (N_12174,N_11451,N_11968);
nand U12175 (N_12175,N_10721,N_10744);
xnor U12176 (N_12176,N_10021,N_11482);
and U12177 (N_12177,N_10601,N_10256);
or U12178 (N_12178,N_10023,N_11700);
nor U12179 (N_12179,N_11469,N_11881);
or U12180 (N_12180,N_11610,N_11697);
xnor U12181 (N_12181,N_10203,N_10546);
and U12182 (N_12182,N_11722,N_11477);
or U12183 (N_12183,N_11151,N_10451);
nand U12184 (N_12184,N_10383,N_11561);
nand U12185 (N_12185,N_10146,N_10327);
nor U12186 (N_12186,N_10102,N_11133);
nor U12187 (N_12187,N_11427,N_10307);
xor U12188 (N_12188,N_11864,N_11084);
and U12189 (N_12189,N_11732,N_11698);
nor U12190 (N_12190,N_10301,N_11432);
and U12191 (N_12191,N_10880,N_11322);
or U12192 (N_12192,N_10308,N_10994);
nand U12193 (N_12193,N_10624,N_11306);
xor U12194 (N_12194,N_11445,N_10748);
and U12195 (N_12195,N_11572,N_11422);
xnor U12196 (N_12196,N_10941,N_11955);
xor U12197 (N_12197,N_10801,N_10179);
nand U12198 (N_12198,N_10534,N_11905);
nor U12199 (N_12199,N_10450,N_11247);
and U12200 (N_12200,N_11876,N_11270);
and U12201 (N_12201,N_10466,N_10917);
or U12202 (N_12202,N_11254,N_10381);
and U12203 (N_12203,N_10370,N_10528);
and U12204 (N_12204,N_10531,N_11966);
nor U12205 (N_12205,N_11942,N_10782);
nand U12206 (N_12206,N_11661,N_11974);
and U12207 (N_12207,N_11090,N_11943);
or U12208 (N_12208,N_11499,N_11765);
or U12209 (N_12209,N_10746,N_11490);
or U12210 (N_12210,N_11636,N_11846);
xor U12211 (N_12211,N_11300,N_10648);
xnor U12212 (N_12212,N_10341,N_11253);
xnor U12213 (N_12213,N_10897,N_10802);
xnor U12214 (N_12214,N_10870,N_10653);
nor U12215 (N_12215,N_10898,N_10185);
nor U12216 (N_12216,N_11196,N_11025);
and U12217 (N_12217,N_10375,N_11574);
and U12218 (N_12218,N_10258,N_10889);
xor U12219 (N_12219,N_10142,N_10233);
nand U12220 (N_12220,N_10552,N_11497);
nand U12221 (N_12221,N_10296,N_11407);
nor U12222 (N_12222,N_10060,N_11586);
and U12223 (N_12223,N_11179,N_11712);
nor U12224 (N_12224,N_10357,N_10079);
xnor U12225 (N_12225,N_11332,N_10833);
and U12226 (N_12226,N_11272,N_11728);
nand U12227 (N_12227,N_10796,N_10540);
nor U12228 (N_12228,N_11439,N_10895);
nand U12229 (N_12229,N_10309,N_11114);
xor U12230 (N_12230,N_10664,N_11788);
xor U12231 (N_12231,N_11766,N_11169);
and U12232 (N_12232,N_10583,N_10220);
or U12233 (N_12233,N_10928,N_10145);
nor U12234 (N_12234,N_10270,N_10410);
and U12235 (N_12235,N_11269,N_11390);
or U12236 (N_12236,N_10362,N_11893);
xnor U12237 (N_12237,N_10686,N_11771);
xor U12238 (N_12238,N_10717,N_11900);
xor U12239 (N_12239,N_11240,N_10166);
or U12240 (N_12240,N_11791,N_11461);
nand U12241 (N_12241,N_11138,N_11148);
and U12242 (N_12242,N_10537,N_11930);
or U12243 (N_12243,N_10636,N_10975);
or U12244 (N_12244,N_10003,N_11057);
nand U12245 (N_12245,N_10382,N_11317);
nor U12246 (N_12246,N_11542,N_10535);
or U12247 (N_12247,N_11202,N_10872);
or U12248 (N_12248,N_10218,N_11232);
nand U12249 (N_12249,N_10558,N_10056);
nor U12250 (N_12250,N_10862,N_11146);
nand U12251 (N_12251,N_10891,N_11739);
and U12252 (N_12252,N_10186,N_10884);
and U12253 (N_12253,N_10886,N_10282);
nor U12254 (N_12254,N_10793,N_10835);
nand U12255 (N_12255,N_11438,N_11437);
or U12256 (N_12256,N_10476,N_11066);
or U12257 (N_12257,N_11687,N_11004);
nand U12258 (N_12258,N_10167,N_11537);
nor U12259 (N_12259,N_10103,N_11374);
nor U12260 (N_12260,N_10501,N_11033);
xnor U12261 (N_12261,N_11067,N_11007);
xor U12262 (N_12262,N_10467,N_11068);
and U12263 (N_12263,N_10691,N_11054);
and U12264 (N_12264,N_10016,N_10810);
or U12265 (N_12265,N_11673,N_11710);
xor U12266 (N_12266,N_11838,N_10311);
or U12267 (N_12267,N_10367,N_11668);
nand U12268 (N_12268,N_11425,N_10789);
nand U12269 (N_12269,N_11426,N_10246);
or U12270 (N_12270,N_11635,N_11837);
or U12271 (N_12271,N_10979,N_11279);
nand U12272 (N_12272,N_10665,N_10911);
xor U12273 (N_12273,N_11396,N_11089);
xnor U12274 (N_12274,N_11579,N_11544);
and U12275 (N_12275,N_11883,N_10318);
nor U12276 (N_12276,N_11431,N_11032);
nor U12277 (N_12277,N_10245,N_10210);
nor U12278 (N_12278,N_10768,N_11380);
nand U12279 (N_12279,N_10732,N_11549);
and U12280 (N_12280,N_11517,N_11450);
nand U12281 (N_12281,N_10280,N_10930);
and U12282 (N_12282,N_10193,N_11449);
nand U12283 (N_12283,N_10002,N_11793);
xor U12284 (N_12284,N_10779,N_11395);
and U12285 (N_12285,N_10143,N_11053);
and U12286 (N_12286,N_10513,N_10495);
and U12287 (N_12287,N_11170,N_10940);
and U12288 (N_12288,N_11956,N_10431);
nand U12289 (N_12289,N_10460,N_11563);
nor U12290 (N_12290,N_11373,N_10936);
xnor U12291 (N_12291,N_10758,N_11518);
nor U12292 (N_12292,N_11748,N_10794);
and U12293 (N_12293,N_11372,N_10472);
and U12294 (N_12294,N_11293,N_11597);
xor U12295 (N_12295,N_11062,N_11760);
nor U12296 (N_12296,N_11460,N_10803);
nor U12297 (N_12297,N_11180,N_11239);
nor U12298 (N_12298,N_11070,N_10078);
nor U12299 (N_12299,N_11377,N_11606);
xnor U12300 (N_12300,N_10398,N_11014);
and U12301 (N_12301,N_11529,N_11531);
or U12302 (N_12302,N_11847,N_10548);
nand U12303 (N_12303,N_10971,N_11304);
xor U12304 (N_12304,N_11783,N_10477);
and U12305 (N_12305,N_11161,N_11284);
and U12306 (N_12306,N_10639,N_11604);
or U12307 (N_12307,N_11158,N_11486);
or U12308 (N_12308,N_11631,N_10961);
xnor U12309 (N_12309,N_10688,N_11391);
nor U12310 (N_12310,N_10883,N_10800);
or U12311 (N_12311,N_10418,N_11654);
nand U12312 (N_12312,N_11657,N_11602);
and U12313 (N_12313,N_11255,N_10300);
nor U12314 (N_12314,N_11491,N_10443);
or U12315 (N_12315,N_11371,N_11267);
nor U12316 (N_12316,N_11435,N_11790);
nor U12317 (N_12317,N_10832,N_10095);
or U12318 (N_12318,N_10606,N_10485);
or U12319 (N_12319,N_10916,N_10599);
nand U12320 (N_12320,N_10253,N_11524);
xor U12321 (N_12321,N_11902,N_11002);
and U12322 (N_12322,N_11500,N_10494);
or U12323 (N_12323,N_10168,N_10903);
and U12324 (N_12324,N_11118,N_11857);
xnor U12325 (N_12325,N_10286,N_10879);
nand U12326 (N_12326,N_10973,N_11556);
nor U12327 (N_12327,N_10608,N_11470);
nor U12328 (N_12328,N_11674,N_11489);
nor U12329 (N_12329,N_11096,N_11249);
xor U12330 (N_12330,N_11315,N_10247);
and U12331 (N_12331,N_10662,N_10271);
and U12332 (N_12332,N_11237,N_10824);
nand U12333 (N_12333,N_11861,N_11222);
and U12334 (N_12334,N_11029,N_11796);
nand U12335 (N_12335,N_11963,N_10695);
nor U12336 (N_12336,N_11620,N_10702);
nor U12337 (N_12337,N_10350,N_10937);
xor U12338 (N_12338,N_11323,N_11869);
nor U12339 (N_12339,N_11743,N_11099);
nand U12340 (N_12340,N_11005,N_11069);
xnor U12341 (N_12341,N_11034,N_11757);
xnor U12342 (N_12342,N_10014,N_11221);
or U12343 (N_12343,N_10983,N_10180);
nor U12344 (N_12344,N_10575,N_11965);
or U12345 (N_12345,N_11849,N_10181);
nor U12346 (N_12346,N_11774,N_10727);
nor U12347 (N_12347,N_11740,N_11077);
nor U12348 (N_12348,N_10814,N_11924);
nand U12349 (N_12349,N_11534,N_10943);
or U12350 (N_12350,N_10533,N_10128);
nand U12351 (N_12351,N_10605,N_10808);
nor U12352 (N_12352,N_11195,N_11211);
or U12353 (N_12353,N_11850,N_11844);
nor U12354 (N_12354,N_10678,N_11649);
nand U12355 (N_12355,N_10703,N_11696);
nor U12356 (N_12356,N_10150,N_11481);
or U12357 (N_12357,N_10330,N_11271);
nand U12358 (N_12358,N_11286,N_10087);
nor U12359 (N_12359,N_10493,N_11115);
or U12360 (N_12360,N_11685,N_11185);
nand U12361 (N_12361,N_10856,N_10959);
and U12362 (N_12362,N_11527,N_10197);
nor U12363 (N_12363,N_11828,N_10419);
or U12364 (N_12364,N_11839,N_10121);
nor U12365 (N_12365,N_11860,N_11820);
nor U12366 (N_12366,N_11807,N_11629);
or U12367 (N_12367,N_10038,N_11353);
nand U12368 (N_12368,N_11464,N_11389);
and U12369 (N_12369,N_10813,N_11016);
and U12370 (N_12370,N_11873,N_11088);
or U12371 (N_12371,N_10524,N_10266);
and U12372 (N_12372,N_11565,N_11953);
nand U12373 (N_12373,N_11018,N_11152);
or U12374 (N_12374,N_11896,N_10454);
nor U12375 (N_12375,N_11733,N_10868);
nand U12376 (N_12376,N_11199,N_10577);
xnor U12377 (N_12377,N_10734,N_11935);
nor U12378 (N_12378,N_10390,N_10644);
xnor U12379 (N_12379,N_11513,N_10596);
and U12380 (N_12380,N_11782,N_11201);
or U12381 (N_12381,N_11815,N_10314);
xnor U12382 (N_12382,N_11063,N_11403);
and U12383 (N_12383,N_10332,N_11746);
xnor U12384 (N_12384,N_10522,N_10407);
xnor U12385 (N_12385,N_11823,N_11419);
or U12386 (N_12386,N_10484,N_11208);
xor U12387 (N_12387,N_11494,N_11176);
nand U12388 (N_12388,N_11383,N_11679);
nand U12389 (N_12389,N_11150,N_10337);
and U12390 (N_12390,N_10999,N_11472);
or U12391 (N_12391,N_10434,N_10863);
xor U12392 (N_12392,N_10622,N_11725);
nor U12393 (N_12393,N_11612,N_10265);
nand U12394 (N_12394,N_10015,N_11910);
xor U12395 (N_12395,N_11141,N_11637);
and U12396 (N_12396,N_11412,N_10209);
or U12397 (N_12397,N_10469,N_10176);
nand U12398 (N_12398,N_11064,N_11659);
xnor U12399 (N_12399,N_11212,N_11496);
or U12400 (N_12400,N_11980,N_10208);
xnor U12401 (N_12401,N_11547,N_10361);
nand U12402 (N_12402,N_10458,N_11205);
nand U12403 (N_12403,N_10061,N_11749);
nand U12404 (N_12404,N_10076,N_11305);
nand U12405 (N_12405,N_11149,N_10051);
xor U12406 (N_12406,N_10499,N_11806);
xor U12407 (N_12407,N_10384,N_10138);
nor U12408 (N_12408,N_11360,N_10385);
xor U12409 (N_12409,N_11994,N_11075);
and U12410 (N_12410,N_11785,N_10853);
and U12411 (N_12411,N_11552,N_10212);
nand U12412 (N_12412,N_10175,N_11670);
and U12413 (N_12413,N_11799,N_10798);
and U12414 (N_12414,N_11350,N_10843);
and U12415 (N_12415,N_11727,N_11609);
nor U12416 (N_12416,N_11442,N_11804);
nor U12417 (N_12417,N_11607,N_11404);
and U12418 (N_12418,N_10547,N_11520);
nor U12419 (N_12419,N_10525,N_11471);
nor U12420 (N_12420,N_10706,N_10840);
nand U12421 (N_12421,N_10304,N_11140);
or U12422 (N_12422,N_11726,N_11701);
nand U12423 (N_12423,N_10553,N_11920);
nor U12424 (N_12424,N_10784,N_10630);
xnor U12425 (N_12425,N_11632,N_11625);
or U12426 (N_12426,N_11566,N_11441);
nand U12427 (N_12427,N_10427,N_10012);
xnor U12428 (N_12428,N_10338,N_10355);
nor U12429 (N_12429,N_10026,N_11081);
nor U12430 (N_12430,N_11867,N_10506);
nor U12431 (N_12431,N_10440,N_11095);
or U12432 (N_12432,N_11540,N_10963);
nand U12433 (N_12433,N_10675,N_10389);
xnor U12434 (N_12434,N_11393,N_10710);
nand U12435 (N_12435,N_11921,N_10353);
or U12436 (N_12436,N_11776,N_11144);
or U12437 (N_12437,N_10215,N_11358);
and U12438 (N_12438,N_11238,N_10640);
and U12439 (N_12439,N_10559,N_11250);
and U12440 (N_12440,N_10643,N_11648);
nand U12441 (N_12441,N_11059,N_11307);
xnor U12442 (N_12442,N_11626,N_10037);
or U12443 (N_12443,N_11593,N_11683);
xor U12444 (N_12444,N_11397,N_11406);
xnor U12445 (N_12445,N_11767,N_11724);
or U12446 (N_12446,N_11261,N_11826);
xor U12447 (N_12447,N_10590,N_11264);
nor U12448 (N_12448,N_11040,N_11555);
nand U12449 (N_12449,N_11265,N_10114);
and U12450 (N_12450,N_11756,N_11908);
nand U12451 (N_12451,N_11209,N_11452);
nor U12452 (N_12452,N_11015,N_10876);
xnor U12453 (N_12453,N_10754,N_10086);
xnor U12454 (N_12454,N_10790,N_11694);
and U12455 (N_12455,N_10171,N_11065);
xnor U12456 (N_12456,N_11017,N_11567);
nor U12457 (N_12457,N_11339,N_11362);
nor U12458 (N_12458,N_10614,N_10251);
and U12459 (N_12459,N_10068,N_10050);
and U12460 (N_12460,N_11311,N_11947);
xnor U12461 (N_12461,N_10683,N_11361);
nand U12462 (N_12462,N_11230,N_11190);
and U12463 (N_12463,N_11971,N_11171);
nand U12464 (N_12464,N_11041,N_10055);
nor U12465 (N_12465,N_10767,N_10036);
and U12466 (N_12466,N_10731,N_10761);
nand U12467 (N_12467,N_10433,N_10687);
or U12468 (N_12468,N_11506,N_11074);
and U12469 (N_12469,N_10229,N_11553);
nor U12470 (N_12470,N_11266,N_10487);
xnor U12471 (N_12471,N_11695,N_10083);
and U12472 (N_12472,N_10955,N_11618);
nand U12473 (N_12473,N_10272,N_10523);
xor U12474 (N_12474,N_10267,N_10371);
or U12475 (N_12475,N_10312,N_11268);
nand U12476 (N_12476,N_10752,N_11937);
xnor U12477 (N_12477,N_11559,N_10742);
nand U12478 (N_12478,N_11851,N_11367);
xnor U12479 (N_12479,N_10255,N_11024);
nand U12480 (N_12480,N_10243,N_11026);
xnor U12481 (N_12481,N_10298,N_10765);
nand U12482 (N_12482,N_10910,N_11758);
nand U12483 (N_12483,N_11502,N_10236);
and U12484 (N_12484,N_11928,N_10697);
xnor U12485 (N_12485,N_10887,N_11925);
and U12486 (N_12486,N_11186,N_10762);
nand U12487 (N_12487,N_11343,N_10222);
nand U12488 (N_12488,N_11582,N_10399);
nand U12489 (N_12489,N_11011,N_10749);
and U12490 (N_12490,N_11137,N_11871);
and U12491 (N_12491,N_11294,N_10257);
and U12492 (N_12492,N_11379,N_11164);
nor U12493 (N_12493,N_10908,N_11630);
and U12494 (N_12494,N_10649,N_10654);
or U12495 (N_12495,N_11689,N_10421);
or U12496 (N_12496,N_11172,N_11365);
nand U12497 (N_12497,N_10725,N_11251);
and U12498 (N_12498,N_10402,N_10646);
or U12499 (N_12499,N_10230,N_11892);
xor U12500 (N_12500,N_10773,N_11759);
nand U12501 (N_12501,N_11462,N_11564);
nor U12502 (N_12502,N_11291,N_11591);
and U12503 (N_12503,N_10741,N_11351);
nor U12504 (N_12504,N_10225,N_11988);
and U12505 (N_12505,N_10323,N_10631);
xnor U12506 (N_12506,N_11507,N_10806);
and U12507 (N_12507,N_10694,N_10029);
or U12508 (N_12508,N_11510,N_10574);
nor U12509 (N_12509,N_11006,N_10099);
and U12510 (N_12510,N_11001,N_11933);
or U12511 (N_12511,N_10254,N_10584);
nand U12512 (N_12512,N_10269,N_10865);
or U12513 (N_12513,N_11344,N_11111);
nor U12514 (N_12514,N_11680,N_10924);
and U12515 (N_12515,N_10320,N_11123);
nand U12516 (N_12516,N_10632,N_10600);
xor U12517 (N_12517,N_10566,N_11278);
and U12518 (N_12518,N_10455,N_11055);
nand U12519 (N_12519,N_11012,N_11931);
nor U12520 (N_12520,N_11259,N_10935);
and U12521 (N_12521,N_11833,N_11713);
nor U12522 (N_12522,N_10560,N_10809);
and U12523 (N_12523,N_10521,N_11459);
nor U12524 (N_12524,N_10010,N_10032);
or U12525 (N_12525,N_10290,N_10403);
nand U12526 (N_12526,N_10588,N_10475);
nand U12527 (N_12527,N_11327,N_10446);
nand U12528 (N_12528,N_11803,N_10200);
or U12529 (N_12529,N_10855,N_10080);
nor U12530 (N_12530,N_11720,N_10339);
nand U12531 (N_12531,N_11652,N_10722);
or U12532 (N_12532,N_11856,N_10745);
and U12533 (N_12533,N_10395,N_10618);
and U12534 (N_12534,N_11157,N_10827);
nand U12535 (N_12535,N_11299,N_10124);
and U12536 (N_12536,N_11418,N_10988);
or U12537 (N_12537,N_10445,N_11967);
xnor U12538 (N_12538,N_11982,N_11175);
or U12539 (N_12539,N_10130,N_10169);
xor U12540 (N_12540,N_11210,N_11792);
and U12541 (N_12541,N_11402,N_10815);
or U12542 (N_12542,N_10031,N_10536);
or U12543 (N_12543,N_11976,N_11447);
and U12544 (N_12544,N_10516,N_11303);
nand U12545 (N_12545,N_10595,N_10638);
nand U12546 (N_12546,N_10945,N_11789);
nand U12547 (N_12547,N_11309,N_10343);
nand U12548 (N_12548,N_10259,N_10094);
nor U12549 (N_12549,N_10689,N_11800);
and U12550 (N_12550,N_11797,N_10163);
or U12551 (N_12551,N_10310,N_10604);
nand U12552 (N_12552,N_10344,N_10771);
nor U12553 (N_12553,N_11049,N_11045);
nand U12554 (N_12554,N_11901,N_11203);
xnor U12555 (N_12555,N_10581,N_10738);
or U12556 (N_12556,N_10066,N_11539);
and U12557 (N_12557,N_10968,N_10615);
and U12558 (N_12558,N_11048,N_11458);
or U12559 (N_12559,N_10223,N_10405);
xnor U12560 (N_12560,N_11975,N_11047);
xor U12561 (N_12561,N_10008,N_10117);
xor U12562 (N_12562,N_10529,N_10195);
xnor U12563 (N_12563,N_10578,N_10406);
or U12564 (N_12564,N_11424,N_10033);
and U12565 (N_12565,N_10668,N_11312);
nor U12566 (N_12566,N_10962,N_10349);
xnor U12567 (N_12567,N_10561,N_10989);
nand U12568 (N_12568,N_10562,N_11275);
nor U12569 (N_12569,N_11087,N_11415);
xor U12570 (N_12570,N_11204,N_10030);
xor U12571 (N_12571,N_11821,N_10471);
xor U12572 (N_12572,N_11723,N_10942);
nor U12573 (N_12573,N_10132,N_10364);
or U12574 (N_12574,N_11560,N_10849);
xnor U12575 (N_12575,N_10241,N_11824);
or U12576 (N_12576,N_10125,N_11200);
nand U12577 (N_12577,N_10657,N_11370);
or U12578 (N_12578,N_10077,N_10116);
or U12579 (N_12579,N_11699,N_11817);
nand U12580 (N_12580,N_10579,N_11972);
or U12581 (N_12581,N_10439,N_11541);
nand U12582 (N_12582,N_11108,N_10551);
and U12583 (N_12583,N_11886,N_11198);
or U12584 (N_12584,N_11962,N_11573);
or U12585 (N_12585,N_10156,N_10217);
and U12586 (N_12586,N_10923,N_10635);
and U12587 (N_12587,N_11936,N_10567);
or U12588 (N_12588,N_11061,N_11781);
and U12589 (N_12589,N_10660,N_11718);
and U12590 (N_12590,N_10572,N_11155);
or U12591 (N_12591,N_11483,N_10894);
or U12592 (N_12592,N_10420,N_11242);
or U12593 (N_12593,N_10847,N_10221);
and U12594 (N_12594,N_11236,N_10004);
and U12595 (N_12595,N_11126,N_10733);
nand U12596 (N_12596,N_11139,N_10348);
or U12597 (N_12597,N_11605,N_10953);
nand U12598 (N_12598,N_11127,N_11214);
or U12599 (N_12599,N_11245,N_11944);
and U12600 (N_12600,N_10747,N_11484);
or U12601 (N_12601,N_10831,N_10262);
xnor U12602 (N_12602,N_10224,N_10609);
nand U12603 (N_12603,N_10869,N_10667);
xnor U12604 (N_12604,N_10518,N_10610);
and U12605 (N_12605,N_10035,N_11256);
or U12606 (N_12606,N_11744,N_10104);
nor U12607 (N_12607,N_10650,N_11669);
or U12608 (N_12608,N_11117,N_10679);
or U12609 (N_12609,N_10661,N_10619);
nor U12610 (N_12610,N_10177,N_11302);
or U12611 (N_12611,N_10556,N_10415);
and U12612 (N_12612,N_11342,N_11809);
and U12613 (N_12613,N_11979,N_11721);
nor U12614 (N_12614,N_11603,N_11855);
nand U12615 (N_12615,N_10995,N_10183);
nor U12616 (N_12616,N_10845,N_11870);
and U12617 (N_12617,N_11808,N_10069);
or U12618 (N_12618,N_11206,N_11434);
xor U12619 (N_12619,N_11193,N_10666);
xnor U12620 (N_12620,N_11958,N_11289);
nand U12621 (N_12621,N_10064,N_10696);
and U12622 (N_12622,N_11142,N_11858);
xnor U12623 (N_12623,N_11105,N_11429);
and U12624 (N_12624,N_11388,N_10411);
or U12625 (N_12625,N_11097,N_10020);
nor U12626 (N_12626,N_10718,N_10275);
nand U12627 (N_12627,N_11923,N_11640);
or U12628 (N_12628,N_11455,N_11887);
xor U12629 (N_12629,N_11811,N_11135);
and U12630 (N_12630,N_11592,N_11188);
or U12631 (N_12631,N_11865,N_10641);
xnor U12632 (N_12632,N_10818,N_11030);
or U12633 (N_12633,N_10751,N_10478);
or U12634 (N_12634,N_11655,N_11341);
nand U12635 (N_12635,N_10866,N_10805);
or U12636 (N_12636,N_11627,N_11110);
or U12637 (N_12637,N_11646,N_10755);
xnor U12638 (N_12638,N_10059,N_11189);
and U12639 (N_12639,N_11569,N_11691);
or U12640 (N_12640,N_10712,N_11862);
or U12641 (N_12641,N_10157,N_11243);
nand U12642 (N_12642,N_10047,N_11587);
xnor U12643 (N_12643,N_11394,N_10226);
or U12644 (N_12644,N_11446,N_10491);
xnor U12645 (N_12645,N_11316,N_11463);
or U12646 (N_12646,N_11708,N_11987);
and U12647 (N_12647,N_11877,N_11914);
nor U12648 (N_12648,N_10938,N_11101);
nand U12649 (N_12649,N_11308,N_11031);
xor U12650 (N_12650,N_10429,N_11915);
nor U12651 (N_12651,N_11511,N_11709);
xnor U12652 (N_12652,N_10992,N_10159);
nor U12653 (N_12653,N_10792,N_10096);
or U12654 (N_12654,N_10511,N_11638);
nor U12655 (N_12655,N_10656,N_10416);
xor U12656 (N_12656,N_10274,N_10854);
nor U12657 (N_12657,N_11939,N_10013);
xnor U12658 (N_12658,N_10873,N_11703);
nand U12659 (N_12659,N_11509,N_10359);
and U12660 (N_12660,N_11872,N_11895);
and U12661 (N_12661,N_10283,N_11836);
nor U12662 (N_12662,N_10118,N_11145);
nor U12663 (N_12663,N_11369,N_10081);
or U12664 (N_12664,N_11046,N_10877);
nor U12665 (N_12665,N_11515,N_11546);
or U12666 (N_12666,N_11121,N_10261);
and U12667 (N_12667,N_10907,N_10424);
nand U12668 (N_12668,N_11167,N_10432);
or U12669 (N_12669,N_10512,N_11829);
and U12670 (N_12670,N_11665,N_11381);
nand U12671 (N_12671,N_11220,N_10685);
or U12672 (N_12672,N_10669,N_10034);
xnor U12673 (N_12673,N_11366,N_11409);
xnor U12674 (N_12674,N_10196,N_11819);
xnor U12675 (N_12675,N_11010,N_10160);
or U12676 (N_12676,N_10006,N_10001);
nand U12677 (N_12677,N_11356,N_11634);
xor U12678 (N_12678,N_10915,N_10461);
and U12679 (N_12679,N_10302,N_10670);
nor U12680 (N_12680,N_10658,N_10607);
nand U12681 (N_12681,N_11401,N_10227);
xnor U12682 (N_12682,N_11642,N_11577);
xor U12683 (N_12683,N_11854,N_10954);
and U12684 (N_12684,N_10673,N_11948);
nand U12685 (N_12685,N_10115,N_11106);
or U12686 (N_12686,N_11473,N_10541);
xnor U12687 (N_12687,N_11677,N_11052);
or U12688 (N_12688,N_11349,N_10781);
or U12689 (N_12689,N_10264,N_10284);
and U12690 (N_12690,N_11617,N_11585);
xnor U12691 (N_12691,N_11083,N_11174);
nor U12692 (N_12692,N_11990,N_10334);
nand U12693 (N_12693,N_11794,N_10199);
xor U12694 (N_12694,N_10019,N_11218);
and U12695 (N_12695,N_11173,N_10182);
xor U12696 (N_12696,N_11009,N_10829);
xnor U12697 (N_12697,N_10374,N_10090);
or U12698 (N_12698,N_11751,N_10690);
xnor U12699 (N_12699,N_10396,N_10925);
or U12700 (N_12700,N_10154,N_11227);
nor U12701 (N_12701,N_11961,N_10515);
nor U12702 (N_12702,N_10890,N_11690);
nor U12703 (N_12703,N_11954,N_10391);
and U12704 (N_12704,N_11246,N_11735);
or U12705 (N_12705,N_11112,N_10603);
xnor U12706 (N_12706,N_11535,N_10007);
xor U12707 (N_12707,N_11551,N_10039);
nand U12708 (N_12708,N_11448,N_10198);
xor U12709 (N_12709,N_11523,N_10295);
or U12710 (N_12710,N_10902,N_11779);
and U12711 (N_12711,N_11187,N_10067);
xnor U12712 (N_12712,N_11197,N_11233);
nor U12713 (N_12713,N_10071,N_10325);
and U12714 (N_12714,N_11543,N_11023);
or U12715 (N_12715,N_11938,N_11827);
xor U12716 (N_12716,N_11950,N_10441);
nor U12717 (N_12717,N_10888,N_10483);
or U12718 (N_12718,N_10376,N_10586);
nand U12719 (N_12719,N_11613,N_10239);
xnor U12720 (N_12720,N_11346,N_10140);
xnor U12721 (N_12721,N_11408,N_11813);
nand U12722 (N_12722,N_10715,N_10947);
xnor U12723 (N_12723,N_11378,N_11922);
nor U12724 (N_12724,N_10763,N_10369);
xor U12725 (N_12725,N_10834,N_10278);
and U12726 (N_12726,N_10207,N_10958);
nor U12727 (N_12727,N_11898,N_11651);
and U12728 (N_12728,N_10465,N_11340);
and U12729 (N_12729,N_11020,N_11736);
xnor U12730 (N_12730,N_10293,N_10438);
and U12731 (N_12731,N_11706,N_10120);
nor U12732 (N_12732,N_10092,N_11485);
xnor U12733 (N_12733,N_10352,N_11775);
and U12734 (N_12734,N_11675,N_11879);
and U12735 (N_12735,N_10819,N_11787);
nand U12736 (N_12736,N_10372,N_10980);
nor U12737 (N_12737,N_10602,N_11436);
nand U12738 (N_12738,N_11282,N_11623);
xor U12739 (N_12739,N_10448,N_11364);
nor U12740 (N_12740,N_10634,N_11440);
nand U12741 (N_12741,N_10652,N_11410);
xor U12742 (N_12742,N_10234,N_10899);
xor U12743 (N_12743,N_10049,N_10354);
or U12744 (N_12744,N_10113,N_11073);
nor U12745 (N_12745,N_11338,N_11124);
nand U12746 (N_12746,N_11413,N_10786);
xor U12747 (N_12747,N_10950,N_11624);
or U12748 (N_12748,N_11676,N_11681);
or U12749 (N_12749,N_11795,N_10131);
nand U12750 (N_12750,N_11318,N_11092);
nand U12751 (N_12751,N_11260,N_10373);
or U12752 (N_12752,N_10838,N_10881);
or U12753 (N_12753,N_10776,N_10072);
xor U12754 (N_12754,N_11805,N_10740);
or U12755 (N_12755,N_10571,N_11042);
nand U12756 (N_12756,N_10288,N_10457);
and U12757 (N_12757,N_10136,N_11545);
and U12758 (N_12758,N_10122,N_10743);
or U12759 (N_12759,N_11050,N_11747);
nor U12760 (N_12760,N_10281,N_10127);
and U12761 (N_12761,N_10914,N_11753);
nand U12762 (N_12762,N_10151,N_11276);
or U12763 (N_12763,N_10841,N_10587);
nand U12764 (N_12764,N_10336,N_10739);
nand U12765 (N_12765,N_10098,N_10412);
nand U12766 (N_12766,N_10428,N_10085);
xor U12767 (N_12767,N_10042,N_11750);
nand U12768 (N_12768,N_10520,N_10321);
and U12769 (N_12769,N_11104,N_11964);
and U12770 (N_12770,N_10394,N_11044);
or U12771 (N_12771,N_11207,N_11336);
or U12772 (N_12772,N_11538,N_10502);
nor U12773 (N_12773,N_11688,N_11568);
xnor U12774 (N_12774,N_10927,N_10864);
and U12775 (N_12775,N_10949,N_10393);
xnor U12776 (N_12776,N_10414,N_11730);
xor U12777 (N_12777,N_10045,N_10093);
and U12778 (N_12778,N_11848,N_10985);
nor U12779 (N_12779,N_10075,N_10462);
nand U12780 (N_12780,N_11768,N_10997);
or U12781 (N_12781,N_11280,N_10351);
xor U12782 (N_12782,N_10324,N_10387);
nand U12783 (N_12783,N_11263,N_10137);
and U12784 (N_12784,N_10589,N_10097);
nor U12785 (N_12785,N_10054,N_10240);
nor U12786 (N_12786,N_11588,N_11581);
nor U12787 (N_12787,N_11595,N_10972);
and U12788 (N_12788,N_11345,N_10244);
nor U12789 (N_12789,N_11611,N_10713);
or U12790 (N_12790,N_10939,N_11021);
nor U12791 (N_12791,N_10857,N_11834);
nand U12792 (N_12792,N_11035,N_11100);
nor U12793 (N_12793,N_11329,N_11131);
and U12794 (N_12794,N_11769,N_11252);
xor U12795 (N_12795,N_10555,N_11376);
and U12796 (N_12796,N_11443,N_10677);
xnor U12797 (N_12797,N_10048,N_10292);
or U12798 (N_12798,N_11241,N_11229);
nor U12799 (N_12799,N_11298,N_11830);
nor U12800 (N_12800,N_11907,N_11129);
nand U12801 (N_12801,N_10046,N_10164);
or U12802 (N_12802,N_11616,N_10564);
nand U12803 (N_12803,N_11132,N_10504);
nor U12804 (N_12804,N_11147,N_11989);
or U12805 (N_12805,N_11355,N_11880);
and U12806 (N_12806,N_10126,N_11091);
or U12807 (N_12807,N_10642,N_11183);
nand U12808 (N_12808,N_11125,N_10736);
nor U12809 (N_12809,N_10909,N_10929);
nor U12810 (N_12810,N_11622,N_10289);
and U12811 (N_12811,N_11414,N_10582);
or U12812 (N_12812,N_10112,N_10011);
nor U12813 (N_12813,N_11798,N_10617);
xor U12814 (N_12814,N_10017,N_11741);
and U12815 (N_12815,N_11234,N_11224);
and U12816 (N_12816,N_10388,N_10896);
and U12817 (N_12817,N_11528,N_11777);
and U12818 (N_12818,N_11600,N_11704);
and U12819 (N_12819,N_10437,N_10317);
nor U12820 (N_12820,N_10313,N_10682);
or U12821 (N_12821,N_10655,N_11058);
xnor U12822 (N_12822,N_11262,N_10335);
nor U12823 (N_12823,N_10397,N_11119);
xnor U12824 (N_12824,N_10040,N_11313);
xnor U12825 (N_12825,N_10753,N_10700);
nand U12826 (N_12826,N_10473,N_10944);
or U12827 (N_12827,N_11731,N_11274);
nor U12828 (N_12828,N_10623,N_10490);
and U12829 (N_12829,N_10871,N_11714);
nand U12830 (N_12830,N_11043,N_10970);
nand U12831 (N_12831,N_10659,N_10974);
nand U12832 (N_12832,N_11184,N_10062);
xnor U12833 (N_12833,N_10468,N_11832);
nand U12834 (N_12834,N_11368,N_11430);
nor U12835 (N_12835,N_10920,N_10637);
or U12836 (N_12836,N_11755,N_10277);
and U12837 (N_12837,N_11319,N_11498);
nor U12838 (N_12838,N_10100,N_10621);
nor U12839 (N_12839,N_11719,N_11773);
nor U12840 (N_12840,N_10449,N_10285);
or U12841 (N_12841,N_11522,N_11906);
and U12842 (N_12842,N_10787,N_11530);
nand U12843 (N_12843,N_10345,N_11386);
nor U12844 (N_12844,N_11940,N_10303);
nor U12845 (N_12845,N_10161,N_10204);
nor U12846 (N_12846,N_10459,N_10934);
nand U12847 (N_12847,N_10882,N_11078);
nand U12848 (N_12848,N_11993,N_11608);
and U12849 (N_12849,N_10987,N_10165);
and U12850 (N_12850,N_10500,N_10009);
xnor U12851 (N_12851,N_11382,N_10025);
xor U12852 (N_12852,N_10505,N_10444);
nand U12853 (N_12853,N_11526,N_11416);
or U12854 (N_12854,N_10986,N_10447);
nor U12855 (N_12855,N_11666,N_11056);
nand U12856 (N_12856,N_11153,N_11331);
xor U12857 (N_12857,N_10867,N_10027);
nor U12858 (N_12858,N_10737,N_10684);
and U12859 (N_12859,N_11868,N_11536);
and U12860 (N_12860,N_11178,N_11177);
and U12861 (N_12861,N_11762,N_10173);
nand U12862 (N_12862,N_10998,N_11945);
or U12863 (N_12863,N_11257,N_10252);
nor U12864 (N_12864,N_10101,N_10316);
nor U12865 (N_12865,N_11970,N_10543);
nor U12866 (N_12866,N_10918,N_10978);
xnor U12867 (N_12867,N_11525,N_11985);
and U12868 (N_12868,N_10053,N_10720);
or U12869 (N_12869,N_10496,N_10851);
xor U12870 (N_12870,N_11693,N_10328);
xnor U12871 (N_12871,N_11598,N_10481);
nand U12872 (N_12872,N_11160,N_11181);
or U12873 (N_12873,N_11466,N_11457);
or U12874 (N_12874,N_11288,N_11894);
xor U12875 (N_12875,N_10593,N_11516);
nand U12876 (N_12876,N_10368,N_11831);
and U12877 (N_12877,N_10201,N_10698);
nand U12878 (N_12878,N_11786,N_10435);
xor U12879 (N_12879,N_10913,N_10107);
xor U12880 (N_12880,N_11128,N_10074);
or U12881 (N_12881,N_10627,N_11764);
and U12882 (N_12882,N_11216,N_11996);
nand U12883 (N_12883,N_10489,N_11487);
nor U12884 (N_12884,N_11619,N_10232);
nand U12885 (N_12885,N_11320,N_11957);
or U12886 (N_12886,N_11321,N_10106);
nand U12887 (N_12887,N_11554,N_10365);
or U12888 (N_12888,N_10996,N_10797);
xor U12889 (N_12889,N_10052,N_10380);
xor U12890 (N_12890,N_11863,N_10598);
or U12891 (N_12891,N_11660,N_10728);
nor U12892 (N_12892,N_11589,N_11072);
xnor U12893 (N_12893,N_11325,N_10268);
or U12894 (N_12894,N_10724,N_10235);
or U12895 (N_12895,N_11594,N_10812);
xor U12896 (N_12896,N_11476,N_11909);
nand U12897 (N_12897,N_10358,N_11639);
or U12898 (N_12898,N_11392,N_11548);
nor U12899 (N_12899,N_11326,N_10549);
nor U12900 (N_12900,N_11752,N_10960);
nor U12901 (N_12901,N_11456,N_10807);
nor U12902 (N_12902,N_11615,N_10152);
and U12903 (N_12903,N_11981,N_10279);
xnor U12904 (N_12904,N_10363,N_10263);
and U12905 (N_12905,N_11330,N_10024);
nor U12906 (N_12906,N_11562,N_11584);
nand U12907 (N_12907,N_11656,N_10701);
nor U12908 (N_12908,N_10430,N_10820);
xor U12909 (N_12909,N_10569,N_11086);
and U12910 (N_12910,N_11998,N_11917);
nor U12911 (N_12911,N_11995,N_10613);
nor U12912 (N_12912,N_11165,N_11845);
and U12913 (N_12913,N_10952,N_10250);
nor U12914 (N_12914,N_10932,N_10671);
nand U12915 (N_12915,N_11601,N_10088);
xnor U12916 (N_12916,N_10453,N_10216);
or U12917 (N_12917,N_11532,N_11159);
nand U12918 (N_12918,N_11465,N_10906);
nor U12919 (N_12919,N_10189,N_10134);
or U12920 (N_12920,N_10219,N_10919);
or U12921 (N_12921,N_11423,N_10844);
or U12922 (N_12922,N_10205,N_11853);
nor U12923 (N_12923,N_11363,N_10680);
and U12924 (N_12924,N_11763,N_11223);
or U12925 (N_12925,N_10231,N_10594);
nor U12926 (N_12926,N_10672,N_11888);
or U12927 (N_12927,N_11295,N_10816);
nand U12928 (N_12928,N_11841,N_11163);
nor U12929 (N_12929,N_11999,N_10479);
nor U12930 (N_12930,N_11028,N_10057);
or U12931 (N_12931,N_10526,N_10497);
nor U12932 (N_12932,N_11878,N_10342);
nand U12933 (N_12933,N_10772,N_11287);
nor U12934 (N_12934,N_10726,N_10550);
and U12935 (N_12935,N_10859,N_11488);
nand U12936 (N_12936,N_10778,N_10969);
or U12937 (N_12937,N_11653,N_10291);
nand U12938 (N_12938,N_10842,N_10681);
or U12939 (N_12939,N_10729,N_11822);
nand U12940 (N_12940,N_11596,N_10597);
and U12941 (N_12941,N_10322,N_10823);
xnor U12942 (N_12942,N_11281,N_10170);
nand U12943 (N_12943,N_10766,N_11784);
nor U12944 (N_12944,N_11614,N_10663);
and U12945 (N_12945,N_11884,N_10519);
or U12946 (N_12946,N_10129,N_10611);
or U12947 (N_12947,N_11076,N_10206);
xnor U12948 (N_12948,N_10760,N_10147);
and U12949 (N_12949,N_10401,N_10329);
xnor U12950 (N_12950,N_10105,N_10858);
nor U12951 (N_12951,N_11590,N_11359);
or U12952 (N_12952,N_10347,N_11986);
xor U12953 (N_12953,N_10545,N_11580);
xor U12954 (N_12954,N_11134,N_10400);
xor U12955 (N_12955,N_11929,N_11818);
or U12956 (N_12956,N_10379,N_11166);
nor U12957 (N_12957,N_10693,N_10276);
nor U12958 (N_12958,N_10591,N_10162);
nand U12959 (N_12959,N_11454,N_11103);
or U12960 (N_12960,N_10509,N_10532);
and U12961 (N_12961,N_10539,N_11780);
or U12962 (N_12962,N_11891,N_10242);
nor U12963 (N_12963,N_11810,N_11899);
nand U12964 (N_12964,N_10777,N_11400);
or U12965 (N_12965,N_10456,N_11039);
xnor U12966 (N_12966,N_11816,N_10830);
nand U12967 (N_12967,N_11913,N_11570);
xor U12968 (N_12968,N_11503,N_10628);
nor U12969 (N_12969,N_11027,N_11558);
nor U12970 (N_12970,N_11036,N_10005);
nand U12971 (N_12971,N_11051,N_11478);
and U12972 (N_12972,N_10791,N_11628);
or U12973 (N_12973,N_10836,N_11801);
xnor U12974 (N_12974,N_10775,N_11384);
xor U12975 (N_12975,N_11143,N_11866);
and U12976 (N_12976,N_11417,N_10922);
xor U12977 (N_12977,N_11228,N_10699);
or U12978 (N_12978,N_11997,N_11226);
nor U12979 (N_12979,N_10110,N_10089);
and U12980 (N_12980,N_10065,N_10616);
or U12981 (N_12981,N_10508,N_11191);
nand U12982 (N_12982,N_11959,N_10413);
xor U12983 (N_12983,N_11983,N_10951);
xnor U12984 (N_12984,N_11314,N_11918);
nand U12985 (N_12985,N_11008,N_10612);
nand U12986 (N_12986,N_11911,N_11678);
and U12987 (N_12987,N_11835,N_11682);
xor U12988 (N_12988,N_10237,N_11495);
and U12989 (N_12989,N_11882,N_11578);
xor U12990 (N_12990,N_10647,N_11113);
nor U12991 (N_12991,N_10861,N_10580);
and U12992 (N_12992,N_10507,N_11387);
nor U12993 (N_12993,N_10426,N_10977);
and U12994 (N_12994,N_10735,N_10860);
xnor U12995 (N_12995,N_11192,N_11761);
nand U12996 (N_12996,N_11385,N_10287);
nand U12997 (N_12997,N_11716,N_11984);
or U12998 (N_12998,N_11912,N_10991);
and U12999 (N_12999,N_11663,N_10780);
xnor U13000 (N_13000,N_10469,N_11398);
and U13001 (N_13001,N_11637,N_10891);
nor U13002 (N_13002,N_10080,N_10965);
or U13003 (N_13003,N_10499,N_10207);
nand U13004 (N_13004,N_11453,N_11562);
nand U13005 (N_13005,N_11829,N_11460);
nor U13006 (N_13006,N_11422,N_11745);
xor U13007 (N_13007,N_10806,N_11275);
nand U13008 (N_13008,N_11408,N_11219);
and U13009 (N_13009,N_10224,N_11395);
nor U13010 (N_13010,N_10083,N_10226);
xor U13011 (N_13011,N_11599,N_11672);
nand U13012 (N_13012,N_11752,N_11018);
nor U13013 (N_13013,N_10594,N_10603);
or U13014 (N_13014,N_10991,N_11481);
nand U13015 (N_13015,N_11311,N_10383);
nand U13016 (N_13016,N_10235,N_11654);
xnor U13017 (N_13017,N_11491,N_10059);
nand U13018 (N_13018,N_11984,N_10334);
and U13019 (N_13019,N_11845,N_10947);
xor U13020 (N_13020,N_11035,N_10264);
nand U13021 (N_13021,N_11195,N_10874);
nor U13022 (N_13022,N_10184,N_11019);
nor U13023 (N_13023,N_11304,N_11626);
xnor U13024 (N_13024,N_10735,N_10370);
nor U13025 (N_13025,N_10575,N_10716);
nor U13026 (N_13026,N_10685,N_11589);
nor U13027 (N_13027,N_11653,N_10771);
or U13028 (N_13028,N_10270,N_10695);
xnor U13029 (N_13029,N_11466,N_10684);
nand U13030 (N_13030,N_10586,N_11188);
nor U13031 (N_13031,N_11465,N_10178);
nand U13032 (N_13032,N_11056,N_10788);
nor U13033 (N_13033,N_11720,N_11666);
xnor U13034 (N_13034,N_10817,N_10611);
nor U13035 (N_13035,N_10438,N_10469);
nor U13036 (N_13036,N_11811,N_10621);
and U13037 (N_13037,N_11781,N_11104);
nor U13038 (N_13038,N_10459,N_10820);
or U13039 (N_13039,N_10229,N_11043);
nand U13040 (N_13040,N_11037,N_11388);
xnor U13041 (N_13041,N_10327,N_11773);
xor U13042 (N_13042,N_11642,N_11530);
nor U13043 (N_13043,N_11282,N_11388);
xnor U13044 (N_13044,N_10350,N_11582);
and U13045 (N_13045,N_11408,N_11850);
nand U13046 (N_13046,N_11647,N_10333);
nand U13047 (N_13047,N_11008,N_11605);
nand U13048 (N_13048,N_10278,N_10454);
or U13049 (N_13049,N_10321,N_11811);
nand U13050 (N_13050,N_11116,N_10736);
nor U13051 (N_13051,N_10939,N_11697);
and U13052 (N_13052,N_11722,N_11308);
nor U13053 (N_13053,N_11740,N_11946);
nand U13054 (N_13054,N_11991,N_11318);
xor U13055 (N_13055,N_11378,N_11129);
xor U13056 (N_13056,N_11160,N_11212);
nand U13057 (N_13057,N_11086,N_10459);
xnor U13058 (N_13058,N_11613,N_10312);
nand U13059 (N_13059,N_10168,N_10091);
and U13060 (N_13060,N_10366,N_10360);
xor U13061 (N_13061,N_10906,N_11286);
nand U13062 (N_13062,N_11428,N_10927);
nand U13063 (N_13063,N_10531,N_10411);
and U13064 (N_13064,N_10214,N_11520);
nand U13065 (N_13065,N_11728,N_11951);
xnor U13066 (N_13066,N_10081,N_10682);
xor U13067 (N_13067,N_11572,N_10998);
or U13068 (N_13068,N_11166,N_11976);
and U13069 (N_13069,N_11898,N_11995);
xnor U13070 (N_13070,N_10977,N_10547);
nand U13071 (N_13071,N_10275,N_11669);
nor U13072 (N_13072,N_10874,N_10588);
nand U13073 (N_13073,N_11854,N_10635);
xnor U13074 (N_13074,N_10586,N_11249);
nor U13075 (N_13075,N_10755,N_10145);
and U13076 (N_13076,N_10710,N_10508);
nand U13077 (N_13077,N_10708,N_11275);
and U13078 (N_13078,N_10795,N_11230);
xnor U13079 (N_13079,N_11125,N_10082);
xnor U13080 (N_13080,N_11553,N_10195);
and U13081 (N_13081,N_11434,N_10175);
or U13082 (N_13082,N_11988,N_11370);
xnor U13083 (N_13083,N_10685,N_11988);
xnor U13084 (N_13084,N_10242,N_11916);
nand U13085 (N_13085,N_10201,N_11626);
nor U13086 (N_13086,N_11552,N_10057);
and U13087 (N_13087,N_10028,N_10296);
or U13088 (N_13088,N_10141,N_11905);
nor U13089 (N_13089,N_11153,N_10847);
and U13090 (N_13090,N_11805,N_11389);
xnor U13091 (N_13091,N_10264,N_11521);
nor U13092 (N_13092,N_11865,N_10311);
and U13093 (N_13093,N_11988,N_11537);
xor U13094 (N_13094,N_10604,N_10994);
nand U13095 (N_13095,N_11920,N_10643);
and U13096 (N_13096,N_10597,N_10109);
xor U13097 (N_13097,N_11629,N_10653);
and U13098 (N_13098,N_10623,N_11474);
nor U13099 (N_13099,N_11786,N_10070);
nand U13100 (N_13100,N_11403,N_10541);
or U13101 (N_13101,N_10073,N_10440);
or U13102 (N_13102,N_11612,N_10093);
nor U13103 (N_13103,N_10474,N_10439);
nor U13104 (N_13104,N_11014,N_11923);
or U13105 (N_13105,N_10139,N_10788);
or U13106 (N_13106,N_10017,N_10091);
nand U13107 (N_13107,N_10226,N_11424);
or U13108 (N_13108,N_11768,N_11520);
nor U13109 (N_13109,N_10154,N_11325);
and U13110 (N_13110,N_11151,N_11028);
xnor U13111 (N_13111,N_10768,N_11208);
nand U13112 (N_13112,N_11056,N_11654);
or U13113 (N_13113,N_10497,N_11076);
nor U13114 (N_13114,N_11041,N_11102);
and U13115 (N_13115,N_10590,N_10736);
and U13116 (N_13116,N_11583,N_11212);
nor U13117 (N_13117,N_10704,N_11690);
xor U13118 (N_13118,N_10312,N_10823);
or U13119 (N_13119,N_11516,N_10174);
or U13120 (N_13120,N_10338,N_11176);
or U13121 (N_13121,N_10973,N_11992);
and U13122 (N_13122,N_11437,N_10558);
and U13123 (N_13123,N_10719,N_10830);
and U13124 (N_13124,N_10976,N_10525);
or U13125 (N_13125,N_10849,N_11041);
xnor U13126 (N_13126,N_10012,N_11762);
nor U13127 (N_13127,N_11983,N_10170);
and U13128 (N_13128,N_11423,N_11368);
nand U13129 (N_13129,N_11225,N_11518);
nand U13130 (N_13130,N_10698,N_10318);
xnor U13131 (N_13131,N_11844,N_10316);
and U13132 (N_13132,N_10860,N_10000);
and U13133 (N_13133,N_10159,N_10589);
xor U13134 (N_13134,N_11315,N_10083);
nor U13135 (N_13135,N_11791,N_11142);
nor U13136 (N_13136,N_11947,N_11894);
nand U13137 (N_13137,N_11036,N_10085);
or U13138 (N_13138,N_10235,N_11496);
nor U13139 (N_13139,N_10029,N_10015);
or U13140 (N_13140,N_10317,N_11028);
and U13141 (N_13141,N_10467,N_11235);
or U13142 (N_13142,N_11898,N_11583);
or U13143 (N_13143,N_11328,N_11311);
and U13144 (N_13144,N_11053,N_11565);
nor U13145 (N_13145,N_11879,N_11176);
nor U13146 (N_13146,N_11518,N_10971);
and U13147 (N_13147,N_11850,N_10209);
and U13148 (N_13148,N_11164,N_10957);
xnor U13149 (N_13149,N_11483,N_10448);
and U13150 (N_13150,N_10505,N_11094);
nor U13151 (N_13151,N_11244,N_11697);
nand U13152 (N_13152,N_11161,N_11428);
and U13153 (N_13153,N_10083,N_11169);
nor U13154 (N_13154,N_11234,N_11076);
nand U13155 (N_13155,N_11357,N_11410);
or U13156 (N_13156,N_11435,N_11428);
or U13157 (N_13157,N_10639,N_11705);
and U13158 (N_13158,N_10358,N_11551);
or U13159 (N_13159,N_11461,N_10145);
nand U13160 (N_13160,N_11180,N_11345);
nor U13161 (N_13161,N_10203,N_11758);
xor U13162 (N_13162,N_11181,N_11452);
nand U13163 (N_13163,N_10198,N_11948);
nor U13164 (N_13164,N_10915,N_11778);
and U13165 (N_13165,N_10759,N_11394);
xnor U13166 (N_13166,N_11407,N_11977);
xor U13167 (N_13167,N_10021,N_11773);
nor U13168 (N_13168,N_10673,N_10000);
and U13169 (N_13169,N_11304,N_11203);
nor U13170 (N_13170,N_11145,N_11450);
or U13171 (N_13171,N_11551,N_11363);
nand U13172 (N_13172,N_10986,N_10523);
or U13173 (N_13173,N_10021,N_10627);
xnor U13174 (N_13174,N_10062,N_11011);
and U13175 (N_13175,N_10359,N_10900);
and U13176 (N_13176,N_10795,N_10667);
or U13177 (N_13177,N_11065,N_10325);
nand U13178 (N_13178,N_11453,N_11568);
xnor U13179 (N_13179,N_11334,N_11555);
xor U13180 (N_13180,N_10554,N_11187);
xnor U13181 (N_13181,N_10628,N_10122);
or U13182 (N_13182,N_10760,N_11354);
nand U13183 (N_13183,N_11007,N_11733);
and U13184 (N_13184,N_10388,N_10864);
xor U13185 (N_13185,N_10459,N_11130);
or U13186 (N_13186,N_11852,N_10488);
nor U13187 (N_13187,N_10737,N_10675);
nor U13188 (N_13188,N_10761,N_11748);
and U13189 (N_13189,N_11083,N_11483);
nor U13190 (N_13190,N_10704,N_11013);
or U13191 (N_13191,N_10538,N_10295);
nor U13192 (N_13192,N_10041,N_11343);
and U13193 (N_13193,N_10652,N_10878);
xor U13194 (N_13194,N_10861,N_11576);
xor U13195 (N_13195,N_10870,N_10575);
xor U13196 (N_13196,N_10865,N_11220);
nor U13197 (N_13197,N_11723,N_11346);
and U13198 (N_13198,N_11451,N_10342);
nand U13199 (N_13199,N_10929,N_10999);
or U13200 (N_13200,N_10048,N_10587);
xnor U13201 (N_13201,N_11638,N_10620);
or U13202 (N_13202,N_10667,N_10543);
nor U13203 (N_13203,N_10445,N_10577);
nor U13204 (N_13204,N_10505,N_11189);
xor U13205 (N_13205,N_11836,N_11639);
nor U13206 (N_13206,N_11919,N_11998);
nand U13207 (N_13207,N_11830,N_10311);
or U13208 (N_13208,N_11438,N_10297);
and U13209 (N_13209,N_10701,N_11587);
or U13210 (N_13210,N_11596,N_10906);
and U13211 (N_13211,N_10125,N_11417);
and U13212 (N_13212,N_11070,N_11122);
xor U13213 (N_13213,N_10017,N_11123);
nand U13214 (N_13214,N_10574,N_10035);
xnor U13215 (N_13215,N_11452,N_11356);
xnor U13216 (N_13216,N_11941,N_11156);
nand U13217 (N_13217,N_10943,N_10603);
nor U13218 (N_13218,N_11167,N_10749);
nand U13219 (N_13219,N_11260,N_10210);
nor U13220 (N_13220,N_11016,N_10561);
nor U13221 (N_13221,N_11272,N_11994);
and U13222 (N_13222,N_11431,N_10946);
nor U13223 (N_13223,N_11286,N_11990);
xnor U13224 (N_13224,N_10311,N_11516);
xor U13225 (N_13225,N_11184,N_11604);
or U13226 (N_13226,N_10947,N_10090);
nand U13227 (N_13227,N_10079,N_11593);
and U13228 (N_13228,N_10519,N_11127);
nand U13229 (N_13229,N_11080,N_11082);
xnor U13230 (N_13230,N_10121,N_10176);
and U13231 (N_13231,N_10746,N_10179);
and U13232 (N_13232,N_10371,N_11225);
and U13233 (N_13233,N_11590,N_11737);
nor U13234 (N_13234,N_11576,N_11682);
or U13235 (N_13235,N_10154,N_10045);
and U13236 (N_13236,N_10674,N_10886);
xor U13237 (N_13237,N_10679,N_10450);
nand U13238 (N_13238,N_11559,N_11931);
and U13239 (N_13239,N_11550,N_11667);
nand U13240 (N_13240,N_10040,N_11801);
nor U13241 (N_13241,N_10832,N_11463);
xnor U13242 (N_13242,N_11831,N_10383);
and U13243 (N_13243,N_10281,N_10280);
or U13244 (N_13244,N_11883,N_10093);
nor U13245 (N_13245,N_11494,N_10661);
or U13246 (N_13246,N_10666,N_11413);
or U13247 (N_13247,N_10368,N_11141);
and U13248 (N_13248,N_10877,N_11237);
xnor U13249 (N_13249,N_11609,N_10542);
or U13250 (N_13250,N_11534,N_11192);
or U13251 (N_13251,N_10745,N_11480);
nor U13252 (N_13252,N_10505,N_11146);
nand U13253 (N_13253,N_10897,N_10694);
and U13254 (N_13254,N_10329,N_11089);
xor U13255 (N_13255,N_10842,N_11676);
xor U13256 (N_13256,N_10083,N_11157);
nor U13257 (N_13257,N_10366,N_10356);
and U13258 (N_13258,N_11212,N_10271);
nand U13259 (N_13259,N_11403,N_11722);
or U13260 (N_13260,N_11997,N_11464);
nor U13261 (N_13261,N_10493,N_10250);
nor U13262 (N_13262,N_11202,N_10202);
nor U13263 (N_13263,N_10049,N_10587);
or U13264 (N_13264,N_11289,N_11986);
xor U13265 (N_13265,N_10036,N_11283);
nand U13266 (N_13266,N_10757,N_10736);
or U13267 (N_13267,N_11214,N_11166);
xnor U13268 (N_13268,N_10699,N_10593);
nand U13269 (N_13269,N_11037,N_10301);
nor U13270 (N_13270,N_11003,N_10099);
nand U13271 (N_13271,N_10564,N_10263);
xor U13272 (N_13272,N_10312,N_10035);
xor U13273 (N_13273,N_11769,N_11484);
or U13274 (N_13274,N_10848,N_10341);
nand U13275 (N_13275,N_11820,N_11650);
xor U13276 (N_13276,N_11092,N_10561);
xnor U13277 (N_13277,N_10598,N_10657);
nand U13278 (N_13278,N_10534,N_11598);
nor U13279 (N_13279,N_11172,N_11021);
or U13280 (N_13280,N_10116,N_11686);
or U13281 (N_13281,N_11083,N_11302);
or U13282 (N_13282,N_11985,N_10661);
and U13283 (N_13283,N_10802,N_11987);
or U13284 (N_13284,N_11724,N_10108);
and U13285 (N_13285,N_10910,N_11469);
or U13286 (N_13286,N_10668,N_11671);
nor U13287 (N_13287,N_10091,N_11931);
and U13288 (N_13288,N_10270,N_10373);
or U13289 (N_13289,N_10809,N_11409);
xor U13290 (N_13290,N_11809,N_10519);
and U13291 (N_13291,N_11690,N_11048);
or U13292 (N_13292,N_10930,N_10301);
nand U13293 (N_13293,N_10551,N_11591);
and U13294 (N_13294,N_10900,N_11469);
xor U13295 (N_13295,N_11097,N_10722);
and U13296 (N_13296,N_10604,N_10796);
nand U13297 (N_13297,N_10648,N_10677);
or U13298 (N_13298,N_11725,N_11029);
xnor U13299 (N_13299,N_10176,N_10766);
or U13300 (N_13300,N_11872,N_10849);
nor U13301 (N_13301,N_10197,N_10587);
and U13302 (N_13302,N_11078,N_10123);
nand U13303 (N_13303,N_10654,N_11066);
or U13304 (N_13304,N_11600,N_11495);
nor U13305 (N_13305,N_11416,N_10987);
nor U13306 (N_13306,N_10412,N_10477);
and U13307 (N_13307,N_11769,N_11370);
nand U13308 (N_13308,N_11907,N_11809);
xnor U13309 (N_13309,N_10288,N_10066);
nor U13310 (N_13310,N_11174,N_10980);
nor U13311 (N_13311,N_10064,N_11968);
or U13312 (N_13312,N_10807,N_10190);
nor U13313 (N_13313,N_11635,N_11985);
or U13314 (N_13314,N_10168,N_10046);
nand U13315 (N_13315,N_10775,N_11824);
xnor U13316 (N_13316,N_10256,N_10204);
xnor U13317 (N_13317,N_11851,N_10248);
nand U13318 (N_13318,N_11065,N_10917);
xnor U13319 (N_13319,N_11424,N_11496);
nor U13320 (N_13320,N_11268,N_10589);
or U13321 (N_13321,N_10072,N_10484);
nand U13322 (N_13322,N_11523,N_10202);
nand U13323 (N_13323,N_11606,N_11980);
nor U13324 (N_13324,N_11592,N_11039);
and U13325 (N_13325,N_11076,N_10552);
xnor U13326 (N_13326,N_11995,N_11538);
and U13327 (N_13327,N_11381,N_10378);
and U13328 (N_13328,N_11894,N_10802);
xor U13329 (N_13329,N_10212,N_10192);
nand U13330 (N_13330,N_10466,N_11061);
and U13331 (N_13331,N_10957,N_11157);
nor U13332 (N_13332,N_11826,N_10657);
and U13333 (N_13333,N_11956,N_11285);
or U13334 (N_13334,N_10696,N_11673);
nand U13335 (N_13335,N_10009,N_11455);
nor U13336 (N_13336,N_10912,N_10993);
and U13337 (N_13337,N_10758,N_11312);
or U13338 (N_13338,N_10491,N_10376);
nand U13339 (N_13339,N_11747,N_10011);
nand U13340 (N_13340,N_11413,N_11740);
xor U13341 (N_13341,N_11185,N_10766);
nor U13342 (N_13342,N_11987,N_10216);
nor U13343 (N_13343,N_11064,N_10687);
and U13344 (N_13344,N_11781,N_10482);
xnor U13345 (N_13345,N_11828,N_11208);
or U13346 (N_13346,N_10148,N_10810);
xor U13347 (N_13347,N_10166,N_11212);
xor U13348 (N_13348,N_10908,N_11092);
nand U13349 (N_13349,N_11388,N_10939);
or U13350 (N_13350,N_11254,N_11121);
or U13351 (N_13351,N_10489,N_10018);
nand U13352 (N_13352,N_11345,N_10914);
nand U13353 (N_13353,N_11944,N_11812);
xor U13354 (N_13354,N_11217,N_11245);
and U13355 (N_13355,N_10983,N_10414);
nand U13356 (N_13356,N_10946,N_10926);
xnor U13357 (N_13357,N_11393,N_11088);
nor U13358 (N_13358,N_11537,N_11011);
or U13359 (N_13359,N_10403,N_10242);
nor U13360 (N_13360,N_10001,N_10173);
and U13361 (N_13361,N_10551,N_10245);
nor U13362 (N_13362,N_10348,N_11782);
nand U13363 (N_13363,N_10867,N_10342);
or U13364 (N_13364,N_11563,N_11357);
or U13365 (N_13365,N_10920,N_11470);
or U13366 (N_13366,N_10388,N_11678);
xor U13367 (N_13367,N_11436,N_11579);
xor U13368 (N_13368,N_11151,N_11372);
and U13369 (N_13369,N_10329,N_10025);
xor U13370 (N_13370,N_10112,N_10842);
nand U13371 (N_13371,N_10238,N_10785);
and U13372 (N_13372,N_10110,N_10049);
nand U13373 (N_13373,N_10912,N_11045);
xor U13374 (N_13374,N_11129,N_10689);
or U13375 (N_13375,N_10175,N_10981);
nand U13376 (N_13376,N_11183,N_10279);
xor U13377 (N_13377,N_10843,N_11290);
or U13378 (N_13378,N_11518,N_11116);
nand U13379 (N_13379,N_10356,N_11709);
nand U13380 (N_13380,N_11333,N_11734);
xor U13381 (N_13381,N_11853,N_10510);
nor U13382 (N_13382,N_11078,N_10129);
or U13383 (N_13383,N_11219,N_10087);
nor U13384 (N_13384,N_11152,N_11038);
and U13385 (N_13385,N_10347,N_11818);
xnor U13386 (N_13386,N_10206,N_10902);
and U13387 (N_13387,N_11503,N_10220);
nand U13388 (N_13388,N_10278,N_10224);
nand U13389 (N_13389,N_10045,N_10519);
and U13390 (N_13390,N_11867,N_11780);
and U13391 (N_13391,N_11777,N_10021);
and U13392 (N_13392,N_11005,N_10255);
and U13393 (N_13393,N_11585,N_11733);
and U13394 (N_13394,N_10450,N_11611);
or U13395 (N_13395,N_11815,N_11476);
xor U13396 (N_13396,N_10448,N_11747);
or U13397 (N_13397,N_11752,N_11438);
xnor U13398 (N_13398,N_11077,N_11007);
or U13399 (N_13399,N_10124,N_10131);
xor U13400 (N_13400,N_11568,N_10697);
and U13401 (N_13401,N_10532,N_10955);
nand U13402 (N_13402,N_10509,N_11625);
or U13403 (N_13403,N_11663,N_11654);
and U13404 (N_13404,N_11342,N_11460);
xor U13405 (N_13405,N_10367,N_10001);
and U13406 (N_13406,N_11865,N_11731);
xnor U13407 (N_13407,N_11949,N_11725);
and U13408 (N_13408,N_10568,N_11687);
nor U13409 (N_13409,N_10483,N_10576);
nor U13410 (N_13410,N_11092,N_10356);
and U13411 (N_13411,N_10815,N_10134);
nor U13412 (N_13412,N_10997,N_11273);
or U13413 (N_13413,N_10565,N_10614);
and U13414 (N_13414,N_11745,N_10686);
and U13415 (N_13415,N_10295,N_11884);
or U13416 (N_13416,N_11501,N_11141);
or U13417 (N_13417,N_11731,N_10251);
and U13418 (N_13418,N_10654,N_10952);
or U13419 (N_13419,N_10392,N_11121);
xor U13420 (N_13420,N_10856,N_11189);
xnor U13421 (N_13421,N_10046,N_11664);
nand U13422 (N_13422,N_11001,N_11192);
or U13423 (N_13423,N_11286,N_11468);
nand U13424 (N_13424,N_10397,N_11674);
or U13425 (N_13425,N_11397,N_11761);
or U13426 (N_13426,N_11884,N_11488);
or U13427 (N_13427,N_10462,N_11972);
nor U13428 (N_13428,N_11473,N_10846);
or U13429 (N_13429,N_11534,N_11986);
nand U13430 (N_13430,N_10434,N_10979);
nand U13431 (N_13431,N_10430,N_10630);
nand U13432 (N_13432,N_11298,N_10538);
nor U13433 (N_13433,N_11432,N_11081);
xnor U13434 (N_13434,N_11153,N_11123);
xor U13435 (N_13435,N_10696,N_11867);
xor U13436 (N_13436,N_10750,N_11302);
nor U13437 (N_13437,N_10417,N_11659);
and U13438 (N_13438,N_11843,N_11890);
and U13439 (N_13439,N_10182,N_10906);
or U13440 (N_13440,N_10218,N_11500);
or U13441 (N_13441,N_10131,N_10410);
xnor U13442 (N_13442,N_11607,N_10565);
xor U13443 (N_13443,N_11001,N_11433);
and U13444 (N_13444,N_11775,N_11536);
or U13445 (N_13445,N_10467,N_11365);
nor U13446 (N_13446,N_11990,N_11482);
and U13447 (N_13447,N_11167,N_11475);
or U13448 (N_13448,N_11904,N_10228);
and U13449 (N_13449,N_11954,N_11487);
and U13450 (N_13450,N_11458,N_11039);
and U13451 (N_13451,N_10477,N_10584);
nor U13452 (N_13452,N_10662,N_10767);
nand U13453 (N_13453,N_11796,N_11481);
nor U13454 (N_13454,N_10204,N_10224);
nand U13455 (N_13455,N_11498,N_11460);
and U13456 (N_13456,N_11857,N_10220);
and U13457 (N_13457,N_11888,N_11870);
nand U13458 (N_13458,N_10265,N_10068);
and U13459 (N_13459,N_10715,N_10091);
xnor U13460 (N_13460,N_10282,N_10332);
and U13461 (N_13461,N_11624,N_11364);
or U13462 (N_13462,N_10167,N_11706);
xnor U13463 (N_13463,N_10219,N_11879);
xor U13464 (N_13464,N_11406,N_11369);
and U13465 (N_13465,N_10125,N_10887);
and U13466 (N_13466,N_11572,N_11623);
nor U13467 (N_13467,N_10579,N_11602);
nand U13468 (N_13468,N_11714,N_11753);
nor U13469 (N_13469,N_11797,N_10525);
and U13470 (N_13470,N_11749,N_10422);
xor U13471 (N_13471,N_11927,N_11385);
xnor U13472 (N_13472,N_10986,N_11511);
xor U13473 (N_13473,N_11123,N_11793);
or U13474 (N_13474,N_11676,N_10024);
xnor U13475 (N_13475,N_10398,N_11625);
and U13476 (N_13476,N_10972,N_10414);
nor U13477 (N_13477,N_10375,N_10745);
and U13478 (N_13478,N_10764,N_11906);
nor U13479 (N_13479,N_11898,N_10744);
and U13480 (N_13480,N_10367,N_10958);
and U13481 (N_13481,N_10660,N_11889);
nand U13482 (N_13482,N_11421,N_10925);
and U13483 (N_13483,N_10936,N_10673);
or U13484 (N_13484,N_11821,N_11777);
and U13485 (N_13485,N_10273,N_10928);
and U13486 (N_13486,N_10344,N_10728);
nor U13487 (N_13487,N_10968,N_10899);
and U13488 (N_13488,N_11862,N_11227);
or U13489 (N_13489,N_10081,N_10613);
nand U13490 (N_13490,N_11015,N_11012);
nand U13491 (N_13491,N_10140,N_11508);
and U13492 (N_13492,N_11115,N_10679);
and U13493 (N_13493,N_11188,N_11384);
and U13494 (N_13494,N_11773,N_11930);
nor U13495 (N_13495,N_11525,N_11964);
nor U13496 (N_13496,N_11800,N_10684);
and U13497 (N_13497,N_11881,N_11709);
and U13498 (N_13498,N_10572,N_11264);
xor U13499 (N_13499,N_11851,N_11266);
and U13500 (N_13500,N_11199,N_11866);
and U13501 (N_13501,N_10798,N_10589);
nand U13502 (N_13502,N_11016,N_11259);
and U13503 (N_13503,N_11678,N_10493);
nand U13504 (N_13504,N_10886,N_11483);
and U13505 (N_13505,N_10471,N_10030);
or U13506 (N_13506,N_11123,N_10831);
xor U13507 (N_13507,N_10224,N_11259);
or U13508 (N_13508,N_11181,N_10072);
nor U13509 (N_13509,N_11541,N_10060);
xnor U13510 (N_13510,N_11410,N_11551);
nor U13511 (N_13511,N_10844,N_10979);
nand U13512 (N_13512,N_10239,N_10680);
or U13513 (N_13513,N_10150,N_10052);
and U13514 (N_13514,N_10309,N_11955);
or U13515 (N_13515,N_11960,N_11135);
xor U13516 (N_13516,N_10126,N_10197);
nand U13517 (N_13517,N_10380,N_11206);
nor U13518 (N_13518,N_11189,N_10806);
and U13519 (N_13519,N_11194,N_11422);
xor U13520 (N_13520,N_10162,N_10321);
nor U13521 (N_13521,N_10069,N_11001);
xor U13522 (N_13522,N_10891,N_11168);
nand U13523 (N_13523,N_10635,N_10524);
nand U13524 (N_13524,N_10376,N_11659);
nor U13525 (N_13525,N_10843,N_10254);
xor U13526 (N_13526,N_11733,N_11869);
xor U13527 (N_13527,N_11804,N_10184);
nor U13528 (N_13528,N_10216,N_10665);
nand U13529 (N_13529,N_11102,N_11812);
or U13530 (N_13530,N_11505,N_11877);
and U13531 (N_13531,N_11823,N_11275);
nand U13532 (N_13532,N_11181,N_10469);
xor U13533 (N_13533,N_11804,N_11910);
and U13534 (N_13534,N_10031,N_10882);
or U13535 (N_13535,N_11154,N_11156);
and U13536 (N_13536,N_11930,N_10471);
and U13537 (N_13537,N_10822,N_10141);
xnor U13538 (N_13538,N_11274,N_11091);
and U13539 (N_13539,N_11888,N_11441);
nor U13540 (N_13540,N_11491,N_11912);
nand U13541 (N_13541,N_11620,N_10682);
or U13542 (N_13542,N_10868,N_11725);
nand U13543 (N_13543,N_11282,N_11286);
and U13544 (N_13544,N_11536,N_10556);
nor U13545 (N_13545,N_10364,N_11385);
xnor U13546 (N_13546,N_11144,N_11347);
or U13547 (N_13547,N_11047,N_11228);
nand U13548 (N_13548,N_11329,N_11716);
xor U13549 (N_13549,N_11437,N_10885);
xnor U13550 (N_13550,N_10564,N_10965);
or U13551 (N_13551,N_10537,N_11722);
nand U13552 (N_13552,N_11437,N_10887);
or U13553 (N_13553,N_10945,N_11028);
nor U13554 (N_13554,N_10527,N_11096);
nor U13555 (N_13555,N_10125,N_10415);
or U13556 (N_13556,N_10251,N_10566);
and U13557 (N_13557,N_10836,N_10719);
nor U13558 (N_13558,N_10877,N_11882);
nand U13559 (N_13559,N_11179,N_11592);
nand U13560 (N_13560,N_11909,N_11105);
nor U13561 (N_13561,N_11423,N_11891);
xor U13562 (N_13562,N_11230,N_10542);
nand U13563 (N_13563,N_10533,N_11526);
nor U13564 (N_13564,N_10859,N_11719);
and U13565 (N_13565,N_11680,N_11106);
xnor U13566 (N_13566,N_10842,N_11462);
or U13567 (N_13567,N_10193,N_10553);
xnor U13568 (N_13568,N_11513,N_11575);
nand U13569 (N_13569,N_10768,N_11728);
xnor U13570 (N_13570,N_11866,N_11505);
and U13571 (N_13571,N_11422,N_10609);
xnor U13572 (N_13572,N_10463,N_11798);
or U13573 (N_13573,N_11174,N_11720);
nand U13574 (N_13574,N_11420,N_10523);
and U13575 (N_13575,N_11856,N_10402);
xor U13576 (N_13576,N_10199,N_10745);
nand U13577 (N_13577,N_10173,N_11393);
xor U13578 (N_13578,N_10804,N_11302);
xor U13579 (N_13579,N_11568,N_10912);
nand U13580 (N_13580,N_10831,N_10713);
or U13581 (N_13581,N_10535,N_11134);
xnor U13582 (N_13582,N_11035,N_10951);
xor U13583 (N_13583,N_10355,N_11581);
nor U13584 (N_13584,N_10132,N_11877);
nor U13585 (N_13585,N_10123,N_11573);
nand U13586 (N_13586,N_11631,N_10582);
nor U13587 (N_13587,N_10250,N_11823);
or U13588 (N_13588,N_10080,N_10732);
nor U13589 (N_13589,N_11970,N_10582);
xor U13590 (N_13590,N_11771,N_10863);
nand U13591 (N_13591,N_11803,N_10091);
and U13592 (N_13592,N_10941,N_11979);
xor U13593 (N_13593,N_11223,N_11832);
xnor U13594 (N_13594,N_10435,N_10900);
nand U13595 (N_13595,N_10004,N_10354);
and U13596 (N_13596,N_10934,N_10736);
nor U13597 (N_13597,N_10442,N_10577);
xnor U13598 (N_13598,N_11010,N_10372);
or U13599 (N_13599,N_10379,N_10689);
or U13600 (N_13600,N_10145,N_10636);
nand U13601 (N_13601,N_10392,N_10020);
and U13602 (N_13602,N_10452,N_10253);
xor U13603 (N_13603,N_10327,N_11186);
xnor U13604 (N_13604,N_10473,N_11306);
nor U13605 (N_13605,N_11368,N_10352);
or U13606 (N_13606,N_10948,N_10014);
nand U13607 (N_13607,N_10024,N_11530);
or U13608 (N_13608,N_11609,N_11150);
and U13609 (N_13609,N_11964,N_10389);
xnor U13610 (N_13610,N_10291,N_11384);
nand U13611 (N_13611,N_11500,N_11720);
or U13612 (N_13612,N_10399,N_11131);
nor U13613 (N_13613,N_11492,N_10677);
xnor U13614 (N_13614,N_11110,N_10775);
xnor U13615 (N_13615,N_10966,N_11519);
and U13616 (N_13616,N_10006,N_11057);
nand U13617 (N_13617,N_11649,N_10765);
and U13618 (N_13618,N_10357,N_11930);
or U13619 (N_13619,N_11425,N_10229);
nand U13620 (N_13620,N_10620,N_11155);
or U13621 (N_13621,N_11262,N_11464);
nand U13622 (N_13622,N_10619,N_10703);
and U13623 (N_13623,N_10797,N_11269);
and U13624 (N_13624,N_11369,N_10192);
and U13625 (N_13625,N_10973,N_10743);
or U13626 (N_13626,N_11159,N_10989);
xnor U13627 (N_13627,N_11666,N_11188);
nand U13628 (N_13628,N_10825,N_11324);
and U13629 (N_13629,N_11388,N_10819);
nor U13630 (N_13630,N_10912,N_10094);
or U13631 (N_13631,N_11540,N_10787);
nand U13632 (N_13632,N_10048,N_10995);
nand U13633 (N_13633,N_11985,N_11137);
or U13634 (N_13634,N_10823,N_10791);
nand U13635 (N_13635,N_11064,N_10939);
and U13636 (N_13636,N_11010,N_11186);
nand U13637 (N_13637,N_10549,N_10389);
or U13638 (N_13638,N_11797,N_11745);
or U13639 (N_13639,N_11885,N_10522);
and U13640 (N_13640,N_11032,N_10276);
xnor U13641 (N_13641,N_11779,N_10662);
and U13642 (N_13642,N_10877,N_11417);
xnor U13643 (N_13643,N_11571,N_11103);
nor U13644 (N_13644,N_11024,N_11368);
xor U13645 (N_13645,N_11559,N_10666);
and U13646 (N_13646,N_11452,N_10120);
nand U13647 (N_13647,N_10885,N_10681);
xor U13648 (N_13648,N_11054,N_10265);
and U13649 (N_13649,N_10040,N_11914);
nor U13650 (N_13650,N_11704,N_10204);
and U13651 (N_13651,N_11243,N_11918);
and U13652 (N_13652,N_10405,N_10939);
xnor U13653 (N_13653,N_10884,N_11319);
and U13654 (N_13654,N_11235,N_10798);
or U13655 (N_13655,N_10272,N_10886);
nor U13656 (N_13656,N_10168,N_11648);
or U13657 (N_13657,N_10431,N_11048);
xor U13658 (N_13658,N_10733,N_10081);
xnor U13659 (N_13659,N_10140,N_11183);
and U13660 (N_13660,N_11340,N_11653);
nand U13661 (N_13661,N_10183,N_11067);
and U13662 (N_13662,N_10650,N_10026);
xor U13663 (N_13663,N_10026,N_11651);
or U13664 (N_13664,N_11534,N_10826);
nand U13665 (N_13665,N_10840,N_11064);
xor U13666 (N_13666,N_11752,N_11425);
nor U13667 (N_13667,N_10133,N_11307);
nor U13668 (N_13668,N_11727,N_11916);
or U13669 (N_13669,N_11586,N_11951);
xnor U13670 (N_13670,N_11948,N_10352);
xnor U13671 (N_13671,N_11138,N_11505);
nand U13672 (N_13672,N_10959,N_10052);
nor U13673 (N_13673,N_11810,N_10201);
nor U13674 (N_13674,N_10144,N_11808);
xnor U13675 (N_13675,N_10958,N_11336);
nor U13676 (N_13676,N_11821,N_11443);
xor U13677 (N_13677,N_11620,N_11428);
xnor U13678 (N_13678,N_11728,N_11120);
nand U13679 (N_13679,N_11918,N_11440);
and U13680 (N_13680,N_10612,N_10703);
or U13681 (N_13681,N_11997,N_10475);
and U13682 (N_13682,N_10095,N_11911);
and U13683 (N_13683,N_11566,N_11282);
or U13684 (N_13684,N_11916,N_11841);
xor U13685 (N_13685,N_10419,N_10889);
and U13686 (N_13686,N_10064,N_11624);
nand U13687 (N_13687,N_10513,N_11945);
nand U13688 (N_13688,N_11796,N_10716);
and U13689 (N_13689,N_11698,N_10249);
nor U13690 (N_13690,N_11646,N_10247);
nand U13691 (N_13691,N_11878,N_11367);
nand U13692 (N_13692,N_11783,N_10053);
or U13693 (N_13693,N_10078,N_10448);
or U13694 (N_13694,N_10248,N_11076);
nand U13695 (N_13695,N_10526,N_11861);
and U13696 (N_13696,N_10594,N_10918);
xor U13697 (N_13697,N_11011,N_10399);
xnor U13698 (N_13698,N_11329,N_10079);
or U13699 (N_13699,N_10736,N_11931);
and U13700 (N_13700,N_11740,N_10772);
and U13701 (N_13701,N_10575,N_11811);
or U13702 (N_13702,N_11593,N_10968);
xnor U13703 (N_13703,N_10111,N_11450);
nand U13704 (N_13704,N_10986,N_10448);
nand U13705 (N_13705,N_10877,N_11408);
or U13706 (N_13706,N_11607,N_11419);
or U13707 (N_13707,N_11954,N_11089);
nor U13708 (N_13708,N_10058,N_11643);
or U13709 (N_13709,N_10459,N_11123);
and U13710 (N_13710,N_10519,N_11655);
or U13711 (N_13711,N_10551,N_11038);
and U13712 (N_13712,N_11390,N_10697);
nor U13713 (N_13713,N_10826,N_10199);
xor U13714 (N_13714,N_10041,N_11419);
nand U13715 (N_13715,N_11473,N_11173);
xor U13716 (N_13716,N_11500,N_10881);
xor U13717 (N_13717,N_11132,N_10625);
xor U13718 (N_13718,N_11418,N_10305);
nand U13719 (N_13719,N_10368,N_10553);
nor U13720 (N_13720,N_10409,N_10044);
nor U13721 (N_13721,N_10499,N_11330);
nand U13722 (N_13722,N_11848,N_11567);
nor U13723 (N_13723,N_10574,N_10990);
and U13724 (N_13724,N_11537,N_10371);
and U13725 (N_13725,N_11336,N_11013);
nor U13726 (N_13726,N_10739,N_10869);
xnor U13727 (N_13727,N_10160,N_11152);
nand U13728 (N_13728,N_10212,N_10772);
nand U13729 (N_13729,N_10395,N_10010);
xnor U13730 (N_13730,N_11177,N_11562);
or U13731 (N_13731,N_11442,N_11178);
xnor U13732 (N_13732,N_10430,N_11667);
nand U13733 (N_13733,N_11444,N_10737);
or U13734 (N_13734,N_10372,N_11219);
xnor U13735 (N_13735,N_10290,N_10155);
or U13736 (N_13736,N_11114,N_10975);
nor U13737 (N_13737,N_11269,N_10878);
or U13738 (N_13738,N_10602,N_10336);
xnor U13739 (N_13739,N_10783,N_10796);
nand U13740 (N_13740,N_10504,N_10863);
xnor U13741 (N_13741,N_10133,N_11102);
xnor U13742 (N_13742,N_10206,N_10443);
nand U13743 (N_13743,N_11896,N_10634);
nor U13744 (N_13744,N_10473,N_10579);
nor U13745 (N_13745,N_10017,N_10842);
xor U13746 (N_13746,N_10472,N_11155);
or U13747 (N_13747,N_11576,N_10257);
nand U13748 (N_13748,N_10779,N_10894);
xnor U13749 (N_13749,N_10286,N_10312);
nor U13750 (N_13750,N_10348,N_10051);
nand U13751 (N_13751,N_11530,N_10611);
nor U13752 (N_13752,N_11225,N_11731);
or U13753 (N_13753,N_11769,N_10882);
or U13754 (N_13754,N_10971,N_11493);
xnor U13755 (N_13755,N_11713,N_11875);
or U13756 (N_13756,N_10355,N_10057);
and U13757 (N_13757,N_11144,N_10669);
nand U13758 (N_13758,N_10861,N_11723);
xor U13759 (N_13759,N_11686,N_10222);
nor U13760 (N_13760,N_10513,N_10477);
or U13761 (N_13761,N_10935,N_11948);
xor U13762 (N_13762,N_10841,N_10685);
and U13763 (N_13763,N_11481,N_11042);
nor U13764 (N_13764,N_10522,N_10152);
or U13765 (N_13765,N_10199,N_10540);
nand U13766 (N_13766,N_10312,N_10556);
nor U13767 (N_13767,N_11660,N_11375);
nand U13768 (N_13768,N_11740,N_11463);
or U13769 (N_13769,N_10270,N_11533);
nand U13770 (N_13770,N_11704,N_10222);
xor U13771 (N_13771,N_11874,N_11233);
nand U13772 (N_13772,N_10223,N_11325);
xnor U13773 (N_13773,N_10228,N_10115);
xor U13774 (N_13774,N_11174,N_10762);
xnor U13775 (N_13775,N_11863,N_10135);
nand U13776 (N_13776,N_11758,N_10820);
xor U13777 (N_13777,N_10004,N_10289);
and U13778 (N_13778,N_10566,N_10209);
nor U13779 (N_13779,N_11474,N_11159);
and U13780 (N_13780,N_11213,N_11537);
nand U13781 (N_13781,N_10453,N_10464);
or U13782 (N_13782,N_11968,N_11298);
or U13783 (N_13783,N_11698,N_11776);
nor U13784 (N_13784,N_10077,N_10012);
or U13785 (N_13785,N_11980,N_10686);
and U13786 (N_13786,N_10765,N_10683);
or U13787 (N_13787,N_10327,N_10147);
and U13788 (N_13788,N_10123,N_10425);
and U13789 (N_13789,N_10436,N_11776);
nor U13790 (N_13790,N_10360,N_10992);
xnor U13791 (N_13791,N_10408,N_11215);
xnor U13792 (N_13792,N_10274,N_11684);
or U13793 (N_13793,N_10553,N_10386);
and U13794 (N_13794,N_11387,N_10014);
xor U13795 (N_13795,N_11026,N_11486);
or U13796 (N_13796,N_10264,N_10570);
or U13797 (N_13797,N_11109,N_11866);
or U13798 (N_13798,N_10447,N_10954);
xor U13799 (N_13799,N_11236,N_10300);
nand U13800 (N_13800,N_11095,N_10334);
and U13801 (N_13801,N_10392,N_11439);
and U13802 (N_13802,N_10930,N_11391);
xor U13803 (N_13803,N_10458,N_10806);
xor U13804 (N_13804,N_11041,N_11543);
nand U13805 (N_13805,N_10794,N_11179);
nand U13806 (N_13806,N_10299,N_10108);
xnor U13807 (N_13807,N_10669,N_10687);
xnor U13808 (N_13808,N_11682,N_10595);
and U13809 (N_13809,N_10874,N_11896);
nand U13810 (N_13810,N_11061,N_10833);
nand U13811 (N_13811,N_10800,N_10918);
nand U13812 (N_13812,N_10107,N_11890);
nand U13813 (N_13813,N_10533,N_10593);
nand U13814 (N_13814,N_11619,N_11162);
xnor U13815 (N_13815,N_11173,N_10027);
or U13816 (N_13816,N_11384,N_11668);
xor U13817 (N_13817,N_10448,N_10809);
or U13818 (N_13818,N_11109,N_10638);
nand U13819 (N_13819,N_10903,N_11027);
xor U13820 (N_13820,N_11593,N_11361);
xor U13821 (N_13821,N_11124,N_11303);
xnor U13822 (N_13822,N_10611,N_11923);
nand U13823 (N_13823,N_11971,N_10746);
or U13824 (N_13824,N_11516,N_10373);
xnor U13825 (N_13825,N_10108,N_10236);
or U13826 (N_13826,N_10393,N_10317);
or U13827 (N_13827,N_10583,N_10089);
xor U13828 (N_13828,N_10388,N_11478);
nor U13829 (N_13829,N_10271,N_11336);
xor U13830 (N_13830,N_11370,N_11621);
or U13831 (N_13831,N_10719,N_11858);
or U13832 (N_13832,N_10573,N_10280);
nor U13833 (N_13833,N_10772,N_10008);
or U13834 (N_13834,N_10909,N_10089);
or U13835 (N_13835,N_10158,N_10268);
xnor U13836 (N_13836,N_11441,N_11637);
nand U13837 (N_13837,N_10043,N_10940);
and U13838 (N_13838,N_10912,N_11457);
xor U13839 (N_13839,N_10281,N_10004);
nor U13840 (N_13840,N_11439,N_11829);
and U13841 (N_13841,N_10678,N_11152);
and U13842 (N_13842,N_11277,N_10468);
or U13843 (N_13843,N_10932,N_11887);
nand U13844 (N_13844,N_11939,N_11342);
nand U13845 (N_13845,N_10515,N_10364);
or U13846 (N_13846,N_10605,N_10469);
nand U13847 (N_13847,N_11283,N_11591);
xor U13848 (N_13848,N_11991,N_11965);
and U13849 (N_13849,N_11234,N_11702);
and U13850 (N_13850,N_10252,N_10413);
or U13851 (N_13851,N_10561,N_11265);
and U13852 (N_13852,N_10504,N_10880);
nand U13853 (N_13853,N_11377,N_10707);
or U13854 (N_13854,N_10152,N_11461);
and U13855 (N_13855,N_11103,N_10163);
and U13856 (N_13856,N_10876,N_11763);
xor U13857 (N_13857,N_10605,N_10248);
nand U13858 (N_13858,N_11826,N_11581);
nand U13859 (N_13859,N_10749,N_10816);
or U13860 (N_13860,N_11773,N_10373);
or U13861 (N_13861,N_10953,N_10226);
nor U13862 (N_13862,N_10422,N_11610);
nor U13863 (N_13863,N_10614,N_11020);
nand U13864 (N_13864,N_11297,N_10429);
and U13865 (N_13865,N_10836,N_11152);
and U13866 (N_13866,N_11078,N_11342);
and U13867 (N_13867,N_11810,N_11325);
and U13868 (N_13868,N_11860,N_11777);
nor U13869 (N_13869,N_10273,N_10256);
xnor U13870 (N_13870,N_11437,N_11068);
nand U13871 (N_13871,N_11538,N_11893);
xnor U13872 (N_13872,N_10323,N_10739);
or U13873 (N_13873,N_10469,N_11709);
xnor U13874 (N_13874,N_11625,N_11830);
xnor U13875 (N_13875,N_11652,N_10661);
xor U13876 (N_13876,N_11761,N_11936);
nor U13877 (N_13877,N_10561,N_10024);
nor U13878 (N_13878,N_10649,N_11003);
nor U13879 (N_13879,N_11528,N_10712);
nand U13880 (N_13880,N_10679,N_11258);
nor U13881 (N_13881,N_11805,N_10755);
and U13882 (N_13882,N_10127,N_10382);
nand U13883 (N_13883,N_10233,N_11819);
and U13884 (N_13884,N_11085,N_10190);
or U13885 (N_13885,N_10325,N_10981);
or U13886 (N_13886,N_10164,N_10502);
and U13887 (N_13887,N_11991,N_11050);
and U13888 (N_13888,N_11145,N_10047);
and U13889 (N_13889,N_11601,N_10473);
xor U13890 (N_13890,N_10939,N_11837);
or U13891 (N_13891,N_11327,N_10702);
xnor U13892 (N_13892,N_11455,N_10639);
and U13893 (N_13893,N_11313,N_10357);
nor U13894 (N_13894,N_10838,N_10630);
nand U13895 (N_13895,N_10030,N_10096);
and U13896 (N_13896,N_11289,N_11459);
nand U13897 (N_13897,N_10039,N_11948);
xor U13898 (N_13898,N_10064,N_11926);
or U13899 (N_13899,N_11683,N_11665);
nor U13900 (N_13900,N_10212,N_10600);
or U13901 (N_13901,N_11271,N_10899);
or U13902 (N_13902,N_11473,N_11180);
and U13903 (N_13903,N_11352,N_10377);
or U13904 (N_13904,N_10698,N_10639);
nor U13905 (N_13905,N_11427,N_11171);
or U13906 (N_13906,N_10293,N_11170);
nor U13907 (N_13907,N_10639,N_11950);
nor U13908 (N_13908,N_10661,N_10558);
nand U13909 (N_13909,N_10159,N_11389);
or U13910 (N_13910,N_10400,N_10101);
xnor U13911 (N_13911,N_10646,N_11804);
xor U13912 (N_13912,N_11226,N_10710);
nor U13913 (N_13913,N_11044,N_10087);
nand U13914 (N_13914,N_10945,N_10785);
xor U13915 (N_13915,N_11395,N_11029);
nor U13916 (N_13916,N_10388,N_10989);
and U13917 (N_13917,N_10676,N_11758);
and U13918 (N_13918,N_10374,N_11490);
or U13919 (N_13919,N_11921,N_11285);
nand U13920 (N_13920,N_10391,N_11549);
xor U13921 (N_13921,N_11843,N_10622);
xnor U13922 (N_13922,N_11534,N_11542);
and U13923 (N_13923,N_11018,N_11708);
nand U13924 (N_13924,N_10344,N_10343);
and U13925 (N_13925,N_11063,N_11507);
xor U13926 (N_13926,N_10505,N_11280);
nand U13927 (N_13927,N_10811,N_11143);
or U13928 (N_13928,N_11584,N_11648);
or U13929 (N_13929,N_10540,N_10072);
or U13930 (N_13930,N_10382,N_10601);
xor U13931 (N_13931,N_11972,N_11005);
xnor U13932 (N_13932,N_11234,N_10298);
and U13933 (N_13933,N_10836,N_10460);
and U13934 (N_13934,N_10041,N_11601);
and U13935 (N_13935,N_11702,N_11838);
and U13936 (N_13936,N_11626,N_10785);
and U13937 (N_13937,N_10178,N_11820);
xnor U13938 (N_13938,N_10576,N_11044);
or U13939 (N_13939,N_11632,N_10278);
and U13940 (N_13940,N_10163,N_10302);
nand U13941 (N_13941,N_10972,N_11605);
xor U13942 (N_13942,N_10366,N_10475);
xor U13943 (N_13943,N_11761,N_11946);
or U13944 (N_13944,N_10669,N_11922);
and U13945 (N_13945,N_11324,N_10873);
nor U13946 (N_13946,N_11256,N_11836);
or U13947 (N_13947,N_10159,N_11922);
and U13948 (N_13948,N_10910,N_10946);
xnor U13949 (N_13949,N_10989,N_11855);
xnor U13950 (N_13950,N_10860,N_11777);
nand U13951 (N_13951,N_10804,N_10813);
xor U13952 (N_13952,N_10825,N_11559);
and U13953 (N_13953,N_10893,N_10826);
nor U13954 (N_13954,N_11595,N_11637);
nand U13955 (N_13955,N_10280,N_10882);
and U13956 (N_13956,N_11958,N_11414);
xor U13957 (N_13957,N_10345,N_10149);
nor U13958 (N_13958,N_11093,N_11270);
nor U13959 (N_13959,N_11800,N_10810);
or U13960 (N_13960,N_10080,N_11757);
and U13961 (N_13961,N_11941,N_10521);
nor U13962 (N_13962,N_11970,N_10013);
nand U13963 (N_13963,N_11433,N_11046);
and U13964 (N_13964,N_10488,N_11552);
xor U13965 (N_13965,N_10361,N_10988);
nor U13966 (N_13966,N_10186,N_11921);
xnor U13967 (N_13967,N_11033,N_10163);
or U13968 (N_13968,N_10254,N_11727);
and U13969 (N_13969,N_11582,N_11618);
or U13970 (N_13970,N_11836,N_10128);
nand U13971 (N_13971,N_11070,N_10215);
nor U13972 (N_13972,N_11112,N_10197);
or U13973 (N_13973,N_10279,N_11323);
or U13974 (N_13974,N_10004,N_11386);
or U13975 (N_13975,N_10700,N_10800);
and U13976 (N_13976,N_10809,N_10098);
nor U13977 (N_13977,N_10901,N_10697);
nand U13978 (N_13978,N_11501,N_10640);
and U13979 (N_13979,N_11362,N_10436);
or U13980 (N_13980,N_10161,N_10914);
nor U13981 (N_13981,N_10566,N_11640);
or U13982 (N_13982,N_10157,N_10848);
and U13983 (N_13983,N_10249,N_11515);
or U13984 (N_13984,N_10723,N_10773);
xnor U13985 (N_13985,N_10914,N_11073);
xor U13986 (N_13986,N_10974,N_10159);
nand U13987 (N_13987,N_11205,N_11728);
xnor U13988 (N_13988,N_10696,N_11860);
nor U13989 (N_13989,N_11248,N_10342);
xor U13990 (N_13990,N_10212,N_11791);
nor U13991 (N_13991,N_10451,N_10484);
nand U13992 (N_13992,N_11313,N_11236);
and U13993 (N_13993,N_11391,N_10027);
nor U13994 (N_13994,N_10635,N_10056);
or U13995 (N_13995,N_10579,N_10824);
nor U13996 (N_13996,N_11583,N_10156);
nand U13997 (N_13997,N_10307,N_11929);
nor U13998 (N_13998,N_10504,N_10453);
or U13999 (N_13999,N_10245,N_11940);
xnor U14000 (N_14000,N_12247,N_12656);
nor U14001 (N_14001,N_13200,N_12837);
xnor U14002 (N_14002,N_13108,N_13503);
or U14003 (N_14003,N_13506,N_12791);
and U14004 (N_14004,N_12955,N_13550);
nor U14005 (N_14005,N_12331,N_13653);
nor U14006 (N_14006,N_12415,N_12567);
nor U14007 (N_14007,N_12764,N_13368);
nor U14008 (N_14008,N_12281,N_13651);
or U14009 (N_14009,N_12217,N_13773);
nor U14010 (N_14010,N_13131,N_13976);
nand U14011 (N_14011,N_13458,N_13135);
and U14012 (N_14012,N_12362,N_12352);
nand U14013 (N_14013,N_13968,N_12034);
xor U14014 (N_14014,N_13327,N_13879);
nand U14015 (N_14015,N_12580,N_13222);
nor U14016 (N_14016,N_12702,N_12111);
or U14017 (N_14017,N_13897,N_12798);
nand U14018 (N_14018,N_12389,N_12280);
nand U14019 (N_14019,N_13679,N_13054);
nand U14020 (N_14020,N_12070,N_13628);
and U14021 (N_14021,N_13514,N_12860);
and U14022 (N_14022,N_12479,N_12598);
or U14023 (N_14023,N_12967,N_13875);
and U14024 (N_14024,N_12525,N_12035);
nand U14025 (N_14025,N_12768,N_13067);
nand U14026 (N_14026,N_13584,N_13310);
and U14027 (N_14027,N_12164,N_13500);
xnor U14028 (N_14028,N_12369,N_13640);
nor U14029 (N_14029,N_13943,N_13918);
and U14030 (N_14030,N_13055,N_12265);
nor U14031 (N_14031,N_12549,N_12098);
or U14032 (N_14032,N_13595,N_13161);
and U14033 (N_14033,N_12646,N_13644);
or U14034 (N_14034,N_13190,N_13507);
xnor U14035 (N_14035,N_12948,N_13895);
or U14036 (N_14036,N_13780,N_13112);
xor U14037 (N_14037,N_12543,N_12480);
nand U14038 (N_14038,N_12729,N_13206);
xnor U14039 (N_14039,N_12212,N_13949);
nor U14040 (N_14040,N_12855,N_13659);
nand U14041 (N_14041,N_13303,N_13522);
xnor U14042 (N_14042,N_13304,N_12260);
or U14043 (N_14043,N_12895,N_13607);
nor U14044 (N_14044,N_13936,N_13165);
xnor U14045 (N_14045,N_12533,N_12752);
or U14046 (N_14046,N_13255,N_13818);
xnor U14047 (N_14047,N_12856,N_12706);
or U14048 (N_14048,N_13034,N_12541);
and U14049 (N_14049,N_12686,N_12645);
nand U14050 (N_14050,N_13783,N_13591);
and U14051 (N_14051,N_13297,N_13151);
and U14052 (N_14052,N_12202,N_13878);
xnor U14053 (N_14053,N_12232,N_13233);
nor U14054 (N_14054,N_13865,N_13967);
nor U14055 (N_14055,N_13900,N_13366);
or U14056 (N_14056,N_13828,N_13863);
nor U14057 (N_14057,N_12565,N_12441);
xnor U14058 (N_14058,N_12340,N_12169);
nand U14059 (N_14059,N_12896,N_13612);
nor U14060 (N_14060,N_12078,N_13502);
nand U14061 (N_14061,N_12172,N_13927);
xnor U14062 (N_14062,N_13431,N_13349);
nor U14063 (N_14063,N_12501,N_12294);
or U14064 (N_14064,N_12476,N_13642);
or U14065 (N_14065,N_13429,N_12321);
nand U14066 (N_14066,N_12296,N_13844);
xnor U14067 (N_14067,N_13602,N_12507);
nand U14068 (N_14068,N_12277,N_13469);
nand U14069 (N_14069,N_12603,N_12100);
or U14070 (N_14070,N_13238,N_12150);
xor U14071 (N_14071,N_12890,N_12724);
or U14072 (N_14072,N_13701,N_12670);
nor U14073 (N_14073,N_12960,N_12191);
nand U14074 (N_14074,N_12809,N_13555);
nor U14075 (N_14075,N_13258,N_13717);
nor U14076 (N_14076,N_13080,N_13561);
nor U14077 (N_14077,N_12511,N_13559);
or U14078 (N_14078,N_13951,N_13164);
and U14079 (N_14079,N_12651,N_12385);
xnor U14080 (N_14080,N_13107,N_12317);
xnor U14081 (N_14081,N_13339,N_12931);
xnor U14082 (N_14082,N_12332,N_12721);
and U14083 (N_14083,N_13988,N_12137);
xnor U14084 (N_14084,N_13808,N_13925);
xor U14085 (N_14085,N_12159,N_12965);
and U14086 (N_14086,N_13075,N_13660);
or U14087 (N_14087,N_13434,N_12526);
or U14088 (N_14088,N_12003,N_13053);
and U14089 (N_14089,N_12915,N_12971);
nand U14090 (N_14090,N_13243,N_12263);
nand U14091 (N_14091,N_12400,N_13630);
nand U14092 (N_14092,N_12840,N_12887);
nor U14093 (N_14093,N_13914,N_12311);
or U14094 (N_14094,N_13296,N_12826);
and U14095 (N_14095,N_12088,N_12066);
and U14096 (N_14096,N_12341,N_12395);
and U14097 (N_14097,N_12658,N_12155);
nor U14098 (N_14098,N_12545,N_12313);
xnor U14099 (N_14099,N_12393,N_13641);
or U14100 (N_14100,N_13025,N_13188);
nor U14101 (N_14101,N_12818,N_13722);
xor U14102 (N_14102,N_12858,N_12685);
and U14103 (N_14103,N_12118,N_12322);
and U14104 (N_14104,N_13718,N_13420);
or U14105 (N_14105,N_12287,N_13216);
xnor U14106 (N_14106,N_12166,N_12816);
nor U14107 (N_14107,N_12142,N_13299);
nor U14108 (N_14108,N_12167,N_13669);
nand U14109 (N_14109,N_13713,N_13741);
or U14110 (N_14110,N_12497,N_13472);
and U14111 (N_14111,N_13197,N_13372);
or U14112 (N_14112,N_12741,N_12097);
or U14113 (N_14113,N_13770,N_12197);
and U14114 (N_14114,N_13110,N_13113);
and U14115 (N_14115,N_12367,N_13556);
nand U14116 (N_14116,N_12380,N_13204);
and U14117 (N_14117,N_12410,N_12170);
or U14118 (N_14118,N_13891,N_13913);
or U14119 (N_14119,N_12248,N_12176);
nand U14120 (N_14120,N_13769,N_12128);
and U14121 (N_14121,N_12359,N_12740);
nor U14122 (N_14122,N_13427,N_13235);
nand U14123 (N_14123,N_12929,N_13163);
nand U14124 (N_14124,N_12508,N_12772);
nand U14125 (N_14125,N_13646,N_12119);
nor U14126 (N_14126,N_12368,N_13426);
and U14127 (N_14127,N_13511,N_12730);
nand U14128 (N_14128,N_12534,N_12786);
or U14129 (N_14129,N_12889,N_13333);
nor U14130 (N_14130,N_12490,N_13470);
nand U14131 (N_14131,N_12274,N_12671);
and U14132 (N_14132,N_12151,N_13886);
nand U14133 (N_14133,N_12981,N_12987);
nand U14134 (N_14134,N_13744,N_12950);
nand U14135 (N_14135,N_13811,N_13829);
nand U14136 (N_14136,N_12186,N_13390);
and U14137 (N_14137,N_13589,N_12596);
nand U14138 (N_14138,N_13980,N_12920);
nand U14139 (N_14139,N_12355,N_13767);
xnor U14140 (N_14140,N_12440,N_12102);
and U14141 (N_14141,N_12267,N_13010);
nand U14142 (N_14142,N_13089,N_12584);
xor U14143 (N_14143,N_12329,N_12949);
or U14144 (N_14144,N_12214,N_12503);
nand U14145 (N_14145,N_12835,N_12160);
or U14146 (N_14146,N_13298,N_13248);
xor U14147 (N_14147,N_12973,N_13850);
nor U14148 (N_14148,N_12557,N_13564);
xnor U14149 (N_14149,N_12897,N_13130);
nor U14150 (N_14150,N_13144,N_12831);
or U14151 (N_14151,N_13379,N_13497);
xnor U14152 (N_14152,N_12956,N_12778);
nand U14153 (N_14153,N_12796,N_12140);
nand U14154 (N_14154,N_12423,N_13708);
nor U14155 (N_14155,N_12374,N_13521);
and U14156 (N_14156,N_12001,N_13187);
and U14157 (N_14157,N_12917,N_12623);
and U14158 (N_14158,N_12542,N_12455);
xor U14159 (N_14159,N_12631,N_12813);
or U14160 (N_14160,N_12642,N_13457);
or U14161 (N_14161,N_12802,N_12841);
or U14162 (N_14162,N_13068,N_12141);
or U14163 (N_14163,N_13202,N_13726);
nor U14164 (N_14164,N_12624,N_13292);
nor U14165 (N_14165,N_13421,N_12854);
nand U14166 (N_14166,N_13237,N_13905);
nor U14167 (N_14167,N_12282,N_12201);
and U14168 (N_14168,N_13035,N_12095);
xnor U14169 (N_14169,N_12607,N_13986);
nand U14170 (N_14170,N_13317,N_12975);
xor U14171 (N_14171,N_13320,N_13389);
or U14172 (N_14172,N_13162,N_13450);
and U14173 (N_14173,N_13846,N_13795);
or U14174 (N_14174,N_12643,N_12418);
xnor U14175 (N_14175,N_12587,N_13479);
xor U14176 (N_14176,N_13820,N_13854);
xnor U14177 (N_14177,N_13051,N_13186);
and U14178 (N_14178,N_12581,N_13170);
nand U14179 (N_14179,N_13388,N_12273);
xor U14180 (N_14180,N_12062,N_13734);
or U14181 (N_14181,N_13154,N_12583);
xnor U14182 (N_14182,N_12928,N_13690);
nor U14183 (N_14183,N_13313,N_12306);
nor U14184 (N_14184,N_13785,N_12892);
xnor U14185 (N_14185,N_13894,N_13580);
and U14186 (N_14186,N_12024,N_12420);
xor U14187 (N_14187,N_12614,N_13592);
nand U14188 (N_14188,N_12774,N_13417);
nand U14189 (N_14189,N_12943,N_13856);
and U14190 (N_14190,N_12983,N_12751);
nand U14191 (N_14191,N_12424,N_12653);
or U14192 (N_14192,N_13563,N_13308);
nand U14193 (N_14193,N_13625,N_13181);
xor U14194 (N_14194,N_12980,N_12015);
or U14195 (N_14195,N_13953,N_13833);
nand U14196 (N_14196,N_13413,N_13684);
nand U14197 (N_14197,N_13316,N_13945);
nor U14198 (N_14198,N_12077,N_12032);
xnor U14199 (N_14199,N_13490,N_12731);
nand U14200 (N_14200,N_12438,N_13733);
xnor U14201 (N_14201,N_12822,N_13473);
nand U14202 (N_14202,N_13843,N_12944);
or U14203 (N_14203,N_12207,N_12789);
nor U14204 (N_14204,N_13066,N_12254);
or U14205 (N_14205,N_13280,N_12365);
nand U14206 (N_14206,N_13582,N_13146);
nor U14207 (N_14207,N_13015,N_12055);
nor U14208 (N_14208,N_12152,N_13018);
xor U14209 (N_14209,N_12022,N_12688);
nor U14210 (N_14210,N_12237,N_13750);
nor U14211 (N_14211,N_12635,N_13096);
xor U14212 (N_14212,N_13452,N_13937);
or U14213 (N_14213,N_13645,N_12605);
or U14214 (N_14214,N_13888,N_12712);
nand U14215 (N_14215,N_13610,N_13736);
and U14216 (N_14216,N_13209,N_13959);
nand U14217 (N_14217,N_12597,N_12958);
nor U14218 (N_14218,N_12448,N_12269);
nor U14219 (N_14219,N_12617,N_12315);
nand U14220 (N_14220,N_12211,N_12402);
or U14221 (N_14221,N_12450,N_12904);
or U14222 (N_14222,N_13069,N_13391);
nor U14223 (N_14223,N_12397,N_12569);
and U14224 (N_14224,N_12761,N_12222);
nand U14225 (N_14225,N_12372,N_12947);
xor U14226 (N_14226,N_12057,N_13562);
nor U14227 (N_14227,N_12832,N_12349);
nand U14228 (N_14228,N_13172,N_13957);
nor U14229 (N_14229,N_12486,N_13230);
and U14230 (N_14230,N_13590,N_13743);
nand U14231 (N_14231,N_12117,N_12551);
and U14232 (N_14232,N_13337,N_13902);
or U14233 (N_14233,N_13070,N_13513);
and U14234 (N_14234,N_12283,N_12168);
and U14235 (N_14235,N_12116,N_12901);
or U14236 (N_14236,N_13754,N_12819);
nand U14237 (N_14237,N_12732,N_13682);
xor U14238 (N_14238,N_13868,N_13175);
nand U14239 (N_14239,N_12820,N_12447);
nor U14240 (N_14240,N_12622,N_13143);
nand U14241 (N_14241,N_13903,N_12964);
or U14242 (N_14242,N_12991,N_12870);
or U14243 (N_14243,N_12249,N_13159);
or U14244 (N_14244,N_12330,N_13899);
nor U14245 (N_14245,N_12690,N_13127);
or U14246 (N_14246,N_13254,N_12316);
nand U14247 (N_14247,N_12694,N_13459);
and U14248 (N_14248,N_13005,N_12675);
xnor U14249 (N_14249,N_13674,N_12318);
xnor U14250 (N_14250,N_12370,N_13823);
xnor U14251 (N_14251,N_12019,N_13853);
nand U14252 (N_14252,N_13841,N_13376);
xnor U14253 (N_14253,N_12080,N_12229);
nand U14254 (N_14254,N_13964,N_13825);
xor U14255 (N_14255,N_12271,N_13821);
or U14256 (N_14256,N_13685,N_13753);
nor U14257 (N_14257,N_13282,N_13665);
and U14258 (N_14258,N_12518,N_12233);
xnor U14259 (N_14259,N_12358,N_13656);
and U14260 (N_14260,N_13023,N_12210);
nor U14261 (N_14261,N_12952,N_13740);
nand U14262 (N_14262,N_12154,N_13885);
or U14263 (N_14263,N_12759,N_12488);
or U14264 (N_14264,N_12909,N_13527);
and U14265 (N_14265,N_12465,N_12376);
nand U14266 (N_14266,N_12184,N_12682);
and U14267 (N_14267,N_12163,N_13948);
or U14268 (N_14268,N_13542,N_13570);
nor U14269 (N_14269,N_12193,N_12572);
xnor U14270 (N_14270,N_13737,N_13752);
nand U14271 (N_14271,N_13194,N_12912);
xnor U14272 (N_14272,N_13267,N_12284);
nor U14273 (N_14273,N_13003,N_13613);
nand U14274 (N_14274,N_13007,N_12988);
xnor U14275 (N_14275,N_12309,N_13956);
nor U14276 (N_14276,N_12737,N_13691);
nor U14277 (N_14277,N_13789,N_13673);
nand U14278 (N_14278,N_13627,N_12454);
xnor U14279 (N_14279,N_13764,N_12788);
and U14280 (N_14280,N_12428,N_12869);
xnor U14281 (N_14281,N_12068,N_12113);
or U14282 (N_14282,N_12231,N_13822);
and U14283 (N_14283,N_12242,N_12110);
nor U14284 (N_14284,N_13924,N_13771);
or U14285 (N_14285,N_12801,N_13571);
xor U14286 (N_14286,N_12037,N_12328);
xnor U14287 (N_14287,N_13496,N_13179);
xnor U14288 (N_14288,N_12325,N_13756);
or U14289 (N_14289,N_12027,N_12907);
or U14290 (N_14290,N_12961,N_13488);
nand U14291 (N_14291,N_12941,N_13762);
xor U14292 (N_14292,N_12481,N_13765);
nand U14293 (N_14293,N_12388,N_13404);
and U14294 (N_14294,N_13881,N_12373);
nor U14295 (N_14295,N_13779,N_13412);
and U14296 (N_14296,N_13453,N_13932);
nor U14297 (N_14297,N_13848,N_13499);
xnor U14298 (N_14298,N_13467,N_13073);
or U14299 (N_14299,N_12698,N_13078);
xnor U14300 (N_14300,N_13537,N_12482);
xor U14301 (N_14301,N_12512,N_12054);
or U14302 (N_14302,N_12305,N_12836);
xor U14303 (N_14303,N_12262,N_12787);
nand U14304 (N_14304,N_12143,N_12290);
and U14305 (N_14305,N_12416,N_13361);
and U14306 (N_14306,N_13742,N_12701);
and U14307 (N_14307,N_13082,N_12379);
nor U14308 (N_14308,N_13300,N_13704);
nor U14309 (N_14309,N_13203,N_12195);
nand U14310 (N_14310,N_13336,N_12205);
nor U14311 (N_14311,N_12408,N_12437);
or U14312 (N_14312,N_12986,N_13583);
and U14313 (N_14313,N_12071,N_12711);
and U14314 (N_14314,N_12667,N_13100);
or U14315 (N_14315,N_12748,N_12435);
and U14316 (N_14316,N_13965,N_12916);
or U14317 (N_14317,N_13864,N_12338);
nor U14318 (N_14318,N_13534,N_13911);
or U14319 (N_14319,N_13977,N_12226);
nand U14320 (N_14320,N_13598,N_13797);
nand U14321 (N_14321,N_13454,N_12219);
nand U14322 (N_14322,N_12431,N_12829);
nand U14323 (N_14323,N_13287,N_13124);
and U14324 (N_14324,N_12521,N_12502);
or U14325 (N_14325,N_13597,N_13901);
or U14326 (N_14326,N_12046,N_13263);
or U14327 (N_14327,N_12064,N_13947);
nand U14328 (N_14328,N_13405,N_12250);
nor U14329 (N_14329,N_13156,N_12606);
nand U14330 (N_14330,N_12135,N_13374);
xnor U14331 (N_14331,N_12382,N_12570);
or U14332 (N_14332,N_13435,N_13451);
nand U14333 (N_14333,N_13476,N_12585);
or U14334 (N_14334,N_12995,N_13227);
and U14335 (N_14335,N_13411,N_12705);
or U14336 (N_14336,N_13788,N_13681);
and U14337 (N_14337,N_12496,N_12735);
or U14338 (N_14338,N_12898,N_12187);
or U14339 (N_14339,N_13763,N_13271);
or U14340 (N_14340,N_13283,N_13636);
or U14341 (N_14341,N_12843,N_13371);
and U14342 (N_14342,N_12519,N_12464);
or U14343 (N_14343,N_12746,N_13505);
or U14344 (N_14344,N_13973,N_12673);
and U14345 (N_14345,N_13538,N_12056);
and U14346 (N_14346,N_13168,N_12620);
or U14347 (N_14347,N_13877,N_13442);
xnor U14348 (N_14348,N_13623,N_13192);
xnor U14349 (N_14349,N_12074,N_13781);
or U14350 (N_14350,N_12560,N_12576);
nor U14351 (N_14351,N_13353,N_13676);
nand U14352 (N_14352,N_13133,N_13824);
nor U14353 (N_14353,N_13138,N_13044);
and U14354 (N_14354,N_12378,N_13326);
xnor U14355 (N_14355,N_13579,N_13926);
or U14356 (N_14356,N_13362,N_12272);
xor U14357 (N_14357,N_12149,N_12087);
or U14358 (N_14358,N_13091,N_12086);
or U14359 (N_14359,N_13528,N_12532);
and U14360 (N_14360,N_13354,N_12510);
or U14361 (N_14361,N_12173,N_13975);
nand U14362 (N_14362,N_13046,N_12180);
xor U14363 (N_14363,N_13128,N_12153);
nor U14364 (N_14364,N_12880,N_12830);
xnor U14365 (N_14365,N_12256,N_13251);
nor U14366 (N_14366,N_12783,N_12523);
nand U14367 (N_14367,N_12553,N_13184);
and U14368 (N_14368,N_13861,N_13639);
nand U14369 (N_14369,N_12157,N_12963);
xnor U14370 (N_14370,N_13777,N_13608);
nand U14371 (N_14371,N_12723,N_13152);
nor U14372 (N_14372,N_12505,N_12865);
xor U14373 (N_14373,N_13540,N_12939);
or U14374 (N_14374,N_12794,N_13306);
or U14375 (N_14375,N_12800,N_13061);
nand U14376 (N_14376,N_13847,N_13862);
nor U14377 (N_14377,N_13385,N_13804);
xnor U14378 (N_14378,N_12555,N_13027);
nand U14379 (N_14379,N_12903,N_12300);
nand U14380 (N_14380,N_12769,N_12756);
nor U14381 (N_14381,N_13778,N_13835);
xor U14382 (N_14382,N_13401,N_12319);
and U14383 (N_14383,N_12921,N_12013);
nand U14384 (N_14384,N_12299,N_12208);
nor U14385 (N_14385,N_13557,N_12619);
nand U14386 (N_14386,N_13461,N_12695);
and U14387 (N_14387,N_12517,N_13698);
xor U14388 (N_14388,N_12595,N_12857);
or U14389 (N_14389,N_12806,N_13483);
and U14390 (N_14390,N_12000,N_13437);
and U14391 (N_14391,N_12289,N_13011);
and U14392 (N_14392,N_12090,N_13360);
or U14393 (N_14393,N_12578,N_13766);
or U14394 (N_14394,N_13761,N_12334);
xnor U14395 (N_14395,N_13896,N_13275);
or U14396 (N_14396,N_13760,N_12324);
nor U14397 (N_14397,N_12894,N_12381);
nand U14398 (N_14398,N_13272,N_12717);
nand U14399 (N_14399,N_13849,N_12396);
or U14400 (N_14400,N_13288,N_12033);
xor U14401 (N_14401,N_13056,N_12323);
or U14402 (N_14402,N_12942,N_13009);
nor U14403 (N_14403,N_12767,N_12236);
xnor U14404 (N_14404,N_12198,N_13436);
xnor U14405 (N_14405,N_12725,N_13890);
or U14406 (N_14406,N_13626,N_12879);
xor U14407 (N_14407,N_13052,N_12878);
or U14408 (N_14408,N_13291,N_12047);
and U14409 (N_14409,N_13594,N_13149);
xnor U14410 (N_14410,N_13573,N_13615);
and U14411 (N_14411,N_12720,N_12839);
or U14412 (N_14412,N_13358,N_12105);
and U14413 (N_14413,N_12266,N_12383);
nor U14414 (N_14414,N_13745,N_12185);
and U14415 (N_14415,N_12457,N_13565);
xnor U14416 (N_14416,N_12647,N_12776);
or U14417 (N_14417,N_13637,N_13805);
nand U14418 (N_14418,N_13065,N_13578);
xor U14419 (N_14419,N_13738,N_12085);
or U14420 (N_14420,N_13099,N_13572);
xor U14421 (N_14421,N_13040,N_12474);
nor U14422 (N_14422,N_12132,N_13338);
and U14423 (N_14423,N_13920,N_12270);
and U14424 (N_14424,N_13077,N_12782);
xor U14425 (N_14425,N_12676,N_12312);
or U14426 (N_14426,N_12101,N_12966);
xnor U14427 (N_14427,N_13111,N_13662);
and U14428 (N_14428,N_13776,N_12221);
and U14429 (N_14429,N_12888,N_12743);
and U14430 (N_14430,N_12021,N_13974);
or U14431 (N_14431,N_12902,N_12344);
nand U14432 (N_14432,N_12763,N_13801);
xor U14433 (N_14433,N_12905,N_12082);
and U14434 (N_14434,N_12770,N_13262);
nor U14435 (N_14435,N_12337,N_12246);
or U14436 (N_14436,N_13851,N_13981);
nand U14437 (N_14437,N_13972,N_13515);
nand U14438 (N_14438,N_13464,N_13382);
or U14439 (N_14439,N_12684,N_13893);
nor U14440 (N_14440,N_12278,N_13687);
xor U14441 (N_14441,N_13575,N_13305);
or U14442 (N_14442,N_12020,N_12072);
or U14443 (N_14443,N_13342,N_13001);
and U14444 (N_14444,N_13871,N_13244);
nor U14445 (N_14445,N_13475,N_12491);
nand U14446 (N_14446,N_13116,N_13587);
xor U14447 (N_14447,N_12710,N_12392);
and U14448 (N_14448,N_12028,N_13620);
xor U14449 (N_14449,N_12815,N_12876);
and U14450 (N_14450,N_13517,N_12183);
nand U14451 (N_14451,N_12850,N_12131);
xnor U14452 (N_14452,N_13699,N_12308);
xor U14453 (N_14453,N_13285,N_12120);
and U14454 (N_14454,N_12421,N_13208);
xor U14455 (N_14455,N_13101,N_12680);
nor U14456 (N_14456,N_12969,N_12473);
nand U14457 (N_14457,N_12548,N_12932);
nand U14458 (N_14458,N_12703,N_12608);
and U14459 (N_14459,N_12536,N_13399);
nor U14460 (N_14460,N_12599,N_12121);
and U14461 (N_14461,N_13508,N_13631);
nor U14462 (N_14462,N_13880,N_12471);
nor U14463 (N_14463,N_12638,N_13799);
nor U14464 (N_14464,N_13739,N_12343);
and U14465 (N_14465,N_13955,N_12825);
and U14466 (N_14466,N_12683,N_13599);
nor U14467 (N_14467,N_12458,N_12045);
or U14468 (N_14468,N_12133,N_12594);
xor U14469 (N_14469,N_12405,N_12257);
or U14470 (N_14470,N_12707,N_12547);
or U14471 (N_14471,N_13794,N_12251);
nor U14472 (N_14472,N_13495,N_13158);
or U14473 (N_14473,N_13774,N_12484);
and U14474 (N_14474,N_13616,N_13939);
nor U14475 (N_14475,N_12529,N_12199);
nor U14476 (N_14476,N_13484,N_12384);
nor U14477 (N_14477,N_13109,N_13006);
xor U14478 (N_14478,N_13567,N_12862);
xor U14479 (N_14479,N_13525,N_12433);
nor U14480 (N_14480,N_12348,N_12182);
nand U14481 (N_14481,N_13480,N_13471);
and U14482 (N_14482,N_12639,N_12018);
nand U14483 (N_14483,N_13249,N_13869);
xnor U14484 (N_14484,N_13443,N_12461);
xnor U14485 (N_14485,N_12094,N_13845);
or U14486 (N_14486,N_13606,N_12220);
and U14487 (N_14487,N_13934,N_13700);
or U14488 (N_14488,N_13730,N_13148);
nor U14489 (N_14489,N_13482,N_12811);
nand U14490 (N_14490,N_13735,N_13104);
or U14491 (N_14491,N_12978,N_12719);
nor U14492 (N_14492,N_13373,N_13294);
xor U14493 (N_14493,N_12407,N_13812);
and U14494 (N_14494,N_12893,N_12773);
or U14495 (N_14495,N_12592,N_12010);
or U14496 (N_14496,N_12970,N_13970);
nor U14497 (N_14497,N_12012,N_13512);
or U14498 (N_14498,N_13072,N_13678);
nor U14499 (N_14499,N_12425,N_13102);
and U14500 (N_14500,N_12336,N_13566);
nor U14501 (N_14501,N_13402,N_12342);
and U14502 (N_14502,N_12738,N_12008);
xnor U14503 (N_14503,N_12494,N_12749);
xnor U14504 (N_14504,N_13671,N_12716);
xnor U14505 (N_14505,N_13322,N_12129);
or U14506 (N_14506,N_12634,N_12734);
xnor U14507 (N_14507,N_12394,N_12432);
nand U14508 (N_14508,N_13942,N_12586);
nand U14509 (N_14509,N_12398,N_13171);
or U14510 (N_14510,N_12333,N_13201);
or U14511 (N_14511,N_12573,N_12030);
xor U14512 (N_14512,N_12722,N_12861);
nor U14513 (N_14513,N_12403,N_12877);
xnor U14514 (N_14514,N_13195,N_12874);
and U14515 (N_14515,N_13241,N_13191);
and U14516 (N_14516,N_13132,N_12564);
xnor U14517 (N_14517,N_12042,N_12899);
nor U14518 (N_14518,N_12279,N_12530);
nand U14519 (N_14519,N_12713,N_12842);
or U14520 (N_14520,N_12439,N_13919);
or U14521 (N_14521,N_13466,N_12371);
nand U14522 (N_14522,N_12546,N_13004);
xor U14523 (N_14523,N_13870,N_12636);
xnor U14524 (N_14524,N_12652,N_12377);
and U14525 (N_14525,N_12002,N_12808);
or U14526 (N_14526,N_13428,N_13960);
nor U14527 (N_14527,N_12445,N_12785);
and U14528 (N_14528,N_13348,N_13239);
nor U14529 (N_14529,N_13692,N_12051);
xnor U14530 (N_14530,N_12951,N_12851);
nand U14531 (N_14531,N_12793,N_13295);
or U14532 (N_14532,N_13624,N_12616);
or U14533 (N_14533,N_13137,N_13093);
and U14534 (N_14534,N_12130,N_13221);
and U14535 (N_14535,N_12123,N_13058);
nor U14536 (N_14536,N_13876,N_12468);
and U14537 (N_14537,N_13830,N_13632);
and U14538 (N_14538,N_12446,N_13649);
or U14539 (N_14539,N_13544,N_12245);
or U14540 (N_14540,N_13548,N_12814);
or U14541 (N_14541,N_12538,N_13039);
or U14542 (N_14542,N_13859,N_13906);
nor U14543 (N_14543,N_12412,N_13438);
or U14544 (N_14544,N_12192,N_12115);
nor U14545 (N_14545,N_13087,N_12419);
or U14546 (N_14546,N_12061,N_13240);
nand U14547 (N_14547,N_13874,N_12657);
nor U14548 (N_14548,N_13126,N_13330);
nand U14549 (N_14549,N_13635,N_13486);
nand U14550 (N_14550,N_12659,N_13793);
nor U14551 (N_14551,N_13922,N_13481);
nand U14552 (N_14552,N_13601,N_13439);
nor U14553 (N_14553,N_13994,N_13551);
nor U14554 (N_14554,N_12356,N_12792);
and U14555 (N_14555,N_13029,N_12346);
and U14556 (N_14556,N_13315,N_13983);
nor U14557 (N_14557,N_12363,N_13460);
xor U14558 (N_14558,N_13214,N_13520);
and U14559 (N_14559,N_13524,N_12936);
or U14560 (N_14560,N_12844,N_13680);
nand U14561 (N_14561,N_13393,N_13751);
and U14562 (N_14562,N_12609,N_12228);
xnor U14563 (N_14563,N_12327,N_12075);
nor U14564 (N_14564,N_13406,N_13634);
xor U14565 (N_14565,N_12753,N_13638);
nand U14566 (N_14566,N_13654,N_12189);
and U14567 (N_14567,N_12812,N_12354);
or U14568 (N_14568,N_12672,N_13539);
nor U14569 (N_14569,N_12919,N_12114);
and U14570 (N_14570,N_13289,N_12320);
or U14571 (N_14571,N_12668,N_12810);
nand U14572 (N_14572,N_13036,N_12562);
nor U14573 (N_14573,N_13997,N_12817);
and U14574 (N_14574,N_12859,N_12615);
and U14575 (N_14575,N_13064,N_12999);
or U14576 (N_14576,N_13759,N_13213);
nand U14577 (N_14577,N_12345,N_12453);
xnor U14578 (N_14578,N_12718,N_13677);
or U14579 (N_14579,N_12727,N_13232);
nand U14580 (N_14580,N_12871,N_13695);
nor U14581 (N_14581,N_13817,N_13013);
xnor U14582 (N_14582,N_13324,N_13908);
nor U14583 (N_14583,N_12509,N_13840);
nand U14584 (N_14584,N_13560,N_13487);
xor U14585 (N_14585,N_12007,N_12216);
nand U14586 (N_14586,N_13519,N_12558);
nor U14587 (N_14587,N_13396,N_12460);
nand U14588 (N_14588,N_12165,N_12449);
and U14589 (N_14589,N_12200,N_12884);
xnor U14590 (N_14590,N_13931,N_12882);
and U14591 (N_14591,N_12689,N_13883);
and U14592 (N_14592,N_12190,N_12103);
nand U14593 (N_14593,N_13558,N_13605);
xnor U14594 (N_14594,N_13952,N_13923);
and U14595 (N_14595,N_12240,N_13842);
and U14596 (N_14596,N_12456,N_13860);
or U14597 (N_14597,N_13648,N_13433);
and U14598 (N_14598,N_12016,N_12241);
nor U14599 (N_14599,N_12011,N_13043);
xnor U14600 (N_14600,N_13302,N_12364);
or U14601 (N_14601,N_13492,N_12847);
nor U14602 (N_14602,N_12833,N_13543);
nor U14603 (N_14603,N_12297,N_13020);
nand U14604 (N_14604,N_12805,N_13386);
nand U14605 (N_14605,N_12938,N_12261);
xor U14606 (N_14606,N_13904,N_13554);
xnor U14607 (N_14607,N_13418,N_12708);
and U14608 (N_14608,N_13278,N_13219);
or U14609 (N_14609,N_12700,N_13141);
or U14610 (N_14610,N_13266,N_13652);
nor U14611 (N_14611,N_13530,N_13334);
nor U14612 (N_14612,N_12790,N_12539);
nor U14613 (N_14613,N_13086,N_12177);
xor U14614 (N_14614,N_13022,N_12426);
nand U14615 (N_14615,N_13060,N_13408);
nor U14616 (N_14616,N_12873,N_12968);
xor U14617 (N_14617,N_13501,N_13916);
nand U14618 (N_14618,N_12109,N_13837);
nor U14619 (N_14619,N_13600,N_12937);
and U14620 (N_14620,N_12544,N_13915);
nor U14621 (N_14621,N_13062,N_13693);
xor U14622 (N_14622,N_13253,N_12757);
nand U14623 (N_14623,N_12303,N_12739);
nor U14624 (N_14624,N_13274,N_13318);
and U14625 (N_14625,N_13657,N_13910);
nor U14626 (N_14626,N_13369,N_13129);
xor U14627 (N_14627,N_12014,N_13547);
nor U14628 (N_14628,N_12025,N_12664);
xnor U14629 (N_14629,N_13729,N_13782);
nor U14630 (N_14630,N_12107,N_12292);
and U14631 (N_14631,N_12036,N_12687);
and U14632 (N_14632,N_13585,N_13242);
xnor U14633 (N_14633,N_13323,N_13415);
nor U14634 (N_14634,N_12301,N_13593);
nand U14635 (N_14635,N_13045,N_13758);
xor U14636 (N_14636,N_13423,N_12083);
or U14637 (N_14637,N_12314,N_12145);
or U14638 (N_14638,N_12528,N_12041);
nand U14639 (N_14639,N_13341,N_13270);
or U14640 (N_14640,N_13356,N_12601);
and U14641 (N_14641,N_13290,N_13617);
or U14642 (N_14642,N_13033,N_12838);
nand U14643 (N_14643,N_12239,N_12522);
or U14644 (N_14644,N_12285,N_12477);
and U14645 (N_14645,N_13145,N_13992);
nand U14646 (N_14646,N_13686,N_13407);
or U14647 (N_14647,N_12495,N_13331);
xor U14648 (N_14648,N_13816,N_13712);
nor U14649 (N_14649,N_13344,N_12867);
nand U14650 (N_14650,N_12158,N_12933);
or U14651 (N_14651,N_12026,N_12775);
or U14652 (N_14652,N_13395,N_12666);
nand U14653 (N_14653,N_12691,N_13629);
xnor U14654 (N_14654,N_13311,N_12006);
or U14655 (N_14655,N_13647,N_12275);
xnor U14656 (N_14656,N_13211,N_12625);
or U14657 (N_14657,N_13688,N_13802);
nand U14658 (N_14658,N_12582,N_13935);
or U14659 (N_14659,N_13588,N_13990);
nor U14660 (N_14660,N_12048,N_13094);
and U14661 (N_14661,N_13403,N_12404);
and U14662 (N_14662,N_12993,N_13568);
xor U14663 (N_14663,N_12059,N_12563);
or U14664 (N_14664,N_13536,N_12678);
xnor U14665 (N_14665,N_12696,N_12076);
nor U14666 (N_14666,N_12179,N_13422);
nand U14667 (N_14667,N_13574,N_13803);
nor U14668 (N_14668,N_12589,N_13301);
xnor U14669 (N_14669,N_12784,N_13719);
nor U14670 (N_14670,N_13226,N_13328);
or U14671 (N_14671,N_13177,N_13655);
nor U14672 (N_14672,N_13982,N_12602);
or U14673 (N_14673,N_13889,N_13150);
nor U14674 (N_14674,N_13703,N_13314);
and U14675 (N_14675,N_12067,N_12611);
and U14676 (N_14676,N_13265,N_13448);
nor U14677 (N_14677,N_12733,N_12807);
or U14678 (N_14678,N_13958,N_12681);
xor U14679 (N_14679,N_13012,N_13489);
nand U14680 (N_14680,N_12875,N_13790);
xnor U14681 (N_14681,N_13084,N_13732);
and U14682 (N_14682,N_13545,N_13016);
nor U14683 (N_14683,N_12399,N_12411);
and U14684 (N_14684,N_12554,N_12144);
nand U14685 (N_14685,N_12934,N_12413);
nand U14686 (N_14686,N_13357,N_12335);
xnor U14687 (N_14687,N_12750,N_13791);
xor U14688 (N_14688,N_13419,N_13463);
nor U14689 (N_14689,N_12339,N_13755);
and U14690 (N_14690,N_12618,N_13961);
or U14691 (N_14691,N_12663,N_13727);
or U14692 (N_14692,N_12754,N_13609);
xnor U14693 (N_14693,N_13944,N_13098);
and U14694 (N_14694,N_13552,N_13553);
nand U14695 (N_14695,N_13940,N_12828);
or U14696 (N_14696,N_13335,N_13182);
nand U14697 (N_14697,N_12174,N_13731);
and U14698 (N_14698,N_13122,N_12766);
and U14699 (N_14699,N_12604,N_12079);
nand U14700 (N_14700,N_13279,N_13346);
nand U14701 (N_14701,N_12627,N_13260);
nor U14702 (N_14702,N_13347,N_12744);
and U14703 (N_14703,N_12516,N_13085);
and U14704 (N_14704,N_13954,N_12946);
or U14705 (N_14705,N_12629,N_13351);
or U14706 (N_14706,N_12864,N_13074);
and U14707 (N_14707,N_13991,N_13352);
nor U14708 (N_14708,N_13667,N_13092);
or U14709 (N_14709,N_13966,N_12058);
xnor U14710 (N_14710,N_13989,N_13746);
nand U14711 (N_14711,N_13710,N_13498);
nor U14712 (N_14712,N_12922,N_13720);
nand U14713 (N_14713,N_13397,N_13455);
and U14714 (N_14714,N_13689,N_12360);
xnor U14715 (N_14715,N_13008,N_12930);
or U14716 (N_14716,N_12568,N_12906);
and U14717 (N_14717,N_13670,N_13350);
nand U14718 (N_14718,N_12626,N_12765);
nor U14719 (N_14719,N_13409,N_12574);
and U14720 (N_14720,N_13810,N_12662);
xor U14721 (N_14721,N_13026,N_12927);
nor U14722 (N_14722,N_12699,N_13441);
nor U14723 (N_14723,N_13815,N_12957);
xnor U14724 (N_14724,N_13178,N_13205);
xor U14725 (N_14725,N_12591,N_13526);
or U14726 (N_14726,N_13160,N_13387);
xnor U14727 (N_14727,N_13933,N_12593);
and U14728 (N_14728,N_13229,N_12227);
and U14729 (N_14729,N_12575,N_12409);
xnor U14730 (N_14730,N_12612,N_13217);
xnor U14731 (N_14731,N_12206,N_13196);
nor U14732 (N_14732,N_12023,N_12571);
or U14733 (N_14733,N_13917,N_12224);
or U14734 (N_14734,N_13462,N_13813);
nand U14735 (N_14735,N_12994,N_12654);
xnor U14736 (N_14736,N_12982,N_13709);
and U14737 (N_14737,N_13032,N_13277);
nand U14738 (N_14738,N_12531,N_12863);
nand U14739 (N_14739,N_12535,N_12276);
nand U14740 (N_14740,N_12953,N_13839);
nor U14741 (N_14741,N_13445,N_13050);
and U14742 (N_14742,N_12146,N_13985);
xnor U14743 (N_14743,N_12485,N_13969);
xnor U14744 (N_14744,N_12891,N_12430);
and U14745 (N_14745,N_13118,N_13416);
xnor U14746 (N_14746,N_12162,N_12552);
or U14747 (N_14747,N_12781,N_13697);
or U14748 (N_14748,N_12442,N_13836);
and U14749 (N_14749,N_12498,N_12258);
or U14750 (N_14750,N_13478,N_13728);
xor U14751 (N_14751,N_13224,N_12704);
nand U14752 (N_14752,N_13456,N_12900);
and U14753 (N_14753,N_13549,N_13134);
or U14754 (N_14754,N_13928,N_13000);
and U14755 (N_14755,N_13749,N_13807);
nand U14756 (N_14756,N_12139,N_12452);
xnor U14757 (N_14757,N_12005,N_13963);
and U14758 (N_14758,N_13873,N_13504);
nand U14759 (N_14759,N_12996,N_12081);
or U14760 (N_14760,N_13041,N_12427);
nand U14761 (N_14761,N_13999,N_12660);
nand U14762 (N_14762,N_13978,N_13533);
nor U14763 (N_14763,N_12295,N_13702);
or U14764 (N_14764,N_13042,N_12053);
and U14765 (N_14765,N_12665,N_12225);
xor U14766 (N_14766,N_13716,N_12194);
and U14767 (N_14767,N_12914,N_13268);
nor U14768 (N_14768,N_12302,N_13907);
and U14769 (N_14769,N_12366,N_13392);
xnor U14770 (N_14770,N_12483,N_12213);
or U14771 (N_14771,N_13621,N_12127);
and U14772 (N_14772,N_13449,N_13225);
or U14773 (N_14773,N_13979,N_13115);
or U14774 (N_14774,N_12091,N_12017);
nor U14775 (N_14775,N_13663,N_13228);
or U14776 (N_14776,N_13207,N_13509);
nand U14777 (N_14777,N_13622,N_13153);
and U14778 (N_14778,N_12655,N_13139);
and U14779 (N_14779,N_12134,N_12935);
nand U14780 (N_14780,N_13198,N_12218);
or U14781 (N_14781,N_12697,N_12715);
nor U14782 (N_14782,N_12777,N_12998);
xor U14783 (N_14783,N_13892,N_13319);
xor U14784 (N_14784,N_13028,N_13136);
nand U14785 (N_14785,N_13485,N_12976);
xnor U14786 (N_14786,N_13340,N_13586);
nor U14787 (N_14787,N_13174,N_12353);
nand U14788 (N_14788,N_13325,N_13367);
nand U14789 (N_14789,N_13048,N_13707);
and U14790 (N_14790,N_12138,N_12467);
nor U14791 (N_14791,N_12632,N_12092);
nand U14792 (N_14792,N_12475,N_12063);
nor U14793 (N_14793,N_12977,N_12444);
nand U14794 (N_14794,N_13030,N_13912);
nand U14795 (N_14795,N_13364,N_13183);
and U14796 (N_14796,N_12096,N_13095);
nor U14797 (N_14797,N_13650,N_12556);
and U14798 (N_14798,N_13024,N_12728);
nor U14799 (N_14799,N_12462,N_12500);
nand U14800 (N_14800,N_12171,N_12848);
and U14801 (N_14801,N_12122,N_13281);
xor U14802 (N_14802,N_13246,N_13796);
xor U14803 (N_14803,N_13332,N_13611);
nand U14804 (N_14804,N_12253,N_12881);
xnor U14805 (N_14805,N_13380,N_12108);
nand U14806 (N_14806,N_12630,N_13711);
xor U14807 (N_14807,N_13014,N_12540);
and U14808 (N_14808,N_12099,N_13212);
or U14809 (N_14809,N_12669,N_13493);
xor U14810 (N_14810,N_13576,N_13097);
or U14811 (N_14811,N_13474,N_12613);
or U14812 (N_14812,N_13658,N_12747);
nor U14813 (N_14813,N_13581,N_12803);
nor U14814 (N_14814,N_13950,N_12979);
nor U14815 (N_14815,N_12924,N_13220);
xor U14816 (N_14816,N_13383,N_12989);
or U14817 (N_14817,N_13264,N_13987);
or U14818 (N_14818,N_12714,N_12291);
nor U14819 (N_14819,N_12992,N_12422);
nor U14820 (N_14820,N_13355,N_12908);
nand U14821 (N_14821,N_12679,N_12386);
nor U14822 (N_14822,N_13432,N_13866);
and U14823 (N_14823,N_13273,N_13798);
and U14824 (N_14824,N_12758,N_12326);
or U14825 (N_14825,N_12600,N_12268);
or U14826 (N_14826,N_13345,N_13772);
and U14827 (N_14827,N_13276,N_12196);
xor U14828 (N_14828,N_12674,N_13215);
or U14829 (N_14829,N_13664,N_12188);
or U14830 (N_14830,N_12692,N_13444);
and U14831 (N_14831,N_12401,N_13125);
nor U14832 (N_14832,N_13683,N_12885);
xor U14833 (N_14833,N_13169,N_13792);
and U14834 (N_14834,N_13017,N_13193);
and U14835 (N_14835,N_13814,N_12779);
and U14836 (N_14836,N_12648,N_12628);
xor U14837 (N_14837,N_13993,N_12052);
xor U14838 (N_14838,N_13834,N_12709);
and U14839 (N_14839,N_13114,N_13021);
nand U14840 (N_14840,N_12043,N_12472);
nor U14841 (N_14841,N_12489,N_13787);
or U14842 (N_14842,N_13218,N_12997);
nor U14843 (N_14843,N_13725,N_12417);
or U14844 (N_14844,N_12559,N_12824);
and U14845 (N_14845,N_13668,N_13468);
nor U14846 (N_14846,N_12588,N_13057);
or U14847 (N_14847,N_12795,N_13858);
or U14848 (N_14848,N_13259,N_13516);
nor U14849 (N_14849,N_12985,N_12039);
xnor U14850 (N_14850,N_12972,N_13996);
xnor U14851 (N_14851,N_12940,N_12661);
xnor U14852 (N_14852,N_12470,N_12060);
and U14853 (N_14853,N_12923,N_12846);
or U14854 (N_14854,N_13826,N_12361);
nand U14855 (N_14855,N_12181,N_13898);
nor U14856 (N_14856,N_13414,N_13715);
nor U14857 (N_14857,N_13185,N_12883);
xor U14858 (N_14858,N_13106,N_13661);
or U14859 (N_14859,N_13757,N_12990);
or U14860 (N_14860,N_13430,N_12579);
nand U14861 (N_14861,N_13123,N_12742);
and U14862 (N_14862,N_13929,N_13806);
or U14863 (N_14863,N_12524,N_12387);
nand U14864 (N_14864,N_13666,N_12499);
xnor U14865 (N_14865,N_12304,N_13832);
and U14866 (N_14866,N_12515,N_12590);
or U14867 (N_14867,N_12463,N_13223);
or U14868 (N_14868,N_13819,N_13531);
nand U14869 (N_14869,N_12633,N_13307);
and U14870 (N_14870,N_13604,N_13867);
xnor U14871 (N_14871,N_12823,N_13838);
nand U14872 (N_14872,N_13809,N_12726);
xnor U14873 (N_14873,N_13394,N_13494);
and U14874 (N_14874,N_12357,N_13465);
nor U14875 (N_14875,N_12493,N_13962);
or U14876 (N_14876,N_12203,N_13105);
and U14877 (N_14877,N_12307,N_13855);
nand U14878 (N_14878,N_13400,N_13596);
nor U14879 (N_14879,N_12204,N_13199);
xor U14880 (N_14880,N_13076,N_12125);
and U14881 (N_14881,N_12925,N_13257);
nand U14882 (N_14882,N_13440,N_13984);
or U14883 (N_14883,N_13410,N_12350);
nor U14884 (N_14884,N_13343,N_13250);
nor U14885 (N_14885,N_13252,N_13518);
xnor U14886 (N_14886,N_13614,N_13142);
nand U14887 (N_14887,N_13930,N_12147);
nor U14888 (N_14888,N_13800,N_13786);
nand U14889 (N_14889,N_13312,N_13748);
and U14890 (N_14890,N_13775,N_12238);
xnor U14891 (N_14891,N_12049,N_12911);
nor U14892 (N_14892,N_12235,N_12136);
or U14893 (N_14893,N_12561,N_12009);
xnor U14894 (N_14894,N_13619,N_13672);
xor U14895 (N_14895,N_13381,N_12252);
and U14896 (N_14896,N_13523,N_13921);
nand U14897 (N_14897,N_12215,N_13284);
xnor U14898 (N_14898,N_13176,N_13675);
nand U14899 (N_14899,N_12293,N_13286);
nor U14900 (N_14900,N_13852,N_13071);
nand U14901 (N_14901,N_12347,N_13261);
or U14902 (N_14902,N_13995,N_12577);
xnor U14903 (N_14903,N_12106,N_13329);
and U14904 (N_14904,N_12637,N_12414);
or U14905 (N_14905,N_13090,N_12390);
nand U14906 (N_14906,N_13618,N_12745);
nor U14907 (N_14907,N_12566,N_13083);
or U14908 (N_14908,N_13378,N_13705);
or U14909 (N_14909,N_12849,N_13375);
nand U14910 (N_14910,N_12175,N_13887);
and U14911 (N_14911,N_13059,N_13147);
or U14912 (N_14912,N_12209,N_12504);
nor U14913 (N_14913,N_12621,N_12298);
and U14914 (N_14914,N_13446,N_12550);
xnor U14915 (N_14915,N_13425,N_12029);
nor U14916 (N_14916,N_13882,N_12073);
and U14917 (N_14917,N_12112,N_13363);
xor U14918 (N_14918,N_12375,N_12487);
nand U14919 (N_14919,N_12886,N_13541);
nand U14920 (N_14920,N_13872,N_12310);
xnor U14921 (N_14921,N_13079,N_13577);
xor U14922 (N_14922,N_12962,N_13269);
xnor U14923 (N_14923,N_12089,N_13309);
nor U14924 (N_14924,N_12044,N_12760);
or U14925 (N_14925,N_12780,N_12852);
nor U14926 (N_14926,N_12244,N_12038);
nor U14927 (N_14927,N_12469,N_12537);
nand U14928 (N_14928,N_13359,N_12755);
nor U14929 (N_14929,N_13569,N_12124);
nand U14930 (N_14930,N_13535,N_12945);
and U14931 (N_14931,N_12821,N_13643);
nor U14932 (N_14932,N_13049,N_13857);
xnor U14933 (N_14933,N_12868,N_13245);
or U14934 (N_14934,N_12126,N_13831);
or U14935 (N_14935,N_12004,N_12640);
nor U14936 (N_14936,N_12084,N_12834);
or U14937 (N_14937,N_12845,N_12065);
nor U14938 (N_14938,N_13532,N_12093);
nand U14939 (N_14939,N_12436,N_12069);
nand U14940 (N_14940,N_12264,N_13236);
nand U14941 (N_14941,N_13603,N_13424);
or U14942 (N_14942,N_12799,N_12926);
nand U14943 (N_14943,N_13189,N_13173);
and U14944 (N_14944,N_12148,N_13971);
nor U14945 (N_14945,N_13510,N_13721);
nor U14946 (N_14946,N_13447,N_12959);
nand U14947 (N_14947,N_13491,N_12156);
or U14948 (N_14948,N_12918,N_13909);
or U14949 (N_14949,N_13140,N_12984);
nand U14950 (N_14950,N_12853,N_12954);
and U14951 (N_14951,N_13155,N_12492);
nor U14952 (N_14952,N_13210,N_13377);
xor U14953 (N_14953,N_12234,N_13784);
nand U14954 (N_14954,N_13157,N_12104);
xor U14955 (N_14955,N_13002,N_12223);
and U14956 (N_14956,N_12259,N_12827);
nand U14957 (N_14957,N_12910,N_13384);
nand U14958 (N_14958,N_13247,N_12466);
nor U14959 (N_14959,N_13706,N_13694);
nor U14960 (N_14960,N_12178,N_12736);
and U14961 (N_14961,N_13231,N_12050);
xnor U14962 (N_14962,N_13723,N_13063);
nor U14963 (N_14963,N_12443,N_13946);
or U14964 (N_14964,N_12286,N_13884);
and U14965 (N_14965,N_12230,N_13714);
nor U14966 (N_14966,N_12514,N_12649);
xnor U14967 (N_14967,N_12797,N_13998);
xnor U14968 (N_14968,N_12391,N_13696);
and U14969 (N_14969,N_13037,N_12434);
or U14970 (N_14970,N_12351,N_13827);
and U14971 (N_14971,N_12641,N_13081);
nand U14972 (N_14972,N_12913,N_12520);
or U14973 (N_14973,N_12527,N_13633);
xnor U14974 (N_14974,N_13256,N_12161);
or U14975 (N_14975,N_12677,N_13370);
and U14976 (N_14976,N_13398,N_12255);
xor U14977 (N_14977,N_13724,N_12974);
nor U14978 (N_14978,N_12804,N_13019);
xnor U14979 (N_14979,N_13477,N_12644);
xor U14980 (N_14980,N_12243,N_12478);
or U14981 (N_14981,N_13768,N_13941);
and U14982 (N_14982,N_13166,N_12288);
or U14983 (N_14983,N_13180,N_12406);
xor U14984 (N_14984,N_12650,N_13117);
or U14985 (N_14985,N_12693,N_13938);
and U14986 (N_14986,N_12506,N_13234);
or U14987 (N_14987,N_12610,N_13747);
xnor U14988 (N_14988,N_12031,N_13038);
nand U14989 (N_14989,N_13121,N_13119);
or U14990 (N_14990,N_13047,N_13167);
and U14991 (N_14991,N_13103,N_12451);
xor U14992 (N_14992,N_13031,N_12762);
nor U14993 (N_14993,N_12040,N_13365);
and U14994 (N_14994,N_12872,N_12513);
nor U14995 (N_14995,N_13120,N_13293);
or U14996 (N_14996,N_13546,N_13321);
nand U14997 (N_14997,N_13088,N_12866);
nor U14998 (N_14998,N_12459,N_13529);
nand U14999 (N_14999,N_12429,N_12771);
nor U15000 (N_15000,N_13078,N_13479);
or U15001 (N_15001,N_13569,N_13847);
and U15002 (N_15002,N_13701,N_13684);
and U15003 (N_15003,N_12634,N_12121);
nand U15004 (N_15004,N_12496,N_12597);
xor U15005 (N_15005,N_13390,N_12083);
and U15006 (N_15006,N_12998,N_12038);
nand U15007 (N_15007,N_12409,N_13297);
and U15008 (N_15008,N_13155,N_13941);
xor U15009 (N_15009,N_12278,N_12291);
xnor U15010 (N_15010,N_12644,N_12467);
nor U15011 (N_15011,N_13885,N_13304);
xnor U15012 (N_15012,N_12395,N_12633);
and U15013 (N_15013,N_12916,N_12314);
xnor U15014 (N_15014,N_12024,N_13722);
nand U15015 (N_15015,N_12955,N_13733);
xor U15016 (N_15016,N_12141,N_12296);
or U15017 (N_15017,N_13947,N_12542);
xnor U15018 (N_15018,N_13655,N_13870);
or U15019 (N_15019,N_12724,N_12330);
nor U15020 (N_15020,N_13672,N_12992);
and U15021 (N_15021,N_12508,N_13826);
xor U15022 (N_15022,N_13977,N_12443);
and U15023 (N_15023,N_13129,N_12350);
nor U15024 (N_15024,N_13046,N_12028);
or U15025 (N_15025,N_13580,N_13401);
or U15026 (N_15026,N_12089,N_13758);
nor U15027 (N_15027,N_12845,N_13090);
and U15028 (N_15028,N_13031,N_12360);
nor U15029 (N_15029,N_12682,N_12126);
or U15030 (N_15030,N_12995,N_12873);
xnor U15031 (N_15031,N_13656,N_12535);
and U15032 (N_15032,N_12159,N_13000);
nor U15033 (N_15033,N_12758,N_12692);
nand U15034 (N_15034,N_12726,N_12629);
and U15035 (N_15035,N_12436,N_13814);
and U15036 (N_15036,N_13789,N_13773);
and U15037 (N_15037,N_13774,N_13773);
and U15038 (N_15038,N_13345,N_13175);
or U15039 (N_15039,N_13452,N_13238);
xnor U15040 (N_15040,N_13777,N_12401);
and U15041 (N_15041,N_13975,N_13744);
and U15042 (N_15042,N_13915,N_13672);
xor U15043 (N_15043,N_12806,N_13520);
and U15044 (N_15044,N_12489,N_12445);
or U15045 (N_15045,N_13709,N_13100);
or U15046 (N_15046,N_13567,N_12825);
nand U15047 (N_15047,N_13953,N_13575);
nor U15048 (N_15048,N_12948,N_13713);
and U15049 (N_15049,N_12334,N_13916);
xnor U15050 (N_15050,N_13173,N_13812);
xnor U15051 (N_15051,N_13001,N_12756);
nand U15052 (N_15052,N_12503,N_13482);
and U15053 (N_15053,N_13410,N_13032);
and U15054 (N_15054,N_13761,N_12217);
xnor U15055 (N_15055,N_12899,N_12072);
nor U15056 (N_15056,N_12918,N_13818);
and U15057 (N_15057,N_12803,N_12992);
nor U15058 (N_15058,N_13768,N_13586);
nor U15059 (N_15059,N_12700,N_13674);
xnor U15060 (N_15060,N_13801,N_13042);
xor U15061 (N_15061,N_13467,N_12841);
and U15062 (N_15062,N_13506,N_13859);
and U15063 (N_15063,N_12105,N_12819);
nand U15064 (N_15064,N_13034,N_13710);
xnor U15065 (N_15065,N_12067,N_12589);
nor U15066 (N_15066,N_12837,N_13421);
nand U15067 (N_15067,N_12064,N_13193);
and U15068 (N_15068,N_12252,N_12491);
and U15069 (N_15069,N_12935,N_13474);
and U15070 (N_15070,N_13364,N_13898);
and U15071 (N_15071,N_12290,N_13270);
or U15072 (N_15072,N_13603,N_13811);
and U15073 (N_15073,N_13814,N_12948);
or U15074 (N_15074,N_13473,N_12956);
and U15075 (N_15075,N_12410,N_13176);
xor U15076 (N_15076,N_13015,N_13345);
xor U15077 (N_15077,N_13462,N_12224);
and U15078 (N_15078,N_13181,N_13318);
nand U15079 (N_15079,N_13267,N_13654);
nand U15080 (N_15080,N_12764,N_12906);
or U15081 (N_15081,N_13595,N_13817);
nor U15082 (N_15082,N_13695,N_13438);
xnor U15083 (N_15083,N_13005,N_13622);
and U15084 (N_15084,N_13366,N_12237);
xor U15085 (N_15085,N_12464,N_12601);
or U15086 (N_15086,N_12862,N_12655);
xnor U15087 (N_15087,N_12710,N_12489);
and U15088 (N_15088,N_12211,N_12150);
and U15089 (N_15089,N_13384,N_12727);
or U15090 (N_15090,N_13377,N_12235);
or U15091 (N_15091,N_13195,N_13150);
nand U15092 (N_15092,N_12043,N_13137);
nor U15093 (N_15093,N_12889,N_13948);
xor U15094 (N_15094,N_12836,N_13841);
xor U15095 (N_15095,N_13216,N_12200);
xor U15096 (N_15096,N_13576,N_12656);
and U15097 (N_15097,N_12474,N_13218);
xnor U15098 (N_15098,N_13349,N_12248);
nor U15099 (N_15099,N_12797,N_13010);
or U15100 (N_15100,N_12565,N_12466);
nor U15101 (N_15101,N_12447,N_13135);
nor U15102 (N_15102,N_13206,N_12328);
xor U15103 (N_15103,N_12565,N_13324);
nand U15104 (N_15104,N_13410,N_12148);
nand U15105 (N_15105,N_12362,N_13258);
xnor U15106 (N_15106,N_13319,N_12320);
nand U15107 (N_15107,N_12441,N_12231);
nand U15108 (N_15108,N_13695,N_12405);
and U15109 (N_15109,N_12439,N_12754);
nand U15110 (N_15110,N_13276,N_12575);
xnor U15111 (N_15111,N_12340,N_13084);
nor U15112 (N_15112,N_12269,N_12526);
or U15113 (N_15113,N_13791,N_12941);
xnor U15114 (N_15114,N_13103,N_12735);
or U15115 (N_15115,N_13999,N_12679);
or U15116 (N_15116,N_13493,N_12660);
nor U15117 (N_15117,N_12515,N_13005);
and U15118 (N_15118,N_13313,N_12151);
nor U15119 (N_15119,N_13949,N_12678);
nor U15120 (N_15120,N_13013,N_13931);
nor U15121 (N_15121,N_12815,N_13318);
nand U15122 (N_15122,N_12989,N_13302);
xor U15123 (N_15123,N_12233,N_12081);
or U15124 (N_15124,N_13552,N_13594);
or U15125 (N_15125,N_12456,N_12894);
nor U15126 (N_15126,N_12060,N_12327);
xnor U15127 (N_15127,N_12034,N_12411);
nor U15128 (N_15128,N_13880,N_13328);
xor U15129 (N_15129,N_12824,N_12282);
or U15130 (N_15130,N_12613,N_13434);
xor U15131 (N_15131,N_12012,N_13013);
nand U15132 (N_15132,N_13213,N_13300);
and U15133 (N_15133,N_12854,N_12524);
or U15134 (N_15134,N_13229,N_13536);
nor U15135 (N_15135,N_13446,N_12636);
nand U15136 (N_15136,N_13782,N_13913);
and U15137 (N_15137,N_13309,N_13429);
xor U15138 (N_15138,N_13402,N_13595);
xor U15139 (N_15139,N_12636,N_13618);
nor U15140 (N_15140,N_12264,N_12924);
nor U15141 (N_15141,N_13321,N_12086);
or U15142 (N_15142,N_13407,N_13348);
nand U15143 (N_15143,N_12466,N_13986);
or U15144 (N_15144,N_13825,N_12739);
nand U15145 (N_15145,N_12463,N_13576);
xnor U15146 (N_15146,N_12609,N_12258);
nor U15147 (N_15147,N_12599,N_13295);
xor U15148 (N_15148,N_13129,N_12514);
nand U15149 (N_15149,N_13637,N_13159);
and U15150 (N_15150,N_12708,N_13483);
xnor U15151 (N_15151,N_13103,N_12621);
xor U15152 (N_15152,N_13132,N_13048);
nor U15153 (N_15153,N_12745,N_13895);
or U15154 (N_15154,N_13914,N_12336);
or U15155 (N_15155,N_12185,N_13296);
nand U15156 (N_15156,N_12872,N_13950);
nand U15157 (N_15157,N_13414,N_12538);
and U15158 (N_15158,N_12237,N_12202);
nand U15159 (N_15159,N_13747,N_13443);
and U15160 (N_15160,N_12419,N_12014);
and U15161 (N_15161,N_13176,N_12961);
or U15162 (N_15162,N_12978,N_12435);
or U15163 (N_15163,N_13135,N_12114);
xnor U15164 (N_15164,N_13668,N_12743);
nor U15165 (N_15165,N_12630,N_13866);
xor U15166 (N_15166,N_12954,N_13438);
and U15167 (N_15167,N_13548,N_12647);
and U15168 (N_15168,N_12191,N_13030);
xor U15169 (N_15169,N_12805,N_13662);
and U15170 (N_15170,N_12020,N_12172);
xor U15171 (N_15171,N_12507,N_13760);
nand U15172 (N_15172,N_13968,N_12312);
nand U15173 (N_15173,N_12823,N_13152);
nand U15174 (N_15174,N_13474,N_13601);
nand U15175 (N_15175,N_13079,N_13331);
xnor U15176 (N_15176,N_13054,N_12681);
or U15177 (N_15177,N_13151,N_13101);
nand U15178 (N_15178,N_12359,N_12684);
xor U15179 (N_15179,N_12337,N_13989);
nor U15180 (N_15180,N_12466,N_12411);
xor U15181 (N_15181,N_13868,N_12168);
or U15182 (N_15182,N_12513,N_13667);
or U15183 (N_15183,N_12364,N_12273);
nor U15184 (N_15184,N_13663,N_12588);
xor U15185 (N_15185,N_13887,N_12160);
xor U15186 (N_15186,N_12062,N_13168);
xor U15187 (N_15187,N_12039,N_13350);
nor U15188 (N_15188,N_12652,N_13847);
nor U15189 (N_15189,N_13250,N_12368);
and U15190 (N_15190,N_13216,N_12378);
and U15191 (N_15191,N_13944,N_13926);
xor U15192 (N_15192,N_12261,N_12399);
or U15193 (N_15193,N_13772,N_12615);
nor U15194 (N_15194,N_13584,N_12780);
nand U15195 (N_15195,N_13974,N_12431);
nand U15196 (N_15196,N_13592,N_13775);
xor U15197 (N_15197,N_12697,N_12645);
xnor U15198 (N_15198,N_12853,N_13695);
nand U15199 (N_15199,N_12636,N_13184);
and U15200 (N_15200,N_13785,N_12660);
nand U15201 (N_15201,N_12897,N_13762);
nand U15202 (N_15202,N_13941,N_12948);
nand U15203 (N_15203,N_13274,N_13774);
xnor U15204 (N_15204,N_13000,N_13160);
nor U15205 (N_15205,N_13783,N_12644);
or U15206 (N_15206,N_12744,N_12366);
nand U15207 (N_15207,N_12766,N_13527);
xor U15208 (N_15208,N_12727,N_13032);
xnor U15209 (N_15209,N_13318,N_13523);
or U15210 (N_15210,N_12889,N_13537);
or U15211 (N_15211,N_13878,N_12935);
nand U15212 (N_15212,N_12922,N_13011);
xor U15213 (N_15213,N_13947,N_12351);
or U15214 (N_15214,N_12252,N_12302);
or U15215 (N_15215,N_13051,N_13241);
or U15216 (N_15216,N_13253,N_12233);
or U15217 (N_15217,N_13725,N_12724);
and U15218 (N_15218,N_12040,N_13665);
nor U15219 (N_15219,N_12265,N_12912);
xnor U15220 (N_15220,N_12705,N_12052);
nor U15221 (N_15221,N_12154,N_13819);
nor U15222 (N_15222,N_12290,N_13621);
and U15223 (N_15223,N_12653,N_12287);
and U15224 (N_15224,N_12937,N_13024);
and U15225 (N_15225,N_12892,N_12997);
or U15226 (N_15226,N_12297,N_12857);
nor U15227 (N_15227,N_12984,N_12089);
and U15228 (N_15228,N_12463,N_13618);
or U15229 (N_15229,N_12940,N_13071);
xor U15230 (N_15230,N_12446,N_13359);
and U15231 (N_15231,N_12416,N_13878);
or U15232 (N_15232,N_12644,N_13941);
nand U15233 (N_15233,N_12804,N_13951);
nor U15234 (N_15234,N_12790,N_12755);
nor U15235 (N_15235,N_13125,N_12186);
or U15236 (N_15236,N_13471,N_12460);
or U15237 (N_15237,N_12269,N_12978);
nand U15238 (N_15238,N_12439,N_13791);
xnor U15239 (N_15239,N_13232,N_12007);
or U15240 (N_15240,N_13989,N_13392);
nand U15241 (N_15241,N_12456,N_13220);
nor U15242 (N_15242,N_13471,N_12083);
nor U15243 (N_15243,N_13516,N_13521);
nand U15244 (N_15244,N_13305,N_12310);
xnor U15245 (N_15245,N_13964,N_13783);
or U15246 (N_15246,N_13629,N_13962);
xor U15247 (N_15247,N_12583,N_13738);
nor U15248 (N_15248,N_13479,N_12683);
and U15249 (N_15249,N_12870,N_13875);
nand U15250 (N_15250,N_13203,N_12956);
or U15251 (N_15251,N_13486,N_13820);
or U15252 (N_15252,N_12127,N_12552);
and U15253 (N_15253,N_12876,N_13240);
or U15254 (N_15254,N_12195,N_12610);
or U15255 (N_15255,N_13323,N_12825);
xor U15256 (N_15256,N_13629,N_12348);
or U15257 (N_15257,N_12349,N_13542);
and U15258 (N_15258,N_12154,N_13354);
nor U15259 (N_15259,N_13199,N_13066);
nor U15260 (N_15260,N_12964,N_12259);
nor U15261 (N_15261,N_12475,N_12938);
nand U15262 (N_15262,N_12215,N_12657);
nor U15263 (N_15263,N_13596,N_12133);
nand U15264 (N_15264,N_12385,N_13351);
and U15265 (N_15265,N_12568,N_12339);
and U15266 (N_15266,N_12796,N_13802);
nor U15267 (N_15267,N_13805,N_13745);
nand U15268 (N_15268,N_12154,N_13882);
xor U15269 (N_15269,N_12123,N_13675);
xnor U15270 (N_15270,N_13421,N_12793);
or U15271 (N_15271,N_12540,N_13235);
and U15272 (N_15272,N_12268,N_12672);
xnor U15273 (N_15273,N_13099,N_13648);
nand U15274 (N_15274,N_13286,N_12340);
and U15275 (N_15275,N_12693,N_12125);
nor U15276 (N_15276,N_12129,N_12134);
or U15277 (N_15277,N_13317,N_13278);
nor U15278 (N_15278,N_13036,N_12688);
and U15279 (N_15279,N_12255,N_13251);
xnor U15280 (N_15280,N_12139,N_12362);
xor U15281 (N_15281,N_13640,N_13759);
and U15282 (N_15282,N_13630,N_12660);
and U15283 (N_15283,N_13813,N_12498);
xnor U15284 (N_15284,N_13803,N_13662);
nor U15285 (N_15285,N_12315,N_12975);
xnor U15286 (N_15286,N_13020,N_12333);
and U15287 (N_15287,N_12150,N_12705);
nand U15288 (N_15288,N_12741,N_12822);
or U15289 (N_15289,N_13134,N_12909);
and U15290 (N_15290,N_12119,N_12897);
or U15291 (N_15291,N_13010,N_13740);
and U15292 (N_15292,N_13176,N_12087);
nor U15293 (N_15293,N_13945,N_13707);
nor U15294 (N_15294,N_13322,N_13787);
nor U15295 (N_15295,N_13256,N_13130);
nor U15296 (N_15296,N_12571,N_13098);
xor U15297 (N_15297,N_13035,N_13028);
nor U15298 (N_15298,N_13675,N_12747);
or U15299 (N_15299,N_12194,N_12786);
nor U15300 (N_15300,N_12353,N_13728);
nand U15301 (N_15301,N_13002,N_13276);
nor U15302 (N_15302,N_12520,N_12528);
or U15303 (N_15303,N_12148,N_12760);
xnor U15304 (N_15304,N_12883,N_12863);
xor U15305 (N_15305,N_13503,N_13459);
xor U15306 (N_15306,N_13955,N_13931);
nor U15307 (N_15307,N_12901,N_13876);
and U15308 (N_15308,N_13156,N_12527);
nor U15309 (N_15309,N_12997,N_12226);
xor U15310 (N_15310,N_12269,N_12083);
or U15311 (N_15311,N_12096,N_13600);
nand U15312 (N_15312,N_12264,N_13909);
xnor U15313 (N_15313,N_12427,N_12931);
xor U15314 (N_15314,N_13215,N_12877);
or U15315 (N_15315,N_13714,N_12430);
and U15316 (N_15316,N_13765,N_13138);
nand U15317 (N_15317,N_12447,N_13835);
nor U15318 (N_15318,N_12096,N_13940);
or U15319 (N_15319,N_13871,N_12289);
nand U15320 (N_15320,N_12984,N_12549);
xor U15321 (N_15321,N_12797,N_13667);
and U15322 (N_15322,N_12348,N_12534);
nor U15323 (N_15323,N_13406,N_12743);
nand U15324 (N_15324,N_12263,N_13143);
nand U15325 (N_15325,N_12203,N_12362);
and U15326 (N_15326,N_13367,N_12850);
or U15327 (N_15327,N_12140,N_12533);
nand U15328 (N_15328,N_13250,N_13008);
nor U15329 (N_15329,N_13499,N_13880);
nand U15330 (N_15330,N_13835,N_13305);
and U15331 (N_15331,N_13475,N_12726);
nand U15332 (N_15332,N_13079,N_12405);
nand U15333 (N_15333,N_13747,N_13116);
or U15334 (N_15334,N_13032,N_12781);
xor U15335 (N_15335,N_12330,N_13686);
xor U15336 (N_15336,N_13499,N_13817);
xnor U15337 (N_15337,N_12465,N_12500);
xnor U15338 (N_15338,N_12969,N_12331);
nand U15339 (N_15339,N_13060,N_12901);
nor U15340 (N_15340,N_13370,N_12636);
or U15341 (N_15341,N_12372,N_13924);
or U15342 (N_15342,N_12401,N_12032);
nor U15343 (N_15343,N_13767,N_12242);
and U15344 (N_15344,N_13161,N_13659);
xor U15345 (N_15345,N_13083,N_12382);
nand U15346 (N_15346,N_13100,N_12601);
xnor U15347 (N_15347,N_13361,N_13947);
or U15348 (N_15348,N_12767,N_12704);
xor U15349 (N_15349,N_13188,N_13523);
xnor U15350 (N_15350,N_12093,N_12933);
nand U15351 (N_15351,N_12551,N_12613);
nand U15352 (N_15352,N_12491,N_13099);
nor U15353 (N_15353,N_13993,N_13425);
xnor U15354 (N_15354,N_13054,N_13406);
xor U15355 (N_15355,N_13256,N_13717);
nand U15356 (N_15356,N_12498,N_13622);
and U15357 (N_15357,N_12025,N_13490);
nor U15358 (N_15358,N_13663,N_13863);
nand U15359 (N_15359,N_13905,N_12907);
or U15360 (N_15360,N_12902,N_12171);
xnor U15361 (N_15361,N_12552,N_13160);
nand U15362 (N_15362,N_13973,N_12017);
and U15363 (N_15363,N_13433,N_13111);
nor U15364 (N_15364,N_12527,N_12536);
xnor U15365 (N_15365,N_12850,N_13085);
or U15366 (N_15366,N_13170,N_12448);
nor U15367 (N_15367,N_12210,N_13333);
or U15368 (N_15368,N_13101,N_13820);
nor U15369 (N_15369,N_12244,N_13005);
nor U15370 (N_15370,N_13446,N_13281);
nand U15371 (N_15371,N_12695,N_13293);
nand U15372 (N_15372,N_12017,N_12235);
nand U15373 (N_15373,N_13269,N_12306);
and U15374 (N_15374,N_13063,N_13060);
or U15375 (N_15375,N_13953,N_12745);
or U15376 (N_15376,N_12215,N_13412);
or U15377 (N_15377,N_13961,N_13312);
xnor U15378 (N_15378,N_12944,N_13097);
or U15379 (N_15379,N_12819,N_12907);
or U15380 (N_15380,N_13801,N_13035);
and U15381 (N_15381,N_13557,N_13190);
and U15382 (N_15382,N_12034,N_12232);
nor U15383 (N_15383,N_13034,N_13468);
nand U15384 (N_15384,N_12065,N_12773);
nor U15385 (N_15385,N_13432,N_12762);
xor U15386 (N_15386,N_12937,N_12733);
and U15387 (N_15387,N_12613,N_13519);
and U15388 (N_15388,N_13036,N_13035);
or U15389 (N_15389,N_12142,N_12703);
nand U15390 (N_15390,N_13605,N_12896);
nor U15391 (N_15391,N_13560,N_13177);
and U15392 (N_15392,N_13292,N_12400);
nor U15393 (N_15393,N_13338,N_13259);
nand U15394 (N_15394,N_13847,N_13809);
or U15395 (N_15395,N_12642,N_12654);
xor U15396 (N_15396,N_12055,N_12814);
and U15397 (N_15397,N_13316,N_12316);
and U15398 (N_15398,N_12774,N_12088);
nor U15399 (N_15399,N_13933,N_13174);
or U15400 (N_15400,N_13991,N_13935);
nor U15401 (N_15401,N_13019,N_12278);
nand U15402 (N_15402,N_13585,N_13230);
and U15403 (N_15403,N_13556,N_12899);
or U15404 (N_15404,N_13577,N_12478);
nor U15405 (N_15405,N_13594,N_12886);
and U15406 (N_15406,N_13712,N_13300);
and U15407 (N_15407,N_13643,N_13237);
and U15408 (N_15408,N_13955,N_12724);
xnor U15409 (N_15409,N_13056,N_12768);
and U15410 (N_15410,N_12980,N_12068);
xnor U15411 (N_15411,N_12127,N_12007);
xnor U15412 (N_15412,N_13499,N_13868);
xor U15413 (N_15413,N_13427,N_13080);
or U15414 (N_15414,N_12942,N_12257);
or U15415 (N_15415,N_13806,N_13103);
xnor U15416 (N_15416,N_12310,N_13560);
and U15417 (N_15417,N_12346,N_13568);
xnor U15418 (N_15418,N_12546,N_13130);
nor U15419 (N_15419,N_12973,N_13677);
nand U15420 (N_15420,N_12304,N_12477);
and U15421 (N_15421,N_12632,N_13775);
or U15422 (N_15422,N_13232,N_13819);
xnor U15423 (N_15423,N_12823,N_12410);
nor U15424 (N_15424,N_12797,N_12966);
or U15425 (N_15425,N_13147,N_13963);
nor U15426 (N_15426,N_12189,N_13849);
or U15427 (N_15427,N_12415,N_13855);
nor U15428 (N_15428,N_13795,N_13002);
nand U15429 (N_15429,N_13074,N_12975);
nor U15430 (N_15430,N_13461,N_13826);
and U15431 (N_15431,N_12036,N_13912);
nor U15432 (N_15432,N_13255,N_12279);
nor U15433 (N_15433,N_13327,N_13646);
nand U15434 (N_15434,N_12718,N_12222);
and U15435 (N_15435,N_13481,N_13552);
and U15436 (N_15436,N_12277,N_12337);
nor U15437 (N_15437,N_12301,N_12758);
and U15438 (N_15438,N_13780,N_13421);
xnor U15439 (N_15439,N_13058,N_12627);
nor U15440 (N_15440,N_13434,N_13717);
nor U15441 (N_15441,N_12673,N_12192);
nor U15442 (N_15442,N_12362,N_13117);
and U15443 (N_15443,N_13182,N_13490);
or U15444 (N_15444,N_12985,N_12208);
nand U15445 (N_15445,N_13718,N_13150);
or U15446 (N_15446,N_13563,N_12358);
and U15447 (N_15447,N_12794,N_13212);
xor U15448 (N_15448,N_13114,N_12457);
nand U15449 (N_15449,N_12500,N_13318);
nand U15450 (N_15450,N_12178,N_12606);
or U15451 (N_15451,N_12706,N_13549);
and U15452 (N_15452,N_12187,N_13695);
nor U15453 (N_15453,N_13535,N_13942);
nand U15454 (N_15454,N_12723,N_13186);
and U15455 (N_15455,N_12698,N_13162);
and U15456 (N_15456,N_13953,N_13670);
or U15457 (N_15457,N_12734,N_12530);
nor U15458 (N_15458,N_13917,N_13192);
and U15459 (N_15459,N_13109,N_13038);
nor U15460 (N_15460,N_13195,N_12900);
nor U15461 (N_15461,N_13868,N_13515);
nor U15462 (N_15462,N_12737,N_12449);
and U15463 (N_15463,N_13110,N_13375);
xnor U15464 (N_15464,N_12402,N_12769);
nand U15465 (N_15465,N_12083,N_13982);
and U15466 (N_15466,N_12179,N_13114);
and U15467 (N_15467,N_12823,N_12775);
and U15468 (N_15468,N_13703,N_13546);
or U15469 (N_15469,N_12586,N_13624);
nor U15470 (N_15470,N_12945,N_12761);
and U15471 (N_15471,N_13133,N_12447);
nor U15472 (N_15472,N_12379,N_13346);
or U15473 (N_15473,N_12611,N_12653);
nand U15474 (N_15474,N_13146,N_13746);
nand U15475 (N_15475,N_12877,N_13808);
and U15476 (N_15476,N_12822,N_12927);
xor U15477 (N_15477,N_13833,N_13160);
nand U15478 (N_15478,N_12404,N_13250);
and U15479 (N_15479,N_12042,N_12693);
or U15480 (N_15480,N_13293,N_12200);
and U15481 (N_15481,N_13871,N_13323);
nand U15482 (N_15482,N_12119,N_12161);
nand U15483 (N_15483,N_13098,N_12712);
or U15484 (N_15484,N_13263,N_12357);
nand U15485 (N_15485,N_13129,N_13927);
xnor U15486 (N_15486,N_13797,N_13548);
or U15487 (N_15487,N_13086,N_13640);
xor U15488 (N_15488,N_13686,N_12518);
xnor U15489 (N_15489,N_12215,N_12413);
and U15490 (N_15490,N_12250,N_13686);
xnor U15491 (N_15491,N_12598,N_13915);
nand U15492 (N_15492,N_13674,N_13349);
and U15493 (N_15493,N_13330,N_13278);
and U15494 (N_15494,N_12867,N_13799);
or U15495 (N_15495,N_13184,N_12441);
xor U15496 (N_15496,N_12826,N_12229);
or U15497 (N_15497,N_13205,N_13839);
and U15498 (N_15498,N_13028,N_12844);
and U15499 (N_15499,N_12167,N_12633);
nand U15500 (N_15500,N_13741,N_12916);
xnor U15501 (N_15501,N_12002,N_13522);
or U15502 (N_15502,N_12723,N_12096);
nand U15503 (N_15503,N_13371,N_12181);
nand U15504 (N_15504,N_12192,N_13562);
nand U15505 (N_15505,N_12616,N_13106);
nor U15506 (N_15506,N_12005,N_12273);
nand U15507 (N_15507,N_13641,N_12062);
and U15508 (N_15508,N_13482,N_13874);
or U15509 (N_15509,N_12085,N_12342);
nor U15510 (N_15510,N_12248,N_12356);
xor U15511 (N_15511,N_12207,N_12390);
xnor U15512 (N_15512,N_12582,N_13810);
nor U15513 (N_15513,N_12113,N_13319);
nor U15514 (N_15514,N_12770,N_13129);
and U15515 (N_15515,N_12808,N_12529);
xnor U15516 (N_15516,N_13379,N_12949);
xnor U15517 (N_15517,N_13249,N_12892);
nor U15518 (N_15518,N_13150,N_12372);
and U15519 (N_15519,N_12718,N_12103);
and U15520 (N_15520,N_12452,N_12285);
xnor U15521 (N_15521,N_13653,N_13256);
xnor U15522 (N_15522,N_13140,N_13802);
or U15523 (N_15523,N_13314,N_12396);
xor U15524 (N_15524,N_13238,N_12642);
nor U15525 (N_15525,N_12365,N_13021);
or U15526 (N_15526,N_12122,N_13656);
nor U15527 (N_15527,N_12865,N_12722);
and U15528 (N_15528,N_12508,N_13768);
nor U15529 (N_15529,N_13881,N_12123);
xor U15530 (N_15530,N_12388,N_13974);
nor U15531 (N_15531,N_13550,N_13912);
and U15532 (N_15532,N_13512,N_12502);
xnor U15533 (N_15533,N_13954,N_13701);
nor U15534 (N_15534,N_12624,N_12830);
xnor U15535 (N_15535,N_12509,N_13082);
xor U15536 (N_15536,N_13012,N_12677);
xnor U15537 (N_15537,N_12923,N_13214);
nor U15538 (N_15538,N_12752,N_13923);
nor U15539 (N_15539,N_12206,N_13709);
nor U15540 (N_15540,N_12099,N_13803);
or U15541 (N_15541,N_12572,N_12944);
or U15542 (N_15542,N_12973,N_13793);
or U15543 (N_15543,N_12603,N_12122);
xor U15544 (N_15544,N_12210,N_13986);
xor U15545 (N_15545,N_12189,N_12893);
and U15546 (N_15546,N_12790,N_13485);
or U15547 (N_15547,N_13651,N_13963);
nor U15548 (N_15548,N_13057,N_13083);
nand U15549 (N_15549,N_12209,N_12430);
nand U15550 (N_15550,N_12033,N_13645);
nand U15551 (N_15551,N_12554,N_13030);
or U15552 (N_15552,N_13253,N_12372);
or U15553 (N_15553,N_13367,N_12649);
nor U15554 (N_15554,N_12707,N_12092);
nor U15555 (N_15555,N_13308,N_13271);
nor U15556 (N_15556,N_12103,N_13501);
and U15557 (N_15557,N_13682,N_12723);
nand U15558 (N_15558,N_13061,N_13142);
xnor U15559 (N_15559,N_13065,N_13904);
nand U15560 (N_15560,N_13700,N_12362);
nand U15561 (N_15561,N_13873,N_13792);
nor U15562 (N_15562,N_12260,N_13072);
or U15563 (N_15563,N_13527,N_13407);
xor U15564 (N_15564,N_13938,N_13648);
nand U15565 (N_15565,N_13688,N_12341);
or U15566 (N_15566,N_12553,N_13123);
xor U15567 (N_15567,N_12924,N_13720);
xor U15568 (N_15568,N_12267,N_12498);
or U15569 (N_15569,N_12332,N_13584);
nand U15570 (N_15570,N_13061,N_13156);
xnor U15571 (N_15571,N_12122,N_13415);
nor U15572 (N_15572,N_12309,N_13517);
nand U15573 (N_15573,N_13621,N_12426);
nor U15574 (N_15574,N_12989,N_13866);
and U15575 (N_15575,N_12322,N_12988);
nor U15576 (N_15576,N_13180,N_13352);
xor U15577 (N_15577,N_13620,N_12221);
xor U15578 (N_15578,N_13669,N_12394);
nor U15579 (N_15579,N_13282,N_13131);
xnor U15580 (N_15580,N_12934,N_12692);
or U15581 (N_15581,N_13419,N_12206);
or U15582 (N_15582,N_13824,N_12650);
nor U15583 (N_15583,N_12687,N_13742);
xor U15584 (N_15584,N_13553,N_12546);
nor U15585 (N_15585,N_12764,N_13633);
or U15586 (N_15586,N_12090,N_12232);
nand U15587 (N_15587,N_12134,N_12617);
xor U15588 (N_15588,N_13511,N_12249);
xor U15589 (N_15589,N_13708,N_13675);
nand U15590 (N_15590,N_12409,N_13308);
and U15591 (N_15591,N_13017,N_13403);
nand U15592 (N_15592,N_13817,N_12672);
xor U15593 (N_15593,N_12764,N_12133);
nand U15594 (N_15594,N_12352,N_12122);
nor U15595 (N_15595,N_13544,N_13255);
nand U15596 (N_15596,N_12555,N_12771);
or U15597 (N_15597,N_12362,N_12840);
and U15598 (N_15598,N_13997,N_13085);
or U15599 (N_15599,N_12850,N_12280);
or U15600 (N_15600,N_12962,N_12639);
nand U15601 (N_15601,N_13936,N_13243);
and U15602 (N_15602,N_13836,N_12392);
nand U15603 (N_15603,N_12684,N_12985);
or U15604 (N_15604,N_12114,N_12756);
or U15605 (N_15605,N_12484,N_13780);
nand U15606 (N_15606,N_12431,N_12807);
and U15607 (N_15607,N_13852,N_12875);
nand U15608 (N_15608,N_12712,N_13775);
nand U15609 (N_15609,N_13152,N_13838);
and U15610 (N_15610,N_13112,N_13166);
xor U15611 (N_15611,N_12903,N_12967);
or U15612 (N_15612,N_12280,N_12780);
nand U15613 (N_15613,N_13945,N_12171);
nand U15614 (N_15614,N_13030,N_12481);
or U15615 (N_15615,N_12505,N_12583);
and U15616 (N_15616,N_12494,N_12737);
and U15617 (N_15617,N_13819,N_13521);
or U15618 (N_15618,N_13684,N_13705);
or U15619 (N_15619,N_13050,N_13078);
or U15620 (N_15620,N_12569,N_12387);
nand U15621 (N_15621,N_13012,N_13001);
nor U15622 (N_15622,N_13337,N_13067);
xor U15623 (N_15623,N_12349,N_12318);
nor U15624 (N_15624,N_12742,N_13721);
or U15625 (N_15625,N_12966,N_12607);
and U15626 (N_15626,N_12307,N_12479);
nor U15627 (N_15627,N_13142,N_12586);
nor U15628 (N_15628,N_13260,N_13437);
nor U15629 (N_15629,N_12052,N_12291);
nand U15630 (N_15630,N_12244,N_12824);
nand U15631 (N_15631,N_13828,N_13641);
xor U15632 (N_15632,N_12996,N_13290);
and U15633 (N_15633,N_12941,N_13882);
and U15634 (N_15634,N_12746,N_13879);
xor U15635 (N_15635,N_13091,N_13429);
xnor U15636 (N_15636,N_12913,N_13793);
nor U15637 (N_15637,N_13827,N_12336);
nand U15638 (N_15638,N_13953,N_12524);
xor U15639 (N_15639,N_12329,N_12385);
nand U15640 (N_15640,N_13703,N_13015);
nor U15641 (N_15641,N_13227,N_12653);
nand U15642 (N_15642,N_12100,N_13723);
and U15643 (N_15643,N_12053,N_12378);
xor U15644 (N_15644,N_13584,N_13325);
and U15645 (N_15645,N_13010,N_13240);
or U15646 (N_15646,N_12408,N_12700);
nand U15647 (N_15647,N_13359,N_13315);
nor U15648 (N_15648,N_12865,N_12911);
xor U15649 (N_15649,N_12760,N_12716);
xor U15650 (N_15650,N_13474,N_13974);
nand U15651 (N_15651,N_13811,N_13322);
or U15652 (N_15652,N_12056,N_13340);
and U15653 (N_15653,N_13628,N_13530);
and U15654 (N_15654,N_12519,N_13439);
xor U15655 (N_15655,N_13151,N_12404);
nor U15656 (N_15656,N_13761,N_13691);
xnor U15657 (N_15657,N_13258,N_13828);
nand U15658 (N_15658,N_13179,N_12636);
nand U15659 (N_15659,N_12341,N_13269);
or U15660 (N_15660,N_13936,N_13002);
nor U15661 (N_15661,N_12111,N_13146);
or U15662 (N_15662,N_12570,N_13052);
nand U15663 (N_15663,N_13049,N_12637);
nor U15664 (N_15664,N_12387,N_12605);
nor U15665 (N_15665,N_13714,N_12223);
xnor U15666 (N_15666,N_12714,N_13544);
and U15667 (N_15667,N_12939,N_12409);
and U15668 (N_15668,N_13606,N_12883);
and U15669 (N_15669,N_12828,N_12647);
and U15670 (N_15670,N_13492,N_12673);
and U15671 (N_15671,N_13309,N_12229);
nand U15672 (N_15672,N_12777,N_13335);
nand U15673 (N_15673,N_12394,N_13654);
and U15674 (N_15674,N_13112,N_12000);
and U15675 (N_15675,N_13772,N_12658);
or U15676 (N_15676,N_13650,N_13111);
nor U15677 (N_15677,N_12678,N_12921);
or U15678 (N_15678,N_12970,N_13179);
and U15679 (N_15679,N_12315,N_12276);
and U15680 (N_15680,N_13808,N_13796);
nor U15681 (N_15681,N_12051,N_12041);
nand U15682 (N_15682,N_13182,N_12633);
xor U15683 (N_15683,N_13210,N_12034);
nand U15684 (N_15684,N_12929,N_12946);
xnor U15685 (N_15685,N_12904,N_12296);
xnor U15686 (N_15686,N_12156,N_13180);
nand U15687 (N_15687,N_12113,N_12627);
nand U15688 (N_15688,N_12794,N_13155);
and U15689 (N_15689,N_13001,N_13869);
or U15690 (N_15690,N_12674,N_13138);
nand U15691 (N_15691,N_13655,N_13270);
nand U15692 (N_15692,N_13321,N_13835);
nand U15693 (N_15693,N_13504,N_13042);
and U15694 (N_15694,N_13268,N_13725);
nor U15695 (N_15695,N_12438,N_12365);
nor U15696 (N_15696,N_12128,N_13748);
or U15697 (N_15697,N_13437,N_13225);
or U15698 (N_15698,N_13975,N_13513);
or U15699 (N_15699,N_12032,N_12235);
xnor U15700 (N_15700,N_13368,N_13000);
and U15701 (N_15701,N_12174,N_12785);
nand U15702 (N_15702,N_12858,N_12933);
nand U15703 (N_15703,N_13957,N_13066);
xor U15704 (N_15704,N_12657,N_12404);
nand U15705 (N_15705,N_12072,N_12755);
and U15706 (N_15706,N_13760,N_12124);
nand U15707 (N_15707,N_13281,N_12568);
and U15708 (N_15708,N_13215,N_13050);
xnor U15709 (N_15709,N_12243,N_12721);
xnor U15710 (N_15710,N_12836,N_13709);
and U15711 (N_15711,N_13531,N_13885);
nand U15712 (N_15712,N_13585,N_13288);
or U15713 (N_15713,N_12341,N_13222);
xnor U15714 (N_15714,N_13237,N_12462);
nand U15715 (N_15715,N_13122,N_13118);
nand U15716 (N_15716,N_13561,N_12885);
or U15717 (N_15717,N_13704,N_13409);
and U15718 (N_15718,N_12989,N_12182);
or U15719 (N_15719,N_12406,N_13153);
or U15720 (N_15720,N_12764,N_12183);
nor U15721 (N_15721,N_13041,N_12817);
nor U15722 (N_15722,N_12466,N_13773);
xnor U15723 (N_15723,N_13617,N_12866);
and U15724 (N_15724,N_13003,N_12299);
xor U15725 (N_15725,N_13615,N_13184);
or U15726 (N_15726,N_12052,N_12737);
xor U15727 (N_15727,N_12880,N_12409);
xor U15728 (N_15728,N_13642,N_12732);
nor U15729 (N_15729,N_12808,N_12274);
and U15730 (N_15730,N_12461,N_12797);
nor U15731 (N_15731,N_13067,N_13644);
nand U15732 (N_15732,N_12693,N_12273);
or U15733 (N_15733,N_13989,N_12135);
xnor U15734 (N_15734,N_12197,N_13760);
nand U15735 (N_15735,N_13381,N_13705);
xor U15736 (N_15736,N_13852,N_13701);
and U15737 (N_15737,N_12867,N_12293);
or U15738 (N_15738,N_12053,N_13472);
and U15739 (N_15739,N_13449,N_13074);
nor U15740 (N_15740,N_12508,N_13646);
nor U15741 (N_15741,N_12059,N_13054);
xor U15742 (N_15742,N_13642,N_12778);
nor U15743 (N_15743,N_13377,N_12849);
xor U15744 (N_15744,N_12542,N_12282);
or U15745 (N_15745,N_12013,N_12091);
and U15746 (N_15746,N_12001,N_13169);
xor U15747 (N_15747,N_13077,N_12289);
nor U15748 (N_15748,N_12700,N_12687);
or U15749 (N_15749,N_13492,N_12752);
or U15750 (N_15750,N_12436,N_12049);
nand U15751 (N_15751,N_13227,N_13816);
nor U15752 (N_15752,N_13615,N_13772);
and U15753 (N_15753,N_12505,N_13044);
or U15754 (N_15754,N_13174,N_13675);
xnor U15755 (N_15755,N_12349,N_13872);
or U15756 (N_15756,N_12480,N_12555);
nand U15757 (N_15757,N_12463,N_12423);
xor U15758 (N_15758,N_13523,N_13972);
and U15759 (N_15759,N_13809,N_13385);
or U15760 (N_15760,N_12710,N_13461);
nor U15761 (N_15761,N_13322,N_12834);
or U15762 (N_15762,N_12360,N_12726);
nor U15763 (N_15763,N_12685,N_13238);
nor U15764 (N_15764,N_12621,N_12658);
or U15765 (N_15765,N_12787,N_12972);
xnor U15766 (N_15766,N_13047,N_13373);
nand U15767 (N_15767,N_13325,N_13378);
nor U15768 (N_15768,N_13247,N_13170);
xor U15769 (N_15769,N_13922,N_12315);
xnor U15770 (N_15770,N_13593,N_12825);
nor U15771 (N_15771,N_13173,N_13143);
nor U15772 (N_15772,N_13562,N_12133);
and U15773 (N_15773,N_13810,N_13843);
xnor U15774 (N_15774,N_12384,N_13245);
or U15775 (N_15775,N_12354,N_12391);
nand U15776 (N_15776,N_13794,N_12861);
nand U15777 (N_15777,N_12422,N_13190);
nand U15778 (N_15778,N_13753,N_12717);
nand U15779 (N_15779,N_12893,N_12820);
or U15780 (N_15780,N_12128,N_13762);
nand U15781 (N_15781,N_13638,N_12841);
or U15782 (N_15782,N_13175,N_12208);
xnor U15783 (N_15783,N_12217,N_12025);
or U15784 (N_15784,N_12948,N_12727);
or U15785 (N_15785,N_13027,N_13096);
nand U15786 (N_15786,N_13521,N_12738);
nand U15787 (N_15787,N_12354,N_12614);
nand U15788 (N_15788,N_13712,N_13597);
xor U15789 (N_15789,N_12526,N_12847);
nor U15790 (N_15790,N_13082,N_12370);
xnor U15791 (N_15791,N_12262,N_12589);
and U15792 (N_15792,N_12921,N_12624);
and U15793 (N_15793,N_12053,N_12474);
nor U15794 (N_15794,N_13764,N_13221);
and U15795 (N_15795,N_12569,N_13851);
or U15796 (N_15796,N_13379,N_12495);
xor U15797 (N_15797,N_13640,N_12197);
xor U15798 (N_15798,N_13249,N_13130);
nor U15799 (N_15799,N_13487,N_12035);
nand U15800 (N_15800,N_13038,N_12607);
nand U15801 (N_15801,N_12959,N_12242);
and U15802 (N_15802,N_12407,N_12142);
nand U15803 (N_15803,N_13459,N_13044);
xnor U15804 (N_15804,N_13869,N_13407);
nand U15805 (N_15805,N_12626,N_13919);
xor U15806 (N_15806,N_13856,N_13621);
and U15807 (N_15807,N_12289,N_13137);
and U15808 (N_15808,N_12182,N_13214);
and U15809 (N_15809,N_13799,N_13744);
nand U15810 (N_15810,N_13492,N_12696);
or U15811 (N_15811,N_12907,N_13405);
or U15812 (N_15812,N_12712,N_12578);
or U15813 (N_15813,N_12194,N_12262);
nor U15814 (N_15814,N_13747,N_12388);
nand U15815 (N_15815,N_13736,N_13148);
nor U15816 (N_15816,N_12274,N_12389);
xnor U15817 (N_15817,N_12611,N_12141);
nand U15818 (N_15818,N_12625,N_13082);
nand U15819 (N_15819,N_12139,N_13400);
nand U15820 (N_15820,N_13486,N_12252);
xnor U15821 (N_15821,N_12807,N_13592);
xor U15822 (N_15822,N_12914,N_13705);
nor U15823 (N_15823,N_12089,N_12860);
xnor U15824 (N_15824,N_13686,N_13186);
xor U15825 (N_15825,N_13511,N_12750);
nor U15826 (N_15826,N_13029,N_13619);
xnor U15827 (N_15827,N_12090,N_12697);
and U15828 (N_15828,N_12253,N_13362);
and U15829 (N_15829,N_12440,N_12909);
or U15830 (N_15830,N_13826,N_13770);
and U15831 (N_15831,N_13844,N_12889);
xnor U15832 (N_15832,N_12736,N_12371);
and U15833 (N_15833,N_13739,N_13152);
or U15834 (N_15834,N_12831,N_12445);
nand U15835 (N_15835,N_12032,N_12755);
nor U15836 (N_15836,N_12895,N_13862);
nor U15837 (N_15837,N_12408,N_13216);
or U15838 (N_15838,N_13066,N_12293);
xnor U15839 (N_15839,N_12316,N_13284);
or U15840 (N_15840,N_13731,N_13298);
nor U15841 (N_15841,N_13532,N_13076);
and U15842 (N_15842,N_12570,N_12660);
xnor U15843 (N_15843,N_12470,N_13848);
xor U15844 (N_15844,N_12928,N_13707);
and U15845 (N_15845,N_12871,N_13231);
or U15846 (N_15846,N_13368,N_13169);
nor U15847 (N_15847,N_12452,N_13912);
xnor U15848 (N_15848,N_13384,N_13284);
xnor U15849 (N_15849,N_12280,N_12329);
nand U15850 (N_15850,N_12416,N_12602);
or U15851 (N_15851,N_13996,N_12645);
and U15852 (N_15852,N_12407,N_12208);
nand U15853 (N_15853,N_13042,N_13867);
nand U15854 (N_15854,N_12962,N_12748);
and U15855 (N_15855,N_12201,N_13593);
nand U15856 (N_15856,N_13141,N_13487);
nand U15857 (N_15857,N_13964,N_13622);
xor U15858 (N_15858,N_12656,N_13495);
nor U15859 (N_15859,N_12850,N_12929);
nand U15860 (N_15860,N_12099,N_12708);
and U15861 (N_15861,N_12973,N_13580);
and U15862 (N_15862,N_12766,N_13730);
nand U15863 (N_15863,N_12359,N_12228);
xor U15864 (N_15864,N_13304,N_13438);
and U15865 (N_15865,N_13823,N_12207);
xor U15866 (N_15866,N_13443,N_12112);
or U15867 (N_15867,N_13355,N_12695);
nor U15868 (N_15868,N_12017,N_13758);
nor U15869 (N_15869,N_12066,N_13867);
or U15870 (N_15870,N_12159,N_12453);
nor U15871 (N_15871,N_12414,N_12710);
nor U15872 (N_15872,N_12532,N_12091);
xor U15873 (N_15873,N_12062,N_13856);
or U15874 (N_15874,N_12179,N_13141);
xor U15875 (N_15875,N_13135,N_12756);
xor U15876 (N_15876,N_13446,N_13457);
nor U15877 (N_15877,N_13908,N_12307);
nor U15878 (N_15878,N_12385,N_13799);
nor U15879 (N_15879,N_12874,N_13935);
xor U15880 (N_15880,N_12472,N_12770);
and U15881 (N_15881,N_12662,N_13937);
nor U15882 (N_15882,N_12660,N_13869);
or U15883 (N_15883,N_12184,N_13904);
or U15884 (N_15884,N_12093,N_12484);
nor U15885 (N_15885,N_12619,N_12439);
and U15886 (N_15886,N_13490,N_13492);
nor U15887 (N_15887,N_12672,N_13706);
nand U15888 (N_15888,N_13657,N_12927);
nor U15889 (N_15889,N_13251,N_13215);
nor U15890 (N_15890,N_12948,N_12401);
and U15891 (N_15891,N_13382,N_13825);
nor U15892 (N_15892,N_13831,N_12450);
nand U15893 (N_15893,N_13429,N_13694);
nand U15894 (N_15894,N_12374,N_12908);
or U15895 (N_15895,N_13619,N_12089);
and U15896 (N_15896,N_12293,N_13869);
xor U15897 (N_15897,N_12751,N_13960);
and U15898 (N_15898,N_12849,N_12880);
or U15899 (N_15899,N_12616,N_13580);
xor U15900 (N_15900,N_13986,N_13880);
or U15901 (N_15901,N_13833,N_12087);
and U15902 (N_15902,N_13815,N_13198);
or U15903 (N_15903,N_13618,N_13315);
nand U15904 (N_15904,N_13951,N_12190);
xnor U15905 (N_15905,N_13242,N_13426);
or U15906 (N_15906,N_13729,N_12279);
or U15907 (N_15907,N_12430,N_12850);
xnor U15908 (N_15908,N_13963,N_13924);
xnor U15909 (N_15909,N_12776,N_12905);
nand U15910 (N_15910,N_13452,N_13279);
xor U15911 (N_15911,N_13942,N_13558);
or U15912 (N_15912,N_12620,N_13821);
xnor U15913 (N_15913,N_12294,N_13893);
or U15914 (N_15914,N_12586,N_12474);
nand U15915 (N_15915,N_13555,N_12210);
nand U15916 (N_15916,N_13374,N_13267);
nand U15917 (N_15917,N_13556,N_13127);
and U15918 (N_15918,N_13928,N_13003);
nand U15919 (N_15919,N_12252,N_13348);
xnor U15920 (N_15920,N_12928,N_13148);
and U15921 (N_15921,N_12947,N_13269);
and U15922 (N_15922,N_12331,N_12415);
or U15923 (N_15923,N_12632,N_12659);
or U15924 (N_15924,N_13152,N_13930);
nor U15925 (N_15925,N_13730,N_13934);
or U15926 (N_15926,N_13917,N_13831);
or U15927 (N_15927,N_12210,N_13296);
or U15928 (N_15928,N_12428,N_12202);
nor U15929 (N_15929,N_13494,N_13615);
or U15930 (N_15930,N_13315,N_12865);
nand U15931 (N_15931,N_12480,N_13071);
nor U15932 (N_15932,N_13122,N_12455);
and U15933 (N_15933,N_12033,N_12711);
nor U15934 (N_15934,N_12098,N_13673);
or U15935 (N_15935,N_13437,N_13364);
nand U15936 (N_15936,N_12234,N_12889);
and U15937 (N_15937,N_13095,N_12686);
nand U15938 (N_15938,N_13618,N_13226);
nor U15939 (N_15939,N_13728,N_13248);
nor U15940 (N_15940,N_13437,N_12726);
xnor U15941 (N_15941,N_13082,N_13307);
or U15942 (N_15942,N_12006,N_12627);
nor U15943 (N_15943,N_13200,N_12178);
nor U15944 (N_15944,N_13121,N_13263);
nand U15945 (N_15945,N_12639,N_12008);
xnor U15946 (N_15946,N_13578,N_13334);
or U15947 (N_15947,N_13588,N_13043);
nand U15948 (N_15948,N_13225,N_13891);
nor U15949 (N_15949,N_13893,N_13535);
nand U15950 (N_15950,N_13930,N_12200);
nor U15951 (N_15951,N_13473,N_12060);
nor U15952 (N_15952,N_12007,N_13922);
nand U15953 (N_15953,N_13477,N_13819);
nor U15954 (N_15954,N_12566,N_12408);
xnor U15955 (N_15955,N_13640,N_12615);
nand U15956 (N_15956,N_13511,N_12928);
and U15957 (N_15957,N_12984,N_12084);
and U15958 (N_15958,N_13663,N_13319);
nand U15959 (N_15959,N_12279,N_12730);
xnor U15960 (N_15960,N_13057,N_12248);
xnor U15961 (N_15961,N_12606,N_12841);
xor U15962 (N_15962,N_12860,N_13338);
nor U15963 (N_15963,N_13105,N_13856);
xnor U15964 (N_15964,N_12416,N_12165);
nor U15965 (N_15965,N_12361,N_13841);
nor U15966 (N_15966,N_13054,N_13720);
nor U15967 (N_15967,N_13563,N_12216);
nor U15968 (N_15968,N_12062,N_12587);
xor U15969 (N_15969,N_13750,N_13993);
nor U15970 (N_15970,N_13488,N_13073);
nor U15971 (N_15971,N_12947,N_12097);
nor U15972 (N_15972,N_12759,N_13564);
nor U15973 (N_15973,N_13733,N_12510);
or U15974 (N_15974,N_13532,N_12229);
xnor U15975 (N_15975,N_12915,N_12756);
xor U15976 (N_15976,N_13783,N_12281);
nand U15977 (N_15977,N_13037,N_12826);
nand U15978 (N_15978,N_13720,N_12508);
and U15979 (N_15979,N_13173,N_12460);
nor U15980 (N_15980,N_12109,N_12360);
nor U15981 (N_15981,N_13329,N_12317);
nor U15982 (N_15982,N_12480,N_12551);
or U15983 (N_15983,N_12694,N_13140);
and U15984 (N_15984,N_12522,N_12626);
nor U15985 (N_15985,N_13714,N_13486);
or U15986 (N_15986,N_12629,N_12731);
and U15987 (N_15987,N_13729,N_13724);
nand U15988 (N_15988,N_13444,N_13307);
or U15989 (N_15989,N_12001,N_13911);
xor U15990 (N_15990,N_13831,N_12433);
and U15991 (N_15991,N_13714,N_12870);
and U15992 (N_15992,N_13375,N_13625);
nor U15993 (N_15993,N_13072,N_13342);
xnor U15994 (N_15994,N_13914,N_13171);
nor U15995 (N_15995,N_12340,N_13338);
or U15996 (N_15996,N_12764,N_13908);
nand U15997 (N_15997,N_12249,N_12099);
nor U15998 (N_15998,N_12118,N_13437);
nand U15999 (N_15999,N_13103,N_12328);
nand U16000 (N_16000,N_15929,N_14310);
nand U16001 (N_16001,N_15652,N_15090);
and U16002 (N_16002,N_14886,N_14269);
and U16003 (N_16003,N_14607,N_15196);
xor U16004 (N_16004,N_14194,N_15354);
or U16005 (N_16005,N_15857,N_15717);
nand U16006 (N_16006,N_15100,N_14105);
xor U16007 (N_16007,N_15879,N_15595);
nand U16008 (N_16008,N_15638,N_15553);
nand U16009 (N_16009,N_15157,N_15637);
xnor U16010 (N_16010,N_14390,N_15561);
or U16011 (N_16011,N_15451,N_14075);
xor U16012 (N_16012,N_14327,N_15645);
nand U16013 (N_16013,N_14610,N_14147);
nor U16014 (N_16014,N_14500,N_15710);
nand U16015 (N_16015,N_15082,N_15377);
or U16016 (N_16016,N_14080,N_14704);
xnor U16017 (N_16017,N_15886,N_14170);
and U16018 (N_16018,N_15881,N_14553);
and U16019 (N_16019,N_14861,N_15084);
or U16020 (N_16020,N_14707,N_14256);
xnor U16021 (N_16021,N_14863,N_15726);
nor U16022 (N_16022,N_15935,N_15365);
nand U16023 (N_16023,N_15471,N_15011);
or U16024 (N_16024,N_14044,N_15620);
nor U16025 (N_16025,N_15441,N_15701);
or U16026 (N_16026,N_14841,N_14539);
and U16027 (N_16027,N_15756,N_14814);
or U16028 (N_16028,N_14839,N_14909);
nor U16029 (N_16029,N_14868,N_14017);
or U16030 (N_16030,N_14238,N_15842);
or U16031 (N_16031,N_15721,N_15640);
nand U16032 (N_16032,N_15831,N_14339);
nor U16033 (N_16033,N_14775,N_15765);
xnor U16034 (N_16034,N_14733,N_14838);
or U16035 (N_16035,N_15642,N_15329);
xnor U16036 (N_16036,N_14217,N_15577);
or U16037 (N_16037,N_15811,N_14006);
xor U16038 (N_16038,N_15630,N_14290);
nand U16039 (N_16039,N_14005,N_15657);
and U16040 (N_16040,N_15078,N_14699);
nand U16041 (N_16041,N_14320,N_15407);
and U16042 (N_16042,N_14904,N_15653);
nor U16043 (N_16043,N_14350,N_14959);
nor U16044 (N_16044,N_14621,N_14282);
and U16045 (N_16045,N_15161,N_15439);
or U16046 (N_16046,N_15192,N_14656);
nand U16047 (N_16047,N_15963,N_14203);
or U16048 (N_16048,N_14905,N_14422);
xnor U16049 (N_16049,N_14537,N_15564);
or U16050 (N_16050,N_14362,N_14204);
and U16051 (N_16051,N_14735,N_14094);
nand U16052 (N_16052,N_14358,N_14802);
nor U16053 (N_16053,N_14039,N_15506);
and U16054 (N_16054,N_15367,N_14109);
xor U16055 (N_16055,N_14564,N_15509);
and U16056 (N_16056,N_15076,N_14205);
or U16057 (N_16057,N_14074,N_15818);
or U16058 (N_16058,N_14948,N_15228);
nand U16059 (N_16059,N_14193,N_14288);
nand U16060 (N_16060,N_15650,N_14262);
or U16061 (N_16061,N_15624,N_14215);
or U16062 (N_16062,N_15415,N_14368);
nor U16063 (N_16063,N_14963,N_15074);
nor U16064 (N_16064,N_14450,N_14121);
nand U16065 (N_16065,N_14561,N_14908);
or U16066 (N_16066,N_15708,N_14465);
and U16067 (N_16067,N_14071,N_14442);
or U16068 (N_16068,N_15408,N_14030);
or U16069 (N_16069,N_14991,N_15562);
nand U16070 (N_16070,N_14898,N_14662);
and U16071 (N_16071,N_15641,N_15602);
nand U16072 (N_16072,N_14603,N_14344);
and U16073 (N_16073,N_14062,N_14411);
nor U16074 (N_16074,N_14661,N_14003);
and U16075 (N_16075,N_14558,N_15116);
or U16076 (N_16076,N_15080,N_14095);
or U16077 (N_16077,N_15573,N_14859);
nor U16078 (N_16078,N_15865,N_14509);
nand U16079 (N_16079,N_15212,N_14754);
xnor U16080 (N_16080,N_15413,N_14867);
and U16081 (N_16081,N_14323,N_14515);
nor U16082 (N_16082,N_14976,N_14043);
nand U16083 (N_16083,N_15837,N_14059);
nor U16084 (N_16084,N_14178,N_15675);
nand U16085 (N_16085,N_14294,N_15584);
xnor U16086 (N_16086,N_15284,N_15846);
xor U16087 (N_16087,N_15106,N_14984);
or U16088 (N_16088,N_14319,N_15986);
nor U16089 (N_16089,N_14950,N_15512);
or U16090 (N_16090,N_15085,N_14123);
and U16091 (N_16091,N_15753,N_14326);
nor U16092 (N_16092,N_14053,N_14389);
or U16093 (N_16093,N_15751,N_14789);
nand U16094 (N_16094,N_15282,N_14804);
nor U16095 (N_16095,N_15055,N_14126);
xnor U16096 (N_16096,N_15111,N_14514);
xor U16097 (N_16097,N_14918,N_14490);
xor U16098 (N_16098,N_15098,N_15950);
or U16099 (N_16099,N_15558,N_15022);
nand U16100 (N_16100,N_14703,N_15387);
nor U16101 (N_16101,N_15006,N_14932);
nand U16102 (N_16102,N_14201,N_14835);
xnor U16103 (N_16103,N_14190,N_14945);
nor U16104 (N_16104,N_15582,N_15121);
xnor U16105 (N_16105,N_15045,N_14919);
nor U16106 (N_16106,N_14493,N_14988);
nor U16107 (N_16107,N_15031,N_15548);
nor U16108 (N_16108,N_14025,N_15610);
and U16109 (N_16109,N_14400,N_14040);
and U16110 (N_16110,N_14793,N_15406);
nor U16111 (N_16111,N_15166,N_15515);
xor U16112 (N_16112,N_15936,N_15679);
nor U16113 (N_16113,N_14641,N_15016);
and U16114 (N_16114,N_14158,N_14923);
nor U16115 (N_16115,N_15146,N_14710);
and U16116 (N_16116,N_15958,N_15040);
xor U16117 (N_16117,N_14504,N_14535);
or U16118 (N_16118,N_14482,N_14391);
xor U16119 (N_16119,N_15030,N_14419);
and U16120 (N_16120,N_14765,N_14278);
or U16121 (N_16121,N_14873,N_15421);
or U16122 (N_16122,N_15829,N_15547);
nand U16123 (N_16123,N_15903,N_15976);
nand U16124 (N_16124,N_14027,N_14745);
and U16125 (N_16125,N_15418,N_15800);
nand U16126 (N_16126,N_14018,N_14554);
and U16127 (N_16127,N_14732,N_14881);
and U16128 (N_16128,N_14267,N_14674);
nand U16129 (N_16129,N_15430,N_15005);
nor U16130 (N_16130,N_15783,N_15681);
nand U16131 (N_16131,N_14488,N_15945);
nand U16132 (N_16132,N_14675,N_15609);
nor U16133 (N_16133,N_15817,N_15165);
nor U16134 (N_16134,N_14229,N_15479);
xor U16135 (N_16135,N_15394,N_15779);
xnor U16136 (N_16136,N_15919,N_14336);
xnor U16137 (N_16137,N_14851,N_14370);
nand U16138 (N_16138,N_15646,N_15442);
nand U16139 (N_16139,N_15019,N_14525);
nor U16140 (N_16140,N_14041,N_14879);
nor U16141 (N_16141,N_14542,N_14133);
xor U16142 (N_16142,N_14616,N_15426);
nand U16143 (N_16143,N_14101,N_15771);
nor U16144 (N_16144,N_14737,N_15793);
and U16145 (N_16145,N_14401,N_14944);
nor U16146 (N_16146,N_14461,N_15521);
xnor U16147 (N_16147,N_14404,N_14246);
nand U16148 (N_16148,N_15156,N_15494);
xor U16149 (N_16149,N_14545,N_14716);
xor U16150 (N_16150,N_15921,N_14129);
or U16151 (N_16151,N_15676,N_15073);
and U16152 (N_16152,N_15974,N_15768);
or U16153 (N_16153,N_14372,N_14993);
and U16154 (N_16154,N_14629,N_15239);
xor U16155 (N_16155,N_14253,N_14533);
or U16156 (N_16156,N_15890,N_14806);
nand U16157 (N_16157,N_15238,N_15036);
and U16158 (N_16158,N_14314,N_15887);
xor U16159 (N_16159,N_14852,N_14785);
xor U16160 (N_16160,N_15320,N_15697);
nor U16161 (N_16161,N_14854,N_14882);
nand U16162 (N_16162,N_15330,N_15613);
or U16163 (N_16163,N_14477,N_14046);
and U16164 (N_16164,N_14956,N_15896);
or U16165 (N_16165,N_15917,N_14531);
nor U16166 (N_16166,N_14184,N_15245);
nor U16167 (N_16167,N_14305,N_14518);
and U16168 (N_16168,N_15568,N_15816);
or U16169 (N_16169,N_15601,N_15296);
nor U16170 (N_16170,N_14657,N_14495);
or U16171 (N_16171,N_15002,N_14055);
or U16172 (N_16172,N_15205,N_15062);
xor U16173 (N_16173,N_15826,N_14567);
nand U16174 (N_16174,N_15252,N_15782);
xnor U16175 (N_16175,N_14388,N_15464);
xor U16176 (N_16176,N_15511,N_15948);
or U16177 (N_16177,N_14432,N_15338);
and U16178 (N_16178,N_14066,N_14242);
xnor U16179 (N_16179,N_15105,N_15133);
and U16180 (N_16180,N_15627,N_14408);
nand U16181 (N_16181,N_14077,N_14611);
nand U16182 (N_16182,N_15142,N_15434);
xnor U16183 (N_16183,N_14165,N_15749);
nand U16184 (N_16184,N_15889,N_14632);
or U16185 (N_16185,N_14056,N_14568);
xor U16186 (N_16186,N_14740,N_14763);
nor U16187 (N_16187,N_15026,N_14148);
or U16188 (N_16188,N_15249,N_14683);
nor U16189 (N_16189,N_15836,N_15323);
nor U16190 (N_16190,N_15486,N_14520);
and U16191 (N_16191,N_15674,N_14110);
nor U16192 (N_16192,N_14702,N_14787);
or U16193 (N_16193,N_14125,N_15206);
nor U16194 (N_16194,N_15195,N_14605);
or U16195 (N_16195,N_14715,N_15064);
nor U16196 (N_16196,N_14840,N_15762);
xnor U16197 (N_16197,N_15004,N_14858);
and U16198 (N_16198,N_15550,N_14717);
or U16199 (N_16199,N_14576,N_15979);
nor U16200 (N_16200,N_15712,N_14188);
xor U16201 (N_16201,N_14255,N_14916);
nand U16202 (N_16202,N_15563,N_14414);
and U16203 (N_16203,N_14550,N_15096);
nor U16204 (N_16204,N_15199,N_15844);
nor U16205 (N_16205,N_15507,N_15869);
or U16206 (N_16206,N_14690,N_14070);
xnor U16207 (N_16207,N_14397,N_14503);
and U16208 (N_16208,N_14471,N_14777);
xnor U16209 (N_16209,N_15028,N_15220);
xor U16210 (N_16210,N_15764,N_14354);
or U16211 (N_16211,N_14087,N_14770);
and U16212 (N_16212,N_15566,N_15218);
nor U16213 (N_16213,N_15739,N_14272);
or U16214 (N_16214,N_15221,N_15549);
nand U16215 (N_16215,N_15557,N_15314);
nor U16216 (N_16216,N_15207,N_15589);
xnor U16217 (N_16217,N_15757,N_15923);
or U16218 (N_16218,N_15361,N_14325);
nor U16219 (N_16219,N_14136,N_14824);
nor U16220 (N_16220,N_14163,N_14214);
xor U16221 (N_16221,N_15885,N_14334);
nand U16222 (N_16222,N_15301,N_15944);
xnor U16223 (N_16223,N_15417,N_15713);
or U16224 (N_16224,N_15532,N_15385);
and U16225 (N_16225,N_15001,N_15801);
or U16226 (N_16226,N_14175,N_14132);
nand U16227 (N_16227,N_15286,N_15079);
nand U16228 (N_16228,N_15457,N_14197);
nor U16229 (N_16229,N_15216,N_15305);
nor U16230 (N_16230,N_14228,N_15876);
nor U16231 (N_16231,N_14399,N_14659);
nor U16232 (N_16232,N_14687,N_15194);
or U16233 (N_16233,N_15290,N_15786);
nor U16234 (N_16234,N_15174,N_15344);
nor U16235 (N_16235,N_14751,N_15389);
or U16236 (N_16236,N_14731,N_15469);
nand U16237 (N_16237,N_14052,N_15898);
and U16238 (N_16238,N_15141,N_15503);
nand U16239 (N_16239,N_14009,N_14106);
and U16240 (N_16240,N_15346,N_14577);
and U16241 (N_16241,N_15812,N_14357);
xor U16242 (N_16242,N_14393,N_15672);
or U16243 (N_16243,N_15924,N_14973);
xnor U16244 (N_16244,N_15233,N_14206);
xnor U16245 (N_16245,N_15694,N_15705);
xnor U16246 (N_16246,N_15902,N_14845);
and U16247 (N_16247,N_14625,N_14251);
xor U16248 (N_16248,N_15119,N_14795);
nor U16249 (N_16249,N_14124,N_15139);
and U16250 (N_16250,N_14816,N_14938);
and U16251 (N_16251,N_15127,N_15404);
or U16252 (N_16252,N_14478,N_15353);
nor U16253 (N_16253,N_15787,N_14930);
nor U16254 (N_16254,N_14402,N_14591);
nor U16255 (N_16255,N_14713,N_15696);
nor U16256 (N_16256,N_15908,N_15840);
and U16257 (N_16257,N_15470,N_15242);
and U16258 (N_16258,N_15414,N_14324);
nand U16259 (N_16259,N_15411,N_14889);
xor U16260 (N_16260,N_15488,N_15773);
and U16261 (N_16261,N_15667,N_15796);
nand U16262 (N_16262,N_14613,N_15853);
nand U16263 (N_16263,N_14036,N_14068);
and U16264 (N_16264,N_15163,N_15134);
or U16265 (N_16265,N_14250,N_15372);
nand U16266 (N_16266,N_14646,N_14031);
and U16267 (N_16267,N_15049,N_15689);
or U16268 (N_16268,N_15256,N_14364);
or U16269 (N_16269,N_14494,N_15302);
nor U16270 (N_16270,N_14534,N_14021);
and U16271 (N_16271,N_14318,N_15032);
and U16272 (N_16272,N_14363,N_15682);
and U16273 (N_16273,N_14423,N_15677);
nor U16274 (N_16274,N_15476,N_14647);
nand U16275 (N_16275,N_15491,N_14437);
nand U16276 (N_16276,N_15784,N_14002);
nand U16277 (N_16277,N_14417,N_14977);
xnor U16278 (N_16278,N_14834,N_15000);
nand U16279 (N_16279,N_15743,N_15477);
nor U16280 (N_16280,N_15215,N_15043);
nand U16281 (N_16281,N_14634,N_15120);
nor U16282 (N_16282,N_14596,N_14640);
nand U16283 (N_16283,N_14670,N_15519);
and U16284 (N_16284,N_15160,N_14492);
or U16285 (N_16285,N_15147,N_14086);
and U16286 (N_16286,N_14752,N_14821);
or U16287 (N_16287,N_14586,N_14013);
nor U16288 (N_16288,N_15190,N_15525);
xor U16289 (N_16289,N_14639,N_14883);
xnor U16290 (N_16290,N_15292,N_15093);
nor U16291 (N_16291,N_14521,N_15536);
xor U16292 (N_16292,N_14971,N_14454);
xor U16293 (N_16293,N_14407,N_15861);
nand U16294 (N_16294,N_15883,N_14676);
or U16295 (N_16295,N_14928,N_15877);
nor U16296 (N_16296,N_15744,N_15483);
and U16297 (N_16297,N_15187,N_14612);
or U16298 (N_16298,N_14578,N_14947);
nor U16299 (N_16299,N_14297,N_15395);
and U16300 (N_16300,N_15775,N_15524);
nand U16301 (N_16301,N_15961,N_14580);
nand U16302 (N_16302,N_15665,N_15799);
nor U16303 (N_16303,N_15048,N_15734);
nor U16304 (N_16304,N_14857,N_14375);
and U16305 (N_16305,N_15268,N_15149);
and U16306 (N_16306,N_14642,N_14679);
nand U16307 (N_16307,N_15342,N_15695);
and U16308 (N_16308,N_14736,N_15820);
and U16309 (N_16309,N_14760,N_15226);
xnor U16310 (N_16310,N_15311,N_15358);
nand U16311 (N_16311,N_14549,N_14037);
or U16312 (N_16312,N_14058,N_15356);
nand U16313 (N_16313,N_15605,N_15254);
nand U16314 (N_16314,N_15189,N_14896);
nand U16315 (N_16315,N_14146,N_15067);
and U16316 (N_16316,N_15746,N_15438);
nor U16317 (N_16317,N_14540,N_15656);
nand U16318 (N_16318,N_15918,N_14665);
nand U16319 (N_16319,N_14669,N_15214);
or U16320 (N_16320,N_14694,N_15213);
or U16321 (N_16321,N_14221,N_15151);
nor U16322 (N_16322,N_14466,N_14063);
xnor U16323 (N_16323,N_15447,N_14933);
xnor U16324 (N_16324,N_14078,N_14870);
xor U16325 (N_16325,N_15153,N_15433);
nand U16326 (N_16326,N_14556,N_15843);
and U16327 (N_16327,N_15900,N_14748);
nor U16328 (N_16328,N_15537,N_14292);
or U16329 (N_16329,N_15044,N_15496);
and U16330 (N_16330,N_15845,N_15091);
or U16331 (N_16331,N_15643,N_14219);
and U16332 (N_16332,N_14594,N_15684);
nor U16333 (N_16333,N_14572,N_15991);
nor U16334 (N_16334,N_14952,N_14380);
or U16335 (N_16335,N_14780,N_15170);
or U16336 (N_16336,N_15698,N_14968);
nor U16337 (N_16337,N_14377,N_15838);
xnor U16338 (N_16338,N_15915,N_15018);
nor U16339 (N_16339,N_15378,N_15864);
xnor U16340 (N_16340,N_14579,N_15403);
nand U16341 (N_16341,N_14428,N_15209);
xnor U16342 (N_16342,N_15299,N_14379);
and U16343 (N_16343,N_15020,N_15419);
nand U16344 (N_16344,N_14090,N_15485);
or U16345 (N_16345,N_15273,N_14457);
nand U16346 (N_16346,N_14869,N_15224);
xor U16347 (N_16347,N_14277,N_15014);
or U16348 (N_16348,N_15530,N_14626);
xnor U16349 (N_16349,N_15130,N_15914);
nor U16350 (N_16350,N_15115,N_15244);
or U16351 (N_16351,N_14864,N_15352);
nand U16352 (N_16352,N_15009,N_14911);
and U16353 (N_16353,N_14664,N_15939);
nand U16354 (N_16354,N_15114,N_15453);
or U16355 (N_16355,N_14098,N_15855);
nand U16356 (N_16356,N_14452,N_15964);
or U16357 (N_16357,N_14783,N_14724);
nand U16358 (N_16358,N_15308,N_14330);
xor U16359 (N_16359,N_14501,N_14987);
and U16360 (N_16360,N_15970,N_15790);
or U16361 (N_16361,N_15599,N_15087);
or U16362 (N_16362,N_14912,N_14943);
or U16363 (N_16363,N_15535,N_14487);
nand U16364 (N_16364,N_14706,N_15989);
nand U16365 (N_16365,N_15882,N_14774);
nor U16366 (N_16366,N_15380,N_14744);
and U16367 (N_16367,N_15980,N_15270);
nor U16368 (N_16368,N_15628,N_14532);
xor U16369 (N_16369,N_15456,N_15359);
and U16370 (N_16370,N_15440,N_14143);
nor U16371 (N_16371,N_14469,N_15412);
xnor U16372 (N_16372,N_15303,N_15973);
and U16373 (N_16373,N_15673,N_15825);
and U16374 (N_16374,N_15992,N_14722);
nor U16375 (N_16375,N_14949,N_15998);
nand U16376 (N_16376,N_14569,N_15813);
nor U16377 (N_16377,N_15789,N_14620);
or U16378 (N_16378,N_15962,N_15193);
and U16379 (N_16379,N_14920,N_15219);
nor U16380 (N_16380,N_15899,N_14114);
xnor U16381 (N_16381,N_14903,N_15081);
and U16382 (N_16382,N_15051,N_14892);
and U16383 (N_16383,N_14196,N_14524);
nand U16384 (N_16384,N_14243,N_15475);
or U16385 (N_16385,N_15386,N_15135);
nor U16386 (N_16386,N_15092,N_15155);
nor U16387 (N_16387,N_15545,N_15904);
nor U16388 (N_16388,N_14047,N_15579);
and U16389 (N_16389,N_14874,N_15452);
nand U16390 (N_16390,N_14983,N_14711);
xor U16391 (N_16391,N_14805,N_14853);
and U16392 (N_16392,N_15671,N_14479);
nand U16393 (N_16393,N_15835,N_14972);
nor U16394 (N_16394,N_15017,N_14798);
nor U16395 (N_16395,N_15603,N_14624);
or U16396 (N_16396,N_15655,N_15508);
or U16397 (N_16397,N_15586,N_15232);
or U16398 (N_16398,N_15607,N_15815);
nand U16399 (N_16399,N_15578,N_15592);
nor U16400 (N_16400,N_15052,N_14028);
nand U16401 (N_16401,N_14181,N_15481);
and U16402 (N_16402,N_14833,N_15490);
nand U16403 (N_16403,N_14637,N_14343);
xor U16404 (N_16404,N_14067,N_14446);
nor U16405 (N_16405,N_14060,N_14307);
nand U16406 (N_16406,N_14672,N_15666);
or U16407 (N_16407,N_14876,N_14742);
and U16408 (N_16408,N_15928,N_15913);
xnor U16409 (N_16409,N_15388,N_14684);
xnor U16410 (N_16410,N_14225,N_15828);
or U16411 (N_16411,N_15247,N_14489);
nand U16412 (N_16412,N_15740,N_15446);
xnor U16413 (N_16413,N_15333,N_15288);
xnor U16414 (N_16414,N_15791,N_15747);
xor U16415 (N_16415,N_14803,N_15693);
xor U16416 (N_16416,N_15391,N_15347);
and U16417 (N_16417,N_14321,N_14222);
and U16418 (N_16418,N_14440,N_14979);
nor U16419 (N_16419,N_15878,N_15651);
xnor U16420 (N_16420,N_15331,N_15162);
or U16421 (N_16421,N_14131,N_14570);
or U16422 (N_16422,N_14552,N_15229);
and U16423 (N_16423,N_14555,N_15294);
nand U16424 (N_16424,N_15594,N_14384);
nand U16425 (N_16425,N_14207,N_14937);
nand U16426 (N_16426,N_14599,N_15523);
nor U16427 (N_16427,N_14154,N_15042);
or U16428 (N_16428,N_14517,N_15183);
or U16429 (N_16429,N_14788,N_14510);
and U16430 (N_16430,N_14915,N_14273);
and U16431 (N_16431,N_14316,N_15738);
xnor U16432 (N_16432,N_15178,N_15619);
nand U16433 (N_16433,N_15350,N_14476);
nand U16434 (N_16434,N_15383,N_14913);
or U16435 (N_16435,N_14796,N_15806);
nand U16436 (N_16436,N_15851,N_14198);
nand U16437 (N_16437,N_15266,N_15501);
nand U16438 (N_16438,N_15546,N_15179);
and U16439 (N_16439,N_15704,N_15678);
or U16440 (N_16440,N_14790,N_14387);
nand U16441 (N_16441,N_15988,N_14054);
and U16442 (N_16442,N_14447,N_14000);
xnor U16443 (N_16443,N_14152,N_15720);
or U16444 (N_16444,N_15943,N_14072);
or U16445 (N_16445,N_14420,N_14781);
and U16446 (N_16446,N_14223,N_14140);
xnor U16447 (N_16447,N_14906,N_15137);
or U16448 (N_16448,N_15176,N_15200);
nand U16449 (N_16449,N_14275,N_14692);
nor U16450 (N_16450,N_14990,N_15122);
nor U16451 (N_16451,N_14429,N_15322);
nand U16452 (N_16452,N_15171,N_15083);
xor U16453 (N_16453,N_14921,N_15763);
nand U16454 (N_16454,N_15542,N_15965);
xnor U16455 (N_16455,N_14563,N_15072);
or U16456 (N_16456,N_15466,N_15099);
nand U16457 (N_16457,N_14069,N_15262);
nand U16458 (N_16458,N_14871,N_15321);
xor U16459 (N_16459,N_15054,N_14015);
nor U16460 (N_16460,N_15136,N_15208);
xnor U16461 (N_16461,N_14264,N_14955);
nand U16462 (N_16462,N_15066,N_14523);
and U16463 (N_16463,N_14232,N_15222);
xnor U16464 (N_16464,N_14268,N_15852);
nor U16465 (N_16465,N_14485,N_14019);
nand U16466 (N_16466,N_14584,N_15117);
nand U16467 (N_16467,N_14022,N_14199);
or U16468 (N_16468,N_15324,N_14828);
and U16469 (N_16469,N_14931,N_14210);
and U16470 (N_16470,N_14274,N_14271);
xor U16471 (N_16471,N_14011,N_15326);
and U16472 (N_16472,N_15699,N_14213);
or U16473 (N_16473,N_15692,N_14239);
nand U16474 (N_16474,N_14666,N_14942);
nand U16475 (N_16475,N_15856,N_14872);
and U16476 (N_16476,N_15996,N_15364);
and U16477 (N_16477,N_15809,N_14827);
and U16478 (N_16478,N_15180,N_15658);
or U16479 (N_16479,N_14439,N_15425);
and U16480 (N_16480,N_14499,N_14741);
xnor U16481 (N_16481,N_14813,N_15248);
nand U16482 (N_16482,N_15410,N_15849);
xnor U16483 (N_16483,N_15969,N_14285);
nand U16484 (N_16484,N_15925,N_15567);
or U16485 (N_16485,N_14922,N_15381);
or U16486 (N_16486,N_15150,N_15947);
nand U16487 (N_16487,N_15258,N_15770);
or U16488 (N_16488,N_14888,N_14761);
xnor U16489 (N_16489,N_15010,N_14311);
nand U16490 (N_16490,N_14496,N_14801);
or U16491 (N_16491,N_14712,N_14866);
xor U16492 (N_16492,N_14506,N_14951);
or U16493 (N_16493,N_15858,N_14162);
and U16494 (N_16494,N_15423,N_15422);
and U16495 (N_16495,N_14601,N_14786);
or U16496 (N_16496,N_15934,N_15777);
nor U16497 (N_16497,N_14257,N_14463);
xnor U16498 (N_16498,N_15158,N_14455);
and U16499 (N_16499,N_15369,N_15987);
or U16500 (N_16500,N_15772,N_15873);
nor U16501 (N_16501,N_14527,N_15057);
or U16502 (N_16502,N_15716,N_14519);
and U16503 (N_16503,N_14161,N_15867);
and U16504 (N_16504,N_14574,N_14901);
nand U16505 (N_16505,N_15482,N_15614);
or U16506 (N_16506,N_15866,N_14116);
and U16507 (N_16507,N_15736,N_14588);
and U16508 (N_16508,N_14636,N_15396);
and U16509 (N_16509,N_14598,N_15709);
nand U16510 (N_16510,N_14346,N_14186);
or U16511 (N_16511,N_15502,N_14831);
nand U16512 (N_16512,N_14341,N_15400);
or U16513 (N_16513,N_14293,N_15175);
and U16514 (N_16514,N_15527,N_15937);
or U16515 (N_16515,N_14929,N_14260);
xor U16516 (N_16516,N_15754,N_14811);
nor U16517 (N_16517,N_15071,N_14144);
or U16518 (N_16518,N_14122,N_15468);
and U16519 (N_16519,N_15590,N_15204);
xor U16520 (N_16520,N_15217,N_15495);
nand U16521 (N_16521,N_14491,N_15382);
nand U16522 (N_16522,N_15907,N_15824);
and U16523 (N_16523,N_15718,N_14966);
xnor U16524 (N_16524,N_14317,N_15926);
and U16525 (N_16525,N_15587,N_15304);
xnor U16526 (N_16526,N_14927,N_14700);
or U16527 (N_16527,N_14638,N_14048);
or U16528 (N_16528,N_14978,N_14042);
or U16529 (N_16529,N_15008,N_14696);
and U16530 (N_16530,N_15341,N_15465);
nor U16531 (N_16531,N_14369,N_14528);
nand U16532 (N_16532,N_14571,N_14753);
nand U16533 (N_16533,N_14529,N_15235);
nor U16534 (N_16534,N_14050,N_15443);
and U16535 (N_16535,N_15448,N_14686);
nand U16536 (N_16536,N_14436,N_15870);
and U16537 (N_16537,N_14459,N_15240);
xor U16538 (N_16538,N_15690,N_14899);
xor U16539 (N_16539,N_15253,N_15059);
xor U16540 (N_16540,N_14998,N_14355);
nor U16541 (N_16541,N_14082,N_14604);
nand U16542 (N_16542,N_14815,N_15894);
xor U16543 (N_16543,N_14836,N_15225);
xnor U16544 (N_16544,N_14356,N_15688);
nor U16545 (N_16545,N_15376,N_14231);
nor U16546 (N_16546,N_15184,N_14995);
xnor U16547 (N_16547,N_15621,N_14103);
and U16548 (N_16548,N_14832,N_15529);
or U16549 (N_16549,N_15803,N_14128);
nor U16550 (N_16550,N_15618,N_14791);
xnor U16551 (N_16551,N_14980,N_15280);
and U16552 (N_16552,N_15363,N_15999);
nand U16553 (N_16553,N_15393,N_15794);
nor U16554 (N_16554,N_15168,N_15355);
or U16555 (N_16555,N_14079,N_15776);
nand U16556 (N_16556,N_15390,N_15922);
nor U16557 (N_16557,N_15629,N_14374);
and U16558 (N_16558,N_14254,N_14960);
nand U16559 (N_16559,N_14734,N_15289);
and U16560 (N_16560,N_14538,N_14141);
or U16561 (N_16561,N_15260,N_14089);
nand U16562 (N_16562,N_15325,N_15862);
nor U16563 (N_16563,N_15373,N_15340);
xor U16564 (N_16564,N_15104,N_14409);
or U16565 (N_16565,N_15683,N_14284);
nor U16566 (N_16566,N_14530,N_15345);
nor U16567 (N_16567,N_14200,N_14032);
nor U16568 (N_16568,N_15731,N_15140);
or U16569 (N_16569,N_14023,N_15328);
and U16570 (N_16570,N_15649,N_14654);
or U16571 (N_16571,N_14299,N_15234);
nand U16572 (N_16572,N_14997,N_15360);
nand U16573 (N_16573,N_14812,N_15102);
and U16574 (N_16574,N_15409,N_14925);
nand U16575 (N_16575,N_14029,N_15435);
xnor U16576 (N_16576,N_14313,N_15474);
or U16577 (N_16577,N_14348,N_14727);
and U16578 (N_16578,N_14381,N_14279);
nor U16579 (N_16579,N_14671,N_15060);
and U16580 (N_16580,N_14166,N_14398);
xnor U16581 (N_16581,N_14695,N_14349);
nand U16582 (N_16582,N_14230,N_15792);
xnor U16583 (N_16583,N_14758,N_14227);
and U16584 (N_16584,N_14064,N_15251);
or U16585 (N_16585,N_14189,N_14705);
or U16586 (N_16586,N_15250,N_14291);
or U16587 (N_16587,N_15297,N_14547);
nand U16588 (N_16588,N_14191,N_15644);
and U16589 (N_16589,N_15990,N_15203);
or U16590 (N_16590,N_15428,N_14894);
nand U16591 (N_16591,N_14513,N_14467);
xnor U16592 (N_16592,N_14914,N_15972);
or U16593 (N_16593,N_15668,N_14771);
or U16594 (N_16594,N_14195,N_15905);
nand U16595 (N_16595,N_14982,N_15893);
nand U16596 (N_16596,N_15349,N_15131);
nor U16597 (N_16597,N_15901,N_15795);
nand U16598 (N_16598,N_14137,N_14335);
nand U16599 (N_16599,N_15752,N_15035);
or U16600 (N_16600,N_14309,N_15778);
xor U16601 (N_16601,N_14680,N_14038);
nand U16602 (N_16602,N_14443,N_14810);
nor U16603 (N_16603,N_15198,N_15021);
or U16604 (N_16604,N_15571,N_14958);
xor U16605 (N_16605,N_15231,N_15730);
or U16606 (N_16606,N_15110,N_15368);
and U16607 (N_16607,N_14885,N_14139);
nand U16608 (N_16608,N_15516,N_15255);
and U16609 (N_16609,N_15037,N_14653);
or U16610 (N_16610,N_14507,N_14051);
or U16611 (N_16611,N_15337,N_15334);
xor U16612 (N_16612,N_14807,N_14648);
or U16613 (N_16613,N_14725,N_14460);
xor U16614 (N_16614,N_15863,N_15808);
nor U16615 (N_16615,N_14677,N_14091);
nand U16616 (N_16616,N_15277,N_14371);
nor U16617 (N_16617,N_14630,N_14746);
or U16618 (N_16618,N_15500,N_15371);
nand U16619 (N_16619,N_15246,N_15598);
xnor U16620 (N_16620,N_15920,N_15202);
or U16621 (N_16621,N_15554,N_15633);
nor U16622 (N_16622,N_14663,N_14847);
or U16623 (N_16623,N_14365,N_15729);
or U16624 (N_16624,N_14138,N_15761);
xor U16625 (N_16625,N_15534,N_14340);
or U16626 (N_16626,N_15741,N_15661);
nand U16627 (N_16627,N_15462,N_14176);
or U16628 (N_16628,N_14111,N_14145);
xnor U16629 (N_16629,N_15538,N_14403);
nor U16630 (N_16630,N_14855,N_15544);
nor U16631 (N_16631,N_14218,N_14286);
xor U16632 (N_16632,N_15402,N_14652);
nor U16633 (N_16633,N_15181,N_15436);
xnor U16634 (N_16634,N_14415,N_15197);
and U16635 (N_16635,N_14595,N_15480);
nor U16636 (N_16636,N_14104,N_15201);
nor U16637 (N_16637,N_15703,N_14164);
and U16638 (N_16638,N_14606,N_15445);
xor U16639 (N_16639,N_14012,N_15617);
xor U16640 (N_16640,N_15143,N_14234);
nor U16641 (N_16641,N_14249,N_14470);
or U16642 (N_16642,N_14302,N_15985);
nand U16643 (N_16643,N_15543,N_14842);
and U16644 (N_16644,N_15132,N_14486);
xnor U16645 (N_16645,N_14057,N_15927);
nand U16646 (N_16646,N_15050,N_15583);
or U16647 (N_16647,N_14280,N_14153);
nand U16648 (N_16648,N_14738,N_14259);
nor U16649 (N_16649,N_14185,N_14689);
or U16650 (N_16650,N_15938,N_14953);
or U16651 (N_16651,N_14682,N_15993);
xnor U16652 (N_16652,N_14764,N_15847);
nand U16653 (N_16653,N_15068,N_14244);
nand U16654 (N_16654,N_14985,N_14261);
nand U16655 (N_16655,N_14236,N_14497);
or U16656 (N_16656,N_14315,N_14435);
nand U16657 (N_16657,N_14092,N_15138);
nand U16658 (N_16658,N_14473,N_14155);
nor U16659 (N_16659,N_14209,N_15805);
and U16660 (N_16660,N_14797,N_14602);
nand U16661 (N_16661,N_15572,N_14592);
nor U16662 (N_16662,N_14800,N_15261);
or U16663 (N_16663,N_15785,N_15063);
nor U16664 (N_16664,N_15946,N_14880);
nor U16665 (N_16665,N_15461,N_14328);
nor U16666 (N_16666,N_15854,N_15070);
and U16667 (N_16667,N_15484,N_15715);
and U16668 (N_16668,N_14544,N_15145);
and U16669 (N_16669,N_15291,N_14808);
nor U16670 (N_16670,N_15351,N_14035);
xnor U16671 (N_16671,N_14081,N_14970);
or U16672 (N_16672,N_15780,N_14296);
nor U16673 (N_16673,N_15097,N_15897);
and U16674 (N_16674,N_15956,N_15967);
and U16675 (N_16675,N_14421,N_15397);
nor U16676 (N_16676,N_14614,N_15177);
or U16677 (N_16677,N_15518,N_14720);
nor U16678 (N_16678,N_14333,N_15188);
and U16679 (N_16679,N_15264,N_15186);
xor U16680 (N_16680,N_14135,N_14739);
and U16681 (N_16681,N_14655,N_14149);
and U16682 (N_16682,N_14505,N_15392);
nand U16683 (N_16683,N_15024,N_15719);
and U16684 (N_16684,N_15570,N_15424);
nand U16685 (N_16685,N_14719,N_15648);
and U16686 (N_16686,N_15267,N_15807);
or U16687 (N_16687,N_15472,N_14295);
nor U16688 (N_16688,N_15295,N_14981);
xor U16689 (N_16689,N_14010,N_15332);
xor U16690 (N_16690,N_14924,N_14448);
xor U16691 (N_16691,N_14378,N_15504);
and U16692 (N_16692,N_14843,N_14438);
nand U16693 (N_16693,N_15848,N_15039);
xor U16694 (N_16694,N_15275,N_14224);
nand U16695 (N_16695,N_15949,N_15427);
nor U16696 (N_16696,N_14667,N_15565);
nor U16697 (N_16697,N_15822,N_14252);
or U16698 (N_16698,N_14856,N_15473);
and U16699 (N_16699,N_15522,N_15552);
nor U16700 (N_16700,N_15265,N_15129);
or U16701 (N_16701,N_15880,N_15318);
nand U16702 (N_16702,N_14668,N_14825);
nand U16703 (N_16703,N_14799,N_14784);
and U16704 (N_16704,N_15348,N_15497);
nand U16705 (N_16705,N_15103,N_15012);
nor U16706 (N_16706,N_14220,N_15025);
nand U16707 (N_16707,N_14100,N_14895);
nor U16708 (N_16708,N_14265,N_14512);
nand U16709 (N_16709,N_14008,N_15541);
nand U16710 (N_16710,N_14337,N_14890);
nand U16711 (N_16711,N_15499,N_15429);
nand U16712 (N_16712,N_14430,N_14559);
xor U16713 (N_16713,N_14768,N_14749);
or U16714 (N_16714,N_14846,N_14893);
xor U16715 (N_16715,N_15366,N_15278);
or U16716 (N_16716,N_15874,N_15298);
xnor U16717 (N_16717,N_15559,N_15003);
nor U16718 (N_16718,N_15513,N_14860);
nor U16719 (N_16719,N_14940,N_14373);
and U16720 (N_16720,N_15995,N_15269);
xor U16721 (N_16721,N_14287,N_14458);
nand U16722 (N_16722,N_14160,N_15966);
or U16723 (N_16723,N_15125,N_14772);
or U16724 (N_16724,N_14453,N_14757);
or U16725 (N_16725,N_14212,N_15802);
nor U16726 (N_16726,N_15023,N_15118);
or U16727 (N_16727,N_14936,N_15959);
and U16728 (N_16728,N_14216,N_14351);
and U16729 (N_16729,N_14329,N_14511);
xnor U16730 (N_16730,N_14117,N_15293);
nand U16731 (N_16731,N_15274,N_14156);
or U16732 (N_16732,N_14130,N_14548);
nand U16733 (N_16733,N_15531,N_15401);
nor U16734 (N_16734,N_15971,N_14406);
nor U16735 (N_16735,N_14405,N_15574);
and U16736 (N_16736,N_14386,N_15910);
nand U16737 (N_16737,N_14635,N_15580);
and U16738 (N_16738,N_14729,N_15834);
nor U16739 (N_16739,N_15033,N_15173);
or U16740 (N_16740,N_14994,N_14792);
xor U16741 (N_16741,N_15622,N_14875);
and U16742 (N_16742,N_15727,N_15312);
nand U16743 (N_16743,N_15210,N_14891);
xnor U16744 (N_16744,N_14410,N_15526);
and U16745 (N_16745,N_15639,N_14721);
nor U16746 (N_16746,N_15953,N_14974);
or U16747 (N_16747,N_14502,N_15047);
and U16748 (N_16748,N_15555,N_14300);
and U16749 (N_16749,N_15317,N_14967);
nor U16750 (N_16750,N_15569,N_14566);
xnor U16751 (N_16751,N_15069,N_14173);
nand U16752 (N_16752,N_14877,N_14522);
nor U16753 (N_16753,N_14045,N_15977);
nor U16754 (N_16754,N_15767,N_14150);
xnor U16755 (N_16755,N_15309,N_14434);
and U16756 (N_16756,N_14688,N_15237);
xor U16757 (N_16757,N_14084,N_14681);
nand U16758 (N_16758,N_14989,N_14266);
xnor U16759 (N_16759,N_14444,N_15094);
and U16760 (N_16760,N_14172,N_14975);
or U16761 (N_16761,N_15517,N_14941);
xnor U16762 (N_16762,N_14617,N_15895);
and U16763 (N_16763,N_14157,N_14134);
or U16764 (N_16764,N_14829,N_14427);
nor U16765 (N_16765,N_15591,N_14312);
xnor U16766 (N_16766,N_14819,N_14247);
or U16767 (N_16767,N_15615,N_15823);
and U16768 (N_16768,N_14332,N_14396);
and U16769 (N_16769,N_14308,N_14474);
nor U16770 (N_16770,N_15169,N_14142);
xor U16771 (N_16771,N_14033,N_15933);
nand U16772 (N_16772,N_15706,N_15612);
nand U16773 (N_16773,N_14917,N_15659);
xnor U16774 (N_16774,N_14283,N_14992);
xor U16775 (N_16775,N_15660,N_14708);
or U16776 (N_16776,N_15339,N_14543);
or U16777 (N_16777,N_14168,N_14644);
and U16778 (N_16778,N_14969,N_15733);
or U16779 (N_16779,N_15257,N_14096);
nand U16780 (N_16780,N_14301,N_14769);
and U16781 (N_16781,N_14759,N_15750);
nor U16782 (N_16782,N_15191,N_14120);
or U16783 (N_16783,N_14004,N_14850);
nor U16784 (N_16784,N_14910,N_15788);
xor U16785 (N_16785,N_15850,N_14897);
xor U16786 (N_16786,N_14127,N_15259);
nand U16787 (N_16787,N_15343,N_14907);
or U16788 (N_16788,N_15975,N_14433);
or U16789 (N_16789,N_15126,N_15034);
and U16790 (N_16790,N_15123,N_14281);
and U16791 (N_16791,N_14600,N_15560);
nand U16792 (N_16792,N_14112,N_14830);
nand U16793 (N_16793,N_15398,N_15832);
nand U16794 (N_16794,N_15575,N_14240);
xor U16795 (N_16795,N_14823,N_15830);
nor U16796 (N_16796,N_14065,N_14557);
and U16797 (N_16797,N_14360,N_15046);
nor U16798 (N_16798,N_15013,N_15432);
and U16799 (N_16799,N_15774,N_15860);
xor U16800 (N_16800,N_14649,N_15276);
nand U16801 (N_16801,N_15588,N_14608);
or U16802 (N_16802,N_15113,N_15038);
xnor U16803 (N_16803,N_15634,N_14169);
nor U16804 (N_16804,N_15611,N_14441);
nand U16805 (N_16805,N_15281,N_14582);
and U16806 (N_16806,N_15626,N_14298);
nor U16807 (N_16807,N_15960,N_15431);
xnor U16808 (N_16808,N_15460,N_15662);
or U16809 (N_16809,N_15781,N_14822);
or U16810 (N_16810,N_14551,N_14088);
nand U16811 (N_16811,N_15596,N_15891);
nor U16812 (N_16812,N_14159,N_15604);
or U16813 (N_16813,N_14151,N_14276);
or U16814 (N_16814,N_14776,N_14049);
or U16815 (N_16815,N_15379,N_14233);
nor U16816 (N_16816,N_15983,N_14762);
xnor U16817 (N_16817,N_15271,N_14383);
and U16818 (N_16818,N_15841,N_15399);
nand U16819 (N_16819,N_14416,N_14026);
nor U16820 (N_16820,N_15148,N_15061);
xnor U16821 (N_16821,N_15940,N_15095);
xor U16822 (N_16822,N_14723,N_15152);
nor U16823 (N_16823,N_14750,N_15185);
nand U16824 (N_16824,N_15663,N_15336);
nor U16825 (N_16825,N_15909,N_15804);
or U16826 (N_16826,N_14961,N_14202);
xor U16827 (N_16827,N_14445,N_14179);
nand U16828 (N_16828,N_14107,N_15814);
nand U16829 (N_16829,N_14862,N_14536);
xor U16830 (N_16830,N_15892,N_14187);
nand U16831 (N_16831,N_14208,N_15172);
or U16832 (N_16832,N_15597,N_14865);
and U16833 (N_16833,N_15514,N_14167);
xnor U16834 (N_16834,N_14418,N_15335);
and U16835 (N_16835,N_14456,N_15144);
nand U16836 (N_16836,N_14211,N_15015);
and U16837 (N_16837,N_15623,N_15313);
nor U16838 (N_16838,N_15285,N_15230);
xor U16839 (N_16839,N_15700,N_15467);
and U16840 (N_16840,N_14102,N_14394);
nand U16841 (N_16841,N_15510,N_15711);
xor U16842 (N_16842,N_15606,N_14589);
nand U16843 (N_16843,N_14962,N_15714);
xor U16844 (N_16844,N_14878,N_14820);
nand U16845 (N_16845,N_14585,N_15307);
nor U16846 (N_16846,N_15287,N_14622);
and U16847 (N_16847,N_14498,N_14347);
or U16848 (N_16848,N_15724,N_14270);
or U16849 (N_16849,N_15821,N_14235);
xor U16850 (N_16850,N_14817,N_15951);
nand U16851 (N_16851,N_15978,N_15086);
or U16852 (N_16852,N_14226,N_14560);
nor U16853 (N_16853,N_14014,N_14174);
or U16854 (N_16854,N_14061,N_15487);
or U16855 (N_16855,N_14424,N_15551);
nor U16856 (N_16856,N_15691,N_14965);
nor U16857 (N_16857,N_15089,N_15608);
nand U16858 (N_16858,N_15459,N_14818);
nand U16859 (N_16859,N_14900,N_14192);
nand U16860 (N_16860,N_14113,N_15533);
nand U16861 (N_16861,N_15540,N_14481);
and U16862 (N_16862,N_15478,N_14884);
or U16863 (N_16863,N_14714,N_14083);
nor U16864 (N_16864,N_14698,N_15759);
nor U16865 (N_16865,N_14593,N_14693);
or U16866 (N_16866,N_15374,N_14623);
xnor U16867 (N_16867,N_15888,N_15981);
xnor U16868 (N_16868,N_15670,N_14645);
and U16869 (N_16869,N_14837,N_14076);
and U16870 (N_16870,N_14743,N_14472);
nor U16871 (N_16871,N_15315,N_15124);
nor U16872 (N_16872,N_15616,N_14338);
xnor U16873 (N_16873,N_15370,N_14887);
and U16874 (N_16874,N_14996,N_14902);
nor U16875 (N_16875,N_14345,N_15300);
xnor U16876 (N_16876,N_14633,N_15942);
nor U16877 (N_16877,N_15243,N_14526);
xnor U16878 (N_16878,N_15450,N_15722);
or U16879 (N_16879,N_14619,N_14001);
xnor U16880 (N_16880,N_15327,N_15416);
nor U16881 (N_16881,N_14660,N_14464);
nand U16882 (N_16882,N_15875,N_14007);
nor U16883 (N_16883,N_14954,N_14755);
nor U16884 (N_16884,N_15437,N_14590);
or U16885 (N_16885,N_14245,N_14119);
and U16886 (N_16886,N_14726,N_14848);
nand U16887 (N_16887,N_15859,N_14016);
nor U16888 (N_16888,N_15758,N_14747);
or U16889 (N_16889,N_14392,N_14794);
xnor U16890 (N_16890,N_14183,N_14756);
xnor U16891 (N_16891,N_15797,N_14946);
and U16892 (N_16892,N_15007,N_14462);
nor U16893 (N_16893,N_14115,N_15310);
or U16894 (N_16894,N_14957,N_14615);
or U16895 (N_16895,N_14628,N_15952);
nand U16896 (N_16896,N_15241,N_15263);
nand U16897 (N_16897,N_14581,N_14475);
and U16898 (N_16898,N_14651,N_14352);
and U16899 (N_16899,N_15760,N_15405);
or U16900 (N_16900,N_15272,N_14631);
nor U16901 (N_16901,N_14425,N_15463);
xor U16902 (N_16902,N_14964,N_15029);
or U16903 (N_16903,N_15982,N_14431);
xor U16904 (N_16904,N_15128,N_15654);
nand U16905 (N_16905,N_14361,N_15236);
nand U16906 (N_16906,N_15027,N_15912);
nand U16907 (N_16907,N_15868,N_15053);
and U16908 (N_16908,N_14573,N_15227);
or U16909 (N_16909,N_14844,N_14180);
xor U16910 (N_16910,N_14376,N_14650);
and U16911 (N_16911,N_14709,N_14289);
nand U16912 (N_16912,N_15420,N_14986);
nor U16913 (N_16913,N_15077,N_15455);
and U16914 (N_16914,N_15685,N_14643);
nand U16915 (N_16915,N_14773,N_14020);
xnor U16916 (N_16916,N_15755,N_15669);
or U16917 (N_16917,N_15941,N_15159);
or U16918 (N_16918,N_15725,N_14782);
nor U16919 (N_16919,N_15505,N_15997);
xnor U16920 (N_16920,N_15319,N_14809);
xor U16921 (N_16921,N_14565,N_15819);
and U16922 (N_16922,N_14182,N_15916);
or U16923 (N_16923,N_15745,N_15954);
and U16924 (N_16924,N_15766,N_15164);
xnor U16925 (N_16925,N_15906,N_15182);
nor U16926 (N_16926,N_14587,N_15932);
xor U16927 (N_16927,N_15109,N_15625);
nand U16928 (N_16928,N_14678,N_14583);
or U16929 (N_16929,N_15707,N_14778);
nor U16930 (N_16930,N_15931,N_15058);
nor U16931 (N_16931,N_14934,N_15498);
nand U16932 (N_16932,N_15223,N_15748);
xor U16933 (N_16933,N_14099,N_15955);
nor U16934 (N_16934,N_15167,N_15075);
or U16935 (N_16935,N_15680,N_14673);
nand U16936 (N_16936,N_15585,N_14171);
xnor U16937 (N_16937,N_14697,N_14258);
xor U16938 (N_16938,N_14849,N_14999);
or U16939 (N_16939,N_15454,N_15957);
nand U16940 (N_16940,N_14480,N_15686);
nand U16941 (N_16941,N_14342,N_14034);
nor U16942 (N_16942,N_15632,N_15056);
and U16943 (N_16943,N_15581,N_15631);
or U16944 (N_16944,N_15576,N_15593);
and U16945 (N_16945,N_15742,N_15994);
nand U16946 (N_16946,N_14701,N_14241);
or U16947 (N_16947,N_15283,N_14627);
nand U16948 (N_16948,N_14935,N_14108);
xor U16949 (N_16949,N_14093,N_14508);
or U16950 (N_16950,N_14597,N_14073);
or U16951 (N_16951,N_14359,N_15154);
nand U16952 (N_16952,N_15306,N_15375);
nand U16953 (N_16953,N_15687,N_14451);
xnor U16954 (N_16954,N_14766,N_14412);
or U16955 (N_16955,N_15723,N_14926);
xor U16956 (N_16956,N_15279,N_14767);
xnor U16957 (N_16957,N_14449,N_14562);
and U16958 (N_16958,N_15107,N_15735);
or U16959 (N_16959,N_14779,N_14609);
or U16960 (N_16960,N_14263,N_15664);
or U16961 (N_16961,N_15635,N_15449);
xnor U16962 (N_16962,N_15357,N_15520);
nand U16963 (N_16963,N_14728,N_15211);
nand U16964 (N_16964,N_14718,N_14618);
or U16965 (N_16965,N_14826,N_15384);
nor U16966 (N_16966,N_15528,N_14413);
and U16967 (N_16967,N_14097,N_15539);
xor U16968 (N_16968,N_15769,N_15362);
xnor U16969 (N_16969,N_15968,N_15884);
or U16970 (N_16970,N_15112,N_15798);
nand U16971 (N_16971,N_14395,N_15493);
xnor U16972 (N_16972,N_14024,N_14516);
nand U16973 (N_16973,N_14322,N_14575);
or U16974 (N_16974,N_15444,N_14484);
nand U16975 (N_16975,N_15728,N_15489);
and U16976 (N_16976,N_14483,N_14939);
nand U16977 (N_16977,N_15458,N_15101);
nor U16978 (N_16978,N_14382,N_14303);
and U16979 (N_16979,N_15810,N_15827);
xnor U16980 (N_16980,N_15088,N_15636);
nand U16981 (N_16981,N_15911,N_14366);
and U16982 (N_16982,N_15737,N_14691);
xnor U16983 (N_16983,N_14468,N_14367);
xor U16984 (N_16984,N_14331,N_14248);
and U16985 (N_16985,N_14426,N_15872);
and U16986 (N_16986,N_14353,N_15647);
nor U16987 (N_16987,N_14546,N_14730);
and U16988 (N_16988,N_15600,N_15930);
or U16989 (N_16989,N_15065,N_14304);
or U16990 (N_16990,N_15833,N_14658);
nand U16991 (N_16991,N_15732,N_14118);
and U16992 (N_16992,N_15839,N_15316);
xor U16993 (N_16993,N_14177,N_15871);
xnor U16994 (N_16994,N_14385,N_15702);
and U16995 (N_16995,N_14306,N_15041);
or U16996 (N_16996,N_15984,N_14085);
or U16997 (N_16997,N_14541,N_14685);
xor U16998 (N_16998,N_15556,N_15492);
nand U16999 (N_16999,N_14237,N_15108);
and U17000 (N_17000,N_15044,N_14136);
nor U17001 (N_17001,N_14149,N_15266);
or U17002 (N_17002,N_14103,N_14074);
nor U17003 (N_17003,N_14890,N_15740);
and U17004 (N_17004,N_14151,N_15942);
or U17005 (N_17005,N_14600,N_15549);
and U17006 (N_17006,N_14549,N_14096);
and U17007 (N_17007,N_15033,N_15908);
nand U17008 (N_17008,N_15537,N_15512);
nor U17009 (N_17009,N_15067,N_15176);
nor U17010 (N_17010,N_15794,N_14928);
nor U17011 (N_17011,N_15436,N_14249);
or U17012 (N_17012,N_14996,N_15092);
nand U17013 (N_17013,N_14730,N_15742);
xnor U17014 (N_17014,N_15648,N_14167);
nand U17015 (N_17015,N_15449,N_14181);
xnor U17016 (N_17016,N_14133,N_14071);
or U17017 (N_17017,N_15716,N_15026);
xor U17018 (N_17018,N_15983,N_15381);
nor U17019 (N_17019,N_14150,N_14289);
nor U17020 (N_17020,N_15272,N_14645);
and U17021 (N_17021,N_15390,N_14339);
and U17022 (N_17022,N_15669,N_14453);
xor U17023 (N_17023,N_14660,N_14701);
nand U17024 (N_17024,N_14506,N_15857);
xor U17025 (N_17025,N_14026,N_15942);
nor U17026 (N_17026,N_14045,N_15972);
and U17027 (N_17027,N_15993,N_15803);
xnor U17028 (N_17028,N_15235,N_14903);
xnor U17029 (N_17029,N_15028,N_15659);
nor U17030 (N_17030,N_14686,N_15846);
nor U17031 (N_17031,N_14037,N_14626);
nor U17032 (N_17032,N_15961,N_14839);
xor U17033 (N_17033,N_14964,N_14606);
or U17034 (N_17034,N_14180,N_15942);
or U17035 (N_17035,N_15316,N_14656);
or U17036 (N_17036,N_15164,N_14381);
xor U17037 (N_17037,N_15141,N_15450);
or U17038 (N_17038,N_15748,N_14808);
or U17039 (N_17039,N_15098,N_14115);
xor U17040 (N_17040,N_15237,N_14788);
and U17041 (N_17041,N_15809,N_15742);
nor U17042 (N_17042,N_15593,N_14201);
nor U17043 (N_17043,N_14549,N_15352);
nand U17044 (N_17044,N_14164,N_14439);
and U17045 (N_17045,N_14090,N_15135);
xnor U17046 (N_17046,N_14400,N_15464);
xor U17047 (N_17047,N_14739,N_15126);
or U17048 (N_17048,N_15394,N_14595);
nand U17049 (N_17049,N_15207,N_14554);
xor U17050 (N_17050,N_14663,N_15045);
and U17051 (N_17051,N_14160,N_15226);
nand U17052 (N_17052,N_15199,N_14372);
and U17053 (N_17053,N_15334,N_15384);
xnor U17054 (N_17054,N_15841,N_14186);
and U17055 (N_17055,N_15605,N_15438);
and U17056 (N_17056,N_14781,N_15814);
nor U17057 (N_17057,N_15966,N_14593);
nor U17058 (N_17058,N_15418,N_15232);
nand U17059 (N_17059,N_15301,N_15264);
nor U17060 (N_17060,N_15081,N_15639);
or U17061 (N_17061,N_14225,N_15695);
nand U17062 (N_17062,N_15201,N_14442);
xnor U17063 (N_17063,N_15529,N_15591);
nor U17064 (N_17064,N_14793,N_15634);
nor U17065 (N_17065,N_15685,N_15155);
and U17066 (N_17066,N_15452,N_15953);
or U17067 (N_17067,N_15989,N_15326);
or U17068 (N_17068,N_14411,N_14304);
xor U17069 (N_17069,N_15305,N_15062);
xor U17070 (N_17070,N_14037,N_14375);
or U17071 (N_17071,N_15987,N_15185);
xnor U17072 (N_17072,N_14297,N_15778);
xor U17073 (N_17073,N_15216,N_14604);
nand U17074 (N_17074,N_14080,N_15403);
xor U17075 (N_17075,N_15703,N_15483);
xor U17076 (N_17076,N_15603,N_14806);
nand U17077 (N_17077,N_15002,N_15830);
or U17078 (N_17078,N_14939,N_15331);
nor U17079 (N_17079,N_14259,N_15846);
nor U17080 (N_17080,N_14709,N_15786);
and U17081 (N_17081,N_14130,N_15436);
and U17082 (N_17082,N_14114,N_15048);
or U17083 (N_17083,N_15462,N_15366);
and U17084 (N_17084,N_14114,N_15923);
or U17085 (N_17085,N_15930,N_15806);
xnor U17086 (N_17086,N_14846,N_15991);
nor U17087 (N_17087,N_15096,N_14804);
nor U17088 (N_17088,N_15855,N_14470);
or U17089 (N_17089,N_15701,N_14955);
nand U17090 (N_17090,N_14824,N_15400);
and U17091 (N_17091,N_15947,N_14904);
xnor U17092 (N_17092,N_14902,N_15856);
or U17093 (N_17093,N_15265,N_15699);
xnor U17094 (N_17094,N_15832,N_14247);
xor U17095 (N_17095,N_15963,N_15006);
and U17096 (N_17096,N_15839,N_14379);
or U17097 (N_17097,N_14563,N_14596);
and U17098 (N_17098,N_15998,N_14910);
nand U17099 (N_17099,N_14360,N_14755);
or U17100 (N_17100,N_15658,N_14593);
and U17101 (N_17101,N_14903,N_15045);
xnor U17102 (N_17102,N_14798,N_15937);
and U17103 (N_17103,N_15690,N_14670);
and U17104 (N_17104,N_15921,N_15859);
xor U17105 (N_17105,N_15131,N_15628);
nor U17106 (N_17106,N_15609,N_14869);
nor U17107 (N_17107,N_15913,N_15425);
nor U17108 (N_17108,N_14054,N_14975);
and U17109 (N_17109,N_14001,N_14512);
and U17110 (N_17110,N_15491,N_14551);
nand U17111 (N_17111,N_15490,N_14457);
nor U17112 (N_17112,N_14274,N_15537);
or U17113 (N_17113,N_15252,N_15845);
xor U17114 (N_17114,N_15372,N_15130);
and U17115 (N_17115,N_14945,N_14801);
xnor U17116 (N_17116,N_15574,N_15420);
nand U17117 (N_17117,N_15661,N_15424);
nand U17118 (N_17118,N_14885,N_15250);
nand U17119 (N_17119,N_14338,N_14343);
xnor U17120 (N_17120,N_14285,N_15946);
nand U17121 (N_17121,N_14812,N_15903);
xor U17122 (N_17122,N_15810,N_14939);
and U17123 (N_17123,N_15049,N_15740);
nand U17124 (N_17124,N_15272,N_14881);
nand U17125 (N_17125,N_15331,N_14689);
nor U17126 (N_17126,N_14299,N_15244);
nor U17127 (N_17127,N_14945,N_15539);
or U17128 (N_17128,N_14448,N_14041);
nand U17129 (N_17129,N_14345,N_14043);
or U17130 (N_17130,N_14543,N_14494);
xnor U17131 (N_17131,N_14884,N_14957);
nand U17132 (N_17132,N_14791,N_14298);
nand U17133 (N_17133,N_15269,N_14291);
nand U17134 (N_17134,N_15919,N_15560);
nor U17135 (N_17135,N_15300,N_15174);
nand U17136 (N_17136,N_15850,N_14436);
and U17137 (N_17137,N_15058,N_14319);
nand U17138 (N_17138,N_14085,N_15765);
or U17139 (N_17139,N_15140,N_15250);
and U17140 (N_17140,N_15304,N_14536);
and U17141 (N_17141,N_14920,N_14973);
nand U17142 (N_17142,N_15907,N_14342);
nor U17143 (N_17143,N_15783,N_14906);
and U17144 (N_17144,N_14368,N_14932);
xnor U17145 (N_17145,N_15497,N_14295);
and U17146 (N_17146,N_15141,N_14138);
or U17147 (N_17147,N_15193,N_14782);
xor U17148 (N_17148,N_15813,N_15401);
xnor U17149 (N_17149,N_15207,N_15390);
nand U17150 (N_17150,N_15027,N_14521);
or U17151 (N_17151,N_15569,N_15896);
xnor U17152 (N_17152,N_15334,N_15980);
nor U17153 (N_17153,N_15633,N_15119);
or U17154 (N_17154,N_15856,N_14376);
or U17155 (N_17155,N_15959,N_14174);
or U17156 (N_17156,N_15622,N_14944);
xor U17157 (N_17157,N_14719,N_15263);
nand U17158 (N_17158,N_14615,N_15266);
nand U17159 (N_17159,N_14667,N_14790);
xor U17160 (N_17160,N_15545,N_14044);
nand U17161 (N_17161,N_15685,N_15462);
or U17162 (N_17162,N_14981,N_14053);
xnor U17163 (N_17163,N_15142,N_14443);
nor U17164 (N_17164,N_14686,N_14894);
xnor U17165 (N_17165,N_15982,N_15537);
xor U17166 (N_17166,N_14103,N_14723);
xor U17167 (N_17167,N_14452,N_14389);
nand U17168 (N_17168,N_14628,N_14153);
nand U17169 (N_17169,N_14403,N_14659);
and U17170 (N_17170,N_15057,N_14005);
nor U17171 (N_17171,N_15297,N_14829);
nor U17172 (N_17172,N_14325,N_14766);
nor U17173 (N_17173,N_15311,N_14332);
nor U17174 (N_17174,N_14318,N_15675);
xor U17175 (N_17175,N_15950,N_14734);
and U17176 (N_17176,N_15490,N_14434);
nor U17177 (N_17177,N_15896,N_14055);
nor U17178 (N_17178,N_14470,N_14186);
nand U17179 (N_17179,N_14538,N_15441);
or U17180 (N_17180,N_15629,N_14760);
and U17181 (N_17181,N_15664,N_15612);
and U17182 (N_17182,N_14509,N_14053);
and U17183 (N_17183,N_15663,N_15324);
and U17184 (N_17184,N_14567,N_14058);
nor U17185 (N_17185,N_15708,N_14588);
xor U17186 (N_17186,N_14430,N_14261);
nand U17187 (N_17187,N_14660,N_15296);
xnor U17188 (N_17188,N_15203,N_15253);
nor U17189 (N_17189,N_15276,N_15742);
and U17190 (N_17190,N_15008,N_15362);
and U17191 (N_17191,N_14340,N_15686);
nor U17192 (N_17192,N_15603,N_15856);
nand U17193 (N_17193,N_14104,N_14072);
or U17194 (N_17194,N_15191,N_14634);
nor U17195 (N_17195,N_15603,N_15162);
nand U17196 (N_17196,N_15815,N_14488);
nor U17197 (N_17197,N_15641,N_15358);
nand U17198 (N_17198,N_15563,N_14375);
and U17199 (N_17199,N_14517,N_14113);
xnor U17200 (N_17200,N_15833,N_14739);
and U17201 (N_17201,N_15630,N_15750);
or U17202 (N_17202,N_15980,N_15016);
and U17203 (N_17203,N_15280,N_15869);
nand U17204 (N_17204,N_15797,N_14062);
and U17205 (N_17205,N_15379,N_15758);
nor U17206 (N_17206,N_15722,N_14411);
nor U17207 (N_17207,N_15445,N_15041);
nand U17208 (N_17208,N_14535,N_15776);
nor U17209 (N_17209,N_14135,N_15664);
xnor U17210 (N_17210,N_14917,N_14955);
xor U17211 (N_17211,N_14009,N_15091);
xnor U17212 (N_17212,N_14191,N_15868);
xor U17213 (N_17213,N_15377,N_15111);
nand U17214 (N_17214,N_14305,N_15354);
nor U17215 (N_17215,N_14074,N_14472);
or U17216 (N_17216,N_14093,N_15688);
or U17217 (N_17217,N_14985,N_15139);
xor U17218 (N_17218,N_15731,N_14606);
or U17219 (N_17219,N_14561,N_14888);
or U17220 (N_17220,N_15017,N_15996);
nand U17221 (N_17221,N_15771,N_14808);
xnor U17222 (N_17222,N_15545,N_15633);
xnor U17223 (N_17223,N_15851,N_15496);
nor U17224 (N_17224,N_14258,N_14480);
xnor U17225 (N_17225,N_15657,N_14422);
xor U17226 (N_17226,N_15250,N_15630);
nor U17227 (N_17227,N_15228,N_15893);
or U17228 (N_17228,N_15991,N_15792);
or U17229 (N_17229,N_15981,N_14187);
xor U17230 (N_17230,N_14440,N_14024);
or U17231 (N_17231,N_15502,N_15553);
nand U17232 (N_17232,N_15169,N_14841);
nor U17233 (N_17233,N_15473,N_15630);
nand U17234 (N_17234,N_15304,N_15799);
nand U17235 (N_17235,N_14909,N_14319);
nor U17236 (N_17236,N_14245,N_15182);
or U17237 (N_17237,N_14505,N_15981);
nand U17238 (N_17238,N_15987,N_14869);
nor U17239 (N_17239,N_14199,N_14851);
and U17240 (N_17240,N_14371,N_14621);
nor U17241 (N_17241,N_14579,N_14867);
nor U17242 (N_17242,N_14851,N_14681);
nor U17243 (N_17243,N_15785,N_14900);
and U17244 (N_17244,N_15561,N_15198);
nand U17245 (N_17245,N_15862,N_15895);
and U17246 (N_17246,N_15014,N_14322);
or U17247 (N_17247,N_14648,N_15352);
nand U17248 (N_17248,N_15200,N_15390);
or U17249 (N_17249,N_15939,N_14388);
xor U17250 (N_17250,N_15494,N_15251);
nand U17251 (N_17251,N_14279,N_15089);
nor U17252 (N_17252,N_14593,N_14080);
or U17253 (N_17253,N_15093,N_14295);
or U17254 (N_17254,N_15162,N_15822);
nand U17255 (N_17255,N_14150,N_15207);
xnor U17256 (N_17256,N_14443,N_14436);
and U17257 (N_17257,N_15651,N_14921);
nand U17258 (N_17258,N_15636,N_14655);
and U17259 (N_17259,N_15489,N_14509);
nor U17260 (N_17260,N_14253,N_15893);
nor U17261 (N_17261,N_15051,N_15159);
or U17262 (N_17262,N_15876,N_14309);
xor U17263 (N_17263,N_15012,N_14237);
nor U17264 (N_17264,N_14831,N_15513);
xor U17265 (N_17265,N_15610,N_14935);
xnor U17266 (N_17266,N_14578,N_15223);
or U17267 (N_17267,N_14944,N_14488);
nand U17268 (N_17268,N_14919,N_15696);
xnor U17269 (N_17269,N_14959,N_15351);
or U17270 (N_17270,N_14687,N_15425);
nor U17271 (N_17271,N_15889,N_15770);
nor U17272 (N_17272,N_14458,N_14226);
or U17273 (N_17273,N_15105,N_14808);
xnor U17274 (N_17274,N_15448,N_14184);
nor U17275 (N_17275,N_15284,N_15729);
and U17276 (N_17276,N_14797,N_14210);
or U17277 (N_17277,N_15038,N_15852);
or U17278 (N_17278,N_14853,N_14392);
xor U17279 (N_17279,N_15589,N_14696);
nor U17280 (N_17280,N_15628,N_15045);
nand U17281 (N_17281,N_15903,N_14908);
xnor U17282 (N_17282,N_15542,N_15575);
or U17283 (N_17283,N_15296,N_14054);
or U17284 (N_17284,N_14559,N_15525);
and U17285 (N_17285,N_15686,N_15737);
nor U17286 (N_17286,N_15449,N_14985);
nand U17287 (N_17287,N_14038,N_14479);
xnor U17288 (N_17288,N_14287,N_14026);
and U17289 (N_17289,N_14006,N_14556);
nand U17290 (N_17290,N_15292,N_15981);
and U17291 (N_17291,N_14181,N_14008);
xnor U17292 (N_17292,N_14731,N_15944);
or U17293 (N_17293,N_14463,N_15596);
and U17294 (N_17294,N_14100,N_15403);
nor U17295 (N_17295,N_15449,N_15622);
xor U17296 (N_17296,N_14786,N_14625);
nand U17297 (N_17297,N_14476,N_14872);
or U17298 (N_17298,N_15382,N_15779);
nand U17299 (N_17299,N_14018,N_15412);
and U17300 (N_17300,N_15949,N_15607);
and U17301 (N_17301,N_14582,N_15598);
nand U17302 (N_17302,N_15031,N_15578);
nor U17303 (N_17303,N_14103,N_15287);
and U17304 (N_17304,N_15082,N_14576);
xor U17305 (N_17305,N_15251,N_15691);
and U17306 (N_17306,N_14853,N_14965);
and U17307 (N_17307,N_15586,N_15037);
nor U17308 (N_17308,N_15816,N_14820);
and U17309 (N_17309,N_15171,N_14195);
and U17310 (N_17310,N_15260,N_15214);
xnor U17311 (N_17311,N_14380,N_14531);
nand U17312 (N_17312,N_14571,N_14416);
or U17313 (N_17313,N_15432,N_14639);
and U17314 (N_17314,N_14580,N_15379);
or U17315 (N_17315,N_14395,N_14569);
nand U17316 (N_17316,N_15089,N_14976);
or U17317 (N_17317,N_15258,N_14478);
nand U17318 (N_17318,N_15206,N_15661);
nand U17319 (N_17319,N_15438,N_14857);
xnor U17320 (N_17320,N_14818,N_14605);
nand U17321 (N_17321,N_15372,N_14028);
and U17322 (N_17322,N_14148,N_14682);
nor U17323 (N_17323,N_14548,N_15187);
nand U17324 (N_17324,N_14063,N_15883);
nand U17325 (N_17325,N_15363,N_15950);
or U17326 (N_17326,N_14379,N_14697);
nand U17327 (N_17327,N_15580,N_15989);
nor U17328 (N_17328,N_14872,N_15845);
nand U17329 (N_17329,N_14695,N_14138);
and U17330 (N_17330,N_14339,N_15755);
and U17331 (N_17331,N_15488,N_15564);
nand U17332 (N_17332,N_14894,N_14287);
nor U17333 (N_17333,N_15630,N_14452);
xnor U17334 (N_17334,N_14704,N_14604);
nor U17335 (N_17335,N_15736,N_15359);
and U17336 (N_17336,N_14164,N_14881);
nor U17337 (N_17337,N_14685,N_15421);
or U17338 (N_17338,N_14986,N_14377);
nand U17339 (N_17339,N_15428,N_15205);
nand U17340 (N_17340,N_14843,N_14372);
xnor U17341 (N_17341,N_15434,N_14607);
xor U17342 (N_17342,N_14269,N_15660);
and U17343 (N_17343,N_14207,N_15778);
nor U17344 (N_17344,N_15430,N_14207);
nor U17345 (N_17345,N_14917,N_14478);
or U17346 (N_17346,N_14511,N_15454);
and U17347 (N_17347,N_15075,N_14640);
nand U17348 (N_17348,N_15659,N_15438);
xor U17349 (N_17349,N_15169,N_15215);
nor U17350 (N_17350,N_14335,N_14745);
xor U17351 (N_17351,N_15524,N_14786);
and U17352 (N_17352,N_14492,N_14168);
or U17353 (N_17353,N_14611,N_15786);
nor U17354 (N_17354,N_14579,N_14280);
xor U17355 (N_17355,N_14273,N_15196);
xor U17356 (N_17356,N_14797,N_14960);
nor U17357 (N_17357,N_15504,N_14241);
nor U17358 (N_17358,N_15094,N_15947);
nor U17359 (N_17359,N_15733,N_15199);
xor U17360 (N_17360,N_15223,N_14099);
or U17361 (N_17361,N_14839,N_14671);
nand U17362 (N_17362,N_15701,N_15370);
or U17363 (N_17363,N_14763,N_14788);
nand U17364 (N_17364,N_15301,N_14731);
nor U17365 (N_17365,N_15441,N_15553);
nand U17366 (N_17366,N_15616,N_14522);
nand U17367 (N_17367,N_15827,N_15603);
nand U17368 (N_17368,N_15293,N_15000);
nor U17369 (N_17369,N_15868,N_15861);
or U17370 (N_17370,N_14440,N_15435);
xnor U17371 (N_17371,N_14739,N_15803);
nor U17372 (N_17372,N_15748,N_14386);
nand U17373 (N_17373,N_14895,N_15107);
nand U17374 (N_17374,N_14779,N_15721);
or U17375 (N_17375,N_14533,N_15475);
or U17376 (N_17376,N_14275,N_14461);
or U17377 (N_17377,N_14775,N_14186);
and U17378 (N_17378,N_15700,N_15073);
or U17379 (N_17379,N_14796,N_15910);
nor U17380 (N_17380,N_15791,N_14065);
and U17381 (N_17381,N_15529,N_14772);
or U17382 (N_17382,N_15421,N_15039);
nor U17383 (N_17383,N_14240,N_14119);
nor U17384 (N_17384,N_15468,N_14292);
or U17385 (N_17385,N_14991,N_15931);
nand U17386 (N_17386,N_14147,N_14682);
and U17387 (N_17387,N_15715,N_15737);
nor U17388 (N_17388,N_14182,N_15106);
or U17389 (N_17389,N_14329,N_15224);
nand U17390 (N_17390,N_15249,N_15869);
nor U17391 (N_17391,N_15179,N_15751);
xnor U17392 (N_17392,N_15654,N_14342);
xnor U17393 (N_17393,N_15032,N_15125);
xnor U17394 (N_17394,N_15279,N_14871);
and U17395 (N_17395,N_15353,N_15785);
or U17396 (N_17396,N_14294,N_14384);
nand U17397 (N_17397,N_14263,N_14795);
xor U17398 (N_17398,N_14323,N_15120);
or U17399 (N_17399,N_15336,N_15785);
or U17400 (N_17400,N_15876,N_15833);
and U17401 (N_17401,N_15587,N_15388);
nand U17402 (N_17402,N_14161,N_15057);
and U17403 (N_17403,N_15333,N_14195);
and U17404 (N_17404,N_14998,N_15911);
nand U17405 (N_17405,N_14592,N_15760);
nor U17406 (N_17406,N_15042,N_15144);
nor U17407 (N_17407,N_14080,N_14545);
nor U17408 (N_17408,N_14752,N_15047);
nand U17409 (N_17409,N_14072,N_15850);
nor U17410 (N_17410,N_14119,N_14169);
nand U17411 (N_17411,N_15936,N_14272);
nand U17412 (N_17412,N_15309,N_14516);
or U17413 (N_17413,N_15008,N_14745);
and U17414 (N_17414,N_14145,N_15622);
and U17415 (N_17415,N_15813,N_14860);
nor U17416 (N_17416,N_15494,N_14996);
or U17417 (N_17417,N_14666,N_15559);
or U17418 (N_17418,N_15719,N_15390);
nor U17419 (N_17419,N_14478,N_15957);
nand U17420 (N_17420,N_14979,N_14276);
nand U17421 (N_17421,N_15494,N_14804);
or U17422 (N_17422,N_14988,N_14911);
nor U17423 (N_17423,N_14026,N_14389);
nor U17424 (N_17424,N_14658,N_15116);
or U17425 (N_17425,N_15764,N_14884);
nand U17426 (N_17426,N_15924,N_15641);
nor U17427 (N_17427,N_15819,N_14370);
and U17428 (N_17428,N_15583,N_14795);
nand U17429 (N_17429,N_15439,N_14575);
nand U17430 (N_17430,N_14076,N_15037);
nand U17431 (N_17431,N_15864,N_14580);
nand U17432 (N_17432,N_14417,N_14651);
or U17433 (N_17433,N_14326,N_14415);
and U17434 (N_17434,N_14277,N_14757);
nor U17435 (N_17435,N_14990,N_14921);
or U17436 (N_17436,N_15551,N_15626);
or U17437 (N_17437,N_14193,N_14435);
or U17438 (N_17438,N_15019,N_15655);
or U17439 (N_17439,N_15559,N_14515);
and U17440 (N_17440,N_15112,N_15239);
nand U17441 (N_17441,N_14355,N_15583);
and U17442 (N_17442,N_15392,N_15126);
nor U17443 (N_17443,N_14276,N_15515);
xor U17444 (N_17444,N_15761,N_14816);
and U17445 (N_17445,N_15816,N_15800);
nand U17446 (N_17446,N_15516,N_14750);
or U17447 (N_17447,N_15473,N_15184);
xnor U17448 (N_17448,N_14320,N_15635);
and U17449 (N_17449,N_15903,N_14739);
and U17450 (N_17450,N_15363,N_15089);
nand U17451 (N_17451,N_14963,N_14108);
xor U17452 (N_17452,N_14800,N_14235);
or U17453 (N_17453,N_15237,N_15219);
and U17454 (N_17454,N_15794,N_15361);
xor U17455 (N_17455,N_14013,N_15146);
xnor U17456 (N_17456,N_15920,N_14064);
nand U17457 (N_17457,N_15471,N_14238);
and U17458 (N_17458,N_15523,N_14982);
and U17459 (N_17459,N_15364,N_14980);
and U17460 (N_17460,N_15565,N_15629);
nor U17461 (N_17461,N_14845,N_15873);
and U17462 (N_17462,N_15524,N_14155);
nor U17463 (N_17463,N_14782,N_15504);
or U17464 (N_17464,N_14721,N_14873);
and U17465 (N_17465,N_14164,N_14039);
nand U17466 (N_17466,N_14534,N_14488);
xnor U17467 (N_17467,N_15860,N_15465);
and U17468 (N_17468,N_14832,N_15516);
xor U17469 (N_17469,N_15532,N_14127);
nand U17470 (N_17470,N_14914,N_14057);
nand U17471 (N_17471,N_14962,N_14922);
nand U17472 (N_17472,N_14944,N_14743);
nor U17473 (N_17473,N_14505,N_15724);
or U17474 (N_17474,N_15617,N_15194);
nor U17475 (N_17475,N_14293,N_14553);
nand U17476 (N_17476,N_14685,N_15496);
xnor U17477 (N_17477,N_15475,N_14750);
or U17478 (N_17478,N_14162,N_15032);
nor U17479 (N_17479,N_14210,N_14787);
or U17480 (N_17480,N_14019,N_15587);
and U17481 (N_17481,N_15831,N_15294);
nor U17482 (N_17482,N_14378,N_14112);
and U17483 (N_17483,N_14110,N_14146);
xor U17484 (N_17484,N_14613,N_14597);
and U17485 (N_17485,N_15556,N_15408);
xor U17486 (N_17486,N_15844,N_14887);
nand U17487 (N_17487,N_15303,N_15524);
nor U17488 (N_17488,N_14997,N_14315);
xor U17489 (N_17489,N_15140,N_15849);
and U17490 (N_17490,N_14434,N_14274);
nor U17491 (N_17491,N_14450,N_15142);
nand U17492 (N_17492,N_14713,N_15939);
and U17493 (N_17493,N_14470,N_15220);
nor U17494 (N_17494,N_15648,N_14215);
nand U17495 (N_17495,N_14429,N_14017);
and U17496 (N_17496,N_15837,N_14916);
xor U17497 (N_17497,N_14860,N_14137);
nor U17498 (N_17498,N_15841,N_14035);
and U17499 (N_17499,N_15669,N_14681);
and U17500 (N_17500,N_14850,N_14596);
xor U17501 (N_17501,N_15656,N_14494);
xor U17502 (N_17502,N_15380,N_14024);
nand U17503 (N_17503,N_15608,N_15499);
nand U17504 (N_17504,N_14897,N_15394);
xnor U17505 (N_17505,N_14456,N_15819);
or U17506 (N_17506,N_14281,N_15487);
nor U17507 (N_17507,N_15367,N_15067);
nor U17508 (N_17508,N_14927,N_14632);
nor U17509 (N_17509,N_14739,N_15682);
or U17510 (N_17510,N_15678,N_15017);
and U17511 (N_17511,N_14340,N_15381);
xnor U17512 (N_17512,N_14749,N_14935);
and U17513 (N_17513,N_14456,N_14236);
and U17514 (N_17514,N_15981,N_14424);
xor U17515 (N_17515,N_15763,N_15089);
xnor U17516 (N_17516,N_15499,N_14531);
xnor U17517 (N_17517,N_15118,N_15525);
and U17518 (N_17518,N_14297,N_15569);
nor U17519 (N_17519,N_14091,N_15198);
xnor U17520 (N_17520,N_15105,N_14784);
and U17521 (N_17521,N_14422,N_15561);
or U17522 (N_17522,N_15111,N_14066);
or U17523 (N_17523,N_15589,N_15043);
or U17524 (N_17524,N_15490,N_14017);
nor U17525 (N_17525,N_15736,N_15389);
and U17526 (N_17526,N_15418,N_15249);
nor U17527 (N_17527,N_14863,N_14420);
or U17528 (N_17528,N_15169,N_14764);
or U17529 (N_17529,N_15361,N_14396);
nand U17530 (N_17530,N_14668,N_14271);
xnor U17531 (N_17531,N_15664,N_15002);
or U17532 (N_17532,N_15248,N_15164);
nor U17533 (N_17533,N_14690,N_15358);
and U17534 (N_17534,N_15324,N_15849);
or U17535 (N_17535,N_14921,N_15579);
nand U17536 (N_17536,N_15457,N_14650);
and U17537 (N_17537,N_14164,N_14233);
nor U17538 (N_17538,N_15879,N_15687);
nor U17539 (N_17539,N_15602,N_14785);
nand U17540 (N_17540,N_15878,N_14359);
nor U17541 (N_17541,N_14745,N_15523);
or U17542 (N_17542,N_14429,N_14505);
and U17543 (N_17543,N_14713,N_14355);
nand U17544 (N_17544,N_15000,N_15279);
nor U17545 (N_17545,N_15479,N_15876);
xor U17546 (N_17546,N_14855,N_14579);
xnor U17547 (N_17547,N_14129,N_15534);
or U17548 (N_17548,N_14694,N_14924);
nor U17549 (N_17549,N_15302,N_15672);
nand U17550 (N_17550,N_14226,N_14225);
nor U17551 (N_17551,N_15426,N_15266);
nor U17552 (N_17552,N_15765,N_14739);
nor U17553 (N_17553,N_14366,N_14786);
xnor U17554 (N_17554,N_14782,N_15519);
nor U17555 (N_17555,N_15875,N_15407);
nand U17556 (N_17556,N_15141,N_15207);
xnor U17557 (N_17557,N_14959,N_15462);
or U17558 (N_17558,N_14702,N_15185);
nand U17559 (N_17559,N_15040,N_15370);
xor U17560 (N_17560,N_14020,N_14851);
nor U17561 (N_17561,N_14197,N_15107);
nor U17562 (N_17562,N_14514,N_14433);
or U17563 (N_17563,N_14000,N_15302);
xor U17564 (N_17564,N_15095,N_14944);
nand U17565 (N_17565,N_15645,N_14892);
xnor U17566 (N_17566,N_14951,N_15940);
nor U17567 (N_17567,N_15724,N_15488);
nand U17568 (N_17568,N_14666,N_14576);
nand U17569 (N_17569,N_15245,N_15534);
or U17570 (N_17570,N_15472,N_14968);
nor U17571 (N_17571,N_15289,N_14548);
and U17572 (N_17572,N_14079,N_15649);
or U17573 (N_17573,N_14055,N_15313);
or U17574 (N_17574,N_15265,N_14557);
and U17575 (N_17575,N_15024,N_15441);
nand U17576 (N_17576,N_15113,N_15078);
nand U17577 (N_17577,N_15575,N_14384);
nor U17578 (N_17578,N_15176,N_15120);
nor U17579 (N_17579,N_15172,N_15850);
nor U17580 (N_17580,N_15626,N_15121);
and U17581 (N_17581,N_14195,N_15013);
nor U17582 (N_17582,N_15152,N_14124);
nor U17583 (N_17583,N_15124,N_14957);
or U17584 (N_17584,N_15078,N_15214);
xnor U17585 (N_17585,N_14260,N_14690);
xnor U17586 (N_17586,N_15434,N_14098);
and U17587 (N_17587,N_15388,N_15569);
xor U17588 (N_17588,N_14081,N_14603);
nor U17589 (N_17589,N_14186,N_15423);
xor U17590 (N_17590,N_14810,N_14493);
or U17591 (N_17591,N_15737,N_14835);
nand U17592 (N_17592,N_15752,N_15091);
and U17593 (N_17593,N_15511,N_15170);
and U17594 (N_17594,N_14549,N_14552);
xor U17595 (N_17595,N_15939,N_15547);
xnor U17596 (N_17596,N_15786,N_14265);
nor U17597 (N_17597,N_15459,N_14178);
nand U17598 (N_17598,N_14170,N_15690);
and U17599 (N_17599,N_15428,N_14991);
and U17600 (N_17600,N_15960,N_15684);
or U17601 (N_17601,N_14456,N_14615);
or U17602 (N_17602,N_14302,N_15367);
and U17603 (N_17603,N_14527,N_14494);
nand U17604 (N_17604,N_15995,N_14080);
and U17605 (N_17605,N_15079,N_14106);
nor U17606 (N_17606,N_15979,N_15314);
xor U17607 (N_17607,N_14509,N_15829);
nand U17608 (N_17608,N_14399,N_14781);
and U17609 (N_17609,N_15275,N_14779);
nand U17610 (N_17610,N_15875,N_14618);
or U17611 (N_17611,N_14216,N_14639);
nor U17612 (N_17612,N_15038,N_14585);
nand U17613 (N_17613,N_15160,N_15815);
nand U17614 (N_17614,N_15387,N_15174);
nand U17615 (N_17615,N_15863,N_14844);
xor U17616 (N_17616,N_14434,N_15893);
nand U17617 (N_17617,N_14702,N_14797);
xnor U17618 (N_17618,N_15094,N_14724);
nor U17619 (N_17619,N_15812,N_15847);
and U17620 (N_17620,N_15830,N_14877);
nand U17621 (N_17621,N_14934,N_15785);
or U17622 (N_17622,N_15971,N_15405);
xor U17623 (N_17623,N_14935,N_14687);
and U17624 (N_17624,N_14843,N_15618);
xor U17625 (N_17625,N_15787,N_14570);
nor U17626 (N_17626,N_14787,N_14166);
xor U17627 (N_17627,N_14756,N_15956);
nand U17628 (N_17628,N_14834,N_15733);
nor U17629 (N_17629,N_14612,N_15446);
xor U17630 (N_17630,N_14709,N_15952);
xor U17631 (N_17631,N_15811,N_15606);
nor U17632 (N_17632,N_15404,N_14144);
or U17633 (N_17633,N_15700,N_15850);
nor U17634 (N_17634,N_14462,N_15682);
xnor U17635 (N_17635,N_15433,N_15735);
nand U17636 (N_17636,N_15391,N_15843);
or U17637 (N_17637,N_14413,N_14930);
and U17638 (N_17638,N_14219,N_15944);
nand U17639 (N_17639,N_14489,N_14748);
and U17640 (N_17640,N_14542,N_14768);
nor U17641 (N_17641,N_15997,N_14612);
xnor U17642 (N_17642,N_15803,N_15887);
nor U17643 (N_17643,N_14166,N_15015);
nor U17644 (N_17644,N_14214,N_14697);
or U17645 (N_17645,N_14611,N_14297);
or U17646 (N_17646,N_15234,N_15047);
nand U17647 (N_17647,N_15457,N_14239);
and U17648 (N_17648,N_14372,N_14818);
xnor U17649 (N_17649,N_14786,N_14967);
xor U17650 (N_17650,N_14215,N_15628);
or U17651 (N_17651,N_15330,N_14012);
xor U17652 (N_17652,N_15938,N_14834);
nand U17653 (N_17653,N_14518,N_14883);
nor U17654 (N_17654,N_15675,N_14462);
and U17655 (N_17655,N_14753,N_15748);
xor U17656 (N_17656,N_15278,N_14151);
nor U17657 (N_17657,N_14934,N_15259);
nand U17658 (N_17658,N_14447,N_15192);
and U17659 (N_17659,N_15400,N_15600);
nand U17660 (N_17660,N_14142,N_14442);
and U17661 (N_17661,N_15218,N_14245);
nand U17662 (N_17662,N_15423,N_15920);
and U17663 (N_17663,N_15204,N_15657);
or U17664 (N_17664,N_14950,N_15752);
xnor U17665 (N_17665,N_15927,N_14201);
xnor U17666 (N_17666,N_14884,N_14024);
xor U17667 (N_17667,N_14205,N_15533);
or U17668 (N_17668,N_15937,N_14722);
and U17669 (N_17669,N_15812,N_15025);
or U17670 (N_17670,N_14274,N_14226);
nor U17671 (N_17671,N_14275,N_14571);
and U17672 (N_17672,N_14460,N_15590);
xor U17673 (N_17673,N_14448,N_15293);
or U17674 (N_17674,N_15566,N_15663);
nor U17675 (N_17675,N_14137,N_14945);
or U17676 (N_17676,N_15426,N_14828);
xor U17677 (N_17677,N_14190,N_15788);
xor U17678 (N_17678,N_14532,N_14671);
and U17679 (N_17679,N_15416,N_14564);
and U17680 (N_17680,N_15369,N_14134);
nor U17681 (N_17681,N_15018,N_15979);
nand U17682 (N_17682,N_15460,N_15579);
and U17683 (N_17683,N_14909,N_15200);
nor U17684 (N_17684,N_14870,N_14789);
nand U17685 (N_17685,N_15968,N_14464);
nand U17686 (N_17686,N_14508,N_14913);
and U17687 (N_17687,N_14715,N_15093);
xor U17688 (N_17688,N_14723,N_15959);
and U17689 (N_17689,N_14810,N_14086);
or U17690 (N_17690,N_15229,N_15644);
xnor U17691 (N_17691,N_14243,N_15603);
xor U17692 (N_17692,N_14516,N_15526);
xnor U17693 (N_17693,N_14050,N_14692);
nor U17694 (N_17694,N_14119,N_14809);
xnor U17695 (N_17695,N_14982,N_14018);
xor U17696 (N_17696,N_15664,N_14415);
nor U17697 (N_17697,N_14154,N_14433);
xnor U17698 (N_17698,N_15989,N_15306);
nand U17699 (N_17699,N_14219,N_15094);
or U17700 (N_17700,N_15796,N_14448);
or U17701 (N_17701,N_15200,N_15504);
and U17702 (N_17702,N_15390,N_14654);
and U17703 (N_17703,N_14598,N_14025);
xnor U17704 (N_17704,N_15973,N_14649);
and U17705 (N_17705,N_15089,N_15952);
nor U17706 (N_17706,N_15028,N_15319);
and U17707 (N_17707,N_15187,N_14674);
nor U17708 (N_17708,N_14936,N_14942);
or U17709 (N_17709,N_14553,N_15090);
nor U17710 (N_17710,N_15339,N_14686);
xor U17711 (N_17711,N_15837,N_14960);
or U17712 (N_17712,N_15873,N_14239);
xor U17713 (N_17713,N_15292,N_15100);
xnor U17714 (N_17714,N_15392,N_15792);
xnor U17715 (N_17715,N_15879,N_15634);
and U17716 (N_17716,N_15881,N_15039);
and U17717 (N_17717,N_15403,N_15136);
xor U17718 (N_17718,N_15725,N_15633);
nand U17719 (N_17719,N_15526,N_15033);
or U17720 (N_17720,N_14599,N_15749);
nand U17721 (N_17721,N_15070,N_14900);
and U17722 (N_17722,N_14947,N_14362);
xor U17723 (N_17723,N_14527,N_14658);
and U17724 (N_17724,N_14321,N_15141);
nor U17725 (N_17725,N_15588,N_14315);
and U17726 (N_17726,N_14707,N_14037);
and U17727 (N_17727,N_14087,N_14518);
or U17728 (N_17728,N_15083,N_14888);
xnor U17729 (N_17729,N_15950,N_15990);
and U17730 (N_17730,N_14756,N_14814);
xor U17731 (N_17731,N_15593,N_15153);
xnor U17732 (N_17732,N_15821,N_14747);
xor U17733 (N_17733,N_14869,N_14650);
nor U17734 (N_17734,N_14045,N_14211);
and U17735 (N_17735,N_14821,N_15440);
nor U17736 (N_17736,N_14303,N_15520);
xnor U17737 (N_17737,N_14116,N_15937);
nand U17738 (N_17738,N_14429,N_15442);
nand U17739 (N_17739,N_15731,N_14534);
nand U17740 (N_17740,N_14902,N_14018);
xor U17741 (N_17741,N_14545,N_15457);
xnor U17742 (N_17742,N_14100,N_14816);
and U17743 (N_17743,N_14096,N_15074);
nand U17744 (N_17744,N_14643,N_15852);
and U17745 (N_17745,N_14184,N_15037);
xor U17746 (N_17746,N_15865,N_15458);
nor U17747 (N_17747,N_14443,N_14405);
nand U17748 (N_17748,N_14657,N_14471);
nand U17749 (N_17749,N_14620,N_14141);
or U17750 (N_17750,N_15610,N_15250);
and U17751 (N_17751,N_15323,N_15086);
or U17752 (N_17752,N_14354,N_15360);
nor U17753 (N_17753,N_15316,N_15577);
nor U17754 (N_17754,N_15538,N_14123);
or U17755 (N_17755,N_14593,N_14662);
nor U17756 (N_17756,N_15960,N_15186);
nand U17757 (N_17757,N_15771,N_14737);
or U17758 (N_17758,N_15418,N_15421);
xor U17759 (N_17759,N_15388,N_15108);
or U17760 (N_17760,N_15594,N_15589);
or U17761 (N_17761,N_15063,N_15119);
nand U17762 (N_17762,N_15284,N_15753);
or U17763 (N_17763,N_14351,N_15581);
nand U17764 (N_17764,N_15574,N_15228);
xor U17765 (N_17765,N_14226,N_14562);
or U17766 (N_17766,N_15036,N_14084);
or U17767 (N_17767,N_15370,N_14545);
and U17768 (N_17768,N_15389,N_14822);
xnor U17769 (N_17769,N_15760,N_15042);
nor U17770 (N_17770,N_15800,N_15346);
or U17771 (N_17771,N_14755,N_14846);
nor U17772 (N_17772,N_15755,N_14256);
or U17773 (N_17773,N_15211,N_14146);
nand U17774 (N_17774,N_15049,N_15615);
and U17775 (N_17775,N_14841,N_14621);
or U17776 (N_17776,N_15120,N_14099);
nor U17777 (N_17777,N_14135,N_14903);
nand U17778 (N_17778,N_15269,N_15129);
nor U17779 (N_17779,N_15871,N_14683);
and U17780 (N_17780,N_14059,N_14248);
xnor U17781 (N_17781,N_14164,N_15997);
xor U17782 (N_17782,N_14033,N_14553);
and U17783 (N_17783,N_14245,N_14603);
or U17784 (N_17784,N_14567,N_15033);
nand U17785 (N_17785,N_15419,N_15873);
xor U17786 (N_17786,N_15084,N_14891);
xnor U17787 (N_17787,N_15975,N_14613);
or U17788 (N_17788,N_15867,N_14506);
or U17789 (N_17789,N_15277,N_14299);
xor U17790 (N_17790,N_15388,N_15622);
xor U17791 (N_17791,N_15083,N_14806);
nor U17792 (N_17792,N_15128,N_15398);
and U17793 (N_17793,N_15857,N_15147);
or U17794 (N_17794,N_15072,N_15346);
and U17795 (N_17795,N_14741,N_15448);
nand U17796 (N_17796,N_15671,N_15211);
and U17797 (N_17797,N_15910,N_15314);
and U17798 (N_17798,N_15678,N_14367);
or U17799 (N_17799,N_15103,N_15286);
nand U17800 (N_17800,N_14448,N_14664);
and U17801 (N_17801,N_15477,N_14202);
nand U17802 (N_17802,N_15507,N_15653);
nand U17803 (N_17803,N_14066,N_14674);
xor U17804 (N_17804,N_14247,N_14078);
xor U17805 (N_17805,N_14280,N_14454);
or U17806 (N_17806,N_15055,N_14320);
xor U17807 (N_17807,N_15003,N_14359);
nor U17808 (N_17808,N_15574,N_15783);
nand U17809 (N_17809,N_15460,N_14684);
nor U17810 (N_17810,N_14616,N_15443);
nand U17811 (N_17811,N_15175,N_15376);
and U17812 (N_17812,N_15518,N_15026);
and U17813 (N_17813,N_15116,N_14214);
nand U17814 (N_17814,N_15649,N_14896);
nand U17815 (N_17815,N_14844,N_15782);
nor U17816 (N_17816,N_15627,N_15472);
and U17817 (N_17817,N_15646,N_15324);
nand U17818 (N_17818,N_14628,N_14551);
nor U17819 (N_17819,N_15584,N_14669);
or U17820 (N_17820,N_15983,N_15546);
or U17821 (N_17821,N_15143,N_14183);
or U17822 (N_17822,N_15407,N_14384);
nand U17823 (N_17823,N_15531,N_15521);
nor U17824 (N_17824,N_14940,N_15248);
xnor U17825 (N_17825,N_14964,N_15544);
or U17826 (N_17826,N_14639,N_15416);
and U17827 (N_17827,N_15223,N_14075);
xor U17828 (N_17828,N_15068,N_14078);
or U17829 (N_17829,N_14102,N_15100);
or U17830 (N_17830,N_15607,N_15111);
or U17831 (N_17831,N_15619,N_14362);
nor U17832 (N_17832,N_14902,N_15813);
nand U17833 (N_17833,N_14926,N_15435);
nor U17834 (N_17834,N_14274,N_15479);
nor U17835 (N_17835,N_14078,N_15165);
nand U17836 (N_17836,N_15669,N_15801);
nor U17837 (N_17837,N_14593,N_14079);
or U17838 (N_17838,N_15646,N_14890);
and U17839 (N_17839,N_15275,N_14802);
and U17840 (N_17840,N_14445,N_15247);
nand U17841 (N_17841,N_14787,N_14231);
and U17842 (N_17842,N_14007,N_14089);
nor U17843 (N_17843,N_14969,N_15663);
nor U17844 (N_17844,N_14925,N_15863);
nand U17845 (N_17845,N_14082,N_14741);
and U17846 (N_17846,N_15834,N_14232);
nor U17847 (N_17847,N_15972,N_15279);
nor U17848 (N_17848,N_14928,N_15914);
or U17849 (N_17849,N_15108,N_15236);
xnor U17850 (N_17850,N_14922,N_15298);
xor U17851 (N_17851,N_15098,N_14779);
nor U17852 (N_17852,N_15495,N_15107);
xnor U17853 (N_17853,N_14683,N_15137);
and U17854 (N_17854,N_14590,N_14564);
or U17855 (N_17855,N_14955,N_14233);
xor U17856 (N_17856,N_15361,N_15422);
and U17857 (N_17857,N_15334,N_15412);
nor U17858 (N_17858,N_15688,N_15525);
nand U17859 (N_17859,N_15306,N_14773);
xnor U17860 (N_17860,N_15160,N_14724);
nor U17861 (N_17861,N_15865,N_15482);
or U17862 (N_17862,N_15281,N_14095);
and U17863 (N_17863,N_15866,N_14803);
nand U17864 (N_17864,N_14366,N_14257);
or U17865 (N_17865,N_15140,N_15643);
nand U17866 (N_17866,N_15909,N_14578);
and U17867 (N_17867,N_15898,N_14343);
nand U17868 (N_17868,N_15871,N_14427);
or U17869 (N_17869,N_14139,N_14765);
and U17870 (N_17870,N_14408,N_14960);
nor U17871 (N_17871,N_15743,N_14448);
nor U17872 (N_17872,N_15119,N_15380);
xor U17873 (N_17873,N_14844,N_15413);
xor U17874 (N_17874,N_14316,N_14718);
nand U17875 (N_17875,N_15970,N_15367);
and U17876 (N_17876,N_14629,N_14676);
or U17877 (N_17877,N_14086,N_15761);
or U17878 (N_17878,N_14857,N_14310);
and U17879 (N_17879,N_15860,N_14060);
xor U17880 (N_17880,N_14361,N_15172);
nand U17881 (N_17881,N_14269,N_14047);
xnor U17882 (N_17882,N_14656,N_15545);
and U17883 (N_17883,N_15954,N_15383);
or U17884 (N_17884,N_15756,N_15331);
and U17885 (N_17885,N_15451,N_15549);
and U17886 (N_17886,N_14137,N_15257);
and U17887 (N_17887,N_15350,N_14162);
xnor U17888 (N_17888,N_14551,N_15733);
nor U17889 (N_17889,N_14173,N_15942);
nand U17890 (N_17890,N_14639,N_15967);
xor U17891 (N_17891,N_15012,N_15205);
or U17892 (N_17892,N_15778,N_14197);
nor U17893 (N_17893,N_14985,N_14837);
nor U17894 (N_17894,N_15166,N_14931);
nand U17895 (N_17895,N_15207,N_15710);
nand U17896 (N_17896,N_15813,N_14519);
nor U17897 (N_17897,N_15422,N_14306);
nand U17898 (N_17898,N_15434,N_14209);
xor U17899 (N_17899,N_14497,N_15789);
nor U17900 (N_17900,N_15838,N_14613);
nor U17901 (N_17901,N_15361,N_14345);
nor U17902 (N_17902,N_15782,N_15113);
or U17903 (N_17903,N_14929,N_15470);
or U17904 (N_17904,N_15881,N_15499);
nand U17905 (N_17905,N_14797,N_14598);
xor U17906 (N_17906,N_14155,N_15641);
or U17907 (N_17907,N_15987,N_15364);
xor U17908 (N_17908,N_15299,N_14537);
xor U17909 (N_17909,N_14000,N_15655);
or U17910 (N_17910,N_14788,N_14430);
and U17911 (N_17911,N_15759,N_15312);
nor U17912 (N_17912,N_15533,N_15921);
xor U17913 (N_17913,N_15939,N_15441);
nor U17914 (N_17914,N_15256,N_14988);
nand U17915 (N_17915,N_14808,N_14328);
nor U17916 (N_17916,N_15925,N_15444);
xnor U17917 (N_17917,N_14088,N_15718);
nand U17918 (N_17918,N_15236,N_14344);
nand U17919 (N_17919,N_14459,N_14717);
nor U17920 (N_17920,N_15722,N_14278);
nor U17921 (N_17921,N_15407,N_15301);
and U17922 (N_17922,N_14395,N_15275);
and U17923 (N_17923,N_14836,N_15042);
or U17924 (N_17924,N_14121,N_15132);
nand U17925 (N_17925,N_14478,N_14546);
nand U17926 (N_17926,N_15873,N_15703);
xnor U17927 (N_17927,N_14213,N_15844);
nand U17928 (N_17928,N_15563,N_14781);
nor U17929 (N_17929,N_15795,N_15906);
nand U17930 (N_17930,N_14748,N_15778);
or U17931 (N_17931,N_15767,N_14483);
or U17932 (N_17932,N_14074,N_15198);
and U17933 (N_17933,N_14812,N_15630);
xnor U17934 (N_17934,N_15856,N_15610);
xnor U17935 (N_17935,N_15092,N_14593);
and U17936 (N_17936,N_14013,N_14333);
and U17937 (N_17937,N_15227,N_15487);
nand U17938 (N_17938,N_15897,N_15059);
nand U17939 (N_17939,N_14491,N_15319);
nand U17940 (N_17940,N_14651,N_14363);
and U17941 (N_17941,N_15941,N_15142);
xor U17942 (N_17942,N_15102,N_14339);
nand U17943 (N_17943,N_15940,N_15298);
and U17944 (N_17944,N_15888,N_14797);
and U17945 (N_17945,N_15081,N_15995);
nand U17946 (N_17946,N_15905,N_15709);
and U17947 (N_17947,N_14925,N_14648);
xor U17948 (N_17948,N_15277,N_14718);
or U17949 (N_17949,N_14708,N_14078);
or U17950 (N_17950,N_14694,N_14289);
or U17951 (N_17951,N_15858,N_15736);
nand U17952 (N_17952,N_15440,N_14056);
or U17953 (N_17953,N_14655,N_14401);
or U17954 (N_17954,N_14597,N_14454);
xnor U17955 (N_17955,N_15606,N_15747);
and U17956 (N_17956,N_14798,N_14947);
and U17957 (N_17957,N_15382,N_14604);
or U17958 (N_17958,N_15450,N_15368);
and U17959 (N_17959,N_15004,N_14279);
xor U17960 (N_17960,N_15715,N_14204);
or U17961 (N_17961,N_14203,N_15364);
xnor U17962 (N_17962,N_15967,N_15866);
and U17963 (N_17963,N_14624,N_14839);
nor U17964 (N_17964,N_14466,N_14917);
nor U17965 (N_17965,N_14179,N_15645);
nand U17966 (N_17966,N_15177,N_15787);
xnor U17967 (N_17967,N_14437,N_14680);
and U17968 (N_17968,N_15006,N_14910);
nand U17969 (N_17969,N_15318,N_15432);
nand U17970 (N_17970,N_14166,N_14772);
nor U17971 (N_17971,N_14218,N_15202);
nand U17972 (N_17972,N_15822,N_14546);
or U17973 (N_17973,N_15006,N_15453);
nand U17974 (N_17974,N_14591,N_14650);
xor U17975 (N_17975,N_15088,N_15376);
xnor U17976 (N_17976,N_14194,N_14914);
nand U17977 (N_17977,N_14380,N_14885);
and U17978 (N_17978,N_14442,N_14846);
nand U17979 (N_17979,N_15135,N_15284);
and U17980 (N_17980,N_14436,N_14316);
nand U17981 (N_17981,N_14846,N_15177);
or U17982 (N_17982,N_14265,N_15252);
nand U17983 (N_17983,N_15768,N_14600);
or U17984 (N_17984,N_14088,N_14346);
nor U17985 (N_17985,N_15653,N_15151);
or U17986 (N_17986,N_14569,N_14815);
nand U17987 (N_17987,N_15082,N_14756);
or U17988 (N_17988,N_15808,N_14552);
xnor U17989 (N_17989,N_15840,N_14063);
or U17990 (N_17990,N_15272,N_14138);
nor U17991 (N_17991,N_14781,N_15896);
nand U17992 (N_17992,N_14714,N_15738);
nand U17993 (N_17993,N_14998,N_14876);
xor U17994 (N_17994,N_15055,N_15507);
xnor U17995 (N_17995,N_14687,N_14647);
or U17996 (N_17996,N_14090,N_15532);
nand U17997 (N_17997,N_15183,N_15321);
nand U17998 (N_17998,N_14766,N_15914);
and U17999 (N_17999,N_14062,N_14334);
nand U18000 (N_18000,N_16696,N_16131);
and U18001 (N_18001,N_16975,N_16938);
and U18002 (N_18002,N_17046,N_16235);
xnor U18003 (N_18003,N_16650,N_16399);
nor U18004 (N_18004,N_17169,N_17265);
or U18005 (N_18005,N_16047,N_17054);
and U18006 (N_18006,N_16619,N_17631);
xnor U18007 (N_18007,N_17803,N_17780);
or U18008 (N_18008,N_17412,N_16206);
nand U18009 (N_18009,N_17355,N_16651);
nor U18010 (N_18010,N_17326,N_16655);
nand U18011 (N_18011,N_16200,N_17321);
nor U18012 (N_18012,N_17986,N_16703);
or U18013 (N_18013,N_16970,N_17354);
and U18014 (N_18014,N_16254,N_17301);
or U18015 (N_18015,N_17651,N_17995);
xnor U18016 (N_18016,N_16036,N_16972);
or U18017 (N_18017,N_17347,N_17077);
xnor U18018 (N_18018,N_17550,N_17450);
nand U18019 (N_18019,N_17055,N_17204);
nand U18020 (N_18020,N_17339,N_16075);
xor U18021 (N_18021,N_16923,N_17726);
nand U18022 (N_18022,N_16705,N_16714);
xor U18023 (N_18023,N_17615,N_16884);
and U18024 (N_18024,N_17741,N_16828);
and U18025 (N_18025,N_17661,N_16546);
nand U18026 (N_18026,N_16679,N_17443);
xnor U18027 (N_18027,N_17068,N_16199);
and U18028 (N_18028,N_17989,N_16327);
xnor U18029 (N_18029,N_17244,N_16357);
and U18030 (N_18030,N_16516,N_17334);
or U18031 (N_18031,N_16486,N_16548);
and U18032 (N_18032,N_17649,N_16997);
and U18033 (N_18033,N_17267,N_17132);
nand U18034 (N_18034,N_17013,N_16067);
nor U18035 (N_18035,N_16168,N_17778);
nand U18036 (N_18036,N_16164,N_16937);
and U18037 (N_18037,N_17150,N_16996);
or U18038 (N_18038,N_17319,N_17369);
xnor U18039 (N_18039,N_16373,N_17496);
and U18040 (N_18040,N_16897,N_17987);
nand U18041 (N_18041,N_16847,N_17205);
xor U18042 (N_18042,N_17019,N_17036);
or U18043 (N_18043,N_17922,N_16228);
or U18044 (N_18044,N_17112,N_16919);
or U18045 (N_18045,N_17647,N_17826);
xnor U18046 (N_18046,N_16121,N_16894);
or U18047 (N_18047,N_17634,N_16999);
nor U18048 (N_18048,N_16402,N_16282);
and U18049 (N_18049,N_17910,N_17302);
xnor U18050 (N_18050,N_17609,N_16858);
and U18051 (N_18051,N_16885,N_17892);
xor U18052 (N_18052,N_16429,N_17870);
xor U18053 (N_18053,N_16032,N_16761);
nand U18054 (N_18054,N_16185,N_16571);
xor U18055 (N_18055,N_16754,N_17291);
xnor U18056 (N_18056,N_17537,N_16807);
xor U18057 (N_18057,N_16447,N_16393);
xnor U18058 (N_18058,N_16215,N_16946);
nand U18059 (N_18059,N_16944,N_16818);
xor U18060 (N_18060,N_16415,N_16125);
or U18061 (N_18061,N_16718,N_17970);
and U18062 (N_18062,N_17900,N_16234);
and U18063 (N_18063,N_16717,N_17610);
or U18064 (N_18064,N_16798,N_17600);
and U18065 (N_18065,N_16671,N_16272);
and U18066 (N_18066,N_16311,N_17784);
or U18067 (N_18067,N_17697,N_17236);
or U18068 (N_18068,N_16560,N_16715);
or U18069 (N_18069,N_16343,N_16670);
nor U18070 (N_18070,N_17133,N_17084);
and U18071 (N_18071,N_16502,N_17116);
or U18072 (N_18072,N_16680,N_17191);
nor U18073 (N_18073,N_16621,N_17297);
xor U18074 (N_18074,N_17493,N_16458);
or U18075 (N_18075,N_17795,N_17747);
nand U18076 (N_18076,N_16806,N_16732);
nand U18077 (N_18077,N_17215,N_17078);
or U18078 (N_18078,N_17269,N_16635);
nand U18079 (N_18079,N_17119,N_16893);
nand U18080 (N_18080,N_16735,N_17536);
nand U18081 (N_18081,N_17771,N_16222);
nor U18082 (N_18082,N_16500,N_16252);
xor U18083 (N_18083,N_17225,N_16437);
nor U18084 (N_18084,N_16287,N_16823);
nand U18085 (N_18085,N_17156,N_16154);
nand U18086 (N_18086,N_17488,N_17394);
xor U18087 (N_18087,N_16531,N_16600);
xnor U18088 (N_18088,N_17271,N_16250);
xnor U18089 (N_18089,N_16641,N_17501);
nand U18090 (N_18090,N_16266,N_16766);
xnor U18091 (N_18091,N_17263,N_16904);
and U18092 (N_18092,N_16618,N_17681);
xnor U18093 (N_18093,N_16793,N_17375);
nor U18094 (N_18094,N_17325,N_16450);
or U18095 (N_18095,N_16179,N_16787);
nor U18096 (N_18096,N_17294,N_16935);
nor U18097 (N_18097,N_17272,N_17854);
nor U18098 (N_18098,N_16167,N_16589);
nor U18099 (N_18099,N_16508,N_16095);
nand U18100 (N_18100,N_17690,N_16720);
xnor U18101 (N_18101,N_17274,N_17599);
nor U18102 (N_18102,N_17814,N_17466);
nor U18103 (N_18103,N_16265,N_17528);
xor U18104 (N_18104,N_16666,N_16066);
or U18105 (N_18105,N_17492,N_17833);
xnor U18106 (N_18106,N_17613,N_16941);
xnor U18107 (N_18107,N_16379,N_16640);
nor U18108 (N_18108,N_17903,N_17167);
and U18109 (N_18109,N_17961,N_16190);
or U18110 (N_18110,N_16637,N_17040);
nor U18111 (N_18111,N_17024,N_17101);
xor U18112 (N_18112,N_17473,N_16054);
or U18113 (N_18113,N_16449,N_16607);
and U18114 (N_18114,N_17070,N_16033);
or U18115 (N_18115,N_17658,N_17308);
nor U18116 (N_18116,N_17632,N_17823);
nor U18117 (N_18117,N_17117,N_16009);
nand U18118 (N_18118,N_16340,N_16656);
xor U18119 (N_18119,N_17606,N_17149);
nand U18120 (N_18120,N_17885,N_17650);
nand U18121 (N_18121,N_16202,N_17923);
and U18122 (N_18122,N_17785,N_16826);
or U18123 (N_18123,N_16109,N_16021);
nand U18124 (N_18124,N_16601,N_16479);
nand U18125 (N_18125,N_17999,N_16588);
nand U18126 (N_18126,N_16139,N_17221);
and U18127 (N_18127,N_17305,N_17762);
nand U18128 (N_18128,N_17232,N_17901);
nor U18129 (N_18129,N_16734,N_17282);
or U18130 (N_18130,N_17009,N_16940);
nor U18131 (N_18131,N_17688,N_17505);
nand U18132 (N_18132,N_17226,N_16976);
or U18133 (N_18133,N_16845,N_17500);
xor U18134 (N_18134,N_17283,N_17640);
and U18135 (N_18135,N_17597,N_16183);
nand U18136 (N_18136,N_16647,N_17927);
and U18137 (N_18137,N_17947,N_16196);
or U18138 (N_18138,N_16323,N_16603);
or U18139 (N_18139,N_16662,N_17855);
xnor U18140 (N_18140,N_17593,N_17454);
nand U18141 (N_18141,N_17011,N_17968);
xnor U18142 (N_18142,N_17994,N_16321);
and U18143 (N_18143,N_17779,N_16470);
xor U18144 (N_18144,N_17813,N_17285);
nor U18145 (N_18145,N_17094,N_17745);
nor U18146 (N_18146,N_17086,N_16256);
nand U18147 (N_18147,N_17715,N_16989);
nand U18148 (N_18148,N_16043,N_17468);
xor U18149 (N_18149,N_16553,N_17194);
nor U18150 (N_18150,N_17007,N_17908);
or U18151 (N_18151,N_16281,N_16163);
and U18152 (N_18152,N_17769,N_17476);
or U18153 (N_18153,N_17208,N_16140);
and U18154 (N_18154,N_17003,N_17139);
or U18155 (N_18155,N_16104,N_16969);
or U18156 (N_18156,N_16060,N_16188);
nand U18157 (N_18157,N_17792,N_16003);
xor U18158 (N_18158,N_17256,N_16042);
nor U18159 (N_18159,N_16342,N_17017);
and U18160 (N_18160,N_16055,N_16028);
xnor U18161 (N_18161,N_17012,N_16263);
nand U18162 (N_18162,N_16332,N_17320);
xnor U18163 (N_18163,N_16676,N_17462);
nor U18164 (N_18164,N_16118,N_16752);
xor U18165 (N_18165,N_17393,N_17368);
xor U18166 (N_18166,N_16848,N_16518);
nor U18167 (N_18167,N_17856,N_17577);
xor U18168 (N_18168,N_17783,N_16750);
xnor U18169 (N_18169,N_16690,N_16669);
nand U18170 (N_18170,N_16472,N_17033);
xnor U18171 (N_18171,N_16280,N_16182);
nor U18172 (N_18172,N_17975,N_17273);
nor U18173 (N_18173,N_16368,N_17703);
and U18174 (N_18174,N_17941,N_17158);
nand U18175 (N_18175,N_17936,N_17511);
nor U18176 (N_18176,N_16305,N_16581);
xnor U18177 (N_18177,N_16499,N_16051);
or U18178 (N_18178,N_17674,N_16704);
and U18179 (N_18179,N_16741,N_16172);
nor U18180 (N_18180,N_16000,N_16902);
and U18181 (N_18181,N_16024,N_17620);
nand U18182 (N_18182,N_17031,N_16451);
and U18183 (N_18183,N_16425,N_16934);
nor U18184 (N_18184,N_17211,N_17281);
or U18185 (N_18185,N_17638,N_16008);
or U18186 (N_18186,N_17956,N_16924);
xnor U18187 (N_18187,N_16347,N_16089);
nand U18188 (N_18188,N_17381,N_17136);
xor U18189 (N_18189,N_16722,N_16391);
xnor U18190 (N_18190,N_16420,N_17755);
or U18191 (N_18191,N_16632,N_16294);
nor U18192 (N_18192,N_16503,N_17085);
nor U18193 (N_18193,N_16563,N_17526);
xor U18194 (N_18194,N_17045,N_17948);
xnor U18195 (N_18195,N_16356,N_17881);
nand U18196 (N_18196,N_16638,N_16709);
and U18197 (N_18197,N_16874,N_17406);
nand U18198 (N_18198,N_17092,N_17564);
nor U18199 (N_18199,N_16951,N_17918);
or U18200 (N_18200,N_17126,N_16817);
xor U18201 (N_18201,N_17764,N_16881);
or U18202 (N_18202,N_16537,N_16105);
and U18203 (N_18203,N_17965,N_17341);
xor U18204 (N_18204,N_17382,N_16314);
xnor U18205 (N_18205,N_17372,N_16112);
nor U18206 (N_18206,N_16697,N_17023);
nand U18207 (N_18207,N_17853,N_16865);
nor U18208 (N_18208,N_17617,N_17777);
nand U18209 (N_18209,N_17644,N_17125);
and U18210 (N_18210,N_17818,N_17370);
nand U18211 (N_18211,N_17246,N_16137);
or U18212 (N_18212,N_16731,N_17098);
and U18213 (N_18213,N_17423,N_17641);
and U18214 (N_18214,N_16466,N_17852);
nand U18215 (N_18215,N_16478,N_17736);
or U18216 (N_18216,N_16918,N_17952);
xnor U18217 (N_18217,N_17653,N_17008);
nor U18218 (N_18218,N_16275,N_16617);
and U18219 (N_18219,N_16257,N_17891);
and U18220 (N_18220,N_16273,N_17489);
or U18221 (N_18221,N_16046,N_16952);
and U18222 (N_18222,N_16065,N_17800);
or U18223 (N_18223,N_17485,N_17127);
nor U18224 (N_18224,N_16496,N_16339);
nor U18225 (N_18225,N_16728,N_17477);
xor U18226 (N_18226,N_16044,N_16261);
and U18227 (N_18227,N_16905,N_16076);
nor U18228 (N_18228,N_17432,N_16219);
nor U18229 (N_18229,N_17160,N_16433);
or U18230 (N_18230,N_17974,N_17866);
xnor U18231 (N_18231,N_16031,N_16476);
xnor U18232 (N_18232,N_16296,N_17479);
nand U18233 (N_18233,N_17560,N_16221);
or U18234 (N_18234,N_17626,N_17893);
xnor U18235 (N_18235,N_16099,N_17206);
nor U18236 (N_18236,N_16528,N_17907);
and U18237 (N_18237,N_16783,N_16128);
and U18238 (N_18238,N_16879,N_17574);
or U18239 (N_18239,N_17464,N_16041);
nor U18240 (N_18240,N_16930,N_16156);
and U18241 (N_18241,N_16568,N_16570);
nor U18242 (N_18242,N_17707,N_16485);
or U18243 (N_18243,N_16233,N_17746);
nor U18244 (N_18244,N_17234,N_17237);
and U18245 (N_18245,N_16812,N_16763);
nor U18246 (N_18246,N_16522,N_17310);
and U18247 (N_18247,N_17129,N_17794);
nor U18248 (N_18248,N_17679,N_17992);
nor U18249 (N_18249,N_16428,N_17721);
nand U18250 (N_18250,N_17004,N_16710);
xnor U18251 (N_18251,N_17686,N_17134);
or U18252 (N_18252,N_17482,N_16757);
and U18253 (N_18253,N_17403,N_17587);
nand U18254 (N_18254,N_16802,N_16507);
and U18255 (N_18255,N_16362,N_16557);
nor U18256 (N_18256,N_17904,N_17220);
xor U18257 (N_18257,N_17239,N_16313);
or U18258 (N_18258,N_16114,N_17197);
or U18259 (N_18259,N_17839,N_17719);
xnor U18260 (N_18260,N_16595,N_16844);
and U18261 (N_18261,N_16835,N_17449);
and U18262 (N_18262,N_16630,N_16404);
and U18263 (N_18263,N_17962,N_17201);
xor U18264 (N_18264,N_16910,N_16290);
nand U18265 (N_18265,N_16446,N_17774);
xor U18266 (N_18266,N_16441,N_16226);
xor U18267 (N_18267,N_16903,N_17603);
xnor U18268 (N_18268,N_17034,N_17635);
or U18269 (N_18269,N_17228,N_16867);
nor U18270 (N_18270,N_17152,N_16577);
nand U18271 (N_18271,N_16096,N_17612);
or U18272 (N_18272,N_16611,N_17619);
or U18273 (N_18273,N_17512,N_17434);
and U18274 (N_18274,N_16085,N_17481);
nor U18275 (N_18275,N_16334,N_16539);
and U18276 (N_18276,N_16816,N_17331);
nand U18277 (N_18277,N_16438,N_16130);
or U18278 (N_18278,N_17105,N_16231);
nor U18279 (N_18279,N_16369,N_17396);
nand U18280 (N_18280,N_16771,N_16077);
xnor U18281 (N_18281,N_16376,N_16832);
xor U18282 (N_18282,N_17309,N_16108);
nor U18283 (N_18283,N_16074,N_16346);
and U18284 (N_18284,N_17932,N_17595);
and U18285 (N_18285,N_17937,N_16573);
nand U18286 (N_18286,N_17317,N_16587);
nor U18287 (N_18287,N_17542,N_17486);
xor U18288 (N_18288,N_16338,N_16187);
nand U18289 (N_18289,N_17407,N_17812);
or U18290 (N_18290,N_17032,N_16120);
or U18291 (N_18291,N_17867,N_17959);
or U18292 (N_18292,N_17580,N_17342);
nor U18293 (N_18293,N_16634,N_17804);
and U18294 (N_18294,N_17295,N_17151);
nor U18295 (N_18295,N_16901,N_16691);
and U18296 (N_18296,N_16749,N_17628);
xor U18297 (N_18297,N_17765,N_16431);
nor U18298 (N_18298,N_17541,N_16210);
and U18299 (N_18299,N_17336,N_16963);
nand U18300 (N_18300,N_16310,N_17413);
nor U18301 (N_18301,N_16291,N_16981);
nor U18302 (N_18302,N_16020,N_17664);
nand U18303 (N_18303,N_17060,N_16015);
and U18304 (N_18304,N_16469,N_16141);
and U18305 (N_18305,N_17039,N_17251);
nor U18306 (N_18306,N_16132,N_17914);
nor U18307 (N_18307,N_17422,N_17386);
or U18308 (N_18308,N_17805,N_16492);
or U18309 (N_18309,N_17524,N_17497);
xnor U18310 (N_18310,N_16360,N_17383);
nand U18311 (N_18311,N_17076,N_17109);
nand U18312 (N_18312,N_16877,N_17447);
or U18313 (N_18313,N_17984,N_16053);
nand U18314 (N_18314,N_16318,N_16796);
and U18315 (N_18315,N_17731,N_16861);
nor U18316 (N_18316,N_17038,N_17988);
nor U18317 (N_18317,N_16465,N_17598);
nand U18318 (N_18318,N_17364,N_16336);
xnor U18319 (N_18319,N_17581,N_17346);
xnor U18320 (N_18320,N_17416,N_16383);
nor U18321 (N_18321,N_16724,N_16688);
nor U18322 (N_18322,N_16255,N_16958);
and U18323 (N_18323,N_17583,N_17453);
nor U18324 (N_18324,N_17047,N_16948);
xor U18325 (N_18325,N_16126,N_17171);
and U18326 (N_18326,N_17335,N_16058);
nor U18327 (N_18327,N_16532,N_17071);
nor U18328 (N_18328,N_17035,N_17535);
nor U18329 (N_18329,N_16358,N_16035);
nand U18330 (N_18330,N_16837,N_16295);
nand U18331 (N_18331,N_17672,N_16390);
xor U18332 (N_18332,N_16019,N_16138);
xnor U18333 (N_18333,N_16061,N_17090);
nand U18334 (N_18334,N_17278,N_16913);
nand U18335 (N_18335,N_16361,N_17062);
nor U18336 (N_18336,N_17155,N_17808);
and U18337 (N_18337,N_16983,N_17063);
xor U18338 (N_18338,N_17058,N_16652);
nor U18339 (N_18339,N_17685,N_16682);
and U18340 (N_18340,N_16153,N_16609);
xnor U18341 (N_18341,N_16134,N_17967);
or U18342 (N_18342,N_16925,N_16950);
nor U18343 (N_18343,N_16224,N_16544);
xnor U18344 (N_18344,N_17056,N_16349);
nand U18345 (N_18345,N_17157,N_17519);
xnor U18346 (N_18346,N_16922,N_17380);
nand U18347 (N_18347,N_17825,N_17217);
xor U18348 (N_18348,N_17569,N_16567);
nor U18349 (N_18349,N_17388,N_16216);
nor U18350 (N_18350,N_17875,N_17130);
nand U18351 (N_18351,N_16536,N_17872);
xnor U18352 (N_18352,N_17973,N_16100);
nor U18353 (N_18353,N_16527,N_17521);
xnor U18354 (N_18354,N_17053,N_17052);
nor U18355 (N_18355,N_16283,N_16864);
and U18356 (N_18356,N_16755,N_17292);
and U18357 (N_18357,N_17820,N_17270);
xor U18358 (N_18358,N_16514,N_16953);
nand U18359 (N_18359,N_17576,N_17934);
nor U18360 (N_18360,N_16916,N_16227);
nand U18361 (N_18361,N_16027,N_17358);
xor U18362 (N_18362,N_17378,N_17895);
or U18363 (N_18363,N_16460,N_16162);
xor U18364 (N_18364,N_17314,N_17884);
nand U18365 (N_18365,N_16191,N_16062);
nand U18366 (N_18366,N_16464,N_16145);
or U18367 (N_18367,N_16454,N_17349);
nand U18368 (N_18368,N_16456,N_16685);
and U18369 (N_18369,N_17057,N_16333);
xor U18370 (N_18370,N_16423,N_16700);
and U18371 (N_18371,N_17337,N_16980);
nor U18372 (N_18372,N_17773,N_16194);
and U18373 (N_18373,N_16056,N_16088);
nor U18374 (N_18374,N_16010,N_17452);
and U18375 (N_18375,N_16928,N_16474);
nor U18376 (N_18376,N_16029,N_16914);
or U18377 (N_18377,N_17689,N_17142);
nand U18378 (N_18378,N_17093,N_17680);
xor U18379 (N_18379,N_16253,N_16768);
nor U18380 (N_18380,N_17427,N_17182);
nor U18381 (N_18381,N_17700,N_17328);
and U18382 (N_18382,N_16551,N_17522);
xnor U18383 (N_18383,N_17671,N_16473);
nand U18384 (N_18384,N_16344,N_17607);
and U18385 (N_18385,N_16876,N_16288);
nand U18386 (N_18386,N_16598,N_17520);
nand U18387 (N_18387,N_17103,N_17656);
xor U18388 (N_18388,N_16098,N_17508);
xnor U18389 (N_18389,N_16049,N_17100);
xnor U18390 (N_18390,N_17556,N_16052);
or U18391 (N_18391,N_17426,N_17252);
and U18392 (N_18392,N_16094,N_17742);
or U18393 (N_18393,N_16022,N_16330);
nand U18394 (N_18394,N_16013,N_16986);
or U18395 (N_18395,N_16026,N_17801);
or U18396 (N_18396,N_17280,N_16303);
and U18397 (N_18397,N_16808,N_17192);
or U18398 (N_18398,N_16854,N_16401);
xnor U18399 (N_18399,N_16827,N_17327);
nand U18400 (N_18400,N_17663,N_17706);
or U18401 (N_18401,N_16048,N_16737);
or U18402 (N_18402,N_16960,N_16775);
nand U18403 (N_18403,N_16284,N_16648);
or U18404 (N_18404,N_16912,N_17161);
or U18405 (N_18405,N_16248,N_16564);
xor U18406 (N_18406,N_16180,N_16378);
xnor U18407 (N_18407,N_17200,N_17879);
nor U18408 (N_18408,N_16961,N_17289);
xnor U18409 (N_18409,N_16899,N_17111);
and U18410 (N_18410,N_17919,N_17738);
xnor U18411 (N_18411,N_17623,N_16488);
and U18412 (N_18412,N_16736,N_16444);
or U18413 (N_18413,N_17869,N_17193);
and U18414 (N_18414,N_17163,N_16435);
nor U18415 (N_18415,N_17441,N_17475);
nor U18416 (N_18416,N_16157,N_16487);
nand U18417 (N_18417,N_16471,N_16891);
nand U18418 (N_18418,N_17629,N_16880);
nor U18419 (N_18419,N_16413,N_17873);
nand U18420 (N_18420,N_17323,N_16663);
nand U18421 (N_18421,N_16805,N_17916);
nand U18422 (N_18422,N_16278,N_17250);
xnor U18423 (N_18423,N_16947,N_17123);
and U18424 (N_18424,N_16626,N_17570);
nor U18425 (N_18425,N_16374,N_16405);
and U18426 (N_18426,N_16968,N_17397);
and U18427 (N_18427,N_16307,N_16629);
and U18428 (N_18428,N_16875,N_16364);
nor U18429 (N_18429,N_16590,N_17750);
xor U18430 (N_18430,N_16610,N_16302);
and U18431 (N_18431,N_16448,N_17436);
and U18432 (N_18432,N_16723,N_17859);
xnor U18433 (N_18433,N_17333,N_16151);
nor U18434 (N_18434,N_17425,N_16515);
nor U18435 (N_18435,N_16057,N_17392);
nor U18436 (N_18436,N_16417,N_17042);
xnor U18437 (N_18437,N_17490,N_17389);
or U18438 (N_18438,N_17313,N_16385);
nand U18439 (N_18439,N_16069,N_16707);
or U18440 (N_18440,N_16606,N_17954);
or U18441 (N_18441,N_16101,N_16247);
or U18442 (N_18442,N_17041,N_16301);
and U18443 (N_18443,N_17049,N_17311);
and U18444 (N_18444,N_16037,N_16942);
and U18445 (N_18445,N_17811,N_16160);
nor U18446 (N_18446,N_16025,N_17074);
nand U18447 (N_18447,N_17790,N_16921);
and U18448 (N_18448,N_16834,N_16073);
nor U18449 (N_18449,N_16774,N_16887);
and U18450 (N_18450,N_16803,N_16006);
nand U18451 (N_18451,N_16646,N_16214);
nand U18452 (N_18452,N_17964,N_16561);
nor U18453 (N_18453,N_17248,N_17979);
and U18454 (N_18454,N_16790,N_17467);
xor U18455 (N_18455,N_16445,N_16936);
nor U18456 (N_18456,N_16692,N_16135);
nand U18457 (N_18457,N_16576,N_16838);
or U18458 (N_18458,N_16142,N_16389);
or U18459 (N_18459,N_16543,N_17022);
or U18460 (N_18460,N_16974,N_17050);
nand U18461 (N_18461,N_17245,N_17940);
or U18462 (N_18462,N_17474,N_16122);
nor U18463 (N_18463,N_17082,N_16195);
nor U18464 (N_18464,N_17376,N_17530);
nand U18465 (N_18465,N_17409,N_16945);
or U18466 (N_18466,N_17568,N_17400);
nor U18467 (N_18467,N_17431,N_16239);
nor U18468 (N_18468,N_17601,N_16149);
or U18469 (N_18469,N_17911,N_16767);
nor U18470 (N_18470,N_17165,N_16993);
xor U18471 (N_18471,N_16966,N_16298);
xnor U18472 (N_18472,N_16242,N_16208);
nor U18473 (N_18473,N_16493,N_16007);
nand U18474 (N_18474,N_17072,N_17361);
or U18475 (N_18475,N_16186,N_16730);
nand U18476 (N_18476,N_16729,N_16434);
and U18477 (N_18477,N_16534,N_16501);
or U18478 (N_18478,N_16932,N_16505);
or U18479 (N_18479,N_16395,N_17566);
nand U18480 (N_18480,N_16129,N_16841);
nand U18481 (N_18481,N_17455,N_16773);
nand U18482 (N_18482,N_16240,N_17164);
and U18483 (N_18483,N_17945,N_16566);
and U18484 (N_18484,N_17075,N_17714);
nor U18485 (N_18485,N_16353,N_17770);
xor U18486 (N_18486,N_16494,N_16843);
nand U18487 (N_18487,N_17740,N_17287);
nor U18488 (N_18488,N_16594,N_17749);
and U18489 (N_18489,N_16939,N_16713);
xor U18490 (N_18490,N_16529,N_17976);
and U18491 (N_18491,N_16907,N_16034);
xor U18492 (N_18492,N_17531,N_16331);
and U18493 (N_18493,N_16672,N_17099);
or U18494 (N_18494,N_16579,N_16982);
and U18495 (N_18495,N_17643,N_17448);
nand U18496 (N_18496,N_16269,N_16675);
xor U18497 (N_18497,N_16512,N_17831);
xor U18498 (N_18498,N_16205,N_16929);
nor U18499 (N_18499,N_16427,N_17212);
or U18500 (N_18500,N_16329,N_17258);
or U18501 (N_18501,N_16770,N_16926);
xnor U18502 (N_18502,N_16558,N_17224);
and U18503 (N_18503,N_17909,N_16987);
or U18504 (N_18504,N_16800,N_16315);
nor U18505 (N_18505,N_16397,N_16335);
nor U18506 (N_18506,N_17459,N_16213);
xor U18507 (N_18507,N_16070,N_17588);
and U18508 (N_18508,N_17878,N_16649);
nand U18509 (N_18509,N_17356,N_16764);
nand U18510 (N_18510,N_16517,N_17666);
nand U18511 (N_18511,N_17137,N_16915);
xnor U18512 (N_18512,N_17065,N_16687);
xnor U18513 (N_18513,N_16545,N_17478);
nand U18514 (N_18514,N_16900,N_16799);
xnor U18515 (N_18515,N_17757,N_16538);
nor U18516 (N_18516,N_16127,N_17418);
or U18517 (N_18517,N_16204,N_17010);
nor U18518 (N_18518,N_17398,N_17648);
or U18519 (N_18519,N_16554,N_17828);
or U18520 (N_18520,N_17027,N_16059);
and U18521 (N_18521,N_16259,N_17353);
or U18522 (N_18522,N_17000,N_17307);
nor U18523 (N_18523,N_17614,N_16860);
nor U18524 (N_18524,N_17782,N_17787);
or U18525 (N_18525,N_16398,N_17510);
xnor U18526 (N_18526,N_17079,N_16738);
nor U18527 (N_18527,N_17938,N_17737);
or U18528 (N_18528,N_17145,N_16521);
nor U18529 (N_18529,N_17379,N_17678);
or U18530 (N_18530,N_17391,N_17696);
and U18531 (N_18531,N_17147,N_17028);
nand U18532 (N_18532,N_17238,N_16836);
nand U18533 (N_18533,N_17095,N_17642);
nor U18534 (N_18534,N_17214,N_17266);
and U18535 (N_18535,N_17636,N_16276);
and U18536 (N_18536,N_16481,N_16964);
or U18537 (N_18537,N_16596,N_17827);
xor U18538 (N_18538,N_17405,N_17429);
nor U18539 (N_18539,N_17442,N_17720);
nand U18540 (N_18540,N_16150,N_17516);
and U18541 (N_18541,N_16184,N_16674);
and U18542 (N_18542,N_16147,N_16819);
xor U18543 (N_18543,N_17759,N_16830);
xnor U18544 (N_18544,N_17179,N_16023);
xnor U18545 (N_18545,N_17766,N_17229);
xor U18546 (N_18546,N_16372,N_17360);
nand U18547 (N_18547,N_16985,N_16642);
and U18548 (N_18548,N_16384,N_16480);
nor U18549 (N_18549,N_16462,N_16562);
nor U18550 (N_18550,N_16744,N_17073);
xnor U18551 (N_18551,N_17861,N_17153);
nor U18552 (N_18552,N_16326,N_17920);
and U18553 (N_18553,N_17016,N_17487);
nor U18554 (N_18554,N_16751,N_17835);
or U18555 (N_18555,N_16578,N_16063);
or U18556 (N_18556,N_16811,N_17915);
xnor U18557 (N_18557,N_16984,N_17699);
nor U18558 (N_18558,N_16371,N_16612);
and U18559 (N_18559,N_16176,N_16559);
or U18560 (N_18560,N_16778,N_17676);
nor U18561 (N_18561,N_17154,N_16956);
and U18562 (N_18562,N_17222,N_16068);
nand U18563 (N_18563,N_16461,N_17458);
nand U18564 (N_18564,N_16739,N_17768);
xnor U18565 (N_18565,N_16856,N_17202);
nor U18566 (N_18566,N_16795,N_17340);
or U18567 (N_18567,N_16249,N_17841);
nor U18568 (N_18568,N_17517,N_17437);
nand U18569 (N_18569,N_16238,N_17868);
xor U18570 (N_18570,N_16236,N_16971);
nor U18571 (N_18571,N_16657,N_17563);
or U18572 (N_18572,N_16086,N_17338);
or U18573 (N_18573,N_16244,N_16959);
or U18574 (N_18574,N_17728,N_16178);
nand U18575 (N_18575,N_16394,N_16863);
nor U18576 (N_18576,N_16177,N_17752);
and U18577 (N_18577,N_16477,N_16866);
xor U18578 (N_18578,N_17618,N_17020);
or U18579 (N_18579,N_17926,N_17877);
nor U18580 (N_18580,N_16591,N_16695);
and U18581 (N_18581,N_17815,N_16359);
nor U18582 (N_18582,N_17513,N_16246);
or U18583 (N_18583,N_17332,N_17404);
xor U18584 (N_18584,N_17824,N_16092);
nor U18585 (N_18585,N_16898,N_16794);
or U18586 (N_18586,N_17865,N_17655);
and U18587 (N_18587,N_16117,N_16082);
xnor U18588 (N_18588,N_17083,N_17791);
nor U18589 (N_18589,N_16804,N_16490);
and U18590 (N_18590,N_17509,N_17207);
and U18591 (N_18591,N_17440,N_16616);
or U18592 (N_18592,N_17763,N_16631);
and U18593 (N_18593,N_17633,N_17138);
xor U18594 (N_18594,N_16143,N_17604);
nor U18595 (N_18595,N_17798,N_16004);
xor U18596 (N_18596,N_16223,N_17716);
nand U18597 (N_18597,N_16541,N_16158);
or U18598 (N_18598,N_16605,N_17514);
or U18599 (N_18599,N_17363,N_16345);
and U18600 (N_18600,N_16664,N_16526);
xor U18601 (N_18601,N_17898,N_16583);
xnor U18602 (N_18602,N_17359,N_17141);
nor U18603 (N_18603,N_17743,N_16842);
nand U18604 (N_18604,N_17844,N_17639);
or U18605 (N_18605,N_17748,N_16762);
nand U18606 (N_18606,N_16319,N_17367);
and U18607 (N_18607,N_17351,N_16801);
and U18608 (N_18608,N_17709,N_17924);
nand U18609 (N_18609,N_16643,N_17876);
or U18610 (N_18610,N_17717,N_17438);
or U18611 (N_18611,N_16859,N_17203);
xor U18612 (N_18612,N_17590,N_16556);
nand U18613 (N_18613,N_17415,N_17573);
or U18614 (N_18614,N_16103,N_16524);
and U18615 (N_18615,N_17420,N_16230);
xor U18616 (N_18616,N_17106,N_17495);
xnor U18617 (N_18617,N_17494,N_17387);
or U18618 (N_18618,N_16872,N_16467);
nor U18619 (N_18619,N_17887,N_16719);
nand U18620 (N_18620,N_17122,N_16645);
and U18621 (N_18621,N_16781,N_17761);
xor U18622 (N_18622,N_16426,N_16853);
nor U18623 (N_18623,N_17983,N_16949);
nor U18624 (N_18624,N_17469,N_17849);
nand U18625 (N_18625,N_16742,N_16322);
xnor U18626 (N_18626,N_17776,N_16377);
and U18627 (N_18627,N_16777,N_16155);
xnor U18628 (N_18628,N_17554,N_17611);
nand U18629 (N_18629,N_16355,N_16113);
xnor U18630 (N_18630,N_17539,N_16119);
and U18631 (N_18631,N_17857,N_17502);
nand U18632 (N_18632,N_16366,N_17518);
or U18633 (N_18633,N_17960,N_17842);
nand U18634 (N_18634,N_16878,N_17277);
nor U18635 (N_18635,N_17148,N_16686);
xnor U18636 (N_18636,N_16251,N_17279);
nor U18637 (N_18637,N_17433,N_17064);
xnor U18638 (N_18638,N_16171,N_16038);
nand U18639 (N_18639,N_17515,N_17435);
and U18640 (N_18640,N_16604,N_17963);
nor U18641 (N_18641,N_17061,N_16822);
or U18642 (N_18642,N_17602,N_16584);
or U18643 (N_18643,N_17991,N_16325);
xor U18644 (N_18644,N_17993,N_16908);
nor U18645 (N_18645,N_17286,N_17410);
nand U18646 (N_18646,N_16442,N_17713);
nor U18647 (N_18647,N_16721,N_17659);
nand U18648 (N_18648,N_17411,N_16277);
xor U18649 (N_18649,N_17107,N_16418);
and U18650 (N_18650,N_17753,N_16549);
xor U18651 (N_18651,N_16779,N_16565);
and U18652 (N_18652,N_17616,N_17390);
and U18653 (N_18653,N_16599,N_17365);
xor U18654 (N_18654,N_17847,N_17044);
xnor U18655 (N_18655,N_17586,N_16484);
nand U18656 (N_18656,N_17181,N_16258);
and U18657 (N_18657,N_17725,N_17128);
xor U18658 (N_18658,N_17732,N_16825);
and U18659 (N_18659,N_17548,N_17980);
nor U18660 (N_18660,N_17385,N_17977);
and U18661 (N_18661,N_17860,N_16659);
and U18662 (N_18662,N_17195,N_17544);
or U18663 (N_18663,N_16833,N_16896);
or U18664 (N_18664,N_17622,N_16840);
and U18665 (N_18665,N_16745,N_17786);
xnor U18666 (N_18666,N_16772,N_17582);
or U18667 (N_18667,N_16110,N_17662);
and U18668 (N_18668,N_17553,N_17694);
and U18669 (N_18669,N_16593,N_16030);
or U18670 (N_18670,N_16574,N_17471);
nor U18671 (N_18671,N_16297,N_16513);
xor U18672 (N_18672,N_17727,N_17730);
nand U18673 (N_18673,N_16765,N_16855);
xnor U18674 (N_18674,N_17978,N_16979);
xor U18675 (N_18675,N_16388,N_17704);
nand U18676 (N_18676,N_17373,N_17646);
or U18677 (N_18677,N_17931,N_17444);
nor U18678 (N_18678,N_16888,N_17990);
and U18679 (N_18679,N_17293,N_16625);
and U18680 (N_18680,N_16821,N_17559);
or U18681 (N_18681,N_17087,N_16743);
xor U18682 (N_18682,N_16270,N_17624);
and U18683 (N_18683,N_17470,N_16653);
nor U18684 (N_18684,N_17871,N_16852);
nand U18685 (N_18685,N_16712,N_16575);
nor U18686 (N_18686,N_16181,N_17682);
nor U18687 (N_18687,N_17858,N_16994);
nand U18688 (N_18688,N_17175,N_16170);
or U18689 (N_18689,N_16483,N_16873);
or U18690 (N_18690,N_16608,N_17037);
and U18691 (N_18691,N_17178,N_16279);
or U18692 (N_18692,N_16525,N_17874);
and U18693 (N_18693,N_17846,N_17081);
and U18694 (N_18694,N_16192,N_16520);
xor U18695 (N_18695,N_17143,N_16628);
xnor U18696 (N_18696,N_16491,N_16146);
xor U18697 (N_18697,N_16102,N_16620);
nor U18698 (N_18698,N_17110,N_17230);
and U18699 (N_18699,N_16133,N_16727);
and U18700 (N_18700,N_16463,N_17675);
xnor U18701 (N_18701,N_16400,N_17080);
nand U18702 (N_18702,N_17558,N_17144);
xnor U18703 (N_18703,N_17660,N_17575);
and U18704 (N_18704,N_17097,N_17480);
nor U18705 (N_18705,N_16211,N_17735);
xnor U18706 (N_18706,N_16232,N_16582);
or U18707 (N_18707,N_16497,N_16716);
and U18708 (N_18708,N_16407,N_17943);
and U18709 (N_18709,N_16124,N_16857);
xnor U18710 (N_18710,N_17925,N_16016);
nor U18711 (N_18711,N_17834,N_17837);
nand U18712 (N_18712,N_16998,N_17929);
or U18713 (N_18713,N_16965,N_17950);
nor U18714 (N_18714,N_16410,N_16482);
nor U18715 (N_18715,N_17669,N_17702);
and U18716 (N_18716,N_17249,N_17957);
and U18717 (N_18717,N_17316,N_17185);
nand U18718 (N_18718,N_16011,N_17210);
nand U18719 (N_18719,N_16375,N_17504);
xor U18720 (N_18720,N_16991,N_16111);
nor U18721 (N_18721,N_16954,N_17775);
or U18722 (N_18722,N_16014,N_16789);
xor U18723 (N_18723,N_17329,N_16530);
nand U18724 (N_18724,N_17951,N_17018);
nor U18725 (N_18725,N_16592,N_16078);
and U18726 (N_18726,N_17625,N_16850);
xnor U18727 (N_18727,N_17668,N_16668);
nand U18728 (N_18728,N_17933,N_16203);
or U18729 (N_18729,N_16436,N_16824);
nand U18730 (N_18730,N_16906,N_17419);
xor U18731 (N_18731,N_16694,N_16312);
xnor U18732 (N_18732,N_17756,N_16889);
nor U18733 (N_18733,N_17417,N_17001);
and U18734 (N_18734,N_16175,N_16453);
or U18735 (N_18735,N_16320,N_16990);
or U18736 (N_18736,N_17118,N_17949);
xor U18737 (N_18737,N_17525,N_17089);
nor U18738 (N_18738,N_16623,N_17348);
or U18739 (N_18739,N_16636,N_16308);
nand U18740 (N_18740,N_16622,N_16106);
nand U18741 (N_18741,N_17722,N_16681);
nand U18742 (N_18742,N_17461,N_17772);
nand U18743 (N_18743,N_16509,N_17114);
xor U18744 (N_18744,N_16173,N_17567);
xor U18745 (N_18745,N_17491,N_17781);
nor U18746 (N_18746,N_17767,N_16784);
and U18747 (N_18747,N_17465,N_16689);
nor U18748 (N_18748,N_17902,N_16408);
nand U18749 (N_18749,N_16012,N_17789);
xnor U18750 (N_18750,N_17029,N_17821);
nand U18751 (N_18751,N_16758,N_16869);
xnor U18752 (N_18752,N_17677,N_16911);
nor U18753 (N_18753,N_16309,N_16148);
xor U18754 (N_18754,N_17330,N_17843);
xor U18755 (N_18755,N_16161,N_16093);
nand U18756 (N_18756,N_17135,N_16699);
nand U18757 (N_18757,N_17188,N_17235);
and U18758 (N_18758,N_16300,N_16274);
xor U18759 (N_18759,N_17711,N_17026);
or U18760 (N_18760,N_17850,N_16489);
or U18761 (N_18761,N_17484,N_16396);
and U18762 (N_18762,N_17255,N_16498);
xnor U18763 (N_18763,N_16430,N_17276);
and U18764 (N_18764,N_17264,N_16039);
and U18765 (N_18765,N_17268,N_17971);
and U18766 (N_18766,N_17572,N_17905);
nand U18767 (N_18767,N_17712,N_17802);
xor U18768 (N_18768,N_16381,N_16665);
nor U18769 (N_18769,N_16849,N_16973);
xnor U18770 (N_18770,N_16776,N_16683);
or U18771 (N_18771,N_16411,N_16851);
nand U18772 (N_18772,N_16677,N_17503);
nor U18773 (N_18773,N_17166,N_17534);
and U18774 (N_18774,N_17845,N_16769);
and U18775 (N_18775,N_16432,N_17921);
nand U18776 (N_18776,N_16005,N_17691);
and U18777 (N_18777,N_16292,N_16040);
and U18778 (N_18778,N_17315,N_17810);
or U18779 (N_18779,N_16123,N_17944);
and U18780 (N_18780,N_16870,N_16271);
or U18781 (N_18781,N_17533,N_17708);
nand U18782 (N_18782,N_16733,N_16189);
and U18783 (N_18783,N_16698,N_17888);
or U18784 (N_18784,N_17043,N_17189);
and U18785 (N_18785,N_16387,N_16661);
nor U18786 (N_18786,N_16920,N_17591);
and U18787 (N_18787,N_17608,N_16909);
nor U18788 (N_18788,N_17673,N_17168);
and U18789 (N_18789,N_16107,N_17162);
or U18790 (N_18790,N_17897,N_17829);
nor U18791 (N_18791,N_16245,N_16569);
xnor U18792 (N_18792,N_16090,N_16422);
or U18793 (N_18793,N_16455,N_17701);
nor U18794 (N_18794,N_16613,N_17399);
and U18795 (N_18795,N_17190,N_17240);
xor U18796 (N_18796,N_16370,N_17247);
or U18797 (N_18797,N_17463,N_17131);
nand U18798 (N_18798,N_16159,N_17733);
xnor U18799 (N_18799,N_16785,N_17692);
or U18800 (N_18800,N_17067,N_16580);
xor U18801 (N_18801,N_17159,N_16091);
xor U18802 (N_18802,N_16002,N_17693);
or U18803 (N_18803,N_16706,N_16813);
xnor U18804 (N_18804,N_16627,N_17840);
nor U18805 (N_18805,N_16083,N_17832);
nor U18806 (N_18806,N_16726,N_16931);
or U18807 (N_18807,N_17241,N_16995);
or U18808 (N_18808,N_17928,N_17350);
nor U18809 (N_18809,N_17483,N_17578);
nand U18810 (N_18810,N_16392,N_16693);
nand U18811 (N_18811,N_17414,N_17366);
nand U18812 (N_18812,N_16443,N_16615);
and U18813 (N_18813,N_17817,N_16382);
nand U18814 (N_18814,N_17562,N_16064);
or U18815 (N_18815,N_16748,N_16585);
xnor U18816 (N_18816,N_16380,N_17705);
nand U18817 (N_18817,N_17529,N_17946);
nor U18818 (N_18818,N_16955,N_17472);
and U18819 (N_18819,N_16136,N_16829);
xnor U18820 (N_18820,N_16352,N_16839);
and U18821 (N_18821,N_16207,N_17687);
or U18822 (N_18822,N_17343,N_17362);
and U18823 (N_18823,N_17571,N_16639);
xnor U18824 (N_18824,N_17304,N_17499);
and U18825 (N_18825,N_17439,N_17894);
or U18826 (N_18826,N_17140,N_16684);
and U18827 (N_18827,N_17890,N_16797);
xor U18828 (N_18828,N_17395,N_17751);
and U18829 (N_18829,N_17300,N_16927);
or U18830 (N_18830,N_16711,N_17066);
nand U18831 (N_18831,N_16962,N_16406);
nand U18832 (N_18832,N_16786,N_16363);
nand U18833 (N_18833,N_17899,N_16050);
nor U18834 (N_18834,N_17421,N_16409);
xnor U18835 (N_18835,N_17030,N_17710);
nand U18836 (N_18836,N_17322,N_16572);
and U18837 (N_18837,N_16440,N_17935);
nand U18838 (N_18838,N_17788,N_17665);
nand U18839 (N_18839,N_17917,N_17985);
nor U18840 (N_18840,N_17630,N_17180);
xor U18841 (N_18841,N_16614,N_17547);
nand U18842 (N_18842,N_17170,N_17549);
xor U18843 (N_18843,N_16535,N_16324);
nor U18844 (N_18844,N_17981,N_17059);
or U18845 (N_18845,N_17953,N_17882);
or U18846 (N_18846,N_17579,N_17374);
xnor U18847 (N_18847,N_17864,N_17262);
xor U18848 (N_18848,N_16678,N_17048);
and U18849 (N_18849,N_17552,N_17257);
and U18850 (N_18850,N_17242,N_16882);
nor U18851 (N_18851,N_17371,N_17428);
nand U18852 (N_18852,N_17445,N_16658);
nand U18853 (N_18853,N_16791,N_16814);
or U18854 (N_18854,N_17966,N_16350);
xor U18855 (N_18855,N_16071,N_17532);
or U18856 (N_18856,N_16633,N_16225);
nand U18857 (N_18857,N_17997,N_16523);
nand U18858 (N_18858,N_16087,N_17108);
nand U18859 (N_18859,N_17124,N_17969);
nor U18860 (N_18860,N_16419,N_16892);
or U18861 (N_18861,N_17146,N_16316);
nor U18862 (N_18862,N_16533,N_16495);
or U18863 (N_18863,N_17557,N_16220);
xor U18864 (N_18864,N_17121,N_17793);
nand U18865 (N_18865,N_16586,N_16299);
and U18866 (N_18866,N_17758,N_17889);
nand U18867 (N_18867,N_16988,N_17718);
xor U18868 (N_18868,N_17654,N_17069);
and U18869 (N_18869,N_17913,N_16317);
and U18870 (N_18870,N_17284,N_17408);
and U18871 (N_18871,N_17972,N_17760);
nor U18872 (N_18872,N_17357,N_17015);
xnor U18873 (N_18873,N_17290,N_17187);
nor U18874 (N_18874,N_17739,N_17734);
nand U18875 (N_18875,N_17657,N_17507);
nand U18876 (N_18876,N_17506,N_17807);
and U18877 (N_18877,N_16831,N_17880);
nor U18878 (N_18878,N_17199,N_17806);
nand U18879 (N_18879,N_16367,N_16237);
nor U18880 (N_18880,N_16304,N_17177);
xnor U18881 (N_18881,N_17809,N_17998);
and U18882 (N_18882,N_16193,N_16209);
nor U18883 (N_18883,N_16890,N_16602);
and U18884 (N_18884,N_16386,N_16416);
and U18885 (N_18885,N_16540,N_17596);
xor U18886 (N_18886,N_16212,N_16511);
nor U18887 (N_18887,N_16289,N_17621);
xor U18888 (N_18888,N_17296,N_16229);
and U18889 (N_18889,N_17223,N_17863);
xor U18890 (N_18890,N_17822,N_17312);
nand U18891 (N_18891,N_16597,N_17695);
or U18892 (N_18892,N_17401,N_17113);
xor U18893 (N_18893,N_17176,N_17172);
nor U18894 (N_18894,N_17561,N_17430);
nand U18895 (N_18895,N_17724,N_17498);
and U18896 (N_18896,N_17698,N_16267);
nand U18897 (N_18897,N_16753,N_16262);
and U18898 (N_18898,N_16201,N_17352);
and U18899 (N_18899,N_17594,N_17088);
or U18900 (N_18900,N_16788,N_16883);
nor U18901 (N_18901,N_16782,N_17830);
or U18902 (N_18902,N_16072,N_16756);
nand U18903 (N_18903,N_17384,N_17799);
nor U18904 (N_18904,N_17585,N_17173);
nand U18905 (N_18905,N_16510,N_16917);
nand U18906 (N_18906,N_17115,N_16475);
nor U18907 (N_18907,N_16943,N_16977);
nor U18908 (N_18908,N_17684,N_17198);
nor U18909 (N_18909,N_17836,N_16165);
nor U18910 (N_18910,N_16759,N_17424);
nand U18911 (N_18911,N_17344,N_16660);
or U18912 (N_18912,N_17538,N_17848);
nand U18913 (N_18913,N_17233,N_17021);
or U18914 (N_18914,N_16268,N_16452);
nand U18915 (N_18915,N_17627,N_17218);
xnor U18916 (N_18916,N_16459,N_17527);
or U18917 (N_18917,N_16354,N_16017);
or U18918 (N_18918,N_17838,N_17014);
and U18919 (N_18919,N_16895,N_17942);
or U18920 (N_18920,N_17796,N_16702);
or U18921 (N_18921,N_17862,N_17670);
nor U18922 (N_18922,N_16846,N_17955);
and U18923 (N_18923,N_16116,N_16439);
xnor U18924 (N_18924,N_17005,N_16701);
xnor U18925 (N_18925,N_17584,N_16644);
and U18926 (N_18926,N_16341,N_17051);
nor U18927 (N_18927,N_16552,N_16080);
xor U18928 (N_18928,N_16351,N_17523);
nand U18929 (N_18929,N_17652,N_17797);
and U18930 (N_18930,N_17592,N_16152);
xnor U18931 (N_18931,N_17605,N_17120);
or U18932 (N_18932,N_17551,N_17259);
and U18933 (N_18933,N_17213,N_16217);
or U18934 (N_18934,N_17216,N_16306);
nor U18935 (N_18935,N_17219,N_17209);
nor U18936 (N_18936,N_17104,N_16933);
xor U18937 (N_18937,N_17645,N_17896);
nand U18938 (N_18938,N_17555,N_17851);
or U18939 (N_18939,N_16624,N_16673);
or U18940 (N_18940,N_16746,N_17451);
and U18941 (N_18941,N_17637,N_17183);
nor U18942 (N_18942,N_17939,N_16654);
xor U18943 (N_18943,N_16115,N_16264);
or U18944 (N_18944,N_16747,N_16957);
nand U18945 (N_18945,N_16550,N_16169);
nor U18946 (N_18946,N_16260,N_16542);
xor U18947 (N_18947,N_17096,N_16218);
or U18948 (N_18948,N_17540,N_16871);
and U18949 (N_18949,N_17227,N_16243);
nand U18950 (N_18950,N_17261,N_17883);
xor U18951 (N_18951,N_17460,N_17303);
nor U18952 (N_18952,N_16414,N_17260);
and U18953 (N_18953,N_16241,N_17184);
xor U18954 (N_18954,N_16547,N_17253);
and U18955 (N_18955,N_16198,N_16967);
nor U18956 (N_18956,N_17819,N_16740);
or U18957 (N_18957,N_16780,N_16457);
nor U18958 (N_18958,N_16293,N_17543);
and U18959 (N_18959,N_16809,N_16820);
or U18960 (N_18960,N_16868,N_16337);
nor U18961 (N_18961,N_17545,N_17243);
and U18962 (N_18962,N_17816,N_17457);
xnor U18963 (N_18963,N_16555,N_17288);
or U18964 (N_18964,N_16197,N_17546);
or U18965 (N_18965,N_17958,N_16079);
nor U18966 (N_18966,N_17996,N_17589);
or U18967 (N_18967,N_16725,N_16403);
nand U18968 (N_18968,N_16708,N_17456);
nor U18969 (N_18969,N_16424,N_16421);
nand U18970 (N_18970,N_16412,N_17565);
nor U18971 (N_18971,N_16166,N_16862);
xnor U18972 (N_18972,N_16097,N_16081);
or U18973 (N_18973,N_16018,N_17306);
or U18974 (N_18974,N_17377,N_17402);
and U18975 (N_18975,N_17231,N_17345);
nor U18976 (N_18976,N_16328,N_16810);
or U18977 (N_18977,N_17744,N_17299);
nor U18978 (N_18978,N_17723,N_17982);
xor U18979 (N_18979,N_17446,N_16504);
or U18980 (N_18980,N_16978,N_17196);
nand U18981 (N_18981,N_17102,N_17318);
and U18982 (N_18982,N_16519,N_16667);
nor U18983 (N_18983,N_16285,N_16144);
nor U18984 (N_18984,N_17254,N_17324);
nand U18985 (N_18985,N_17091,N_17906);
nand U18986 (N_18986,N_16815,N_17275);
nand U18987 (N_18987,N_16506,N_16045);
xnor U18988 (N_18988,N_17886,N_17729);
and U18989 (N_18989,N_16760,N_17186);
xnor U18990 (N_18990,N_16174,N_16886);
or U18991 (N_18991,N_16992,N_17298);
or U18992 (N_18992,N_16286,N_17006);
and U18993 (N_18993,N_16001,N_17667);
nand U18994 (N_18994,N_17683,N_17754);
nor U18995 (N_18995,N_17002,N_16792);
nor U18996 (N_18996,N_17930,N_17912);
xnor U18997 (N_18997,N_17174,N_16348);
xor U18998 (N_18998,N_17025,N_16468);
or U18999 (N_18999,N_16365,N_16084);
or U19000 (N_19000,N_17362,N_16644);
nor U19001 (N_19001,N_17689,N_17638);
nand U19002 (N_19002,N_16018,N_17334);
and U19003 (N_19003,N_16021,N_16306);
nand U19004 (N_19004,N_16541,N_16338);
nand U19005 (N_19005,N_16602,N_17027);
nand U19006 (N_19006,N_17543,N_17823);
xnor U19007 (N_19007,N_17208,N_17835);
xor U19008 (N_19008,N_17156,N_16975);
nand U19009 (N_19009,N_17940,N_16067);
and U19010 (N_19010,N_16686,N_17885);
and U19011 (N_19011,N_17459,N_16170);
nor U19012 (N_19012,N_16170,N_17953);
and U19013 (N_19013,N_16752,N_16663);
or U19014 (N_19014,N_16062,N_17904);
nand U19015 (N_19015,N_16621,N_17348);
nor U19016 (N_19016,N_16731,N_17777);
nor U19017 (N_19017,N_17974,N_16376);
xnor U19018 (N_19018,N_16127,N_16680);
and U19019 (N_19019,N_16906,N_16272);
nand U19020 (N_19020,N_17392,N_16721);
and U19021 (N_19021,N_17627,N_17259);
nor U19022 (N_19022,N_17612,N_16651);
nand U19023 (N_19023,N_16932,N_16824);
nor U19024 (N_19024,N_16438,N_17440);
or U19025 (N_19025,N_17012,N_16898);
nand U19026 (N_19026,N_16265,N_16156);
or U19027 (N_19027,N_16802,N_16488);
and U19028 (N_19028,N_16967,N_17631);
xnor U19029 (N_19029,N_16319,N_17700);
nand U19030 (N_19030,N_16744,N_17274);
xor U19031 (N_19031,N_16897,N_16089);
and U19032 (N_19032,N_16625,N_17118);
or U19033 (N_19033,N_16088,N_16842);
nand U19034 (N_19034,N_17113,N_16329);
or U19035 (N_19035,N_16450,N_17502);
nand U19036 (N_19036,N_17316,N_17806);
and U19037 (N_19037,N_17182,N_17050);
nor U19038 (N_19038,N_17089,N_17671);
xor U19039 (N_19039,N_16414,N_16193);
xor U19040 (N_19040,N_16070,N_16784);
and U19041 (N_19041,N_16422,N_16209);
and U19042 (N_19042,N_17998,N_17060);
and U19043 (N_19043,N_17792,N_16451);
nor U19044 (N_19044,N_16034,N_16047);
nand U19045 (N_19045,N_16595,N_17116);
and U19046 (N_19046,N_16223,N_16432);
nand U19047 (N_19047,N_17640,N_17065);
nand U19048 (N_19048,N_17021,N_17762);
nand U19049 (N_19049,N_17558,N_16881);
xor U19050 (N_19050,N_17241,N_17290);
and U19051 (N_19051,N_17703,N_16120);
and U19052 (N_19052,N_17569,N_17807);
xor U19053 (N_19053,N_16399,N_16966);
xor U19054 (N_19054,N_17160,N_16243);
or U19055 (N_19055,N_17889,N_17715);
nand U19056 (N_19056,N_16524,N_16955);
or U19057 (N_19057,N_17648,N_17213);
or U19058 (N_19058,N_16786,N_16795);
and U19059 (N_19059,N_17048,N_17958);
nor U19060 (N_19060,N_16325,N_17391);
nor U19061 (N_19061,N_16637,N_17437);
and U19062 (N_19062,N_17372,N_16356);
nand U19063 (N_19063,N_17691,N_17398);
and U19064 (N_19064,N_17998,N_16934);
nand U19065 (N_19065,N_16301,N_16163);
nand U19066 (N_19066,N_17115,N_16776);
and U19067 (N_19067,N_17721,N_17417);
or U19068 (N_19068,N_16114,N_16677);
nor U19069 (N_19069,N_16117,N_16777);
nor U19070 (N_19070,N_17714,N_16820);
nand U19071 (N_19071,N_16807,N_16766);
xor U19072 (N_19072,N_17572,N_16116);
and U19073 (N_19073,N_17991,N_17748);
xnor U19074 (N_19074,N_16264,N_16005);
or U19075 (N_19075,N_16218,N_16793);
nor U19076 (N_19076,N_16303,N_17569);
nor U19077 (N_19077,N_16884,N_16278);
xnor U19078 (N_19078,N_16448,N_16800);
and U19079 (N_19079,N_17454,N_17549);
xnor U19080 (N_19080,N_16529,N_16482);
or U19081 (N_19081,N_17418,N_17851);
xnor U19082 (N_19082,N_16655,N_17798);
xor U19083 (N_19083,N_17843,N_17636);
nor U19084 (N_19084,N_17522,N_17149);
xor U19085 (N_19085,N_16319,N_16154);
and U19086 (N_19086,N_17341,N_16076);
and U19087 (N_19087,N_17458,N_17469);
or U19088 (N_19088,N_17127,N_17826);
nor U19089 (N_19089,N_17177,N_16823);
nand U19090 (N_19090,N_16601,N_16152);
and U19091 (N_19091,N_17165,N_17791);
and U19092 (N_19092,N_17201,N_17849);
or U19093 (N_19093,N_17445,N_16158);
and U19094 (N_19094,N_17583,N_16772);
or U19095 (N_19095,N_17183,N_17895);
and U19096 (N_19096,N_17140,N_16966);
or U19097 (N_19097,N_17616,N_16166);
or U19098 (N_19098,N_17368,N_17251);
or U19099 (N_19099,N_16324,N_17713);
or U19100 (N_19100,N_17471,N_16325);
xnor U19101 (N_19101,N_17000,N_17512);
nor U19102 (N_19102,N_17695,N_17078);
and U19103 (N_19103,N_16044,N_17571);
nor U19104 (N_19104,N_16826,N_17314);
and U19105 (N_19105,N_16573,N_17176);
nor U19106 (N_19106,N_17208,N_17621);
and U19107 (N_19107,N_17147,N_17696);
or U19108 (N_19108,N_17798,N_17641);
nand U19109 (N_19109,N_16730,N_17135);
and U19110 (N_19110,N_17221,N_16658);
nor U19111 (N_19111,N_17601,N_16480);
xnor U19112 (N_19112,N_17852,N_16497);
nand U19113 (N_19113,N_17811,N_16095);
or U19114 (N_19114,N_16656,N_17153);
and U19115 (N_19115,N_17298,N_16262);
nor U19116 (N_19116,N_17321,N_16017);
xor U19117 (N_19117,N_17490,N_17465);
or U19118 (N_19118,N_17075,N_17550);
or U19119 (N_19119,N_17299,N_16267);
xor U19120 (N_19120,N_16439,N_17388);
nand U19121 (N_19121,N_16785,N_17407);
nand U19122 (N_19122,N_17589,N_17076);
xnor U19123 (N_19123,N_17048,N_16543);
xnor U19124 (N_19124,N_16579,N_16741);
or U19125 (N_19125,N_16235,N_16595);
and U19126 (N_19126,N_17345,N_17116);
nor U19127 (N_19127,N_16933,N_17419);
nor U19128 (N_19128,N_17760,N_17711);
nor U19129 (N_19129,N_16094,N_17390);
nand U19130 (N_19130,N_17781,N_16219);
nand U19131 (N_19131,N_17685,N_17758);
and U19132 (N_19132,N_16225,N_16648);
and U19133 (N_19133,N_16115,N_17722);
and U19134 (N_19134,N_17277,N_16786);
nor U19135 (N_19135,N_16336,N_16181);
and U19136 (N_19136,N_16123,N_16640);
nor U19137 (N_19137,N_16003,N_16745);
nand U19138 (N_19138,N_17904,N_16584);
nor U19139 (N_19139,N_16405,N_16252);
nor U19140 (N_19140,N_16172,N_17432);
and U19141 (N_19141,N_17743,N_17455);
nor U19142 (N_19142,N_17362,N_16863);
or U19143 (N_19143,N_16323,N_17030);
or U19144 (N_19144,N_17994,N_16435);
nand U19145 (N_19145,N_17139,N_17022);
and U19146 (N_19146,N_16784,N_16648);
or U19147 (N_19147,N_16480,N_16831);
xnor U19148 (N_19148,N_16132,N_17302);
or U19149 (N_19149,N_16883,N_16930);
or U19150 (N_19150,N_16112,N_17609);
xor U19151 (N_19151,N_16563,N_16129);
and U19152 (N_19152,N_16624,N_17549);
nand U19153 (N_19153,N_17758,N_16496);
xor U19154 (N_19154,N_16665,N_17593);
nor U19155 (N_19155,N_16304,N_16284);
xnor U19156 (N_19156,N_17775,N_16879);
xor U19157 (N_19157,N_16412,N_17634);
or U19158 (N_19158,N_17797,N_17046);
or U19159 (N_19159,N_17255,N_17870);
nand U19160 (N_19160,N_17087,N_17579);
xor U19161 (N_19161,N_16787,N_16098);
nor U19162 (N_19162,N_17457,N_16659);
nor U19163 (N_19163,N_16174,N_17336);
and U19164 (N_19164,N_17953,N_16768);
and U19165 (N_19165,N_16986,N_16425);
xor U19166 (N_19166,N_16177,N_16822);
xor U19167 (N_19167,N_16119,N_17294);
or U19168 (N_19168,N_16343,N_16562);
or U19169 (N_19169,N_16070,N_17264);
and U19170 (N_19170,N_17281,N_17223);
nand U19171 (N_19171,N_17780,N_17945);
nor U19172 (N_19172,N_16369,N_16757);
nand U19173 (N_19173,N_17975,N_16018);
nand U19174 (N_19174,N_17585,N_17714);
xor U19175 (N_19175,N_17321,N_16778);
and U19176 (N_19176,N_16642,N_16532);
nand U19177 (N_19177,N_17190,N_16824);
xor U19178 (N_19178,N_17095,N_17304);
and U19179 (N_19179,N_17364,N_16307);
and U19180 (N_19180,N_17410,N_17762);
nand U19181 (N_19181,N_16732,N_17533);
xor U19182 (N_19182,N_16351,N_16812);
and U19183 (N_19183,N_17742,N_17457);
nor U19184 (N_19184,N_16340,N_17462);
or U19185 (N_19185,N_17883,N_16521);
xor U19186 (N_19186,N_17125,N_17273);
and U19187 (N_19187,N_17038,N_17499);
nand U19188 (N_19188,N_17611,N_17378);
xnor U19189 (N_19189,N_17923,N_16638);
xor U19190 (N_19190,N_16802,N_17773);
or U19191 (N_19191,N_16022,N_16640);
nand U19192 (N_19192,N_16070,N_16848);
nor U19193 (N_19193,N_17246,N_16872);
and U19194 (N_19194,N_16289,N_17345);
nand U19195 (N_19195,N_16930,N_16707);
nand U19196 (N_19196,N_17650,N_16709);
nand U19197 (N_19197,N_16160,N_17094);
or U19198 (N_19198,N_16091,N_17993);
nand U19199 (N_19199,N_17321,N_17514);
and U19200 (N_19200,N_17390,N_17370);
or U19201 (N_19201,N_16208,N_17622);
nor U19202 (N_19202,N_16925,N_17551);
nand U19203 (N_19203,N_16017,N_16062);
xor U19204 (N_19204,N_17302,N_17358);
nor U19205 (N_19205,N_16585,N_16698);
nand U19206 (N_19206,N_16109,N_16424);
or U19207 (N_19207,N_17516,N_17265);
and U19208 (N_19208,N_16571,N_16970);
or U19209 (N_19209,N_17741,N_17014);
and U19210 (N_19210,N_16434,N_16660);
nand U19211 (N_19211,N_16993,N_16440);
nand U19212 (N_19212,N_17457,N_17285);
or U19213 (N_19213,N_16617,N_17149);
or U19214 (N_19214,N_17184,N_17606);
nor U19215 (N_19215,N_17284,N_16278);
nor U19216 (N_19216,N_17631,N_17070);
nor U19217 (N_19217,N_16923,N_17015);
and U19218 (N_19218,N_17340,N_16335);
or U19219 (N_19219,N_17360,N_16311);
or U19220 (N_19220,N_16392,N_16756);
and U19221 (N_19221,N_16153,N_17153);
and U19222 (N_19222,N_17703,N_17130);
or U19223 (N_19223,N_16642,N_17876);
and U19224 (N_19224,N_16160,N_16915);
xnor U19225 (N_19225,N_16418,N_17834);
xnor U19226 (N_19226,N_16870,N_16970);
xnor U19227 (N_19227,N_16587,N_17671);
nor U19228 (N_19228,N_17496,N_16790);
nand U19229 (N_19229,N_16472,N_17448);
and U19230 (N_19230,N_16925,N_17847);
nor U19231 (N_19231,N_17585,N_17906);
or U19232 (N_19232,N_17174,N_17203);
or U19233 (N_19233,N_17575,N_17462);
or U19234 (N_19234,N_16404,N_17033);
nor U19235 (N_19235,N_17373,N_16910);
nand U19236 (N_19236,N_17974,N_17957);
and U19237 (N_19237,N_16995,N_17011);
nor U19238 (N_19238,N_17271,N_17639);
and U19239 (N_19239,N_17560,N_17427);
or U19240 (N_19240,N_17165,N_17511);
nand U19241 (N_19241,N_16553,N_17195);
or U19242 (N_19242,N_16882,N_17253);
or U19243 (N_19243,N_16114,N_17685);
xnor U19244 (N_19244,N_17792,N_16257);
nand U19245 (N_19245,N_17211,N_16887);
nand U19246 (N_19246,N_17869,N_16025);
and U19247 (N_19247,N_16816,N_16575);
xor U19248 (N_19248,N_16262,N_17249);
and U19249 (N_19249,N_16478,N_16533);
nor U19250 (N_19250,N_16855,N_17729);
xnor U19251 (N_19251,N_16718,N_16630);
xnor U19252 (N_19252,N_16688,N_17052);
nor U19253 (N_19253,N_16422,N_16538);
xor U19254 (N_19254,N_16910,N_17866);
nand U19255 (N_19255,N_17115,N_16302);
nand U19256 (N_19256,N_17468,N_16035);
xnor U19257 (N_19257,N_16837,N_16678);
and U19258 (N_19258,N_16136,N_17279);
or U19259 (N_19259,N_17434,N_16571);
nand U19260 (N_19260,N_17159,N_17774);
or U19261 (N_19261,N_16765,N_16012);
or U19262 (N_19262,N_16327,N_16937);
xor U19263 (N_19263,N_17505,N_17337);
nand U19264 (N_19264,N_16827,N_17192);
nand U19265 (N_19265,N_17050,N_16386);
nand U19266 (N_19266,N_17990,N_17324);
and U19267 (N_19267,N_17745,N_16268);
xor U19268 (N_19268,N_16002,N_17521);
nand U19269 (N_19269,N_17038,N_17714);
nand U19270 (N_19270,N_17819,N_17031);
xnor U19271 (N_19271,N_16461,N_17407);
or U19272 (N_19272,N_17488,N_16127);
or U19273 (N_19273,N_16900,N_17949);
and U19274 (N_19274,N_17183,N_17899);
xnor U19275 (N_19275,N_16927,N_16202);
nand U19276 (N_19276,N_16083,N_16923);
nand U19277 (N_19277,N_17405,N_16876);
or U19278 (N_19278,N_17883,N_17851);
and U19279 (N_19279,N_16656,N_16188);
nor U19280 (N_19280,N_16629,N_16363);
nand U19281 (N_19281,N_16371,N_17227);
or U19282 (N_19282,N_17935,N_16102);
or U19283 (N_19283,N_17364,N_16635);
nor U19284 (N_19284,N_16831,N_17147);
or U19285 (N_19285,N_17855,N_16597);
and U19286 (N_19286,N_17940,N_17615);
and U19287 (N_19287,N_16153,N_16526);
or U19288 (N_19288,N_17490,N_16831);
or U19289 (N_19289,N_16378,N_16016);
nor U19290 (N_19290,N_16771,N_16247);
and U19291 (N_19291,N_17999,N_17921);
xnor U19292 (N_19292,N_16791,N_17380);
xnor U19293 (N_19293,N_16604,N_17590);
nor U19294 (N_19294,N_17881,N_16346);
or U19295 (N_19295,N_16860,N_16934);
nand U19296 (N_19296,N_16304,N_16006);
nor U19297 (N_19297,N_16604,N_16432);
xor U19298 (N_19298,N_16107,N_17991);
xor U19299 (N_19299,N_17330,N_16366);
nor U19300 (N_19300,N_17924,N_16989);
and U19301 (N_19301,N_16718,N_16807);
or U19302 (N_19302,N_16653,N_16315);
or U19303 (N_19303,N_17629,N_17344);
xor U19304 (N_19304,N_16076,N_17894);
nor U19305 (N_19305,N_16314,N_16340);
xor U19306 (N_19306,N_16368,N_16504);
xor U19307 (N_19307,N_16956,N_16316);
nor U19308 (N_19308,N_17877,N_17068);
nand U19309 (N_19309,N_16034,N_17669);
or U19310 (N_19310,N_16178,N_17367);
nand U19311 (N_19311,N_17192,N_16625);
or U19312 (N_19312,N_16520,N_17104);
and U19313 (N_19313,N_17117,N_16860);
nor U19314 (N_19314,N_17491,N_16676);
and U19315 (N_19315,N_16535,N_17643);
nand U19316 (N_19316,N_16817,N_17033);
xor U19317 (N_19317,N_17176,N_17280);
or U19318 (N_19318,N_16644,N_16303);
or U19319 (N_19319,N_16166,N_16217);
nor U19320 (N_19320,N_17607,N_16661);
and U19321 (N_19321,N_17127,N_16614);
xor U19322 (N_19322,N_16176,N_17937);
nand U19323 (N_19323,N_17346,N_16208);
xor U19324 (N_19324,N_16756,N_16720);
and U19325 (N_19325,N_17163,N_17581);
and U19326 (N_19326,N_17544,N_16219);
nor U19327 (N_19327,N_17271,N_16906);
nor U19328 (N_19328,N_16239,N_16653);
nand U19329 (N_19329,N_17179,N_17524);
nand U19330 (N_19330,N_17747,N_16207);
or U19331 (N_19331,N_16802,N_17953);
or U19332 (N_19332,N_17842,N_16630);
and U19333 (N_19333,N_17896,N_16784);
nor U19334 (N_19334,N_17814,N_17210);
and U19335 (N_19335,N_17619,N_16955);
and U19336 (N_19336,N_17326,N_17660);
nor U19337 (N_19337,N_17531,N_17395);
nand U19338 (N_19338,N_16471,N_17161);
and U19339 (N_19339,N_16138,N_17271);
nand U19340 (N_19340,N_16259,N_16428);
xnor U19341 (N_19341,N_17468,N_17115);
or U19342 (N_19342,N_17015,N_16691);
and U19343 (N_19343,N_16358,N_17561);
xnor U19344 (N_19344,N_17172,N_17000);
and U19345 (N_19345,N_17479,N_17501);
or U19346 (N_19346,N_16826,N_17090);
nor U19347 (N_19347,N_16733,N_16990);
and U19348 (N_19348,N_17070,N_17953);
nand U19349 (N_19349,N_16595,N_16598);
and U19350 (N_19350,N_17074,N_17533);
xor U19351 (N_19351,N_16508,N_16845);
and U19352 (N_19352,N_17273,N_16955);
and U19353 (N_19353,N_17864,N_16557);
or U19354 (N_19354,N_16423,N_17165);
nor U19355 (N_19355,N_17773,N_16964);
or U19356 (N_19356,N_17070,N_17656);
nor U19357 (N_19357,N_17726,N_17845);
xor U19358 (N_19358,N_17191,N_17722);
and U19359 (N_19359,N_16069,N_16775);
and U19360 (N_19360,N_17015,N_17866);
xnor U19361 (N_19361,N_16277,N_17506);
nand U19362 (N_19362,N_17866,N_16779);
and U19363 (N_19363,N_17702,N_17649);
and U19364 (N_19364,N_16908,N_17020);
or U19365 (N_19365,N_17010,N_17393);
or U19366 (N_19366,N_16757,N_17686);
or U19367 (N_19367,N_16349,N_16582);
nand U19368 (N_19368,N_17340,N_17365);
xor U19369 (N_19369,N_17549,N_17373);
and U19370 (N_19370,N_16272,N_17993);
or U19371 (N_19371,N_17657,N_17588);
xnor U19372 (N_19372,N_16256,N_17894);
nor U19373 (N_19373,N_17768,N_17207);
or U19374 (N_19374,N_16136,N_17150);
and U19375 (N_19375,N_16091,N_16219);
nor U19376 (N_19376,N_16066,N_16211);
nor U19377 (N_19377,N_17166,N_17919);
nor U19378 (N_19378,N_16520,N_16987);
nor U19379 (N_19379,N_17607,N_17277);
nor U19380 (N_19380,N_17352,N_16166);
or U19381 (N_19381,N_16400,N_17209);
nand U19382 (N_19382,N_17965,N_17400);
or U19383 (N_19383,N_16953,N_17017);
xnor U19384 (N_19384,N_16755,N_17464);
and U19385 (N_19385,N_17256,N_16248);
xor U19386 (N_19386,N_17961,N_16747);
nor U19387 (N_19387,N_16805,N_17975);
nor U19388 (N_19388,N_17998,N_17292);
or U19389 (N_19389,N_16201,N_17673);
or U19390 (N_19390,N_17634,N_17980);
and U19391 (N_19391,N_17573,N_17826);
nand U19392 (N_19392,N_16210,N_17583);
and U19393 (N_19393,N_16368,N_16207);
xnor U19394 (N_19394,N_17203,N_17196);
and U19395 (N_19395,N_16401,N_17988);
nor U19396 (N_19396,N_17014,N_16869);
nand U19397 (N_19397,N_16373,N_16813);
xnor U19398 (N_19398,N_16591,N_16919);
nor U19399 (N_19399,N_17641,N_16470);
nand U19400 (N_19400,N_17269,N_16140);
and U19401 (N_19401,N_16389,N_16865);
xnor U19402 (N_19402,N_17194,N_17710);
and U19403 (N_19403,N_16117,N_16339);
nand U19404 (N_19404,N_17964,N_16121);
nor U19405 (N_19405,N_17730,N_16863);
and U19406 (N_19406,N_17299,N_17761);
and U19407 (N_19407,N_17227,N_16241);
or U19408 (N_19408,N_17801,N_17321);
xnor U19409 (N_19409,N_16939,N_17178);
nand U19410 (N_19410,N_16035,N_17799);
xnor U19411 (N_19411,N_17357,N_17812);
or U19412 (N_19412,N_16168,N_17420);
and U19413 (N_19413,N_17191,N_17023);
nor U19414 (N_19414,N_17354,N_16948);
and U19415 (N_19415,N_17801,N_16307);
xnor U19416 (N_19416,N_17559,N_17992);
nor U19417 (N_19417,N_17942,N_17525);
or U19418 (N_19418,N_16828,N_16582);
or U19419 (N_19419,N_17636,N_16637);
nand U19420 (N_19420,N_16202,N_16634);
and U19421 (N_19421,N_16227,N_17870);
nand U19422 (N_19422,N_17618,N_16087);
xor U19423 (N_19423,N_16346,N_17613);
nor U19424 (N_19424,N_16185,N_16332);
and U19425 (N_19425,N_16330,N_17407);
xor U19426 (N_19426,N_17764,N_17737);
xnor U19427 (N_19427,N_17396,N_16293);
xor U19428 (N_19428,N_16863,N_17336);
nor U19429 (N_19429,N_16200,N_17555);
xor U19430 (N_19430,N_17766,N_17902);
and U19431 (N_19431,N_17961,N_17739);
or U19432 (N_19432,N_17485,N_16150);
and U19433 (N_19433,N_17727,N_17934);
nand U19434 (N_19434,N_16510,N_17448);
xor U19435 (N_19435,N_16216,N_16874);
nand U19436 (N_19436,N_17248,N_16502);
nand U19437 (N_19437,N_16283,N_16543);
nor U19438 (N_19438,N_17735,N_17236);
nor U19439 (N_19439,N_17251,N_17040);
or U19440 (N_19440,N_17672,N_16560);
xor U19441 (N_19441,N_16312,N_17755);
or U19442 (N_19442,N_16421,N_17918);
nor U19443 (N_19443,N_17498,N_16928);
or U19444 (N_19444,N_16787,N_16367);
and U19445 (N_19445,N_17220,N_17473);
nand U19446 (N_19446,N_17621,N_17667);
or U19447 (N_19447,N_17722,N_17085);
xor U19448 (N_19448,N_17553,N_16623);
or U19449 (N_19449,N_17577,N_17748);
nand U19450 (N_19450,N_17877,N_17194);
or U19451 (N_19451,N_16513,N_16207);
nand U19452 (N_19452,N_16959,N_17253);
nand U19453 (N_19453,N_17259,N_17106);
nor U19454 (N_19454,N_16166,N_16614);
nand U19455 (N_19455,N_16761,N_17266);
nor U19456 (N_19456,N_17838,N_16737);
or U19457 (N_19457,N_16424,N_16008);
or U19458 (N_19458,N_17083,N_17973);
or U19459 (N_19459,N_16208,N_16266);
nand U19460 (N_19460,N_16773,N_17731);
nand U19461 (N_19461,N_17126,N_16381);
or U19462 (N_19462,N_17101,N_16775);
xor U19463 (N_19463,N_16508,N_16556);
xor U19464 (N_19464,N_16552,N_16672);
nand U19465 (N_19465,N_17318,N_16616);
xnor U19466 (N_19466,N_16147,N_16342);
or U19467 (N_19467,N_16049,N_16790);
or U19468 (N_19468,N_17430,N_16274);
or U19469 (N_19469,N_17516,N_17666);
and U19470 (N_19470,N_16101,N_16367);
nand U19471 (N_19471,N_16860,N_16114);
nand U19472 (N_19472,N_17880,N_16640);
nand U19473 (N_19473,N_16716,N_16111);
xnor U19474 (N_19474,N_17943,N_16465);
xor U19475 (N_19475,N_16615,N_16881);
xor U19476 (N_19476,N_16162,N_17654);
or U19477 (N_19477,N_17994,N_17945);
xnor U19478 (N_19478,N_16149,N_17196);
or U19479 (N_19479,N_17527,N_17229);
nor U19480 (N_19480,N_16025,N_16982);
and U19481 (N_19481,N_17210,N_16240);
xnor U19482 (N_19482,N_17769,N_17447);
xnor U19483 (N_19483,N_16299,N_16567);
nand U19484 (N_19484,N_16403,N_16244);
xnor U19485 (N_19485,N_16853,N_16245);
nand U19486 (N_19486,N_17505,N_17102);
xor U19487 (N_19487,N_17943,N_17642);
nor U19488 (N_19488,N_16144,N_16598);
or U19489 (N_19489,N_16996,N_17343);
nand U19490 (N_19490,N_17115,N_17726);
xnor U19491 (N_19491,N_16567,N_17213);
xor U19492 (N_19492,N_16620,N_16715);
nand U19493 (N_19493,N_16721,N_16124);
xor U19494 (N_19494,N_17410,N_16368);
and U19495 (N_19495,N_16766,N_16931);
nor U19496 (N_19496,N_17927,N_17178);
xnor U19497 (N_19497,N_16252,N_16739);
nor U19498 (N_19498,N_16193,N_17924);
or U19499 (N_19499,N_16994,N_16631);
nand U19500 (N_19500,N_17229,N_17779);
xnor U19501 (N_19501,N_17947,N_17133);
nand U19502 (N_19502,N_17413,N_16441);
and U19503 (N_19503,N_17683,N_17076);
xor U19504 (N_19504,N_16154,N_16923);
or U19505 (N_19505,N_17220,N_16617);
and U19506 (N_19506,N_16835,N_17078);
xor U19507 (N_19507,N_17802,N_16723);
xnor U19508 (N_19508,N_16204,N_16269);
nand U19509 (N_19509,N_16852,N_17864);
xnor U19510 (N_19510,N_17120,N_17969);
nor U19511 (N_19511,N_17400,N_16081);
or U19512 (N_19512,N_17260,N_16091);
xor U19513 (N_19513,N_16542,N_16088);
nor U19514 (N_19514,N_16040,N_16063);
and U19515 (N_19515,N_16274,N_16685);
and U19516 (N_19516,N_16646,N_17516);
nand U19517 (N_19517,N_16417,N_17298);
and U19518 (N_19518,N_16611,N_16987);
and U19519 (N_19519,N_16591,N_16510);
or U19520 (N_19520,N_16140,N_16205);
and U19521 (N_19521,N_16636,N_17680);
nor U19522 (N_19522,N_16268,N_17622);
and U19523 (N_19523,N_16112,N_17102);
xor U19524 (N_19524,N_16758,N_17656);
nand U19525 (N_19525,N_17848,N_16153);
and U19526 (N_19526,N_17514,N_16280);
or U19527 (N_19527,N_16844,N_16543);
and U19528 (N_19528,N_17356,N_17484);
nor U19529 (N_19529,N_17595,N_17415);
and U19530 (N_19530,N_16067,N_16896);
nand U19531 (N_19531,N_16213,N_17461);
nor U19532 (N_19532,N_17569,N_16957);
nor U19533 (N_19533,N_16607,N_17479);
and U19534 (N_19534,N_16970,N_17812);
nor U19535 (N_19535,N_16074,N_17409);
and U19536 (N_19536,N_16226,N_16748);
and U19537 (N_19537,N_16770,N_17758);
and U19538 (N_19538,N_16958,N_17578);
xnor U19539 (N_19539,N_17828,N_17734);
or U19540 (N_19540,N_17882,N_17601);
and U19541 (N_19541,N_16012,N_16100);
and U19542 (N_19542,N_17458,N_16692);
and U19543 (N_19543,N_17700,N_16961);
and U19544 (N_19544,N_16041,N_17462);
xnor U19545 (N_19545,N_16598,N_16120);
or U19546 (N_19546,N_16011,N_16478);
nor U19547 (N_19547,N_16382,N_16502);
xnor U19548 (N_19548,N_16539,N_16549);
nor U19549 (N_19549,N_16214,N_17604);
or U19550 (N_19550,N_17428,N_16639);
or U19551 (N_19551,N_17277,N_16207);
xnor U19552 (N_19552,N_17701,N_17209);
nor U19553 (N_19553,N_16380,N_16900);
and U19554 (N_19554,N_16818,N_16582);
xnor U19555 (N_19555,N_17356,N_17276);
or U19556 (N_19556,N_16520,N_16304);
xor U19557 (N_19557,N_17691,N_16331);
nand U19558 (N_19558,N_16161,N_16085);
nand U19559 (N_19559,N_16530,N_17000);
nor U19560 (N_19560,N_16412,N_17624);
nand U19561 (N_19561,N_17169,N_16219);
nand U19562 (N_19562,N_16591,N_16523);
nor U19563 (N_19563,N_16143,N_16091);
nand U19564 (N_19564,N_17123,N_17521);
and U19565 (N_19565,N_17418,N_16508);
or U19566 (N_19566,N_17305,N_17468);
nor U19567 (N_19567,N_16717,N_17431);
or U19568 (N_19568,N_17435,N_16098);
nand U19569 (N_19569,N_17831,N_16017);
xor U19570 (N_19570,N_16918,N_16175);
and U19571 (N_19571,N_16724,N_17536);
nand U19572 (N_19572,N_16876,N_17585);
or U19573 (N_19573,N_16665,N_16167);
or U19574 (N_19574,N_17083,N_16681);
and U19575 (N_19575,N_16089,N_16769);
or U19576 (N_19576,N_17143,N_17931);
nor U19577 (N_19577,N_16815,N_16765);
and U19578 (N_19578,N_17646,N_16740);
nand U19579 (N_19579,N_16920,N_17759);
and U19580 (N_19580,N_16341,N_17775);
nand U19581 (N_19581,N_17526,N_17302);
nand U19582 (N_19582,N_16222,N_16068);
nand U19583 (N_19583,N_17382,N_16310);
nand U19584 (N_19584,N_17588,N_17326);
xnor U19585 (N_19585,N_17818,N_17145);
and U19586 (N_19586,N_16800,N_16719);
xnor U19587 (N_19587,N_16070,N_16147);
nand U19588 (N_19588,N_17936,N_17132);
nor U19589 (N_19589,N_16739,N_16730);
and U19590 (N_19590,N_16032,N_17746);
and U19591 (N_19591,N_17985,N_16396);
nand U19592 (N_19592,N_16030,N_17962);
nor U19593 (N_19593,N_17244,N_17829);
xnor U19594 (N_19594,N_16356,N_17924);
nor U19595 (N_19595,N_16141,N_17271);
or U19596 (N_19596,N_17671,N_17819);
nor U19597 (N_19597,N_16653,N_16995);
nor U19598 (N_19598,N_16741,N_16187);
nand U19599 (N_19599,N_17266,N_16641);
xor U19600 (N_19600,N_16060,N_17661);
xor U19601 (N_19601,N_17448,N_17544);
and U19602 (N_19602,N_16648,N_17552);
or U19603 (N_19603,N_17081,N_16826);
nor U19604 (N_19604,N_16954,N_16920);
xor U19605 (N_19605,N_17233,N_17241);
xnor U19606 (N_19606,N_17033,N_17282);
nor U19607 (N_19607,N_17585,N_17823);
or U19608 (N_19608,N_17441,N_17357);
nand U19609 (N_19609,N_16695,N_16954);
and U19610 (N_19610,N_17247,N_17311);
or U19611 (N_19611,N_17040,N_17538);
xor U19612 (N_19612,N_17472,N_16954);
or U19613 (N_19613,N_17715,N_17042);
and U19614 (N_19614,N_17898,N_16773);
and U19615 (N_19615,N_17649,N_17060);
xor U19616 (N_19616,N_16794,N_16177);
or U19617 (N_19617,N_16123,N_16038);
or U19618 (N_19618,N_17657,N_16056);
nor U19619 (N_19619,N_16555,N_16128);
xor U19620 (N_19620,N_16610,N_17629);
nand U19621 (N_19621,N_17800,N_16102);
and U19622 (N_19622,N_17724,N_16083);
or U19623 (N_19623,N_16774,N_17380);
or U19624 (N_19624,N_17420,N_17095);
xnor U19625 (N_19625,N_17725,N_16979);
xnor U19626 (N_19626,N_17939,N_16033);
xor U19627 (N_19627,N_16360,N_16191);
and U19628 (N_19628,N_17383,N_16394);
or U19629 (N_19629,N_17086,N_17071);
nand U19630 (N_19630,N_17397,N_17381);
nor U19631 (N_19631,N_17411,N_16742);
nor U19632 (N_19632,N_16024,N_17398);
or U19633 (N_19633,N_16495,N_17765);
or U19634 (N_19634,N_16927,N_16877);
nand U19635 (N_19635,N_17461,N_16828);
or U19636 (N_19636,N_17565,N_16011);
or U19637 (N_19637,N_17274,N_17721);
xnor U19638 (N_19638,N_17201,N_17435);
nor U19639 (N_19639,N_16892,N_16001);
or U19640 (N_19640,N_16160,N_17466);
xor U19641 (N_19641,N_17363,N_17568);
and U19642 (N_19642,N_17314,N_17973);
and U19643 (N_19643,N_17294,N_17810);
and U19644 (N_19644,N_16630,N_17982);
nor U19645 (N_19645,N_16857,N_17414);
or U19646 (N_19646,N_17235,N_16306);
xnor U19647 (N_19647,N_16828,N_16371);
and U19648 (N_19648,N_16850,N_17772);
and U19649 (N_19649,N_17308,N_16474);
nor U19650 (N_19650,N_17608,N_17953);
nand U19651 (N_19651,N_17852,N_17998);
and U19652 (N_19652,N_17368,N_17161);
nand U19653 (N_19653,N_17268,N_16315);
nor U19654 (N_19654,N_16422,N_16565);
nand U19655 (N_19655,N_17868,N_16984);
and U19656 (N_19656,N_17485,N_17969);
or U19657 (N_19657,N_16575,N_17800);
nor U19658 (N_19658,N_17353,N_16408);
or U19659 (N_19659,N_17048,N_17293);
and U19660 (N_19660,N_17116,N_16653);
xnor U19661 (N_19661,N_16318,N_16936);
or U19662 (N_19662,N_16982,N_17527);
or U19663 (N_19663,N_17726,N_17195);
xor U19664 (N_19664,N_17985,N_16651);
nor U19665 (N_19665,N_17727,N_17446);
nand U19666 (N_19666,N_16591,N_16886);
and U19667 (N_19667,N_16775,N_16770);
xor U19668 (N_19668,N_16803,N_16929);
or U19669 (N_19669,N_16748,N_16593);
xnor U19670 (N_19670,N_16653,N_17035);
nand U19671 (N_19671,N_16409,N_17452);
or U19672 (N_19672,N_17650,N_16424);
nor U19673 (N_19673,N_17304,N_17212);
and U19674 (N_19674,N_17070,N_16059);
and U19675 (N_19675,N_17567,N_17147);
and U19676 (N_19676,N_16883,N_16995);
xor U19677 (N_19677,N_16438,N_17391);
xnor U19678 (N_19678,N_16710,N_17595);
nor U19679 (N_19679,N_16060,N_17032);
nand U19680 (N_19680,N_16210,N_17462);
and U19681 (N_19681,N_17397,N_16054);
nor U19682 (N_19682,N_17348,N_17514);
and U19683 (N_19683,N_17861,N_17000);
xor U19684 (N_19684,N_17414,N_17460);
xor U19685 (N_19685,N_16991,N_16975);
nor U19686 (N_19686,N_16496,N_16970);
or U19687 (N_19687,N_16111,N_17674);
nand U19688 (N_19688,N_17758,N_16587);
and U19689 (N_19689,N_17005,N_17724);
nand U19690 (N_19690,N_16181,N_16334);
and U19691 (N_19691,N_16022,N_16270);
nand U19692 (N_19692,N_17181,N_17467);
nand U19693 (N_19693,N_17404,N_17823);
or U19694 (N_19694,N_17293,N_16448);
nor U19695 (N_19695,N_17336,N_17970);
and U19696 (N_19696,N_17471,N_16385);
xnor U19697 (N_19697,N_16075,N_16146);
xnor U19698 (N_19698,N_16349,N_16139);
or U19699 (N_19699,N_16650,N_16615);
or U19700 (N_19700,N_16736,N_17033);
nor U19701 (N_19701,N_16295,N_16122);
xor U19702 (N_19702,N_16492,N_16760);
xor U19703 (N_19703,N_16216,N_16721);
xnor U19704 (N_19704,N_16032,N_16493);
nand U19705 (N_19705,N_16511,N_17311);
nand U19706 (N_19706,N_17846,N_16665);
nor U19707 (N_19707,N_17032,N_16792);
nand U19708 (N_19708,N_17043,N_17723);
or U19709 (N_19709,N_16705,N_17576);
and U19710 (N_19710,N_16826,N_17385);
nor U19711 (N_19711,N_17830,N_17389);
nand U19712 (N_19712,N_17410,N_16108);
xnor U19713 (N_19713,N_17679,N_17139);
nor U19714 (N_19714,N_17213,N_16348);
nor U19715 (N_19715,N_16173,N_16883);
or U19716 (N_19716,N_16153,N_17316);
nor U19717 (N_19717,N_16005,N_16438);
or U19718 (N_19718,N_17005,N_17223);
and U19719 (N_19719,N_17016,N_16271);
xnor U19720 (N_19720,N_16660,N_16422);
nand U19721 (N_19721,N_16499,N_16309);
or U19722 (N_19722,N_16010,N_16422);
and U19723 (N_19723,N_16136,N_16065);
and U19724 (N_19724,N_17594,N_16745);
or U19725 (N_19725,N_16000,N_16645);
and U19726 (N_19726,N_16782,N_16648);
or U19727 (N_19727,N_16261,N_17330);
or U19728 (N_19728,N_16524,N_17587);
or U19729 (N_19729,N_16747,N_16222);
nand U19730 (N_19730,N_16551,N_16662);
nand U19731 (N_19731,N_16535,N_16671);
xor U19732 (N_19732,N_16084,N_17959);
nor U19733 (N_19733,N_16123,N_17048);
and U19734 (N_19734,N_16424,N_17949);
xor U19735 (N_19735,N_16693,N_17502);
xnor U19736 (N_19736,N_17591,N_16536);
xor U19737 (N_19737,N_17812,N_17330);
nor U19738 (N_19738,N_16197,N_17894);
and U19739 (N_19739,N_17380,N_16097);
nand U19740 (N_19740,N_17194,N_16581);
nand U19741 (N_19741,N_16482,N_16540);
nor U19742 (N_19742,N_17833,N_16933);
and U19743 (N_19743,N_16150,N_17315);
xnor U19744 (N_19744,N_17023,N_17110);
and U19745 (N_19745,N_16211,N_17722);
and U19746 (N_19746,N_17796,N_17226);
nor U19747 (N_19747,N_17479,N_17123);
xor U19748 (N_19748,N_17618,N_16957);
and U19749 (N_19749,N_16133,N_16953);
or U19750 (N_19750,N_16452,N_17788);
nor U19751 (N_19751,N_16889,N_16460);
nor U19752 (N_19752,N_16974,N_16037);
or U19753 (N_19753,N_17247,N_17667);
or U19754 (N_19754,N_16057,N_16846);
xor U19755 (N_19755,N_17982,N_17493);
xnor U19756 (N_19756,N_17871,N_16090);
xor U19757 (N_19757,N_17736,N_16463);
nor U19758 (N_19758,N_16797,N_16565);
and U19759 (N_19759,N_16653,N_17067);
or U19760 (N_19760,N_17472,N_17021);
nand U19761 (N_19761,N_17212,N_17068);
and U19762 (N_19762,N_16679,N_17318);
and U19763 (N_19763,N_17369,N_17730);
nor U19764 (N_19764,N_16666,N_17008);
or U19765 (N_19765,N_16641,N_17683);
or U19766 (N_19766,N_16364,N_16527);
xnor U19767 (N_19767,N_16883,N_17699);
and U19768 (N_19768,N_17150,N_17970);
nand U19769 (N_19769,N_17385,N_16528);
nand U19770 (N_19770,N_16472,N_17642);
or U19771 (N_19771,N_17367,N_16336);
xor U19772 (N_19772,N_17990,N_17793);
nor U19773 (N_19773,N_17615,N_17181);
nand U19774 (N_19774,N_17510,N_16637);
or U19775 (N_19775,N_16492,N_16763);
nor U19776 (N_19776,N_17033,N_17063);
and U19777 (N_19777,N_17238,N_17246);
nand U19778 (N_19778,N_17595,N_17241);
or U19779 (N_19779,N_17610,N_17160);
xnor U19780 (N_19780,N_16139,N_17181);
and U19781 (N_19781,N_16694,N_17330);
xnor U19782 (N_19782,N_17097,N_17131);
and U19783 (N_19783,N_17589,N_17781);
or U19784 (N_19784,N_16305,N_16068);
nand U19785 (N_19785,N_16408,N_16681);
xor U19786 (N_19786,N_17441,N_17035);
or U19787 (N_19787,N_16349,N_16557);
nand U19788 (N_19788,N_17116,N_17966);
xnor U19789 (N_19789,N_17096,N_16800);
nor U19790 (N_19790,N_16285,N_17838);
nand U19791 (N_19791,N_16255,N_16664);
or U19792 (N_19792,N_16846,N_17043);
nor U19793 (N_19793,N_17511,N_17120);
nor U19794 (N_19794,N_17381,N_16742);
or U19795 (N_19795,N_17703,N_16198);
nor U19796 (N_19796,N_16795,N_17762);
xor U19797 (N_19797,N_16666,N_16357);
xnor U19798 (N_19798,N_17379,N_16984);
and U19799 (N_19799,N_17129,N_17966);
nand U19800 (N_19800,N_16163,N_16371);
and U19801 (N_19801,N_17312,N_16371);
and U19802 (N_19802,N_16733,N_17221);
nand U19803 (N_19803,N_16800,N_16284);
xnor U19804 (N_19804,N_17909,N_17910);
and U19805 (N_19805,N_16679,N_16189);
nand U19806 (N_19806,N_17770,N_17400);
nor U19807 (N_19807,N_17871,N_16377);
nand U19808 (N_19808,N_16783,N_16740);
and U19809 (N_19809,N_17248,N_17647);
nand U19810 (N_19810,N_17945,N_16233);
and U19811 (N_19811,N_17011,N_16032);
and U19812 (N_19812,N_17793,N_16524);
or U19813 (N_19813,N_17733,N_17382);
nand U19814 (N_19814,N_17874,N_17601);
xor U19815 (N_19815,N_17857,N_17471);
nor U19816 (N_19816,N_16121,N_16041);
and U19817 (N_19817,N_17256,N_16728);
xor U19818 (N_19818,N_16959,N_16914);
nor U19819 (N_19819,N_16362,N_17279);
xor U19820 (N_19820,N_17248,N_17077);
nor U19821 (N_19821,N_17240,N_16792);
and U19822 (N_19822,N_16882,N_17387);
or U19823 (N_19823,N_17727,N_17846);
nor U19824 (N_19824,N_16158,N_16939);
or U19825 (N_19825,N_16511,N_17759);
nor U19826 (N_19826,N_17671,N_16022);
xor U19827 (N_19827,N_17827,N_17419);
xor U19828 (N_19828,N_17968,N_17484);
nor U19829 (N_19829,N_17167,N_16123);
nand U19830 (N_19830,N_17158,N_17505);
nand U19831 (N_19831,N_17269,N_17704);
xnor U19832 (N_19832,N_16492,N_17345);
or U19833 (N_19833,N_17979,N_17656);
nand U19834 (N_19834,N_16466,N_17770);
nor U19835 (N_19835,N_17770,N_17902);
nand U19836 (N_19836,N_17526,N_16534);
nor U19837 (N_19837,N_17435,N_16099);
nand U19838 (N_19838,N_17445,N_16562);
xnor U19839 (N_19839,N_16368,N_16482);
nand U19840 (N_19840,N_16889,N_17917);
xor U19841 (N_19841,N_17583,N_16370);
and U19842 (N_19842,N_16703,N_16867);
xnor U19843 (N_19843,N_16245,N_17159);
or U19844 (N_19844,N_17406,N_16347);
or U19845 (N_19845,N_17089,N_16951);
xor U19846 (N_19846,N_17810,N_16366);
and U19847 (N_19847,N_17645,N_17704);
nor U19848 (N_19848,N_17749,N_17053);
xor U19849 (N_19849,N_16440,N_16535);
nand U19850 (N_19850,N_16578,N_17546);
nor U19851 (N_19851,N_17013,N_17100);
nor U19852 (N_19852,N_16026,N_16608);
nand U19853 (N_19853,N_17700,N_16741);
or U19854 (N_19854,N_16469,N_16156);
nand U19855 (N_19855,N_16514,N_16503);
and U19856 (N_19856,N_17549,N_16084);
or U19857 (N_19857,N_17220,N_17785);
nor U19858 (N_19858,N_17330,N_17846);
nor U19859 (N_19859,N_17817,N_17090);
nor U19860 (N_19860,N_16808,N_16371);
nand U19861 (N_19861,N_16968,N_16423);
nand U19862 (N_19862,N_16984,N_17752);
xor U19863 (N_19863,N_17532,N_16040);
and U19864 (N_19864,N_16142,N_17581);
and U19865 (N_19865,N_16156,N_17831);
xnor U19866 (N_19866,N_17002,N_16424);
and U19867 (N_19867,N_17096,N_16761);
xnor U19868 (N_19868,N_17680,N_17461);
nand U19869 (N_19869,N_16540,N_16657);
nand U19870 (N_19870,N_16382,N_16282);
nand U19871 (N_19871,N_17946,N_16573);
and U19872 (N_19872,N_16432,N_16424);
nand U19873 (N_19873,N_16851,N_17165);
or U19874 (N_19874,N_17119,N_16965);
or U19875 (N_19875,N_17994,N_16607);
xnor U19876 (N_19876,N_17574,N_16817);
and U19877 (N_19877,N_17880,N_17356);
xnor U19878 (N_19878,N_17924,N_16686);
nor U19879 (N_19879,N_16108,N_16899);
xor U19880 (N_19880,N_16571,N_16372);
xor U19881 (N_19881,N_17984,N_16041);
and U19882 (N_19882,N_16268,N_17047);
nor U19883 (N_19883,N_16721,N_16170);
nor U19884 (N_19884,N_17434,N_16643);
nand U19885 (N_19885,N_17330,N_16403);
nor U19886 (N_19886,N_16489,N_16418);
and U19887 (N_19887,N_17732,N_17604);
nor U19888 (N_19888,N_17063,N_16246);
and U19889 (N_19889,N_16707,N_16153);
or U19890 (N_19890,N_16175,N_17053);
or U19891 (N_19891,N_16713,N_17128);
xnor U19892 (N_19892,N_17966,N_17982);
xnor U19893 (N_19893,N_17546,N_16497);
or U19894 (N_19894,N_17872,N_17793);
or U19895 (N_19895,N_17300,N_17528);
xor U19896 (N_19896,N_17421,N_16421);
nor U19897 (N_19897,N_17126,N_17885);
or U19898 (N_19898,N_16235,N_17502);
nor U19899 (N_19899,N_16940,N_16158);
nor U19900 (N_19900,N_17657,N_17802);
nor U19901 (N_19901,N_16486,N_17198);
and U19902 (N_19902,N_16463,N_16963);
nand U19903 (N_19903,N_17899,N_16156);
or U19904 (N_19904,N_17386,N_17402);
or U19905 (N_19905,N_17138,N_16379);
xor U19906 (N_19906,N_17588,N_17414);
nor U19907 (N_19907,N_17096,N_16771);
or U19908 (N_19908,N_17660,N_16674);
nand U19909 (N_19909,N_17962,N_17535);
xnor U19910 (N_19910,N_17310,N_17991);
or U19911 (N_19911,N_16414,N_17052);
nor U19912 (N_19912,N_17610,N_17408);
nand U19913 (N_19913,N_16955,N_16764);
and U19914 (N_19914,N_16170,N_16359);
nor U19915 (N_19915,N_16781,N_16261);
xor U19916 (N_19916,N_17178,N_16058);
nand U19917 (N_19917,N_17796,N_16281);
and U19918 (N_19918,N_16584,N_16779);
xnor U19919 (N_19919,N_17124,N_16164);
nor U19920 (N_19920,N_17091,N_17992);
and U19921 (N_19921,N_16649,N_16409);
nor U19922 (N_19922,N_17654,N_17917);
nand U19923 (N_19923,N_16528,N_16023);
or U19924 (N_19924,N_16580,N_16161);
xor U19925 (N_19925,N_17615,N_17750);
and U19926 (N_19926,N_16124,N_17409);
or U19927 (N_19927,N_17029,N_17253);
and U19928 (N_19928,N_16733,N_16796);
nand U19929 (N_19929,N_16350,N_17720);
or U19930 (N_19930,N_17653,N_16449);
xor U19931 (N_19931,N_17358,N_16480);
nor U19932 (N_19932,N_17681,N_16051);
nor U19933 (N_19933,N_16749,N_17026);
xnor U19934 (N_19934,N_16407,N_17744);
nor U19935 (N_19935,N_16881,N_16078);
nand U19936 (N_19936,N_17782,N_16529);
and U19937 (N_19937,N_16289,N_17083);
xor U19938 (N_19938,N_17847,N_17061);
nor U19939 (N_19939,N_17280,N_17553);
nor U19940 (N_19940,N_16228,N_17304);
and U19941 (N_19941,N_17153,N_17320);
xor U19942 (N_19942,N_16602,N_17129);
or U19943 (N_19943,N_17936,N_17172);
xor U19944 (N_19944,N_16212,N_17619);
nand U19945 (N_19945,N_17018,N_16270);
or U19946 (N_19946,N_17674,N_16513);
nand U19947 (N_19947,N_16431,N_17848);
or U19948 (N_19948,N_16880,N_16996);
and U19949 (N_19949,N_16750,N_16409);
and U19950 (N_19950,N_16807,N_16621);
or U19951 (N_19951,N_17596,N_16395);
and U19952 (N_19952,N_17950,N_17174);
nand U19953 (N_19953,N_17804,N_16969);
nor U19954 (N_19954,N_16063,N_17723);
nand U19955 (N_19955,N_17228,N_16619);
and U19956 (N_19956,N_17153,N_17048);
xnor U19957 (N_19957,N_17476,N_17876);
or U19958 (N_19958,N_17698,N_16751);
or U19959 (N_19959,N_17296,N_16844);
xor U19960 (N_19960,N_16817,N_17929);
nor U19961 (N_19961,N_16278,N_17914);
nor U19962 (N_19962,N_16717,N_16630);
or U19963 (N_19963,N_17368,N_16642);
nor U19964 (N_19964,N_16956,N_17610);
or U19965 (N_19965,N_16195,N_17600);
xnor U19966 (N_19966,N_16692,N_16403);
nor U19967 (N_19967,N_17811,N_17694);
or U19968 (N_19968,N_17743,N_16435);
or U19969 (N_19969,N_17841,N_17990);
and U19970 (N_19970,N_16226,N_17122);
nand U19971 (N_19971,N_17670,N_16000);
nor U19972 (N_19972,N_17033,N_16909);
and U19973 (N_19973,N_16687,N_16610);
and U19974 (N_19974,N_17411,N_17674);
nand U19975 (N_19975,N_16091,N_16243);
xor U19976 (N_19976,N_16174,N_17183);
xnor U19977 (N_19977,N_16915,N_16450);
and U19978 (N_19978,N_17719,N_17744);
and U19979 (N_19979,N_16025,N_16468);
xor U19980 (N_19980,N_16975,N_17299);
nor U19981 (N_19981,N_16215,N_17304);
and U19982 (N_19982,N_16211,N_17795);
and U19983 (N_19983,N_17655,N_17753);
or U19984 (N_19984,N_16992,N_17223);
xnor U19985 (N_19985,N_17346,N_16894);
nor U19986 (N_19986,N_16960,N_16759);
and U19987 (N_19987,N_17541,N_17026);
nand U19988 (N_19988,N_17169,N_17385);
nand U19989 (N_19989,N_16651,N_16578);
and U19990 (N_19990,N_16258,N_17498);
nand U19991 (N_19991,N_16976,N_17553);
nand U19992 (N_19992,N_17471,N_16364);
nand U19993 (N_19993,N_16522,N_16531);
and U19994 (N_19994,N_16760,N_17625);
xnor U19995 (N_19995,N_17084,N_17054);
and U19996 (N_19996,N_17564,N_17278);
nor U19997 (N_19997,N_17867,N_16638);
nand U19998 (N_19998,N_17962,N_17211);
nand U19999 (N_19999,N_17961,N_16076);
nand U20000 (N_20000,N_19780,N_19980);
xnor U20001 (N_20001,N_19066,N_18008);
xor U20002 (N_20002,N_18745,N_19298);
nand U20003 (N_20003,N_18566,N_19046);
and U20004 (N_20004,N_18575,N_18472);
nand U20005 (N_20005,N_18957,N_19366);
xor U20006 (N_20006,N_18191,N_19147);
nor U20007 (N_20007,N_19671,N_18609);
and U20008 (N_20008,N_19747,N_19941);
nand U20009 (N_20009,N_18145,N_19678);
nand U20010 (N_20010,N_19617,N_18089);
xor U20011 (N_20011,N_19981,N_18372);
nor U20012 (N_20012,N_18662,N_18031);
xnor U20013 (N_20013,N_18080,N_18385);
nand U20014 (N_20014,N_19216,N_19084);
and U20015 (N_20015,N_19207,N_19561);
nor U20016 (N_20016,N_19319,N_18898);
xor U20017 (N_20017,N_18610,N_18862);
and U20018 (N_20018,N_18180,N_18787);
nand U20019 (N_20019,N_19797,N_19406);
and U20020 (N_20020,N_18932,N_19894);
nor U20021 (N_20021,N_18311,N_18552);
or U20022 (N_20022,N_19338,N_18348);
or U20023 (N_20023,N_19200,N_19361);
xnor U20024 (N_20024,N_19015,N_19988);
and U20025 (N_20025,N_19893,N_18707);
xor U20026 (N_20026,N_18785,N_18933);
nor U20027 (N_20027,N_18087,N_18593);
nand U20028 (N_20028,N_18510,N_19533);
and U20029 (N_20029,N_18527,N_19815);
xor U20030 (N_20030,N_19859,N_19189);
nor U20031 (N_20031,N_18751,N_18377);
xor U20032 (N_20032,N_18924,N_19929);
nor U20033 (N_20033,N_19841,N_18734);
and U20034 (N_20034,N_18847,N_19494);
nor U20035 (N_20035,N_18749,N_19399);
xnor U20036 (N_20036,N_18840,N_19590);
and U20037 (N_20037,N_18339,N_19737);
nor U20038 (N_20038,N_18220,N_18367);
or U20039 (N_20039,N_18615,N_18402);
nand U20040 (N_20040,N_18403,N_18506);
nand U20041 (N_20041,N_19769,N_18284);
nand U20042 (N_20042,N_19685,N_18845);
nor U20043 (N_20043,N_18926,N_18194);
xnor U20044 (N_20044,N_18184,N_18052);
nor U20045 (N_20045,N_18897,N_19720);
and U20046 (N_20046,N_19902,N_18571);
and U20047 (N_20047,N_19208,N_18303);
xor U20048 (N_20048,N_18318,N_19595);
xor U20049 (N_20049,N_18490,N_18717);
xnor U20050 (N_20050,N_18990,N_18783);
or U20051 (N_20051,N_18983,N_19693);
and U20052 (N_20052,N_18873,N_19805);
nor U20053 (N_20053,N_18190,N_19257);
xnor U20054 (N_20054,N_19967,N_19479);
nand U20055 (N_20055,N_19295,N_18305);
nor U20056 (N_20056,N_18193,N_18138);
or U20057 (N_20057,N_19634,N_18558);
nor U20058 (N_20058,N_18005,N_19175);
xnor U20059 (N_20059,N_18657,N_19477);
and U20060 (N_20060,N_18442,N_18480);
xnor U20061 (N_20061,N_18432,N_19545);
xor U20062 (N_20062,N_18117,N_18820);
nand U20063 (N_20063,N_19370,N_18248);
or U20064 (N_20064,N_18104,N_19122);
nand U20065 (N_20065,N_18386,N_18391);
nor U20066 (N_20066,N_18469,N_19924);
nor U20067 (N_20067,N_18896,N_18221);
nor U20068 (N_20068,N_19497,N_19485);
or U20069 (N_20069,N_18178,N_19936);
xor U20070 (N_20070,N_19251,N_19622);
xor U20071 (N_20071,N_19717,N_18400);
nand U20072 (N_20072,N_18369,N_18226);
nand U20073 (N_20073,N_19968,N_19708);
nand U20074 (N_20074,N_18353,N_19254);
xnor U20075 (N_20075,N_18186,N_19184);
or U20076 (N_20076,N_18078,N_19198);
xor U20077 (N_20077,N_19349,N_19410);
and U20078 (N_20078,N_19726,N_19882);
or U20079 (N_20079,N_18539,N_19703);
and U20080 (N_20080,N_18054,N_19579);
or U20081 (N_20081,N_19195,N_19362);
or U20082 (N_20082,N_19935,N_19178);
or U20083 (N_20083,N_18109,N_19445);
nand U20084 (N_20084,N_19713,N_18895);
nand U20085 (N_20085,N_19812,N_18635);
or U20086 (N_20086,N_19912,N_18413);
xnor U20087 (N_20087,N_18953,N_19526);
and U20088 (N_20088,N_18972,N_19984);
nor U20089 (N_20089,N_18686,N_19647);
nor U20090 (N_20090,N_18202,N_19067);
nand U20091 (N_20091,N_19193,N_19766);
or U20092 (N_20092,N_19762,N_19773);
xor U20093 (N_20093,N_19456,N_18766);
or U20094 (N_20094,N_19017,N_19138);
nand U20095 (N_20095,N_19746,N_19256);
xor U20096 (N_20096,N_19642,N_19565);
nand U20097 (N_20097,N_19356,N_19413);
nor U20098 (N_20098,N_19297,N_18324);
or U20099 (N_20099,N_18126,N_19055);
and U20100 (N_20100,N_18894,N_19520);
xor U20101 (N_20101,N_19679,N_18482);
nand U20102 (N_20102,N_18904,N_19652);
or U20103 (N_20103,N_18863,N_19172);
nor U20104 (N_20104,N_18310,N_19846);
or U20105 (N_20105,N_19644,N_18028);
or U20106 (N_20106,N_19457,N_18146);
nand U20107 (N_20107,N_18498,N_19990);
and U20108 (N_20108,N_18656,N_18546);
nand U20109 (N_20109,N_19535,N_18105);
or U20110 (N_20110,N_19306,N_19111);
xnor U20111 (N_20111,N_19329,N_19684);
xnor U20112 (N_20112,N_19016,N_19830);
nand U20113 (N_20113,N_19415,N_18663);
and U20114 (N_20114,N_19301,N_19408);
or U20115 (N_20115,N_19896,N_19355);
or U20116 (N_20116,N_19618,N_18670);
nor U20117 (N_20117,N_18010,N_19752);
xnor U20118 (N_20118,N_19978,N_18659);
xor U20119 (N_20119,N_18815,N_18633);
xor U20120 (N_20120,N_18965,N_19538);
or U20121 (N_20121,N_19222,N_19441);
nor U20122 (N_20122,N_18450,N_19630);
nand U20123 (N_20123,N_18712,N_19887);
or U20124 (N_20124,N_19788,N_19648);
and U20125 (N_20125,N_19043,N_19664);
and U20126 (N_20126,N_19464,N_18974);
or U20127 (N_20127,N_18903,N_19710);
and U20128 (N_20128,N_19613,N_18411);
nand U20129 (N_20129,N_18379,N_19059);
xnor U20130 (N_20130,N_19435,N_18286);
and U20131 (N_20131,N_18959,N_19164);
and U20132 (N_20132,N_19916,N_19691);
and U20133 (N_20133,N_18017,N_19080);
nor U20134 (N_20134,N_19921,N_18298);
or U20135 (N_20135,N_18042,N_19280);
or U20136 (N_20136,N_18595,N_19637);
nor U20137 (N_20137,N_18487,N_19285);
xnor U20138 (N_20138,N_18878,N_19834);
or U20139 (N_20139,N_19753,N_18503);
or U20140 (N_20140,N_18362,N_18338);
nand U20141 (N_20141,N_18171,N_19099);
and U20142 (N_20142,N_19000,N_19476);
nor U20143 (N_20143,N_19816,N_18619);
nand U20144 (N_20144,N_18134,N_18790);
xnor U20145 (N_20145,N_19144,N_19194);
xor U20146 (N_20146,N_18922,N_18465);
nor U20147 (N_20147,N_19422,N_19934);
nor U20148 (N_20148,N_19471,N_19865);
or U20149 (N_20149,N_18777,N_18299);
nand U20150 (N_20150,N_18557,N_19149);
and U20151 (N_20151,N_19969,N_18130);
nor U20152 (N_20152,N_18927,N_19230);
nand U20153 (N_20153,N_19312,N_19885);
and U20154 (N_20154,N_19872,N_18312);
and U20155 (N_20155,N_18053,N_19548);
and U20156 (N_20156,N_18675,N_18810);
or U20157 (N_20157,N_18817,N_18275);
xor U20158 (N_20158,N_18750,N_19959);
nor U20159 (N_20159,N_19250,N_18660);
nand U20160 (N_20160,N_18113,N_18481);
or U20161 (N_20161,N_18405,N_19443);
nor U20162 (N_20162,N_19334,N_19440);
or U20163 (N_20163,N_19442,N_19363);
nand U20164 (N_20164,N_18233,N_19377);
nand U20165 (N_20165,N_19542,N_18131);
xnor U20166 (N_20166,N_19819,N_18024);
nor U20167 (N_20167,N_18292,N_18531);
nand U20168 (N_20168,N_19150,N_18371);
xnor U20169 (N_20169,N_19009,N_19465);
and U20170 (N_20170,N_19192,N_19234);
xor U20171 (N_20171,N_19392,N_18097);
nand U20172 (N_20172,N_18996,N_19369);
nor U20173 (N_20173,N_19789,N_18437);
nor U20174 (N_20174,N_19086,N_18685);
xnor U20175 (N_20175,N_19578,N_18910);
or U20176 (N_20176,N_19202,N_18645);
or U20177 (N_20177,N_19263,N_18611);
and U20178 (N_20178,N_19657,N_18860);
nor U20179 (N_20179,N_19970,N_19026);
and U20180 (N_20180,N_19877,N_18940);
xor U20181 (N_20181,N_18003,N_19601);
nor U20182 (N_20182,N_18929,N_19725);
nand U20183 (N_20183,N_18501,N_18175);
nand U20184 (N_20184,N_19448,N_18524);
nand U20185 (N_20185,N_18417,N_19236);
or U20186 (N_20186,N_19845,N_18401);
nand U20187 (N_20187,N_19426,N_18759);
xnor U20188 (N_20188,N_19958,N_19418);
or U20189 (N_20189,N_19231,N_18197);
nand U20190 (N_20190,N_18522,N_19760);
xnor U20191 (N_20191,N_19564,N_18889);
nand U20192 (N_20192,N_19809,N_18573);
xor U20193 (N_20193,N_19499,N_19032);
and U20194 (N_20194,N_18466,N_18364);
nand U20195 (N_20195,N_18781,N_19927);
or U20196 (N_20196,N_19472,N_19770);
and U20197 (N_20197,N_18692,N_19714);
nand U20198 (N_20198,N_19566,N_19531);
nand U20199 (N_20199,N_19719,N_19417);
xnor U20200 (N_20200,N_19856,N_19640);
nand U20201 (N_20201,N_19955,N_19358);
and U20202 (N_20202,N_18051,N_19064);
and U20203 (N_20203,N_19239,N_18690);
nor U20204 (N_20204,N_18969,N_18628);
or U20205 (N_20205,N_19274,N_18512);
or U20206 (N_20206,N_18560,N_19555);
or U20207 (N_20207,N_19133,N_19300);
xnor U20208 (N_20208,N_18828,N_18136);
or U20209 (N_20209,N_18824,N_19534);
xor U20210 (N_20210,N_19090,N_18947);
nor U20211 (N_20211,N_18276,N_18746);
nand U20212 (N_20212,N_18906,N_19848);
nand U20213 (N_20213,N_19906,N_18551);
and U20214 (N_20214,N_19028,N_18326);
nand U20215 (N_20215,N_18673,N_19748);
nand U20216 (N_20216,N_19022,N_18971);
and U20217 (N_20217,N_18687,N_19074);
nor U20218 (N_20218,N_18913,N_18306);
and U20219 (N_20219,N_19658,N_19179);
or U20220 (N_20220,N_19718,N_19271);
nor U20221 (N_20221,N_19705,N_18638);
nand U20222 (N_20222,N_18916,N_19614);
xnor U20223 (N_20223,N_19842,N_19326);
or U20224 (N_20224,N_19911,N_19414);
nand U20225 (N_20225,N_19076,N_19977);
nor U20226 (N_20226,N_18963,N_18977);
and U20227 (N_20227,N_19488,N_19143);
xnor U20228 (N_20228,N_19284,N_18547);
xnor U20229 (N_20229,N_18398,N_19145);
xor U20230 (N_20230,N_19732,N_18647);
nand U20231 (N_20231,N_18223,N_19134);
nor U20232 (N_20232,N_19563,N_18095);
and U20233 (N_20233,N_18128,N_18544);
or U20234 (N_20234,N_18714,N_18370);
nand U20235 (N_20235,N_19556,N_19128);
or U20236 (N_20236,N_19123,N_18960);
and U20237 (N_20237,N_18949,N_18020);
nand U20238 (N_20238,N_18701,N_19518);
nor U20239 (N_20239,N_19467,N_19591);
nor U20240 (N_20240,N_18049,N_18899);
and U20241 (N_20241,N_19768,N_19828);
or U20242 (N_20242,N_19003,N_19330);
or U20243 (N_20243,N_19574,N_19930);
nor U20244 (N_20244,N_18945,N_19690);
and U20245 (N_20245,N_18259,N_18718);
xnor U20246 (N_20246,N_19480,N_18724);
and U20247 (N_20247,N_18112,N_19135);
xor U20248 (N_20248,N_19757,N_18076);
or U20249 (N_20249,N_18967,N_19100);
or U20250 (N_20250,N_19940,N_18943);
or U20251 (N_20251,N_18637,N_19381);
xnor U20252 (N_20252,N_19082,N_19754);
xnor U20253 (N_20253,N_19651,N_18846);
or U20254 (N_20254,N_18856,N_18827);
and U20255 (N_20255,N_18300,N_18640);
xor U20256 (N_20256,N_18597,N_18886);
and U20257 (N_20257,N_18606,N_18302);
nor U20258 (N_20258,N_19199,N_18954);
and U20259 (N_20259,N_18388,N_18731);
nor U20260 (N_20260,N_18858,N_19077);
nor U20261 (N_20261,N_18537,N_19108);
and U20262 (N_20262,N_19364,N_18604);
nand U20263 (N_20263,N_19779,N_19458);
nor U20264 (N_20264,N_18463,N_19552);
and U20265 (N_20265,N_18309,N_18448);
and U20266 (N_20266,N_18564,N_19801);
or U20267 (N_20267,N_18956,N_19455);
nand U20268 (N_20268,N_19982,N_19851);
xor U20269 (N_20269,N_19901,N_19771);
nor U20270 (N_20270,N_18885,N_18019);
or U20271 (N_20271,N_19037,N_18681);
and U20272 (N_20272,N_19079,N_18151);
or U20273 (N_20273,N_19504,N_19127);
xnor U20274 (N_20274,N_18455,N_19947);
nand U20275 (N_20275,N_18941,N_19803);
or U20276 (N_20276,N_18639,N_18703);
and U20277 (N_20277,N_19822,N_18509);
nand U20278 (N_20278,N_19148,N_18819);
xnor U20279 (N_20279,N_19394,N_19174);
xor U20280 (N_20280,N_18587,N_18525);
nand U20281 (N_20281,N_18380,N_18617);
nand U20282 (N_20282,N_19191,N_19107);
and U20283 (N_20283,N_19683,N_19359);
and U20284 (N_20284,N_18409,N_19914);
xor U20285 (N_20285,N_18110,N_19873);
and U20286 (N_20286,N_19162,N_19142);
nor U20287 (N_20287,N_18037,N_18174);
nand U20288 (N_20288,N_19867,N_18461);
or U20289 (N_20289,N_19058,N_18278);
nand U20290 (N_20290,N_19811,N_19049);
nor U20291 (N_20291,N_18211,N_19689);
or U20292 (N_20292,N_18453,N_19129);
nand U20293 (N_20293,N_19633,N_19573);
nand U20294 (N_20294,N_18156,N_18540);
and U20295 (N_20295,N_18315,N_18073);
or U20296 (N_20296,N_18142,N_18082);
nand U20297 (N_20297,N_18358,N_19875);
nor U20298 (N_20298,N_18242,N_19273);
nand U20299 (N_20299,N_19351,N_19692);
and U20300 (N_20300,N_19840,N_18561);
and U20301 (N_20301,N_18317,N_19081);
nor U20302 (N_20302,N_18901,N_19165);
and U20303 (N_20303,N_19388,N_19506);
nand U20304 (N_20304,N_18767,N_19401);
and U20305 (N_20305,N_19020,N_19511);
nor U20306 (N_20306,N_18804,N_18022);
and U20307 (N_20307,N_18231,N_19806);
nand U20308 (N_20308,N_19034,N_19201);
or U20309 (N_20309,N_19772,N_18255);
and U20310 (N_20310,N_18955,N_18702);
and U20311 (N_20311,N_18486,N_18296);
nand U20312 (N_20312,N_19068,N_18252);
or U20313 (N_20313,N_19957,N_18986);
or U20314 (N_20314,N_19728,N_19209);
or U20315 (N_20315,N_18050,N_19831);
nand U20316 (N_20316,N_18599,N_19682);
xnor U20317 (N_20317,N_18664,N_18631);
or U20318 (N_20318,N_19814,N_19006);
or U20319 (N_20319,N_19843,N_18260);
nand U20320 (N_20320,N_18406,N_18327);
and U20321 (N_20321,N_19001,N_18241);
nor U20322 (N_20322,N_18500,N_18594);
nand U20323 (N_20323,N_18934,N_18596);
nand U20324 (N_20324,N_18213,N_18891);
and U20325 (N_20325,N_18267,N_19949);
xnor U20326 (N_20326,N_18449,N_19764);
nand U20327 (N_20327,N_19599,N_18313);
or U20328 (N_20328,N_19153,N_19701);
or U20329 (N_20329,N_19227,N_19668);
nand U20330 (N_20330,N_19268,N_19821);
xor U20331 (N_20331,N_18133,N_18307);
and U20332 (N_20332,N_18835,N_19343);
and U20333 (N_20333,N_19745,N_19289);
and U20334 (N_20334,N_18834,N_18408);
and U20335 (N_20335,N_18568,N_18565);
or U20336 (N_20336,N_18581,N_19093);
nand U20337 (N_20337,N_18736,N_18928);
nand U20338 (N_20338,N_19986,N_18484);
xor U20339 (N_20339,N_19501,N_18875);
xor U20340 (N_20340,N_19791,N_19562);
nor U20341 (N_20341,N_18550,N_19375);
nand U20342 (N_20342,N_19372,N_18841);
or U20343 (N_20343,N_19795,N_19242);
and U20344 (N_20344,N_19182,N_19557);
nand U20345 (N_20345,N_19799,N_18396);
or U20346 (N_20346,N_19808,N_18980);
or U20347 (N_20347,N_19196,N_19505);
or U20348 (N_20348,N_19035,N_19804);
xor U20349 (N_20349,N_18011,N_18813);
or U20350 (N_20350,N_19010,N_19054);
xor U20351 (N_20351,N_19489,N_18948);
xnor U20352 (N_20352,N_19224,N_19669);
or U20353 (N_20353,N_19405,N_18084);
or U20354 (N_20354,N_19248,N_19121);
nand U20355 (N_20355,N_18831,N_18458);
or U20356 (N_20356,N_18798,N_18730);
nor U20357 (N_20357,N_18061,N_18789);
nand U20358 (N_20358,N_18739,N_19181);
nand U20359 (N_20359,N_18009,N_19004);
xor U20360 (N_20360,N_19785,N_18602);
xnor U20361 (N_20361,N_19519,N_19626);
and U20362 (N_20362,N_19249,N_18183);
nand U20363 (N_20363,N_19204,N_19582);
nand U20364 (N_20364,N_19820,N_18689);
and U20365 (N_20365,N_18976,N_18648);
nor U20366 (N_20366,N_18691,N_19641);
and U20367 (N_20367,N_19083,N_18607);
xnor U20368 (N_20368,N_19400,N_18880);
nor U20369 (N_20369,N_19558,N_19491);
xnor U20370 (N_20370,N_18902,N_18538);
nor U20371 (N_20371,N_18429,N_19989);
nor U20372 (N_20372,N_18496,N_18874);
xor U20373 (N_20373,N_19992,N_18535);
or U20374 (N_20374,N_19736,N_19320);
and U20375 (N_20375,N_18048,N_18058);
nand U20376 (N_20376,N_19844,N_19765);
nor U20377 (N_20377,N_19120,N_19695);
nor U20378 (N_20378,N_19470,N_18268);
or U20379 (N_20379,N_18705,N_19378);
nor U20380 (N_20380,N_18438,N_19011);
xor U20381 (N_20381,N_18066,N_19849);
and U20382 (N_20382,N_19146,N_18144);
or U20383 (N_20383,N_19152,N_19215);
nand U20384 (N_20384,N_18584,N_18794);
xnor U20385 (N_20385,N_18366,N_19596);
nand U20386 (N_20386,N_19778,N_18658);
nand U20387 (N_20387,N_19905,N_18964);
nor U20388 (N_20388,N_19125,N_18290);
nand U20389 (N_20389,N_18613,N_18279);
nand U20390 (N_20390,N_18882,N_19987);
xor U20391 (N_20391,N_18427,N_18341);
xor U20392 (N_20392,N_18788,N_18281);
nor U20393 (N_20393,N_18478,N_19246);
and U20394 (N_20394,N_18340,N_19952);
nor U20395 (N_20395,N_19151,N_19975);
nand U20396 (N_20396,N_19281,N_19266);
or U20397 (N_20397,N_19782,N_19917);
and U20398 (N_20398,N_19880,N_19098);
nand U20399 (N_20399,N_18711,N_18572);
nor U20400 (N_20400,N_18556,N_19836);
nand U20401 (N_20401,N_18164,N_18425);
or U20402 (N_20402,N_19498,N_19365);
nand U20403 (N_20403,N_18839,N_18649);
nor U20404 (N_20404,N_19238,N_18548);
and U20405 (N_20405,N_19995,N_18129);
nor U20406 (N_20406,N_18100,N_18950);
xor U20407 (N_20407,N_19659,N_18814);
nand U20408 (N_20408,N_18944,N_18654);
or U20409 (N_20409,N_18853,N_19317);
xnor U20410 (N_20410,N_18688,N_18651);
and U20411 (N_20411,N_19159,N_18262);
and U20412 (N_20412,N_18001,N_18395);
or U20413 (N_20413,N_19462,N_19933);
xnor U20414 (N_20414,N_18735,N_18579);
nand U20415 (N_20415,N_19180,N_18919);
nor U20416 (N_20416,N_19420,N_18209);
xnor U20417 (N_20417,N_19884,N_19939);
nand U20418 (N_20418,N_19052,N_18529);
nor U20419 (N_20419,N_19089,N_19963);
nor U20420 (N_20420,N_19267,N_19862);
or U20421 (N_20421,N_18137,N_18426);
or U20422 (N_20422,N_19225,N_19247);
and U20423 (N_20423,N_18832,N_19221);
or U20424 (N_20424,N_19047,N_18792);
xnor U20425 (N_20425,N_18301,N_18504);
xor U20426 (N_20426,N_18256,N_19743);
and U20427 (N_20427,N_18114,N_18838);
or U20428 (N_20428,N_19007,N_19807);
xor U20429 (N_20429,N_18289,N_19523);
and U20430 (N_20430,N_18471,N_19459);
xnor U20431 (N_20431,N_18023,N_19106);
xor U20432 (N_20432,N_18476,N_18614);
or U20433 (N_20433,N_19724,N_18232);
xnor U20434 (N_20434,N_18243,N_18987);
or U20435 (N_20435,N_19155,N_18111);
nor U20436 (N_20436,N_18418,N_18779);
nor U20437 (N_20437,N_18060,N_19632);
nand U20438 (N_20438,N_18376,N_19681);
or U20439 (N_20439,N_18422,N_18070);
and U20440 (N_20440,N_19069,N_18764);
nand U20441 (N_20441,N_18752,N_18999);
nand U20442 (N_20442,N_19384,N_18021);
xor U20443 (N_20443,N_19881,N_19730);
xor U20444 (N_20444,N_19352,N_18684);
nand U20445 (N_20445,N_18018,N_18297);
nor U20446 (N_20446,N_18187,N_18074);
xor U20447 (N_20447,N_18713,N_19071);
nor U20448 (N_20448,N_19444,N_19620);
and U20449 (N_20449,N_19864,N_18125);
xor U20450 (N_20450,N_18770,N_18452);
and U20451 (N_20451,N_19876,N_18784);
nor U20452 (N_20452,N_18799,N_18773);
or U20453 (N_20453,N_19676,N_18592);
nand U20454 (N_20454,N_18586,N_19904);
nor U20455 (N_20455,N_18716,N_19437);
nand U20456 (N_20456,N_18454,N_19419);
or U20457 (N_20457,N_18680,N_19291);
and U20458 (N_20458,N_18696,N_18542);
nor U20459 (N_20459,N_18368,N_18672);
xor U20460 (N_20460,N_19985,N_19585);
nand U20461 (N_20461,N_19292,N_18605);
xnor U20462 (N_20462,N_18855,N_18756);
nor U20463 (N_20463,N_19721,N_19702);
xor U20464 (N_20464,N_18630,N_19275);
or U20465 (N_20465,N_19385,N_18122);
and U20466 (N_20466,N_18041,N_18811);
or U20467 (N_20467,N_18181,N_18758);
nor U20468 (N_20468,N_19508,N_18727);
and U20469 (N_20469,N_18570,N_19767);
xnor U20470 (N_20470,N_19354,N_18869);
xor U20471 (N_20471,N_18365,N_18287);
xor U20472 (N_20472,N_19907,N_19056);
nor U20473 (N_20473,N_18920,N_18332);
nand U20474 (N_20474,N_19265,N_19070);
nand U20475 (N_20475,N_19237,N_19979);
xor U20476 (N_20476,N_18189,N_18007);
nor U20477 (N_20477,N_19466,N_18182);
and U20478 (N_20478,N_19166,N_19516);
and U20479 (N_20479,N_18322,N_18765);
and U20480 (N_20480,N_19451,N_18253);
nor U20481 (N_20481,N_18536,N_19603);
nor U20482 (N_20482,N_18837,N_19367);
or U20483 (N_20483,N_19232,N_18936);
or U20484 (N_20484,N_19802,N_19438);
or U20485 (N_20485,N_18473,N_19889);
and U20486 (N_20486,N_19088,N_19097);
nand U20487 (N_20487,N_19991,N_19203);
nor U20488 (N_20488,N_18795,N_19002);
nand U20489 (N_20489,N_18493,N_18169);
and U20490 (N_20490,N_19091,N_18387);
nor U20491 (N_20491,N_19600,N_18098);
or U20492 (N_20492,N_19296,N_19560);
and U20493 (N_20493,N_18264,N_19299);
and U20494 (N_20494,N_19589,N_19217);
nor U20495 (N_20495,N_18555,N_19829);
and U20496 (N_20496,N_19858,N_18890);
nand U20497 (N_20497,N_18304,N_18728);
nor U20498 (N_20498,N_19604,N_19433);
nand U20499 (N_20499,N_19272,N_19117);
nand U20500 (N_20500,N_19183,N_18079);
nor U20501 (N_20501,N_19739,N_18966);
xnor U20502 (N_20502,N_19813,N_18600);
nor U20503 (N_20503,N_18830,N_19328);
nor U20504 (N_20504,N_18195,N_19750);
and U20505 (N_20505,N_19116,N_18188);
nand U20506 (N_20506,N_18135,N_19774);
and U20507 (N_20507,N_19387,N_19468);
and U20508 (N_20508,N_18295,N_18859);
nor U20509 (N_20509,N_18622,N_19629);
xor U20510 (N_20510,N_18545,N_18033);
or U20511 (N_20511,N_19439,N_18650);
nand U20512 (N_20512,N_18375,N_18598);
xor U20513 (N_20513,N_18179,N_18644);
nor U20514 (N_20514,N_18392,N_19169);
and U20515 (N_20515,N_18293,N_18147);
xor U20516 (N_20516,N_19241,N_18055);
and U20517 (N_20517,N_18763,N_19962);
xor U20518 (N_20518,N_18612,N_19707);
and U20519 (N_20519,N_18250,N_19348);
xnor U20520 (N_20520,N_19428,N_18970);
xnor U20521 (N_20521,N_18217,N_18323);
xnor U20522 (N_20522,N_18985,N_18120);
nand U20523 (N_20523,N_18363,N_19551);
xor U20524 (N_20524,N_18908,N_19339);
and U20525 (N_20525,N_19950,N_19700);
or U20526 (N_20526,N_19283,N_18938);
xnor U20527 (N_20527,N_19853,N_19403);
or U20528 (N_20528,N_18775,N_18468);
or U20529 (N_20529,N_18826,N_18534);
nand U20530 (N_20530,N_19960,N_19592);
nand U20531 (N_20531,N_18474,N_19461);
nand U20532 (N_20532,N_19983,N_18930);
nor U20533 (N_20533,N_18237,N_18797);
nor U20534 (N_20534,N_19625,N_19493);
nand U20535 (N_20535,N_18439,N_19030);
xor U20536 (N_20536,N_19276,N_19219);
nor U20537 (N_20537,N_18805,N_19677);
or U20538 (N_20538,N_18870,N_19734);
xnor U20539 (N_20539,N_18962,N_19639);
nand U20540 (N_20540,N_19672,N_19576);
or U20541 (N_20541,N_19478,N_19624);
xnor U20542 (N_20542,N_18769,N_19926);
and U20543 (N_20543,N_18096,N_18888);
or U20544 (N_20544,N_18523,N_19696);
and U20545 (N_20545,N_18210,N_18068);
or U20546 (N_20546,N_19609,N_19389);
or U20547 (N_20547,N_19240,N_18270);
nor U20548 (N_20548,N_18939,N_18721);
xor U20549 (N_20549,N_18747,N_19602);
or U20550 (N_20550,N_18240,N_18034);
nor U20551 (N_20551,N_18266,N_19500);
nand U20552 (N_20552,N_18445,N_19374);
and U20553 (N_20553,N_18710,N_18754);
nand U20554 (N_20554,N_19965,N_19449);
xnor U20555 (N_20555,N_18103,N_19167);
nand U20556 (N_20556,N_19946,N_19956);
nor U20557 (N_20557,N_18868,N_18329);
xor U20558 (N_20558,N_19638,N_19758);
nand U20559 (N_20559,N_18803,N_18912);
xor U20560 (N_20560,N_19447,N_19278);
xor U20561 (N_20561,N_19948,N_19663);
nor U20562 (N_20562,N_19024,N_18723);
or U20563 (N_20563,N_19852,N_19065);
or U20564 (N_20564,N_18337,N_19130);
or U20565 (N_20565,N_19103,N_19158);
and U20566 (N_20566,N_18988,N_19645);
nand U20567 (N_20567,N_19027,N_18532);
xnor U20568 (N_20568,N_19966,N_19549);
and U20569 (N_20569,N_19587,N_19096);
and U20570 (N_20570,N_18871,N_18069);
and U20571 (N_20571,N_18099,N_19008);
xor U20572 (N_20572,N_18554,N_19512);
nor U20573 (N_20573,N_18352,N_18771);
xor U20574 (N_20574,N_19817,N_18559);
nand U20575 (N_20575,N_19235,N_19544);
or U20576 (N_20576,N_18517,N_19176);
nor U20577 (N_20577,N_18748,N_18416);
or U20578 (N_20578,N_19396,N_19655);
nand U20579 (N_20579,N_19206,N_19335);
or U20580 (N_20580,N_18271,N_19255);
xnor U20581 (N_20581,N_18513,N_19997);
or U20582 (N_20582,N_19460,N_19742);
and U20583 (N_20583,N_18591,N_19863);
and U20584 (N_20584,N_19569,N_18433);
and U20585 (N_20585,N_18695,N_18700);
or U20586 (N_20586,N_18744,N_19888);
and U20587 (N_20587,N_18045,N_19550);
and U20588 (N_20588,N_18520,N_19018);
or U20589 (N_20589,N_19105,N_19612);
nand U20590 (N_20590,N_19755,N_19796);
or U20591 (N_20591,N_18325,N_19673);
or U20592 (N_20592,N_18434,N_18778);
or U20593 (N_20593,N_18911,N_18992);
nor U20594 (N_20594,N_19391,N_19131);
and U20595 (N_20595,N_18047,N_19908);
nand U20596 (N_20596,N_18015,N_19537);
xnor U20597 (N_20597,N_18239,N_18244);
nand U20598 (N_20598,N_19072,N_19163);
and U20599 (N_20599,N_18163,N_19340);
or U20600 (N_20600,N_18984,N_18900);
xnor U20601 (N_20601,N_18753,N_19214);
nor U20602 (N_20602,N_18444,N_18978);
xnor U20603 (N_20603,N_19104,N_19434);
xnor U20604 (N_20604,N_18004,N_19416);
nand U20605 (N_20605,N_19492,N_18308);
xor U20606 (N_20606,N_19621,N_19656);
and U20607 (N_20607,N_18374,N_18567);
nor U20608 (N_20608,N_18343,N_18616);
nor U20609 (N_20609,N_18822,N_18646);
and U20610 (N_20610,N_18743,N_18415);
xnor U20611 (N_20611,N_18065,N_18722);
or U20612 (N_20612,N_19794,N_19218);
nor U20613 (N_20613,N_18479,N_18321);
nand U20614 (N_20614,N_19139,N_19514);
or U20615 (N_20615,N_19706,N_19373);
xnor U20616 (N_20616,N_18085,N_19704);
xor U20617 (N_20617,N_19973,N_19094);
nor U20618 (N_20618,N_19309,N_18115);
and U20619 (N_20619,N_18291,N_18669);
and U20620 (N_20620,N_19302,N_18549);
nand U20621 (N_20621,N_19662,N_18335);
xnor U20622 (N_20622,N_18139,N_19711);
and U20623 (N_20623,N_19910,N_19021);
xnor U20624 (N_20624,N_19357,N_19213);
and U20625 (N_20625,N_18121,N_18225);
and U20626 (N_20626,N_18075,N_18153);
and U20627 (N_20627,N_19044,N_18698);
nand U20628 (N_20628,N_18116,N_18732);
nor U20629 (N_20629,N_19744,N_18801);
nand U20630 (N_20630,N_19051,N_18014);
xor U20631 (N_20631,N_18505,N_18032);
and U20632 (N_20632,N_19976,N_19342);
xor U20633 (N_20633,N_18585,N_18807);
or U20634 (N_20634,N_19453,N_18488);
nor U20635 (N_20635,N_19322,N_18982);
and U20636 (N_20636,N_19810,N_18729);
xor U20637 (N_20637,N_19315,N_18627);
nand U20638 (N_20638,N_18958,N_18516);
nand U20639 (N_20639,N_18872,N_18314);
and U20640 (N_20640,N_19323,N_19109);
nand U20641 (N_20641,N_19210,N_19818);
and U20642 (N_20642,N_18350,N_18351);
nand U20643 (N_20643,N_19115,N_18219);
xnor U20644 (N_20644,N_19029,N_18699);
nand U20645 (N_20645,N_18282,N_18907);
nand U20646 (N_20646,N_18198,N_19486);
nand U20647 (N_20647,N_18257,N_19532);
or U20648 (N_20648,N_18697,N_18247);
or U20649 (N_20649,N_18774,N_19536);
and U20650 (N_20650,N_18578,N_18173);
nand U20651 (N_20651,N_19961,N_18277);
and U20652 (N_20652,N_19729,N_19345);
and U20653 (N_20653,N_19972,N_18483);
xor U20654 (N_20654,N_19727,N_18285);
and U20655 (N_20655,N_19943,N_18216);
and U20656 (N_20656,N_19577,N_19891);
nand U20657 (N_20657,N_19463,N_18204);
xnor U20658 (N_20658,N_18850,N_18761);
or U20659 (N_20659,N_18854,N_18410);
and U20660 (N_20660,N_19756,N_18108);
nand U20661 (N_20661,N_18973,N_18123);
or U20662 (N_20662,N_19660,N_19793);
xnor U20663 (N_20663,N_18328,N_19897);
nand U20664 (N_20664,N_18553,N_19040);
nor U20665 (N_20665,N_19776,N_19025);
nor U20666 (N_20666,N_18119,N_18064);
xnor U20667 (N_20667,N_19050,N_19436);
nor U20668 (N_20668,N_19871,N_19124);
xor U20669 (N_20669,N_19136,N_18347);
and U20670 (N_20670,N_18043,N_19429);
nand U20671 (N_20671,N_18674,N_19919);
or U20672 (N_20672,N_19376,N_18562);
and U20673 (N_20673,N_19546,N_19371);
xor U20674 (N_20674,N_19344,N_19407);
xnor U20675 (N_20675,N_18808,N_19775);
xnor U20676 (N_20676,N_18331,N_19909);
and U20677 (N_20677,N_19383,N_18269);
nor U20678 (N_20678,N_18230,N_19261);
xor U20679 (N_20679,N_18720,N_19866);
and U20680 (N_20680,N_18489,N_19048);
and U20681 (N_20681,N_19495,N_18632);
and U20682 (N_20682,N_18979,N_18677);
or U20683 (N_20683,N_18201,N_18543);
xnor U20684 (N_20684,N_19786,N_19932);
nand U20685 (N_20685,N_18935,N_18981);
nand U20686 (N_20686,N_19826,N_18475);
nand U20687 (N_20687,N_18013,N_18682);
or U20688 (N_20688,N_19085,N_19211);
nand U20689 (N_20689,N_18200,N_18254);
nand U20690 (N_20690,N_19398,N_18521);
and U20691 (N_20691,N_19540,N_19784);
nand U20692 (N_20692,N_19735,N_18038);
and U20693 (N_20693,N_18212,N_18218);
and U20694 (N_20694,N_19269,N_18086);
nor U20695 (N_20695,N_19790,N_18884);
or U20696 (N_20696,N_18124,N_18161);
or U20697 (N_20697,N_19738,N_18508);
nor U20698 (N_20698,N_18849,N_19262);
and U20699 (N_20699,N_19277,N_19892);
nor U20700 (N_20700,N_19931,N_19543);
or U20701 (N_20701,N_19584,N_18057);
nand U20702 (N_20702,N_19228,N_18235);
nand U20703 (N_20703,N_19321,N_19883);
and U20704 (N_20704,N_18921,N_18655);
nor U20705 (N_20705,N_18742,N_19608);
nand U20706 (N_20706,N_19140,N_18208);
nor U20707 (N_20707,N_19229,N_19060);
nor U20708 (N_20708,N_18283,N_18741);
nor U20709 (N_20709,N_19279,N_19974);
xnor U20710 (N_20710,N_19316,N_19838);
nor U20711 (N_20711,N_19928,N_18419);
or U20712 (N_20712,N_19686,N_19350);
or U20713 (N_20713,N_19318,N_18851);
nor U20714 (N_20714,N_18265,N_18668);
xnor U20715 (N_20715,N_19581,N_19636);
and U20716 (N_20716,N_18447,N_19333);
or U20717 (N_20717,N_19870,N_18083);
xor U20718 (N_20718,N_18373,N_18192);
nand U20719 (N_20719,N_19627,N_18892);
nand U20720 (N_20720,N_18738,N_18246);
nand U20721 (N_20721,N_19605,N_18816);
or U20722 (N_20722,N_19431,N_18107);
nand U20723 (N_20723,N_19697,N_19308);
nor U20724 (N_20724,N_18848,N_19220);
nand U20725 (N_20725,N_18495,N_19857);
nor U20726 (N_20726,N_19687,N_18384);
and U20727 (N_20727,N_18514,N_19597);
nor U20728 (N_20728,N_18062,N_19304);
and U20729 (N_20729,N_19078,N_18390);
or U20730 (N_20730,N_19095,N_18582);
nand U20731 (N_20731,N_19999,N_19825);
xor U20732 (N_20732,N_19837,N_19347);
or U20733 (N_20733,N_18263,N_18006);
and U20734 (N_20734,N_18046,N_18404);
nor U20735 (N_20735,N_18917,N_18272);
and U20736 (N_20736,N_18608,N_19404);
or U20737 (N_20737,N_18274,N_19855);
nand U20738 (N_20738,N_18563,N_18881);
or U20739 (N_20739,N_19270,N_18642);
or U20740 (N_20740,N_19137,N_18000);
xor U20741 (N_20741,N_19580,N_19530);
nand U20742 (N_20742,N_18737,N_18165);
xor U20743 (N_20743,N_18626,N_19452);
xnor U20744 (N_20744,N_18518,N_19287);
nand U20745 (N_20745,N_18791,N_18238);
or U20746 (N_20746,N_19890,N_19964);
nand U20747 (N_20747,N_18666,N_18914);
nor U20748 (N_20748,N_19469,N_18588);
nand U20749 (N_20749,N_19341,N_18989);
and U20750 (N_20750,N_19923,N_18762);
nand U20751 (N_20751,N_19553,N_18876);
xnor U20752 (N_20752,N_18316,N_18185);
or U20753 (N_20753,N_19869,N_18867);
and U20754 (N_20754,N_18224,N_19101);
or U20755 (N_20755,N_18378,N_19325);
or U20756 (N_20756,N_19033,N_19539);
nor U20757 (N_20757,N_19264,N_19653);
or U20758 (N_20758,N_19053,N_18203);
or U20759 (N_20759,N_18704,N_18909);
nand U20760 (N_20760,N_18507,N_19792);
xnor U20761 (N_20761,N_19517,N_18251);
or U20762 (N_20762,N_18796,N_19019);
nand U20763 (N_20763,N_19154,N_19827);
or U20764 (N_20764,N_19607,N_19188);
nand U20765 (N_20765,N_18029,N_19953);
and U20766 (N_20766,N_19393,N_19861);
and U20767 (N_20767,N_19588,N_18423);
and U20768 (N_20768,N_18991,N_19570);
or U20769 (N_20769,N_18160,N_18360);
or U20770 (N_20770,N_19619,N_19113);
xnor U20771 (N_20771,N_19430,N_18653);
and U20772 (N_20772,N_19868,N_18821);
nand U20773 (N_20773,N_19205,N_19733);
or U20774 (N_20774,N_19005,N_19484);
or U20775 (N_20775,N_19895,N_18446);
xor U20776 (N_20776,N_18072,N_18683);
or U20777 (N_20777,N_19346,N_19994);
and U20778 (N_20778,N_18412,N_19454);
nor U20779 (N_20779,N_18740,N_18497);
and U20780 (N_20780,N_19014,N_18923);
xnor U20781 (N_20781,N_19631,N_19998);
or U20782 (N_20782,N_19310,N_18222);
nand U20783 (N_20783,N_19132,N_18127);
and U20784 (N_20784,N_19654,N_18877);
nor U20785 (N_20785,N_18320,N_18025);
nor U20786 (N_20786,N_18354,N_19258);
and U20787 (N_20787,N_18149,N_18526);
and U20788 (N_20788,N_19643,N_18421);
or U20789 (N_20789,N_19226,N_19878);
xnor U20790 (N_20790,N_19313,N_19835);
and U20791 (N_20791,N_19397,N_19379);
nand U20792 (N_20792,N_18424,N_18951);
nand U20793 (N_20793,N_19039,N_18101);
nand U20794 (N_20794,N_18994,N_18414);
or U20795 (N_20795,N_18383,N_19709);
nor U20796 (N_20796,N_18229,N_18725);
nand U20797 (N_20797,N_18915,N_19187);
and U20798 (N_20798,N_18931,N_19409);
nand U20799 (N_20799,N_18168,N_19759);
or U20800 (N_20800,N_19509,N_19698);
or U20801 (N_20801,N_18942,N_18071);
nand U20802 (N_20802,N_18207,N_18883);
nor U20803 (N_20803,N_18772,N_19118);
nand U20804 (N_20804,N_19763,N_18625);
or U20805 (N_20805,N_18825,N_18528);
nor U20806 (N_20806,N_18952,N_18459);
or U20807 (N_20807,N_18780,N_19395);
or U20808 (N_20808,N_18294,N_19740);
nand U20809 (N_20809,N_18726,N_18515);
or U20810 (N_20810,N_18800,N_18843);
nor U20811 (N_20811,N_18056,N_18407);
or U20812 (N_20812,N_18887,N_19327);
nor U20813 (N_20813,N_18968,N_18925);
and U20814 (N_20814,N_18818,N_19042);
and U20815 (N_20815,N_18118,N_18206);
and U20816 (N_20816,N_18420,N_18389);
nand U20817 (N_20817,N_18059,N_18541);
and U20818 (N_20818,N_18760,N_19903);
nand U20819 (N_20819,N_18215,N_18249);
xnor U20820 (N_20820,N_19332,N_19119);
and U20821 (N_20821,N_19616,N_19314);
nand U20822 (N_20822,N_19023,N_19110);
xor U20823 (N_20823,N_18485,N_18852);
and U20824 (N_20824,N_19087,N_19311);
and U20825 (N_20825,N_18576,N_19324);
nand U20826 (N_20826,N_19503,N_19751);
xor U20827 (N_20827,N_18618,N_19541);
and U20828 (N_20828,N_18467,N_18157);
or U20829 (N_20829,N_18158,N_19586);
nand U20830 (N_20830,N_18460,N_19450);
nand U20831 (N_20831,N_18693,N_18492);
xor U20832 (N_20832,N_19223,N_18998);
xor U20833 (N_20833,N_18706,N_19993);
xor U20834 (N_20834,N_18665,N_18162);
or U20835 (N_20835,N_19850,N_19521);
xor U20836 (N_20836,N_19898,N_18937);
nand U20837 (N_20837,N_18393,N_18671);
xnor U20838 (N_20838,N_18829,N_18709);
or U20839 (N_20839,N_18694,N_18574);
nor U20840 (N_20840,N_18757,N_19212);
xor U20841 (N_20841,N_19899,N_19554);
nor U20842 (N_20842,N_19649,N_19411);
nor U20843 (N_20843,N_18199,N_18776);
nand U20844 (N_20844,N_19502,N_19938);
or U20845 (N_20845,N_19839,N_19102);
and U20846 (N_20846,N_18861,N_19675);
nor U20847 (N_20847,N_19847,N_19073);
or U20848 (N_20848,N_18381,N_19944);
or U20849 (N_20849,N_18623,N_18345);
xnor U20850 (N_20850,N_18319,N_19386);
and U20851 (N_20851,N_18167,N_18918);
xor U20852 (N_20852,N_18502,N_18634);
xnor U20853 (N_20853,N_19860,N_19036);
nand U20854 (N_20854,N_19446,N_18397);
or U20855 (N_20855,N_18802,N_19307);
nand U20856 (N_20856,N_18067,N_19062);
or U20857 (N_20857,N_18879,N_19925);
nand U20858 (N_20858,N_19527,N_18441);
nand U20859 (N_20859,N_19293,N_18842);
or U20860 (N_20860,N_18865,N_19197);
nor U20861 (N_20861,N_18258,N_19723);
or U20862 (N_20862,N_18793,N_19915);
nand U20863 (N_20863,N_19161,N_18159);
nor U20864 (N_20864,N_19661,N_18806);
and U20865 (N_20865,N_19432,N_19650);
and U20866 (N_20866,N_18470,N_19012);
xnor U20867 (N_20867,N_19382,N_18652);
or U20868 (N_20868,N_19474,N_19606);
xnor U20869 (N_20869,N_18090,N_19336);
nand U20870 (N_20870,N_19171,N_19522);
nor U20871 (N_20871,N_18177,N_18451);
nor U20872 (N_20872,N_19170,N_19922);
nand U20873 (N_20873,N_19777,N_18629);
or U20874 (N_20874,N_19824,N_19594);
xor U20875 (N_20875,N_18081,N_19942);
or U20876 (N_20876,N_18708,N_19487);
xor U20877 (N_20877,N_19781,N_18864);
nor U20878 (N_20878,N_18357,N_19305);
or U20879 (N_20879,N_19045,N_18533);
nor U20880 (N_20880,N_19252,N_19286);
and U20881 (N_20881,N_18620,N_18580);
xnor U20882 (N_20882,N_18039,N_19031);
xor U20883 (N_20883,N_19996,N_19061);
nand U20884 (N_20884,N_18336,N_18946);
or U20885 (N_20885,N_18667,N_18477);
nand U20886 (N_20886,N_18755,N_19572);
or U20887 (N_20887,N_18601,N_19360);
or U20888 (N_20888,N_19920,N_19173);
nand U20889 (N_20889,N_19368,N_18356);
xor U20890 (N_20890,N_19245,N_19126);
and U20891 (N_20891,N_18273,N_18589);
and U20892 (N_20892,N_18196,N_18679);
nor U20893 (N_20893,N_19390,N_18016);
or U20894 (N_20894,N_18150,N_18044);
nor U20895 (N_20895,N_19057,N_19593);
xnor U20896 (N_20896,N_18036,N_18333);
and U20897 (N_20897,N_18893,N_18280);
nand U20898 (N_20898,N_19900,N_18002);
and U20899 (N_20899,N_19524,N_18511);
xor U20900 (N_20900,N_18430,N_18590);
nor U20901 (N_20901,N_18027,N_19156);
xor U20902 (N_20902,N_18261,N_19674);
nor U20903 (N_20903,N_19559,N_19141);
xor U20904 (N_20904,N_18678,N_18040);
nand U20905 (N_20905,N_18344,N_18661);
nand U20906 (N_20906,N_19787,N_18012);
and U20907 (N_20907,N_18102,N_19665);
nand U20908 (N_20908,N_19635,N_19823);
nand U20909 (N_20909,N_18833,N_18997);
and U20910 (N_20910,N_18435,N_19749);
xnor U20911 (N_20911,N_18809,N_19157);
or U20912 (N_20912,N_18088,N_19337);
and U20913 (N_20913,N_19854,N_18812);
nand U20914 (N_20914,N_18519,N_19918);
xnor U20915 (N_20915,N_19670,N_19699);
or U20916 (N_20916,N_18443,N_19568);
nor U20917 (N_20917,N_19177,N_19186);
or U20918 (N_20918,N_19761,N_19623);
or U20919 (N_20919,N_19547,N_18245);
nor U20920 (N_20920,N_18836,N_18715);
and U20921 (N_20921,N_18719,N_19666);
xor U20922 (N_20922,N_18094,N_18382);
nand U20923 (N_20923,N_19507,N_19114);
nand U20924 (N_20924,N_19913,N_18170);
xor U20925 (N_20925,N_18491,N_19513);
nand U20926 (N_20926,N_19832,N_18214);
nor U20927 (N_20927,N_18462,N_18091);
xor U20928 (N_20928,N_18768,N_19886);
xor U20929 (N_20929,N_19722,N_18236);
or U20930 (N_20930,N_18457,N_18975);
xnor U20931 (N_20931,N_18172,N_18234);
or U20932 (N_20932,N_19496,N_19160);
and U20933 (N_20933,N_19185,N_18026);
or U20934 (N_20934,N_19615,N_18030);
nor U20935 (N_20935,N_18603,N_19243);
and U20936 (N_20936,N_19425,N_18641);
nor U20937 (N_20937,N_19667,N_18624);
xor U20938 (N_20938,N_19041,N_18621);
nor U20939 (N_20939,N_18063,N_19741);
nor U20940 (N_20940,N_18394,N_18993);
or U20941 (N_20941,N_19427,N_19610);
and U20942 (N_20942,N_19331,N_18428);
and U20943 (N_20943,N_18361,N_18092);
nand U20944 (N_20944,N_19954,N_19971);
nor U20945 (N_20945,N_18205,N_19731);
and U20946 (N_20946,N_18866,N_19190);
or U20947 (N_20947,N_19598,N_19879);
nor U20948 (N_20948,N_19951,N_18844);
and U20949 (N_20949,N_19038,N_19611);
nand U20950 (N_20950,N_19694,N_18140);
xnor U20951 (N_20951,N_19092,N_18636);
nor U20952 (N_20952,N_18583,N_19583);
nand U20953 (N_20953,N_18155,N_19571);
xor U20954 (N_20954,N_19628,N_19482);
xor U20955 (N_20955,N_19481,N_19063);
or U20956 (N_20956,N_19244,N_18330);
nor U20957 (N_20957,N_18132,N_18154);
xnor U20958 (N_20958,N_19112,N_19402);
xnor U20959 (N_20959,N_18288,N_19294);
nor U20960 (N_20960,N_18995,N_18464);
or U20961 (N_20961,N_18905,N_18961);
nand U20962 (N_20962,N_19833,N_18436);
and U20963 (N_20963,N_18499,N_18359);
xor U20964 (N_20964,N_19412,N_18643);
nand U20965 (N_20965,N_18342,N_19937);
nand U20966 (N_20966,N_18334,N_19798);
or U20967 (N_20967,N_18733,N_18494);
or U20968 (N_20968,N_19421,N_18141);
nand U20969 (N_20969,N_19282,N_19253);
nand U20970 (N_20970,N_19715,N_19259);
nor U20971 (N_20971,N_18456,N_18093);
xnor U20972 (N_20972,N_19260,N_18676);
or U20973 (N_20973,N_19529,N_18857);
xor U20974 (N_20974,N_19525,N_19483);
xor U20975 (N_20975,N_19688,N_18530);
and U20976 (N_20976,N_19515,N_18227);
nand U20977 (N_20977,N_19353,N_18346);
nor U20978 (N_20978,N_19528,N_18148);
nor U20979 (N_20979,N_19380,N_18166);
xor U20980 (N_20980,N_18569,N_19712);
and U20981 (N_20981,N_19075,N_18431);
xnor U20982 (N_20982,N_19716,N_19680);
or U20983 (N_20983,N_18786,N_19290);
nor U20984 (N_20984,N_19510,N_18106);
and U20985 (N_20985,N_19646,N_19945);
or U20986 (N_20986,N_19473,N_19800);
xor U20987 (N_20987,N_19303,N_19490);
xnor U20988 (N_20988,N_19424,N_19233);
nand U20989 (N_20989,N_18077,N_19423);
or U20990 (N_20990,N_18152,N_19575);
and U20991 (N_20991,N_18143,N_18399);
nand U20992 (N_20992,N_18440,N_19783);
and U20993 (N_20993,N_18355,N_19288);
xor U20994 (N_20994,N_18176,N_18228);
or U20995 (N_20995,N_18782,N_18823);
xor U20996 (N_20996,N_19013,N_18577);
xor U20997 (N_20997,N_18349,N_19874);
or U20998 (N_20998,N_19475,N_18035);
nand U20999 (N_20999,N_19168,N_19567);
nor U21000 (N_21000,N_18487,N_19414);
xor U21001 (N_21001,N_18955,N_18415);
nor U21002 (N_21002,N_18967,N_19127);
nor U21003 (N_21003,N_19670,N_18677);
xnor U21004 (N_21004,N_19992,N_18910);
and U21005 (N_21005,N_19034,N_19047);
xnor U21006 (N_21006,N_18612,N_19535);
xor U21007 (N_21007,N_19069,N_18007);
or U21008 (N_21008,N_18754,N_18452);
xnor U21009 (N_21009,N_19558,N_18121);
or U21010 (N_21010,N_18135,N_19565);
nor U21011 (N_21011,N_18658,N_18026);
and U21012 (N_21012,N_19244,N_19998);
and U21013 (N_21013,N_19828,N_19039);
or U21014 (N_21014,N_19337,N_19940);
nor U21015 (N_21015,N_19113,N_19126);
nand U21016 (N_21016,N_18585,N_18989);
or U21017 (N_21017,N_19430,N_18863);
or U21018 (N_21018,N_18040,N_18905);
nand U21019 (N_21019,N_19458,N_19517);
or U21020 (N_21020,N_18452,N_19836);
and U21021 (N_21021,N_18784,N_18496);
nand U21022 (N_21022,N_18322,N_19432);
nand U21023 (N_21023,N_18658,N_19766);
nor U21024 (N_21024,N_18296,N_19701);
xnor U21025 (N_21025,N_19617,N_18288);
nor U21026 (N_21026,N_18904,N_18109);
nor U21027 (N_21027,N_19375,N_18455);
nand U21028 (N_21028,N_19394,N_19850);
or U21029 (N_21029,N_18823,N_19093);
nor U21030 (N_21030,N_18831,N_18084);
and U21031 (N_21031,N_19059,N_18657);
or U21032 (N_21032,N_19047,N_19378);
nand U21033 (N_21033,N_18090,N_18367);
and U21034 (N_21034,N_18645,N_19462);
xnor U21035 (N_21035,N_19459,N_18999);
xor U21036 (N_21036,N_19387,N_19258);
xnor U21037 (N_21037,N_19259,N_18381);
xor U21038 (N_21038,N_18101,N_18331);
nor U21039 (N_21039,N_18579,N_19566);
or U21040 (N_21040,N_19879,N_19875);
and U21041 (N_21041,N_19798,N_19012);
or U21042 (N_21042,N_19203,N_19331);
and U21043 (N_21043,N_19324,N_19928);
xnor U21044 (N_21044,N_19902,N_18846);
and U21045 (N_21045,N_18264,N_18298);
xor U21046 (N_21046,N_19932,N_18209);
nand U21047 (N_21047,N_18538,N_19389);
or U21048 (N_21048,N_18405,N_18501);
nor U21049 (N_21049,N_18996,N_18134);
or U21050 (N_21050,N_19553,N_18914);
nor U21051 (N_21051,N_18609,N_18469);
or U21052 (N_21052,N_18129,N_19239);
xor U21053 (N_21053,N_19865,N_18052);
nor U21054 (N_21054,N_19185,N_19923);
xor U21055 (N_21055,N_19945,N_18906);
nor U21056 (N_21056,N_19457,N_18676);
and U21057 (N_21057,N_18019,N_19924);
xor U21058 (N_21058,N_18876,N_18167);
nor U21059 (N_21059,N_18884,N_18455);
and U21060 (N_21060,N_19381,N_19361);
nor U21061 (N_21061,N_19792,N_18590);
or U21062 (N_21062,N_18004,N_19241);
nor U21063 (N_21063,N_19852,N_18562);
or U21064 (N_21064,N_18350,N_18015);
and U21065 (N_21065,N_19258,N_19188);
xnor U21066 (N_21066,N_18639,N_19796);
and U21067 (N_21067,N_19749,N_18045);
or U21068 (N_21068,N_19573,N_18136);
and U21069 (N_21069,N_18984,N_18845);
nand U21070 (N_21070,N_19587,N_19138);
xor U21071 (N_21071,N_18697,N_18950);
and U21072 (N_21072,N_19244,N_18484);
xnor U21073 (N_21073,N_19095,N_19962);
xnor U21074 (N_21074,N_18732,N_19104);
and U21075 (N_21075,N_19676,N_19280);
xor U21076 (N_21076,N_19181,N_19947);
or U21077 (N_21077,N_18816,N_19364);
or U21078 (N_21078,N_18360,N_18836);
nor U21079 (N_21079,N_19255,N_19149);
nor U21080 (N_21080,N_18026,N_19255);
nand U21081 (N_21081,N_19832,N_19907);
xor U21082 (N_21082,N_19002,N_18241);
and U21083 (N_21083,N_18705,N_18830);
or U21084 (N_21084,N_18250,N_18573);
or U21085 (N_21085,N_18744,N_19765);
nor U21086 (N_21086,N_18136,N_18557);
nor U21087 (N_21087,N_19761,N_19441);
nor U21088 (N_21088,N_19661,N_18717);
xor U21089 (N_21089,N_19818,N_19259);
or U21090 (N_21090,N_18261,N_18509);
nor U21091 (N_21091,N_19020,N_18492);
and U21092 (N_21092,N_19203,N_19732);
or U21093 (N_21093,N_19083,N_19551);
nand U21094 (N_21094,N_18055,N_18136);
xnor U21095 (N_21095,N_19796,N_18022);
or U21096 (N_21096,N_19839,N_19946);
nand U21097 (N_21097,N_18187,N_19890);
and U21098 (N_21098,N_18635,N_18828);
nor U21099 (N_21099,N_18640,N_18333);
or U21100 (N_21100,N_19621,N_18812);
or U21101 (N_21101,N_19571,N_19268);
nand U21102 (N_21102,N_18313,N_18851);
xnor U21103 (N_21103,N_18090,N_19055);
and U21104 (N_21104,N_19631,N_19175);
nand U21105 (N_21105,N_19501,N_19893);
nor U21106 (N_21106,N_19255,N_18681);
nand U21107 (N_21107,N_19115,N_19389);
xnor U21108 (N_21108,N_19199,N_19677);
nand U21109 (N_21109,N_18196,N_19179);
xor U21110 (N_21110,N_18937,N_19662);
nand U21111 (N_21111,N_18878,N_18974);
nand U21112 (N_21112,N_18979,N_19809);
xnor U21113 (N_21113,N_18649,N_19501);
xnor U21114 (N_21114,N_18850,N_19610);
and U21115 (N_21115,N_19602,N_18086);
and U21116 (N_21116,N_19258,N_18532);
nor U21117 (N_21117,N_18907,N_19334);
and U21118 (N_21118,N_18598,N_18179);
and U21119 (N_21119,N_19326,N_19315);
nand U21120 (N_21120,N_18632,N_18134);
xnor U21121 (N_21121,N_18393,N_19404);
and U21122 (N_21122,N_18537,N_19254);
nor U21123 (N_21123,N_18982,N_18567);
nand U21124 (N_21124,N_18489,N_18657);
nor U21125 (N_21125,N_19619,N_18457);
nand U21126 (N_21126,N_18519,N_19976);
and U21127 (N_21127,N_18590,N_18272);
and U21128 (N_21128,N_19773,N_19325);
and U21129 (N_21129,N_19447,N_19114);
nor U21130 (N_21130,N_18891,N_19302);
xnor U21131 (N_21131,N_19626,N_19086);
nand U21132 (N_21132,N_19228,N_19893);
and U21133 (N_21133,N_18142,N_18897);
or U21134 (N_21134,N_18698,N_19205);
nand U21135 (N_21135,N_18529,N_18227);
xnor U21136 (N_21136,N_18538,N_19973);
and U21137 (N_21137,N_18666,N_19418);
or U21138 (N_21138,N_19518,N_18794);
nor U21139 (N_21139,N_18619,N_18497);
nand U21140 (N_21140,N_19521,N_19623);
xor U21141 (N_21141,N_18127,N_19947);
or U21142 (N_21142,N_19246,N_18471);
or U21143 (N_21143,N_19523,N_19065);
nor U21144 (N_21144,N_18225,N_19595);
nor U21145 (N_21145,N_18407,N_19879);
nand U21146 (N_21146,N_19143,N_19116);
xor U21147 (N_21147,N_19409,N_18139);
nor U21148 (N_21148,N_19568,N_19499);
or U21149 (N_21149,N_18634,N_18837);
or U21150 (N_21150,N_19621,N_18501);
nand U21151 (N_21151,N_19501,N_18507);
nand U21152 (N_21152,N_19589,N_19031);
nand U21153 (N_21153,N_18377,N_19913);
nor U21154 (N_21154,N_18853,N_19521);
and U21155 (N_21155,N_18823,N_19651);
nand U21156 (N_21156,N_19361,N_18015);
and U21157 (N_21157,N_19954,N_19668);
and U21158 (N_21158,N_18854,N_18820);
or U21159 (N_21159,N_18950,N_18531);
nand U21160 (N_21160,N_18859,N_18694);
and U21161 (N_21161,N_18550,N_18566);
or U21162 (N_21162,N_19924,N_19472);
nand U21163 (N_21163,N_19963,N_18281);
xnor U21164 (N_21164,N_18858,N_19235);
xor U21165 (N_21165,N_19399,N_19002);
nand U21166 (N_21166,N_19732,N_18531);
and U21167 (N_21167,N_19097,N_19246);
or U21168 (N_21168,N_19599,N_18126);
or U21169 (N_21169,N_19558,N_19532);
and U21170 (N_21170,N_18280,N_19025);
and U21171 (N_21171,N_18675,N_18133);
or U21172 (N_21172,N_18333,N_19247);
and U21173 (N_21173,N_19396,N_19157);
or U21174 (N_21174,N_19227,N_19474);
xor U21175 (N_21175,N_18299,N_19783);
nor U21176 (N_21176,N_19119,N_18453);
or U21177 (N_21177,N_19765,N_18963);
or U21178 (N_21178,N_19601,N_18068);
and U21179 (N_21179,N_19959,N_18171);
nor U21180 (N_21180,N_19867,N_19695);
nor U21181 (N_21181,N_18125,N_18916);
xnor U21182 (N_21182,N_18269,N_18185);
or U21183 (N_21183,N_18700,N_18197);
and U21184 (N_21184,N_18021,N_19557);
or U21185 (N_21185,N_19787,N_18070);
xor U21186 (N_21186,N_18823,N_19999);
or U21187 (N_21187,N_18302,N_19193);
and U21188 (N_21188,N_19363,N_19016);
or U21189 (N_21189,N_19575,N_19629);
xnor U21190 (N_21190,N_18407,N_18134);
and U21191 (N_21191,N_18216,N_18182);
and U21192 (N_21192,N_19313,N_19766);
nor U21193 (N_21193,N_19155,N_19505);
or U21194 (N_21194,N_18695,N_18891);
xnor U21195 (N_21195,N_18609,N_19282);
nand U21196 (N_21196,N_18540,N_18996);
xnor U21197 (N_21197,N_19084,N_18713);
and U21198 (N_21198,N_18477,N_18378);
and U21199 (N_21199,N_19060,N_19611);
nand U21200 (N_21200,N_19369,N_19519);
and U21201 (N_21201,N_18108,N_19295);
nand U21202 (N_21202,N_19041,N_19140);
and U21203 (N_21203,N_19822,N_18612);
xor U21204 (N_21204,N_18939,N_19298);
and U21205 (N_21205,N_18622,N_19894);
xor U21206 (N_21206,N_18091,N_18401);
nand U21207 (N_21207,N_19908,N_18823);
xor U21208 (N_21208,N_19491,N_19592);
nand U21209 (N_21209,N_19594,N_18588);
and U21210 (N_21210,N_18410,N_19901);
nand U21211 (N_21211,N_19498,N_19690);
and U21212 (N_21212,N_19218,N_18469);
or U21213 (N_21213,N_18412,N_19959);
or U21214 (N_21214,N_18635,N_18535);
nor U21215 (N_21215,N_19767,N_18598);
xor U21216 (N_21216,N_18534,N_18240);
nand U21217 (N_21217,N_19574,N_18161);
and U21218 (N_21218,N_19259,N_18457);
or U21219 (N_21219,N_18927,N_18719);
nand U21220 (N_21220,N_18110,N_18090);
xnor U21221 (N_21221,N_18864,N_19204);
or U21222 (N_21222,N_19896,N_19789);
nor U21223 (N_21223,N_18780,N_18648);
or U21224 (N_21224,N_19346,N_19805);
and U21225 (N_21225,N_18583,N_19922);
nand U21226 (N_21226,N_19829,N_18126);
and U21227 (N_21227,N_19297,N_19319);
nand U21228 (N_21228,N_18278,N_18415);
or U21229 (N_21229,N_18039,N_18993);
nand U21230 (N_21230,N_19927,N_18542);
and U21231 (N_21231,N_18548,N_18279);
xor U21232 (N_21232,N_18172,N_18629);
nand U21233 (N_21233,N_19993,N_18321);
nand U21234 (N_21234,N_18655,N_19745);
and U21235 (N_21235,N_19867,N_19323);
and U21236 (N_21236,N_19702,N_18123);
nor U21237 (N_21237,N_19142,N_19453);
or U21238 (N_21238,N_18429,N_18213);
xnor U21239 (N_21239,N_19254,N_19916);
and U21240 (N_21240,N_18743,N_19390);
xor U21241 (N_21241,N_18678,N_19776);
or U21242 (N_21242,N_19267,N_18021);
nand U21243 (N_21243,N_19223,N_18623);
nor U21244 (N_21244,N_18791,N_18550);
nor U21245 (N_21245,N_18410,N_18524);
and U21246 (N_21246,N_18721,N_18274);
and U21247 (N_21247,N_18846,N_19559);
and U21248 (N_21248,N_19332,N_19573);
xnor U21249 (N_21249,N_18034,N_19486);
nor U21250 (N_21250,N_18969,N_19790);
and U21251 (N_21251,N_19591,N_19205);
nor U21252 (N_21252,N_18735,N_19281);
xnor U21253 (N_21253,N_18430,N_19854);
nand U21254 (N_21254,N_18249,N_19809);
nor U21255 (N_21255,N_18053,N_18597);
nand U21256 (N_21256,N_18836,N_18202);
or U21257 (N_21257,N_19555,N_19679);
xor U21258 (N_21258,N_19265,N_19601);
nand U21259 (N_21259,N_18550,N_19711);
and U21260 (N_21260,N_18946,N_18691);
or U21261 (N_21261,N_19201,N_19334);
and U21262 (N_21262,N_19250,N_19266);
xor U21263 (N_21263,N_18055,N_18314);
xnor U21264 (N_21264,N_18107,N_18687);
or U21265 (N_21265,N_19869,N_19693);
nand U21266 (N_21266,N_18822,N_19306);
nand U21267 (N_21267,N_18018,N_19111);
and U21268 (N_21268,N_19647,N_19785);
nor U21269 (N_21269,N_18428,N_18543);
and U21270 (N_21270,N_19319,N_19535);
nor U21271 (N_21271,N_19451,N_19692);
or U21272 (N_21272,N_18490,N_19754);
xor U21273 (N_21273,N_18806,N_18295);
nand U21274 (N_21274,N_18302,N_19884);
and U21275 (N_21275,N_19225,N_18536);
or U21276 (N_21276,N_18189,N_19369);
nand U21277 (N_21277,N_18813,N_19335);
or U21278 (N_21278,N_18091,N_19722);
and U21279 (N_21279,N_19687,N_18492);
nand U21280 (N_21280,N_19761,N_18742);
nor U21281 (N_21281,N_18637,N_19222);
nor U21282 (N_21282,N_18815,N_19626);
xnor U21283 (N_21283,N_18910,N_19707);
nand U21284 (N_21284,N_19104,N_18518);
or U21285 (N_21285,N_18663,N_19411);
or U21286 (N_21286,N_18945,N_19763);
nor U21287 (N_21287,N_19014,N_18421);
and U21288 (N_21288,N_18349,N_18811);
or U21289 (N_21289,N_19065,N_18925);
nor U21290 (N_21290,N_19557,N_19834);
and U21291 (N_21291,N_19175,N_18799);
nor U21292 (N_21292,N_18214,N_19429);
or U21293 (N_21293,N_18109,N_18520);
or U21294 (N_21294,N_18330,N_18040);
xor U21295 (N_21295,N_18672,N_19088);
xnor U21296 (N_21296,N_18005,N_19395);
xnor U21297 (N_21297,N_18483,N_18391);
nor U21298 (N_21298,N_18022,N_19807);
nand U21299 (N_21299,N_18834,N_19266);
nand U21300 (N_21300,N_19265,N_19707);
nand U21301 (N_21301,N_18802,N_19905);
or U21302 (N_21302,N_19103,N_18287);
or U21303 (N_21303,N_19267,N_18382);
nor U21304 (N_21304,N_19134,N_19290);
nand U21305 (N_21305,N_19668,N_19583);
xor U21306 (N_21306,N_19168,N_19985);
or U21307 (N_21307,N_18075,N_19818);
nand U21308 (N_21308,N_18288,N_18366);
nand U21309 (N_21309,N_18139,N_19945);
and U21310 (N_21310,N_18875,N_19092);
xor U21311 (N_21311,N_18731,N_19379);
and U21312 (N_21312,N_18844,N_18475);
nand U21313 (N_21313,N_18325,N_18875);
nand U21314 (N_21314,N_19441,N_18242);
xor U21315 (N_21315,N_19367,N_19569);
and U21316 (N_21316,N_18561,N_18835);
and U21317 (N_21317,N_18733,N_19818);
nand U21318 (N_21318,N_19363,N_18925);
xor U21319 (N_21319,N_19452,N_18863);
nand U21320 (N_21320,N_18642,N_18135);
and U21321 (N_21321,N_18014,N_19470);
nor U21322 (N_21322,N_19657,N_19823);
or U21323 (N_21323,N_19300,N_19685);
and U21324 (N_21324,N_19218,N_19644);
and U21325 (N_21325,N_18228,N_19807);
nand U21326 (N_21326,N_18783,N_19401);
or U21327 (N_21327,N_18622,N_19637);
xnor U21328 (N_21328,N_18730,N_19958);
nand U21329 (N_21329,N_18898,N_18093);
or U21330 (N_21330,N_18021,N_18966);
xor U21331 (N_21331,N_18010,N_19322);
and U21332 (N_21332,N_19646,N_18596);
xnor U21333 (N_21333,N_19513,N_18977);
nand U21334 (N_21334,N_18758,N_18416);
xnor U21335 (N_21335,N_18449,N_18392);
or U21336 (N_21336,N_19338,N_19387);
nand U21337 (N_21337,N_18755,N_19058);
nand U21338 (N_21338,N_18876,N_18282);
or U21339 (N_21339,N_18529,N_19224);
xnor U21340 (N_21340,N_18295,N_19061);
or U21341 (N_21341,N_18615,N_18867);
nor U21342 (N_21342,N_19443,N_18206);
nand U21343 (N_21343,N_18072,N_18971);
xnor U21344 (N_21344,N_18842,N_19168);
xnor U21345 (N_21345,N_18558,N_19883);
nand U21346 (N_21346,N_18379,N_19878);
nand U21347 (N_21347,N_18002,N_18237);
xnor U21348 (N_21348,N_18058,N_19640);
xnor U21349 (N_21349,N_18395,N_18997);
xnor U21350 (N_21350,N_19060,N_19382);
and U21351 (N_21351,N_18311,N_19117);
nor U21352 (N_21352,N_19094,N_19802);
nand U21353 (N_21353,N_18802,N_19008);
and U21354 (N_21354,N_19686,N_18150);
nand U21355 (N_21355,N_18793,N_19861);
or U21356 (N_21356,N_19721,N_18613);
xnor U21357 (N_21357,N_18668,N_18941);
nor U21358 (N_21358,N_18960,N_18173);
or U21359 (N_21359,N_18637,N_18531);
nor U21360 (N_21360,N_18535,N_19354);
nand U21361 (N_21361,N_18139,N_19962);
and U21362 (N_21362,N_18368,N_19123);
and U21363 (N_21363,N_19024,N_19808);
or U21364 (N_21364,N_19935,N_19613);
nand U21365 (N_21365,N_19202,N_18675);
nand U21366 (N_21366,N_19117,N_18709);
nand U21367 (N_21367,N_19131,N_19666);
or U21368 (N_21368,N_19559,N_18191);
or U21369 (N_21369,N_19356,N_18972);
xnor U21370 (N_21370,N_19988,N_19538);
xnor U21371 (N_21371,N_19798,N_19991);
xor U21372 (N_21372,N_19646,N_19890);
nor U21373 (N_21373,N_19020,N_19556);
xnor U21374 (N_21374,N_18864,N_18870);
nand U21375 (N_21375,N_19812,N_19149);
nor U21376 (N_21376,N_18942,N_18902);
nor U21377 (N_21377,N_19794,N_19297);
xor U21378 (N_21378,N_19122,N_18962);
and U21379 (N_21379,N_18512,N_19633);
xor U21380 (N_21380,N_18241,N_18606);
and U21381 (N_21381,N_19198,N_18853);
and U21382 (N_21382,N_19217,N_18981);
xor U21383 (N_21383,N_19786,N_19236);
xor U21384 (N_21384,N_19424,N_18080);
xnor U21385 (N_21385,N_19128,N_19224);
or U21386 (N_21386,N_18202,N_18190);
xor U21387 (N_21387,N_18058,N_18180);
xor U21388 (N_21388,N_19734,N_18192);
nand U21389 (N_21389,N_19867,N_18865);
nor U21390 (N_21390,N_19177,N_19385);
and U21391 (N_21391,N_19511,N_18502);
xor U21392 (N_21392,N_18464,N_19866);
nand U21393 (N_21393,N_19981,N_18052);
nand U21394 (N_21394,N_19238,N_18652);
nand U21395 (N_21395,N_19353,N_18659);
nand U21396 (N_21396,N_19731,N_18705);
nand U21397 (N_21397,N_19185,N_18391);
nand U21398 (N_21398,N_18108,N_19227);
nor U21399 (N_21399,N_18603,N_19762);
nor U21400 (N_21400,N_18195,N_19745);
xor U21401 (N_21401,N_18256,N_19629);
or U21402 (N_21402,N_18244,N_19188);
nand U21403 (N_21403,N_18838,N_19688);
nor U21404 (N_21404,N_18912,N_18433);
and U21405 (N_21405,N_19781,N_19840);
xnor U21406 (N_21406,N_18425,N_18535);
nor U21407 (N_21407,N_19341,N_19005);
nor U21408 (N_21408,N_19944,N_19143);
and U21409 (N_21409,N_18002,N_19745);
nand U21410 (N_21410,N_18349,N_19626);
or U21411 (N_21411,N_19449,N_19291);
and U21412 (N_21412,N_19651,N_19327);
nand U21413 (N_21413,N_18218,N_18859);
nor U21414 (N_21414,N_18041,N_18326);
and U21415 (N_21415,N_18069,N_18120);
and U21416 (N_21416,N_19463,N_19334);
or U21417 (N_21417,N_19745,N_19750);
or U21418 (N_21418,N_19978,N_18083);
nor U21419 (N_21419,N_18196,N_18728);
nor U21420 (N_21420,N_18779,N_18424);
nand U21421 (N_21421,N_19164,N_18856);
or U21422 (N_21422,N_19729,N_18428);
or U21423 (N_21423,N_19053,N_18483);
xor U21424 (N_21424,N_18894,N_19657);
xnor U21425 (N_21425,N_18222,N_18997);
nor U21426 (N_21426,N_18628,N_19216);
or U21427 (N_21427,N_18863,N_18667);
nand U21428 (N_21428,N_18620,N_18009);
xor U21429 (N_21429,N_18923,N_18671);
nor U21430 (N_21430,N_18710,N_19788);
or U21431 (N_21431,N_19368,N_18586);
xnor U21432 (N_21432,N_18011,N_19110);
or U21433 (N_21433,N_18945,N_19774);
xnor U21434 (N_21434,N_18946,N_19376);
nor U21435 (N_21435,N_19452,N_19032);
nand U21436 (N_21436,N_18497,N_19897);
nand U21437 (N_21437,N_19668,N_18495);
nor U21438 (N_21438,N_18587,N_18367);
nand U21439 (N_21439,N_18650,N_18027);
and U21440 (N_21440,N_18682,N_18272);
or U21441 (N_21441,N_19455,N_19483);
and U21442 (N_21442,N_18539,N_19720);
xor U21443 (N_21443,N_19595,N_19676);
or U21444 (N_21444,N_18579,N_18503);
nand U21445 (N_21445,N_19532,N_19432);
xor U21446 (N_21446,N_19379,N_18734);
nand U21447 (N_21447,N_18180,N_19309);
xor U21448 (N_21448,N_18654,N_19386);
and U21449 (N_21449,N_19468,N_19593);
or U21450 (N_21450,N_19198,N_19560);
or U21451 (N_21451,N_18956,N_19248);
xor U21452 (N_21452,N_19863,N_18284);
or U21453 (N_21453,N_19122,N_19733);
nor U21454 (N_21454,N_18085,N_19807);
xor U21455 (N_21455,N_19702,N_19227);
xnor U21456 (N_21456,N_19722,N_19542);
and U21457 (N_21457,N_18758,N_19823);
xnor U21458 (N_21458,N_19078,N_18254);
and U21459 (N_21459,N_19648,N_18434);
and U21460 (N_21460,N_18685,N_18844);
nor U21461 (N_21461,N_19552,N_19592);
or U21462 (N_21462,N_18409,N_19827);
nor U21463 (N_21463,N_19910,N_19963);
or U21464 (N_21464,N_18579,N_19084);
or U21465 (N_21465,N_18778,N_19957);
nor U21466 (N_21466,N_18811,N_18197);
or U21467 (N_21467,N_19327,N_18361);
nor U21468 (N_21468,N_18886,N_18940);
nand U21469 (N_21469,N_18462,N_19017);
nor U21470 (N_21470,N_18055,N_18722);
nand U21471 (N_21471,N_18123,N_18883);
and U21472 (N_21472,N_18627,N_19515);
or U21473 (N_21473,N_19209,N_19288);
xor U21474 (N_21474,N_18733,N_19952);
or U21475 (N_21475,N_18452,N_18588);
or U21476 (N_21476,N_19179,N_18094);
nor U21477 (N_21477,N_18026,N_18235);
nand U21478 (N_21478,N_19603,N_19244);
nor U21479 (N_21479,N_18359,N_19016);
xnor U21480 (N_21480,N_18786,N_19571);
and U21481 (N_21481,N_18952,N_19955);
or U21482 (N_21482,N_19087,N_19880);
nor U21483 (N_21483,N_18945,N_18193);
xnor U21484 (N_21484,N_19897,N_18075);
nand U21485 (N_21485,N_19365,N_18527);
xor U21486 (N_21486,N_19198,N_18382);
nor U21487 (N_21487,N_18854,N_18554);
nor U21488 (N_21488,N_18229,N_19785);
nand U21489 (N_21489,N_18757,N_18297);
xnor U21490 (N_21490,N_19516,N_18275);
nor U21491 (N_21491,N_19806,N_19773);
nor U21492 (N_21492,N_18760,N_19886);
or U21493 (N_21493,N_18389,N_18415);
nand U21494 (N_21494,N_18920,N_19098);
xnor U21495 (N_21495,N_18009,N_18893);
xnor U21496 (N_21496,N_18270,N_18968);
or U21497 (N_21497,N_18487,N_18928);
nor U21498 (N_21498,N_19145,N_18368);
and U21499 (N_21499,N_19197,N_18266);
and U21500 (N_21500,N_18074,N_18248);
nor U21501 (N_21501,N_19576,N_19151);
nor U21502 (N_21502,N_19997,N_18749);
nor U21503 (N_21503,N_18778,N_19442);
xor U21504 (N_21504,N_18430,N_18352);
nand U21505 (N_21505,N_19326,N_18341);
xnor U21506 (N_21506,N_19917,N_18372);
nand U21507 (N_21507,N_18216,N_19053);
or U21508 (N_21508,N_19186,N_19693);
xor U21509 (N_21509,N_19211,N_18387);
nor U21510 (N_21510,N_19587,N_18546);
and U21511 (N_21511,N_18396,N_18827);
xnor U21512 (N_21512,N_18981,N_19894);
or U21513 (N_21513,N_19414,N_18992);
nand U21514 (N_21514,N_18899,N_19905);
and U21515 (N_21515,N_18407,N_19511);
and U21516 (N_21516,N_19642,N_18208);
nand U21517 (N_21517,N_18277,N_19878);
nor U21518 (N_21518,N_18710,N_18187);
nand U21519 (N_21519,N_19130,N_19235);
and U21520 (N_21520,N_19708,N_19119);
nand U21521 (N_21521,N_19615,N_18939);
nor U21522 (N_21522,N_19232,N_19275);
nand U21523 (N_21523,N_19797,N_19175);
nand U21524 (N_21524,N_19542,N_19515);
nand U21525 (N_21525,N_19745,N_18900);
or U21526 (N_21526,N_19255,N_18169);
nor U21527 (N_21527,N_19797,N_18160);
and U21528 (N_21528,N_18321,N_18456);
nor U21529 (N_21529,N_18431,N_18582);
and U21530 (N_21530,N_18928,N_19847);
and U21531 (N_21531,N_18261,N_18391);
or U21532 (N_21532,N_19385,N_18845);
or U21533 (N_21533,N_19523,N_18309);
nor U21534 (N_21534,N_18266,N_18614);
and U21535 (N_21535,N_18631,N_19398);
nor U21536 (N_21536,N_19610,N_18599);
xor U21537 (N_21537,N_19901,N_18020);
or U21538 (N_21538,N_19972,N_18595);
nand U21539 (N_21539,N_18497,N_19926);
and U21540 (N_21540,N_19868,N_18427);
and U21541 (N_21541,N_19931,N_19785);
nor U21542 (N_21542,N_19884,N_18632);
nor U21543 (N_21543,N_19566,N_19203);
xor U21544 (N_21544,N_18041,N_18779);
and U21545 (N_21545,N_19969,N_19893);
and U21546 (N_21546,N_18198,N_18996);
nor U21547 (N_21547,N_18556,N_18958);
and U21548 (N_21548,N_18006,N_18812);
nor U21549 (N_21549,N_19239,N_18746);
nor U21550 (N_21550,N_18825,N_18193);
and U21551 (N_21551,N_19529,N_19014);
and U21552 (N_21552,N_18019,N_19197);
xnor U21553 (N_21553,N_18686,N_18976);
nand U21554 (N_21554,N_19508,N_19281);
nand U21555 (N_21555,N_18125,N_18054);
and U21556 (N_21556,N_19259,N_19883);
nand U21557 (N_21557,N_19469,N_18657);
xor U21558 (N_21558,N_18422,N_18215);
nor U21559 (N_21559,N_18707,N_18255);
nand U21560 (N_21560,N_18594,N_19756);
xnor U21561 (N_21561,N_18203,N_19670);
xnor U21562 (N_21562,N_18211,N_18072);
or U21563 (N_21563,N_18277,N_18167);
nand U21564 (N_21564,N_19594,N_19702);
and U21565 (N_21565,N_19252,N_18110);
nor U21566 (N_21566,N_19556,N_19196);
nand U21567 (N_21567,N_18517,N_18904);
and U21568 (N_21568,N_18213,N_18498);
nor U21569 (N_21569,N_18510,N_19206);
nand U21570 (N_21570,N_18449,N_19527);
or U21571 (N_21571,N_19749,N_18717);
or U21572 (N_21572,N_19925,N_19534);
or U21573 (N_21573,N_19449,N_18760);
or U21574 (N_21574,N_18696,N_19893);
or U21575 (N_21575,N_18380,N_19630);
and U21576 (N_21576,N_18917,N_18223);
or U21577 (N_21577,N_19627,N_18832);
and U21578 (N_21578,N_18940,N_19530);
nor U21579 (N_21579,N_18690,N_18308);
or U21580 (N_21580,N_19709,N_18969);
nor U21581 (N_21581,N_19492,N_19608);
or U21582 (N_21582,N_18836,N_18916);
or U21583 (N_21583,N_18546,N_19196);
nand U21584 (N_21584,N_19040,N_18440);
and U21585 (N_21585,N_19667,N_19935);
nor U21586 (N_21586,N_19925,N_19185);
nor U21587 (N_21587,N_18570,N_19157);
xor U21588 (N_21588,N_18525,N_18137);
nand U21589 (N_21589,N_18308,N_18036);
nor U21590 (N_21590,N_19105,N_19855);
nor U21591 (N_21591,N_18203,N_19622);
and U21592 (N_21592,N_19894,N_19953);
xnor U21593 (N_21593,N_19921,N_18352);
and U21594 (N_21594,N_19175,N_18598);
and U21595 (N_21595,N_19956,N_19113);
or U21596 (N_21596,N_19401,N_19093);
nor U21597 (N_21597,N_18598,N_19612);
nor U21598 (N_21598,N_19980,N_18969);
and U21599 (N_21599,N_18862,N_18056);
or U21600 (N_21600,N_19363,N_19356);
nand U21601 (N_21601,N_18878,N_19628);
nor U21602 (N_21602,N_19231,N_19338);
xnor U21603 (N_21603,N_19981,N_19545);
nand U21604 (N_21604,N_18141,N_18830);
xnor U21605 (N_21605,N_18300,N_18981);
nand U21606 (N_21606,N_19091,N_18247);
nand U21607 (N_21607,N_19754,N_19931);
and U21608 (N_21608,N_18098,N_18092);
or U21609 (N_21609,N_18259,N_18848);
xor U21610 (N_21610,N_19279,N_19474);
xnor U21611 (N_21611,N_19027,N_19919);
xor U21612 (N_21612,N_19183,N_19155);
or U21613 (N_21613,N_19909,N_18585);
xnor U21614 (N_21614,N_18686,N_19568);
and U21615 (N_21615,N_19500,N_19819);
nand U21616 (N_21616,N_18099,N_19108);
and U21617 (N_21617,N_19276,N_19097);
nor U21618 (N_21618,N_19535,N_18724);
nor U21619 (N_21619,N_18879,N_18291);
and U21620 (N_21620,N_18029,N_18455);
xnor U21621 (N_21621,N_19190,N_18602);
nand U21622 (N_21622,N_19206,N_18429);
and U21623 (N_21623,N_18948,N_19313);
xnor U21624 (N_21624,N_19902,N_19844);
or U21625 (N_21625,N_18457,N_19527);
or U21626 (N_21626,N_19521,N_18532);
and U21627 (N_21627,N_19532,N_19381);
or U21628 (N_21628,N_19342,N_18237);
xor U21629 (N_21629,N_18637,N_18788);
and U21630 (N_21630,N_19925,N_19948);
and U21631 (N_21631,N_18560,N_19659);
xnor U21632 (N_21632,N_18761,N_19683);
and U21633 (N_21633,N_18470,N_18165);
nand U21634 (N_21634,N_18116,N_19563);
or U21635 (N_21635,N_18134,N_18116);
nor U21636 (N_21636,N_18411,N_18511);
or U21637 (N_21637,N_19029,N_19739);
and U21638 (N_21638,N_19213,N_18864);
nor U21639 (N_21639,N_18218,N_18101);
nor U21640 (N_21640,N_18044,N_18408);
xnor U21641 (N_21641,N_19691,N_18291);
and U21642 (N_21642,N_18850,N_18743);
or U21643 (N_21643,N_19927,N_19468);
and U21644 (N_21644,N_18872,N_19735);
and U21645 (N_21645,N_18437,N_18056);
nor U21646 (N_21646,N_19834,N_18700);
nand U21647 (N_21647,N_18969,N_18420);
nor U21648 (N_21648,N_19761,N_18321);
nor U21649 (N_21649,N_19929,N_19235);
nor U21650 (N_21650,N_18852,N_18486);
xor U21651 (N_21651,N_18705,N_19837);
or U21652 (N_21652,N_19544,N_19231);
xor U21653 (N_21653,N_18232,N_18767);
nor U21654 (N_21654,N_19020,N_19636);
xor U21655 (N_21655,N_18489,N_19049);
nand U21656 (N_21656,N_18291,N_18679);
and U21657 (N_21657,N_19581,N_18171);
xor U21658 (N_21658,N_19137,N_18251);
nand U21659 (N_21659,N_19512,N_19392);
and U21660 (N_21660,N_18271,N_19653);
xnor U21661 (N_21661,N_19938,N_18410);
nand U21662 (N_21662,N_18685,N_18102);
or U21663 (N_21663,N_18488,N_18993);
xnor U21664 (N_21664,N_18799,N_19525);
nand U21665 (N_21665,N_19882,N_18331);
nand U21666 (N_21666,N_19652,N_18102);
nor U21667 (N_21667,N_18394,N_18139);
nand U21668 (N_21668,N_18777,N_18207);
and U21669 (N_21669,N_18688,N_19790);
nor U21670 (N_21670,N_19962,N_19823);
nor U21671 (N_21671,N_19152,N_18227);
and U21672 (N_21672,N_18092,N_18731);
nand U21673 (N_21673,N_19630,N_19402);
or U21674 (N_21674,N_19937,N_18121);
nand U21675 (N_21675,N_18357,N_19387);
nor U21676 (N_21676,N_19994,N_19666);
nor U21677 (N_21677,N_19885,N_18235);
nor U21678 (N_21678,N_19619,N_19361);
nor U21679 (N_21679,N_19107,N_18203);
or U21680 (N_21680,N_18660,N_18349);
and U21681 (N_21681,N_19202,N_18381);
nand U21682 (N_21682,N_19565,N_18559);
xor U21683 (N_21683,N_19062,N_19649);
and U21684 (N_21684,N_18455,N_18331);
and U21685 (N_21685,N_18880,N_19872);
and U21686 (N_21686,N_18852,N_18253);
or U21687 (N_21687,N_19857,N_18635);
and U21688 (N_21688,N_18946,N_18114);
and U21689 (N_21689,N_18431,N_18109);
and U21690 (N_21690,N_19863,N_18909);
nand U21691 (N_21691,N_18999,N_19340);
nand U21692 (N_21692,N_19466,N_18000);
xnor U21693 (N_21693,N_19403,N_18927);
and U21694 (N_21694,N_19693,N_19260);
nand U21695 (N_21695,N_19003,N_19376);
and U21696 (N_21696,N_19738,N_19848);
nor U21697 (N_21697,N_18683,N_19990);
nand U21698 (N_21698,N_18142,N_18674);
and U21699 (N_21699,N_18446,N_18405);
xnor U21700 (N_21700,N_18920,N_19489);
nand U21701 (N_21701,N_18405,N_19198);
nor U21702 (N_21702,N_19257,N_18996);
xor U21703 (N_21703,N_18543,N_19049);
xor U21704 (N_21704,N_18280,N_18247);
nand U21705 (N_21705,N_19064,N_19148);
nor U21706 (N_21706,N_19733,N_18394);
nand U21707 (N_21707,N_18595,N_18913);
xnor U21708 (N_21708,N_18308,N_18540);
xor U21709 (N_21709,N_18561,N_18640);
nor U21710 (N_21710,N_19670,N_19942);
nor U21711 (N_21711,N_18386,N_18170);
nand U21712 (N_21712,N_18657,N_19933);
nand U21713 (N_21713,N_18591,N_18347);
nor U21714 (N_21714,N_19626,N_18607);
xor U21715 (N_21715,N_19739,N_19563);
nor U21716 (N_21716,N_19710,N_19495);
or U21717 (N_21717,N_18168,N_18976);
or U21718 (N_21718,N_18790,N_18977);
nand U21719 (N_21719,N_19577,N_19534);
xnor U21720 (N_21720,N_19169,N_19193);
nand U21721 (N_21721,N_18433,N_19533);
nor U21722 (N_21722,N_19373,N_19063);
nand U21723 (N_21723,N_19078,N_19538);
and U21724 (N_21724,N_19759,N_19294);
xor U21725 (N_21725,N_18195,N_19280);
or U21726 (N_21726,N_19086,N_18367);
and U21727 (N_21727,N_18548,N_18736);
nor U21728 (N_21728,N_19456,N_18546);
and U21729 (N_21729,N_18161,N_18882);
and U21730 (N_21730,N_19526,N_18261);
nor U21731 (N_21731,N_19022,N_19163);
and U21732 (N_21732,N_18267,N_18605);
nand U21733 (N_21733,N_18262,N_18946);
xnor U21734 (N_21734,N_19065,N_18943);
and U21735 (N_21735,N_18758,N_19087);
nor U21736 (N_21736,N_19671,N_18886);
xor U21737 (N_21737,N_19639,N_19320);
and U21738 (N_21738,N_19620,N_19567);
xnor U21739 (N_21739,N_19418,N_18497);
xor U21740 (N_21740,N_18179,N_18863);
or U21741 (N_21741,N_18302,N_18297);
nor U21742 (N_21742,N_18095,N_19353);
nand U21743 (N_21743,N_19759,N_18208);
nand U21744 (N_21744,N_18989,N_18318);
xor U21745 (N_21745,N_18635,N_19797);
nand U21746 (N_21746,N_18560,N_19883);
or U21747 (N_21747,N_19837,N_19412);
or U21748 (N_21748,N_19179,N_18897);
and U21749 (N_21749,N_18056,N_18436);
nand U21750 (N_21750,N_18920,N_18867);
and U21751 (N_21751,N_19003,N_18657);
nand U21752 (N_21752,N_18200,N_18264);
xnor U21753 (N_21753,N_18094,N_19048);
and U21754 (N_21754,N_19901,N_19674);
nor U21755 (N_21755,N_18635,N_18188);
and U21756 (N_21756,N_19663,N_19684);
or U21757 (N_21757,N_19274,N_19584);
xnor U21758 (N_21758,N_18764,N_18301);
and U21759 (N_21759,N_18906,N_18265);
nor U21760 (N_21760,N_18837,N_19281);
nand U21761 (N_21761,N_18877,N_19472);
xor U21762 (N_21762,N_18310,N_19748);
xnor U21763 (N_21763,N_18611,N_18884);
nand U21764 (N_21764,N_18030,N_19901);
or U21765 (N_21765,N_18857,N_19071);
nor U21766 (N_21766,N_18697,N_18168);
nand U21767 (N_21767,N_19132,N_19147);
or U21768 (N_21768,N_18205,N_19985);
nor U21769 (N_21769,N_19518,N_19333);
and U21770 (N_21770,N_19363,N_19522);
xnor U21771 (N_21771,N_18995,N_18507);
xor U21772 (N_21772,N_19647,N_19359);
or U21773 (N_21773,N_18979,N_19845);
and U21774 (N_21774,N_18250,N_18230);
xnor U21775 (N_21775,N_18180,N_18733);
or U21776 (N_21776,N_18247,N_19475);
nor U21777 (N_21777,N_18027,N_18627);
and U21778 (N_21778,N_19465,N_19180);
and U21779 (N_21779,N_19197,N_18938);
xnor U21780 (N_21780,N_18934,N_18560);
xor U21781 (N_21781,N_18738,N_19204);
xnor U21782 (N_21782,N_19758,N_19556);
or U21783 (N_21783,N_19531,N_19201);
and U21784 (N_21784,N_19019,N_19272);
nand U21785 (N_21785,N_19583,N_19406);
xnor U21786 (N_21786,N_19312,N_18078);
or U21787 (N_21787,N_18540,N_19002);
nor U21788 (N_21788,N_18951,N_19359);
or U21789 (N_21789,N_19867,N_19582);
nand U21790 (N_21790,N_19955,N_18620);
or U21791 (N_21791,N_19212,N_18540);
or U21792 (N_21792,N_18109,N_18480);
nor U21793 (N_21793,N_19101,N_18281);
xnor U21794 (N_21794,N_18049,N_18749);
and U21795 (N_21795,N_19116,N_18136);
nand U21796 (N_21796,N_18856,N_18665);
nor U21797 (N_21797,N_19135,N_19273);
and U21798 (N_21798,N_19754,N_18635);
nand U21799 (N_21799,N_19850,N_18636);
xor U21800 (N_21800,N_19095,N_19206);
and U21801 (N_21801,N_19493,N_19032);
and U21802 (N_21802,N_18617,N_18351);
xnor U21803 (N_21803,N_19814,N_18847);
and U21804 (N_21804,N_19992,N_19715);
and U21805 (N_21805,N_19583,N_18110);
nor U21806 (N_21806,N_18651,N_18806);
and U21807 (N_21807,N_18098,N_18559);
xnor U21808 (N_21808,N_19695,N_18354);
or U21809 (N_21809,N_19910,N_18230);
nand U21810 (N_21810,N_18754,N_19768);
nor U21811 (N_21811,N_18050,N_19572);
xnor U21812 (N_21812,N_18849,N_18954);
or U21813 (N_21813,N_18143,N_18621);
nand U21814 (N_21814,N_18809,N_19216);
and U21815 (N_21815,N_18402,N_18679);
nor U21816 (N_21816,N_18741,N_18795);
xor U21817 (N_21817,N_18425,N_18594);
xnor U21818 (N_21818,N_18044,N_19775);
or U21819 (N_21819,N_18618,N_19024);
nor U21820 (N_21820,N_19424,N_19608);
nand U21821 (N_21821,N_19292,N_19591);
xor U21822 (N_21822,N_18603,N_18091);
nor U21823 (N_21823,N_19807,N_19394);
nor U21824 (N_21824,N_19475,N_19943);
xnor U21825 (N_21825,N_19298,N_18694);
nor U21826 (N_21826,N_19534,N_18074);
nand U21827 (N_21827,N_19655,N_18874);
xor U21828 (N_21828,N_18334,N_18081);
and U21829 (N_21829,N_18607,N_19349);
nor U21830 (N_21830,N_19333,N_18378);
and U21831 (N_21831,N_18467,N_18676);
xnor U21832 (N_21832,N_18774,N_19610);
nand U21833 (N_21833,N_18653,N_19954);
nor U21834 (N_21834,N_18815,N_19555);
or U21835 (N_21835,N_19242,N_19792);
xnor U21836 (N_21836,N_19170,N_18122);
or U21837 (N_21837,N_18923,N_19427);
nand U21838 (N_21838,N_19251,N_18486);
nand U21839 (N_21839,N_18202,N_19661);
nand U21840 (N_21840,N_19032,N_18549);
xor U21841 (N_21841,N_18512,N_19789);
nand U21842 (N_21842,N_18357,N_19752);
xor U21843 (N_21843,N_18961,N_19496);
nand U21844 (N_21844,N_19597,N_18092);
and U21845 (N_21845,N_19540,N_19586);
or U21846 (N_21846,N_18417,N_18922);
or U21847 (N_21847,N_18857,N_19647);
nor U21848 (N_21848,N_19222,N_18844);
nand U21849 (N_21849,N_18893,N_19559);
nor U21850 (N_21850,N_19637,N_19419);
nand U21851 (N_21851,N_19862,N_18312);
nand U21852 (N_21852,N_19177,N_19163);
nor U21853 (N_21853,N_19133,N_18773);
nand U21854 (N_21854,N_18766,N_18115);
nand U21855 (N_21855,N_19543,N_19425);
nand U21856 (N_21856,N_18614,N_18360);
nor U21857 (N_21857,N_18696,N_19035);
or U21858 (N_21858,N_18724,N_19160);
or U21859 (N_21859,N_18274,N_18800);
xnor U21860 (N_21860,N_18076,N_19072);
xnor U21861 (N_21861,N_19694,N_18053);
xor U21862 (N_21862,N_19405,N_19089);
and U21863 (N_21863,N_19511,N_18911);
nand U21864 (N_21864,N_19989,N_19277);
and U21865 (N_21865,N_18823,N_19284);
and U21866 (N_21866,N_18081,N_19856);
nor U21867 (N_21867,N_18925,N_19187);
and U21868 (N_21868,N_19453,N_19513);
xnor U21869 (N_21869,N_18241,N_18435);
nor U21870 (N_21870,N_18445,N_18385);
xnor U21871 (N_21871,N_18129,N_18191);
nor U21872 (N_21872,N_18033,N_19288);
nor U21873 (N_21873,N_19471,N_18588);
and U21874 (N_21874,N_18353,N_18289);
nor U21875 (N_21875,N_18875,N_18960);
or U21876 (N_21876,N_19832,N_19723);
nor U21877 (N_21877,N_19989,N_18083);
or U21878 (N_21878,N_19786,N_19934);
xnor U21879 (N_21879,N_18246,N_18397);
nor U21880 (N_21880,N_18531,N_19459);
nand U21881 (N_21881,N_19353,N_19034);
xnor U21882 (N_21882,N_19423,N_18416);
or U21883 (N_21883,N_19233,N_18918);
or U21884 (N_21884,N_18146,N_19482);
nand U21885 (N_21885,N_18061,N_18380);
nand U21886 (N_21886,N_19762,N_18156);
and U21887 (N_21887,N_19838,N_18429);
and U21888 (N_21888,N_18548,N_18780);
and U21889 (N_21889,N_19347,N_19627);
xnor U21890 (N_21890,N_18014,N_19006);
nand U21891 (N_21891,N_19177,N_19692);
nand U21892 (N_21892,N_18975,N_19300);
nor U21893 (N_21893,N_19570,N_19413);
or U21894 (N_21894,N_19611,N_18947);
nand U21895 (N_21895,N_18269,N_18178);
or U21896 (N_21896,N_18444,N_18148);
nand U21897 (N_21897,N_18567,N_19154);
and U21898 (N_21898,N_19526,N_18125);
nor U21899 (N_21899,N_18059,N_19197);
xor U21900 (N_21900,N_19528,N_19941);
and U21901 (N_21901,N_18963,N_18856);
or U21902 (N_21902,N_19249,N_18867);
nor U21903 (N_21903,N_18474,N_19074);
or U21904 (N_21904,N_19945,N_19749);
xor U21905 (N_21905,N_19628,N_19309);
or U21906 (N_21906,N_19275,N_19144);
or U21907 (N_21907,N_19372,N_18281);
nor U21908 (N_21908,N_18473,N_19190);
xnor U21909 (N_21909,N_19176,N_19575);
or U21910 (N_21910,N_18160,N_19545);
nand U21911 (N_21911,N_18148,N_18308);
nand U21912 (N_21912,N_19625,N_18258);
nor U21913 (N_21913,N_19751,N_18055);
xor U21914 (N_21914,N_18992,N_18268);
nor U21915 (N_21915,N_19175,N_18314);
nand U21916 (N_21916,N_19384,N_19905);
and U21917 (N_21917,N_19052,N_19669);
and U21918 (N_21918,N_19583,N_18230);
nor U21919 (N_21919,N_19816,N_18348);
nor U21920 (N_21920,N_18822,N_19245);
nor U21921 (N_21921,N_18385,N_18595);
xnor U21922 (N_21922,N_19290,N_19095);
nor U21923 (N_21923,N_19986,N_19298);
nand U21924 (N_21924,N_18037,N_19654);
or U21925 (N_21925,N_19087,N_19266);
and U21926 (N_21926,N_18500,N_18765);
nand U21927 (N_21927,N_19265,N_19266);
nand U21928 (N_21928,N_19335,N_19450);
nand U21929 (N_21929,N_19793,N_19020);
and U21930 (N_21930,N_18796,N_19864);
nor U21931 (N_21931,N_19242,N_18151);
nand U21932 (N_21932,N_19428,N_18790);
nand U21933 (N_21933,N_19529,N_18292);
nand U21934 (N_21934,N_18700,N_19668);
nand U21935 (N_21935,N_19731,N_19117);
and U21936 (N_21936,N_19563,N_19498);
nand U21937 (N_21937,N_18217,N_18766);
or U21938 (N_21938,N_19015,N_19999);
nor U21939 (N_21939,N_18967,N_18322);
and U21940 (N_21940,N_19288,N_19384);
xor U21941 (N_21941,N_18992,N_19539);
nand U21942 (N_21942,N_18524,N_18338);
nor U21943 (N_21943,N_18949,N_19595);
or U21944 (N_21944,N_18073,N_18493);
xor U21945 (N_21945,N_18517,N_18490);
and U21946 (N_21946,N_19797,N_19445);
nor U21947 (N_21947,N_18320,N_19400);
and U21948 (N_21948,N_18144,N_18990);
xor U21949 (N_21949,N_18156,N_19379);
and U21950 (N_21950,N_19679,N_18082);
nand U21951 (N_21951,N_19696,N_19402);
and U21952 (N_21952,N_19484,N_19614);
or U21953 (N_21953,N_18766,N_18456);
nand U21954 (N_21954,N_18565,N_19953);
and U21955 (N_21955,N_18004,N_18076);
nand U21956 (N_21956,N_18832,N_19594);
nor U21957 (N_21957,N_18202,N_19830);
and U21958 (N_21958,N_18421,N_18267);
nand U21959 (N_21959,N_19742,N_19537);
nand U21960 (N_21960,N_19620,N_19735);
xnor U21961 (N_21961,N_18162,N_18848);
and U21962 (N_21962,N_18893,N_19839);
or U21963 (N_21963,N_18138,N_18976);
and U21964 (N_21964,N_19685,N_19705);
nand U21965 (N_21965,N_19093,N_18774);
and U21966 (N_21966,N_19381,N_18513);
nor U21967 (N_21967,N_18891,N_19450);
nand U21968 (N_21968,N_19174,N_18741);
nor U21969 (N_21969,N_18167,N_18598);
and U21970 (N_21970,N_19079,N_19008);
nand U21971 (N_21971,N_19638,N_18935);
or U21972 (N_21972,N_18959,N_18563);
xnor U21973 (N_21973,N_18088,N_19804);
and U21974 (N_21974,N_18641,N_18335);
and U21975 (N_21975,N_19802,N_19130);
nor U21976 (N_21976,N_19133,N_19128);
nor U21977 (N_21977,N_18063,N_19845);
nand U21978 (N_21978,N_18191,N_18167);
xor U21979 (N_21979,N_19758,N_19356);
nand U21980 (N_21980,N_19990,N_19811);
and U21981 (N_21981,N_19185,N_18371);
nor U21982 (N_21982,N_18898,N_18666);
or U21983 (N_21983,N_18941,N_19436);
and U21984 (N_21984,N_19716,N_18527);
or U21985 (N_21985,N_19529,N_18790);
xor U21986 (N_21986,N_19014,N_18781);
and U21987 (N_21987,N_19945,N_18797);
nand U21988 (N_21988,N_18292,N_19093);
or U21989 (N_21989,N_19700,N_18144);
nand U21990 (N_21990,N_18296,N_19027);
or U21991 (N_21991,N_18764,N_19856);
nand U21992 (N_21992,N_18434,N_19195);
xor U21993 (N_21993,N_18160,N_18223);
nor U21994 (N_21994,N_19649,N_18762);
xor U21995 (N_21995,N_19645,N_18771);
nand U21996 (N_21996,N_18199,N_18962);
nor U21997 (N_21997,N_18755,N_19445);
nand U21998 (N_21998,N_19135,N_18329);
or U21999 (N_21999,N_18252,N_18952);
nand U22000 (N_22000,N_20603,N_20531);
nor U22001 (N_22001,N_20889,N_20554);
or U22002 (N_22002,N_20816,N_20944);
nor U22003 (N_22003,N_21901,N_20533);
or U22004 (N_22004,N_20403,N_21695);
xnor U22005 (N_22005,N_20496,N_21944);
and U22006 (N_22006,N_21294,N_20227);
nor U22007 (N_22007,N_20598,N_21021);
or U22008 (N_22008,N_21817,N_21130);
xnor U22009 (N_22009,N_21684,N_20854);
and U22010 (N_22010,N_20855,N_20100);
nand U22011 (N_22011,N_20036,N_20589);
or U22012 (N_22012,N_21401,N_21737);
nand U22013 (N_22013,N_20165,N_20608);
nor U22014 (N_22014,N_21381,N_20753);
xor U22015 (N_22015,N_21201,N_21721);
xor U22016 (N_22016,N_20984,N_21263);
nor U22017 (N_22017,N_21987,N_20459);
and U22018 (N_22018,N_20102,N_21417);
nor U22019 (N_22019,N_20006,N_21945);
and U22020 (N_22020,N_20880,N_20560);
nor U22021 (N_22021,N_21159,N_20260);
nor U22022 (N_22022,N_20966,N_20532);
xor U22023 (N_22023,N_20019,N_21559);
xnor U22024 (N_22024,N_20610,N_21383);
xor U22025 (N_22025,N_20446,N_20926);
nand U22026 (N_22026,N_21956,N_20826);
nand U22027 (N_22027,N_20059,N_21959);
nor U22028 (N_22028,N_21711,N_21606);
nand U22029 (N_22029,N_21533,N_21141);
xnor U22030 (N_22030,N_20520,N_21049);
nor U22031 (N_22031,N_21153,N_21003);
nand U22032 (N_22032,N_20968,N_20229);
and U22033 (N_22033,N_20136,N_21094);
nand U22034 (N_22034,N_21978,N_20699);
nand U22035 (N_22035,N_21477,N_21403);
or U22036 (N_22036,N_20343,N_21147);
xnor U22037 (N_22037,N_21903,N_20048);
or U22038 (N_22038,N_20576,N_21138);
and U22039 (N_22039,N_21667,N_21301);
nor U22040 (N_22040,N_20862,N_20927);
xor U22041 (N_22041,N_20977,N_21551);
nand U22042 (N_22042,N_21856,N_21904);
nor U22043 (N_22043,N_20545,N_20594);
and U22044 (N_22044,N_20461,N_20170);
or U22045 (N_22045,N_20015,N_21190);
or U22046 (N_22046,N_21756,N_20187);
nor U22047 (N_22047,N_21030,N_21079);
nand U22048 (N_22048,N_21665,N_20181);
and U22049 (N_22049,N_21988,N_20108);
or U22050 (N_22050,N_21697,N_21038);
nor U22051 (N_22051,N_20115,N_21523);
or U22052 (N_22052,N_21083,N_21429);
nand U22053 (N_22053,N_21453,N_21719);
nand U22054 (N_22054,N_20524,N_21882);
xnor U22055 (N_22055,N_20718,N_21686);
xnor U22056 (N_22056,N_21984,N_21171);
and U22057 (N_22057,N_21149,N_20592);
and U22058 (N_22058,N_21279,N_20857);
xnor U22059 (N_22059,N_21497,N_20457);
and U22060 (N_22060,N_20099,N_20068);
nor U22061 (N_22061,N_20578,N_20570);
or U22062 (N_22062,N_20482,N_21954);
nand U22063 (N_22063,N_20262,N_20755);
or U22064 (N_22064,N_20067,N_21894);
nor U22065 (N_22065,N_20606,N_21262);
nand U22066 (N_22066,N_20273,N_21860);
nand U22067 (N_22067,N_21179,N_21596);
nor U22068 (N_22068,N_20786,N_20504);
nand U22069 (N_22069,N_21035,N_20191);
xor U22070 (N_22070,N_20700,N_21785);
nand U22071 (N_22071,N_20013,N_21155);
or U22072 (N_22072,N_21034,N_20324);
nand U22073 (N_22073,N_20155,N_21108);
nor U22074 (N_22074,N_21610,N_20128);
nor U22075 (N_22075,N_21783,N_20807);
nor U22076 (N_22076,N_20123,N_21249);
or U22077 (N_22077,N_20991,N_21573);
or U22078 (N_22078,N_21512,N_21742);
nand U22079 (N_22079,N_21986,N_20904);
or U22080 (N_22080,N_20322,N_20963);
and U22081 (N_22081,N_21674,N_20632);
nor U22082 (N_22082,N_21370,N_20012);
or U22083 (N_22083,N_20318,N_21587);
and U22084 (N_22084,N_20618,N_20023);
nand U22085 (N_22085,N_21255,N_20865);
and U22086 (N_22086,N_21208,N_20484);
and U22087 (N_22087,N_20621,N_20667);
xor U22088 (N_22088,N_20039,N_20571);
xor U22089 (N_22089,N_20838,N_21295);
nor U22090 (N_22090,N_20580,N_20245);
or U22091 (N_22091,N_20124,N_21304);
nor U22092 (N_22092,N_20515,N_21656);
and U22093 (N_22093,N_21788,N_20360);
nand U22094 (N_22094,N_21847,N_21808);
and U22095 (N_22095,N_20025,N_21646);
and U22096 (N_22096,N_21603,N_21322);
nor U22097 (N_22097,N_20922,N_21919);
and U22098 (N_22098,N_21471,N_21902);
and U22099 (N_22099,N_20648,N_21963);
xor U22100 (N_22100,N_20134,N_20144);
and U22101 (N_22101,N_21253,N_20710);
xor U22102 (N_22102,N_20467,N_20118);
or U22103 (N_22103,N_21096,N_20351);
nand U22104 (N_22104,N_20693,N_21886);
xnor U22105 (N_22105,N_20595,N_20433);
and U22106 (N_22106,N_20490,N_21122);
nand U22107 (N_22107,N_21770,N_20998);
xor U22108 (N_22108,N_21015,N_20280);
nor U22109 (N_22109,N_20659,N_21617);
xnor U22110 (N_22110,N_20051,N_21811);
xnor U22111 (N_22111,N_20327,N_21259);
xnor U22112 (N_22112,N_20783,N_20089);
xor U22113 (N_22113,N_21273,N_20236);
xnor U22114 (N_22114,N_21728,N_20562);
nor U22115 (N_22115,N_21560,N_21070);
nand U22116 (N_22116,N_21604,N_21710);
and U22117 (N_22117,N_20762,N_20213);
nor U22118 (N_22118,N_21655,N_20691);
or U22119 (N_22119,N_20445,N_21812);
nand U22120 (N_22120,N_21935,N_20154);
and U22121 (N_22121,N_20375,N_21852);
xnor U22122 (N_22122,N_21763,N_20321);
or U22123 (N_22123,N_21082,N_20526);
nor U22124 (N_22124,N_20145,N_21467);
nor U22125 (N_22125,N_21333,N_20701);
nand U22126 (N_22126,N_21715,N_20449);
xnor U22127 (N_22127,N_20217,N_21223);
xnor U22128 (N_22128,N_20081,N_20418);
nand U22129 (N_22129,N_20917,N_21237);
nand U22130 (N_22130,N_21486,N_20787);
xnor U22131 (N_22131,N_20429,N_20483);
and U22132 (N_22132,N_20739,N_20827);
xnor U22133 (N_22133,N_21182,N_20368);
nor U22134 (N_22134,N_20579,N_21880);
nand U22135 (N_22135,N_20480,N_20292);
and U22136 (N_22136,N_21680,N_20822);
xnor U22137 (N_22137,N_20004,N_21806);
nor U22138 (N_22138,N_20702,N_21885);
nor U22139 (N_22139,N_21651,N_20272);
nor U22140 (N_22140,N_21011,N_20934);
nor U22141 (N_22141,N_21853,N_20999);
and U22142 (N_22142,N_21782,N_20831);
or U22143 (N_22143,N_20551,N_20088);
nand U22144 (N_22144,N_21845,N_20703);
nor U22145 (N_22145,N_21535,N_21229);
xor U22146 (N_22146,N_21008,N_20732);
nor U22147 (N_22147,N_21809,N_20597);
or U22148 (N_22148,N_20333,N_21837);
and U22149 (N_22149,N_21058,N_20132);
and U22150 (N_22150,N_20489,N_21996);
nor U22151 (N_22151,N_21396,N_21567);
nand U22152 (N_22152,N_20507,N_20296);
or U22153 (N_22153,N_21462,N_21591);
nand U22154 (N_22154,N_21608,N_21242);
or U22155 (N_22155,N_20736,N_21773);
xor U22156 (N_22156,N_20297,N_20874);
nand U22157 (N_22157,N_21759,N_21772);
xnor U22158 (N_22158,N_20080,N_21009);
nor U22159 (N_22159,N_21464,N_20789);
nand U22160 (N_22160,N_21930,N_21245);
or U22161 (N_22161,N_21946,N_20399);
nand U22162 (N_22162,N_21735,N_21514);
and U22163 (N_22163,N_21064,N_20247);
nor U22164 (N_22164,N_20198,N_20705);
nand U22165 (N_22165,N_20127,N_21906);
and U22166 (N_22166,N_21142,N_20278);
or U22167 (N_22167,N_21394,N_21271);
nor U22168 (N_22168,N_21629,N_20364);
and U22169 (N_22169,N_20546,N_21781);
nand U22170 (N_22170,N_20293,N_20920);
xnor U22171 (N_22171,N_21797,N_21161);
and U22172 (N_22172,N_20239,N_21990);
or U22173 (N_22173,N_20731,N_20176);
nand U22174 (N_22174,N_21572,N_21023);
and U22175 (N_22175,N_20498,N_20042);
and U22176 (N_22176,N_20972,N_21983);
and U22177 (N_22177,N_20211,N_21998);
nand U22178 (N_22178,N_20000,N_21341);
nor U22179 (N_22179,N_20122,N_20210);
nand U22180 (N_22180,N_21795,N_20500);
xor U22181 (N_22181,N_20715,N_20866);
nand U22182 (N_22182,N_21205,N_20335);
xnor U22183 (N_22183,N_21115,N_20848);
nand U22184 (N_22184,N_21579,N_20362);
and U22185 (N_22185,N_21189,N_20923);
nor U22186 (N_22186,N_20689,N_20945);
xor U22187 (N_22187,N_21734,N_20350);
or U22188 (N_22188,N_21713,N_21750);
nor U22189 (N_22189,N_21326,N_20224);
and U22190 (N_22190,N_20508,N_20680);
or U22191 (N_22191,N_21466,N_20312);
or U22192 (N_22192,N_20555,N_20957);
and U22193 (N_22193,N_20394,N_20425);
and U22194 (N_22194,N_20954,N_20331);
xor U22195 (N_22195,N_20558,N_20354);
nand U22196 (N_22196,N_21303,N_21068);
xnor U22197 (N_22197,N_21601,N_21029);
and U22198 (N_22198,N_21169,N_21361);
and U22199 (N_22199,N_21864,N_20810);
xor U22200 (N_22200,N_20682,N_20129);
nor U22201 (N_22201,N_20405,N_21484);
nand U22202 (N_22202,N_20392,N_21553);
nor U22203 (N_22203,N_21164,N_20402);
nand U22204 (N_22204,N_20175,N_20694);
nand U22205 (N_22205,N_21209,N_20502);
nand U22206 (N_22206,N_21185,N_21291);
and U22207 (N_22207,N_21947,N_20567);
nand U22208 (N_22208,N_20076,N_20289);
nor U22209 (N_22209,N_20778,N_20024);
and U22210 (N_22210,N_21283,N_20843);
or U22211 (N_22211,N_21243,N_20381);
xor U22212 (N_22212,N_21200,N_20252);
nor U22213 (N_22213,N_21940,N_21373);
nor U22214 (N_22214,N_21925,N_20269);
xnor U22215 (N_22215,N_21405,N_21236);
or U22216 (N_22216,N_21520,N_21505);
nor U22217 (N_22217,N_20338,N_20714);
nand U22218 (N_22218,N_20665,N_21548);
xnor U22219 (N_22219,N_20883,N_20628);
or U22220 (N_22220,N_21084,N_20591);
nand U22221 (N_22221,N_21432,N_21315);
or U22222 (N_22222,N_21526,N_20650);
and U22223 (N_22223,N_21942,N_21897);
xor U22224 (N_22224,N_21198,N_21004);
and U22225 (N_22225,N_21327,N_20007);
xor U22226 (N_22226,N_20481,N_21356);
nand U22227 (N_22227,N_21430,N_20232);
or U22228 (N_22228,N_21588,N_21324);
nor U22229 (N_22229,N_20879,N_21659);
nand U22230 (N_22230,N_21421,N_21884);
nand U22231 (N_22231,N_20540,N_21445);
and U22232 (N_22232,N_21195,N_21402);
nand U22233 (N_22233,N_20361,N_21632);
xor U22234 (N_22234,N_20468,N_20802);
or U22235 (N_22235,N_21751,N_20427);
or U22236 (N_22236,N_21530,N_20172);
or U22237 (N_22237,N_21335,N_20133);
and U22238 (N_22238,N_20726,N_20918);
and U22239 (N_22239,N_20776,N_21664);
or U22240 (N_22240,N_21826,N_21764);
xnor U22241 (N_22241,N_21865,N_21688);
or U22242 (N_22242,N_21412,N_20887);
xor U22243 (N_22243,N_21057,N_20315);
nor U22244 (N_22244,N_20847,N_20139);
nor U22245 (N_22245,N_21091,N_20743);
and U22246 (N_22246,N_21937,N_21334);
nand U22247 (N_22247,N_21887,N_20426);
nor U22248 (N_22248,N_21148,N_20435);
nor U22249 (N_22249,N_20347,N_21131);
or U22250 (N_22250,N_20738,N_20685);
and U22251 (N_22251,N_21280,N_20065);
xor U22252 (N_22252,N_21225,N_20713);
or U22253 (N_22253,N_20419,N_20975);
xor U22254 (N_22254,N_21689,N_21836);
and U22255 (N_22255,N_21152,N_20541);
xnor U22256 (N_22256,N_20575,N_20043);
nand U22257 (N_22257,N_21515,N_21472);
nor U22258 (N_22258,N_20121,N_21626);
or U22259 (N_22259,N_21392,N_20149);
or U22260 (N_22260,N_21406,N_20267);
or U22261 (N_22261,N_20029,N_21475);
xnor U22262 (N_22262,N_20462,N_21020);
nor U22263 (N_22263,N_21511,N_21036);
or U22264 (N_22264,N_21168,N_20937);
xnor U22265 (N_22265,N_20309,N_20931);
xnor U22266 (N_22266,N_20179,N_20897);
xnor U22267 (N_22267,N_20844,N_21418);
nand U22268 (N_22268,N_20385,N_20030);
or U22269 (N_22269,N_20098,N_21916);
nand U22270 (N_22270,N_20057,N_21855);
nor U22271 (N_22271,N_21972,N_21961);
xnor U22272 (N_22272,N_20661,N_21543);
xnor U22273 (N_22273,N_20298,N_20003);
nand U22274 (N_22274,N_20105,N_21268);
nand U22275 (N_22275,N_21879,N_21849);
xnor U22276 (N_22276,N_20775,N_20219);
and U22277 (N_22277,N_21419,N_20021);
nor U22278 (N_22278,N_21558,N_21144);
and U22279 (N_22279,N_20161,N_21053);
and U22280 (N_22280,N_21000,N_20027);
nand U22281 (N_22281,N_21634,N_21106);
nor U22282 (N_22282,N_20640,N_21639);
xnor U22283 (N_22283,N_20040,N_20241);
nor U22284 (N_22284,N_20183,N_21031);
or U22285 (N_22285,N_21831,N_21816);
nor U22286 (N_22286,N_21720,N_21235);
or U22287 (N_22287,N_20765,N_21687);
or U22288 (N_22288,N_20474,N_20939);
nor U22289 (N_22289,N_21620,N_20050);
xnor U22290 (N_22290,N_21063,N_21092);
or U22291 (N_22291,N_20494,N_21557);
or U22292 (N_22292,N_20537,N_21985);
and U22293 (N_22293,N_21362,N_21896);
nor U22294 (N_22294,N_20517,N_21565);
or U22295 (N_22295,N_20442,N_20463);
or U22296 (N_22296,N_21193,N_20131);
and U22297 (N_22297,N_20248,N_20820);
or U22298 (N_22298,N_21246,N_21460);
and U22299 (N_22299,N_21121,N_21099);
xor U22300 (N_22300,N_20281,N_20987);
xnor U22301 (N_22301,N_20777,N_21823);
and U22302 (N_22302,N_20654,N_20919);
xnor U22303 (N_22303,N_21647,N_21452);
nor U22304 (N_22304,N_21732,N_21834);
nor U22305 (N_22305,N_21873,N_20754);
and U22306 (N_22306,N_21850,N_20861);
and U22307 (N_22307,N_20203,N_20371);
or U22308 (N_22308,N_21910,N_21982);
nand U22309 (N_22309,N_20189,N_21329);
nor U22310 (N_22310,N_20936,N_20670);
or U22311 (N_22311,N_20075,N_20629);
nand U22312 (N_22312,N_20471,N_20573);
nor U22313 (N_22313,N_20649,N_20949);
nor U22314 (N_22314,N_20237,N_20564);
or U22315 (N_22315,N_21256,N_21261);
nand U22316 (N_22316,N_20758,N_20623);
nor U22317 (N_22317,N_20990,N_20274);
xor U22318 (N_22318,N_20216,N_20569);
nand U22319 (N_22319,N_20087,N_20005);
and U22320 (N_22320,N_21156,N_20069);
nor U22321 (N_22321,N_20071,N_21041);
and U22322 (N_22322,N_21499,N_20091);
nand U22323 (N_22323,N_20177,N_20801);
xnor U22324 (N_22324,N_20935,N_21380);
or U22325 (N_22325,N_21747,N_20363);
nand U22326 (N_22326,N_21479,N_21621);
nand U22327 (N_22327,N_21233,N_21891);
nand U22328 (N_22328,N_20994,N_21794);
nand U22329 (N_22329,N_21389,N_21671);
nand U22330 (N_22330,N_21349,N_20858);
and U22331 (N_22331,N_20456,N_21248);
and U22332 (N_22332,N_20645,N_20817);
nor U22333 (N_22333,N_20492,N_21594);
xnor U22334 (N_22334,N_21648,N_21977);
xor U22335 (N_22335,N_20053,N_21490);
nor U22336 (N_22336,N_21739,N_21493);
or U22337 (N_22337,N_20344,N_21012);
nand U22338 (N_22338,N_20891,N_20431);
nor U22339 (N_22339,N_21292,N_21685);
nand U22340 (N_22340,N_20249,N_21024);
xor U22341 (N_22341,N_20959,N_20378);
and U22342 (N_22342,N_21178,N_21563);
nand U22343 (N_22343,N_20358,N_21792);
nor U22344 (N_22344,N_21239,N_20748);
or U22345 (N_22345,N_20141,N_21032);
and U22346 (N_22346,N_20270,N_20107);
nand U22347 (N_22347,N_21939,N_20720);
nand U22348 (N_22348,N_20148,N_21701);
xnor U22349 (N_22349,N_20444,N_20047);
nor U22350 (N_22350,N_20986,N_20448);
or U22351 (N_22351,N_20721,N_20978);
nor U22352 (N_22352,N_20566,N_21638);
nand U22353 (N_22353,N_20464,N_21556);
or U22354 (N_22354,N_21958,N_21397);
nand U22355 (N_22355,N_20214,N_20523);
xnor U22356 (N_22356,N_20353,N_21913);
nor U22357 (N_22357,N_21395,N_21250);
nor U22358 (N_22358,N_20921,N_20008);
nand U22359 (N_22359,N_21272,N_21693);
nor U22360 (N_22360,N_20153,N_20276);
nor U22361 (N_22361,N_21644,N_20653);
and U22362 (N_22362,N_21900,N_20611);
and U22363 (N_22363,N_21677,N_20834);
and U22364 (N_22364,N_20147,N_20782);
nor U22365 (N_22365,N_20259,N_21858);
or U22366 (N_22366,N_20877,N_21247);
nand U22367 (N_22367,N_20208,N_21337);
or U22368 (N_22368,N_21387,N_21230);
nand U22369 (N_22369,N_21344,N_21044);
or U22370 (N_22370,N_21345,N_21448);
nand U22371 (N_22371,N_21502,N_21284);
xor U22372 (N_22372,N_21833,N_20325);
xnor U22373 (N_22373,N_21375,N_20819);
or U22374 (N_22374,N_20372,N_20616);
and U22375 (N_22375,N_21931,N_21458);
xnor U22376 (N_22376,N_20011,N_21574);
xnor U22377 (N_22377,N_21920,N_21267);
and U22378 (N_22378,N_20706,N_20781);
nand U22379 (N_22379,N_20881,N_21727);
nor U22380 (N_22380,N_20723,N_20641);
xor U22381 (N_22381,N_21415,N_20600);
xnor U22382 (N_22382,N_20254,N_20840);
xor U22383 (N_22383,N_20910,N_20791);
nand U22384 (N_22384,N_20319,N_21163);
nand U22385 (N_22385,N_21384,N_20626);
nor U22386 (N_22386,N_20473,N_20976);
and U22387 (N_22387,N_20985,N_21948);
nand U22388 (N_22388,N_20942,N_21481);
and U22389 (N_22389,N_21114,N_21866);
xnor U22390 (N_22390,N_21874,N_20169);
nand U22391 (N_22391,N_21133,N_21595);
and U22392 (N_22392,N_20478,N_20173);
nand U22393 (N_22393,N_21615,N_21150);
nand U22394 (N_22394,N_21895,N_20020);
or U22395 (N_22395,N_20432,N_20989);
nand U22396 (N_22396,N_21909,N_21705);
and U22397 (N_22397,N_21981,N_20180);
xnor U22398 (N_22398,N_21504,N_21760);
nand U22399 (N_22399,N_20014,N_21933);
nand U22400 (N_22400,N_21889,N_20094);
nand U22401 (N_22401,N_20250,N_20398);
and U22402 (N_22402,N_21135,N_21241);
nor U22403 (N_22403,N_20982,N_21577);
or U22404 (N_22404,N_21211,N_20140);
or U22405 (N_22405,N_20636,N_21662);
xnor U22406 (N_22406,N_21605,N_20299);
xor U22407 (N_22407,N_20336,N_21372);
nand U22408 (N_22408,N_20709,N_21364);
and U22409 (N_22409,N_20932,N_20475);
nand U22410 (N_22410,N_20220,N_20406);
nor U22411 (N_22411,N_21700,N_21059);
xor U22412 (N_22412,N_21813,N_21777);
and U22413 (N_22413,N_21854,N_21872);
nor U22414 (N_22414,N_21974,N_21683);
nand U22415 (N_22415,N_21799,N_20915);
or U22416 (N_22416,N_21509,N_21798);
nor U22417 (N_22417,N_20348,N_21314);
xor U22418 (N_22418,N_21966,N_20408);
and U22419 (N_22419,N_21784,N_21410);
nand U22420 (N_22420,N_20757,N_21212);
or U22421 (N_22421,N_21623,N_21413);
and U22422 (N_22422,N_20302,N_21017);
or U22423 (N_22423,N_21277,N_21952);
nand U22424 (N_22424,N_20930,N_21851);
or U22425 (N_22425,N_21431,N_20503);
nor U22426 (N_22426,N_20828,N_20760);
nand U22427 (N_22427,N_20261,N_21226);
nand U22428 (N_22428,N_20717,N_21427);
nand U22429 (N_22429,N_21755,N_21180);
or U22430 (N_22430,N_20407,N_21843);
nor U22431 (N_22431,N_21391,N_20505);
nand U22432 (N_22432,N_21050,N_21580);
nand U22433 (N_22433,N_21582,N_20275);
nand U22434 (N_22434,N_20388,N_21300);
or U22435 (N_22435,N_20958,N_21726);
or U22436 (N_22436,N_21485,N_20642);
nand U22437 (N_22437,N_21654,N_20771);
or U22438 (N_22438,N_21446,N_20607);
xor U22439 (N_22439,N_21822,N_20766);
xnor U22440 (N_22440,N_20867,N_20704);
nor U22441 (N_22441,N_21970,N_21519);
nand U22442 (N_22442,N_21305,N_21332);
and U22443 (N_22443,N_20195,N_20470);
xnor U22444 (N_22444,N_21941,N_20719);
xnor U22445 (N_22445,N_20070,N_21218);
and U22446 (N_22446,N_21411,N_20303);
or U22447 (N_22447,N_20679,N_20192);
xnor U22448 (N_22448,N_21546,N_21359);
xnor U22449 (N_22449,N_20032,N_21488);
and U22450 (N_22450,N_20264,N_21740);
and U22451 (N_22451,N_20521,N_21491);
and U22452 (N_22452,N_20886,N_20202);
nor U22453 (N_22453,N_21143,N_21476);
and U22454 (N_22454,N_21564,N_21167);
and U22455 (N_22455,N_21691,N_21358);
and U22456 (N_22456,N_21881,N_21844);
nand U22457 (N_22457,N_21065,N_20519);
nand U22458 (N_22458,N_20614,N_21093);
nor U22459 (N_22459,N_20770,N_21037);
or U22460 (N_22460,N_20602,N_20750);
xnor U22461 (N_22461,N_21388,N_20599);
or U22462 (N_22462,N_20253,N_21366);
and U22463 (N_22463,N_21382,N_20125);
nand U22464 (N_22464,N_20768,N_21441);
and U22465 (N_22465,N_20946,N_20586);
xor U22466 (N_22466,N_21552,N_20101);
or U22467 (N_22467,N_21597,N_20488);
nand U22468 (N_22468,N_21151,N_20062);
and U22469 (N_22469,N_21602,N_21040);
or U22470 (N_22470,N_21435,N_21328);
nor U22471 (N_22471,N_20314,N_21522);
and U22472 (N_22472,N_21221,N_21501);
and U22473 (N_22473,N_21474,N_20655);
or U22474 (N_22474,N_20876,N_20868);
and U22475 (N_22475,N_21536,N_21213);
nand U22476 (N_22476,N_20619,N_20112);
or U22477 (N_22477,N_21778,N_20178);
nand U22478 (N_22478,N_21754,N_20044);
nor U22479 (N_22479,N_21583,N_20207);
nand U22480 (N_22480,N_21875,N_20633);
and U22481 (N_22481,N_21128,N_21669);
xor U22482 (N_22482,N_20479,N_21331);
nor U22483 (N_22483,N_21675,N_21628);
nor U22484 (N_22484,N_21371,N_20593);
xor U22485 (N_22485,N_21113,N_20962);
or U22486 (N_22486,N_20465,N_21297);
xnor U22487 (N_22487,N_20472,N_20965);
or U22488 (N_22488,N_21960,N_20221);
nor U22489 (N_22489,N_20413,N_21949);
xor U22490 (N_22490,N_20194,N_20251);
nand U22491 (N_22491,N_20522,N_20850);
nor U22492 (N_22492,N_20627,N_21955);
nand U22493 (N_22493,N_20114,N_21224);
nor U22494 (N_22494,N_20773,N_21348);
xnor U22495 (N_22495,N_21166,N_21173);
or U22496 (N_22496,N_21377,N_20662);
or U22497 (N_22497,N_21196,N_20637);
nor U22498 (N_22498,N_20815,N_20767);
nand U22499 (N_22499,N_21480,N_21494);
nand U22500 (N_22500,N_20223,N_21191);
or U22501 (N_22501,N_20041,N_20205);
and U22502 (N_22502,N_21496,N_20215);
xnor U22503 (N_22503,N_21134,N_20761);
or U22504 (N_22504,N_21915,N_21060);
nand U22505 (N_22505,N_21962,N_20342);
nand U22506 (N_22506,N_20676,N_21838);
or U22507 (N_22507,N_21492,N_21257);
nand U22508 (N_22508,N_20677,N_21576);
nand U22509 (N_22509,N_21254,N_20898);
nor U22510 (N_22510,N_20652,N_20400);
xnor U22511 (N_22511,N_21641,N_20895);
nor U22512 (N_22512,N_20851,N_21285);
nand U22513 (N_22513,N_20054,N_20647);
xor U22514 (N_22514,N_21018,N_20416);
xor U22515 (N_22515,N_21652,N_20209);
and U22516 (N_22516,N_20516,N_20103);
xor U22517 (N_22517,N_21336,N_21663);
or U22518 (N_22518,N_20971,N_20544);
xor U22519 (N_22519,N_20414,N_20657);
and U22520 (N_22520,N_20415,N_20357);
or U22521 (N_22521,N_21104,N_21566);
or U22522 (N_22522,N_21709,N_20163);
nor U22523 (N_22523,N_20171,N_20746);
xnor U22524 (N_22524,N_21994,N_21892);
nand U22525 (N_22525,N_20852,N_21821);
xnor U22526 (N_22526,N_20316,N_20231);
or U22527 (N_22527,N_21206,N_20997);
and U22528 (N_22528,N_20692,N_20864);
nand U22529 (N_22529,N_21022,N_21609);
or U22530 (N_22530,N_20981,N_21531);
xnor U22531 (N_22531,N_21805,N_20200);
nor U22532 (N_22532,N_20447,N_20605);
nand U22533 (N_22533,N_20196,N_21658);
xor U22534 (N_22534,N_20130,N_20969);
xnor U22535 (N_22535,N_20311,N_21428);
and U22536 (N_22536,N_21507,N_20234);
xor U22537 (N_22537,N_21433,N_20747);
nor U22538 (N_22538,N_21724,N_20026);
nand U22539 (N_22539,N_21470,N_21202);
and U22540 (N_22540,N_21450,N_21414);
or U22541 (N_22541,N_21635,N_21820);
nor U22542 (N_22542,N_20330,N_20980);
nand U22543 (N_22543,N_21343,N_21712);
or U22544 (N_22544,N_20334,N_20845);
nand U22545 (N_22545,N_21199,N_20093);
or U22546 (N_22546,N_20725,N_21296);
xor U22547 (N_22547,N_21575,N_20870);
xnor U22548 (N_22548,N_21047,N_21210);
xnor U22549 (N_22549,N_20974,N_21918);
nand U22550 (N_22550,N_21269,N_21310);
nand U22551 (N_22551,N_20830,N_20553);
nor U22552 (N_22552,N_20317,N_20117);
nand U22553 (N_22553,N_20332,N_20035);
and U22554 (N_22554,N_21537,N_20116);
xnor U22555 (N_22555,N_20790,N_20370);
or U22556 (N_22556,N_21929,N_20320);
nand U22557 (N_22557,N_21936,N_20695);
and U22558 (N_22558,N_20119,N_21160);
and U22559 (N_22559,N_20907,N_20222);
xor U22560 (N_22560,N_20157,N_20061);
or U22561 (N_22561,N_21863,N_20872);
and U22562 (N_22562,N_20367,N_21181);
nand U22563 (N_22563,N_21042,N_21203);
and U22564 (N_22564,N_21117,N_20443);
nand U22565 (N_22565,N_20450,N_21840);
nand U22566 (N_22566,N_21136,N_20894);
nor U22567 (N_22567,N_21204,N_21824);
nor U22568 (N_22568,N_21748,N_20631);
xor U22569 (N_22569,N_20912,N_21907);
and U22570 (N_22570,N_20792,N_21420);
nor U22571 (N_22571,N_21757,N_20437);
and U22572 (N_22572,N_21016,N_20095);
nand U22573 (N_22573,N_20106,N_20451);
xnor U22574 (N_22574,N_20669,N_21489);
or U22575 (N_22575,N_20993,N_20961);
xnor U22576 (N_22576,N_20441,N_20383);
and U22577 (N_22577,N_21216,N_21637);
xor U22578 (N_22578,N_21922,N_21753);
nand U22579 (N_22579,N_20882,N_21498);
xor U22580 (N_22580,N_20010,N_20785);
nand U22581 (N_22581,N_20587,N_20896);
xnor U22582 (N_22582,N_21101,N_21422);
nand U22583 (N_22583,N_21126,N_20708);
or U22584 (N_22584,N_21771,N_21282);
or U22585 (N_22585,N_20284,N_20411);
xor U22586 (N_22586,N_21733,N_21867);
xor U22587 (N_22587,N_21052,N_20849);
nor U22588 (N_22588,N_20724,N_21730);
nand U22589 (N_22589,N_20109,N_21426);
xor U22590 (N_22590,N_21631,N_20377);
xnor U22591 (N_22591,N_21717,N_20609);
and U22592 (N_22592,N_21692,N_21074);
nand U22593 (N_22593,N_21599,N_21100);
xor U22594 (N_22594,N_21600,N_21468);
or U22595 (N_22595,N_21067,N_20379);
and U22596 (N_22596,N_21815,N_20037);
xor U22597 (N_22597,N_21461,N_20584);
nand U22598 (N_22598,N_20818,N_21964);
xor U22599 (N_22599,N_21991,N_20271);
and U22600 (N_22600,N_21839,N_21527);
nor U22601 (N_22601,N_21473,N_21080);
nand U22602 (N_22602,N_20151,N_20967);
nor U22603 (N_22603,N_21614,N_20612);
nand U22604 (N_22604,N_20058,N_20453);
nor U22605 (N_22605,N_21001,N_20938);
nor U22606 (N_22606,N_21281,N_20733);
nor U22607 (N_22607,N_21616,N_21593);
nand U22608 (N_22608,N_21367,N_20288);
and U22609 (N_22609,N_21398,N_20410);
nand U22610 (N_22610,N_20305,N_20511);
nor U22611 (N_22611,N_20142,N_20613);
and U22612 (N_22612,N_21234,N_21400);
xor U22613 (N_22613,N_20486,N_21908);
xor U22614 (N_22614,N_20097,N_20643);
nor U22615 (N_22615,N_20646,N_20476);
xor U22616 (N_22616,N_21758,N_20563);
and U22617 (N_22617,N_21592,N_20688);
nand U22618 (N_22618,N_20728,N_20017);
nor U22619 (N_22619,N_20823,N_20146);
and U22620 (N_22620,N_21529,N_20730);
nor U22621 (N_22621,N_21718,N_21971);
or U22622 (N_22622,N_21266,N_20941);
or U22623 (N_22623,N_21917,N_20423);
xnor U22624 (N_22624,N_20832,N_20756);
nor U22625 (N_22625,N_21376,N_21877);
and U22626 (N_22626,N_21028,N_21087);
xor U22627 (N_22627,N_20268,N_20328);
nand U22628 (N_22628,N_21165,N_21027);
nor U22629 (N_22629,N_21111,N_21780);
nor U22630 (N_22630,N_20803,N_20635);
or U22631 (N_22631,N_20282,N_20780);
and U22632 (N_22632,N_21207,N_20583);
or U22633 (N_22633,N_20950,N_21129);
xor U22634 (N_22634,N_20525,N_20046);
xnor U22635 (N_22635,N_20814,N_21302);
xnor U22636 (N_22636,N_20916,N_21731);
nand U22637 (N_22637,N_20550,N_21048);
xnor U22638 (N_22638,N_21571,N_20197);
and U22639 (N_22639,N_20875,N_21127);
and U22640 (N_22640,N_21289,N_21706);
nand U22641 (N_22641,N_20956,N_20487);
or U22642 (N_22642,N_21423,N_21791);
or U22643 (N_22643,N_21157,N_21316);
and U22644 (N_22644,N_20345,N_21265);
or U22645 (N_22645,N_21738,N_20620);
xor U22646 (N_22646,N_21500,N_20233);
or U22647 (N_22647,N_20084,N_21832);
nor U22648 (N_22648,N_20434,N_20582);
or U22649 (N_22649,N_20226,N_21365);
nand U22650 (N_22650,N_20326,N_21439);
nand U22651 (N_22651,N_20162,N_21077);
xnor U22652 (N_22652,N_20529,N_20238);
or U22653 (N_22653,N_21924,N_20697);
nand U22654 (N_22654,N_20639,N_20556);
and U22655 (N_22655,N_20300,N_20243);
nand U22656 (N_22656,N_20617,N_21447);
nor U22657 (N_22657,N_21992,N_20016);
nand U22658 (N_22658,N_20668,N_20809);
xnor U22659 (N_22659,N_20346,N_20510);
and U22660 (N_22660,N_21578,N_20064);
nor U22661 (N_22661,N_21075,N_20527);
nor U22662 (N_22662,N_21222,N_21124);
or U22663 (N_22663,N_20382,N_20083);
or U22664 (N_22664,N_21694,N_21890);
xor U22665 (N_22665,N_20349,N_20028);
nand U22666 (N_22666,N_21859,N_21357);
xor U22667 (N_22667,N_20396,N_21926);
and U22668 (N_22668,N_21841,N_21934);
nand U22669 (N_22669,N_21102,N_20795);
xnor U22670 (N_22670,N_20373,N_20846);
or U22671 (N_22671,N_20900,N_20535);
and U22672 (N_22672,N_20513,N_20588);
and U22673 (N_22673,N_20277,N_21319);
or U22674 (N_22674,N_20390,N_20687);
xor U22675 (N_22675,N_20018,N_21555);
xnor U22676 (N_22676,N_21056,N_20577);
and U22677 (N_22677,N_20256,N_21549);
and U22678 (N_22678,N_20286,N_20188);
nand U22679 (N_22679,N_21360,N_20499);
and U22680 (N_22680,N_20369,N_20853);
xor U22681 (N_22681,N_20340,N_21061);
nor U22682 (N_22682,N_21487,N_20455);
xnor U22683 (N_22683,N_20110,N_20049);
or U22684 (N_22684,N_21090,N_21354);
nor U22685 (N_22685,N_20684,N_21274);
and U22686 (N_22686,N_20038,N_20996);
nand U22687 (N_22687,N_20307,N_20509);
nand U22688 (N_22688,N_21633,N_21508);
nand U22689 (N_22689,N_21459,N_20283);
xnor U22690 (N_22690,N_21765,N_21818);
nor U22691 (N_22691,N_20808,N_20824);
nand U22692 (N_22692,N_21624,N_21528);
nor U22693 (N_22693,N_20924,N_21309);
and U22694 (N_22694,N_20892,N_21154);
nand U22695 (N_22695,N_21532,N_20769);
xor U22696 (N_22696,N_20341,N_21682);
nor U22697 (N_22697,N_21089,N_20079);
nand U22698 (N_22698,N_21787,N_20543);
nor U22699 (N_22699,N_21585,N_20784);
nor U22700 (N_22700,N_20512,N_20893);
and U22701 (N_22701,N_20878,N_20077);
xor U22702 (N_22702,N_21869,N_21888);
nor U22703 (N_22703,N_21776,N_20052);
nor U22704 (N_22704,N_20811,N_21386);
or U22705 (N_22705,N_20466,N_21139);
or U22706 (N_22706,N_20111,N_21980);
or U22707 (N_22707,N_21132,N_21215);
and U22708 (N_22708,N_21105,N_20903);
or U22709 (N_22709,N_21550,N_20871);
nand U22710 (N_22710,N_20495,N_21066);
nor U22711 (N_22711,N_20788,N_21339);
or U22712 (N_22712,N_20359,N_20734);
nand U22713 (N_22713,N_20547,N_21095);
or U22714 (N_22714,N_20863,N_20190);
nor U22715 (N_22715,N_21451,N_21270);
xor U22716 (N_22716,N_21162,N_20391);
nor U22717 (N_22717,N_20752,N_20741);
or U22718 (N_22718,N_21989,N_20568);
xor U22719 (N_22719,N_20458,N_20313);
nor U22720 (N_22720,N_21857,N_21340);
nor U22721 (N_22721,N_20304,N_21416);
nor U22722 (N_22722,N_21862,N_21443);
and U22723 (N_22723,N_20841,N_21590);
and U22724 (N_22724,N_21842,N_20228);
nor U22725 (N_22725,N_21352,N_21046);
nor U22726 (N_22726,N_21228,N_21219);
xor U22727 (N_22727,N_21013,N_20266);
and U22728 (N_22728,N_21545,N_21231);
and U22729 (N_22729,N_21010,N_21538);
nand U22730 (N_22730,N_20888,N_21893);
nor U22731 (N_22731,N_21025,N_20159);
or U22732 (N_22732,N_21645,N_21943);
xor U22733 (N_22733,N_21643,N_21927);
xnor U22734 (N_22734,N_20664,N_21723);
nor U22735 (N_22735,N_21408,N_20698);
xnor U22736 (N_22736,N_21800,N_20737);
nand U22737 (N_22737,N_20799,N_21534);
nor U22738 (N_22738,N_20199,N_21118);
or U22739 (N_22739,N_21905,N_21145);
xnor U22740 (N_22740,N_20031,N_20797);
or U22741 (N_22741,N_20242,N_20630);
and U22742 (N_22742,N_20287,N_20074);
and U22743 (N_22743,N_21802,N_20514);
or U22744 (N_22744,N_20212,N_21744);
or U22745 (N_22745,N_21950,N_21478);
and U22746 (N_22746,N_21014,N_21338);
nor U22747 (N_22747,N_21932,N_20542);
and U22748 (N_22748,N_21766,N_21007);
xnor U22749 (N_22749,N_20675,N_20559);
nor U22750 (N_22750,N_21320,N_20913);
nand U22751 (N_22751,N_20420,N_21463);
and U22752 (N_22752,N_21547,N_21969);
or U22753 (N_22753,N_21078,N_20742);
xnor U22754 (N_22754,N_21186,N_21379);
nand U22755 (N_22755,N_20092,N_21673);
nand U22756 (N_22756,N_20301,N_20439);
and U22757 (N_22757,N_20255,N_20156);
or U22758 (N_22758,N_21598,N_21898);
nor U22759 (N_22759,N_21729,N_20120);
nor U22760 (N_22760,N_21137,N_20393);
and U22761 (N_22761,N_20422,N_21506);
or U22762 (N_22762,N_21275,N_21298);
nor U22763 (N_22763,N_20914,N_21404);
xnor U22764 (N_22764,N_20366,N_20909);
xor U22765 (N_22765,N_20951,N_21125);
xnor U22766 (N_22766,N_20240,N_20622);
nor U22767 (N_22767,N_20365,N_21516);
or U22768 (N_22768,N_21636,N_20905);
or U22769 (N_22769,N_20906,N_21790);
or U22770 (N_22770,N_20355,N_20096);
xor U22771 (N_22771,N_21330,N_20988);
nor U22772 (N_22772,N_21146,N_20671);
nor U22773 (N_22773,N_21240,N_21437);
nor U22774 (N_22774,N_20491,N_21584);
and U22775 (N_22775,N_20356,N_20995);
and U22776 (N_22776,N_21870,N_20796);
or U22777 (N_22777,N_21503,N_21979);
or U22778 (N_22778,N_21158,N_20992);
nor U22779 (N_22779,N_20285,N_20835);
xor U22780 (N_22780,N_20663,N_20409);
and U22781 (N_22781,N_20856,N_20160);
and U22782 (N_22782,N_20681,N_20722);
or U22783 (N_22783,N_21217,N_20263);
nor U22784 (N_22784,N_21690,N_20290);
xor U22785 (N_22785,N_20135,N_20970);
nand U22786 (N_22786,N_21581,N_20947);
or U22787 (N_22787,N_21707,N_20150);
nand U22788 (N_22788,N_20184,N_21848);
xnor U22789 (N_22789,N_21220,N_21482);
nand U22790 (N_22790,N_21103,N_20829);
xor U22791 (N_22791,N_21611,N_21539);
xnor U22792 (N_22792,N_21957,N_21188);
or U22793 (N_22793,N_20683,N_21123);
xnor U22794 (N_22794,N_21378,N_21997);
nor U22795 (N_22795,N_21390,N_21438);
xor U22796 (N_22796,N_20022,N_21055);
xor U22797 (N_22797,N_21835,N_20764);
nand U22798 (N_22798,N_20793,N_20666);
nand U22799 (N_22799,N_20644,N_20421);
nor U22800 (N_22800,N_21116,N_21796);
xnor U22801 (N_22801,N_21562,N_21019);
xnor U22802 (N_22802,N_20660,N_21708);
xor U22803 (N_22803,N_21542,N_20983);
nor U22804 (N_22804,N_21912,N_20774);
xor U22805 (N_22805,N_21227,N_20955);
nand U22806 (N_22806,N_20352,N_20066);
and U22807 (N_22807,N_20158,N_20585);
and U22808 (N_22808,N_21752,N_21786);
xnor U22809 (N_22809,N_20800,N_21187);
or U22810 (N_22810,N_20890,N_21561);
xor U22811 (N_22811,N_20979,N_21039);
or U22812 (N_22812,N_21630,N_21676);
and U22813 (N_22813,N_20716,N_20001);
and U22814 (N_22814,N_21434,N_20929);
nor U22815 (N_22815,N_20552,N_20206);
xor U22816 (N_22816,N_21368,N_21803);
or U22817 (N_22817,N_21002,N_20557);
xor U22818 (N_22818,N_20908,N_21071);
xor U22819 (N_22819,N_20574,N_20604);
nand U22820 (N_22820,N_21286,N_21544);
nand U22821 (N_22821,N_21827,N_21871);
nor U22822 (N_22822,N_21653,N_21088);
nor U22823 (N_22823,N_21308,N_20842);
nand U22824 (N_22824,N_21613,N_20174);
nor U22825 (N_22825,N_20310,N_20034);
xnor U22826 (N_22826,N_21440,N_20452);
or U22827 (N_22827,N_21672,N_21625);
nand U22828 (N_22828,N_21975,N_21069);
nand U22829 (N_22829,N_20836,N_20839);
nor U22830 (N_22830,N_20306,N_20063);
or U22831 (N_22831,N_21192,N_21642);
and U22832 (N_22832,N_21666,N_20258);
or U22833 (N_22833,N_20060,N_21085);
and U22834 (N_22834,N_20561,N_21006);
and U22835 (N_22835,N_20678,N_21214);
xnor U22836 (N_22836,N_21923,N_20672);
xor U22837 (N_22837,N_21313,N_20166);
nor U22838 (N_22838,N_20225,N_21456);
or U22839 (N_22839,N_20873,N_21425);
or U22840 (N_22840,N_20601,N_20911);
nor U22841 (N_22841,N_21670,N_21883);
nor U22842 (N_22842,N_21293,N_21846);
nor U22843 (N_22843,N_21681,N_20821);
nand U22844 (N_22844,N_21098,N_20485);
and U22845 (N_22845,N_20590,N_20804);
nand U22846 (N_22846,N_20530,N_20501);
xor U22847 (N_22847,N_21702,N_21678);
or U22848 (N_22848,N_20204,N_21455);
or U22849 (N_22849,N_21789,N_20727);
nand U22850 (N_22850,N_20082,N_20104);
and U22851 (N_22851,N_20902,N_21260);
or U22852 (N_22852,N_21745,N_21569);
or U22853 (N_22853,N_20469,N_21184);
or U22854 (N_22854,N_21311,N_20869);
or U22855 (N_22855,N_20460,N_21868);
or U22856 (N_22856,N_21725,N_20073);
and U22857 (N_22857,N_21825,N_20658);
nand U22858 (N_22858,N_21045,N_21072);
and U22859 (N_22859,N_21176,N_21276);
nand U22860 (N_22860,N_21657,N_21252);
and U22861 (N_22861,N_20235,N_20744);
nor U22862 (N_22862,N_21554,N_20033);
nor U22863 (N_22863,N_21704,N_20090);
and U22864 (N_22864,N_20964,N_21810);
or U22865 (N_22865,N_21351,N_20167);
and U22866 (N_22866,N_21469,N_20002);
nor U22867 (N_22867,N_21649,N_21513);
and U22868 (N_22868,N_20086,N_21465);
nor U22869 (N_22869,N_21876,N_21109);
nand U22870 (N_22870,N_20265,N_21779);
or U22871 (N_22871,N_21140,N_21928);
nand U22872 (N_22872,N_20389,N_20812);
xor U22873 (N_22873,N_21775,N_21172);
xnor U22874 (N_22874,N_20376,N_21568);
nor U22875 (N_22875,N_20596,N_20436);
nand U22876 (N_22876,N_20925,N_20138);
or U22877 (N_22877,N_21973,N_21761);
nor U22878 (N_22878,N_20113,N_21307);
nand U22879 (N_22879,N_20572,N_20440);
nor U22880 (N_22880,N_21703,N_21174);
xor U22881 (N_22881,N_21197,N_21619);
xor U22882 (N_22882,N_20164,N_21807);
or U22883 (N_22883,N_20656,N_20674);
xnor U22884 (N_22884,N_20860,N_20518);
and U22885 (N_22885,N_20143,N_20374);
nor U22886 (N_22886,N_21107,N_20126);
or U22887 (N_22887,N_20885,N_20933);
or U22888 (N_22888,N_20749,N_20960);
nor U22889 (N_22889,N_20948,N_21407);
or U22890 (N_22890,N_21540,N_20696);
nand U22891 (N_22891,N_20901,N_20538);
and U22892 (N_22892,N_20384,N_20045);
or U22893 (N_22893,N_20078,N_21385);
or U22894 (N_22894,N_20686,N_21743);
nor U22895 (N_22895,N_21660,N_20438);
nor U22896 (N_22896,N_20884,N_20056);
xor U22897 (N_22897,N_20707,N_21026);
or U22898 (N_22898,N_20417,N_21342);
and U22899 (N_22899,N_21570,N_20806);
and U22900 (N_22900,N_21442,N_20244);
nand U22901 (N_22901,N_20137,N_20182);
or U22902 (N_22902,N_21668,N_20412);
and U22903 (N_22903,N_21951,N_20493);
and U22904 (N_22904,N_21321,N_20257);
and U22905 (N_22905,N_21622,N_21346);
or U22906 (N_22906,N_21650,N_21495);
nor U22907 (N_22907,N_21741,N_20401);
xor U22908 (N_22908,N_20193,N_20615);
and U22909 (N_22909,N_20740,N_20323);
nand U22910 (N_22910,N_20430,N_20759);
nand U22911 (N_22911,N_20690,N_21244);
nor U22912 (N_22912,N_21793,N_21517);
nor U22913 (N_22913,N_21627,N_21194);
xnor U22914 (N_22914,N_20218,N_21819);
nor U22915 (N_22915,N_21076,N_20928);
or U22916 (N_22916,N_21768,N_20454);
nor U22917 (N_22917,N_21762,N_21399);
and U22918 (N_22918,N_21938,N_20973);
nor U22919 (N_22919,N_20152,N_21170);
or U22920 (N_22920,N_20825,N_20729);
xnor U22921 (N_22921,N_21716,N_20634);
and U22922 (N_22922,N_21238,N_20859);
nand U22923 (N_22923,N_21444,N_20549);
nor U22924 (N_22924,N_20230,N_21804);
nor U22925 (N_22925,N_20952,N_21119);
nor U22926 (N_22926,N_21814,N_20477);
nand U22927 (N_22927,N_20779,N_20339);
nand U22928 (N_22928,N_20085,N_21318);
and U22929 (N_22929,N_21829,N_21288);
nor U22930 (N_22930,N_21525,N_21993);
nor U22931 (N_22931,N_20387,N_20711);
and U22932 (N_22932,N_21510,N_21347);
and U22933 (N_22933,N_21524,N_21921);
or U22934 (N_22934,N_20168,N_20534);
nand U22935 (N_22935,N_20794,N_21112);
xnor U22936 (N_22936,N_20404,N_21054);
xor U22937 (N_22937,N_20581,N_20329);
or U22938 (N_22938,N_20772,N_20751);
nor U22939 (N_22939,N_21177,N_20940);
or U22940 (N_22940,N_21612,N_21454);
nor U22941 (N_22941,N_20625,N_20833);
or U22942 (N_22942,N_21640,N_20539);
nand U22943 (N_22943,N_21911,N_20337);
nand U22944 (N_22944,N_21995,N_21062);
nand U22945 (N_22945,N_20397,N_20386);
xnor U22946 (N_22946,N_20798,N_21878);
nor U22947 (N_22947,N_21086,N_20506);
xnor U22948 (N_22948,N_21968,N_20536);
or U22949 (N_22949,N_21350,N_20837);
xor U22950 (N_22950,N_21589,N_21999);
nand U22951 (N_22951,N_21769,N_20745);
xor U22952 (N_22952,N_21317,N_21698);
nor U22953 (N_22953,N_21830,N_20279);
nor U22954 (N_22954,N_21661,N_20528);
xor U22955 (N_22955,N_21353,N_21120);
and U22956 (N_22956,N_21287,N_20638);
and U22957 (N_22957,N_21251,N_21696);
nor U22958 (N_22958,N_21899,N_21374);
xnor U22959 (N_22959,N_21175,N_21541);
or U22960 (N_22960,N_21457,N_20201);
nor U22961 (N_22961,N_21699,N_21767);
nor U22962 (N_22962,N_21278,N_20813);
xor U22963 (N_22963,N_21409,N_21258);
nor U22964 (N_22964,N_21749,N_21051);
or U22965 (N_22965,N_20424,N_21436);
xor U22966 (N_22966,N_21363,N_20380);
xnor U22967 (N_22967,N_20395,N_21312);
or U22968 (N_22968,N_21965,N_21521);
and U22969 (N_22969,N_21828,N_20246);
nor U22970 (N_22970,N_21369,N_21323);
and U22971 (N_22971,N_21618,N_20712);
nand U22972 (N_22972,N_20548,N_21586);
nand U22973 (N_22973,N_20295,N_21914);
and U22974 (N_22974,N_20805,N_20565);
nand U22975 (N_22975,N_21714,N_21518);
and U22976 (N_22976,N_21097,N_20185);
or U22977 (N_22977,N_21736,N_21393);
or U22978 (N_22978,N_20651,N_21801);
nand U22979 (N_22979,N_21299,N_21033);
nor U22980 (N_22980,N_21043,N_21953);
nand U22981 (N_22981,N_20308,N_20294);
nand U22982 (N_22982,N_20291,N_21306);
nor U22983 (N_22983,N_21005,N_21967);
and U22984 (N_22984,N_21325,N_21449);
or U22985 (N_22985,N_21976,N_21110);
nor U22986 (N_22986,N_21081,N_21722);
nor U22987 (N_22987,N_20428,N_20763);
and U22988 (N_22988,N_20943,N_21290);
nand U22989 (N_22989,N_21183,N_21232);
nand U22990 (N_22990,N_21424,N_21607);
xnor U22991 (N_22991,N_21679,N_20186);
xor U22992 (N_22992,N_21355,N_20735);
or U22993 (N_22993,N_21264,N_21861);
xnor U22994 (N_22994,N_21746,N_20072);
or U22995 (N_22995,N_20055,N_20624);
and U22996 (N_22996,N_20899,N_21073);
or U22997 (N_22997,N_21483,N_20953);
and U22998 (N_22998,N_20009,N_21774);
nand U22999 (N_22999,N_20673,N_20497);
xnor U23000 (N_23000,N_21987,N_20477);
and U23001 (N_23001,N_20610,N_20229);
nand U23002 (N_23002,N_21721,N_20298);
and U23003 (N_23003,N_21371,N_20714);
and U23004 (N_23004,N_20425,N_21775);
nand U23005 (N_23005,N_20658,N_21289);
or U23006 (N_23006,N_21135,N_20385);
nor U23007 (N_23007,N_20340,N_21728);
nor U23008 (N_23008,N_21908,N_21275);
xnor U23009 (N_23009,N_21987,N_21565);
xnor U23010 (N_23010,N_21856,N_21109);
or U23011 (N_23011,N_21473,N_21843);
nor U23012 (N_23012,N_20216,N_20883);
and U23013 (N_23013,N_20823,N_20126);
nor U23014 (N_23014,N_20140,N_20312);
xnor U23015 (N_23015,N_20891,N_20063);
xnor U23016 (N_23016,N_21395,N_21607);
nand U23017 (N_23017,N_20465,N_21943);
or U23018 (N_23018,N_21371,N_21729);
or U23019 (N_23019,N_21186,N_21065);
nor U23020 (N_23020,N_20007,N_20235);
and U23021 (N_23021,N_20796,N_20007);
nor U23022 (N_23022,N_20524,N_20999);
nand U23023 (N_23023,N_21538,N_21268);
and U23024 (N_23024,N_21302,N_20837);
or U23025 (N_23025,N_21504,N_20084);
nand U23026 (N_23026,N_20757,N_20238);
nand U23027 (N_23027,N_21943,N_20847);
or U23028 (N_23028,N_20570,N_20959);
or U23029 (N_23029,N_21220,N_21542);
nor U23030 (N_23030,N_20886,N_20681);
nand U23031 (N_23031,N_20589,N_21015);
nor U23032 (N_23032,N_20974,N_20887);
nand U23033 (N_23033,N_20816,N_21130);
nor U23034 (N_23034,N_21672,N_21762);
or U23035 (N_23035,N_20277,N_20612);
xor U23036 (N_23036,N_20020,N_20642);
nor U23037 (N_23037,N_20389,N_21238);
nand U23038 (N_23038,N_21075,N_21639);
and U23039 (N_23039,N_20994,N_20852);
xor U23040 (N_23040,N_20575,N_20604);
xor U23041 (N_23041,N_20062,N_20645);
and U23042 (N_23042,N_20506,N_20261);
nand U23043 (N_23043,N_20682,N_20411);
nor U23044 (N_23044,N_21794,N_21512);
and U23045 (N_23045,N_20623,N_20246);
and U23046 (N_23046,N_21115,N_21016);
xor U23047 (N_23047,N_20009,N_21173);
nor U23048 (N_23048,N_20453,N_20667);
xor U23049 (N_23049,N_21253,N_21876);
nand U23050 (N_23050,N_20507,N_21888);
nand U23051 (N_23051,N_21494,N_20186);
or U23052 (N_23052,N_20629,N_20110);
nand U23053 (N_23053,N_20893,N_21497);
xor U23054 (N_23054,N_21249,N_21725);
and U23055 (N_23055,N_20545,N_21879);
xnor U23056 (N_23056,N_20953,N_20576);
and U23057 (N_23057,N_21011,N_21226);
or U23058 (N_23058,N_20487,N_21042);
nand U23059 (N_23059,N_21414,N_20324);
and U23060 (N_23060,N_21150,N_20899);
nor U23061 (N_23061,N_20874,N_21070);
nand U23062 (N_23062,N_20446,N_21102);
nor U23063 (N_23063,N_21930,N_20947);
nand U23064 (N_23064,N_21245,N_20486);
nand U23065 (N_23065,N_21919,N_21757);
and U23066 (N_23066,N_20637,N_20853);
xnor U23067 (N_23067,N_20926,N_20764);
and U23068 (N_23068,N_20570,N_20971);
xnor U23069 (N_23069,N_21427,N_21607);
and U23070 (N_23070,N_21493,N_21627);
nand U23071 (N_23071,N_21460,N_21510);
and U23072 (N_23072,N_20534,N_20113);
or U23073 (N_23073,N_20560,N_20123);
xor U23074 (N_23074,N_20914,N_21940);
or U23075 (N_23075,N_21875,N_21009);
nand U23076 (N_23076,N_21209,N_20511);
nand U23077 (N_23077,N_20570,N_20476);
and U23078 (N_23078,N_20087,N_21119);
nor U23079 (N_23079,N_20097,N_21954);
or U23080 (N_23080,N_20354,N_21150);
nand U23081 (N_23081,N_20752,N_20565);
xor U23082 (N_23082,N_20442,N_20167);
nor U23083 (N_23083,N_20914,N_21339);
or U23084 (N_23084,N_21306,N_20820);
and U23085 (N_23085,N_21937,N_20670);
nand U23086 (N_23086,N_20173,N_20191);
xnor U23087 (N_23087,N_20132,N_20039);
xnor U23088 (N_23088,N_20097,N_21396);
xnor U23089 (N_23089,N_20777,N_21834);
xor U23090 (N_23090,N_20802,N_20657);
nand U23091 (N_23091,N_20725,N_21959);
or U23092 (N_23092,N_21352,N_21518);
or U23093 (N_23093,N_21556,N_21973);
nand U23094 (N_23094,N_20317,N_20643);
or U23095 (N_23095,N_21817,N_21451);
nand U23096 (N_23096,N_21800,N_20452);
xnor U23097 (N_23097,N_20785,N_21789);
xnor U23098 (N_23098,N_20747,N_20485);
xnor U23099 (N_23099,N_21359,N_20771);
xor U23100 (N_23100,N_21183,N_21312);
xnor U23101 (N_23101,N_21318,N_20879);
nand U23102 (N_23102,N_21924,N_20002);
and U23103 (N_23103,N_20076,N_20498);
nor U23104 (N_23104,N_21717,N_20616);
and U23105 (N_23105,N_20454,N_21340);
xor U23106 (N_23106,N_21200,N_21565);
or U23107 (N_23107,N_20613,N_21108);
nand U23108 (N_23108,N_21143,N_21377);
or U23109 (N_23109,N_21326,N_20975);
nor U23110 (N_23110,N_20542,N_21309);
and U23111 (N_23111,N_21654,N_21420);
nor U23112 (N_23112,N_21421,N_20043);
nor U23113 (N_23113,N_20853,N_20616);
nor U23114 (N_23114,N_20784,N_20929);
or U23115 (N_23115,N_20798,N_20614);
or U23116 (N_23116,N_20476,N_20157);
xnor U23117 (N_23117,N_20372,N_20915);
or U23118 (N_23118,N_20098,N_20718);
or U23119 (N_23119,N_21726,N_20355);
nor U23120 (N_23120,N_21034,N_20816);
nor U23121 (N_23121,N_20371,N_20350);
and U23122 (N_23122,N_21358,N_21742);
or U23123 (N_23123,N_21591,N_20427);
or U23124 (N_23124,N_20644,N_21456);
xnor U23125 (N_23125,N_20918,N_21447);
nor U23126 (N_23126,N_21626,N_21110);
or U23127 (N_23127,N_20127,N_20377);
nor U23128 (N_23128,N_21276,N_21609);
nor U23129 (N_23129,N_20171,N_21924);
xnor U23130 (N_23130,N_20497,N_21844);
xor U23131 (N_23131,N_20355,N_20470);
nand U23132 (N_23132,N_21043,N_21140);
xor U23133 (N_23133,N_20608,N_21586);
nand U23134 (N_23134,N_21448,N_20826);
xnor U23135 (N_23135,N_20568,N_20186);
and U23136 (N_23136,N_20217,N_20734);
and U23137 (N_23137,N_20597,N_21105);
xor U23138 (N_23138,N_20090,N_21831);
and U23139 (N_23139,N_21862,N_20243);
or U23140 (N_23140,N_21333,N_21002);
nand U23141 (N_23141,N_21304,N_20778);
nor U23142 (N_23142,N_21076,N_21194);
nor U23143 (N_23143,N_21822,N_20981);
or U23144 (N_23144,N_21805,N_20868);
or U23145 (N_23145,N_21309,N_20721);
or U23146 (N_23146,N_21527,N_20411);
or U23147 (N_23147,N_20855,N_21744);
xor U23148 (N_23148,N_21456,N_20582);
nor U23149 (N_23149,N_20260,N_21085);
nor U23150 (N_23150,N_20396,N_20016);
and U23151 (N_23151,N_20803,N_21239);
and U23152 (N_23152,N_21513,N_20809);
xor U23153 (N_23153,N_20456,N_20203);
nor U23154 (N_23154,N_20347,N_21421);
or U23155 (N_23155,N_20478,N_20058);
and U23156 (N_23156,N_20744,N_21270);
and U23157 (N_23157,N_21120,N_20904);
nand U23158 (N_23158,N_21257,N_21557);
and U23159 (N_23159,N_21010,N_21724);
nand U23160 (N_23160,N_21479,N_21782);
nand U23161 (N_23161,N_21828,N_20238);
and U23162 (N_23162,N_20177,N_21460);
nand U23163 (N_23163,N_21572,N_21411);
or U23164 (N_23164,N_20820,N_21681);
nand U23165 (N_23165,N_21061,N_20460);
or U23166 (N_23166,N_21917,N_20119);
or U23167 (N_23167,N_21719,N_21213);
or U23168 (N_23168,N_20149,N_21859);
nand U23169 (N_23169,N_21488,N_20705);
and U23170 (N_23170,N_20492,N_20711);
and U23171 (N_23171,N_20796,N_21847);
xnor U23172 (N_23172,N_20726,N_20877);
nor U23173 (N_23173,N_21719,N_20886);
and U23174 (N_23174,N_20809,N_20929);
or U23175 (N_23175,N_21718,N_21098);
nand U23176 (N_23176,N_21962,N_21943);
nor U23177 (N_23177,N_21289,N_21752);
xnor U23178 (N_23178,N_20971,N_21932);
nor U23179 (N_23179,N_21208,N_20828);
and U23180 (N_23180,N_20877,N_20530);
nor U23181 (N_23181,N_20429,N_21410);
nor U23182 (N_23182,N_20968,N_20941);
nor U23183 (N_23183,N_20218,N_21281);
nand U23184 (N_23184,N_20903,N_20068);
nand U23185 (N_23185,N_20780,N_20795);
nor U23186 (N_23186,N_20515,N_20399);
and U23187 (N_23187,N_21304,N_20933);
nor U23188 (N_23188,N_20575,N_20907);
and U23189 (N_23189,N_20911,N_21199);
nand U23190 (N_23190,N_21932,N_21124);
xor U23191 (N_23191,N_20024,N_20641);
and U23192 (N_23192,N_20749,N_20618);
nor U23193 (N_23193,N_20079,N_21119);
and U23194 (N_23194,N_21688,N_20285);
nor U23195 (N_23195,N_21070,N_20242);
or U23196 (N_23196,N_21278,N_20263);
nand U23197 (N_23197,N_20188,N_20944);
nor U23198 (N_23198,N_21565,N_20985);
and U23199 (N_23199,N_21988,N_20120);
nor U23200 (N_23200,N_20146,N_20043);
xnor U23201 (N_23201,N_21529,N_20596);
and U23202 (N_23202,N_21297,N_20767);
xnor U23203 (N_23203,N_20303,N_21134);
xor U23204 (N_23204,N_21175,N_21460);
and U23205 (N_23205,N_21558,N_21240);
or U23206 (N_23206,N_20326,N_20207);
nand U23207 (N_23207,N_21598,N_20037);
and U23208 (N_23208,N_21850,N_21329);
and U23209 (N_23209,N_21789,N_20705);
xnor U23210 (N_23210,N_21318,N_20546);
and U23211 (N_23211,N_20360,N_21765);
or U23212 (N_23212,N_20114,N_20264);
nor U23213 (N_23213,N_21834,N_21915);
xnor U23214 (N_23214,N_21416,N_21635);
or U23215 (N_23215,N_21949,N_21336);
nor U23216 (N_23216,N_20689,N_20799);
xor U23217 (N_23217,N_20668,N_21212);
or U23218 (N_23218,N_20512,N_21768);
or U23219 (N_23219,N_21769,N_21164);
nor U23220 (N_23220,N_21623,N_21170);
and U23221 (N_23221,N_20936,N_21209);
nand U23222 (N_23222,N_20818,N_20805);
xor U23223 (N_23223,N_21822,N_21106);
nand U23224 (N_23224,N_21886,N_21074);
nor U23225 (N_23225,N_21491,N_21102);
or U23226 (N_23226,N_21248,N_20623);
and U23227 (N_23227,N_21029,N_20151);
or U23228 (N_23228,N_20540,N_21487);
xor U23229 (N_23229,N_21444,N_21072);
nand U23230 (N_23230,N_21742,N_20792);
and U23231 (N_23231,N_20626,N_21744);
and U23232 (N_23232,N_21775,N_21470);
nor U23233 (N_23233,N_20783,N_20423);
xnor U23234 (N_23234,N_21387,N_21333);
or U23235 (N_23235,N_21593,N_21570);
nand U23236 (N_23236,N_21998,N_21584);
nor U23237 (N_23237,N_21846,N_20075);
nand U23238 (N_23238,N_21211,N_20534);
xnor U23239 (N_23239,N_21502,N_21899);
or U23240 (N_23240,N_20045,N_21160);
or U23241 (N_23241,N_20535,N_21411);
xor U23242 (N_23242,N_20683,N_21903);
or U23243 (N_23243,N_21082,N_20858);
nor U23244 (N_23244,N_21158,N_21358);
xor U23245 (N_23245,N_20563,N_20776);
and U23246 (N_23246,N_20672,N_21401);
nor U23247 (N_23247,N_21801,N_20139);
xnor U23248 (N_23248,N_21187,N_20425);
nor U23249 (N_23249,N_20036,N_21704);
nand U23250 (N_23250,N_21197,N_20200);
xor U23251 (N_23251,N_21571,N_20558);
or U23252 (N_23252,N_20962,N_21056);
nor U23253 (N_23253,N_21283,N_21862);
and U23254 (N_23254,N_21613,N_20679);
nand U23255 (N_23255,N_21141,N_20116);
xor U23256 (N_23256,N_20827,N_21428);
and U23257 (N_23257,N_20872,N_20814);
or U23258 (N_23258,N_20861,N_20363);
nor U23259 (N_23259,N_21554,N_21931);
or U23260 (N_23260,N_21048,N_21761);
xor U23261 (N_23261,N_20568,N_20737);
or U23262 (N_23262,N_20099,N_21993);
nor U23263 (N_23263,N_20301,N_20066);
and U23264 (N_23264,N_20947,N_21316);
xor U23265 (N_23265,N_21404,N_21122);
and U23266 (N_23266,N_20173,N_20051);
xnor U23267 (N_23267,N_20920,N_20037);
and U23268 (N_23268,N_21433,N_20841);
xnor U23269 (N_23269,N_20958,N_21069);
xor U23270 (N_23270,N_21090,N_20694);
nand U23271 (N_23271,N_21971,N_21973);
xnor U23272 (N_23272,N_20476,N_21876);
nand U23273 (N_23273,N_20494,N_20923);
nor U23274 (N_23274,N_20062,N_21951);
and U23275 (N_23275,N_21478,N_20931);
nor U23276 (N_23276,N_20238,N_20465);
nor U23277 (N_23277,N_20776,N_20905);
nor U23278 (N_23278,N_21216,N_20835);
nand U23279 (N_23279,N_21273,N_20927);
or U23280 (N_23280,N_20123,N_21678);
nor U23281 (N_23281,N_20294,N_20445);
or U23282 (N_23282,N_20105,N_20799);
and U23283 (N_23283,N_21161,N_21697);
or U23284 (N_23284,N_20020,N_21582);
nand U23285 (N_23285,N_21660,N_21924);
nand U23286 (N_23286,N_20420,N_21395);
nand U23287 (N_23287,N_21445,N_21108);
and U23288 (N_23288,N_21836,N_20653);
xor U23289 (N_23289,N_21543,N_20918);
xor U23290 (N_23290,N_20274,N_21741);
nand U23291 (N_23291,N_20920,N_21446);
nand U23292 (N_23292,N_21039,N_21518);
or U23293 (N_23293,N_21452,N_21094);
nand U23294 (N_23294,N_20815,N_20004);
nand U23295 (N_23295,N_20378,N_20428);
xnor U23296 (N_23296,N_21670,N_21788);
nor U23297 (N_23297,N_21711,N_20341);
xnor U23298 (N_23298,N_21956,N_20610);
and U23299 (N_23299,N_21495,N_21986);
and U23300 (N_23300,N_20478,N_21848);
or U23301 (N_23301,N_20700,N_20956);
nand U23302 (N_23302,N_21586,N_20265);
and U23303 (N_23303,N_21516,N_21919);
xor U23304 (N_23304,N_20894,N_21092);
xor U23305 (N_23305,N_21299,N_20641);
and U23306 (N_23306,N_21088,N_21497);
or U23307 (N_23307,N_21190,N_20696);
nor U23308 (N_23308,N_20076,N_20588);
nor U23309 (N_23309,N_20438,N_21684);
and U23310 (N_23310,N_20230,N_20983);
and U23311 (N_23311,N_21148,N_21957);
or U23312 (N_23312,N_21849,N_20731);
xor U23313 (N_23313,N_20244,N_21967);
nand U23314 (N_23314,N_20865,N_20298);
nand U23315 (N_23315,N_20931,N_20732);
or U23316 (N_23316,N_21256,N_21129);
xnor U23317 (N_23317,N_21298,N_20928);
nor U23318 (N_23318,N_20183,N_21079);
xnor U23319 (N_23319,N_21514,N_20856);
nand U23320 (N_23320,N_21964,N_20165);
xor U23321 (N_23321,N_20702,N_20173);
and U23322 (N_23322,N_20467,N_20279);
or U23323 (N_23323,N_21014,N_21892);
xnor U23324 (N_23324,N_21918,N_21959);
nor U23325 (N_23325,N_20040,N_21941);
and U23326 (N_23326,N_21353,N_21965);
xor U23327 (N_23327,N_21335,N_20741);
nand U23328 (N_23328,N_21470,N_20742);
and U23329 (N_23329,N_21792,N_21113);
nor U23330 (N_23330,N_20513,N_21760);
or U23331 (N_23331,N_21781,N_20521);
or U23332 (N_23332,N_20477,N_21052);
or U23333 (N_23333,N_20308,N_21523);
and U23334 (N_23334,N_21160,N_20872);
or U23335 (N_23335,N_20146,N_20488);
and U23336 (N_23336,N_20579,N_21759);
nand U23337 (N_23337,N_20144,N_20052);
xor U23338 (N_23338,N_21977,N_21876);
nand U23339 (N_23339,N_20630,N_20916);
and U23340 (N_23340,N_21328,N_20012);
nand U23341 (N_23341,N_21855,N_21573);
xor U23342 (N_23342,N_20251,N_20575);
or U23343 (N_23343,N_21655,N_21013);
nand U23344 (N_23344,N_20751,N_20311);
and U23345 (N_23345,N_20512,N_21442);
nand U23346 (N_23346,N_21505,N_20397);
nand U23347 (N_23347,N_21140,N_21045);
and U23348 (N_23348,N_20931,N_20925);
or U23349 (N_23349,N_21583,N_21869);
xnor U23350 (N_23350,N_20037,N_20003);
xor U23351 (N_23351,N_20482,N_20862);
nor U23352 (N_23352,N_21470,N_21496);
xor U23353 (N_23353,N_20759,N_20967);
nand U23354 (N_23354,N_20461,N_21016);
nor U23355 (N_23355,N_20310,N_20441);
and U23356 (N_23356,N_21264,N_21270);
or U23357 (N_23357,N_20315,N_21994);
nor U23358 (N_23358,N_20899,N_20020);
and U23359 (N_23359,N_21755,N_21654);
and U23360 (N_23360,N_20477,N_20309);
and U23361 (N_23361,N_21245,N_20800);
and U23362 (N_23362,N_20139,N_21661);
nand U23363 (N_23363,N_21501,N_21979);
xnor U23364 (N_23364,N_21560,N_21747);
nand U23365 (N_23365,N_21682,N_20966);
and U23366 (N_23366,N_20878,N_20254);
nand U23367 (N_23367,N_20481,N_21681);
and U23368 (N_23368,N_20337,N_21927);
nor U23369 (N_23369,N_20561,N_20806);
and U23370 (N_23370,N_21779,N_21133);
nand U23371 (N_23371,N_20966,N_21338);
and U23372 (N_23372,N_20079,N_20884);
and U23373 (N_23373,N_20450,N_21096);
nand U23374 (N_23374,N_20781,N_20584);
and U23375 (N_23375,N_21657,N_21561);
and U23376 (N_23376,N_20242,N_21881);
and U23377 (N_23377,N_21921,N_20797);
or U23378 (N_23378,N_20322,N_21140);
nor U23379 (N_23379,N_21845,N_20764);
or U23380 (N_23380,N_21142,N_20823);
nor U23381 (N_23381,N_21591,N_20472);
or U23382 (N_23382,N_21617,N_21950);
and U23383 (N_23383,N_20885,N_20069);
or U23384 (N_23384,N_21577,N_20424);
nor U23385 (N_23385,N_21707,N_21735);
nor U23386 (N_23386,N_20401,N_21968);
xnor U23387 (N_23387,N_20956,N_21306);
xor U23388 (N_23388,N_21017,N_21423);
nand U23389 (N_23389,N_21174,N_20817);
and U23390 (N_23390,N_20263,N_21774);
or U23391 (N_23391,N_20614,N_21828);
xor U23392 (N_23392,N_21127,N_20411);
nand U23393 (N_23393,N_20774,N_20043);
and U23394 (N_23394,N_21731,N_20937);
xnor U23395 (N_23395,N_21849,N_20003);
nand U23396 (N_23396,N_21501,N_21532);
xor U23397 (N_23397,N_20222,N_20096);
xor U23398 (N_23398,N_21251,N_20437);
or U23399 (N_23399,N_20009,N_20843);
and U23400 (N_23400,N_20929,N_21890);
xnor U23401 (N_23401,N_20002,N_21180);
or U23402 (N_23402,N_20954,N_20443);
nand U23403 (N_23403,N_21909,N_20511);
or U23404 (N_23404,N_20334,N_21310);
xor U23405 (N_23405,N_21478,N_20801);
nor U23406 (N_23406,N_21909,N_20015);
nand U23407 (N_23407,N_21507,N_21151);
nand U23408 (N_23408,N_21753,N_20764);
xor U23409 (N_23409,N_20258,N_21467);
or U23410 (N_23410,N_20952,N_21624);
or U23411 (N_23411,N_21454,N_21394);
or U23412 (N_23412,N_21177,N_20357);
or U23413 (N_23413,N_20184,N_21408);
and U23414 (N_23414,N_20361,N_21998);
and U23415 (N_23415,N_21091,N_21168);
nor U23416 (N_23416,N_21264,N_20984);
nand U23417 (N_23417,N_21304,N_20475);
xnor U23418 (N_23418,N_21324,N_20619);
nor U23419 (N_23419,N_21043,N_21358);
xnor U23420 (N_23420,N_20525,N_21036);
and U23421 (N_23421,N_20297,N_21560);
nand U23422 (N_23422,N_20842,N_21160);
xor U23423 (N_23423,N_21789,N_20307);
nand U23424 (N_23424,N_20197,N_20093);
or U23425 (N_23425,N_20964,N_21270);
nand U23426 (N_23426,N_20916,N_21293);
and U23427 (N_23427,N_21191,N_21671);
xor U23428 (N_23428,N_21702,N_21636);
or U23429 (N_23429,N_20003,N_20329);
nor U23430 (N_23430,N_20453,N_20425);
or U23431 (N_23431,N_21190,N_20311);
xnor U23432 (N_23432,N_21026,N_20833);
xnor U23433 (N_23433,N_21132,N_21305);
xnor U23434 (N_23434,N_21830,N_21925);
nor U23435 (N_23435,N_20632,N_20522);
nor U23436 (N_23436,N_20801,N_20155);
or U23437 (N_23437,N_20945,N_20268);
nand U23438 (N_23438,N_21034,N_20911);
nand U23439 (N_23439,N_20533,N_21983);
or U23440 (N_23440,N_21772,N_20733);
or U23441 (N_23441,N_20684,N_21891);
and U23442 (N_23442,N_20545,N_21909);
nand U23443 (N_23443,N_20304,N_20275);
xor U23444 (N_23444,N_21656,N_21784);
or U23445 (N_23445,N_20421,N_20214);
nand U23446 (N_23446,N_21148,N_21627);
nor U23447 (N_23447,N_20646,N_21011);
nor U23448 (N_23448,N_20324,N_20826);
or U23449 (N_23449,N_20055,N_20802);
or U23450 (N_23450,N_20683,N_20543);
or U23451 (N_23451,N_20290,N_21050);
xor U23452 (N_23452,N_20213,N_21051);
nand U23453 (N_23453,N_21026,N_21313);
xor U23454 (N_23454,N_20413,N_21825);
xor U23455 (N_23455,N_21040,N_21125);
and U23456 (N_23456,N_21036,N_20806);
or U23457 (N_23457,N_21178,N_21108);
nor U23458 (N_23458,N_21614,N_20551);
or U23459 (N_23459,N_21191,N_21498);
xnor U23460 (N_23460,N_21680,N_21912);
nand U23461 (N_23461,N_21602,N_21014);
and U23462 (N_23462,N_21619,N_20329);
nand U23463 (N_23463,N_21574,N_20185);
xor U23464 (N_23464,N_20810,N_21522);
nor U23465 (N_23465,N_21268,N_20469);
xor U23466 (N_23466,N_21296,N_20401);
or U23467 (N_23467,N_21500,N_21055);
nor U23468 (N_23468,N_20128,N_20941);
xnor U23469 (N_23469,N_20787,N_21028);
nand U23470 (N_23470,N_20518,N_20040);
and U23471 (N_23471,N_20970,N_21141);
or U23472 (N_23472,N_21041,N_21872);
nor U23473 (N_23473,N_20024,N_20754);
or U23474 (N_23474,N_20710,N_21888);
and U23475 (N_23475,N_21045,N_20469);
nor U23476 (N_23476,N_21863,N_21731);
nor U23477 (N_23477,N_20010,N_21270);
or U23478 (N_23478,N_21977,N_20435);
nand U23479 (N_23479,N_21896,N_20267);
nor U23480 (N_23480,N_20522,N_20719);
and U23481 (N_23481,N_20135,N_20907);
and U23482 (N_23482,N_20749,N_21392);
nand U23483 (N_23483,N_21474,N_20736);
xor U23484 (N_23484,N_21463,N_20646);
nand U23485 (N_23485,N_20774,N_21782);
and U23486 (N_23486,N_20150,N_21868);
xor U23487 (N_23487,N_21327,N_20588);
nor U23488 (N_23488,N_21119,N_21570);
nor U23489 (N_23489,N_21051,N_20078);
xnor U23490 (N_23490,N_20550,N_21602);
or U23491 (N_23491,N_21634,N_20631);
and U23492 (N_23492,N_21850,N_21990);
nor U23493 (N_23493,N_21167,N_20293);
and U23494 (N_23494,N_21747,N_20557);
xor U23495 (N_23495,N_20858,N_20309);
nand U23496 (N_23496,N_21300,N_21425);
xnor U23497 (N_23497,N_20097,N_20769);
xnor U23498 (N_23498,N_21497,N_21016);
or U23499 (N_23499,N_21654,N_20340);
xnor U23500 (N_23500,N_21511,N_21202);
nand U23501 (N_23501,N_20954,N_21538);
nor U23502 (N_23502,N_20806,N_20829);
or U23503 (N_23503,N_20494,N_20684);
and U23504 (N_23504,N_21915,N_21541);
and U23505 (N_23505,N_21690,N_20952);
or U23506 (N_23506,N_20515,N_21197);
xnor U23507 (N_23507,N_20264,N_21866);
or U23508 (N_23508,N_21120,N_20452);
and U23509 (N_23509,N_20113,N_21102);
nor U23510 (N_23510,N_21692,N_20169);
or U23511 (N_23511,N_21688,N_20932);
or U23512 (N_23512,N_21094,N_21586);
or U23513 (N_23513,N_20021,N_20441);
nor U23514 (N_23514,N_21794,N_20501);
xnor U23515 (N_23515,N_20664,N_20902);
nor U23516 (N_23516,N_20803,N_21606);
xor U23517 (N_23517,N_20348,N_20376);
and U23518 (N_23518,N_20868,N_21011);
nor U23519 (N_23519,N_20569,N_20232);
nor U23520 (N_23520,N_20222,N_20863);
nand U23521 (N_23521,N_20624,N_21190);
nand U23522 (N_23522,N_21099,N_21141);
nor U23523 (N_23523,N_20323,N_21731);
xor U23524 (N_23524,N_21124,N_20095);
and U23525 (N_23525,N_20964,N_21020);
or U23526 (N_23526,N_20545,N_21740);
nor U23527 (N_23527,N_20523,N_20567);
and U23528 (N_23528,N_20484,N_20573);
and U23529 (N_23529,N_21777,N_21543);
nand U23530 (N_23530,N_21331,N_20808);
and U23531 (N_23531,N_21578,N_21699);
nor U23532 (N_23532,N_20152,N_21752);
nand U23533 (N_23533,N_20211,N_20783);
nor U23534 (N_23534,N_20030,N_21279);
nand U23535 (N_23535,N_20575,N_21702);
xor U23536 (N_23536,N_21741,N_20899);
nor U23537 (N_23537,N_20319,N_20362);
and U23538 (N_23538,N_20183,N_20066);
nand U23539 (N_23539,N_20359,N_21692);
nor U23540 (N_23540,N_21173,N_20489);
or U23541 (N_23541,N_20496,N_20143);
nand U23542 (N_23542,N_20702,N_21118);
and U23543 (N_23543,N_20237,N_21992);
xor U23544 (N_23544,N_21891,N_21061);
or U23545 (N_23545,N_20887,N_20410);
and U23546 (N_23546,N_21099,N_21542);
nand U23547 (N_23547,N_20371,N_21995);
nor U23548 (N_23548,N_21576,N_21154);
and U23549 (N_23549,N_21831,N_21511);
nand U23550 (N_23550,N_20002,N_20013);
and U23551 (N_23551,N_21678,N_21164);
nor U23552 (N_23552,N_20046,N_21302);
xor U23553 (N_23553,N_20897,N_20998);
nand U23554 (N_23554,N_21055,N_21694);
or U23555 (N_23555,N_21296,N_20587);
xor U23556 (N_23556,N_21535,N_20526);
and U23557 (N_23557,N_21078,N_20760);
or U23558 (N_23558,N_20064,N_20103);
nor U23559 (N_23559,N_21133,N_20192);
or U23560 (N_23560,N_21088,N_21146);
xor U23561 (N_23561,N_21690,N_21851);
and U23562 (N_23562,N_21409,N_20898);
and U23563 (N_23563,N_21670,N_20999);
or U23564 (N_23564,N_20891,N_20500);
or U23565 (N_23565,N_21089,N_20747);
and U23566 (N_23566,N_21604,N_20848);
or U23567 (N_23567,N_21958,N_20897);
nor U23568 (N_23568,N_21420,N_20784);
and U23569 (N_23569,N_21657,N_21239);
xor U23570 (N_23570,N_21296,N_21282);
or U23571 (N_23571,N_20501,N_21260);
and U23572 (N_23572,N_21002,N_21311);
nor U23573 (N_23573,N_20528,N_20444);
or U23574 (N_23574,N_21405,N_20035);
nand U23575 (N_23575,N_21086,N_21084);
nor U23576 (N_23576,N_20527,N_20154);
nand U23577 (N_23577,N_21566,N_20775);
and U23578 (N_23578,N_20004,N_21423);
nand U23579 (N_23579,N_21295,N_20699);
or U23580 (N_23580,N_21593,N_20339);
and U23581 (N_23581,N_20098,N_21747);
or U23582 (N_23582,N_20604,N_21739);
or U23583 (N_23583,N_21024,N_20146);
and U23584 (N_23584,N_21027,N_21457);
xnor U23585 (N_23585,N_21137,N_20297);
and U23586 (N_23586,N_20780,N_21455);
nor U23587 (N_23587,N_21906,N_21007);
nor U23588 (N_23588,N_21204,N_20355);
nand U23589 (N_23589,N_20582,N_21443);
or U23590 (N_23590,N_21386,N_20810);
nand U23591 (N_23591,N_21987,N_21799);
and U23592 (N_23592,N_20125,N_21661);
and U23593 (N_23593,N_21823,N_21672);
nand U23594 (N_23594,N_20969,N_21698);
or U23595 (N_23595,N_20369,N_20881);
and U23596 (N_23596,N_21178,N_21103);
nand U23597 (N_23597,N_21805,N_21992);
nand U23598 (N_23598,N_21854,N_21489);
or U23599 (N_23599,N_20070,N_20301);
nor U23600 (N_23600,N_20074,N_21629);
nor U23601 (N_23601,N_20739,N_20719);
nor U23602 (N_23602,N_21929,N_21168);
nand U23603 (N_23603,N_20807,N_21317);
and U23604 (N_23604,N_21616,N_21257);
and U23605 (N_23605,N_21041,N_20672);
xnor U23606 (N_23606,N_20016,N_21155);
xor U23607 (N_23607,N_20690,N_21512);
or U23608 (N_23608,N_20436,N_20001);
nor U23609 (N_23609,N_20403,N_21945);
and U23610 (N_23610,N_21167,N_21517);
nand U23611 (N_23611,N_20324,N_21172);
nand U23612 (N_23612,N_20519,N_21023);
or U23613 (N_23613,N_20417,N_20036);
and U23614 (N_23614,N_20205,N_21003);
nor U23615 (N_23615,N_20559,N_21994);
xnor U23616 (N_23616,N_21482,N_21234);
nor U23617 (N_23617,N_20067,N_21818);
and U23618 (N_23618,N_21904,N_21372);
or U23619 (N_23619,N_21191,N_21209);
nand U23620 (N_23620,N_20278,N_21687);
nor U23621 (N_23621,N_21250,N_20196);
xor U23622 (N_23622,N_20567,N_21260);
and U23623 (N_23623,N_21360,N_21145);
or U23624 (N_23624,N_20175,N_20790);
nor U23625 (N_23625,N_20477,N_21290);
nand U23626 (N_23626,N_21293,N_21388);
and U23627 (N_23627,N_21292,N_20039);
or U23628 (N_23628,N_20280,N_21331);
nand U23629 (N_23629,N_20228,N_21163);
or U23630 (N_23630,N_21048,N_20277);
or U23631 (N_23631,N_20232,N_20067);
xor U23632 (N_23632,N_20225,N_21143);
or U23633 (N_23633,N_21032,N_21808);
xor U23634 (N_23634,N_20752,N_20744);
nand U23635 (N_23635,N_20178,N_20327);
nor U23636 (N_23636,N_21346,N_21603);
xnor U23637 (N_23637,N_20802,N_21824);
xor U23638 (N_23638,N_20516,N_20649);
xor U23639 (N_23639,N_20401,N_21280);
xnor U23640 (N_23640,N_20213,N_21571);
nor U23641 (N_23641,N_20549,N_20137);
nor U23642 (N_23642,N_20920,N_20617);
and U23643 (N_23643,N_20844,N_20427);
nor U23644 (N_23644,N_21904,N_21097);
nand U23645 (N_23645,N_21052,N_20828);
and U23646 (N_23646,N_20733,N_21836);
nand U23647 (N_23647,N_21900,N_20092);
nor U23648 (N_23648,N_21985,N_20949);
nand U23649 (N_23649,N_20286,N_21837);
or U23650 (N_23650,N_21659,N_20023);
xnor U23651 (N_23651,N_20630,N_20709);
and U23652 (N_23652,N_20472,N_21670);
nor U23653 (N_23653,N_20052,N_20232);
xnor U23654 (N_23654,N_21530,N_21152);
xnor U23655 (N_23655,N_20626,N_20731);
xor U23656 (N_23656,N_20485,N_20377);
nand U23657 (N_23657,N_21900,N_20519);
xor U23658 (N_23658,N_20036,N_20093);
and U23659 (N_23659,N_20230,N_21915);
or U23660 (N_23660,N_20920,N_21001);
and U23661 (N_23661,N_20169,N_21629);
or U23662 (N_23662,N_20035,N_21779);
nor U23663 (N_23663,N_20787,N_20283);
nand U23664 (N_23664,N_20364,N_21303);
or U23665 (N_23665,N_20643,N_21698);
nor U23666 (N_23666,N_21257,N_21474);
nor U23667 (N_23667,N_21358,N_21585);
and U23668 (N_23668,N_21578,N_20705);
nor U23669 (N_23669,N_20739,N_20945);
and U23670 (N_23670,N_21704,N_20925);
nor U23671 (N_23671,N_20143,N_20432);
xnor U23672 (N_23672,N_21959,N_20673);
xor U23673 (N_23673,N_20570,N_21975);
and U23674 (N_23674,N_20515,N_21478);
and U23675 (N_23675,N_21367,N_20004);
or U23676 (N_23676,N_20466,N_21764);
or U23677 (N_23677,N_21982,N_20564);
nand U23678 (N_23678,N_20033,N_20752);
xnor U23679 (N_23679,N_20689,N_20095);
nand U23680 (N_23680,N_21590,N_21970);
xor U23681 (N_23681,N_20991,N_21868);
xnor U23682 (N_23682,N_21489,N_21002);
nand U23683 (N_23683,N_20324,N_21136);
and U23684 (N_23684,N_20753,N_21351);
or U23685 (N_23685,N_20143,N_20469);
xnor U23686 (N_23686,N_21560,N_21654);
and U23687 (N_23687,N_21258,N_20717);
nor U23688 (N_23688,N_20907,N_20291);
nor U23689 (N_23689,N_20718,N_20013);
xor U23690 (N_23690,N_20284,N_20034);
nand U23691 (N_23691,N_21398,N_20564);
nand U23692 (N_23692,N_21077,N_21406);
nor U23693 (N_23693,N_20458,N_20766);
xnor U23694 (N_23694,N_20644,N_20259);
or U23695 (N_23695,N_21676,N_21800);
or U23696 (N_23696,N_21060,N_21663);
nor U23697 (N_23697,N_21678,N_20383);
nand U23698 (N_23698,N_21044,N_20537);
nor U23699 (N_23699,N_20596,N_20157);
and U23700 (N_23700,N_21942,N_21201);
nor U23701 (N_23701,N_21049,N_20122);
or U23702 (N_23702,N_21005,N_21206);
xor U23703 (N_23703,N_20243,N_21033);
nand U23704 (N_23704,N_20707,N_20447);
and U23705 (N_23705,N_20432,N_20875);
nand U23706 (N_23706,N_20950,N_21940);
or U23707 (N_23707,N_21658,N_20189);
nor U23708 (N_23708,N_20818,N_20850);
nand U23709 (N_23709,N_21092,N_20360);
nand U23710 (N_23710,N_20717,N_20484);
xnor U23711 (N_23711,N_21832,N_21501);
or U23712 (N_23712,N_21321,N_20553);
xor U23713 (N_23713,N_20050,N_21486);
nand U23714 (N_23714,N_21608,N_20867);
nor U23715 (N_23715,N_21962,N_20359);
nor U23716 (N_23716,N_21287,N_21551);
and U23717 (N_23717,N_21439,N_20636);
nand U23718 (N_23718,N_21830,N_21773);
or U23719 (N_23719,N_21412,N_21024);
nand U23720 (N_23720,N_20248,N_20695);
nand U23721 (N_23721,N_21213,N_21342);
or U23722 (N_23722,N_21754,N_21276);
or U23723 (N_23723,N_21828,N_21115);
nand U23724 (N_23724,N_21684,N_21254);
or U23725 (N_23725,N_21566,N_21298);
and U23726 (N_23726,N_21361,N_20630);
xnor U23727 (N_23727,N_20647,N_21498);
nand U23728 (N_23728,N_21192,N_20915);
or U23729 (N_23729,N_21426,N_20764);
xnor U23730 (N_23730,N_20977,N_20693);
nand U23731 (N_23731,N_20844,N_21857);
xor U23732 (N_23732,N_21465,N_21125);
nor U23733 (N_23733,N_21656,N_21337);
and U23734 (N_23734,N_21524,N_20534);
xnor U23735 (N_23735,N_20901,N_20303);
or U23736 (N_23736,N_21724,N_20576);
or U23737 (N_23737,N_20491,N_21635);
or U23738 (N_23738,N_21719,N_21404);
nor U23739 (N_23739,N_20961,N_20866);
and U23740 (N_23740,N_21439,N_20446);
or U23741 (N_23741,N_20418,N_21735);
or U23742 (N_23742,N_21905,N_21569);
nand U23743 (N_23743,N_20761,N_20089);
or U23744 (N_23744,N_21669,N_20930);
xnor U23745 (N_23745,N_21150,N_21102);
and U23746 (N_23746,N_21780,N_20140);
and U23747 (N_23747,N_21797,N_20960);
and U23748 (N_23748,N_21862,N_20350);
and U23749 (N_23749,N_21941,N_20215);
nand U23750 (N_23750,N_21988,N_21000);
nor U23751 (N_23751,N_21050,N_20997);
and U23752 (N_23752,N_21044,N_21445);
or U23753 (N_23753,N_21277,N_20316);
or U23754 (N_23754,N_21439,N_21676);
or U23755 (N_23755,N_20616,N_20046);
or U23756 (N_23756,N_20841,N_20609);
or U23757 (N_23757,N_21212,N_21481);
nor U23758 (N_23758,N_21756,N_20900);
or U23759 (N_23759,N_21868,N_20054);
or U23760 (N_23760,N_21639,N_20864);
xor U23761 (N_23761,N_20431,N_21297);
or U23762 (N_23762,N_20320,N_20099);
nor U23763 (N_23763,N_21482,N_20396);
or U23764 (N_23764,N_20835,N_20455);
or U23765 (N_23765,N_20278,N_20392);
or U23766 (N_23766,N_21002,N_20291);
or U23767 (N_23767,N_20068,N_21856);
or U23768 (N_23768,N_21128,N_21643);
xor U23769 (N_23769,N_21586,N_21539);
and U23770 (N_23770,N_21769,N_20328);
nor U23771 (N_23771,N_20260,N_20732);
and U23772 (N_23772,N_20812,N_21400);
or U23773 (N_23773,N_20622,N_21740);
nand U23774 (N_23774,N_20212,N_21041);
nor U23775 (N_23775,N_20784,N_21766);
xor U23776 (N_23776,N_20315,N_21292);
and U23777 (N_23777,N_20640,N_21322);
or U23778 (N_23778,N_20818,N_20123);
xor U23779 (N_23779,N_20706,N_21022);
xnor U23780 (N_23780,N_21263,N_20535);
and U23781 (N_23781,N_21157,N_21809);
xnor U23782 (N_23782,N_21664,N_20435);
xnor U23783 (N_23783,N_20633,N_21093);
xnor U23784 (N_23784,N_21524,N_21268);
or U23785 (N_23785,N_20547,N_21453);
xnor U23786 (N_23786,N_21992,N_20111);
nor U23787 (N_23787,N_20179,N_21042);
and U23788 (N_23788,N_20217,N_20917);
and U23789 (N_23789,N_21322,N_21386);
or U23790 (N_23790,N_21478,N_20351);
xor U23791 (N_23791,N_20698,N_20503);
xor U23792 (N_23792,N_20051,N_21900);
xor U23793 (N_23793,N_21862,N_20030);
and U23794 (N_23794,N_20503,N_20828);
nand U23795 (N_23795,N_21448,N_21823);
or U23796 (N_23796,N_20984,N_20352);
nand U23797 (N_23797,N_21497,N_20631);
nor U23798 (N_23798,N_20642,N_20623);
nand U23799 (N_23799,N_20445,N_21579);
xor U23800 (N_23800,N_20881,N_21509);
or U23801 (N_23801,N_21607,N_20365);
and U23802 (N_23802,N_20348,N_21581);
and U23803 (N_23803,N_21285,N_21590);
nor U23804 (N_23804,N_21767,N_20258);
or U23805 (N_23805,N_20662,N_20750);
and U23806 (N_23806,N_20223,N_21454);
or U23807 (N_23807,N_20065,N_20535);
or U23808 (N_23808,N_20348,N_21742);
or U23809 (N_23809,N_21791,N_20277);
or U23810 (N_23810,N_20738,N_20007);
or U23811 (N_23811,N_21223,N_20817);
xor U23812 (N_23812,N_21312,N_20083);
xor U23813 (N_23813,N_21735,N_21791);
nor U23814 (N_23814,N_21182,N_21329);
xor U23815 (N_23815,N_21006,N_21466);
nand U23816 (N_23816,N_21496,N_21999);
nand U23817 (N_23817,N_21677,N_21142);
nand U23818 (N_23818,N_21844,N_21959);
nor U23819 (N_23819,N_21253,N_20591);
nor U23820 (N_23820,N_20305,N_20018);
nand U23821 (N_23821,N_20166,N_20808);
xor U23822 (N_23822,N_21021,N_20272);
or U23823 (N_23823,N_20945,N_20914);
and U23824 (N_23824,N_21725,N_20837);
or U23825 (N_23825,N_20809,N_20464);
xnor U23826 (N_23826,N_20250,N_20411);
or U23827 (N_23827,N_21098,N_21115);
nand U23828 (N_23828,N_20041,N_20337);
xnor U23829 (N_23829,N_20045,N_20783);
xnor U23830 (N_23830,N_21682,N_21060);
and U23831 (N_23831,N_20949,N_21837);
or U23832 (N_23832,N_20832,N_20478);
xnor U23833 (N_23833,N_21956,N_21530);
nand U23834 (N_23834,N_21923,N_21753);
and U23835 (N_23835,N_20201,N_20217);
nand U23836 (N_23836,N_20248,N_21513);
and U23837 (N_23837,N_21773,N_21035);
and U23838 (N_23838,N_21198,N_21463);
xor U23839 (N_23839,N_21807,N_21598);
or U23840 (N_23840,N_20238,N_21582);
nor U23841 (N_23841,N_20539,N_20680);
xor U23842 (N_23842,N_20220,N_20980);
nand U23843 (N_23843,N_20072,N_21053);
nor U23844 (N_23844,N_21062,N_21978);
nand U23845 (N_23845,N_20840,N_21994);
and U23846 (N_23846,N_20653,N_20337);
and U23847 (N_23847,N_20095,N_21863);
or U23848 (N_23848,N_20337,N_20807);
xnor U23849 (N_23849,N_21118,N_21024);
xnor U23850 (N_23850,N_21173,N_21734);
or U23851 (N_23851,N_21401,N_20516);
and U23852 (N_23852,N_21004,N_21911);
nand U23853 (N_23853,N_21342,N_21932);
nor U23854 (N_23854,N_21337,N_20922);
nand U23855 (N_23855,N_20451,N_21532);
nand U23856 (N_23856,N_21379,N_20440);
xor U23857 (N_23857,N_21423,N_21159);
and U23858 (N_23858,N_20090,N_20178);
nand U23859 (N_23859,N_20866,N_20024);
or U23860 (N_23860,N_20956,N_20099);
nand U23861 (N_23861,N_20890,N_20679);
nor U23862 (N_23862,N_20435,N_20274);
or U23863 (N_23863,N_20956,N_20756);
nand U23864 (N_23864,N_20776,N_20087);
or U23865 (N_23865,N_21711,N_21245);
nor U23866 (N_23866,N_21539,N_20874);
xnor U23867 (N_23867,N_21370,N_20210);
or U23868 (N_23868,N_21632,N_20781);
xnor U23869 (N_23869,N_21400,N_21605);
nor U23870 (N_23870,N_21276,N_21534);
or U23871 (N_23871,N_20764,N_20119);
xnor U23872 (N_23872,N_21082,N_20638);
xnor U23873 (N_23873,N_21555,N_21283);
nor U23874 (N_23874,N_21041,N_20313);
nor U23875 (N_23875,N_21127,N_20634);
nand U23876 (N_23876,N_21174,N_20552);
or U23877 (N_23877,N_21773,N_20838);
or U23878 (N_23878,N_20426,N_20388);
xor U23879 (N_23879,N_21154,N_21289);
nor U23880 (N_23880,N_20310,N_20642);
nor U23881 (N_23881,N_21585,N_20932);
nand U23882 (N_23882,N_21521,N_21123);
nand U23883 (N_23883,N_21764,N_20045);
nand U23884 (N_23884,N_21160,N_21618);
nor U23885 (N_23885,N_21876,N_20117);
nor U23886 (N_23886,N_21182,N_20104);
and U23887 (N_23887,N_20684,N_21784);
or U23888 (N_23888,N_20332,N_20594);
xor U23889 (N_23889,N_20973,N_20369);
nor U23890 (N_23890,N_20398,N_20252);
and U23891 (N_23891,N_21425,N_20496);
nor U23892 (N_23892,N_21351,N_21072);
or U23893 (N_23893,N_20171,N_21044);
xnor U23894 (N_23894,N_20070,N_20811);
nor U23895 (N_23895,N_21424,N_21391);
xor U23896 (N_23896,N_21435,N_20103);
nor U23897 (N_23897,N_21854,N_20098);
nor U23898 (N_23898,N_20606,N_21267);
and U23899 (N_23899,N_21354,N_21580);
or U23900 (N_23900,N_20080,N_20444);
xnor U23901 (N_23901,N_21104,N_20912);
and U23902 (N_23902,N_21505,N_21255);
nor U23903 (N_23903,N_21810,N_21138);
nand U23904 (N_23904,N_20986,N_20052);
nand U23905 (N_23905,N_21281,N_21180);
nor U23906 (N_23906,N_20053,N_21036);
or U23907 (N_23907,N_21528,N_21865);
or U23908 (N_23908,N_20550,N_20338);
nand U23909 (N_23909,N_20501,N_21286);
and U23910 (N_23910,N_20259,N_20253);
nand U23911 (N_23911,N_20976,N_21444);
and U23912 (N_23912,N_20115,N_21154);
nand U23913 (N_23913,N_21855,N_20790);
nor U23914 (N_23914,N_21549,N_20540);
xnor U23915 (N_23915,N_20717,N_20136);
xor U23916 (N_23916,N_20367,N_21359);
nor U23917 (N_23917,N_20600,N_20588);
or U23918 (N_23918,N_20817,N_20328);
or U23919 (N_23919,N_20826,N_20277);
nand U23920 (N_23920,N_21544,N_21519);
nand U23921 (N_23921,N_20278,N_20359);
nand U23922 (N_23922,N_21155,N_20488);
or U23923 (N_23923,N_20152,N_20647);
xor U23924 (N_23924,N_21744,N_20211);
xnor U23925 (N_23925,N_20330,N_20183);
or U23926 (N_23926,N_21112,N_21332);
nand U23927 (N_23927,N_20992,N_20886);
xor U23928 (N_23928,N_20600,N_21305);
nor U23929 (N_23929,N_21832,N_21881);
nor U23930 (N_23930,N_21937,N_20463);
or U23931 (N_23931,N_20856,N_20171);
nor U23932 (N_23932,N_20673,N_21360);
and U23933 (N_23933,N_21910,N_20098);
and U23934 (N_23934,N_21228,N_20760);
xor U23935 (N_23935,N_21948,N_21299);
and U23936 (N_23936,N_21178,N_20949);
xor U23937 (N_23937,N_20830,N_21439);
nand U23938 (N_23938,N_21617,N_21165);
or U23939 (N_23939,N_21587,N_20225);
xnor U23940 (N_23940,N_20359,N_21874);
or U23941 (N_23941,N_21591,N_21283);
or U23942 (N_23942,N_20532,N_20005);
xnor U23943 (N_23943,N_21127,N_20547);
nand U23944 (N_23944,N_20812,N_21016);
nor U23945 (N_23945,N_20254,N_20297);
and U23946 (N_23946,N_21514,N_21200);
nand U23947 (N_23947,N_21068,N_20740);
and U23948 (N_23948,N_20005,N_21026);
nand U23949 (N_23949,N_21648,N_20154);
nor U23950 (N_23950,N_21620,N_21584);
nor U23951 (N_23951,N_21292,N_21611);
xnor U23952 (N_23952,N_21256,N_20372);
nor U23953 (N_23953,N_21316,N_21979);
and U23954 (N_23954,N_20174,N_21674);
xnor U23955 (N_23955,N_21234,N_20167);
xnor U23956 (N_23956,N_21021,N_20971);
xnor U23957 (N_23957,N_21250,N_20138);
xnor U23958 (N_23958,N_21057,N_20128);
nand U23959 (N_23959,N_21142,N_21552);
nand U23960 (N_23960,N_20365,N_20460);
nor U23961 (N_23961,N_20142,N_20655);
nand U23962 (N_23962,N_20396,N_20773);
or U23963 (N_23963,N_21540,N_21130);
or U23964 (N_23964,N_21089,N_20380);
xnor U23965 (N_23965,N_21914,N_20617);
nand U23966 (N_23966,N_21602,N_20294);
and U23967 (N_23967,N_21345,N_21865);
and U23968 (N_23968,N_21464,N_21389);
or U23969 (N_23969,N_20275,N_21828);
xor U23970 (N_23970,N_20375,N_21981);
xnor U23971 (N_23971,N_21284,N_21374);
nand U23972 (N_23972,N_20389,N_21923);
xor U23973 (N_23973,N_21413,N_20088);
or U23974 (N_23974,N_20245,N_20879);
nand U23975 (N_23975,N_21131,N_20279);
nand U23976 (N_23976,N_20072,N_20381);
nor U23977 (N_23977,N_21723,N_21664);
and U23978 (N_23978,N_20924,N_21982);
nor U23979 (N_23979,N_20903,N_21590);
nand U23980 (N_23980,N_20461,N_20096);
or U23981 (N_23981,N_20460,N_21558);
and U23982 (N_23982,N_21871,N_21107);
nor U23983 (N_23983,N_20877,N_21368);
and U23984 (N_23984,N_20725,N_20169);
xor U23985 (N_23985,N_21050,N_20202);
xor U23986 (N_23986,N_20445,N_21962);
or U23987 (N_23987,N_21560,N_21187);
or U23988 (N_23988,N_21394,N_20685);
xnor U23989 (N_23989,N_20583,N_20041);
or U23990 (N_23990,N_20674,N_21365);
xor U23991 (N_23991,N_20877,N_20597);
nand U23992 (N_23992,N_21303,N_21464);
nor U23993 (N_23993,N_20562,N_20737);
and U23994 (N_23994,N_20388,N_21393);
nand U23995 (N_23995,N_20401,N_20282);
nand U23996 (N_23996,N_20141,N_21621);
xor U23997 (N_23997,N_21049,N_20022);
or U23998 (N_23998,N_20779,N_21151);
nor U23999 (N_23999,N_21053,N_20200);
xnor U24000 (N_24000,N_22450,N_22559);
xor U24001 (N_24001,N_22648,N_22519);
or U24002 (N_24002,N_23086,N_23771);
nor U24003 (N_24003,N_23661,N_22048);
xor U24004 (N_24004,N_22052,N_22100);
xnor U24005 (N_24005,N_23485,N_22161);
xnor U24006 (N_24006,N_23559,N_22879);
xor U24007 (N_24007,N_22901,N_22794);
nand U24008 (N_24008,N_23344,N_22872);
and U24009 (N_24009,N_23990,N_23563);
and U24010 (N_24010,N_23178,N_22711);
xor U24011 (N_24011,N_23573,N_23108);
xnor U24012 (N_24012,N_22061,N_22494);
or U24013 (N_24013,N_22859,N_23281);
or U24014 (N_24014,N_23273,N_23545);
nor U24015 (N_24015,N_22682,N_22707);
nor U24016 (N_24016,N_22316,N_23277);
nor U24017 (N_24017,N_22262,N_23495);
and U24018 (N_24018,N_23896,N_23535);
nand U24019 (N_24019,N_23246,N_23840);
xor U24020 (N_24020,N_23141,N_22999);
xnor U24021 (N_24021,N_23409,N_22149);
nand U24022 (N_24022,N_22558,N_22168);
xor U24023 (N_24023,N_22775,N_22728);
or U24024 (N_24024,N_23516,N_23911);
nand U24025 (N_24025,N_23403,N_23774);
and U24026 (N_24026,N_22851,N_22553);
or U24027 (N_24027,N_22715,N_23873);
xnor U24028 (N_24028,N_23493,N_22968);
xnor U24029 (N_24029,N_23947,N_22634);
xnor U24030 (N_24030,N_22352,N_23577);
and U24031 (N_24031,N_22001,N_22816);
xor U24032 (N_24032,N_22169,N_22643);
nor U24033 (N_24033,N_23011,N_22414);
nor U24034 (N_24034,N_22265,N_22752);
nor U24035 (N_24035,N_23604,N_23813);
nand U24036 (N_24036,N_23984,N_23471);
nand U24037 (N_24037,N_23490,N_23006);
nand U24038 (N_24038,N_23399,N_23404);
nor U24039 (N_24039,N_23855,N_22111);
nor U24040 (N_24040,N_23864,N_22259);
nand U24041 (N_24041,N_22943,N_22572);
or U24042 (N_24042,N_23870,N_22854);
nand U24043 (N_24043,N_22492,N_23743);
xor U24044 (N_24044,N_23118,N_23519);
or U24045 (N_24045,N_23486,N_22768);
nand U24046 (N_24046,N_23826,N_22633);
and U24047 (N_24047,N_22411,N_22759);
or U24048 (N_24048,N_23369,N_23009);
and U24049 (N_24049,N_22189,N_22490);
xor U24050 (N_24050,N_23394,N_22228);
xnor U24051 (N_24051,N_23123,N_23338);
nand U24052 (N_24052,N_22749,N_23662);
and U24053 (N_24053,N_22120,N_22764);
nand U24054 (N_24054,N_23373,N_23239);
nor U24055 (N_24055,N_23817,N_23620);
and U24056 (N_24056,N_23933,N_23885);
xnor U24057 (N_24057,N_22299,N_22125);
and U24058 (N_24058,N_22446,N_22580);
nand U24059 (N_24059,N_23260,N_22928);
nand U24060 (N_24060,N_23922,N_23224);
nor U24061 (N_24061,N_23455,N_23803);
or U24062 (N_24062,N_22871,N_22565);
nor U24063 (N_24063,N_22680,N_23214);
nor U24064 (N_24064,N_22221,N_23720);
and U24065 (N_24065,N_22391,N_22053);
xor U24066 (N_24066,N_22665,N_23003);
and U24067 (N_24067,N_22886,N_22146);
or U24068 (N_24068,N_23196,N_22119);
and U24069 (N_24069,N_22543,N_22307);
xnor U24070 (N_24070,N_22925,N_22908);
or U24071 (N_24071,N_22508,N_22724);
or U24072 (N_24072,N_22392,N_23127);
and U24073 (N_24073,N_22371,N_23790);
or U24074 (N_24074,N_22351,N_22166);
xnor U24075 (N_24075,N_22888,N_22012);
or U24076 (N_24076,N_23723,N_23905);
nand U24077 (N_24077,N_22095,N_23186);
or U24078 (N_24078,N_23469,N_22842);
nand U24079 (N_24079,N_22704,N_23606);
xor U24080 (N_24080,N_23657,N_22093);
and U24081 (N_24081,N_23320,N_22635);
nand U24082 (N_24082,N_22211,N_23555);
and U24083 (N_24083,N_23358,N_22255);
nor U24084 (N_24084,N_22133,N_23134);
and U24085 (N_24085,N_22396,N_23724);
and U24086 (N_24086,N_22062,N_22023);
or U24087 (N_24087,N_23703,N_22401);
nor U24088 (N_24088,N_23153,N_23889);
and U24089 (N_24089,N_23309,N_22485);
xnor U24090 (N_24090,N_22193,N_22548);
nor U24091 (N_24091,N_22876,N_23100);
xor U24092 (N_24092,N_22698,N_22660);
or U24093 (N_24093,N_23039,N_22757);
nand U24094 (N_24094,N_23090,N_23861);
and U24095 (N_24095,N_23388,N_23435);
nor U24096 (N_24096,N_23776,N_22128);
nor U24097 (N_24097,N_23036,N_22511);
xor U24098 (N_24098,N_23477,N_22388);
nor U24099 (N_24099,N_22448,N_22474);
and U24100 (N_24100,N_23700,N_22174);
and U24101 (N_24101,N_23684,N_23295);
and U24102 (N_24102,N_23801,N_22070);
xnor U24103 (N_24103,N_22393,N_23756);
nor U24104 (N_24104,N_22654,N_23151);
or U24105 (N_24105,N_22455,N_23888);
or U24106 (N_24106,N_22230,N_22240);
or U24107 (N_24107,N_22792,N_22071);
nand U24108 (N_24108,N_22186,N_23694);
nor U24109 (N_24109,N_22849,N_23385);
nor U24110 (N_24110,N_23744,N_23111);
nor U24111 (N_24111,N_22135,N_22719);
xnor U24112 (N_24112,N_22602,N_22845);
nor U24113 (N_24113,N_23112,N_22975);
nor U24114 (N_24114,N_22190,N_22147);
xor U24115 (N_24115,N_23307,N_22079);
nor U24116 (N_24116,N_22720,N_22250);
nor U24117 (N_24117,N_22829,N_22923);
or U24118 (N_24118,N_23441,N_23423);
xnor U24119 (N_24119,N_23007,N_23533);
nor U24120 (N_24120,N_23010,N_22955);
nor U24121 (N_24121,N_22693,N_23759);
or U24122 (N_24122,N_23074,N_23289);
xnor U24123 (N_24123,N_23585,N_23977);
and U24124 (N_24124,N_22131,N_22581);
or U24125 (N_24125,N_22356,N_22231);
nor U24126 (N_24126,N_23576,N_23414);
nand U24127 (N_24127,N_22824,N_23778);
nand U24128 (N_24128,N_22315,N_22463);
xor U24129 (N_24129,N_23627,N_22538);
or U24130 (N_24130,N_22285,N_22354);
xnor U24131 (N_24131,N_22458,N_23938);
and U24132 (N_24132,N_23245,N_22322);
nor U24133 (N_24133,N_23951,N_22932);
and U24134 (N_24134,N_22587,N_23242);
xor U24135 (N_24135,N_23386,N_23880);
nor U24136 (N_24136,N_22298,N_23649);
xnor U24137 (N_24137,N_23439,N_22853);
nand U24138 (N_24138,N_23753,N_23229);
or U24139 (N_24139,N_22279,N_22725);
and U24140 (N_24140,N_22033,N_23042);
nor U24141 (N_24141,N_23928,N_23955);
or U24142 (N_24142,N_23936,N_23702);
xnor U24143 (N_24143,N_23420,N_22954);
nand U24144 (N_24144,N_22054,N_22195);
and U24145 (N_24145,N_22020,N_23304);
xor U24146 (N_24146,N_23467,N_22547);
and U24147 (N_24147,N_23558,N_22469);
xnor U24148 (N_24148,N_22418,N_22918);
nor U24149 (N_24149,N_22308,N_23235);
and U24150 (N_24150,N_23874,N_23047);
and U24151 (N_24151,N_23209,N_23421);
nor U24152 (N_24152,N_22007,N_23590);
or U24153 (N_24153,N_22726,N_23676);
xor U24154 (N_24154,N_22838,N_23331);
nand U24155 (N_24155,N_23267,N_22087);
nor U24156 (N_24156,N_23542,N_23596);
or U24157 (N_24157,N_23809,N_23511);
nand U24158 (N_24158,N_23612,N_22456);
nor U24159 (N_24159,N_23482,N_22056);
xnor U24160 (N_24160,N_22422,N_23121);
nor U24161 (N_24161,N_23601,N_22609);
or U24162 (N_24162,N_22115,N_23664);
nor U24163 (N_24163,N_22475,N_23303);
or U24164 (N_24164,N_23243,N_22625);
nand U24165 (N_24165,N_22107,N_22554);
nand U24166 (N_24166,N_23540,N_22284);
xnor U24167 (N_24167,N_23712,N_23020);
or U24168 (N_24168,N_23730,N_23142);
nand U24169 (N_24169,N_22516,N_22869);
xor U24170 (N_24170,N_23089,N_23191);
xnor U24171 (N_24171,N_22751,N_23652);
and U24172 (N_24172,N_22357,N_23784);
nand U24173 (N_24173,N_22140,N_23155);
nor U24174 (N_24174,N_22342,N_22434);
nor U24175 (N_24175,N_22158,N_22772);
or U24176 (N_24176,N_22536,N_22065);
or U24177 (N_24177,N_23610,N_23937);
or U24178 (N_24178,N_22066,N_22767);
xor U24179 (N_24179,N_23122,N_23717);
xor U24180 (N_24180,N_23898,N_22611);
nor U24181 (N_24181,N_22616,N_23048);
or U24182 (N_24182,N_22394,N_22727);
or U24183 (N_24183,N_23237,N_22229);
xnor U24184 (N_24184,N_23363,N_23525);
or U24185 (N_24185,N_23301,N_23110);
and U24186 (N_24186,N_23865,N_23157);
nor U24187 (N_24187,N_22964,N_23146);
or U24188 (N_24188,N_23154,N_23337);
nor U24189 (N_24189,N_23981,N_23255);
nor U24190 (N_24190,N_23312,N_23250);
and U24191 (N_24191,N_23690,N_22561);
nor U24192 (N_24192,N_22883,N_23806);
xor U24193 (N_24193,N_22462,N_22958);
xor U24194 (N_24194,N_23568,N_23431);
and U24195 (N_24195,N_22527,N_22714);
xor U24196 (N_24196,N_22837,N_23881);
nor U24197 (N_24197,N_23629,N_22897);
nor U24198 (N_24198,N_22758,N_23740);
and U24199 (N_24199,N_23773,N_22591);
and U24200 (N_24200,N_23181,N_23859);
nor U24201 (N_24201,N_23893,N_22438);
nor U24202 (N_24202,N_23923,N_23707);
xnor U24203 (N_24203,N_22914,N_22468);
xnor U24204 (N_24204,N_22623,N_22436);
or U24205 (N_24205,N_22960,N_22971);
nand U24206 (N_24206,N_22427,N_23647);
or U24207 (N_24207,N_22787,N_22733);
and U24208 (N_24208,N_23314,N_22867);
or U24209 (N_24209,N_23347,N_22687);
and U24210 (N_24210,N_22919,N_22713);
nand U24211 (N_24211,N_22151,N_23689);
xnor U24212 (N_24212,N_22215,N_22953);
nand U24213 (N_24213,N_23241,N_23317);
xnor U24214 (N_24214,N_23588,N_22922);
nand U24215 (N_24215,N_22144,N_22477);
nand U24216 (N_24216,N_22185,N_22742);
xor U24217 (N_24217,N_22889,N_23547);
nand U24218 (N_24218,N_22563,N_23901);
xnor U24219 (N_24219,N_23491,N_22175);
or U24220 (N_24220,N_22806,N_23536);
nand U24221 (N_24221,N_22045,N_23965);
and U24222 (N_24222,N_23727,N_22425);
and U24223 (N_24223,N_22831,N_22799);
and U24224 (N_24224,N_23615,N_23549);
and U24225 (N_24225,N_22517,N_22604);
and U24226 (N_24226,N_22077,N_23244);
xnor U24227 (N_24227,N_22499,N_22570);
nor U24228 (N_24228,N_22786,N_22850);
and U24229 (N_24229,N_23838,N_22729);
nor U24230 (N_24230,N_22641,N_23436);
nor U24231 (N_24231,N_22302,N_23512);
nor U24232 (N_24232,N_23472,N_22597);
nand U24233 (N_24233,N_23634,N_23745);
nand U24234 (N_24234,N_22510,N_22176);
or U24235 (N_24235,N_22612,N_22376);
or U24236 (N_24236,N_22137,N_23132);
nor U24237 (N_24237,N_22046,N_22542);
nor U24238 (N_24238,N_23029,N_23302);
xor U24239 (N_24239,N_22333,N_23854);
nand U24240 (N_24240,N_23452,N_23973);
xnor U24241 (N_24241,N_23763,N_22060);
and U24242 (N_24242,N_23262,N_23742);
or U24243 (N_24243,N_23960,N_22945);
nor U24244 (N_24244,N_23150,N_22493);
nor U24245 (N_24245,N_23589,N_22472);
nand U24246 (N_24246,N_22762,N_22900);
nor U24247 (N_24247,N_22172,N_23383);
or U24248 (N_24248,N_22926,N_22246);
xnor U24249 (N_24249,N_22110,N_22607);
or U24250 (N_24250,N_23411,N_22970);
or U24251 (N_24251,N_22486,N_23135);
nand U24252 (N_24252,N_22270,N_23642);
xor U24253 (N_24253,N_22523,N_22802);
and U24254 (N_24254,N_22703,N_22619);
and U24255 (N_24255,N_22798,N_22473);
nor U24256 (N_24256,N_23197,N_23152);
nand U24257 (N_24257,N_23028,N_22873);
or U24258 (N_24258,N_23754,N_22747);
and U24259 (N_24259,N_22583,N_22086);
xnor U24260 (N_24260,N_22483,N_23192);
nor U24261 (N_24261,N_22142,N_23213);
nand U24262 (N_24262,N_22870,N_23942);
nor U24263 (N_24263,N_22721,N_23413);
nor U24264 (N_24264,N_23457,N_23719);
nor U24265 (N_24265,N_22470,N_23619);
xnor U24266 (N_24266,N_23269,N_22332);
nor U24267 (N_24267,N_23379,N_22946);
nor U24268 (N_24268,N_22575,N_22920);
xor U24269 (N_24269,N_22500,N_22909);
nor U24270 (N_24270,N_23376,N_23203);
xor U24271 (N_24271,N_22985,N_23749);
nand U24272 (N_24272,N_23909,N_23052);
xor U24273 (N_24273,N_22126,N_23043);
or U24274 (N_24274,N_23375,N_23367);
or U24275 (N_24275,N_23748,N_22301);
xor U24276 (N_24276,N_23480,N_23501);
and U24277 (N_24277,N_23699,N_22464);
nand U24278 (N_24278,N_23492,N_23066);
and U24279 (N_24279,N_22399,N_22323);
or U24280 (N_24280,N_23920,N_22044);
nand U24281 (N_24281,N_23296,N_23069);
xor U24282 (N_24282,N_23843,N_23024);
or U24283 (N_24283,N_23811,N_22717);
xor U24284 (N_24284,N_22360,N_23875);
nor U24285 (N_24285,N_23561,N_22991);
xor U24286 (N_24286,N_23603,N_23082);
nor U24287 (N_24287,N_23396,N_23232);
nand U24288 (N_24288,N_23483,N_22807);
and U24289 (N_24289,N_22939,N_23695);
and U24290 (N_24290,N_22311,N_22116);
and U24291 (N_24291,N_23292,N_23370);
xor U24292 (N_24292,N_22613,N_22884);
nor U24293 (N_24293,N_22320,N_23425);
xor U24294 (N_24294,N_22813,N_23520);
xor U24295 (N_24295,N_23668,N_23161);
and U24296 (N_24296,N_23321,N_22380);
nand U24297 (N_24297,N_22367,N_22987);
or U24298 (N_24298,N_22670,N_23159);
nor U24299 (N_24299,N_23827,N_23023);
nand U24300 (N_24300,N_22866,N_23410);
or U24301 (N_24301,N_22552,N_23163);
and U24302 (N_24302,N_23625,N_22675);
or U24303 (N_24303,N_23971,N_23497);
and U24304 (N_24304,N_22998,N_23539);
nand U24305 (N_24305,N_22460,N_22588);
or U24306 (N_24306,N_22435,N_22010);
and U24307 (N_24307,N_22329,N_23510);
nand U24308 (N_24308,N_22310,N_22699);
and U24309 (N_24309,N_22618,N_22647);
nor U24310 (N_24310,N_22210,N_22300);
or U24311 (N_24311,N_23631,N_22730);
or U24312 (N_24312,N_22218,N_23081);
or U24313 (N_24313,N_23731,N_22179);
nand U24314 (N_24314,N_22030,N_23957);
nand U24315 (N_24315,N_23655,N_23617);
nor U24316 (N_24316,N_23750,N_23608);
or U24317 (N_24317,N_23355,N_22579);
or U24318 (N_24318,N_22479,N_23475);
or U24319 (N_24319,N_22820,N_22397);
xor U24320 (N_24320,N_23945,N_22754);
nor U24321 (N_24321,N_22557,N_22042);
or U24322 (N_24322,N_23172,N_23966);
nor U24323 (N_24323,N_23459,N_23804);
and U24324 (N_24324,N_22313,N_23919);
and U24325 (N_24325,N_22636,N_23878);
nor U24326 (N_24326,N_23190,N_22819);
nor U24327 (N_24327,N_22835,N_23095);
nor U24328 (N_24328,N_22624,N_22689);
xor U24329 (N_24329,N_23815,N_22642);
nand U24330 (N_24330,N_23902,N_22921);
nor U24331 (N_24331,N_23892,N_23953);
or U24332 (N_24332,N_23114,N_23044);
nor U24333 (N_24333,N_22976,N_22454);
nand U24334 (N_24334,N_23844,N_22614);
and U24335 (N_24335,N_22569,N_22610);
nor U24336 (N_24336,N_22594,N_22031);
or U24337 (N_24337,N_23607,N_23099);
nand U24338 (N_24338,N_23087,N_23538);
and U24339 (N_24339,N_22145,N_22663);
nand U24340 (N_24340,N_23426,N_23174);
xor U24341 (N_24341,N_23286,N_22843);
and U24342 (N_24342,N_23071,N_23348);
or U24343 (N_24343,N_22457,N_22083);
nor U24344 (N_24344,N_23400,N_23504);
and U24345 (N_24345,N_22669,N_22132);
xor U24346 (N_24346,N_22039,N_22788);
nand U24347 (N_24347,N_23967,N_22949);
and U24348 (N_24348,N_23935,N_23941);
nand U24349 (N_24349,N_22387,N_23768);
or U24350 (N_24350,N_22181,N_22567);
and U24351 (N_24351,N_22153,N_22331);
nand U24352 (N_24352,N_23247,N_23798);
nand U24353 (N_24353,N_22162,N_22289);
xnor U24354 (N_24354,N_23671,N_23952);
xnor U24355 (N_24355,N_22109,N_23272);
or U24356 (N_24356,N_22902,N_22826);
nand U24357 (N_24357,N_23210,N_23021);
nor U24358 (N_24358,N_23378,N_22571);
or U24359 (N_24359,N_23049,N_22534);
and U24360 (N_24360,N_22694,N_22716);
and U24361 (N_24361,N_23328,N_23678);
and U24362 (N_24362,N_23532,N_23696);
nor U24363 (N_24363,N_22043,N_22194);
nor U24364 (N_24364,N_23340,N_22375);
xnor U24365 (N_24365,N_22793,N_23517);
xor U24366 (N_24366,N_23033,N_22124);
nor U24367 (N_24367,N_23780,N_23835);
and U24368 (N_24368,N_23143,N_23359);
nor U24369 (N_24369,N_22049,N_22531);
nand U24370 (N_24370,N_23437,N_22488);
nor U24371 (N_24371,N_23406,N_23871);
or U24372 (N_24372,N_22525,N_22513);
nand U24373 (N_24373,N_22688,N_23252);
nand U24374 (N_24374,N_22092,N_22745);
nor U24375 (N_24375,N_22978,N_23544);
and U24376 (N_24376,N_22544,N_23772);
nand U24377 (N_24377,N_23746,N_22520);
and U24378 (N_24378,N_23995,N_22325);
xnor U24379 (N_24379,N_23943,N_23144);
nand U24380 (N_24380,N_23623,N_23323);
nand U24381 (N_24381,N_22709,N_23924);
or U24382 (N_24382,N_23626,N_23884);
or U24383 (N_24383,N_22924,N_23546);
or U24384 (N_24384,N_22327,N_22617);
or U24385 (N_24385,N_22122,N_22216);
xnor U24386 (N_24386,N_22518,N_23663);
or U24387 (N_24387,N_23713,N_22040);
and U24388 (N_24388,N_23681,N_23752);
nand U24389 (N_24389,N_22810,N_22232);
nor U24390 (N_24390,N_23982,N_22522);
or U24391 (N_24391,N_22038,N_22197);
or U24392 (N_24392,N_22738,N_23599);
or U24393 (N_24393,N_22545,N_23781);
nand U24394 (N_24394,N_23877,N_23022);
or U24395 (N_24395,N_23611,N_22372);
nor U24396 (N_24396,N_23339,N_23531);
and U24397 (N_24397,N_22756,N_22860);
nor U24398 (N_24398,N_22041,N_22868);
xnor U24399 (N_24399,N_23921,N_22927);
nand U24400 (N_24400,N_22827,N_22390);
or U24401 (N_24401,N_23377,N_23035);
nand U24402 (N_24402,N_22929,N_23906);
nand U24403 (N_24403,N_23969,N_23079);
xor U24404 (N_24404,N_23553,N_23233);
or U24405 (N_24405,N_23183,N_22088);
or U24406 (N_24406,N_22601,N_23481);
nand U24407 (N_24407,N_23390,N_22200);
and U24408 (N_24408,N_23291,N_23466);
nand U24409 (N_24409,N_23718,N_23758);
or U24410 (N_24410,N_22980,N_22309);
nand U24411 (N_24411,N_22014,N_23993);
nand U24412 (N_24412,N_23518,N_22950);
or U24413 (N_24413,N_23075,N_22503);
nor U24414 (N_24414,N_22551,N_22931);
or U24415 (N_24415,N_23416,N_23998);
and U24416 (N_24416,N_22811,N_22008);
or U24417 (N_24417,N_22415,N_23238);
nand U24418 (N_24418,N_23637,N_23470);
or U24419 (N_24419,N_22303,N_23541);
and U24420 (N_24420,N_22237,N_23867);
and U24421 (N_24421,N_23013,N_23256);
or U24422 (N_24422,N_22121,N_23851);
xor U24423 (N_24423,N_22243,N_23929);
and U24424 (N_24424,N_23633,N_23398);
and U24425 (N_24425,N_23264,N_22606);
and U24426 (N_24426,N_23897,N_22672);
nor U24427 (N_24427,N_23177,N_22576);
or U24428 (N_24428,N_22155,N_22409);
nand U24429 (N_24429,N_23821,N_22848);
xor U24430 (N_24430,N_23357,N_23014);
nor U24431 (N_24431,N_22449,N_23677);
nand U24432 (N_24432,N_22198,N_22273);
xnor U24433 (N_24433,N_23882,N_23476);
xor U24434 (N_24434,N_23948,N_22432);
nor U24435 (N_24435,N_23012,N_23184);
and U24436 (N_24436,N_22058,N_22822);
nor U24437 (N_24437,N_22765,N_23834);
or U24438 (N_24438,N_23939,N_22984);
nand U24439 (N_24439,N_22744,N_23807);
nor U24440 (N_24440,N_23445,N_23119);
and U24441 (N_24441,N_23862,N_23600);
xnor U24442 (N_24442,N_23484,N_23932);
nor U24443 (N_24443,N_23147,N_22700);
xor U24444 (N_24444,N_22287,N_22484);
nand U24445 (N_24445,N_23017,N_23651);
and U24446 (N_24446,N_23001,N_22072);
or U24447 (N_24447,N_22134,N_22421);
nand U24448 (N_24448,N_22318,N_23365);
and U24449 (N_24449,N_23534,N_22334);
or U24450 (N_24450,N_23672,N_23648);
and U24451 (N_24451,N_22814,N_23204);
and U24452 (N_24452,N_22880,N_23254);
nand U24453 (N_24453,N_22212,N_22507);
xnor U24454 (N_24454,N_22533,N_22515);
xnor U24455 (N_24455,N_23961,N_22885);
nand U24456 (N_24456,N_23999,N_23786);
xnor U24457 (N_24457,N_23198,N_22280);
xnor U24458 (N_24458,N_23872,N_22413);
xnor U24459 (N_24459,N_22965,N_23444);
xnor U24460 (N_24460,N_23741,N_23667);
nand U24461 (N_24461,N_23234,N_22277);
xor U24462 (N_24462,N_23353,N_22595);
and U24463 (N_24463,N_23456,N_23635);
or U24464 (N_24464,N_22708,N_23330);
nand U24465 (N_24465,N_22365,N_22136);
nor U24466 (N_24466,N_22948,N_23138);
xnor U24467 (N_24467,N_22407,N_23216);
nand U24468 (N_24468,N_23529,N_23509);
or U24469 (N_24469,N_23894,N_23876);
nor U24470 (N_24470,N_22295,N_22801);
xor U24471 (N_24471,N_22314,N_23787);
xnor U24472 (N_24472,N_22637,N_23770);
xnor U24473 (N_24473,N_22064,N_23986);
nand U24474 (N_24474,N_22163,N_22773);
or U24475 (N_24475,N_23249,N_23329);
xnor U24476 (N_24476,N_23285,N_23226);
or U24477 (N_24477,N_22593,N_23979);
and U24478 (N_24478,N_22102,N_22497);
or U24479 (N_24479,N_23322,N_23751);
and U24480 (N_24480,N_22702,N_22402);
nor U24481 (N_24481,N_22078,N_23714);
or U24482 (N_24482,N_23927,N_22274);
or U24483 (N_24483,N_22398,N_23628);
xnor U24484 (N_24484,N_23737,N_22735);
and U24485 (N_24485,N_22489,N_23507);
nor U24486 (N_24486,N_22769,N_23104);
or U24487 (N_24487,N_23526,N_22973);
or U24488 (N_24488,N_22678,N_23222);
nor U24489 (N_24489,N_22141,N_23211);
xnor U24490 (N_24490,N_22661,N_22057);
nor U24491 (N_24491,N_23124,N_23869);
nand U24492 (N_24492,N_23176,N_23318);
xor U24493 (N_24493,N_23764,N_22073);
nand U24494 (N_24494,N_23293,N_23324);
nor U24495 (N_24495,N_22004,N_22292);
nand U24496 (N_24496,N_22911,N_22481);
xnor U24497 (N_24497,N_23068,N_23890);
nor U24498 (N_24498,N_22546,N_23789);
or U24499 (N_24499,N_23595,N_22874);
xor U24500 (N_24500,N_23288,N_23823);
nand U24501 (N_24501,N_22296,N_22586);
xor U24502 (N_24502,N_23478,N_22555);
or U24503 (N_24503,N_22644,N_22317);
or U24504 (N_24504,N_22346,N_23306);
xnor U24505 (N_24505,N_22021,N_23408);
and U24506 (N_24506,N_22264,N_23372);
or U24507 (N_24507,N_22003,N_22695);
and U24508 (N_24508,N_23158,N_22306);
nor U24509 (N_24509,N_23584,N_22736);
nand U24510 (N_24510,N_23059,N_22138);
nor U24511 (N_24511,N_22384,N_22562);
nor U24512 (N_24512,N_23225,N_23782);
and U24513 (N_24513,N_23424,N_22781);
and U24514 (N_24514,N_23722,N_23450);
and U24515 (N_24515,N_23432,N_23384);
nor U24516 (N_24516,N_22361,N_23785);
nand U24517 (N_24517,N_22467,N_23698);
nor U24518 (N_24518,N_22442,N_23351);
nor U24519 (N_24519,N_23728,N_23822);
xor U24520 (N_24520,N_22800,N_23208);
and U24521 (N_24521,N_23199,N_23463);
or U24522 (N_24522,N_22227,N_23644);
xor U24523 (N_24523,N_23609,N_23061);
xor U24524 (N_24524,N_22344,N_23251);
or U24525 (N_24525,N_23290,N_22271);
xor U24526 (N_24526,N_23653,N_22560);
nor U24527 (N_24527,N_23018,N_23602);
nor U24528 (N_24528,N_23349,N_23056);
xnor U24529 (N_24529,N_23673,N_22620);
nand U24530 (N_24530,N_22205,N_22247);
and U24531 (N_24531,N_22368,N_22374);
nor U24532 (N_24532,N_23765,N_23624);
nand U24533 (N_24533,N_23032,N_23934);
or U24534 (N_24534,N_22505,N_22177);
xor U24535 (N_24535,N_23812,N_22934);
or U24536 (N_24536,N_22217,N_22235);
or U24537 (N_24537,N_23462,N_22164);
nand U24538 (N_24538,N_23716,N_22603);
or U24539 (N_24539,N_22034,N_23230);
nor U24540 (N_24540,N_23579,N_23136);
xnor U24541 (N_24541,N_22480,N_23489);
nand U24542 (N_24542,N_22101,N_23447);
or U24543 (N_24543,N_22220,N_22501);
and U24544 (N_24544,N_22098,N_22015);
or U24545 (N_24545,N_23096,N_22097);
and U24546 (N_24546,N_22667,N_22281);
xnor U24547 (N_24547,N_22364,N_22910);
and U24548 (N_24548,N_22566,N_23051);
or U24549 (N_24549,N_23117,N_23297);
nand U24550 (N_24550,N_23820,N_23221);
or U24551 (N_24551,N_23343,N_22405);
or U24552 (N_24552,N_23739,N_22864);
nor U24553 (N_24553,N_22608,N_23567);
and U24554 (N_24554,N_23800,N_23846);
or U24555 (N_24555,N_23205,N_23959);
nor U24556 (N_24556,N_23311,N_23170);
xnor U24557 (N_24557,N_23395,N_22916);
or U24558 (N_24558,N_22521,N_22487);
nor U24559 (N_24559,N_22096,N_23819);
and U24560 (N_24560,N_22841,N_23810);
xnor U24561 (N_24561,N_22203,N_23473);
nor U24562 (N_24562,N_22653,N_22171);
and U24563 (N_24563,N_22535,N_23125);
nand U24564 (N_24564,N_23828,N_22723);
and U24565 (N_24565,N_23670,N_22741);
xnor U24566 (N_24566,N_22795,N_22117);
nor U24567 (N_24567,N_23674,N_22363);
nand U24568 (N_24568,N_23963,N_22896);
nand U24569 (N_24569,N_22024,N_22912);
or U24570 (N_24570,N_23706,N_23128);
or U24571 (N_24571,N_22234,N_22938);
nor U24572 (N_24572,N_22063,N_22692);
or U24573 (N_24573,N_22790,N_22347);
nand U24574 (N_24574,N_22815,N_23972);
and U24575 (N_24575,N_23775,N_22476);
and U24576 (N_24576,N_23236,N_23895);
nand U24577 (N_24577,N_22887,N_23137);
xor U24578 (N_24578,N_22995,N_22940);
and U24579 (N_24579,N_23000,N_23284);
and U24580 (N_24580,N_22283,N_23098);
nor U24581 (N_24581,N_22657,N_23643);
nand U24582 (N_24582,N_23058,N_23201);
xor U24583 (N_24583,N_22249,N_23332);
nor U24584 (N_24584,N_22664,N_22993);
and U24585 (N_24585,N_22590,N_22679);
and U24586 (N_24586,N_22582,N_23101);
or U24587 (N_24587,N_22783,N_23500);
nor U24588 (N_24588,N_22898,N_23729);
or U24589 (N_24589,N_22192,N_22340);
nor U24590 (N_24590,N_23734,N_23975);
nand U24591 (N_24591,N_23715,N_23464);
xnor U24592 (N_24592,N_22408,N_22540);
or U24593 (N_24593,N_22568,N_23552);
nor U24594 (N_24594,N_22350,N_23053);
and U24595 (N_24595,N_22966,N_22444);
nor U24596 (N_24596,N_23451,N_23983);
and U24597 (N_24597,N_23103,N_23175);
nor U24598 (N_24598,N_23797,N_22429);
and U24599 (N_24599,N_23085,N_22899);
or U24600 (N_24600,N_23002,N_23832);
xor U24601 (N_24601,N_23837,N_23115);
and U24602 (N_24602,N_22905,N_22208);
or U24603 (N_24603,N_22766,N_22532);
and U24604 (N_24604,N_23645,N_22207);
xnor U24605 (N_24605,N_23680,N_23278);
and U24606 (N_24606,N_23836,N_23350);
or U24607 (N_24607,N_22362,N_23853);
or U24608 (N_24608,N_23220,N_23064);
nand U24609 (N_24609,N_23366,N_22882);
nand U24610 (N_24610,N_22293,N_22165);
or U24611 (N_24611,N_23031,N_23614);
or U24612 (N_24612,N_22025,N_23336);
and U24613 (N_24613,N_22337,N_23215);
nor U24614 (N_24614,N_23683,N_22685);
nor U24615 (N_24615,N_23160,N_23916);
or U24616 (N_24616,N_23488,N_23537);
nand U24617 (N_24617,N_22585,N_22502);
or U24618 (N_24618,N_23361,N_22242);
nor U24619 (N_24619,N_22370,N_22671);
and U24620 (N_24620,N_22443,N_23362);
nor U24621 (N_24621,N_23503,N_23757);
nand U24622 (N_24622,N_22369,N_23988);
or U24623 (N_24623,N_23597,N_22893);
xnor U24624 (N_24624,N_23268,N_22782);
and U24625 (N_24625,N_23055,N_23566);
and U24626 (N_24626,N_22424,N_23636);
and U24627 (N_24627,N_22406,N_22537);
nand U24628 (N_24628,N_22417,N_23621);
xnor U24629 (N_24629,N_22903,N_23422);
nor U24630 (N_24630,N_22378,N_22865);
or U24631 (N_24631,N_23156,N_23502);
nand U24632 (N_24632,N_22389,N_22437);
and U24633 (N_24633,N_22646,N_23335);
nand U24634 (N_24634,N_23997,N_23333);
nand U24635 (N_24635,N_23868,N_22026);
nor U24636 (N_24636,N_23258,N_23551);
nor U24637 (N_24637,N_23802,N_23062);
nand U24638 (N_24638,N_23433,N_22750);
and U24639 (N_24639,N_23282,N_23839);
nor U24640 (N_24640,N_23438,N_23976);
xor U24641 (N_24641,N_22059,N_22184);
nor U24642 (N_24642,N_22423,N_23202);
and U24643 (N_24643,N_23097,N_23223);
nand U24644 (N_24644,N_23499,N_22319);
nor U24645 (N_24645,N_23038,N_23460);
xnor U24646 (N_24646,N_22099,N_22839);
xnor U24647 (N_24647,N_22191,N_23393);
and U24648 (N_24648,N_23669,N_23076);
xnor U24649 (N_24649,N_23418,N_22530);
xor U24650 (N_24650,N_22852,N_23283);
xor U24651 (N_24651,N_23387,N_23554);
xnor U24652 (N_24652,N_22482,N_23931);
xnor U24653 (N_24653,N_22662,N_22336);
nand U24654 (N_24654,N_23030,N_22258);
or U24655 (N_24655,N_23557,N_22167);
xor U24656 (N_24656,N_22431,N_23334);
xnor U24657 (N_24657,N_22343,N_22784);
nor U24658 (N_24658,N_22199,N_22214);
nor U24659 (N_24659,N_22209,N_23917);
nand U24660 (N_24660,N_23040,N_22875);
and U24661 (N_24661,N_22666,N_22913);
or U24662 (N_24662,N_22722,N_23968);
and U24663 (N_24663,N_22683,N_22068);
nand U24664 (N_24664,N_23687,N_23083);
and U24665 (N_24665,N_22471,N_23791);
or U24666 (N_24666,N_22676,N_22426);
nand U24667 (N_24667,N_22746,N_23926);
xor U24668 (N_24668,N_23795,N_22005);
and U24669 (N_24669,N_23164,N_22404);
and U24670 (N_24670,N_23259,N_22245);
and U24671 (N_24671,N_22433,N_22383);
nor U24672 (N_24672,N_23442,N_23883);
nand U24673 (N_24673,N_22395,N_23342);
xnor U24674 (N_24674,N_23574,N_23496);
or U24675 (N_24675,N_22818,N_23721);
nand U24676 (N_24676,N_23427,N_22574);
nand U24677 (N_24677,N_23980,N_23050);
and U24678 (N_24678,N_23080,N_22358);
xor U24679 (N_24679,N_23630,N_22659);
nor U24680 (N_24680,N_23298,N_23319);
and U24681 (N_24681,N_22183,N_22178);
nand U24682 (N_24682,N_22143,N_22504);
or U24683 (N_24683,N_23613,N_22832);
xor U24684 (N_24684,N_22936,N_23987);
and U24685 (N_24685,N_22233,N_22051);
nor U24686 (N_24686,N_23569,N_23093);
or U24687 (N_24687,N_22705,N_22272);
nand U24688 (N_24688,N_23833,N_22834);
nand U24689 (N_24689,N_23182,N_22017);
nor U24690 (N_24690,N_22439,N_23130);
xnor U24691 (N_24691,N_23046,N_23261);
or U24692 (N_24692,N_23632,N_23989);
and U24693 (N_24693,N_23316,N_23958);
or U24694 (N_24694,N_23274,N_22269);
and U24695 (N_24695,N_22840,N_23514);
and U24696 (N_24696,N_22596,N_23189);
or U24697 (N_24697,N_23341,N_22118);
xnor U24698 (N_24698,N_23726,N_23570);
xor U24699 (N_24699,N_22027,N_23380);
nand U24700 (N_24700,N_22992,N_23294);
or U24701 (N_24701,N_23300,N_23736);
or U24702 (N_24702,N_22022,N_22514);
xnor U24703 (N_24703,N_22656,N_22400);
nand U24704 (N_24704,N_23686,N_22251);
or U24705 (N_24705,N_22862,N_22821);
and U24706 (N_24706,N_23168,N_23691);
xor U24707 (N_24707,N_22706,N_22182);
and U24708 (N_24708,N_22495,N_22952);
and U24709 (N_24709,N_22556,N_22789);
and U24710 (N_24710,N_23458,N_23994);
nand U24711 (N_24711,N_22011,N_23417);
or U24712 (N_24712,N_23845,N_22681);
xnor U24713 (N_24713,N_23166,N_22150);
nor U24714 (N_24714,N_23985,N_22156);
or U24715 (N_24715,N_23792,N_23078);
or U24716 (N_24716,N_23448,N_23402);
and U24717 (N_24717,N_23522,N_22904);
nand U24718 (N_24718,N_22844,N_23692);
or U24719 (N_24719,N_22846,N_22890);
and U24720 (N_24720,N_22037,N_23915);
or U24721 (N_24721,N_23779,N_23271);
xnor U24722 (N_24722,N_23315,N_22013);
xnor U24723 (N_24723,N_22201,N_22691);
nor U24724 (N_24724,N_23430,N_22906);
and U24725 (N_24725,N_22833,N_23067);
nor U24726 (N_24726,N_23276,N_22204);
nand U24727 (N_24727,N_22895,N_22106);
nand U24728 (N_24728,N_23253,N_22075);
nor U24729 (N_24729,N_22441,N_23705);
nor U24730 (N_24730,N_23063,N_23725);
and U24731 (N_24731,N_22268,N_22731);
nand U24732 (N_24732,N_23027,N_22809);
nor U24733 (N_24733,N_23831,N_22564);
and U24734 (N_24734,N_23265,N_22589);
or U24735 (N_24735,N_23808,N_22359);
nor U24736 (N_24736,N_22202,N_22461);
or U24737 (N_24737,N_23443,N_23374);
and U24738 (N_24738,N_22291,N_22933);
xor U24739 (N_24739,N_22506,N_22416);
and U24740 (N_24740,N_22930,N_22305);
xor U24741 (N_24741,N_23524,N_23710);
and U24742 (N_24742,N_22990,N_23310);
or U24743 (N_24743,N_23842,N_23825);
nand U24744 (N_24744,N_22225,N_23206);
nor U24745 (N_24745,N_22778,N_22348);
nor U24746 (N_24746,N_22805,N_23449);
nor U24747 (N_24747,N_22584,N_23964);
xnor U24748 (N_24748,N_23113,N_22541);
nor U24749 (N_24749,N_22478,N_22668);
and U24750 (N_24750,N_22697,N_23829);
and U24751 (N_24751,N_23910,N_22465);
and U24752 (N_24752,N_23605,N_22892);
or U24753 (N_24753,N_23382,N_22069);
and U24754 (N_24754,N_23944,N_22260);
and U24755 (N_24755,N_22002,N_23352);
nand U24756 (N_24756,N_22094,N_23996);
nor U24757 (N_24757,N_22863,N_22956);
or U24758 (N_24758,N_22382,N_22677);
and U24759 (N_24759,N_22152,N_22777);
and U24760 (N_24760,N_22091,N_23783);
or U24761 (N_24761,N_22631,N_22599);
and U24762 (N_24762,N_23389,N_22297);
or U24763 (N_24763,N_23468,N_22600);
xor U24764 (N_24764,N_23841,N_23105);
xor U24765 (N_24765,N_22381,N_22312);
nor U24766 (N_24766,N_23054,N_22278);
and U24767 (N_24767,N_22989,N_22148);
or U24768 (N_24768,N_23913,N_23991);
or U24769 (N_24769,N_23900,N_22090);
and U24770 (N_24770,N_22047,N_23041);
xnor U24771 (N_24771,N_23346,N_23218);
nand U24772 (N_24772,N_22290,N_22029);
xnor U24773 (N_24773,N_23685,N_23106);
or U24774 (N_24774,N_22649,N_23180);
xnor U24775 (N_24775,N_23816,N_22763);
nor U24776 (N_24776,N_23946,N_22825);
nor U24777 (N_24777,N_23962,N_22881);
nor U24778 (N_24778,N_23228,N_22684);
or U24779 (N_24779,N_23824,N_22373);
and U24780 (N_24780,N_22139,N_23091);
or U24781 (N_24781,N_23693,N_22036);
or U24782 (N_24782,N_23391,N_23970);
nor U24783 (N_24783,N_23440,N_23077);
and U24784 (N_24784,N_22447,N_22817);
xnor U24785 (N_24785,N_22701,N_22578);
nand U24786 (N_24786,N_23429,N_23193);
nor U24787 (N_24787,N_22170,N_23708);
xnor U24788 (N_24788,N_23738,N_23305);
or U24789 (N_24789,N_22776,N_22673);
nand U24790 (N_24790,N_23847,N_22105);
or U24791 (N_24791,N_22951,N_23586);
or U24792 (N_24792,N_22226,N_22857);
nor U24793 (N_24793,N_22962,N_23766);
and U24794 (N_24794,N_22018,N_23194);
or U24795 (N_24795,N_22549,N_23796);
nand U24796 (N_24796,N_22622,N_22830);
nor U24797 (N_24797,N_23102,N_22526);
or U24798 (N_24798,N_22130,N_22937);
nor U24799 (N_24799,N_23498,N_22428);
nand U24800 (N_24800,N_23735,N_23762);
nand U24801 (N_24801,N_23591,N_23852);
or U24802 (N_24802,N_22213,N_22996);
nor U24803 (N_24803,N_22734,N_23654);
nand U24804 (N_24804,N_23407,N_23646);
xnor U24805 (N_24805,N_22276,N_22379);
nand U24806 (N_24806,N_23109,N_23908);
or U24807 (N_24807,N_22009,N_23037);
nor U24808 (N_24808,N_23207,N_23405);
xor U24809 (N_24809,N_23583,N_23326);
xnor U24810 (N_24810,N_23587,N_23145);
and U24811 (N_24811,N_22254,N_22803);
nand U24812 (N_24812,N_22686,N_22129);
nor U24813 (N_24813,N_22420,N_23793);
nor U24814 (N_24814,N_23381,N_23327);
xnor U24815 (N_24815,N_22941,N_23200);
xor U24816 (N_24816,N_23575,N_23026);
or U24817 (N_24817,N_23116,N_22412);
nor U24818 (N_24818,N_22760,N_22935);
nand U24819 (N_24819,N_23325,N_22256);
nand U24820 (N_24820,N_23454,N_22238);
nand U24821 (N_24821,N_22196,N_22304);
and U24822 (N_24822,N_23523,N_22828);
xor U24823 (N_24823,N_23360,N_23592);
nor U24824 (N_24824,N_22718,N_22986);
xor U24825 (N_24825,N_23640,N_23777);
nor U24826 (N_24826,N_22386,N_23688);
and U24827 (N_24827,N_23005,N_22748);
or U24828 (N_24828,N_23550,N_22263);
xnor U24829 (N_24829,N_22324,N_22103);
nand U24830 (N_24830,N_22974,N_23530);
or U24831 (N_24831,N_22804,N_23711);
or U24832 (N_24832,N_22836,N_22419);
xnor U24833 (N_24833,N_23131,N_22187);
and U24834 (N_24834,N_23072,N_22223);
or U24835 (N_24835,N_23679,N_23848);
and U24836 (N_24836,N_22224,N_23446);
nor U24837 (N_24837,N_22257,N_23760);
xnor U24838 (N_24838,N_23371,N_23992);
nor U24839 (N_24839,N_22598,N_23120);
nor U24840 (N_24840,N_22288,N_22385);
nor U24841 (N_24841,N_23248,N_23126);
nand U24842 (N_24842,N_22855,N_23879);
or U24843 (N_24843,N_23185,N_22104);
or U24844 (N_24844,N_23571,N_22055);
nor U24845 (N_24845,N_22550,N_22524);
nand U24846 (N_24846,N_22983,N_22891);
nor U24847 (N_24847,N_23165,N_22696);
nand U24848 (N_24848,N_22089,N_23392);
nand U24849 (N_24849,N_22498,N_22861);
nor U24850 (N_24850,N_22108,N_22774);
or U24851 (N_24851,N_23088,N_23704);
and U24852 (N_24852,N_23299,N_22275);
xor U24853 (N_24853,N_22963,N_22605);
xor U24854 (N_24854,N_23487,N_23240);
nand U24855 (N_24855,N_23453,N_22282);
or U24856 (N_24856,N_22512,N_23925);
or U24857 (N_24857,N_22252,N_22528);
or U24858 (N_24858,N_22770,N_23060);
nor U24859 (N_24859,N_22630,N_22894);
xor U24860 (N_24860,N_22823,N_23219);
and U24861 (N_24861,N_23016,N_22453);
nor U24862 (N_24862,N_23263,N_23818);
nor U24863 (N_24863,N_22377,N_22627);
nor U24864 (N_24864,N_23004,N_22239);
nor U24865 (N_24865,N_22466,N_22157);
nand U24866 (N_24866,N_22074,N_23364);
and U24867 (N_24867,N_23860,N_22573);
and U24868 (N_24868,N_22674,N_23212);
or U24869 (N_24869,N_22113,N_23479);
or U24870 (N_24870,N_23167,N_22961);
xnor U24871 (N_24871,N_23231,N_22739);
xnor U24872 (N_24872,N_22740,N_22459);
nor U24873 (N_24873,N_22430,N_22335);
nand U24874 (N_24874,N_23270,N_23279);
or U24875 (N_24875,N_22529,N_22615);
nand U24876 (N_24876,N_22797,N_23659);
nand U24877 (N_24877,N_22638,N_23799);
nand U24878 (N_24878,N_23622,N_22640);
xnor U24879 (N_24879,N_22028,N_22496);
nand U24880 (N_24880,N_23598,N_23173);
xor U24881 (N_24881,N_23065,N_23412);
xnor U24882 (N_24882,N_23914,N_22248);
nand U24883 (N_24883,N_22286,N_22345);
nand U24884 (N_24884,N_23140,N_23434);
nor U24885 (N_24885,N_23465,N_23562);
nand U24886 (N_24886,N_22907,N_22366);
or U24887 (N_24887,N_23419,N_22967);
and U24888 (N_24888,N_22982,N_22266);
nor U24889 (N_24889,N_22712,N_23594);
nor U24890 (N_24890,N_23904,N_23415);
or U24891 (N_24891,N_23094,N_23767);
nand U24892 (N_24892,N_23515,N_23639);
nand U24893 (N_24893,N_22032,N_22771);
or U24894 (N_24894,N_22222,N_22509);
or U24895 (N_24895,N_23148,N_23227);
nand U24896 (N_24896,N_22330,N_22253);
xnor U24897 (N_24897,N_23073,N_22180);
nor U24898 (N_24898,N_22112,N_22972);
and U24899 (N_24899,N_22629,N_22019);
nand U24900 (N_24900,N_23015,N_23474);
xnor U24901 (N_24901,N_23581,N_23732);
or U24902 (N_24902,N_23701,N_23313);
nor U24903 (N_24903,N_23582,N_22621);
or U24904 (N_24904,N_22000,N_22326);
nor U24905 (N_24905,N_23866,N_23974);
or U24906 (N_24906,N_23697,N_23954);
nand U24907 (N_24907,N_23978,N_22539);
xnor U24908 (N_24908,N_22006,N_23266);
and U24909 (N_24909,N_22877,N_23169);
or U24910 (N_24910,N_23849,N_23092);
nand U24911 (N_24911,N_23580,N_22076);
nand U24912 (N_24912,N_22452,N_22050);
or U24913 (N_24913,N_22114,N_23461);
nand U24914 (N_24914,N_23755,N_23857);
or U24915 (N_24915,N_23084,N_23638);
and U24916 (N_24916,N_22081,N_22451);
and U24917 (N_24917,N_23709,N_22994);
or U24918 (N_24918,N_23171,N_22791);
nand U24919 (N_24919,N_22915,N_23956);
and U24920 (N_24920,N_23527,N_23556);
or U24921 (N_24921,N_23856,N_22997);
xor U24922 (N_24922,N_23940,N_23025);
and U24923 (N_24923,N_23912,N_22796);
and U24924 (N_24924,N_22981,N_23858);
nor U24925 (N_24925,N_22988,N_23769);
nor U24926 (N_24926,N_23428,N_23658);
and U24927 (N_24927,N_22403,N_22154);
and U24928 (N_24928,N_22244,N_23733);
nor U24929 (N_24929,N_22785,N_23356);
nand U24930 (N_24930,N_23179,N_23070);
and U24931 (N_24931,N_22577,N_22206);
xnor U24932 (N_24932,N_23345,N_22942);
nor U24933 (N_24933,N_23891,N_22959);
nor U24934 (N_24934,N_22639,N_22710);
or U24935 (N_24935,N_23572,N_22626);
xor U24936 (N_24936,N_23907,N_22349);
and U24937 (N_24937,N_23887,N_22085);
or U24938 (N_24938,N_23747,N_22341);
nor U24939 (N_24939,N_23618,N_23008);
and U24940 (N_24940,N_23543,N_23107);
nand U24941 (N_24941,N_23505,N_23513);
or U24942 (N_24942,N_23162,N_23788);
xor U24943 (N_24943,N_23616,N_23814);
and U24944 (N_24944,N_22847,N_23188);
nor U24945 (N_24945,N_23308,N_22645);
xor U24946 (N_24946,N_23057,N_23794);
nor U24947 (N_24947,N_22858,N_22080);
and U24948 (N_24948,N_22690,N_22241);
or U24949 (N_24949,N_22808,N_23195);
and U24950 (N_24950,N_23275,N_23280);
nor U24951 (N_24951,N_22016,N_22737);
nor U24952 (N_24952,N_23139,N_22338);
or U24953 (N_24953,N_23863,N_22658);
nand U24954 (N_24954,N_23354,N_22294);
or U24955 (N_24955,N_23761,N_23578);
and U24956 (N_24956,N_23287,N_23903);
nor U24957 (N_24957,N_22779,N_22160);
or U24958 (N_24958,N_23528,N_22339);
nand U24959 (N_24959,N_22267,N_23650);
nor U24960 (N_24960,N_22628,N_23508);
nor U24961 (N_24961,N_23666,N_23129);
or U24962 (N_24962,N_22650,N_23045);
nand U24963 (N_24963,N_22084,N_22947);
and U24964 (N_24964,N_22977,N_22944);
xor U24965 (N_24965,N_22979,N_23899);
or U24966 (N_24966,N_23133,N_23217);
xor U24967 (N_24967,N_23368,N_22082);
or U24968 (N_24968,N_23850,N_22445);
nor U24969 (N_24969,N_22969,N_23886);
or U24970 (N_24970,N_23641,N_23257);
and U24971 (N_24971,N_23675,N_22123);
nor U24972 (N_24972,N_23187,N_23149);
or U24973 (N_24973,N_22219,N_22856);
or U24974 (N_24974,N_22410,N_22732);
and U24975 (N_24975,N_22355,N_22652);
xnor U24976 (N_24976,N_23560,N_23665);
nand U24977 (N_24977,N_22780,N_22173);
or U24978 (N_24978,N_22651,N_22655);
nor U24979 (N_24979,N_22743,N_23930);
and U24980 (N_24980,N_23656,N_22917);
nand U24981 (N_24981,N_22957,N_23682);
xnor U24982 (N_24982,N_23830,N_23506);
nor U24983 (N_24983,N_22632,N_22159);
and U24984 (N_24984,N_22761,N_22067);
xnor U24985 (N_24985,N_23521,N_22353);
or U24986 (N_24986,N_23019,N_22236);
nand U24987 (N_24987,N_23397,N_23548);
xnor U24988 (N_24988,N_22812,N_23949);
or U24989 (N_24989,N_23564,N_23034);
nor U24990 (N_24990,N_22755,N_22328);
xnor U24991 (N_24991,N_23565,N_23950);
nor U24992 (N_24992,N_22188,N_22321);
nand U24993 (N_24993,N_22035,N_22261);
nor U24994 (N_24994,N_23593,N_23805);
nand U24995 (N_24995,N_22592,N_23918);
xor U24996 (N_24996,N_22753,N_23660);
nand U24997 (N_24997,N_22491,N_23494);
xnor U24998 (N_24998,N_22127,N_22440);
and U24999 (N_24999,N_22878,N_23401);
nor U25000 (N_25000,N_23046,N_22313);
nand U25001 (N_25001,N_23756,N_22046);
xor U25002 (N_25002,N_23984,N_23980);
and U25003 (N_25003,N_22883,N_23752);
or U25004 (N_25004,N_23011,N_22976);
and U25005 (N_25005,N_23291,N_22360);
xor U25006 (N_25006,N_23372,N_22759);
or U25007 (N_25007,N_22188,N_22624);
nor U25008 (N_25008,N_23961,N_22929);
or U25009 (N_25009,N_22469,N_23963);
xnor U25010 (N_25010,N_23492,N_22365);
nand U25011 (N_25011,N_22202,N_22000);
or U25012 (N_25012,N_22370,N_23124);
nand U25013 (N_25013,N_23003,N_23774);
and U25014 (N_25014,N_23912,N_23925);
and U25015 (N_25015,N_22417,N_23656);
nor U25016 (N_25016,N_23868,N_23491);
nor U25017 (N_25017,N_22419,N_22847);
or U25018 (N_25018,N_22337,N_22918);
nor U25019 (N_25019,N_23392,N_23184);
xor U25020 (N_25020,N_22678,N_23653);
xor U25021 (N_25021,N_22547,N_23242);
nor U25022 (N_25022,N_23151,N_22149);
nor U25023 (N_25023,N_23100,N_23101);
nor U25024 (N_25024,N_22865,N_23034);
nor U25025 (N_25025,N_23009,N_22292);
and U25026 (N_25026,N_22007,N_22369);
xor U25027 (N_25027,N_23461,N_23655);
and U25028 (N_25028,N_22602,N_22273);
nor U25029 (N_25029,N_23978,N_23995);
or U25030 (N_25030,N_23165,N_22346);
nor U25031 (N_25031,N_23377,N_23728);
nand U25032 (N_25032,N_23932,N_22752);
nor U25033 (N_25033,N_22246,N_23019);
xor U25034 (N_25034,N_22628,N_23548);
xor U25035 (N_25035,N_23709,N_22490);
xnor U25036 (N_25036,N_23361,N_22318);
nand U25037 (N_25037,N_22967,N_22837);
nand U25038 (N_25038,N_23451,N_22009);
and U25039 (N_25039,N_22975,N_23799);
nand U25040 (N_25040,N_23871,N_22888);
or U25041 (N_25041,N_22125,N_22788);
nand U25042 (N_25042,N_22340,N_22402);
nand U25043 (N_25043,N_22519,N_22273);
xor U25044 (N_25044,N_23865,N_22486);
nor U25045 (N_25045,N_22989,N_22570);
or U25046 (N_25046,N_23491,N_22079);
xnor U25047 (N_25047,N_22938,N_22737);
nor U25048 (N_25048,N_23983,N_22229);
or U25049 (N_25049,N_23015,N_23268);
or U25050 (N_25050,N_22600,N_23426);
and U25051 (N_25051,N_22988,N_22014);
nand U25052 (N_25052,N_23629,N_22931);
and U25053 (N_25053,N_23219,N_22010);
nor U25054 (N_25054,N_23157,N_22310);
or U25055 (N_25055,N_22111,N_23243);
xnor U25056 (N_25056,N_22668,N_22881);
nand U25057 (N_25057,N_22454,N_23557);
nand U25058 (N_25058,N_23214,N_23313);
xnor U25059 (N_25059,N_22902,N_23439);
or U25060 (N_25060,N_23617,N_22581);
nor U25061 (N_25061,N_22954,N_22623);
nor U25062 (N_25062,N_23453,N_22149);
and U25063 (N_25063,N_22042,N_22380);
nand U25064 (N_25064,N_23127,N_22538);
and U25065 (N_25065,N_23907,N_22400);
and U25066 (N_25066,N_23211,N_22816);
nor U25067 (N_25067,N_23213,N_23357);
nand U25068 (N_25068,N_22667,N_22622);
and U25069 (N_25069,N_22493,N_22572);
or U25070 (N_25070,N_23622,N_23912);
or U25071 (N_25071,N_23239,N_22906);
nand U25072 (N_25072,N_22020,N_22730);
and U25073 (N_25073,N_23315,N_22419);
xor U25074 (N_25074,N_23238,N_23650);
and U25075 (N_25075,N_22075,N_22628);
nor U25076 (N_25076,N_22910,N_22674);
xor U25077 (N_25077,N_23857,N_23964);
nand U25078 (N_25078,N_22019,N_22230);
nor U25079 (N_25079,N_23800,N_23668);
or U25080 (N_25080,N_23284,N_22320);
or U25081 (N_25081,N_23890,N_23978);
or U25082 (N_25082,N_22490,N_22623);
nand U25083 (N_25083,N_22034,N_22894);
xnor U25084 (N_25084,N_22436,N_23821);
nor U25085 (N_25085,N_23492,N_22230);
or U25086 (N_25086,N_22404,N_23426);
or U25087 (N_25087,N_23677,N_22117);
nor U25088 (N_25088,N_23750,N_22634);
xnor U25089 (N_25089,N_23666,N_23150);
nor U25090 (N_25090,N_22885,N_22256);
or U25091 (N_25091,N_22174,N_22430);
and U25092 (N_25092,N_23372,N_23037);
nand U25093 (N_25093,N_23932,N_22983);
xor U25094 (N_25094,N_23036,N_23117);
and U25095 (N_25095,N_23428,N_23954);
xor U25096 (N_25096,N_22902,N_23620);
nor U25097 (N_25097,N_23359,N_22097);
xor U25098 (N_25098,N_23820,N_22121);
nand U25099 (N_25099,N_22629,N_23241);
and U25100 (N_25100,N_23924,N_23155);
xnor U25101 (N_25101,N_22937,N_23959);
and U25102 (N_25102,N_23687,N_22321);
xnor U25103 (N_25103,N_22401,N_22112);
or U25104 (N_25104,N_22608,N_23601);
nand U25105 (N_25105,N_22249,N_23111);
and U25106 (N_25106,N_23172,N_22237);
and U25107 (N_25107,N_23012,N_23742);
nor U25108 (N_25108,N_23706,N_22798);
and U25109 (N_25109,N_22528,N_22842);
nor U25110 (N_25110,N_22597,N_23856);
and U25111 (N_25111,N_22877,N_22450);
or U25112 (N_25112,N_22541,N_22051);
nor U25113 (N_25113,N_23829,N_22248);
or U25114 (N_25114,N_23196,N_23918);
nor U25115 (N_25115,N_23787,N_22510);
or U25116 (N_25116,N_23796,N_22862);
nand U25117 (N_25117,N_23971,N_22924);
or U25118 (N_25118,N_22626,N_22415);
nor U25119 (N_25119,N_23096,N_23974);
and U25120 (N_25120,N_23311,N_23933);
or U25121 (N_25121,N_22148,N_22753);
nand U25122 (N_25122,N_23629,N_22881);
xnor U25123 (N_25123,N_23631,N_23491);
or U25124 (N_25124,N_23938,N_22384);
nand U25125 (N_25125,N_22849,N_23720);
and U25126 (N_25126,N_22934,N_23077);
nand U25127 (N_25127,N_22133,N_22993);
or U25128 (N_25128,N_22104,N_23340);
nand U25129 (N_25129,N_23128,N_23877);
nand U25130 (N_25130,N_23491,N_23804);
and U25131 (N_25131,N_22349,N_22443);
xnor U25132 (N_25132,N_22653,N_22124);
nand U25133 (N_25133,N_23487,N_23670);
xnor U25134 (N_25134,N_23381,N_23920);
xnor U25135 (N_25135,N_22814,N_22605);
or U25136 (N_25136,N_22042,N_23162);
or U25137 (N_25137,N_22526,N_23497);
and U25138 (N_25138,N_22042,N_22425);
xnor U25139 (N_25139,N_22095,N_22192);
nand U25140 (N_25140,N_23785,N_22179);
xnor U25141 (N_25141,N_23490,N_22345);
or U25142 (N_25142,N_23335,N_23790);
xor U25143 (N_25143,N_22037,N_22076);
or U25144 (N_25144,N_22670,N_22232);
nand U25145 (N_25145,N_22233,N_22555);
or U25146 (N_25146,N_23720,N_22865);
and U25147 (N_25147,N_23193,N_22518);
nand U25148 (N_25148,N_23583,N_22794);
xor U25149 (N_25149,N_23835,N_22229);
nor U25150 (N_25150,N_22329,N_23215);
nand U25151 (N_25151,N_22693,N_22682);
and U25152 (N_25152,N_23231,N_22628);
nor U25153 (N_25153,N_23101,N_22215);
or U25154 (N_25154,N_23683,N_22753);
nor U25155 (N_25155,N_22602,N_23168);
nand U25156 (N_25156,N_23678,N_23839);
and U25157 (N_25157,N_23708,N_22212);
and U25158 (N_25158,N_23398,N_23247);
or U25159 (N_25159,N_23878,N_22626);
and U25160 (N_25160,N_22259,N_23829);
nand U25161 (N_25161,N_23817,N_22854);
and U25162 (N_25162,N_22053,N_22503);
or U25163 (N_25163,N_22577,N_23406);
nand U25164 (N_25164,N_23385,N_23448);
xor U25165 (N_25165,N_22815,N_23939);
and U25166 (N_25166,N_22532,N_23728);
nand U25167 (N_25167,N_22558,N_23211);
nor U25168 (N_25168,N_22486,N_22445);
or U25169 (N_25169,N_23922,N_22922);
and U25170 (N_25170,N_22875,N_22342);
xnor U25171 (N_25171,N_22819,N_22305);
or U25172 (N_25172,N_22981,N_22446);
xnor U25173 (N_25173,N_23789,N_22141);
nor U25174 (N_25174,N_23690,N_23657);
and U25175 (N_25175,N_22703,N_22114);
nand U25176 (N_25176,N_22422,N_22945);
nand U25177 (N_25177,N_23625,N_23460);
or U25178 (N_25178,N_23649,N_23181);
nor U25179 (N_25179,N_23311,N_23918);
or U25180 (N_25180,N_23206,N_22794);
or U25181 (N_25181,N_22627,N_22942);
or U25182 (N_25182,N_23353,N_22110);
nand U25183 (N_25183,N_23735,N_23964);
or U25184 (N_25184,N_22362,N_22653);
or U25185 (N_25185,N_22979,N_22691);
or U25186 (N_25186,N_23794,N_23294);
and U25187 (N_25187,N_22640,N_22176);
and U25188 (N_25188,N_22703,N_22162);
nor U25189 (N_25189,N_22588,N_23076);
nand U25190 (N_25190,N_23054,N_23729);
xnor U25191 (N_25191,N_23835,N_23542);
xnor U25192 (N_25192,N_23767,N_22091);
or U25193 (N_25193,N_22285,N_23251);
nor U25194 (N_25194,N_22529,N_22845);
nor U25195 (N_25195,N_22520,N_22934);
xor U25196 (N_25196,N_23557,N_22039);
nor U25197 (N_25197,N_22110,N_23340);
nor U25198 (N_25198,N_22976,N_23859);
or U25199 (N_25199,N_23376,N_22157);
or U25200 (N_25200,N_22200,N_22342);
nand U25201 (N_25201,N_22363,N_23808);
or U25202 (N_25202,N_22771,N_22670);
or U25203 (N_25203,N_23875,N_23560);
nand U25204 (N_25204,N_22162,N_22566);
nor U25205 (N_25205,N_23670,N_23173);
nor U25206 (N_25206,N_23006,N_22501);
xor U25207 (N_25207,N_23040,N_22564);
xor U25208 (N_25208,N_23275,N_22185);
nand U25209 (N_25209,N_22700,N_23559);
and U25210 (N_25210,N_23125,N_22178);
nor U25211 (N_25211,N_23351,N_22774);
nand U25212 (N_25212,N_22076,N_22252);
or U25213 (N_25213,N_22049,N_22200);
or U25214 (N_25214,N_22402,N_22894);
or U25215 (N_25215,N_23875,N_22801);
nand U25216 (N_25216,N_23226,N_23014);
xor U25217 (N_25217,N_22685,N_22286);
or U25218 (N_25218,N_22341,N_22256);
nor U25219 (N_25219,N_22738,N_22503);
and U25220 (N_25220,N_22687,N_23252);
nand U25221 (N_25221,N_22112,N_22172);
and U25222 (N_25222,N_23808,N_23475);
nor U25223 (N_25223,N_23247,N_23087);
or U25224 (N_25224,N_23016,N_23462);
xor U25225 (N_25225,N_23177,N_23501);
and U25226 (N_25226,N_23742,N_23668);
nor U25227 (N_25227,N_23363,N_23113);
or U25228 (N_25228,N_23747,N_23706);
and U25229 (N_25229,N_22212,N_22279);
and U25230 (N_25230,N_22019,N_23076);
nor U25231 (N_25231,N_22956,N_23362);
nand U25232 (N_25232,N_22239,N_23121);
nor U25233 (N_25233,N_23706,N_23911);
and U25234 (N_25234,N_22685,N_22499);
nand U25235 (N_25235,N_23006,N_23055);
or U25236 (N_25236,N_23582,N_22584);
or U25237 (N_25237,N_23682,N_22026);
nand U25238 (N_25238,N_22013,N_22370);
nor U25239 (N_25239,N_22390,N_22540);
nand U25240 (N_25240,N_22793,N_23546);
nand U25241 (N_25241,N_23485,N_22225);
and U25242 (N_25242,N_23139,N_23311);
or U25243 (N_25243,N_23015,N_23211);
or U25244 (N_25244,N_22192,N_23405);
and U25245 (N_25245,N_22982,N_22190);
or U25246 (N_25246,N_23545,N_23345);
or U25247 (N_25247,N_23024,N_22455);
and U25248 (N_25248,N_23478,N_23968);
xnor U25249 (N_25249,N_22299,N_23650);
nand U25250 (N_25250,N_23914,N_23491);
xor U25251 (N_25251,N_23302,N_22297);
and U25252 (N_25252,N_23689,N_23902);
nand U25253 (N_25253,N_22879,N_23429);
and U25254 (N_25254,N_23356,N_23671);
nor U25255 (N_25255,N_22298,N_23129);
nor U25256 (N_25256,N_22690,N_22940);
nand U25257 (N_25257,N_23395,N_23553);
nor U25258 (N_25258,N_22597,N_22121);
or U25259 (N_25259,N_22870,N_23645);
xnor U25260 (N_25260,N_22569,N_23987);
nand U25261 (N_25261,N_22651,N_23961);
nand U25262 (N_25262,N_22878,N_22332);
nor U25263 (N_25263,N_22866,N_23709);
and U25264 (N_25264,N_22703,N_22902);
or U25265 (N_25265,N_23477,N_23534);
xor U25266 (N_25266,N_23328,N_22199);
or U25267 (N_25267,N_22854,N_22596);
nand U25268 (N_25268,N_23359,N_22252);
and U25269 (N_25269,N_22746,N_23485);
or U25270 (N_25270,N_22320,N_22176);
nor U25271 (N_25271,N_23574,N_23456);
xnor U25272 (N_25272,N_23936,N_23162);
or U25273 (N_25273,N_22049,N_22294);
nand U25274 (N_25274,N_22168,N_22057);
and U25275 (N_25275,N_23041,N_22173);
or U25276 (N_25276,N_23310,N_23445);
xnor U25277 (N_25277,N_23662,N_22788);
nor U25278 (N_25278,N_23540,N_23023);
nand U25279 (N_25279,N_22874,N_23588);
nor U25280 (N_25280,N_23889,N_23815);
or U25281 (N_25281,N_23746,N_23298);
nand U25282 (N_25282,N_23035,N_22298);
nor U25283 (N_25283,N_22793,N_23231);
and U25284 (N_25284,N_22937,N_22181);
or U25285 (N_25285,N_22100,N_22249);
nand U25286 (N_25286,N_22414,N_23905);
or U25287 (N_25287,N_22541,N_22677);
nor U25288 (N_25288,N_23917,N_22011);
nand U25289 (N_25289,N_23061,N_23178);
and U25290 (N_25290,N_23724,N_22193);
or U25291 (N_25291,N_22237,N_23580);
nor U25292 (N_25292,N_22784,N_23665);
xnor U25293 (N_25293,N_23014,N_23679);
and U25294 (N_25294,N_22043,N_23604);
nor U25295 (N_25295,N_23388,N_22084);
and U25296 (N_25296,N_23064,N_23686);
and U25297 (N_25297,N_22909,N_22314);
or U25298 (N_25298,N_22472,N_22339);
and U25299 (N_25299,N_22623,N_23818);
nand U25300 (N_25300,N_22079,N_22700);
or U25301 (N_25301,N_23339,N_23458);
and U25302 (N_25302,N_22671,N_22185);
nor U25303 (N_25303,N_23155,N_23395);
and U25304 (N_25304,N_22763,N_23920);
nor U25305 (N_25305,N_23381,N_22281);
nand U25306 (N_25306,N_22323,N_23312);
or U25307 (N_25307,N_23287,N_23237);
xnor U25308 (N_25308,N_23354,N_23512);
or U25309 (N_25309,N_22390,N_23254);
xnor U25310 (N_25310,N_23294,N_22039);
xnor U25311 (N_25311,N_23569,N_22025);
or U25312 (N_25312,N_23256,N_22856);
or U25313 (N_25313,N_23149,N_23609);
or U25314 (N_25314,N_23789,N_22122);
and U25315 (N_25315,N_23948,N_23530);
nand U25316 (N_25316,N_22133,N_23052);
and U25317 (N_25317,N_22988,N_22997);
xnor U25318 (N_25318,N_23812,N_23726);
nor U25319 (N_25319,N_23870,N_23735);
xnor U25320 (N_25320,N_22677,N_22078);
nor U25321 (N_25321,N_23171,N_22118);
nand U25322 (N_25322,N_23980,N_22865);
or U25323 (N_25323,N_22330,N_22975);
and U25324 (N_25324,N_22645,N_22039);
xor U25325 (N_25325,N_22838,N_22176);
xor U25326 (N_25326,N_22212,N_22976);
and U25327 (N_25327,N_22138,N_22276);
and U25328 (N_25328,N_22636,N_22984);
or U25329 (N_25329,N_22939,N_22891);
or U25330 (N_25330,N_22126,N_23658);
or U25331 (N_25331,N_22961,N_23879);
and U25332 (N_25332,N_22069,N_23611);
or U25333 (N_25333,N_22315,N_22066);
nand U25334 (N_25334,N_22806,N_23366);
nor U25335 (N_25335,N_22434,N_23106);
nand U25336 (N_25336,N_23287,N_23451);
nor U25337 (N_25337,N_23860,N_22626);
or U25338 (N_25338,N_23473,N_22572);
nand U25339 (N_25339,N_23715,N_23140);
nand U25340 (N_25340,N_22876,N_23389);
nor U25341 (N_25341,N_23841,N_23720);
and U25342 (N_25342,N_23612,N_23772);
and U25343 (N_25343,N_22760,N_22866);
or U25344 (N_25344,N_23875,N_22012);
or U25345 (N_25345,N_22612,N_22049);
or U25346 (N_25346,N_22853,N_22258);
nor U25347 (N_25347,N_22777,N_23680);
xnor U25348 (N_25348,N_23097,N_22400);
nor U25349 (N_25349,N_22978,N_22000);
xnor U25350 (N_25350,N_23147,N_22560);
xnor U25351 (N_25351,N_23623,N_22886);
nand U25352 (N_25352,N_22083,N_22087);
nor U25353 (N_25353,N_23039,N_23289);
and U25354 (N_25354,N_22008,N_23156);
nor U25355 (N_25355,N_22307,N_22861);
or U25356 (N_25356,N_23642,N_23342);
or U25357 (N_25357,N_22491,N_23355);
xnor U25358 (N_25358,N_23390,N_22227);
nand U25359 (N_25359,N_22817,N_22780);
or U25360 (N_25360,N_22764,N_22462);
or U25361 (N_25361,N_22653,N_22148);
nor U25362 (N_25362,N_22011,N_23488);
nor U25363 (N_25363,N_23837,N_22087);
xnor U25364 (N_25364,N_22452,N_23007);
xor U25365 (N_25365,N_22137,N_23904);
or U25366 (N_25366,N_22846,N_22942);
and U25367 (N_25367,N_22932,N_22752);
and U25368 (N_25368,N_22850,N_22434);
xor U25369 (N_25369,N_22857,N_23890);
xor U25370 (N_25370,N_22387,N_23204);
nand U25371 (N_25371,N_23798,N_23406);
or U25372 (N_25372,N_22257,N_23803);
or U25373 (N_25373,N_23701,N_23838);
and U25374 (N_25374,N_23007,N_22005);
nand U25375 (N_25375,N_22854,N_22153);
nor U25376 (N_25376,N_22903,N_22595);
nand U25377 (N_25377,N_23887,N_22356);
nand U25378 (N_25378,N_23493,N_22928);
nand U25379 (N_25379,N_23246,N_22069);
nor U25380 (N_25380,N_22634,N_23887);
or U25381 (N_25381,N_23704,N_23389);
nor U25382 (N_25382,N_22894,N_23923);
and U25383 (N_25383,N_23795,N_22983);
xnor U25384 (N_25384,N_22529,N_23335);
or U25385 (N_25385,N_23154,N_22803);
xnor U25386 (N_25386,N_23923,N_23005);
nand U25387 (N_25387,N_22781,N_22726);
xor U25388 (N_25388,N_22945,N_23846);
xor U25389 (N_25389,N_23922,N_23493);
xnor U25390 (N_25390,N_23261,N_22168);
or U25391 (N_25391,N_22162,N_23475);
nor U25392 (N_25392,N_22103,N_22323);
nand U25393 (N_25393,N_22374,N_22525);
nor U25394 (N_25394,N_23613,N_23881);
xnor U25395 (N_25395,N_23035,N_23794);
or U25396 (N_25396,N_23877,N_22940);
and U25397 (N_25397,N_23908,N_23490);
or U25398 (N_25398,N_23909,N_23817);
nor U25399 (N_25399,N_22682,N_23548);
xor U25400 (N_25400,N_22617,N_22746);
nor U25401 (N_25401,N_23915,N_23755);
or U25402 (N_25402,N_22887,N_23006);
nor U25403 (N_25403,N_23210,N_23626);
or U25404 (N_25404,N_22515,N_22396);
and U25405 (N_25405,N_23541,N_23981);
and U25406 (N_25406,N_22326,N_22500);
xnor U25407 (N_25407,N_22473,N_23395);
nand U25408 (N_25408,N_23341,N_23308);
and U25409 (N_25409,N_22000,N_22931);
or U25410 (N_25410,N_22255,N_22027);
or U25411 (N_25411,N_23568,N_22485);
or U25412 (N_25412,N_23799,N_22128);
nand U25413 (N_25413,N_23685,N_23051);
xnor U25414 (N_25414,N_23428,N_22022);
or U25415 (N_25415,N_23613,N_23860);
and U25416 (N_25416,N_22392,N_23270);
nor U25417 (N_25417,N_23476,N_22119);
and U25418 (N_25418,N_22281,N_22795);
or U25419 (N_25419,N_22579,N_23038);
xnor U25420 (N_25420,N_23802,N_23435);
nor U25421 (N_25421,N_23463,N_23943);
nor U25422 (N_25422,N_23535,N_23489);
nor U25423 (N_25423,N_23272,N_22397);
or U25424 (N_25424,N_23149,N_22600);
xnor U25425 (N_25425,N_23671,N_23061);
nor U25426 (N_25426,N_22769,N_23624);
xnor U25427 (N_25427,N_22069,N_23516);
or U25428 (N_25428,N_23250,N_23416);
xnor U25429 (N_25429,N_22974,N_22719);
xnor U25430 (N_25430,N_22356,N_22039);
and U25431 (N_25431,N_22673,N_22900);
or U25432 (N_25432,N_23673,N_23473);
nor U25433 (N_25433,N_22454,N_23897);
and U25434 (N_25434,N_22234,N_22917);
nand U25435 (N_25435,N_23752,N_22598);
xor U25436 (N_25436,N_23725,N_23780);
and U25437 (N_25437,N_23352,N_22420);
nor U25438 (N_25438,N_22270,N_22817);
and U25439 (N_25439,N_23372,N_22786);
and U25440 (N_25440,N_23091,N_22943);
xor U25441 (N_25441,N_22311,N_22980);
nand U25442 (N_25442,N_23454,N_22852);
nor U25443 (N_25443,N_22380,N_22669);
nand U25444 (N_25444,N_22674,N_22010);
or U25445 (N_25445,N_23830,N_23443);
nand U25446 (N_25446,N_22402,N_22584);
xor U25447 (N_25447,N_22312,N_22476);
or U25448 (N_25448,N_22381,N_22361);
xor U25449 (N_25449,N_22987,N_23397);
nand U25450 (N_25450,N_22791,N_23662);
nand U25451 (N_25451,N_23573,N_22994);
and U25452 (N_25452,N_22019,N_22972);
and U25453 (N_25453,N_22804,N_23818);
xnor U25454 (N_25454,N_23936,N_22679);
and U25455 (N_25455,N_22332,N_23109);
or U25456 (N_25456,N_22877,N_22971);
and U25457 (N_25457,N_23308,N_23141);
nand U25458 (N_25458,N_22115,N_22186);
nand U25459 (N_25459,N_23519,N_23611);
xor U25460 (N_25460,N_23566,N_22779);
or U25461 (N_25461,N_22120,N_22892);
and U25462 (N_25462,N_22624,N_23990);
or U25463 (N_25463,N_23686,N_23773);
nand U25464 (N_25464,N_22999,N_22756);
xnor U25465 (N_25465,N_23864,N_23779);
or U25466 (N_25466,N_22375,N_23088);
and U25467 (N_25467,N_22979,N_22466);
or U25468 (N_25468,N_22816,N_23528);
and U25469 (N_25469,N_22252,N_22677);
nand U25470 (N_25470,N_23226,N_23294);
nor U25471 (N_25471,N_23436,N_22016);
or U25472 (N_25472,N_23440,N_23536);
xnor U25473 (N_25473,N_23937,N_22315);
nor U25474 (N_25474,N_23420,N_23357);
or U25475 (N_25475,N_22254,N_23334);
nand U25476 (N_25476,N_22996,N_22544);
xnor U25477 (N_25477,N_22954,N_23338);
nand U25478 (N_25478,N_22486,N_22931);
and U25479 (N_25479,N_22135,N_22481);
and U25480 (N_25480,N_22625,N_23662);
nand U25481 (N_25481,N_23277,N_23951);
xnor U25482 (N_25482,N_23339,N_22019);
nand U25483 (N_25483,N_22080,N_22574);
nor U25484 (N_25484,N_22470,N_22878);
or U25485 (N_25485,N_23152,N_23885);
or U25486 (N_25486,N_22642,N_22385);
nand U25487 (N_25487,N_23144,N_22933);
nand U25488 (N_25488,N_23063,N_22010);
xnor U25489 (N_25489,N_23356,N_22487);
and U25490 (N_25490,N_22156,N_22743);
nor U25491 (N_25491,N_22453,N_22074);
nand U25492 (N_25492,N_22547,N_23900);
nand U25493 (N_25493,N_23669,N_22506);
nor U25494 (N_25494,N_22727,N_23326);
nor U25495 (N_25495,N_23821,N_22121);
xnor U25496 (N_25496,N_23663,N_23400);
nor U25497 (N_25497,N_23523,N_23198);
and U25498 (N_25498,N_23428,N_23109);
xnor U25499 (N_25499,N_22357,N_23731);
nor U25500 (N_25500,N_23701,N_23383);
nand U25501 (N_25501,N_22889,N_23272);
and U25502 (N_25502,N_23579,N_23172);
nand U25503 (N_25503,N_23004,N_22625);
and U25504 (N_25504,N_23931,N_23324);
nor U25505 (N_25505,N_22244,N_22313);
or U25506 (N_25506,N_23609,N_23405);
or U25507 (N_25507,N_23113,N_23803);
or U25508 (N_25508,N_22341,N_22895);
nand U25509 (N_25509,N_23061,N_23295);
or U25510 (N_25510,N_23074,N_23800);
nand U25511 (N_25511,N_22072,N_23565);
nor U25512 (N_25512,N_22111,N_22005);
or U25513 (N_25513,N_23600,N_23157);
or U25514 (N_25514,N_23061,N_23371);
and U25515 (N_25515,N_22611,N_22304);
nand U25516 (N_25516,N_22704,N_23911);
nand U25517 (N_25517,N_23611,N_23880);
nor U25518 (N_25518,N_23465,N_22112);
nor U25519 (N_25519,N_23140,N_22991);
xor U25520 (N_25520,N_22535,N_23517);
and U25521 (N_25521,N_22715,N_23805);
nor U25522 (N_25522,N_23032,N_22846);
xnor U25523 (N_25523,N_23405,N_23113);
or U25524 (N_25524,N_23607,N_22327);
and U25525 (N_25525,N_23879,N_23151);
nor U25526 (N_25526,N_23459,N_22091);
xnor U25527 (N_25527,N_22571,N_22898);
and U25528 (N_25528,N_23391,N_22745);
or U25529 (N_25529,N_22894,N_23295);
xor U25530 (N_25530,N_22814,N_23029);
and U25531 (N_25531,N_22076,N_22417);
nand U25532 (N_25532,N_22442,N_22929);
xor U25533 (N_25533,N_22673,N_22201);
nand U25534 (N_25534,N_22338,N_23953);
or U25535 (N_25535,N_22705,N_23497);
nand U25536 (N_25536,N_22455,N_22896);
nor U25537 (N_25537,N_23886,N_22489);
nand U25538 (N_25538,N_23903,N_23925);
nor U25539 (N_25539,N_23770,N_23862);
and U25540 (N_25540,N_23625,N_22550);
nand U25541 (N_25541,N_22574,N_22713);
xnor U25542 (N_25542,N_22134,N_22060);
nand U25543 (N_25543,N_22639,N_22425);
xor U25544 (N_25544,N_23125,N_23787);
and U25545 (N_25545,N_22766,N_22651);
or U25546 (N_25546,N_23989,N_23056);
nor U25547 (N_25547,N_22071,N_23505);
or U25548 (N_25548,N_23673,N_22319);
and U25549 (N_25549,N_23838,N_22066);
xnor U25550 (N_25550,N_23732,N_22663);
or U25551 (N_25551,N_22792,N_22416);
and U25552 (N_25552,N_22259,N_22940);
and U25553 (N_25553,N_22523,N_23245);
xor U25554 (N_25554,N_23072,N_23836);
and U25555 (N_25555,N_22876,N_22623);
nand U25556 (N_25556,N_23260,N_22466);
xor U25557 (N_25557,N_22638,N_22187);
nand U25558 (N_25558,N_22740,N_22629);
or U25559 (N_25559,N_22027,N_22699);
nand U25560 (N_25560,N_23753,N_22119);
and U25561 (N_25561,N_23055,N_23435);
nor U25562 (N_25562,N_23661,N_22024);
xnor U25563 (N_25563,N_22217,N_22156);
xnor U25564 (N_25564,N_22882,N_22082);
or U25565 (N_25565,N_23371,N_23215);
nor U25566 (N_25566,N_22164,N_23006);
nand U25567 (N_25567,N_23235,N_23457);
or U25568 (N_25568,N_22366,N_23853);
or U25569 (N_25569,N_22921,N_22108);
nand U25570 (N_25570,N_23618,N_22766);
nand U25571 (N_25571,N_23964,N_22437);
xnor U25572 (N_25572,N_22705,N_23583);
xnor U25573 (N_25573,N_22166,N_23561);
nor U25574 (N_25574,N_23295,N_22009);
and U25575 (N_25575,N_22702,N_23883);
nor U25576 (N_25576,N_22383,N_22164);
nor U25577 (N_25577,N_23326,N_22720);
nand U25578 (N_25578,N_22597,N_23170);
and U25579 (N_25579,N_22787,N_22409);
or U25580 (N_25580,N_23998,N_23694);
and U25581 (N_25581,N_22919,N_23799);
and U25582 (N_25582,N_22045,N_22268);
xnor U25583 (N_25583,N_22696,N_22724);
and U25584 (N_25584,N_23413,N_22521);
and U25585 (N_25585,N_23609,N_23810);
nand U25586 (N_25586,N_22369,N_23700);
nor U25587 (N_25587,N_22466,N_23240);
nand U25588 (N_25588,N_22345,N_23836);
and U25589 (N_25589,N_23100,N_22516);
xor U25590 (N_25590,N_23978,N_23203);
or U25591 (N_25591,N_22704,N_23445);
nor U25592 (N_25592,N_22204,N_22764);
or U25593 (N_25593,N_22379,N_23557);
nor U25594 (N_25594,N_23292,N_23859);
xnor U25595 (N_25595,N_23735,N_23012);
and U25596 (N_25596,N_23682,N_22579);
nor U25597 (N_25597,N_23890,N_23135);
and U25598 (N_25598,N_23062,N_22998);
or U25599 (N_25599,N_22560,N_23280);
and U25600 (N_25600,N_23388,N_22412);
nand U25601 (N_25601,N_23069,N_22333);
and U25602 (N_25602,N_23549,N_22853);
or U25603 (N_25603,N_23288,N_22517);
and U25604 (N_25604,N_23702,N_22881);
xnor U25605 (N_25605,N_23855,N_23630);
nor U25606 (N_25606,N_22472,N_23331);
and U25607 (N_25607,N_22911,N_22835);
and U25608 (N_25608,N_23500,N_23189);
and U25609 (N_25609,N_23304,N_23780);
nand U25610 (N_25610,N_23445,N_22577);
xor U25611 (N_25611,N_22549,N_22932);
and U25612 (N_25612,N_23176,N_22282);
nor U25613 (N_25613,N_23205,N_22429);
nor U25614 (N_25614,N_22774,N_23250);
xnor U25615 (N_25615,N_23436,N_22679);
nand U25616 (N_25616,N_23126,N_22261);
xnor U25617 (N_25617,N_23568,N_22567);
xnor U25618 (N_25618,N_22851,N_22637);
nor U25619 (N_25619,N_23299,N_23524);
or U25620 (N_25620,N_22064,N_22600);
nand U25621 (N_25621,N_23861,N_23561);
xnor U25622 (N_25622,N_23368,N_23994);
and U25623 (N_25623,N_22573,N_22275);
nor U25624 (N_25624,N_22395,N_23348);
or U25625 (N_25625,N_22196,N_23315);
nand U25626 (N_25626,N_22242,N_22334);
nor U25627 (N_25627,N_23878,N_23718);
nand U25628 (N_25628,N_23650,N_22025);
xnor U25629 (N_25629,N_22095,N_22574);
or U25630 (N_25630,N_22094,N_23593);
nand U25631 (N_25631,N_23783,N_23782);
nand U25632 (N_25632,N_22791,N_23944);
and U25633 (N_25633,N_23600,N_22609);
or U25634 (N_25634,N_22183,N_22683);
nand U25635 (N_25635,N_22255,N_22706);
and U25636 (N_25636,N_22797,N_23990);
xor U25637 (N_25637,N_23010,N_23218);
or U25638 (N_25638,N_23319,N_22540);
and U25639 (N_25639,N_23918,N_23809);
xnor U25640 (N_25640,N_22947,N_22814);
nand U25641 (N_25641,N_23109,N_23817);
nor U25642 (N_25642,N_22178,N_22276);
nor U25643 (N_25643,N_22447,N_23992);
and U25644 (N_25644,N_23690,N_23875);
xor U25645 (N_25645,N_23175,N_23043);
nand U25646 (N_25646,N_23850,N_22593);
xor U25647 (N_25647,N_22053,N_22256);
or U25648 (N_25648,N_22933,N_23103);
nor U25649 (N_25649,N_23009,N_22669);
and U25650 (N_25650,N_23708,N_23972);
nand U25651 (N_25651,N_23498,N_22067);
nor U25652 (N_25652,N_23960,N_22920);
and U25653 (N_25653,N_22563,N_22774);
and U25654 (N_25654,N_23959,N_22717);
or U25655 (N_25655,N_23617,N_23857);
nand U25656 (N_25656,N_23495,N_22209);
nor U25657 (N_25657,N_23124,N_22381);
xnor U25658 (N_25658,N_23244,N_22441);
or U25659 (N_25659,N_22844,N_22334);
nor U25660 (N_25660,N_22520,N_22356);
nand U25661 (N_25661,N_23893,N_23466);
or U25662 (N_25662,N_23237,N_22715);
and U25663 (N_25663,N_23670,N_23391);
or U25664 (N_25664,N_22560,N_22790);
nand U25665 (N_25665,N_23403,N_23944);
and U25666 (N_25666,N_23812,N_22402);
and U25667 (N_25667,N_23514,N_22309);
xor U25668 (N_25668,N_22855,N_22680);
nand U25669 (N_25669,N_23057,N_23867);
nand U25670 (N_25670,N_22908,N_23565);
xor U25671 (N_25671,N_22203,N_22809);
xnor U25672 (N_25672,N_23143,N_22691);
nand U25673 (N_25673,N_23599,N_22049);
nor U25674 (N_25674,N_22625,N_23225);
and U25675 (N_25675,N_22061,N_23700);
xnor U25676 (N_25676,N_23249,N_23455);
nand U25677 (N_25677,N_22060,N_22678);
xor U25678 (N_25678,N_22647,N_23211);
nand U25679 (N_25679,N_23425,N_23683);
xor U25680 (N_25680,N_22865,N_22141);
and U25681 (N_25681,N_23319,N_23485);
or U25682 (N_25682,N_22115,N_23962);
or U25683 (N_25683,N_22999,N_23106);
nand U25684 (N_25684,N_22990,N_22257);
xor U25685 (N_25685,N_22822,N_23047);
nor U25686 (N_25686,N_23385,N_22594);
xor U25687 (N_25687,N_23826,N_23047);
nor U25688 (N_25688,N_23022,N_23126);
and U25689 (N_25689,N_23188,N_22102);
and U25690 (N_25690,N_22225,N_23014);
and U25691 (N_25691,N_22229,N_22078);
xor U25692 (N_25692,N_23870,N_23945);
and U25693 (N_25693,N_23725,N_23934);
or U25694 (N_25694,N_23138,N_23905);
nand U25695 (N_25695,N_22455,N_23156);
nor U25696 (N_25696,N_23996,N_23406);
or U25697 (N_25697,N_22469,N_22232);
nor U25698 (N_25698,N_22160,N_22007);
xnor U25699 (N_25699,N_22866,N_23538);
xnor U25700 (N_25700,N_22164,N_23126);
and U25701 (N_25701,N_23022,N_23257);
or U25702 (N_25702,N_22109,N_23147);
xor U25703 (N_25703,N_22373,N_23677);
or U25704 (N_25704,N_23153,N_22089);
or U25705 (N_25705,N_22962,N_22733);
xor U25706 (N_25706,N_22824,N_22153);
xor U25707 (N_25707,N_23859,N_23493);
nand U25708 (N_25708,N_22656,N_23934);
and U25709 (N_25709,N_23905,N_23154);
nor U25710 (N_25710,N_23744,N_23846);
xnor U25711 (N_25711,N_23826,N_22251);
and U25712 (N_25712,N_22995,N_22348);
or U25713 (N_25713,N_22847,N_23236);
nor U25714 (N_25714,N_22537,N_22599);
nor U25715 (N_25715,N_23294,N_22858);
or U25716 (N_25716,N_23082,N_22956);
and U25717 (N_25717,N_23966,N_22009);
or U25718 (N_25718,N_23290,N_22715);
nand U25719 (N_25719,N_23799,N_22742);
nor U25720 (N_25720,N_23031,N_22990);
and U25721 (N_25721,N_23297,N_23039);
nand U25722 (N_25722,N_23163,N_23555);
xnor U25723 (N_25723,N_23637,N_23434);
nor U25724 (N_25724,N_22489,N_22364);
or U25725 (N_25725,N_23552,N_22538);
xnor U25726 (N_25726,N_23935,N_22157);
and U25727 (N_25727,N_22291,N_23075);
or U25728 (N_25728,N_23754,N_22630);
nor U25729 (N_25729,N_22944,N_22724);
or U25730 (N_25730,N_23795,N_22208);
or U25731 (N_25731,N_23252,N_23801);
or U25732 (N_25732,N_22583,N_22211);
nor U25733 (N_25733,N_22367,N_22500);
xnor U25734 (N_25734,N_23792,N_23355);
nor U25735 (N_25735,N_22241,N_23085);
and U25736 (N_25736,N_22755,N_23539);
or U25737 (N_25737,N_23255,N_23993);
nand U25738 (N_25738,N_23465,N_22443);
or U25739 (N_25739,N_22450,N_22537);
nor U25740 (N_25740,N_23674,N_22070);
and U25741 (N_25741,N_22718,N_22485);
nand U25742 (N_25742,N_22803,N_23028);
and U25743 (N_25743,N_22098,N_22758);
or U25744 (N_25744,N_23999,N_22892);
and U25745 (N_25745,N_22771,N_22241);
or U25746 (N_25746,N_22879,N_22559);
or U25747 (N_25747,N_22560,N_22531);
and U25748 (N_25748,N_22459,N_23270);
and U25749 (N_25749,N_23142,N_23891);
or U25750 (N_25750,N_22182,N_22290);
or U25751 (N_25751,N_23800,N_23836);
nand U25752 (N_25752,N_22478,N_22797);
xor U25753 (N_25753,N_22940,N_23020);
nor U25754 (N_25754,N_22864,N_23466);
nand U25755 (N_25755,N_23546,N_22642);
or U25756 (N_25756,N_23579,N_23161);
and U25757 (N_25757,N_23086,N_23241);
and U25758 (N_25758,N_22169,N_23117);
and U25759 (N_25759,N_23255,N_23136);
nand U25760 (N_25760,N_23411,N_23646);
nand U25761 (N_25761,N_23958,N_22845);
xor U25762 (N_25762,N_22483,N_22974);
xnor U25763 (N_25763,N_23771,N_22649);
xor U25764 (N_25764,N_23538,N_23549);
and U25765 (N_25765,N_22888,N_22223);
nand U25766 (N_25766,N_22626,N_23327);
nand U25767 (N_25767,N_22009,N_22457);
and U25768 (N_25768,N_23298,N_22390);
nand U25769 (N_25769,N_22927,N_22470);
xnor U25770 (N_25770,N_23394,N_22599);
nor U25771 (N_25771,N_23275,N_23964);
nand U25772 (N_25772,N_22716,N_22012);
nor U25773 (N_25773,N_22502,N_23450);
xnor U25774 (N_25774,N_22359,N_22695);
and U25775 (N_25775,N_22715,N_22285);
or U25776 (N_25776,N_23919,N_23311);
xnor U25777 (N_25777,N_22332,N_22577);
or U25778 (N_25778,N_22546,N_22129);
or U25779 (N_25779,N_23483,N_23595);
nor U25780 (N_25780,N_23613,N_22184);
xnor U25781 (N_25781,N_22234,N_22161);
xor U25782 (N_25782,N_23647,N_22595);
and U25783 (N_25783,N_22686,N_22536);
nor U25784 (N_25784,N_22966,N_22565);
xor U25785 (N_25785,N_23148,N_22545);
nand U25786 (N_25786,N_22115,N_23303);
xor U25787 (N_25787,N_22790,N_23649);
and U25788 (N_25788,N_23984,N_23169);
nor U25789 (N_25789,N_23898,N_23864);
nand U25790 (N_25790,N_23741,N_22266);
nand U25791 (N_25791,N_23652,N_23707);
nand U25792 (N_25792,N_22268,N_22557);
nand U25793 (N_25793,N_22355,N_23726);
nand U25794 (N_25794,N_22715,N_23725);
and U25795 (N_25795,N_23963,N_22724);
xnor U25796 (N_25796,N_23673,N_23298);
and U25797 (N_25797,N_23517,N_23293);
xnor U25798 (N_25798,N_22962,N_22479);
nor U25799 (N_25799,N_23503,N_23557);
or U25800 (N_25800,N_22204,N_22305);
and U25801 (N_25801,N_23312,N_23711);
or U25802 (N_25802,N_23839,N_22539);
xor U25803 (N_25803,N_23082,N_23944);
nor U25804 (N_25804,N_22094,N_22993);
nor U25805 (N_25805,N_22300,N_22882);
or U25806 (N_25806,N_23861,N_23997);
nor U25807 (N_25807,N_22446,N_22700);
nand U25808 (N_25808,N_23933,N_22746);
and U25809 (N_25809,N_23923,N_23096);
xnor U25810 (N_25810,N_23296,N_23054);
and U25811 (N_25811,N_22393,N_23950);
nor U25812 (N_25812,N_22176,N_22795);
nand U25813 (N_25813,N_22631,N_23758);
or U25814 (N_25814,N_22236,N_22209);
or U25815 (N_25815,N_23880,N_23609);
and U25816 (N_25816,N_23646,N_22979);
or U25817 (N_25817,N_22577,N_23854);
or U25818 (N_25818,N_23878,N_22251);
xor U25819 (N_25819,N_23792,N_22705);
xnor U25820 (N_25820,N_23043,N_23612);
nand U25821 (N_25821,N_22562,N_22952);
and U25822 (N_25822,N_23450,N_23572);
nor U25823 (N_25823,N_23298,N_22809);
and U25824 (N_25824,N_23103,N_22724);
and U25825 (N_25825,N_23276,N_23203);
nand U25826 (N_25826,N_23796,N_22486);
nand U25827 (N_25827,N_22871,N_23426);
nand U25828 (N_25828,N_22670,N_23811);
and U25829 (N_25829,N_23848,N_22535);
xnor U25830 (N_25830,N_23946,N_22181);
and U25831 (N_25831,N_23970,N_22182);
and U25832 (N_25832,N_22094,N_23386);
and U25833 (N_25833,N_22026,N_23804);
or U25834 (N_25834,N_22259,N_22694);
or U25835 (N_25835,N_23299,N_22991);
nand U25836 (N_25836,N_22596,N_22125);
xor U25837 (N_25837,N_23764,N_22698);
xor U25838 (N_25838,N_23166,N_23275);
xor U25839 (N_25839,N_22264,N_22796);
nor U25840 (N_25840,N_23605,N_22144);
xnor U25841 (N_25841,N_23233,N_22881);
xor U25842 (N_25842,N_23262,N_22619);
xor U25843 (N_25843,N_23761,N_22394);
xnor U25844 (N_25844,N_22766,N_22155);
and U25845 (N_25845,N_23617,N_22474);
nand U25846 (N_25846,N_22975,N_22114);
nand U25847 (N_25847,N_22605,N_22396);
nor U25848 (N_25848,N_23405,N_22360);
nor U25849 (N_25849,N_22657,N_22811);
nand U25850 (N_25850,N_22368,N_23255);
xor U25851 (N_25851,N_23326,N_23691);
nor U25852 (N_25852,N_22274,N_23998);
or U25853 (N_25853,N_22286,N_22084);
nor U25854 (N_25854,N_23834,N_23374);
xor U25855 (N_25855,N_23542,N_23365);
xnor U25856 (N_25856,N_23717,N_22257);
nor U25857 (N_25857,N_22703,N_23497);
and U25858 (N_25858,N_22053,N_22260);
nor U25859 (N_25859,N_22167,N_23538);
nand U25860 (N_25860,N_22850,N_23567);
xnor U25861 (N_25861,N_22182,N_23697);
xnor U25862 (N_25862,N_22512,N_22680);
or U25863 (N_25863,N_22541,N_22665);
or U25864 (N_25864,N_23098,N_22792);
nor U25865 (N_25865,N_23436,N_22983);
or U25866 (N_25866,N_22119,N_23668);
or U25867 (N_25867,N_22772,N_22663);
or U25868 (N_25868,N_22161,N_23283);
or U25869 (N_25869,N_22579,N_23491);
and U25870 (N_25870,N_22974,N_22425);
and U25871 (N_25871,N_22990,N_23082);
or U25872 (N_25872,N_22299,N_23700);
nor U25873 (N_25873,N_23928,N_23601);
and U25874 (N_25874,N_23249,N_22167);
nand U25875 (N_25875,N_22268,N_23681);
or U25876 (N_25876,N_22311,N_23863);
xnor U25877 (N_25877,N_22978,N_22135);
nor U25878 (N_25878,N_22999,N_23556);
xnor U25879 (N_25879,N_23113,N_22915);
nand U25880 (N_25880,N_23796,N_22200);
nor U25881 (N_25881,N_23686,N_23316);
nand U25882 (N_25882,N_23932,N_23642);
nand U25883 (N_25883,N_22797,N_22442);
or U25884 (N_25884,N_22707,N_23178);
or U25885 (N_25885,N_22619,N_22072);
xor U25886 (N_25886,N_23156,N_23833);
nand U25887 (N_25887,N_23400,N_23858);
nand U25888 (N_25888,N_23935,N_22568);
and U25889 (N_25889,N_23669,N_23596);
or U25890 (N_25890,N_23928,N_22645);
nor U25891 (N_25891,N_23836,N_23401);
xor U25892 (N_25892,N_23706,N_23250);
nor U25893 (N_25893,N_22656,N_22227);
or U25894 (N_25894,N_23536,N_22520);
nand U25895 (N_25895,N_22328,N_22427);
nand U25896 (N_25896,N_22408,N_23813);
xnor U25897 (N_25897,N_22869,N_23939);
nor U25898 (N_25898,N_23339,N_23241);
and U25899 (N_25899,N_23212,N_22519);
and U25900 (N_25900,N_23968,N_23766);
and U25901 (N_25901,N_23213,N_23968);
or U25902 (N_25902,N_23361,N_22268);
nand U25903 (N_25903,N_23957,N_22828);
xor U25904 (N_25904,N_23093,N_23057);
nor U25905 (N_25905,N_23919,N_23283);
or U25906 (N_25906,N_23164,N_22194);
or U25907 (N_25907,N_22991,N_23536);
nor U25908 (N_25908,N_22477,N_23057);
xor U25909 (N_25909,N_23352,N_22081);
and U25910 (N_25910,N_23886,N_22939);
nor U25911 (N_25911,N_22423,N_23542);
xor U25912 (N_25912,N_23289,N_23940);
or U25913 (N_25913,N_22482,N_23682);
nor U25914 (N_25914,N_22381,N_23897);
xor U25915 (N_25915,N_23128,N_23266);
or U25916 (N_25916,N_23872,N_23835);
nor U25917 (N_25917,N_22014,N_23555);
or U25918 (N_25918,N_23633,N_22784);
or U25919 (N_25919,N_23251,N_22763);
and U25920 (N_25920,N_22190,N_22763);
nand U25921 (N_25921,N_23111,N_22153);
xor U25922 (N_25922,N_23826,N_22078);
and U25923 (N_25923,N_23019,N_23281);
and U25924 (N_25924,N_23448,N_22831);
nor U25925 (N_25925,N_22234,N_22227);
and U25926 (N_25926,N_23354,N_23233);
xor U25927 (N_25927,N_22107,N_23938);
nor U25928 (N_25928,N_23031,N_22538);
and U25929 (N_25929,N_22078,N_23851);
or U25930 (N_25930,N_22006,N_23392);
nor U25931 (N_25931,N_23052,N_23127);
nand U25932 (N_25932,N_23608,N_22731);
and U25933 (N_25933,N_22500,N_22682);
xnor U25934 (N_25934,N_22841,N_23997);
nand U25935 (N_25935,N_22803,N_22998);
or U25936 (N_25936,N_23555,N_23963);
and U25937 (N_25937,N_23723,N_22092);
nand U25938 (N_25938,N_22572,N_23136);
xnor U25939 (N_25939,N_22873,N_22973);
nand U25940 (N_25940,N_23829,N_22721);
and U25941 (N_25941,N_22069,N_23295);
or U25942 (N_25942,N_23653,N_22604);
nor U25943 (N_25943,N_22340,N_22736);
and U25944 (N_25944,N_23001,N_22645);
or U25945 (N_25945,N_23468,N_23242);
or U25946 (N_25946,N_22409,N_22523);
nand U25947 (N_25947,N_23613,N_23592);
and U25948 (N_25948,N_23917,N_23102);
xor U25949 (N_25949,N_23636,N_23385);
xor U25950 (N_25950,N_22741,N_23742);
nor U25951 (N_25951,N_22160,N_23711);
nor U25952 (N_25952,N_23856,N_23122);
nand U25953 (N_25953,N_23617,N_23344);
and U25954 (N_25954,N_22453,N_23476);
xor U25955 (N_25955,N_23317,N_22206);
nor U25956 (N_25956,N_22229,N_23019);
nor U25957 (N_25957,N_23385,N_23597);
nand U25958 (N_25958,N_22967,N_22892);
nand U25959 (N_25959,N_22820,N_23252);
xor U25960 (N_25960,N_23525,N_23001);
or U25961 (N_25961,N_22711,N_23681);
nor U25962 (N_25962,N_23818,N_22366);
or U25963 (N_25963,N_23000,N_23392);
nor U25964 (N_25964,N_23314,N_23691);
and U25965 (N_25965,N_23529,N_23678);
nand U25966 (N_25966,N_23581,N_22907);
and U25967 (N_25967,N_22136,N_22321);
or U25968 (N_25968,N_23919,N_22169);
and U25969 (N_25969,N_22862,N_23975);
and U25970 (N_25970,N_23442,N_22716);
and U25971 (N_25971,N_23312,N_22976);
nor U25972 (N_25972,N_23169,N_22113);
or U25973 (N_25973,N_23044,N_23266);
or U25974 (N_25974,N_23516,N_22696);
and U25975 (N_25975,N_22352,N_23348);
nor U25976 (N_25976,N_22800,N_23529);
xor U25977 (N_25977,N_22789,N_23231);
and U25978 (N_25978,N_22545,N_22327);
nand U25979 (N_25979,N_22890,N_22034);
xor U25980 (N_25980,N_22360,N_22673);
and U25981 (N_25981,N_23515,N_23401);
xor U25982 (N_25982,N_23051,N_22532);
nand U25983 (N_25983,N_22558,N_22313);
xnor U25984 (N_25984,N_23619,N_23348);
xnor U25985 (N_25985,N_23166,N_22643);
xnor U25986 (N_25986,N_22117,N_22712);
and U25987 (N_25987,N_22757,N_23189);
nand U25988 (N_25988,N_23952,N_22803);
nor U25989 (N_25989,N_22894,N_23905);
nand U25990 (N_25990,N_22929,N_22421);
or U25991 (N_25991,N_23559,N_23745);
or U25992 (N_25992,N_22580,N_22153);
or U25993 (N_25993,N_22300,N_23328);
or U25994 (N_25994,N_22863,N_23999);
nand U25995 (N_25995,N_22962,N_23106);
nor U25996 (N_25996,N_22080,N_23314);
and U25997 (N_25997,N_22965,N_22527);
nand U25998 (N_25998,N_23018,N_22877);
nand U25999 (N_25999,N_23837,N_22483);
and U26000 (N_26000,N_24876,N_25054);
or U26001 (N_26001,N_24034,N_25421);
nand U26002 (N_26002,N_24239,N_24230);
nand U26003 (N_26003,N_24643,N_25380);
nand U26004 (N_26004,N_25858,N_25624);
or U26005 (N_26005,N_24552,N_24833);
xnor U26006 (N_26006,N_24649,N_24258);
or U26007 (N_26007,N_25664,N_25126);
xor U26008 (N_26008,N_25363,N_25899);
nor U26009 (N_26009,N_25639,N_24314);
xor U26010 (N_26010,N_25963,N_25652);
and U26011 (N_26011,N_24826,N_24768);
nand U26012 (N_26012,N_24322,N_25549);
xor U26013 (N_26013,N_24444,N_24486);
or U26014 (N_26014,N_24187,N_25143);
or U26015 (N_26015,N_24896,N_24645);
nand U26016 (N_26016,N_24677,N_24726);
or U26017 (N_26017,N_25879,N_24959);
and U26018 (N_26018,N_24309,N_25718);
and U26019 (N_26019,N_24722,N_24026);
nand U26020 (N_26020,N_25311,N_24977);
xnor U26021 (N_26021,N_24715,N_25589);
xnor U26022 (N_26022,N_25021,N_24687);
or U26023 (N_26023,N_24146,N_24585);
nand U26024 (N_26024,N_25098,N_24805);
or U26025 (N_26025,N_24899,N_24333);
nor U26026 (N_26026,N_24285,N_25086);
or U26027 (N_26027,N_24582,N_24500);
and U26028 (N_26028,N_25558,N_25807);
and U26029 (N_26029,N_25885,N_24114);
and U26030 (N_26030,N_24459,N_24572);
or U26031 (N_26031,N_24694,N_24029);
and U26032 (N_26032,N_24131,N_25369);
or U26033 (N_26033,N_25790,N_25862);
nand U26034 (N_26034,N_24688,N_24147);
nor U26035 (N_26035,N_25156,N_24583);
xnor U26036 (N_26036,N_25288,N_24743);
xnor U26037 (N_26037,N_24617,N_25484);
and U26038 (N_26038,N_24646,N_24033);
xor U26039 (N_26039,N_24702,N_25239);
nand U26040 (N_26040,N_25111,N_25186);
or U26041 (N_26041,N_24375,N_25348);
or U26042 (N_26042,N_24757,N_24987);
nor U26043 (N_26043,N_24671,N_24893);
xnor U26044 (N_26044,N_25245,N_24592);
or U26045 (N_26045,N_24602,N_24944);
and U26046 (N_26046,N_25112,N_24477);
or U26047 (N_26047,N_24410,N_25185);
or U26048 (N_26048,N_25828,N_24838);
nand U26049 (N_26049,N_24596,N_24797);
xor U26050 (N_26050,N_25141,N_24890);
xor U26051 (N_26051,N_24076,N_24004);
and U26052 (N_26052,N_24228,N_24209);
or U26053 (N_26053,N_24847,N_25124);
xnor U26054 (N_26054,N_25896,N_25903);
or U26055 (N_26055,N_24597,N_25454);
nor U26056 (N_26056,N_25315,N_25961);
or U26057 (N_26057,N_25524,N_24629);
nand U26058 (N_26058,N_24243,N_24053);
and U26059 (N_26059,N_25383,N_25056);
nor U26060 (N_26060,N_25527,N_25880);
or U26061 (N_26061,N_24070,N_24553);
xnor U26062 (N_26062,N_24016,N_25563);
nor U26063 (N_26063,N_25600,N_24675);
nand U26064 (N_26064,N_24164,N_24479);
nor U26065 (N_26065,N_24961,N_24599);
nor U26066 (N_26066,N_24122,N_25485);
and U26067 (N_26067,N_25509,N_24383);
nor U26068 (N_26068,N_25620,N_25629);
nand U26069 (N_26069,N_25654,N_25225);
nand U26070 (N_26070,N_25377,N_24268);
nand U26071 (N_26071,N_25048,N_24811);
nand U26072 (N_26072,N_24773,N_24378);
nor U26073 (N_26073,N_24651,N_25672);
and U26074 (N_26074,N_25188,N_25017);
xor U26075 (N_26075,N_25364,N_25476);
nand U26076 (N_26076,N_24161,N_24861);
or U26077 (N_26077,N_24898,N_25950);
xor U26078 (N_26078,N_24021,N_24974);
and U26079 (N_26079,N_24573,N_24973);
or U26080 (N_26080,N_24863,N_24499);
or U26081 (N_26081,N_25260,N_24173);
and U26082 (N_26082,N_24087,N_25276);
or U26083 (N_26083,N_25473,N_25168);
nor U26084 (N_26084,N_24312,N_24919);
nor U26085 (N_26085,N_25180,N_25166);
nand U26086 (N_26086,N_25971,N_24823);
or U26087 (N_26087,N_25169,N_24766);
nand U26088 (N_26088,N_24384,N_24918);
nor U26089 (N_26089,N_24999,N_24819);
and U26090 (N_26090,N_25058,N_25118);
nand U26091 (N_26091,N_25341,N_25779);
xnor U26092 (N_26092,N_25844,N_24767);
and U26093 (N_26093,N_24222,N_25660);
nor U26094 (N_26094,N_24020,N_24468);
xnor U26095 (N_26095,N_25065,N_24374);
and U26096 (N_26096,N_25516,N_24681);
xnor U26097 (N_26097,N_25131,N_25465);
nor U26098 (N_26098,N_25104,N_25583);
and U26099 (N_26099,N_25955,N_24357);
nor U26100 (N_26100,N_24392,N_24947);
or U26101 (N_26101,N_25511,N_24879);
and U26102 (N_26102,N_24699,N_25217);
nand U26103 (N_26103,N_24614,N_25748);
nor U26104 (N_26104,N_25756,N_25998);
xor U26105 (N_26105,N_25174,N_25740);
nor U26106 (N_26106,N_24754,N_25929);
nor U26107 (N_26107,N_24492,N_25940);
nand U26108 (N_26108,N_25145,N_25344);
nor U26109 (N_26109,N_24178,N_24380);
nor U26110 (N_26110,N_24779,N_24298);
nand U26111 (N_26111,N_24902,N_25890);
and U26112 (N_26112,N_25148,N_24249);
nand U26113 (N_26113,N_25800,N_25269);
xnor U26114 (N_26114,N_24443,N_25373);
or U26115 (N_26115,N_25401,N_25954);
or U26116 (N_26116,N_24104,N_24707);
nor U26117 (N_26117,N_24784,N_25384);
nand U26118 (N_26118,N_25456,N_25044);
and U26119 (N_26119,N_24081,N_24856);
nand U26120 (N_26120,N_25435,N_24551);
nor U26121 (N_26121,N_24657,N_25817);
nand U26122 (N_26122,N_24493,N_24296);
or U26123 (N_26123,N_25477,N_24134);
xnor U26124 (N_26124,N_25713,N_24434);
xor U26125 (N_26125,N_25095,N_24512);
xnor U26126 (N_26126,N_24578,N_24690);
xor U26127 (N_26127,N_24090,N_25888);
xnor U26128 (N_26128,N_24262,N_25229);
or U26129 (N_26129,N_25392,N_25281);
or U26130 (N_26130,N_25760,N_24284);
nor U26131 (N_26131,N_24831,N_24264);
nor U26132 (N_26132,N_24470,N_24858);
nand U26133 (N_26133,N_24611,N_24247);
nor U26134 (N_26134,N_24372,N_24039);
nand U26135 (N_26135,N_24860,N_24825);
nand U26136 (N_26136,N_24608,N_25324);
nand U26137 (N_26137,N_24514,N_24884);
nor U26138 (N_26138,N_25327,N_25925);
and U26139 (N_26139,N_25924,N_25525);
nor U26140 (N_26140,N_24658,N_24320);
and U26141 (N_26141,N_24814,N_24982);
nor U26142 (N_26142,N_25000,N_25182);
nor U26143 (N_26143,N_25317,N_24027);
nor U26144 (N_26144,N_25633,N_24478);
xnor U26145 (N_26145,N_25034,N_25866);
nor U26146 (N_26146,N_24813,N_24742);
nor U26147 (N_26147,N_24108,N_24046);
nand U26148 (N_26148,N_24673,N_25016);
xnor U26149 (N_26149,N_24975,N_25043);
nor U26150 (N_26150,N_24338,N_24442);
nand U26151 (N_26151,N_25627,N_24416);
or U26152 (N_26152,N_25912,N_25486);
or U26153 (N_26153,N_24621,N_25611);
and U26154 (N_26154,N_24267,N_24618);
nand U26155 (N_26155,N_24171,N_24121);
nor U26156 (N_26156,N_24331,N_25191);
nor U26157 (N_26157,N_25948,N_25018);
xor U26158 (N_26158,N_25794,N_25003);
xnor U26159 (N_26159,N_25825,N_25334);
xor U26160 (N_26160,N_25662,N_24462);
or U26161 (N_26161,N_25602,N_25258);
or U26162 (N_26162,N_25496,N_24356);
nor U26163 (N_26163,N_24749,N_25009);
xor U26164 (N_26164,N_25444,N_24855);
xor U26165 (N_26165,N_24849,N_25801);
nor U26166 (N_26166,N_25299,N_25049);
xnor U26167 (N_26167,N_25780,N_24783);
and U26168 (N_26168,N_25962,N_25426);
nor U26169 (N_26169,N_25412,N_25423);
or U26170 (N_26170,N_25855,N_25883);
nor U26171 (N_26171,N_25554,N_25079);
nand U26172 (N_26172,N_25626,N_24865);
xnor U26173 (N_26173,N_25908,N_24349);
nand U26174 (N_26174,N_25920,N_24924);
nor U26175 (N_26175,N_24625,N_25552);
or U26176 (N_26176,N_24463,N_25400);
nor U26177 (N_26177,N_25673,N_25028);
nor U26178 (N_26178,N_25943,N_25262);
and U26179 (N_26179,N_25861,N_25005);
nand U26180 (N_26180,N_25694,N_25247);
or U26181 (N_26181,N_25592,N_24185);
or U26182 (N_26182,N_24613,N_24190);
nand U26183 (N_26183,N_24232,N_25551);
nor U26184 (N_26184,N_24659,N_25804);
nor U26185 (N_26185,N_25041,N_25415);
nand U26186 (N_26186,N_25574,N_24853);
nor U26187 (N_26187,N_24964,N_24841);
xor U26188 (N_26188,N_25622,N_24064);
and U26189 (N_26189,N_24052,N_25455);
or U26190 (N_26190,N_24518,N_24759);
nor U26191 (N_26191,N_24755,N_24691);
and U26192 (N_26192,N_24705,N_24979);
xnor U26193 (N_26193,N_24238,N_24904);
or U26194 (N_26194,N_25538,N_24875);
and U26195 (N_26195,N_25987,N_24438);
or U26196 (N_26196,N_24487,N_25613);
nor U26197 (N_26197,N_24830,N_24246);
xnor U26198 (N_26198,N_25176,N_24288);
xnor U26199 (N_26199,N_24764,N_25766);
nor U26200 (N_26200,N_25046,N_25212);
and U26201 (N_26201,N_25057,N_24778);
or U26202 (N_26202,N_25337,N_25120);
nand U26203 (N_26203,N_24335,N_24516);
nand U26204 (N_26204,N_25936,N_24665);
and U26205 (N_26205,N_25097,N_24397);
xnor U26206 (N_26206,N_25474,N_25750);
or U26207 (N_26207,N_25437,N_25832);
or U26208 (N_26208,N_24686,N_25884);
xnor U26209 (N_26209,N_24195,N_25055);
nor U26210 (N_26210,N_25150,N_25729);
xnor U26211 (N_26211,N_25733,N_25578);
nor U26212 (N_26212,N_25158,N_25062);
and U26213 (N_26213,N_24808,N_24461);
nor U26214 (N_26214,N_24447,N_24120);
or U26215 (N_26215,N_24682,N_25507);
or U26216 (N_26216,N_24054,N_24628);
and U26217 (N_26217,N_25572,N_25906);
or U26218 (N_26218,N_25960,N_24747);
nand U26219 (N_26219,N_25784,N_25234);
nand U26220 (N_26220,N_25264,N_25916);
and U26221 (N_26221,N_24379,N_25209);
and U26222 (N_26222,N_24310,N_25901);
nor U26223 (N_26223,N_25081,N_25585);
nor U26224 (N_26224,N_24940,N_25618);
or U26225 (N_26225,N_25710,N_25036);
nor U26226 (N_26226,N_24005,N_25134);
nand U26227 (N_26227,N_24359,N_24454);
xor U26228 (N_26228,N_24780,N_25952);
or U26229 (N_26229,N_24640,N_25490);
nor U26230 (N_26230,N_24425,N_24086);
or U26231 (N_26231,N_25391,N_24482);
nand U26232 (N_26232,N_24988,N_24736);
nor U26233 (N_26233,N_24012,N_24261);
xnor U26234 (N_26234,N_24018,N_25555);
or U26235 (N_26235,N_25278,N_24801);
nand U26236 (N_26236,N_24377,N_25653);
nor U26237 (N_26237,N_25445,N_25153);
nor U26238 (N_26238,N_25932,N_25214);
and U26239 (N_26239,N_25656,N_24762);
nand U26240 (N_26240,N_25184,N_25202);
and U26241 (N_26241,N_25193,N_24517);
xor U26242 (N_26242,N_25787,N_25067);
xor U26243 (N_26243,N_25997,N_24422);
nor U26244 (N_26244,N_24326,N_25135);
nand U26245 (N_26245,N_25689,N_24174);
and U26246 (N_26246,N_25039,N_24913);
nand U26247 (N_26247,N_25235,N_25601);
nand U26248 (N_26248,N_24827,N_24570);
and U26249 (N_26249,N_25146,N_25501);
or U26250 (N_26250,N_24107,N_24689);
nor U26251 (N_26251,N_24241,N_24935);
xor U26252 (N_26252,N_25568,N_25290);
nand U26253 (N_26253,N_24501,N_25744);
nand U26254 (N_26254,N_25007,N_25181);
nand U26255 (N_26255,N_24221,N_24182);
and U26256 (N_26256,N_25418,N_24450);
or U26257 (N_26257,N_25510,N_25404);
and U26258 (N_26258,N_25138,N_25721);
nor U26259 (N_26259,N_25297,N_25014);
or U26260 (N_26260,N_25390,N_24369);
and U26261 (N_26261,N_25590,N_25667);
nor U26262 (N_26262,N_24166,N_24236);
or U26263 (N_26263,N_25697,N_25408);
and U26264 (N_26264,N_25060,N_25514);
nand U26265 (N_26265,N_24972,N_24844);
nand U26266 (N_26266,N_25597,N_24574);
or U26267 (N_26267,N_24073,N_25941);
nor U26268 (N_26268,N_25416,N_24579);
xor U26269 (N_26269,N_25831,N_25078);
nor U26270 (N_26270,N_24138,N_24231);
and U26271 (N_26271,N_25478,N_25090);
xnor U26272 (N_26272,N_24328,N_24672);
and U26273 (N_26273,N_24539,N_24725);
nand U26274 (N_26274,N_25868,N_24537);
and U26275 (N_26275,N_25252,N_24911);
nor U26276 (N_26276,N_25096,N_25805);
and U26277 (N_26277,N_24002,N_24325);
or U26278 (N_26278,N_24466,N_24734);
and U26279 (N_26279,N_24346,N_25547);
or U26280 (N_26280,N_25215,N_25417);
or U26281 (N_26281,N_24183,N_25244);
and U26282 (N_26282,N_24273,N_25035);
xnor U26283 (N_26283,N_24339,N_25722);
nor U26284 (N_26284,N_25351,N_24216);
nor U26285 (N_26285,N_24943,N_25900);
or U26286 (N_26286,N_25368,N_25686);
nor U26287 (N_26287,N_24215,N_25761);
nor U26288 (N_26288,N_24367,N_24735);
xnor U26289 (N_26289,N_24733,N_24057);
or U26290 (N_26290,N_25342,N_24103);
or U26291 (N_26291,N_24280,N_25882);
or U26292 (N_26292,N_25339,N_25599);
xor U26293 (N_26293,N_25714,N_25848);
nor U26294 (N_26294,N_24269,N_25892);
nand U26295 (N_26295,N_24083,N_24718);
xnor U26296 (N_26296,N_24127,N_24632);
nand U26297 (N_26297,N_24474,N_25038);
or U26298 (N_26298,N_24253,N_24945);
xor U26299 (N_26299,N_24028,N_25999);
and U26300 (N_26300,N_24206,N_25949);
or U26301 (N_26301,N_25372,N_24564);
xnor U26302 (N_26302,N_25291,N_25909);
and U26303 (N_26303,N_24765,N_25399);
nor U26304 (N_26304,N_25468,N_24839);
nor U26305 (N_26305,N_24900,N_24732);
nand U26306 (N_26306,N_25436,N_24561);
nor U26307 (N_26307,N_24914,N_25967);
nand U26308 (N_26308,N_24697,N_24878);
xor U26309 (N_26309,N_24229,N_25641);
xor U26310 (N_26310,N_25438,N_24641);
xnor U26311 (N_26311,N_25091,N_24023);
xnor U26312 (N_26312,N_24199,N_25815);
and U26313 (N_26313,N_25338,N_24740);
xor U26314 (N_26314,N_24398,N_25946);
xor U26315 (N_26315,N_25210,N_25329);
and U26316 (N_26316,N_25797,N_25117);
and U26317 (N_26317,N_25226,N_24006);
nor U26318 (N_26318,N_25811,N_25040);
xnor U26319 (N_26319,N_24106,N_24816);
and U26320 (N_26320,N_25560,N_25764);
nor U26321 (N_26321,N_24361,N_24627);
or U26322 (N_26322,N_25052,N_25647);
xnor U26323 (N_26323,N_24150,N_25576);
xnor U26324 (N_26324,N_25864,N_25521);
nor U26325 (N_26325,N_25777,N_24846);
nor U26326 (N_26326,N_24730,N_24317);
nor U26327 (N_26327,N_25781,N_25991);
xor U26328 (N_26328,N_25984,N_25298);
nor U26329 (N_26329,N_24761,N_24036);
xnor U26330 (N_26330,N_25776,N_25050);
nor U26331 (N_26331,N_25289,N_24927);
xor U26332 (N_26332,N_24109,N_24874);
or U26333 (N_26333,N_25751,N_24154);
nand U26334 (N_26334,N_24311,N_25887);
nor U26335 (N_26335,N_25758,N_25803);
and U26336 (N_26336,N_25856,N_24424);
and U26337 (N_26337,N_24030,N_24414);
and U26338 (N_26338,N_25757,N_24217);
and U26339 (N_26339,N_24967,N_25813);
or U26340 (N_26340,N_25691,N_25282);
nor U26341 (N_26341,N_24031,N_25615);
and U26342 (N_26342,N_24639,N_24817);
or U26343 (N_26343,N_24464,N_25886);
or U26344 (N_26344,N_25237,N_24695);
nor U26345 (N_26345,N_24000,N_25569);
and U26346 (N_26346,N_24556,N_25816);
and U26347 (N_26347,N_25637,N_24044);
nor U26348 (N_26348,N_24213,N_25814);
nand U26349 (N_26349,N_25025,N_24316);
or U26350 (N_26350,N_25587,N_24101);
and U26351 (N_26351,N_24685,N_24297);
nand U26352 (N_26352,N_25575,N_25115);
nor U26353 (N_26353,N_24295,N_25072);
or U26354 (N_26354,N_24786,N_25688);
xnor U26355 (N_26355,N_25254,N_24088);
nand U26356 (N_26356,N_25727,N_25769);
or U26357 (N_26357,N_25499,N_25240);
nor U26358 (N_26358,N_24340,N_25246);
nor U26359 (N_26359,N_24022,N_25361);
nand U26360 (N_26360,N_25645,N_24832);
xor U26361 (N_26361,N_25623,N_25222);
nand U26362 (N_26362,N_25631,N_25434);
and U26363 (N_26363,N_25083,N_24289);
nand U26364 (N_26364,N_25670,N_25846);
nor U26365 (N_26365,N_24144,N_24737);
and U26366 (N_26366,N_25376,N_24452);
nor U26367 (N_26367,N_25671,N_24151);
nand U26368 (N_26368,N_25241,N_24393);
and U26369 (N_26369,N_25253,N_25261);
nand U26370 (N_26370,N_25165,N_25394);
or U26371 (N_26371,N_25989,N_25230);
and U26372 (N_26372,N_24777,N_25544);
nor U26373 (N_26373,N_25894,N_24938);
nand U26374 (N_26374,N_24113,N_24793);
nor U26375 (N_26375,N_24888,N_25959);
and U26376 (N_26376,N_24547,N_24094);
nand U26377 (N_26377,N_25023,N_25658);
nand U26378 (N_26378,N_25649,N_24038);
xor U26379 (N_26379,N_25708,N_24660);
xnor U26380 (N_26380,N_25773,N_25965);
nand U26381 (N_26381,N_25255,N_25783);
nand U26382 (N_26382,N_25518,N_24042);
xor U26383 (N_26383,N_25678,N_25177);
and U26384 (N_26384,N_25251,N_24433);
nand U26385 (N_26385,N_24409,N_24062);
xor U26386 (N_26386,N_25100,N_24214);
and U26387 (N_26387,N_24007,N_25915);
nand U26388 (N_26388,N_24901,N_24746);
xnor U26389 (N_26389,N_25529,N_25318);
or U26390 (N_26390,N_24319,N_25666);
or U26391 (N_26391,N_25319,N_25632);
or U26392 (N_26392,N_25314,N_25405);
and U26393 (N_26393,N_24612,N_24917);
nor U26394 (N_26394,N_25881,N_25810);
xnor U26395 (N_26395,N_25010,N_24491);
xor U26396 (N_26396,N_24403,N_24594);
xnor U26397 (N_26397,N_25119,N_24412);
and U26398 (N_26398,N_25029,N_25735);
or U26399 (N_26399,N_24820,N_25307);
nand U26400 (N_26400,N_24008,N_25231);
nand U26401 (N_26401,N_25731,N_25517);
nor U26402 (N_26402,N_25755,N_25559);
nor U26403 (N_26403,N_24949,N_24413);
nand U26404 (N_26404,N_24197,N_25248);
nand U26405 (N_26405,N_24729,N_24420);
or U26406 (N_26406,N_25681,N_24915);
or U26407 (N_26407,N_25675,N_25788);
nor U26408 (N_26408,N_24644,N_24449);
nand U26409 (N_26409,N_25461,N_25413);
or U26410 (N_26410,N_25995,N_25836);
or U26411 (N_26411,N_24279,N_24652);
and U26412 (N_26412,N_24727,N_24177);
nand U26413 (N_26413,N_25084,N_25063);
nor U26414 (N_26414,N_24345,N_24347);
xnor U26415 (N_26415,N_24948,N_24758);
nand U26416 (N_26416,N_24721,N_24794);
or U26417 (N_26417,N_25316,N_25604);
or U26418 (N_26418,N_24437,N_25108);
nor U26419 (N_26419,N_25266,N_25103);
nor U26420 (N_26420,N_24524,N_25619);
or U26421 (N_26421,N_24664,N_25716);
xor U26422 (N_26422,N_25360,N_24648);
nand U26423 (N_26423,N_25522,N_25020);
or U26424 (N_26424,N_24872,N_24274);
nor U26425 (N_26425,N_24984,N_25492);
xor U26426 (N_26426,N_25355,N_24427);
or U26427 (N_26427,N_24763,N_25481);
and U26428 (N_26428,N_25852,N_24698);
or U26429 (N_26429,N_24489,N_24870);
nor U26430 (N_26430,N_24851,N_24966);
nand U26431 (N_26431,N_25411,N_24490);
xor U26432 (N_26432,N_25580,N_25139);
xnor U26433 (N_26433,N_25132,N_24848);
nor U26434 (N_26434,N_25452,N_25286);
and U26435 (N_26435,N_25957,N_24994);
and U26436 (N_26436,N_25066,N_25699);
xnor U26437 (N_26437,N_25424,N_24877);
nor U26438 (N_26438,N_25889,N_24590);
or U26439 (N_26439,N_24526,N_25487);
and U26440 (N_26440,N_25154,N_24198);
xor U26441 (N_26441,N_24871,N_24511);
nand U26442 (N_26442,N_25616,N_25561);
nand U26443 (N_26443,N_25149,N_24986);
nor U26444 (N_26444,N_24969,N_24277);
or U26445 (N_26445,N_25179,N_25512);
nand U26446 (N_26446,N_25059,N_24061);
and U26447 (N_26447,N_24523,N_24475);
xor U26448 (N_26448,N_24205,N_25853);
nand U26449 (N_26449,N_24857,N_25228);
or U26450 (N_26450,N_25087,N_25388);
xnor U26451 (N_26451,N_25042,N_24591);
and U26452 (N_26452,N_24769,N_25820);
or U26453 (N_26453,N_24250,N_24429);
nor U26454 (N_26454,N_24933,N_25498);
or U26455 (N_26455,N_25533,N_25293);
nand U26456 (N_26456,N_24441,N_24647);
and U26457 (N_26457,N_24287,N_24990);
nand U26458 (N_26458,N_25859,N_24344);
nand U26459 (N_26459,N_25128,N_24674);
nand U26460 (N_26460,N_24162,N_24050);
and U26461 (N_26461,N_25564,N_24668);
xor U26462 (N_26462,N_24436,N_24092);
or U26463 (N_26463,N_24294,N_25593);
nand U26464 (N_26464,N_25717,N_24498);
nor U26465 (N_26465,N_25806,N_25553);
nor U26466 (N_26466,N_24744,N_25596);
or U26467 (N_26467,N_25285,N_25113);
nand U26468 (N_26468,N_25505,N_25579);
or U26469 (N_26469,N_24321,N_25753);
nor U26470 (N_26470,N_25796,N_25284);
nand U26471 (N_26471,N_25294,N_25562);
or U26472 (N_26472,N_24840,N_25431);
xor U26473 (N_26473,N_25819,N_24515);
or U26474 (N_26474,N_25930,N_24510);
or U26475 (N_26475,N_25144,N_25397);
nor U26476 (N_26476,N_25107,N_24428);
and U26477 (N_26477,N_24237,N_24327);
and U26478 (N_26478,N_25199,N_24167);
and U26479 (N_26479,N_24032,N_24983);
nand U26480 (N_26480,N_25459,N_24529);
or U26481 (N_26481,N_24041,N_25875);
or U26482 (N_26482,N_25163,N_24776);
nand U26483 (N_26483,N_24196,N_24824);
or U26484 (N_26484,N_24728,N_24003);
nand U26485 (N_26485,N_24165,N_24318);
xor U26486 (N_26486,N_25292,N_25939);
nand U26487 (N_26487,N_25835,N_24532);
or U26488 (N_26488,N_24502,N_24669);
nor U26489 (N_26489,N_24907,N_25441);
nor U26490 (N_26490,N_25387,N_25798);
and U26491 (N_26491,N_24605,N_24724);
xor U26492 (N_26492,N_24882,N_24191);
and U26493 (N_26493,N_25402,N_25603);
and U26494 (N_26494,N_24388,N_25051);
xor U26495 (N_26495,N_25378,N_24802);
or U26496 (N_26496,N_24105,N_24921);
and U26497 (N_26497,N_24895,N_24624);
nor U26498 (N_26498,N_24139,N_25162);
or U26499 (N_26499,N_24219,N_24148);
or U26500 (N_26500,N_24391,N_25366);
nor U26501 (N_26501,N_25981,N_24152);
or U26502 (N_26502,N_25406,N_25935);
nor U26503 (N_26503,N_24184,N_25271);
and U26504 (N_26504,N_24473,N_24791);
or U26505 (N_26505,N_24928,N_24978);
or U26506 (N_26506,N_24399,N_25674);
nor U26507 (N_26507,N_25427,N_25898);
nor U26508 (N_26508,N_24670,N_25537);
and U26509 (N_26509,N_25546,N_25614);
nor U26510 (N_26510,N_24343,N_24916);
and U26511 (N_26511,N_25871,N_25542);
nand U26512 (N_26512,N_25734,N_25157);
xor U26513 (N_26513,N_25082,N_24804);
or U26514 (N_26514,N_24063,N_24661);
xnor U26515 (N_26515,N_24126,N_24586);
nand U26516 (N_26516,N_25609,N_25565);
nor U26517 (N_26517,N_24263,N_25595);
nor U26518 (N_26518,N_24577,N_25964);
xnor U26519 (N_26519,N_24980,N_24351);
nor U26520 (N_26520,N_25818,N_25792);
and U26521 (N_26521,N_24760,N_25704);
or U26522 (N_26522,N_25515,N_24976);
xor U26523 (N_26523,N_24620,N_25918);
and U26524 (N_26524,N_24019,N_25979);
nor U26525 (N_26525,N_25720,N_25171);
nor U26526 (N_26526,N_24565,N_24130);
nand U26527 (N_26527,N_24534,N_25089);
and U26528 (N_26528,N_24533,N_25470);
nor U26529 (N_26529,N_25543,N_24432);
or U26530 (N_26530,N_24954,N_25743);
and U26531 (N_26531,N_24010,N_24503);
nor U26532 (N_26532,N_25904,N_24955);
xnor U26533 (N_26533,N_25765,N_25302);
or U26534 (N_26534,N_25706,N_24259);
or U26535 (N_26535,N_24204,N_24203);
or U26536 (N_26536,N_24281,N_24275);
or U26537 (N_26537,N_24854,N_25483);
nand U26538 (N_26538,N_25011,N_25243);
and U26539 (N_26539,N_25677,N_25536);
or U26540 (N_26540,N_24157,N_24456);
xor U26541 (N_26541,N_24807,N_24806);
nand U26542 (N_26542,N_25323,N_25545);
nand U26543 (N_26543,N_25775,N_24912);
nand U26544 (N_26544,N_25359,N_25321);
or U26545 (N_26545,N_24623,N_24421);
xor U26546 (N_26546,N_24775,N_24936);
xor U26547 (N_26547,N_25175,N_24024);
nor U26548 (N_26548,N_25187,N_25953);
nor U26549 (N_26549,N_24886,N_25736);
and U26550 (N_26550,N_25114,N_25008);
and U26551 (N_26551,N_24040,N_24226);
nor U26552 (N_26552,N_25102,N_24283);
or U26553 (N_26553,N_24810,N_25869);
and U26554 (N_26554,N_25793,N_25863);
xnor U26555 (N_26555,N_24782,N_25428);
xnor U26556 (N_26556,N_25330,N_25106);
xnor U26557 (N_26557,N_24894,N_24115);
or U26558 (N_26558,N_25080,N_25069);
xnor U26559 (N_26559,N_25197,N_24342);
and U26560 (N_26560,N_24557,N_24772);
nor U26561 (N_26561,N_24607,N_25306);
xor U26562 (N_26562,N_24123,N_24546);
nand U26563 (N_26563,N_24080,N_25914);
and U26564 (N_26564,N_25571,N_24324);
and U26565 (N_26565,N_25480,N_25343);
nor U26566 (N_26566,N_24635,N_24981);
nand U26567 (N_26567,N_24423,N_24371);
or U26568 (N_26568,N_25259,N_25759);
xnor U26569 (N_26569,N_25450,N_25024);
or U26570 (N_26570,N_25208,N_24696);
xor U26571 (N_26571,N_25782,N_24835);
and U26572 (N_26572,N_24352,N_25679);
and U26573 (N_26573,N_24991,N_25636);
or U26574 (N_26574,N_25968,N_25463);
and U26575 (N_26575,N_24926,N_25635);
xor U26576 (N_26576,N_24156,N_24353);
xnor U26577 (N_26577,N_25328,N_25830);
and U26578 (N_26578,N_25370,N_25164);
or U26579 (N_26579,N_24842,N_24234);
nand U26580 (N_26580,N_24852,N_25786);
nor U26581 (N_26581,N_24667,N_24125);
or U26582 (N_26582,N_24227,N_24155);
or U26583 (N_26583,N_24270,N_24606);
and U26584 (N_26584,N_24440,N_25076);
and U26585 (N_26585,N_25471,N_24102);
nor U26586 (N_26586,N_24430,N_25207);
nand U26587 (N_26587,N_24738,N_24713);
or U26588 (N_26588,N_24680,N_25839);
nand U26589 (N_26589,N_25019,N_24941);
nand U26590 (N_26590,N_25206,N_25350);
nor U26591 (N_26591,N_24829,N_25151);
or U26592 (N_26592,N_25745,N_24934);
nor U26593 (N_26593,N_25978,N_24293);
xor U26594 (N_26594,N_24531,N_25194);
and U26595 (N_26595,N_24937,N_24997);
nand U26596 (N_26596,N_24282,N_24548);
xor U26597 (N_26597,N_24058,N_25927);
nor U26598 (N_26598,N_25785,N_25313);
xor U26599 (N_26599,N_24306,N_25687);
nor U26600 (N_26600,N_25396,N_24741);
or U26601 (N_26601,N_24431,N_25466);
nor U26602 (N_26602,N_24223,N_24701);
nand U26603 (N_26603,N_25429,N_25250);
nand U26604 (N_26604,N_24211,N_25335);
nand U26605 (N_26605,N_25870,N_25556);
nor U26606 (N_26606,N_24559,N_25249);
xor U26607 (N_26607,N_25728,N_24480);
nand U26608 (N_26608,N_25448,N_24931);
or U26609 (N_26609,N_25309,N_24542);
nor U26610 (N_26610,N_24993,N_24084);
nand U26611 (N_26611,N_25257,N_24789);
and U26612 (N_26612,N_25723,N_25737);
or U26613 (N_26613,N_24560,N_25502);
nor U26614 (N_26614,N_25500,N_24684);
or U26615 (N_26615,N_24538,N_25488);
and U26616 (N_26616,N_25911,N_25845);
and U26617 (N_26617,N_25030,N_24481);
or U26618 (N_26618,N_25557,N_25274);
nor U26619 (N_26619,N_24530,N_25956);
xnor U26620 (N_26620,N_24111,N_24089);
nand U26621 (N_26621,N_25532,N_25354);
and U26622 (N_26622,N_24909,N_24957);
or U26623 (N_26623,N_24390,N_25389);
nand U26624 (N_26624,N_24601,N_24989);
nor U26625 (N_26625,N_25190,N_24880);
and U26626 (N_26626,N_24001,N_24843);
nand U26627 (N_26627,N_24535,N_24992);
nor U26628 (N_26628,N_25232,N_24129);
nand U26629 (N_26629,N_24809,N_25891);
nand U26630 (N_26630,N_25643,N_24836);
and U26631 (N_26631,N_25178,N_24603);
nor U26632 (N_26632,N_25410,N_24091);
nor U26633 (N_26633,N_25567,N_24400);
nor U26634 (N_26634,N_24364,N_24653);
and U26635 (N_26635,N_25746,N_24567);
nand U26636 (N_26636,N_25926,N_24868);
xor U26637 (N_26637,N_25322,N_24097);
or U26638 (N_26638,N_24488,N_24133);
nor U26639 (N_26639,N_24235,N_25213);
xor U26640 (N_26640,N_24071,N_25917);
xor U26641 (N_26641,N_24099,N_24453);
xor U26642 (N_26642,N_24082,N_24043);
and U26643 (N_26643,N_25850,N_24278);
or U26644 (N_26644,N_24188,N_24469);
nor U26645 (N_26645,N_25218,N_24407);
and U26646 (N_26646,N_25331,N_24971);
nand U26647 (N_26647,N_25287,N_24207);
nor U26648 (N_26648,N_25923,N_24595);
and U26649 (N_26649,N_24355,N_24812);
or U26650 (N_26650,N_25277,N_25447);
and U26651 (N_26651,N_24609,N_25045);
nand U26652 (N_26652,N_24011,N_24093);
nor U26653 (N_26653,N_25129,N_25657);
xor U26654 (N_26654,N_24376,N_25770);
xnor U26655 (N_26655,N_25136,N_24704);
nor U26656 (N_26656,N_25088,N_25340);
and U26657 (N_26657,N_24850,N_25336);
or U26658 (N_26658,N_25742,N_25462);
xnor U26659 (N_26659,N_25665,N_25977);
xor U26660 (N_26660,N_25865,N_25692);
and U26661 (N_26661,N_25655,N_24405);
xnor U26662 (N_26662,N_25910,N_25789);
and U26663 (N_26663,N_24580,N_24785);
xnor U26664 (N_26664,N_25983,N_24569);
nor U26665 (N_26665,N_25548,N_25446);
or U26666 (N_26666,N_24796,N_25305);
nand U26667 (N_26667,N_25715,N_25508);
and U26668 (N_26668,N_24303,N_24159);
xnor U26669 (N_26669,N_25907,N_25774);
and U26670 (N_26670,N_25823,N_24170);
xnor U26671 (N_26671,N_25333,N_24276);
nand U26672 (N_26672,N_25928,N_25192);
nand U26673 (N_26673,N_24859,N_25992);
xnor U26674 (N_26674,N_25771,N_24622);
or U26675 (N_26675,N_24593,N_25607);
xor U26676 (N_26676,N_25256,N_24873);
or U26677 (N_26677,N_24248,N_24394);
nor U26678 (N_26678,N_24458,N_25439);
nand U26679 (N_26679,N_25676,N_24923);
and U26680 (N_26680,N_25125,N_24818);
and U26681 (N_26681,N_24960,N_25283);
and U26682 (N_26682,N_24965,N_25407);
xnor U26683 (N_26683,N_25071,N_24181);
nand U26684 (N_26684,N_25242,N_24096);
nand U26685 (N_26685,N_24451,N_24642);
or U26686 (N_26686,N_25931,N_25094);
nand U26687 (N_26687,N_25709,N_24266);
xor U26688 (N_26688,N_25921,N_25200);
or U26689 (N_26689,N_25986,N_25130);
or U26690 (N_26690,N_24439,N_24956);
and U26691 (N_26691,N_24910,N_24862);
nand U26692 (N_26692,N_24636,N_24068);
xnor U26693 (N_26693,N_24662,N_24562);
or U26694 (N_26694,N_24015,N_25032);
nand U26695 (N_26695,N_25004,N_24619);
and U26696 (N_26696,N_24706,N_24417);
nor U26697 (N_26697,N_24885,N_24717);
nor U26698 (N_26698,N_25061,N_24996);
xor U26699 (N_26699,N_25489,N_24078);
and U26700 (N_26700,N_25534,N_25047);
or U26701 (N_26701,N_25451,N_24903);
nand U26702 (N_26702,N_25074,N_24494);
nor U26703 (N_26703,N_25738,N_25015);
or U26704 (N_26704,N_24571,N_24290);
nand U26705 (N_26705,N_25584,N_25395);
nor U26706 (N_26706,N_24942,N_25006);
and U26707 (N_26707,N_24968,N_25772);
nand U26708 (N_26708,N_24513,N_24970);
or U26709 (N_26709,N_25414,N_24716);
or U26710 (N_26710,N_24710,N_24555);
and U26711 (N_26711,N_25821,N_24098);
or U26712 (N_26712,N_25365,N_25838);
or U26713 (N_26713,N_25160,N_24411);
xor U26714 (N_26714,N_25988,N_24255);
or U26715 (N_26715,N_24370,N_24563);
nand U26716 (N_26716,N_24821,N_25895);
nand U26717 (N_26717,N_24519,N_24953);
nor U26718 (N_26718,N_25523,N_25308);
nor U26719 (N_26719,N_24693,N_25127);
nand U26720 (N_26720,N_25732,N_25588);
and U26721 (N_26721,N_24679,N_24756);
or U26722 (N_26722,N_24549,N_24925);
or U26723 (N_26723,N_25958,N_24066);
and U26724 (N_26724,N_24521,N_24908);
and U26725 (N_26725,N_24077,N_25301);
nand U26726 (N_26726,N_25913,N_25905);
nand U26727 (N_26727,N_25358,N_24055);
nor U26728 (N_26728,N_24252,N_25980);
or U26729 (N_26729,N_24140,N_24815);
or U26730 (N_26730,N_24406,N_24373);
or U26731 (N_26731,N_25012,N_25221);
xnor U26732 (N_26732,N_25077,N_24550);
xor U26733 (N_26733,N_25922,N_25273);
nor U26734 (N_26734,N_25398,N_24201);
and U26735 (N_26735,N_24663,N_24009);
or U26736 (N_26736,N_24224,N_24291);
xor U26737 (N_26737,N_25268,N_25528);
nand U26738 (N_26738,N_24128,N_24210);
nand U26739 (N_26739,N_25829,N_24337);
and U26740 (N_26740,N_24025,N_25122);
or U26741 (N_26741,N_25840,N_24631);
or U26742 (N_26742,N_25778,N_24889);
nand U26743 (N_26743,N_24366,N_25976);
xor U26744 (N_26744,N_24300,N_25938);
and U26745 (N_26745,N_24118,N_24396);
xnor U26746 (N_26746,N_25833,N_25320);
nor U26747 (N_26747,N_24329,N_25577);
xnor U26748 (N_26748,N_25472,N_24800);
or U26749 (N_26749,N_24354,N_24233);
or U26750 (N_26750,N_24598,N_25791);
or U26751 (N_26751,N_25220,N_24748);
nand U26752 (N_26752,N_25109,N_24180);
or U26753 (N_26753,N_24543,N_25795);
nand U26754 (N_26754,N_25205,N_24770);
nor U26755 (N_26755,N_24795,N_25479);
xor U26756 (N_26756,N_25216,N_25204);
and U26757 (N_26757,N_25703,N_25121);
and U26758 (N_26758,N_24951,N_25695);
or U26759 (N_26759,N_24866,N_25822);
nand U26760 (N_26760,N_24666,N_24525);
xor U26761 (N_26761,N_24678,N_25238);
nor U26762 (N_26762,N_24313,N_24589);
and U26763 (N_26763,N_24541,N_25296);
or U26764 (N_26764,N_24708,N_24117);
or U26765 (N_26765,N_25841,N_25847);
or U26766 (N_26766,N_24395,N_25449);
and U26767 (N_26767,N_24341,N_24143);
xor U26768 (N_26768,N_25680,N_24176);
xnor U26769 (N_26769,N_24656,N_25725);
or U26770 (N_26770,N_25026,N_24193);
or U26771 (N_26771,N_25504,N_24251);
and U26772 (N_26772,N_24186,N_25385);
and U26773 (N_26773,N_25458,N_24655);
and U26774 (N_26774,N_24604,N_24483);
nand U26775 (N_26775,N_24256,N_24700);
or U26776 (N_26776,N_24119,N_25605);
and U26777 (N_26777,N_24575,N_25357);
nand U26778 (N_26778,N_25037,N_25442);
nand U26779 (N_26779,N_25834,N_24220);
and U26780 (N_26780,N_24265,N_24906);
and U26781 (N_26781,N_24771,N_25696);
or U26782 (N_26782,N_25183,N_25581);
nor U26783 (N_26783,N_24790,N_24792);
nand U26784 (N_26784,N_24142,N_24638);
nand U26785 (N_26785,N_25075,N_25684);
xnor U26786 (N_26786,N_24404,N_25374);
nand U26787 (N_26787,N_24654,N_25763);
and U26788 (N_26788,N_25203,N_25503);
or U26789 (N_26789,N_24172,N_24952);
nor U26790 (N_26790,N_24145,N_24867);
xor U26791 (N_26791,N_24998,N_25535);
xnor U26792 (N_26792,N_25945,N_25497);
nand U26793 (N_26793,N_24920,N_25842);
or U26794 (N_26794,N_24545,N_25352);
nand U26795 (N_26795,N_24985,N_24100);
nor U26796 (N_26796,N_24419,N_24536);
or U26797 (N_26797,N_24240,N_25349);
xor U26798 (N_26798,N_25236,N_24719);
nor U26799 (N_26799,N_24116,N_24368);
xnor U26800 (N_26800,N_24753,N_24798);
and U26801 (N_26801,N_25195,N_24149);
and U26802 (N_26802,N_25682,N_25419);
nor U26803 (N_26803,N_24950,N_25541);
nand U26804 (N_26804,N_24179,N_24069);
and U26805 (N_26805,N_24471,N_25693);
xnor U26806 (N_26806,N_25304,N_24922);
xor U26807 (N_26807,N_25325,N_24386);
xnor U26808 (N_26808,N_24544,N_24060);
nand U26809 (N_26809,N_25661,N_24527);
and U26810 (N_26810,N_24014,N_24720);
xor U26811 (N_26811,N_25425,N_24883);
and U26812 (N_26812,N_25876,N_25752);
or U26813 (N_26813,N_24506,N_24799);
nor U26814 (N_26814,N_24457,N_25550);
nor U26815 (N_26815,N_25133,N_25469);
and U26816 (N_26816,N_24683,N_25142);
xor U26817 (N_26817,N_24788,N_25982);
and U26818 (N_26818,N_25137,N_24932);
and U26819 (N_26819,N_25970,N_25155);
nand U26820 (N_26820,N_24554,N_25854);
nor U26821 (N_26821,N_25874,N_25707);
nand U26822 (N_26822,N_25702,N_25951);
xor U26823 (N_26823,N_25099,N_25933);
nand U26824 (N_26824,N_25467,N_24299);
and U26825 (N_26825,N_24445,N_24365);
nand U26826 (N_26826,N_25762,N_24302);
or U26827 (N_26827,N_24709,N_25520);
nor U26828 (N_26828,N_25843,N_24124);
or U26829 (N_26829,N_25712,N_24132);
and U26830 (N_26830,N_24803,N_24963);
xor U26831 (N_26831,N_25628,N_25161);
nand U26832 (N_26832,N_24135,N_25711);
and U26833 (N_26833,N_24112,N_25724);
nand U26834 (N_26834,N_24495,N_25942);
nor U26835 (N_26835,N_24085,N_24067);
nand U26836 (N_26836,N_25295,N_24739);
xor U26837 (N_26837,N_25606,N_25700);
xnor U26838 (N_26838,N_24566,N_24787);
xor U26839 (N_26839,N_24616,N_24703);
or U26840 (N_26840,N_24292,N_24079);
and U26841 (N_26841,N_25808,N_25827);
and U26842 (N_26842,N_25768,N_24141);
nand U26843 (N_26843,N_25379,N_24348);
and U26844 (N_26844,N_24192,N_24930);
or U26845 (N_26845,N_24381,N_25749);
or U26846 (N_26846,N_24426,N_25685);
or U26847 (N_26847,N_25453,N_25159);
nor U26848 (N_26848,N_24286,N_25644);
xnor U26849 (N_26849,N_24897,N_25332);
nand U26850 (N_26850,N_24110,N_25280);
nand U26851 (N_26851,N_25031,N_25650);
nand U26852 (N_26852,N_24522,N_25902);
or U26853 (N_26853,N_24751,N_24905);
nand U26854 (N_26854,N_25403,N_24600);
nand U26855 (N_26855,N_24891,N_24065);
or U26856 (N_26856,N_25531,N_25310);
nand U26857 (N_26857,N_25612,N_25211);
and U26858 (N_26858,N_24869,N_25227);
xnor U26859 (N_26859,N_24887,N_25386);
xor U26860 (N_26860,N_24465,N_25726);
and U26861 (N_26861,N_25519,N_25857);
or U26862 (N_26862,N_25919,N_24158);
xor U26863 (N_26863,N_25739,N_25070);
nor U26864 (N_26864,N_24958,N_25506);
xor U26865 (N_26865,N_25173,N_25198);
nor U26866 (N_26866,N_24208,N_24505);
and U26867 (N_26867,N_24095,N_25027);
nor U26868 (N_26868,N_24332,N_24633);
xnor U26869 (N_26869,N_24363,N_25105);
nand U26870 (N_26870,N_24308,N_24305);
or U26871 (N_26871,N_25625,N_25741);
nor U26872 (N_26872,N_25993,N_24189);
xnor U26873 (N_26873,N_25809,N_24509);
xnor U26874 (N_26874,N_24323,N_25648);
nand U26875 (N_26875,N_24168,N_24242);
and U26876 (N_26876,N_24307,N_24892);
or U26877 (N_26877,N_25033,N_25966);
and U26878 (N_26878,N_24271,N_25591);
or U26879 (N_26879,N_25573,N_24446);
nand U26880 (N_26880,N_24745,N_25659);
nand U26881 (N_26881,N_24837,N_25867);
and U26882 (N_26882,N_24137,N_25475);
nand U26883 (N_26883,N_24049,N_24169);
xnor U26884 (N_26884,N_24864,N_24485);
nor U26885 (N_26885,N_24225,N_24072);
nor U26886 (N_26886,N_24260,N_24051);
nor U26887 (N_26887,N_25356,N_25996);
nand U26888 (N_26888,N_24507,N_25375);
and U26889 (N_26889,N_24017,N_25422);
or U26890 (N_26890,N_24750,N_24257);
nor U26891 (N_26891,N_25196,N_25824);
nand U26892 (N_26892,N_25566,N_25651);
or U26893 (N_26893,N_24245,N_24059);
xnor U26894 (N_26894,N_25849,N_25586);
or U26895 (N_26895,N_24528,N_25826);
or U26896 (N_26896,N_25482,N_25270);
or U26897 (N_26897,N_24568,N_24385);
nor U26898 (N_26898,N_25642,N_25460);
nand U26899 (N_26899,N_24476,N_25669);
xor U26900 (N_26900,N_25767,N_25345);
or U26901 (N_26901,N_24508,N_25275);
nor U26902 (N_26902,N_25617,N_24045);
xnor U26903 (N_26903,N_25530,N_25640);
nor U26904 (N_26904,N_24781,N_25152);
xnor U26905 (N_26905,N_25312,N_25367);
xor U26906 (N_26906,N_25974,N_25683);
nand U26907 (N_26907,N_25493,N_24939);
and U26908 (N_26908,N_25877,N_25969);
nor U26909 (N_26909,N_24315,N_24175);
and U26910 (N_26910,N_25985,N_25347);
and U26911 (N_26911,N_25719,N_24712);
xnor U26912 (N_26912,N_25690,N_24401);
xnor U26913 (N_26913,N_24828,N_24160);
nor U26914 (N_26914,N_24610,N_25491);
or U26915 (N_26915,N_25570,N_25973);
xnor U26916 (N_26916,N_24435,N_25167);
xor U26917 (N_26917,N_25430,N_25172);
nor U26918 (N_26918,N_25754,N_24194);
nor U26919 (N_26919,N_24244,N_24330);
or U26920 (N_26920,N_25381,N_24202);
or U26921 (N_26921,N_25224,N_25540);
and U26922 (N_26922,N_25934,N_25663);
xnor U26923 (N_26923,N_24845,N_24212);
nand U26924 (N_26924,N_25123,N_25513);
and U26925 (N_26925,N_25022,N_24484);
nor U26926 (N_26926,N_24650,N_24415);
nor U26927 (N_26927,N_25267,N_25393);
or U26928 (N_26928,N_25300,N_24074);
or U26929 (N_26929,N_25705,N_24946);
and U26930 (N_26930,N_24358,N_24711);
nand U26931 (N_26931,N_24472,N_25265);
nor U26932 (N_26932,N_25634,N_25860);
nand U26933 (N_26933,N_25893,N_25073);
and U26934 (N_26934,N_25093,N_25432);
xor U26935 (N_26935,N_25975,N_24336);
xnor U26936 (N_26936,N_25944,N_24637);
xor U26937 (N_26937,N_25851,N_25812);
and U26938 (N_26938,N_25582,N_24576);
or U26939 (N_26939,N_25002,N_25621);
nor U26940 (N_26940,N_24581,N_25201);
nor U26941 (N_26941,N_25646,N_25872);
nor U26942 (N_26942,N_24418,N_25799);
xor U26943 (N_26943,N_25873,N_25326);
xnor U26944 (N_26944,N_25443,N_25608);
or U26945 (N_26945,N_25279,N_24584);
or U26946 (N_26946,N_25668,N_25990);
xor U26947 (N_26947,N_25147,N_24676);
nand U26948 (N_26948,N_25494,N_24360);
and U26949 (N_26949,N_24163,N_25994);
nor U26950 (N_26950,N_24455,N_25346);
nand U26951 (N_26951,N_24723,N_25382);
and U26952 (N_26952,N_24692,N_24048);
and U26953 (N_26953,N_25420,N_25440);
and U26954 (N_26954,N_24881,N_24588);
nand U26955 (N_26955,N_24408,N_25189);
nand U26956 (N_26956,N_24467,N_24540);
and U26957 (N_26957,N_25526,N_25937);
xnor U26958 (N_26958,N_25837,N_24626);
nand U26959 (N_26959,N_24634,N_24615);
or U26960 (N_26960,N_25698,N_24362);
and U26961 (N_26961,N_24013,N_24448);
nor U26962 (N_26962,N_25539,N_25223);
nand U26963 (N_26963,N_25053,N_24272);
nand U26964 (N_26964,N_25594,N_25263);
xor U26965 (N_26965,N_24304,N_24929);
nand U26966 (N_26966,N_25878,N_24834);
and U26967 (N_26967,N_24497,N_25233);
nor U26968 (N_26968,N_24334,N_25701);
nand U26969 (N_26969,N_25116,N_24520);
nor U26970 (N_26970,N_24382,N_24035);
nand U26971 (N_26971,N_24075,N_24301);
xor U26972 (N_26972,N_25947,N_24387);
nor U26973 (N_26973,N_25064,N_24350);
xnor U26974 (N_26974,N_25610,N_25433);
or U26975 (N_26975,N_24402,N_25598);
nor U26976 (N_26976,N_25272,N_24558);
nand U26977 (N_26977,N_24496,N_25085);
and U26978 (N_26978,N_25013,N_25362);
xor U26979 (N_26979,N_25630,N_25747);
xor U26980 (N_26980,N_25140,N_25371);
or U26981 (N_26981,N_24389,N_24504);
and U26982 (N_26982,N_24200,N_24047);
nor U26983 (N_26983,N_24714,N_25353);
and U26984 (N_26984,N_25001,N_24153);
nor U26985 (N_26985,N_25170,N_24995);
nand U26986 (N_26986,N_24056,N_24218);
xor U26987 (N_26987,N_24460,N_25495);
nor U26988 (N_26988,N_25101,N_24630);
nor U26989 (N_26989,N_25409,N_25638);
and U26990 (N_26990,N_25092,N_24731);
nand U26991 (N_26991,N_24822,N_25457);
nor U26992 (N_26992,N_24037,N_24587);
xor U26993 (N_26993,N_25897,N_25464);
and U26994 (N_26994,N_24254,N_25303);
and U26995 (N_26995,N_24962,N_25110);
or U26996 (N_26996,N_25068,N_24136);
nand U26997 (N_26997,N_25802,N_24774);
nand U26998 (N_26998,N_25972,N_25219);
and U26999 (N_26999,N_25730,N_24752);
nor U27000 (N_27000,N_25457,N_25943);
nand U27001 (N_27001,N_25474,N_25593);
xor U27002 (N_27002,N_24697,N_24464);
or U27003 (N_27003,N_24330,N_24239);
or U27004 (N_27004,N_24293,N_24072);
nand U27005 (N_27005,N_25118,N_24325);
nor U27006 (N_27006,N_24247,N_24248);
and U27007 (N_27007,N_25993,N_24482);
xnor U27008 (N_27008,N_25535,N_24698);
nor U27009 (N_27009,N_25190,N_25794);
nand U27010 (N_27010,N_24200,N_24305);
nand U27011 (N_27011,N_25953,N_24274);
or U27012 (N_27012,N_24977,N_25364);
xnor U27013 (N_27013,N_25161,N_24742);
nand U27014 (N_27014,N_25950,N_25869);
nand U27015 (N_27015,N_24358,N_25814);
or U27016 (N_27016,N_24794,N_25345);
nor U27017 (N_27017,N_24268,N_25497);
xnor U27018 (N_27018,N_25735,N_24214);
or U27019 (N_27019,N_24692,N_24331);
nand U27020 (N_27020,N_25557,N_24449);
xor U27021 (N_27021,N_24470,N_24304);
xnor U27022 (N_27022,N_24342,N_25320);
or U27023 (N_27023,N_25105,N_24033);
nor U27024 (N_27024,N_24529,N_24873);
nand U27025 (N_27025,N_25812,N_24125);
or U27026 (N_27026,N_24078,N_25775);
or U27027 (N_27027,N_24708,N_24724);
nor U27028 (N_27028,N_25687,N_25817);
nand U27029 (N_27029,N_25000,N_24979);
and U27030 (N_27030,N_25195,N_25577);
and U27031 (N_27031,N_25487,N_24496);
or U27032 (N_27032,N_25275,N_24305);
xnor U27033 (N_27033,N_24013,N_25840);
xnor U27034 (N_27034,N_24894,N_25529);
xnor U27035 (N_27035,N_25533,N_25006);
and U27036 (N_27036,N_25626,N_25891);
and U27037 (N_27037,N_25365,N_25708);
and U27038 (N_27038,N_25785,N_25935);
nor U27039 (N_27039,N_24848,N_25531);
and U27040 (N_27040,N_25334,N_24148);
and U27041 (N_27041,N_24996,N_24168);
and U27042 (N_27042,N_24182,N_25598);
and U27043 (N_27043,N_24586,N_24196);
nor U27044 (N_27044,N_24255,N_24813);
xor U27045 (N_27045,N_24600,N_24237);
nor U27046 (N_27046,N_24020,N_25867);
xnor U27047 (N_27047,N_25025,N_24006);
nand U27048 (N_27048,N_24676,N_25698);
nand U27049 (N_27049,N_24893,N_24675);
or U27050 (N_27050,N_25344,N_24332);
xnor U27051 (N_27051,N_24896,N_25870);
nand U27052 (N_27052,N_24500,N_25283);
nor U27053 (N_27053,N_24972,N_25047);
and U27054 (N_27054,N_24882,N_24906);
nor U27055 (N_27055,N_25266,N_24728);
nor U27056 (N_27056,N_25293,N_25154);
nor U27057 (N_27057,N_24310,N_24852);
nand U27058 (N_27058,N_24913,N_25671);
nand U27059 (N_27059,N_25737,N_24716);
xor U27060 (N_27060,N_25972,N_24864);
nand U27061 (N_27061,N_25884,N_25719);
nor U27062 (N_27062,N_25651,N_24287);
nand U27063 (N_27063,N_24243,N_24662);
and U27064 (N_27064,N_25083,N_25238);
xor U27065 (N_27065,N_25279,N_25739);
or U27066 (N_27066,N_25397,N_25955);
and U27067 (N_27067,N_24411,N_24691);
xor U27068 (N_27068,N_25622,N_24101);
nand U27069 (N_27069,N_25878,N_24974);
and U27070 (N_27070,N_25001,N_24731);
nor U27071 (N_27071,N_24030,N_24933);
xnor U27072 (N_27072,N_24652,N_24171);
nor U27073 (N_27073,N_25794,N_25206);
or U27074 (N_27074,N_24302,N_24992);
xnor U27075 (N_27075,N_24608,N_25534);
xnor U27076 (N_27076,N_24460,N_24667);
and U27077 (N_27077,N_25134,N_24144);
or U27078 (N_27078,N_25780,N_25459);
xnor U27079 (N_27079,N_25524,N_25924);
xnor U27080 (N_27080,N_25285,N_24191);
nand U27081 (N_27081,N_24442,N_24585);
and U27082 (N_27082,N_25512,N_25847);
xnor U27083 (N_27083,N_25501,N_24005);
xnor U27084 (N_27084,N_25454,N_24816);
or U27085 (N_27085,N_25156,N_25515);
xnor U27086 (N_27086,N_24641,N_25966);
nand U27087 (N_27087,N_25900,N_24325);
nor U27088 (N_27088,N_24008,N_25811);
nand U27089 (N_27089,N_25945,N_25244);
or U27090 (N_27090,N_24297,N_24630);
and U27091 (N_27091,N_24516,N_25554);
nand U27092 (N_27092,N_24575,N_24654);
nand U27093 (N_27093,N_24987,N_24130);
nor U27094 (N_27094,N_24512,N_25224);
nor U27095 (N_27095,N_25805,N_24264);
and U27096 (N_27096,N_24318,N_25984);
and U27097 (N_27097,N_25800,N_24504);
nand U27098 (N_27098,N_25130,N_24394);
xnor U27099 (N_27099,N_25136,N_25332);
nand U27100 (N_27100,N_25720,N_24783);
nor U27101 (N_27101,N_25382,N_25599);
xnor U27102 (N_27102,N_24106,N_25918);
nand U27103 (N_27103,N_25489,N_24786);
xnor U27104 (N_27104,N_24874,N_24751);
or U27105 (N_27105,N_25830,N_24401);
nor U27106 (N_27106,N_25605,N_24953);
and U27107 (N_27107,N_24473,N_25816);
and U27108 (N_27108,N_25983,N_24641);
and U27109 (N_27109,N_25794,N_25977);
nand U27110 (N_27110,N_24943,N_24967);
xnor U27111 (N_27111,N_25536,N_25025);
nand U27112 (N_27112,N_24427,N_24579);
or U27113 (N_27113,N_24248,N_24861);
or U27114 (N_27114,N_25526,N_25476);
nand U27115 (N_27115,N_24345,N_24749);
nand U27116 (N_27116,N_24224,N_24767);
xor U27117 (N_27117,N_24000,N_25663);
or U27118 (N_27118,N_25471,N_24050);
or U27119 (N_27119,N_25333,N_24454);
xnor U27120 (N_27120,N_25521,N_25931);
xor U27121 (N_27121,N_24049,N_25566);
and U27122 (N_27122,N_24837,N_25677);
or U27123 (N_27123,N_24824,N_25559);
or U27124 (N_27124,N_24474,N_24114);
xnor U27125 (N_27125,N_25176,N_25874);
nor U27126 (N_27126,N_24255,N_24202);
nand U27127 (N_27127,N_24404,N_24379);
and U27128 (N_27128,N_25003,N_25226);
nand U27129 (N_27129,N_24037,N_25273);
or U27130 (N_27130,N_25161,N_25298);
and U27131 (N_27131,N_24140,N_24591);
and U27132 (N_27132,N_24877,N_24688);
and U27133 (N_27133,N_25417,N_25427);
nor U27134 (N_27134,N_25038,N_25941);
xnor U27135 (N_27135,N_25679,N_24823);
and U27136 (N_27136,N_25857,N_24427);
nor U27137 (N_27137,N_24817,N_24599);
nor U27138 (N_27138,N_25090,N_24717);
and U27139 (N_27139,N_25718,N_25903);
or U27140 (N_27140,N_24655,N_24301);
and U27141 (N_27141,N_24116,N_24411);
and U27142 (N_27142,N_25136,N_25380);
nand U27143 (N_27143,N_25457,N_25004);
nor U27144 (N_27144,N_25477,N_25693);
nor U27145 (N_27145,N_24583,N_25376);
xnor U27146 (N_27146,N_24519,N_25731);
xnor U27147 (N_27147,N_25738,N_24566);
or U27148 (N_27148,N_24898,N_25607);
xnor U27149 (N_27149,N_24665,N_24295);
and U27150 (N_27150,N_24210,N_24669);
xor U27151 (N_27151,N_24211,N_25208);
and U27152 (N_27152,N_24543,N_24829);
xnor U27153 (N_27153,N_25009,N_25791);
nor U27154 (N_27154,N_24551,N_25088);
xnor U27155 (N_27155,N_24780,N_25281);
nor U27156 (N_27156,N_25317,N_24946);
nand U27157 (N_27157,N_24167,N_25436);
nand U27158 (N_27158,N_25742,N_24948);
nor U27159 (N_27159,N_24377,N_25908);
nor U27160 (N_27160,N_24571,N_25082);
nor U27161 (N_27161,N_24909,N_25012);
xor U27162 (N_27162,N_25624,N_24083);
and U27163 (N_27163,N_25624,N_24514);
nand U27164 (N_27164,N_25328,N_24622);
or U27165 (N_27165,N_25835,N_24838);
nand U27166 (N_27166,N_24401,N_25218);
xnor U27167 (N_27167,N_24256,N_24328);
nand U27168 (N_27168,N_24050,N_24081);
xor U27169 (N_27169,N_24908,N_25943);
xnor U27170 (N_27170,N_25730,N_24009);
xor U27171 (N_27171,N_25927,N_25391);
nand U27172 (N_27172,N_25819,N_24071);
or U27173 (N_27173,N_24326,N_25880);
or U27174 (N_27174,N_25744,N_25087);
nand U27175 (N_27175,N_25713,N_25461);
xor U27176 (N_27176,N_24560,N_24902);
or U27177 (N_27177,N_25521,N_25138);
and U27178 (N_27178,N_25083,N_24527);
xnor U27179 (N_27179,N_24223,N_24485);
and U27180 (N_27180,N_24168,N_25904);
nand U27181 (N_27181,N_24488,N_25749);
nand U27182 (N_27182,N_24641,N_25997);
or U27183 (N_27183,N_24811,N_24538);
or U27184 (N_27184,N_25499,N_25810);
xnor U27185 (N_27185,N_24165,N_24141);
nand U27186 (N_27186,N_25450,N_25614);
nand U27187 (N_27187,N_25818,N_24119);
xnor U27188 (N_27188,N_25420,N_24742);
nand U27189 (N_27189,N_24476,N_24718);
and U27190 (N_27190,N_24045,N_25076);
or U27191 (N_27191,N_25578,N_25309);
nand U27192 (N_27192,N_24212,N_24040);
or U27193 (N_27193,N_25569,N_25167);
and U27194 (N_27194,N_25155,N_25999);
nand U27195 (N_27195,N_25326,N_25819);
and U27196 (N_27196,N_24432,N_24897);
or U27197 (N_27197,N_24884,N_24320);
or U27198 (N_27198,N_25087,N_25822);
or U27199 (N_27199,N_24887,N_25041);
nand U27200 (N_27200,N_24014,N_25390);
nor U27201 (N_27201,N_25748,N_24012);
and U27202 (N_27202,N_25018,N_25858);
and U27203 (N_27203,N_25393,N_24471);
nand U27204 (N_27204,N_25293,N_25369);
and U27205 (N_27205,N_24412,N_24235);
nand U27206 (N_27206,N_24924,N_24875);
nand U27207 (N_27207,N_24542,N_24798);
nor U27208 (N_27208,N_25241,N_25938);
or U27209 (N_27209,N_24881,N_25796);
or U27210 (N_27210,N_24739,N_25178);
nand U27211 (N_27211,N_25698,N_25396);
xnor U27212 (N_27212,N_25623,N_24114);
and U27213 (N_27213,N_25971,N_25441);
nand U27214 (N_27214,N_25500,N_24820);
or U27215 (N_27215,N_25620,N_25788);
nand U27216 (N_27216,N_24631,N_24873);
or U27217 (N_27217,N_24457,N_25976);
and U27218 (N_27218,N_25954,N_24538);
or U27219 (N_27219,N_24862,N_24784);
nor U27220 (N_27220,N_24480,N_25789);
and U27221 (N_27221,N_25306,N_24836);
and U27222 (N_27222,N_24702,N_25512);
or U27223 (N_27223,N_24868,N_24784);
or U27224 (N_27224,N_25426,N_25926);
nor U27225 (N_27225,N_24924,N_25329);
or U27226 (N_27226,N_24197,N_25202);
xor U27227 (N_27227,N_25525,N_24671);
nand U27228 (N_27228,N_25475,N_24397);
nor U27229 (N_27229,N_25893,N_25795);
nand U27230 (N_27230,N_25314,N_25687);
nor U27231 (N_27231,N_24419,N_24601);
and U27232 (N_27232,N_25646,N_25888);
and U27233 (N_27233,N_25227,N_24072);
or U27234 (N_27234,N_24438,N_24633);
and U27235 (N_27235,N_25816,N_25445);
or U27236 (N_27236,N_24931,N_25963);
nor U27237 (N_27237,N_25960,N_25348);
nor U27238 (N_27238,N_25592,N_24593);
xnor U27239 (N_27239,N_24083,N_24702);
xor U27240 (N_27240,N_25988,N_25207);
xnor U27241 (N_27241,N_25231,N_24112);
and U27242 (N_27242,N_24946,N_24751);
nand U27243 (N_27243,N_25230,N_24257);
nand U27244 (N_27244,N_24813,N_25301);
or U27245 (N_27245,N_24056,N_24879);
nand U27246 (N_27246,N_24244,N_24548);
nand U27247 (N_27247,N_24268,N_25439);
and U27248 (N_27248,N_25556,N_24994);
xor U27249 (N_27249,N_25321,N_25065);
or U27250 (N_27250,N_25547,N_25409);
or U27251 (N_27251,N_25503,N_25815);
or U27252 (N_27252,N_24206,N_24864);
nor U27253 (N_27253,N_25036,N_24991);
and U27254 (N_27254,N_25368,N_25401);
nand U27255 (N_27255,N_24333,N_24779);
and U27256 (N_27256,N_25820,N_24954);
xor U27257 (N_27257,N_24725,N_24489);
and U27258 (N_27258,N_24737,N_25127);
nand U27259 (N_27259,N_25004,N_24351);
nor U27260 (N_27260,N_24737,N_25433);
or U27261 (N_27261,N_24818,N_25696);
and U27262 (N_27262,N_24372,N_25482);
or U27263 (N_27263,N_25385,N_24542);
or U27264 (N_27264,N_24328,N_24443);
nor U27265 (N_27265,N_25852,N_25595);
nor U27266 (N_27266,N_25931,N_24909);
nand U27267 (N_27267,N_25059,N_25854);
and U27268 (N_27268,N_24888,N_24785);
nand U27269 (N_27269,N_24545,N_25961);
nand U27270 (N_27270,N_24623,N_24508);
nor U27271 (N_27271,N_25692,N_25133);
or U27272 (N_27272,N_25072,N_24118);
nor U27273 (N_27273,N_24234,N_24324);
nor U27274 (N_27274,N_24591,N_25452);
nand U27275 (N_27275,N_25806,N_25842);
nor U27276 (N_27276,N_24124,N_24851);
or U27277 (N_27277,N_25952,N_25497);
xor U27278 (N_27278,N_25559,N_24656);
or U27279 (N_27279,N_25030,N_24425);
xnor U27280 (N_27280,N_24399,N_25473);
nor U27281 (N_27281,N_25207,N_24464);
xor U27282 (N_27282,N_25616,N_24480);
xnor U27283 (N_27283,N_25118,N_24869);
nand U27284 (N_27284,N_24790,N_24225);
xor U27285 (N_27285,N_25312,N_25065);
or U27286 (N_27286,N_25649,N_24236);
and U27287 (N_27287,N_24724,N_24878);
nand U27288 (N_27288,N_24764,N_25915);
nor U27289 (N_27289,N_24411,N_24266);
and U27290 (N_27290,N_25204,N_25628);
or U27291 (N_27291,N_24156,N_25186);
and U27292 (N_27292,N_24543,N_25351);
or U27293 (N_27293,N_24831,N_25769);
nor U27294 (N_27294,N_24334,N_24726);
nand U27295 (N_27295,N_25835,N_24021);
nor U27296 (N_27296,N_24449,N_24321);
or U27297 (N_27297,N_25660,N_25729);
nand U27298 (N_27298,N_25320,N_25506);
nand U27299 (N_27299,N_25394,N_25598);
and U27300 (N_27300,N_25372,N_25976);
and U27301 (N_27301,N_25562,N_25109);
and U27302 (N_27302,N_24027,N_24214);
and U27303 (N_27303,N_25510,N_25741);
nand U27304 (N_27304,N_24444,N_24672);
nand U27305 (N_27305,N_24739,N_24525);
nand U27306 (N_27306,N_25475,N_24271);
nor U27307 (N_27307,N_24020,N_24943);
nor U27308 (N_27308,N_25742,N_24347);
xor U27309 (N_27309,N_25040,N_25293);
nor U27310 (N_27310,N_25066,N_25374);
and U27311 (N_27311,N_25082,N_24348);
or U27312 (N_27312,N_24780,N_25866);
nand U27313 (N_27313,N_25631,N_24249);
nand U27314 (N_27314,N_24318,N_24252);
or U27315 (N_27315,N_24870,N_24141);
xnor U27316 (N_27316,N_25253,N_25129);
xnor U27317 (N_27317,N_24782,N_25547);
and U27318 (N_27318,N_24622,N_25749);
and U27319 (N_27319,N_24308,N_24336);
and U27320 (N_27320,N_24987,N_24651);
nand U27321 (N_27321,N_24111,N_24477);
nor U27322 (N_27322,N_25330,N_25255);
nand U27323 (N_27323,N_25204,N_24217);
and U27324 (N_27324,N_25346,N_24293);
and U27325 (N_27325,N_25634,N_24087);
and U27326 (N_27326,N_24690,N_24847);
or U27327 (N_27327,N_25761,N_24480);
nand U27328 (N_27328,N_25159,N_25436);
or U27329 (N_27329,N_25151,N_25348);
nor U27330 (N_27330,N_24015,N_25812);
or U27331 (N_27331,N_24298,N_24106);
or U27332 (N_27332,N_25866,N_24977);
or U27333 (N_27333,N_25938,N_24891);
nor U27334 (N_27334,N_25633,N_25781);
or U27335 (N_27335,N_25318,N_25910);
xor U27336 (N_27336,N_24317,N_25617);
nor U27337 (N_27337,N_25397,N_24933);
nor U27338 (N_27338,N_24006,N_25293);
and U27339 (N_27339,N_24529,N_24848);
and U27340 (N_27340,N_24778,N_25353);
and U27341 (N_27341,N_25039,N_24057);
and U27342 (N_27342,N_24131,N_25556);
and U27343 (N_27343,N_24816,N_25401);
and U27344 (N_27344,N_25555,N_25863);
nand U27345 (N_27345,N_25201,N_24913);
nand U27346 (N_27346,N_25875,N_25200);
or U27347 (N_27347,N_25866,N_25567);
nor U27348 (N_27348,N_24731,N_24440);
nand U27349 (N_27349,N_25053,N_25152);
xnor U27350 (N_27350,N_25341,N_24490);
or U27351 (N_27351,N_24936,N_24151);
nand U27352 (N_27352,N_24960,N_24010);
and U27353 (N_27353,N_24387,N_25496);
nand U27354 (N_27354,N_25324,N_25414);
xor U27355 (N_27355,N_24017,N_25727);
nor U27356 (N_27356,N_25140,N_24814);
nand U27357 (N_27357,N_25075,N_25795);
or U27358 (N_27358,N_24866,N_24120);
xnor U27359 (N_27359,N_24846,N_25552);
and U27360 (N_27360,N_25554,N_25487);
nand U27361 (N_27361,N_25516,N_24981);
and U27362 (N_27362,N_25694,N_25667);
or U27363 (N_27363,N_24078,N_25182);
nor U27364 (N_27364,N_24913,N_25958);
and U27365 (N_27365,N_25986,N_24089);
xnor U27366 (N_27366,N_25095,N_25202);
or U27367 (N_27367,N_25446,N_24631);
nor U27368 (N_27368,N_24541,N_25248);
xnor U27369 (N_27369,N_25985,N_24505);
xor U27370 (N_27370,N_24617,N_25209);
xnor U27371 (N_27371,N_25144,N_24305);
nand U27372 (N_27372,N_25903,N_25139);
or U27373 (N_27373,N_25593,N_24513);
or U27374 (N_27374,N_24670,N_25261);
and U27375 (N_27375,N_25620,N_24428);
xor U27376 (N_27376,N_25173,N_24541);
nor U27377 (N_27377,N_25307,N_25541);
nand U27378 (N_27378,N_24786,N_24752);
xnor U27379 (N_27379,N_25069,N_24680);
and U27380 (N_27380,N_24498,N_25624);
and U27381 (N_27381,N_25205,N_24325);
and U27382 (N_27382,N_25238,N_25579);
nor U27383 (N_27383,N_24095,N_24137);
nor U27384 (N_27384,N_24403,N_24997);
nor U27385 (N_27385,N_24657,N_24631);
and U27386 (N_27386,N_25659,N_24527);
xor U27387 (N_27387,N_24696,N_24154);
and U27388 (N_27388,N_24497,N_24538);
or U27389 (N_27389,N_25139,N_25472);
nor U27390 (N_27390,N_25383,N_25958);
and U27391 (N_27391,N_24751,N_24329);
or U27392 (N_27392,N_25026,N_25630);
or U27393 (N_27393,N_24755,N_24511);
or U27394 (N_27394,N_25808,N_25668);
or U27395 (N_27395,N_24650,N_24617);
and U27396 (N_27396,N_25000,N_24316);
or U27397 (N_27397,N_25767,N_25738);
nor U27398 (N_27398,N_25739,N_25838);
and U27399 (N_27399,N_24162,N_24196);
nor U27400 (N_27400,N_24121,N_25302);
xnor U27401 (N_27401,N_25519,N_24717);
nor U27402 (N_27402,N_25872,N_24114);
or U27403 (N_27403,N_25396,N_24856);
xnor U27404 (N_27404,N_24503,N_24904);
nand U27405 (N_27405,N_24154,N_24273);
or U27406 (N_27406,N_24823,N_24639);
or U27407 (N_27407,N_25109,N_25983);
nor U27408 (N_27408,N_25413,N_24927);
xnor U27409 (N_27409,N_25911,N_24058);
xor U27410 (N_27410,N_24806,N_25789);
xnor U27411 (N_27411,N_24006,N_24655);
nand U27412 (N_27412,N_25120,N_24475);
or U27413 (N_27413,N_24358,N_25542);
or U27414 (N_27414,N_24929,N_25877);
nor U27415 (N_27415,N_25996,N_25478);
nand U27416 (N_27416,N_25600,N_25030);
xnor U27417 (N_27417,N_25100,N_24292);
xnor U27418 (N_27418,N_25993,N_24067);
nor U27419 (N_27419,N_25586,N_25109);
or U27420 (N_27420,N_24174,N_24029);
nand U27421 (N_27421,N_25079,N_25879);
nand U27422 (N_27422,N_25354,N_25711);
nand U27423 (N_27423,N_24096,N_25125);
or U27424 (N_27424,N_24462,N_25256);
nor U27425 (N_27425,N_25221,N_25549);
and U27426 (N_27426,N_24651,N_24869);
nor U27427 (N_27427,N_25913,N_25737);
and U27428 (N_27428,N_25055,N_24775);
nand U27429 (N_27429,N_25716,N_25704);
nand U27430 (N_27430,N_25814,N_25498);
and U27431 (N_27431,N_25520,N_25000);
xor U27432 (N_27432,N_25829,N_25911);
xor U27433 (N_27433,N_25306,N_25447);
and U27434 (N_27434,N_24892,N_25839);
nor U27435 (N_27435,N_24639,N_24981);
nor U27436 (N_27436,N_24420,N_25249);
nand U27437 (N_27437,N_24134,N_24146);
nor U27438 (N_27438,N_25359,N_25610);
xnor U27439 (N_27439,N_24432,N_25892);
or U27440 (N_27440,N_25187,N_24758);
nand U27441 (N_27441,N_25832,N_25226);
nand U27442 (N_27442,N_24377,N_25430);
xnor U27443 (N_27443,N_24618,N_24644);
nor U27444 (N_27444,N_25851,N_25706);
or U27445 (N_27445,N_24957,N_24383);
nor U27446 (N_27446,N_25646,N_25315);
xor U27447 (N_27447,N_25677,N_25836);
xnor U27448 (N_27448,N_24011,N_25410);
nand U27449 (N_27449,N_25457,N_25506);
nand U27450 (N_27450,N_24130,N_24192);
and U27451 (N_27451,N_24654,N_24093);
nand U27452 (N_27452,N_24841,N_24200);
and U27453 (N_27453,N_24171,N_24697);
xnor U27454 (N_27454,N_25140,N_25154);
xor U27455 (N_27455,N_24247,N_24434);
or U27456 (N_27456,N_24722,N_25605);
nand U27457 (N_27457,N_25169,N_25799);
nor U27458 (N_27458,N_25789,N_25038);
xor U27459 (N_27459,N_24645,N_25039);
xnor U27460 (N_27460,N_24212,N_25303);
and U27461 (N_27461,N_25167,N_25745);
or U27462 (N_27462,N_25677,N_24540);
xnor U27463 (N_27463,N_25536,N_25475);
or U27464 (N_27464,N_25247,N_25806);
nand U27465 (N_27465,N_24351,N_24646);
nand U27466 (N_27466,N_24233,N_25314);
nor U27467 (N_27467,N_25904,N_24652);
and U27468 (N_27468,N_25851,N_24306);
and U27469 (N_27469,N_24376,N_24491);
xor U27470 (N_27470,N_25518,N_24612);
nand U27471 (N_27471,N_25153,N_24422);
xor U27472 (N_27472,N_25177,N_24906);
xor U27473 (N_27473,N_25785,N_24233);
nor U27474 (N_27474,N_25465,N_24314);
and U27475 (N_27475,N_24690,N_24662);
or U27476 (N_27476,N_25638,N_25574);
xor U27477 (N_27477,N_24219,N_25045);
nand U27478 (N_27478,N_24659,N_24580);
nand U27479 (N_27479,N_24761,N_24673);
and U27480 (N_27480,N_25934,N_25844);
nor U27481 (N_27481,N_24267,N_25141);
and U27482 (N_27482,N_24912,N_25453);
and U27483 (N_27483,N_24992,N_24938);
xor U27484 (N_27484,N_24658,N_25881);
or U27485 (N_27485,N_25313,N_25400);
nand U27486 (N_27486,N_24141,N_25453);
and U27487 (N_27487,N_25078,N_25679);
or U27488 (N_27488,N_24647,N_24262);
nor U27489 (N_27489,N_25516,N_25453);
and U27490 (N_27490,N_25228,N_24821);
xor U27491 (N_27491,N_24595,N_25632);
nand U27492 (N_27492,N_25442,N_24203);
and U27493 (N_27493,N_24258,N_25345);
nor U27494 (N_27494,N_25020,N_24178);
and U27495 (N_27495,N_25899,N_24883);
nand U27496 (N_27496,N_24995,N_24650);
nand U27497 (N_27497,N_24347,N_25224);
and U27498 (N_27498,N_25240,N_24054);
and U27499 (N_27499,N_24516,N_25918);
nor U27500 (N_27500,N_25418,N_25737);
nand U27501 (N_27501,N_24085,N_24771);
and U27502 (N_27502,N_24563,N_25964);
or U27503 (N_27503,N_25299,N_24559);
or U27504 (N_27504,N_25122,N_24752);
nand U27505 (N_27505,N_25937,N_25649);
nor U27506 (N_27506,N_24065,N_25583);
xnor U27507 (N_27507,N_24945,N_24808);
nor U27508 (N_27508,N_25390,N_24774);
nand U27509 (N_27509,N_24432,N_24831);
nor U27510 (N_27510,N_24556,N_25333);
nor U27511 (N_27511,N_24390,N_24807);
xnor U27512 (N_27512,N_25261,N_24352);
nor U27513 (N_27513,N_25438,N_24446);
and U27514 (N_27514,N_25907,N_24297);
nor U27515 (N_27515,N_24795,N_24006);
and U27516 (N_27516,N_25402,N_25215);
and U27517 (N_27517,N_25953,N_25472);
nor U27518 (N_27518,N_24379,N_24988);
nor U27519 (N_27519,N_25376,N_24546);
xnor U27520 (N_27520,N_25389,N_24671);
xnor U27521 (N_27521,N_24654,N_25660);
nor U27522 (N_27522,N_25485,N_25636);
and U27523 (N_27523,N_25682,N_25667);
nand U27524 (N_27524,N_25187,N_24335);
nand U27525 (N_27525,N_25674,N_25392);
nand U27526 (N_27526,N_25132,N_25224);
xnor U27527 (N_27527,N_24616,N_24987);
nand U27528 (N_27528,N_24975,N_25980);
and U27529 (N_27529,N_25867,N_25468);
nand U27530 (N_27530,N_25541,N_25972);
or U27531 (N_27531,N_24407,N_24219);
xnor U27532 (N_27532,N_25190,N_25829);
nand U27533 (N_27533,N_25632,N_24086);
xor U27534 (N_27534,N_25030,N_25245);
xor U27535 (N_27535,N_24027,N_24598);
and U27536 (N_27536,N_24781,N_25466);
nor U27537 (N_27537,N_24629,N_24135);
nor U27538 (N_27538,N_24430,N_24302);
and U27539 (N_27539,N_24744,N_24679);
or U27540 (N_27540,N_24379,N_25575);
nand U27541 (N_27541,N_25647,N_25058);
or U27542 (N_27542,N_25154,N_24822);
nand U27543 (N_27543,N_25243,N_24555);
nand U27544 (N_27544,N_25268,N_25460);
xnor U27545 (N_27545,N_24233,N_25180);
or U27546 (N_27546,N_24318,N_25318);
and U27547 (N_27547,N_24219,N_25260);
nand U27548 (N_27548,N_24295,N_25449);
nor U27549 (N_27549,N_25379,N_24635);
xnor U27550 (N_27550,N_25288,N_25088);
nor U27551 (N_27551,N_24004,N_24355);
and U27552 (N_27552,N_24164,N_24231);
nand U27553 (N_27553,N_25976,N_25571);
nor U27554 (N_27554,N_24696,N_24187);
and U27555 (N_27555,N_25738,N_25543);
or U27556 (N_27556,N_24448,N_24963);
and U27557 (N_27557,N_24007,N_24584);
nor U27558 (N_27558,N_24883,N_25994);
and U27559 (N_27559,N_25378,N_24223);
nor U27560 (N_27560,N_24813,N_24987);
xor U27561 (N_27561,N_25122,N_24107);
or U27562 (N_27562,N_25845,N_25092);
or U27563 (N_27563,N_24363,N_25844);
xnor U27564 (N_27564,N_24018,N_24445);
nand U27565 (N_27565,N_24358,N_24188);
nand U27566 (N_27566,N_25305,N_24818);
nor U27567 (N_27567,N_24874,N_24547);
or U27568 (N_27568,N_25884,N_24067);
xnor U27569 (N_27569,N_25077,N_24334);
nor U27570 (N_27570,N_25382,N_25924);
xor U27571 (N_27571,N_25709,N_25571);
nor U27572 (N_27572,N_24773,N_24229);
nor U27573 (N_27573,N_24930,N_24000);
xnor U27574 (N_27574,N_25548,N_25783);
or U27575 (N_27575,N_24580,N_24923);
and U27576 (N_27576,N_24118,N_25896);
xnor U27577 (N_27577,N_24090,N_25216);
or U27578 (N_27578,N_25006,N_25174);
xor U27579 (N_27579,N_24224,N_25013);
or U27580 (N_27580,N_24895,N_24386);
or U27581 (N_27581,N_25023,N_24497);
nand U27582 (N_27582,N_24185,N_24553);
nor U27583 (N_27583,N_24245,N_25581);
and U27584 (N_27584,N_25475,N_24284);
nor U27585 (N_27585,N_25817,N_25165);
nor U27586 (N_27586,N_24402,N_24262);
or U27587 (N_27587,N_25032,N_24238);
nor U27588 (N_27588,N_25808,N_24432);
nor U27589 (N_27589,N_24136,N_24383);
nor U27590 (N_27590,N_24447,N_24897);
or U27591 (N_27591,N_24936,N_25124);
or U27592 (N_27592,N_24192,N_24554);
and U27593 (N_27593,N_24180,N_24416);
nor U27594 (N_27594,N_25366,N_25242);
and U27595 (N_27595,N_24017,N_24738);
nor U27596 (N_27596,N_25351,N_25217);
or U27597 (N_27597,N_24948,N_25950);
nand U27598 (N_27598,N_25791,N_24776);
or U27599 (N_27599,N_24911,N_24928);
xnor U27600 (N_27600,N_25682,N_24405);
nand U27601 (N_27601,N_24039,N_24838);
nor U27602 (N_27602,N_24139,N_24400);
nor U27603 (N_27603,N_25540,N_25684);
nand U27604 (N_27604,N_24386,N_25691);
nor U27605 (N_27605,N_25776,N_25495);
nand U27606 (N_27606,N_25891,N_24421);
nand U27607 (N_27607,N_24561,N_24965);
nand U27608 (N_27608,N_25642,N_25790);
nor U27609 (N_27609,N_25690,N_24409);
and U27610 (N_27610,N_24959,N_25999);
nor U27611 (N_27611,N_24807,N_25082);
xor U27612 (N_27612,N_24486,N_24855);
nand U27613 (N_27613,N_25827,N_24275);
nor U27614 (N_27614,N_24986,N_25044);
or U27615 (N_27615,N_25203,N_25345);
or U27616 (N_27616,N_25504,N_25334);
and U27617 (N_27617,N_24715,N_24588);
or U27618 (N_27618,N_24523,N_25523);
and U27619 (N_27619,N_25051,N_25083);
nand U27620 (N_27620,N_24229,N_25681);
or U27621 (N_27621,N_25505,N_25451);
and U27622 (N_27622,N_24740,N_24168);
and U27623 (N_27623,N_24095,N_24706);
nand U27624 (N_27624,N_24649,N_25855);
and U27625 (N_27625,N_24183,N_24954);
nand U27626 (N_27626,N_24296,N_24980);
and U27627 (N_27627,N_25568,N_25516);
or U27628 (N_27628,N_25263,N_24445);
and U27629 (N_27629,N_25479,N_24598);
and U27630 (N_27630,N_24914,N_25893);
xor U27631 (N_27631,N_25848,N_25678);
nand U27632 (N_27632,N_24863,N_24746);
nand U27633 (N_27633,N_25655,N_25291);
xnor U27634 (N_27634,N_25676,N_24296);
nor U27635 (N_27635,N_25664,N_24465);
nand U27636 (N_27636,N_25438,N_24929);
xor U27637 (N_27637,N_24532,N_24861);
xnor U27638 (N_27638,N_25458,N_25005);
nand U27639 (N_27639,N_24216,N_25086);
or U27640 (N_27640,N_25778,N_25578);
and U27641 (N_27641,N_24285,N_25083);
nand U27642 (N_27642,N_24174,N_24479);
and U27643 (N_27643,N_24217,N_25904);
nor U27644 (N_27644,N_24175,N_24789);
xor U27645 (N_27645,N_25127,N_25699);
or U27646 (N_27646,N_25339,N_25286);
xnor U27647 (N_27647,N_25316,N_24453);
and U27648 (N_27648,N_25036,N_25774);
and U27649 (N_27649,N_25475,N_24482);
xnor U27650 (N_27650,N_25471,N_25690);
xnor U27651 (N_27651,N_24420,N_24712);
or U27652 (N_27652,N_24208,N_25709);
nand U27653 (N_27653,N_25858,N_24365);
nor U27654 (N_27654,N_25794,N_25975);
nand U27655 (N_27655,N_24865,N_24779);
and U27656 (N_27656,N_24745,N_24788);
or U27657 (N_27657,N_25948,N_25467);
xor U27658 (N_27658,N_25440,N_24524);
nor U27659 (N_27659,N_25990,N_24784);
and U27660 (N_27660,N_25720,N_24815);
and U27661 (N_27661,N_24155,N_24055);
or U27662 (N_27662,N_24180,N_25256);
nor U27663 (N_27663,N_24639,N_25328);
or U27664 (N_27664,N_25411,N_24776);
xnor U27665 (N_27665,N_25192,N_25097);
xnor U27666 (N_27666,N_24206,N_24475);
and U27667 (N_27667,N_24836,N_25874);
nor U27668 (N_27668,N_24404,N_25560);
nand U27669 (N_27669,N_24122,N_25163);
nor U27670 (N_27670,N_25307,N_25947);
xnor U27671 (N_27671,N_25952,N_25897);
or U27672 (N_27672,N_24979,N_24781);
and U27673 (N_27673,N_24608,N_25118);
and U27674 (N_27674,N_24963,N_25454);
and U27675 (N_27675,N_25622,N_24371);
or U27676 (N_27676,N_24120,N_24357);
nand U27677 (N_27677,N_25807,N_25837);
and U27678 (N_27678,N_24101,N_24237);
xor U27679 (N_27679,N_24265,N_25830);
and U27680 (N_27680,N_24200,N_25114);
xor U27681 (N_27681,N_24081,N_25533);
nor U27682 (N_27682,N_25290,N_25610);
xor U27683 (N_27683,N_25744,N_25192);
nor U27684 (N_27684,N_25424,N_25818);
nor U27685 (N_27685,N_25794,N_25987);
xor U27686 (N_27686,N_24259,N_24351);
or U27687 (N_27687,N_24149,N_25170);
nor U27688 (N_27688,N_25609,N_25026);
nand U27689 (N_27689,N_25900,N_25127);
and U27690 (N_27690,N_25947,N_25968);
nand U27691 (N_27691,N_25799,N_25522);
and U27692 (N_27692,N_25241,N_24060);
and U27693 (N_27693,N_24160,N_25216);
nand U27694 (N_27694,N_25249,N_24067);
or U27695 (N_27695,N_24984,N_25867);
or U27696 (N_27696,N_25979,N_24905);
and U27697 (N_27697,N_25883,N_25650);
nand U27698 (N_27698,N_24701,N_25300);
nor U27699 (N_27699,N_24915,N_24598);
or U27700 (N_27700,N_25945,N_25784);
nand U27701 (N_27701,N_24269,N_25927);
nand U27702 (N_27702,N_25992,N_25599);
and U27703 (N_27703,N_25270,N_25864);
nor U27704 (N_27704,N_25462,N_24463);
nand U27705 (N_27705,N_25331,N_24362);
nor U27706 (N_27706,N_25285,N_24248);
nor U27707 (N_27707,N_25941,N_24109);
nor U27708 (N_27708,N_24447,N_24540);
xor U27709 (N_27709,N_25631,N_24923);
nand U27710 (N_27710,N_25210,N_24958);
nand U27711 (N_27711,N_25942,N_25978);
nand U27712 (N_27712,N_25749,N_24093);
or U27713 (N_27713,N_25089,N_24731);
or U27714 (N_27714,N_24312,N_25645);
or U27715 (N_27715,N_25994,N_24849);
and U27716 (N_27716,N_24397,N_24912);
nand U27717 (N_27717,N_25689,N_25917);
and U27718 (N_27718,N_25310,N_24828);
xor U27719 (N_27719,N_25427,N_25750);
nor U27720 (N_27720,N_24343,N_25393);
nor U27721 (N_27721,N_25565,N_24771);
and U27722 (N_27722,N_24374,N_25472);
nor U27723 (N_27723,N_25460,N_25331);
nor U27724 (N_27724,N_24065,N_25845);
nand U27725 (N_27725,N_25174,N_24120);
or U27726 (N_27726,N_24365,N_24701);
and U27727 (N_27727,N_24615,N_25219);
or U27728 (N_27728,N_24988,N_25616);
or U27729 (N_27729,N_24251,N_25020);
nor U27730 (N_27730,N_24591,N_24560);
or U27731 (N_27731,N_25882,N_25534);
and U27732 (N_27732,N_24285,N_24173);
xnor U27733 (N_27733,N_25786,N_24561);
and U27734 (N_27734,N_24241,N_25518);
nor U27735 (N_27735,N_24868,N_25454);
xnor U27736 (N_27736,N_24044,N_25319);
xnor U27737 (N_27737,N_24124,N_25851);
nor U27738 (N_27738,N_24705,N_25401);
and U27739 (N_27739,N_24893,N_24339);
or U27740 (N_27740,N_24667,N_24346);
or U27741 (N_27741,N_25643,N_24688);
xnor U27742 (N_27742,N_24216,N_25851);
and U27743 (N_27743,N_25903,N_24679);
or U27744 (N_27744,N_24926,N_24458);
nand U27745 (N_27745,N_24850,N_25835);
or U27746 (N_27746,N_25842,N_24918);
and U27747 (N_27747,N_25787,N_24353);
and U27748 (N_27748,N_25962,N_25315);
and U27749 (N_27749,N_24459,N_24773);
and U27750 (N_27750,N_25539,N_25534);
nand U27751 (N_27751,N_24718,N_25443);
or U27752 (N_27752,N_24801,N_24959);
or U27753 (N_27753,N_24598,N_24551);
or U27754 (N_27754,N_25533,N_25794);
or U27755 (N_27755,N_25725,N_25901);
nor U27756 (N_27756,N_25758,N_25751);
nand U27757 (N_27757,N_24409,N_25659);
and U27758 (N_27758,N_24861,N_25838);
and U27759 (N_27759,N_25297,N_24975);
xor U27760 (N_27760,N_25164,N_24824);
nand U27761 (N_27761,N_24967,N_24639);
or U27762 (N_27762,N_24697,N_24306);
nor U27763 (N_27763,N_25956,N_24577);
and U27764 (N_27764,N_24125,N_25515);
xor U27765 (N_27765,N_25812,N_24856);
or U27766 (N_27766,N_25779,N_24821);
xnor U27767 (N_27767,N_24757,N_24898);
xor U27768 (N_27768,N_24671,N_25094);
nor U27769 (N_27769,N_24631,N_25211);
or U27770 (N_27770,N_25363,N_24158);
xor U27771 (N_27771,N_25534,N_24253);
or U27772 (N_27772,N_25487,N_25893);
and U27773 (N_27773,N_24263,N_24180);
and U27774 (N_27774,N_25729,N_25314);
nor U27775 (N_27775,N_24130,N_25949);
nor U27776 (N_27776,N_25474,N_25945);
nor U27777 (N_27777,N_24027,N_25034);
or U27778 (N_27778,N_24777,N_24719);
xor U27779 (N_27779,N_25957,N_24991);
and U27780 (N_27780,N_24041,N_24369);
nor U27781 (N_27781,N_24807,N_24726);
xnor U27782 (N_27782,N_24561,N_24349);
nand U27783 (N_27783,N_25467,N_24909);
nor U27784 (N_27784,N_25520,N_25122);
nand U27785 (N_27785,N_24064,N_24694);
or U27786 (N_27786,N_24822,N_24205);
xor U27787 (N_27787,N_25579,N_24968);
or U27788 (N_27788,N_24054,N_24438);
nand U27789 (N_27789,N_24310,N_25761);
or U27790 (N_27790,N_24534,N_24903);
xnor U27791 (N_27791,N_24903,N_24986);
nor U27792 (N_27792,N_24017,N_25574);
nand U27793 (N_27793,N_24834,N_24238);
nor U27794 (N_27794,N_24543,N_24206);
or U27795 (N_27795,N_24562,N_25861);
and U27796 (N_27796,N_24757,N_25914);
xor U27797 (N_27797,N_25755,N_24354);
and U27798 (N_27798,N_25218,N_25969);
xnor U27799 (N_27799,N_24792,N_25237);
and U27800 (N_27800,N_25755,N_25999);
xor U27801 (N_27801,N_25038,N_24112);
and U27802 (N_27802,N_25444,N_24387);
nand U27803 (N_27803,N_24048,N_25276);
xor U27804 (N_27804,N_25724,N_24261);
or U27805 (N_27805,N_24388,N_25167);
nand U27806 (N_27806,N_24823,N_24615);
or U27807 (N_27807,N_25273,N_25665);
and U27808 (N_27808,N_25475,N_25156);
and U27809 (N_27809,N_25781,N_24674);
and U27810 (N_27810,N_25965,N_24047);
xor U27811 (N_27811,N_25258,N_24807);
or U27812 (N_27812,N_24928,N_25027);
and U27813 (N_27813,N_25895,N_25038);
and U27814 (N_27814,N_25812,N_24281);
nor U27815 (N_27815,N_25005,N_25887);
nor U27816 (N_27816,N_25114,N_25899);
and U27817 (N_27817,N_25736,N_25656);
nand U27818 (N_27818,N_24184,N_24890);
nand U27819 (N_27819,N_24146,N_25034);
xnor U27820 (N_27820,N_24503,N_25604);
or U27821 (N_27821,N_24738,N_25586);
or U27822 (N_27822,N_24780,N_25814);
and U27823 (N_27823,N_24887,N_25190);
and U27824 (N_27824,N_25026,N_25511);
nand U27825 (N_27825,N_25650,N_25994);
or U27826 (N_27826,N_25402,N_25153);
and U27827 (N_27827,N_25029,N_24495);
xor U27828 (N_27828,N_25373,N_24343);
nand U27829 (N_27829,N_24089,N_24397);
xnor U27830 (N_27830,N_25965,N_24702);
and U27831 (N_27831,N_24013,N_24037);
nor U27832 (N_27832,N_24940,N_25492);
nand U27833 (N_27833,N_24010,N_24859);
or U27834 (N_27834,N_25642,N_24301);
or U27835 (N_27835,N_24143,N_25877);
xnor U27836 (N_27836,N_25730,N_25904);
nor U27837 (N_27837,N_25844,N_24194);
or U27838 (N_27838,N_24102,N_25318);
and U27839 (N_27839,N_24215,N_24514);
xor U27840 (N_27840,N_24180,N_25047);
or U27841 (N_27841,N_25334,N_24411);
nand U27842 (N_27842,N_24199,N_24341);
xor U27843 (N_27843,N_25278,N_25727);
or U27844 (N_27844,N_24181,N_25506);
nor U27845 (N_27845,N_25045,N_25508);
and U27846 (N_27846,N_24110,N_24571);
or U27847 (N_27847,N_24899,N_24149);
nor U27848 (N_27848,N_25001,N_25202);
nor U27849 (N_27849,N_24309,N_25352);
xnor U27850 (N_27850,N_24373,N_24510);
nand U27851 (N_27851,N_25219,N_25169);
xor U27852 (N_27852,N_25207,N_24450);
nor U27853 (N_27853,N_24232,N_24222);
or U27854 (N_27854,N_24815,N_24073);
nor U27855 (N_27855,N_25532,N_25759);
nand U27856 (N_27856,N_25375,N_25576);
and U27857 (N_27857,N_25235,N_24866);
or U27858 (N_27858,N_25126,N_25884);
nand U27859 (N_27859,N_24433,N_25898);
xnor U27860 (N_27860,N_24958,N_25228);
xor U27861 (N_27861,N_25720,N_24638);
and U27862 (N_27862,N_25482,N_25069);
nor U27863 (N_27863,N_24245,N_25341);
xnor U27864 (N_27864,N_24203,N_24633);
xnor U27865 (N_27865,N_25412,N_24052);
and U27866 (N_27866,N_24651,N_25113);
or U27867 (N_27867,N_25684,N_25870);
or U27868 (N_27868,N_24041,N_24037);
xnor U27869 (N_27869,N_25946,N_25506);
xnor U27870 (N_27870,N_25708,N_24438);
nor U27871 (N_27871,N_25534,N_24949);
xnor U27872 (N_27872,N_25284,N_24108);
nand U27873 (N_27873,N_24254,N_24734);
nand U27874 (N_27874,N_25996,N_25677);
nand U27875 (N_27875,N_25080,N_25931);
or U27876 (N_27876,N_25344,N_24854);
xor U27877 (N_27877,N_25871,N_25001);
or U27878 (N_27878,N_24914,N_25050);
nand U27879 (N_27879,N_25135,N_24743);
or U27880 (N_27880,N_25135,N_25583);
xnor U27881 (N_27881,N_25183,N_25829);
or U27882 (N_27882,N_25706,N_25513);
nor U27883 (N_27883,N_24813,N_24536);
or U27884 (N_27884,N_24051,N_24176);
nand U27885 (N_27885,N_24251,N_24227);
nand U27886 (N_27886,N_25135,N_24582);
or U27887 (N_27887,N_25934,N_24997);
nor U27888 (N_27888,N_25359,N_24634);
nor U27889 (N_27889,N_25471,N_24560);
and U27890 (N_27890,N_25659,N_24403);
nor U27891 (N_27891,N_25757,N_24115);
and U27892 (N_27892,N_24453,N_25923);
xor U27893 (N_27893,N_25719,N_24472);
or U27894 (N_27894,N_24366,N_24024);
and U27895 (N_27895,N_24590,N_25154);
xnor U27896 (N_27896,N_25665,N_25272);
nor U27897 (N_27897,N_24461,N_25416);
or U27898 (N_27898,N_25409,N_25986);
xor U27899 (N_27899,N_25413,N_25214);
xnor U27900 (N_27900,N_25051,N_25541);
nor U27901 (N_27901,N_24196,N_24961);
or U27902 (N_27902,N_25094,N_24435);
nor U27903 (N_27903,N_25489,N_24306);
and U27904 (N_27904,N_25464,N_25049);
nor U27905 (N_27905,N_25059,N_24992);
and U27906 (N_27906,N_24434,N_25607);
or U27907 (N_27907,N_24643,N_25984);
or U27908 (N_27908,N_24542,N_24035);
or U27909 (N_27909,N_24454,N_25051);
xnor U27910 (N_27910,N_24945,N_25269);
nor U27911 (N_27911,N_24811,N_24019);
xor U27912 (N_27912,N_25492,N_25859);
and U27913 (N_27913,N_24560,N_25265);
xor U27914 (N_27914,N_24431,N_24017);
nand U27915 (N_27915,N_24513,N_24517);
or U27916 (N_27916,N_25913,N_25357);
nor U27917 (N_27917,N_25227,N_25932);
nor U27918 (N_27918,N_25811,N_24104);
nand U27919 (N_27919,N_25154,N_25767);
and U27920 (N_27920,N_25624,N_24930);
xor U27921 (N_27921,N_25595,N_25848);
or U27922 (N_27922,N_24870,N_24659);
nor U27923 (N_27923,N_24516,N_24926);
or U27924 (N_27924,N_24163,N_24818);
nand U27925 (N_27925,N_24718,N_24567);
and U27926 (N_27926,N_24506,N_25234);
xnor U27927 (N_27927,N_24502,N_25657);
and U27928 (N_27928,N_24225,N_25174);
xnor U27929 (N_27929,N_25401,N_24549);
and U27930 (N_27930,N_25271,N_24499);
or U27931 (N_27931,N_25165,N_25334);
nand U27932 (N_27932,N_25013,N_24947);
nand U27933 (N_27933,N_25124,N_24834);
nor U27934 (N_27934,N_24923,N_25931);
nand U27935 (N_27935,N_25315,N_24628);
xor U27936 (N_27936,N_25520,N_25830);
nand U27937 (N_27937,N_24518,N_24467);
xor U27938 (N_27938,N_25160,N_24900);
nor U27939 (N_27939,N_25725,N_24134);
xor U27940 (N_27940,N_25292,N_24928);
xnor U27941 (N_27941,N_24088,N_25004);
xor U27942 (N_27942,N_25151,N_24040);
nand U27943 (N_27943,N_25927,N_25787);
nor U27944 (N_27944,N_24396,N_25095);
xor U27945 (N_27945,N_24415,N_24336);
nand U27946 (N_27946,N_25991,N_25138);
or U27947 (N_27947,N_25856,N_25505);
xnor U27948 (N_27948,N_24870,N_25960);
xor U27949 (N_27949,N_24097,N_24723);
nor U27950 (N_27950,N_25011,N_24091);
nand U27951 (N_27951,N_25550,N_25728);
xor U27952 (N_27952,N_24043,N_25440);
nor U27953 (N_27953,N_24423,N_24923);
nor U27954 (N_27954,N_24452,N_25191);
and U27955 (N_27955,N_24642,N_24793);
or U27956 (N_27956,N_24063,N_25219);
xor U27957 (N_27957,N_24043,N_25944);
nor U27958 (N_27958,N_25249,N_24300);
nand U27959 (N_27959,N_24147,N_24723);
or U27960 (N_27960,N_24279,N_24297);
or U27961 (N_27961,N_25499,N_24768);
or U27962 (N_27962,N_24739,N_25335);
or U27963 (N_27963,N_25573,N_25638);
and U27964 (N_27964,N_24906,N_24386);
nand U27965 (N_27965,N_24332,N_24934);
nor U27966 (N_27966,N_24151,N_24648);
or U27967 (N_27967,N_25913,N_25295);
nand U27968 (N_27968,N_25774,N_24566);
nor U27969 (N_27969,N_25115,N_24050);
xor U27970 (N_27970,N_24065,N_24594);
nand U27971 (N_27971,N_25581,N_25256);
nor U27972 (N_27972,N_24817,N_24627);
nor U27973 (N_27973,N_24348,N_24058);
and U27974 (N_27974,N_25035,N_25731);
nand U27975 (N_27975,N_25366,N_24099);
and U27976 (N_27976,N_24494,N_25261);
and U27977 (N_27977,N_24612,N_25966);
and U27978 (N_27978,N_25605,N_24958);
nand U27979 (N_27979,N_25456,N_24454);
nor U27980 (N_27980,N_25726,N_24113);
nand U27981 (N_27981,N_25976,N_24229);
xor U27982 (N_27982,N_25072,N_24424);
nor U27983 (N_27983,N_25468,N_24279);
nand U27984 (N_27984,N_25915,N_24404);
or U27985 (N_27985,N_24410,N_24243);
and U27986 (N_27986,N_24869,N_25041);
xnor U27987 (N_27987,N_24709,N_24111);
nand U27988 (N_27988,N_24671,N_24280);
nor U27989 (N_27989,N_25382,N_24321);
and U27990 (N_27990,N_24375,N_24147);
nand U27991 (N_27991,N_24378,N_24822);
and U27992 (N_27992,N_25333,N_24951);
nand U27993 (N_27993,N_24447,N_25745);
nor U27994 (N_27994,N_24565,N_24492);
and U27995 (N_27995,N_24845,N_24720);
xnor U27996 (N_27996,N_24127,N_24826);
or U27997 (N_27997,N_24301,N_25224);
and U27998 (N_27998,N_25011,N_24816);
nand U27999 (N_27999,N_25836,N_25980);
nor U28000 (N_28000,N_27490,N_26861);
and U28001 (N_28001,N_26702,N_27952);
and U28002 (N_28002,N_26153,N_26262);
and U28003 (N_28003,N_27603,N_27056);
nand U28004 (N_28004,N_26150,N_26091);
or U28005 (N_28005,N_27895,N_27742);
xnor U28006 (N_28006,N_26652,N_27737);
xnor U28007 (N_28007,N_26825,N_26604);
nor U28008 (N_28008,N_26980,N_26761);
and U28009 (N_28009,N_26574,N_27563);
xor U28010 (N_28010,N_27449,N_27276);
and U28011 (N_28011,N_27736,N_26845);
nor U28012 (N_28012,N_26499,N_27834);
and U28013 (N_28013,N_26847,N_27567);
and U28014 (N_28014,N_26465,N_26720);
nor U28015 (N_28015,N_26594,N_27639);
or U28016 (N_28016,N_27781,N_26459);
xnor U28017 (N_28017,N_27769,N_27804);
or U28018 (N_28018,N_27533,N_27986);
xor U28019 (N_28019,N_27861,N_26225);
nand U28020 (N_28020,N_26068,N_27296);
nand U28021 (N_28021,N_26265,N_27032);
nand U28022 (N_28022,N_26421,N_27470);
or U28023 (N_28023,N_26795,N_27034);
and U28024 (N_28024,N_27434,N_27645);
and U28025 (N_28025,N_26273,N_26081);
or U28026 (N_28026,N_26045,N_26970);
nor U28027 (N_28027,N_27063,N_27049);
and U28028 (N_28028,N_26076,N_27831);
nor U28029 (N_28029,N_26609,N_26138);
and U28030 (N_28030,N_27238,N_26201);
nand U28031 (N_28031,N_26496,N_26532);
nand U28032 (N_28032,N_26900,N_27973);
nor U28033 (N_28033,N_27007,N_27474);
nor U28034 (N_28034,N_27347,N_26555);
xor U28035 (N_28035,N_27424,N_26165);
nor U28036 (N_28036,N_26264,N_27403);
and U28037 (N_28037,N_27260,N_27544);
xnor U28038 (N_28038,N_26056,N_27762);
xnor U28039 (N_28039,N_26893,N_26377);
xnor U28040 (N_28040,N_27362,N_27303);
xor U28041 (N_28041,N_27892,N_27636);
xor U28042 (N_28042,N_26228,N_27024);
nor U28043 (N_28043,N_26101,N_26983);
xor U28044 (N_28044,N_26616,N_27270);
and U28045 (N_28045,N_26935,N_26100);
xor U28046 (N_28046,N_26724,N_27251);
and U28047 (N_28047,N_27874,N_26177);
nor U28048 (N_28048,N_27110,N_27231);
nand U28049 (N_28049,N_27499,N_27314);
or U28050 (N_28050,N_27728,N_27538);
nor U28051 (N_28051,N_26742,N_26820);
or U28052 (N_28052,N_27376,N_27658);
nor U28053 (N_28053,N_26433,N_26011);
or U28054 (N_28054,N_26271,N_27686);
or U28055 (N_28055,N_26454,N_27946);
and U28056 (N_28056,N_27132,N_27333);
xnor U28057 (N_28057,N_26467,N_26188);
nor U28058 (N_28058,N_26318,N_26187);
xor U28059 (N_28059,N_26053,N_27543);
nor U28060 (N_28060,N_27635,N_26489);
nor U28061 (N_28061,N_26600,N_26480);
nand U28062 (N_28062,N_26729,N_26233);
nor U28063 (N_28063,N_26839,N_27890);
xor U28064 (N_28064,N_26482,N_27562);
nor U28065 (N_28065,N_26412,N_27398);
xnor U28066 (N_28066,N_27185,N_27248);
and U28067 (N_28067,N_26577,N_27366);
or U28068 (N_28068,N_26199,N_26017);
or U28069 (N_28069,N_26185,N_26442);
or U28070 (N_28070,N_27628,N_26818);
and U28071 (N_28071,N_26718,N_27922);
xnor U28072 (N_28072,N_27328,N_27319);
or U28073 (N_28073,N_26778,N_27877);
or U28074 (N_28074,N_27534,N_27082);
or U28075 (N_28075,N_27367,N_27167);
and U28076 (N_28076,N_27528,N_26103);
nor U28077 (N_28077,N_27593,N_27439);
or U28078 (N_28078,N_27662,N_26733);
or U28079 (N_28079,N_27318,N_27375);
and U28080 (N_28080,N_27018,N_27710);
and U28081 (N_28081,N_26198,N_26668);
and U28082 (N_28082,N_27400,N_26242);
nor U28083 (N_28083,N_27712,N_27705);
nand U28084 (N_28084,N_26735,N_26678);
and U28085 (N_28085,N_26799,N_27327);
xnor U28086 (N_28086,N_26368,N_27391);
xnor U28087 (N_28087,N_26708,N_27655);
xnor U28088 (N_28088,N_26736,N_27405);
nor U28089 (N_28089,N_26021,N_27661);
nand U28090 (N_28090,N_26329,N_26645);
and U28091 (N_28091,N_26524,N_26420);
nand U28092 (N_28092,N_26682,N_26958);
and U28093 (N_28093,N_27496,N_26022);
nand U28094 (N_28094,N_27141,N_27146);
and U28095 (N_28095,N_27990,N_26737);
and U28096 (N_28096,N_27076,N_26964);
nor U28097 (N_28097,N_26926,N_26922);
nand U28098 (N_28098,N_27878,N_27432);
nand U28099 (N_28099,N_27396,N_26322);
nor U28100 (N_28100,N_27027,N_27390);
nor U28101 (N_28101,N_27226,N_27440);
xor U28102 (N_28102,N_26597,N_26491);
nor U28103 (N_28103,N_27153,N_27531);
xnor U28104 (N_28104,N_26186,N_26064);
or U28105 (N_28105,N_26218,N_26722);
xor U28106 (N_28106,N_26250,N_26413);
xor U28107 (N_28107,N_27682,N_26918);
xnor U28108 (N_28108,N_26407,N_27818);
xor U28109 (N_28109,N_26178,N_27476);
nand U28110 (N_28110,N_27605,N_26208);
and U28111 (N_28111,N_26042,N_26525);
and U28112 (N_28112,N_27600,N_27659);
nand U28113 (N_28113,N_26593,N_26510);
and U28114 (N_28114,N_27237,N_27058);
and U28115 (N_28115,N_26142,N_26074);
xnor U28116 (N_28116,N_27749,N_27981);
xnor U28117 (N_28117,N_27526,N_26578);
nor U28118 (N_28118,N_27671,N_26509);
nand U28119 (N_28119,N_27194,N_26418);
nor U28120 (N_28120,N_26770,N_27217);
and U28121 (N_28121,N_26495,N_27339);
nand U28122 (N_28122,N_27124,N_27075);
or U28123 (N_28123,N_27441,N_27274);
xor U28124 (N_28124,N_27042,N_27967);
nand U28125 (N_28125,N_27936,N_26615);
nand U28126 (N_28126,N_26195,N_26275);
and U28127 (N_28127,N_27989,N_26498);
or U28128 (N_28128,N_27553,N_26289);
xor U28129 (N_28129,N_26288,N_27987);
or U28130 (N_28130,N_27322,N_27999);
nor U28131 (N_28131,N_26429,N_27930);
xnor U28132 (N_28132,N_26695,N_26161);
xnor U28133 (N_28133,N_27340,N_27283);
nand U28134 (N_28134,N_27370,N_27527);
and U28135 (N_28135,N_27115,N_27910);
or U28136 (N_28136,N_26487,N_27865);
xnor U28137 (N_28137,N_27601,N_27297);
nand U28138 (N_28138,N_26332,N_26805);
xor U28139 (N_28139,N_26147,N_27059);
nand U28140 (N_28140,N_27423,N_27951);
nor U28141 (N_28141,N_27569,N_26966);
nand U28142 (N_28142,N_27093,N_27640);
xnor U28143 (N_28143,N_26406,N_26436);
nor U28144 (N_28144,N_26346,N_26950);
and U28145 (N_28145,N_26758,N_26596);
nand U28146 (N_28146,N_26430,N_26865);
xor U28147 (N_28147,N_27155,N_26437);
or U28148 (N_28148,N_26375,N_27037);
xor U28149 (N_28149,N_26913,N_27135);
nor U28150 (N_28150,N_27383,N_27443);
and U28151 (N_28151,N_26019,N_26330);
nor U28152 (N_28152,N_26933,N_27036);
nor U28153 (N_28153,N_26641,N_27939);
or U28154 (N_28154,N_27506,N_27113);
or U28155 (N_28155,N_27897,N_26369);
xnor U28156 (N_28156,N_27255,N_26908);
xor U28157 (N_28157,N_26323,N_26107);
nor U28158 (N_28158,N_26921,N_27698);
or U28159 (N_28159,N_26383,N_26236);
xor U28160 (N_28160,N_26241,N_26889);
nand U28161 (N_28161,N_27358,N_27458);
xor U28162 (N_28162,N_26697,N_26904);
nand U28163 (N_28163,N_27931,N_27656);
xor U28164 (N_28164,N_26326,N_27856);
xor U28165 (N_28165,N_27753,N_26752);
and U28166 (N_28166,N_26083,N_27554);
xnor U28167 (N_28167,N_27004,N_26295);
and U28168 (N_28168,N_27595,N_26376);
nand U28169 (N_28169,N_27843,N_27087);
nor U28170 (N_28170,N_27450,N_27938);
or U28171 (N_28171,N_27719,N_26850);
or U28172 (N_28172,N_26519,N_27262);
xor U28173 (N_28173,N_27883,N_26576);
or U28174 (N_28174,N_26305,N_26469);
and U28175 (N_28175,N_27416,N_27315);
xnor U28176 (N_28176,N_26148,N_27074);
or U28177 (N_28177,N_27859,N_26898);
xnor U28178 (N_28178,N_27565,N_26713);
and U28179 (N_28179,N_26409,N_27077);
nand U28180 (N_28180,N_27670,N_26094);
nor U28181 (N_28181,N_26226,N_26679);
and U28182 (N_28182,N_26540,N_26569);
or U28183 (N_28183,N_26686,N_26144);
or U28184 (N_28184,N_27239,N_26553);
xor U28185 (N_28185,N_27828,N_27876);
and U28186 (N_28186,N_27045,N_27240);
and U28187 (N_28187,N_27862,N_27001);
nor U28188 (N_28188,N_26050,N_27797);
xor U28189 (N_28189,N_26963,N_26456);
nor U28190 (N_28190,N_26961,N_26916);
and U28191 (N_28191,N_27023,N_27166);
nand U28192 (N_28192,N_27970,N_26052);
or U28193 (N_28193,N_27385,N_26631);
nand U28194 (N_28194,N_27128,N_26692);
xnor U28195 (N_28195,N_26215,N_26222);
xor U28196 (N_28196,N_26610,N_27386);
xnor U28197 (N_28197,N_27792,N_27751);
or U28198 (N_28198,N_26629,N_26009);
nor U28199 (N_28199,N_27665,N_27446);
nor U28200 (N_28200,N_26967,N_26632);
and U28201 (N_28201,N_27889,N_27807);
or U28202 (N_28202,N_26872,N_27627);
xnor U28203 (N_28203,N_27566,N_27505);
nand U28204 (N_28204,N_26292,N_27879);
and U28205 (N_28205,N_27105,N_26563);
or U28206 (N_28206,N_26106,N_27752);
or U28207 (N_28207,N_26344,N_26357);
nor U28208 (N_28208,N_27794,N_26183);
nor U28209 (N_28209,N_26987,N_26527);
xor U28210 (N_28210,N_27062,N_26651);
or U28211 (N_28211,N_27522,N_27718);
or U28212 (N_28212,N_27447,N_26352);
nand U28213 (N_28213,N_26356,N_26526);
xnor U28214 (N_28214,N_27184,N_26962);
nand U28215 (N_28215,N_26905,N_26755);
nor U28216 (N_28216,N_26164,N_27057);
or U28217 (N_28217,N_26623,N_26535);
nor U28218 (N_28218,N_26685,N_26723);
or U28219 (N_28219,N_26092,N_27244);
xor U28220 (N_28220,N_26879,N_27891);
and U28221 (N_28221,N_27477,N_26603);
xnor U28222 (N_28222,N_27944,N_26197);
or U28223 (N_28223,N_27279,N_26727);
nor U28224 (N_28224,N_27149,N_27516);
and U28225 (N_28225,N_27469,N_27329);
xor U28226 (N_28226,N_27326,N_26883);
nor U28227 (N_28227,N_27438,N_27332);
xor U28228 (N_28228,N_26015,N_26644);
xnor U28229 (N_28229,N_27501,N_26672);
nand U28230 (N_28230,N_26231,N_27421);
or U28231 (N_28231,N_26364,N_27817);
and U28232 (N_28232,N_27455,N_26281);
xnor U28233 (N_28233,N_27572,N_27955);
nor U28234 (N_28234,N_27551,N_27069);
xnor U28235 (N_28235,N_26080,N_27352);
nand U28236 (N_28236,N_27133,N_27019);
nand U28237 (N_28237,N_26690,N_27485);
xnor U28238 (N_28238,N_26874,N_26530);
and U28239 (N_28239,N_27965,N_27863);
and U28240 (N_28240,N_27183,N_27145);
xnor U28241 (N_28241,N_27591,N_27577);
xor U28242 (N_28242,N_26707,N_27431);
nand U28243 (N_28243,N_27815,N_26367);
nand U28244 (N_28244,N_26804,N_27875);
and U28245 (N_28245,N_27679,N_27151);
xnor U28246 (N_28246,N_26309,N_27508);
nor U28247 (N_28247,N_27882,N_27745);
or U28248 (N_28248,N_27824,N_26440);
and U28249 (N_28249,N_26590,N_27047);
nand U28250 (N_28250,N_26841,N_26739);
or U28251 (N_28251,N_26556,N_26614);
nand U28252 (N_28252,N_27630,N_27893);
and U28253 (N_28253,N_26314,N_26296);
or U28254 (N_28254,N_26771,N_26808);
nand U28255 (N_28255,N_26827,N_27540);
nor U28256 (N_28256,N_26130,N_27191);
nand U28257 (N_28257,N_27933,N_26057);
nor U28258 (N_28258,N_27827,N_26166);
nor U28259 (N_28259,N_26086,N_27678);
or U28260 (N_28260,N_27871,N_26002);
nand U28261 (N_28261,N_27273,N_27812);
or U28262 (N_28262,N_27437,N_27313);
nand U28263 (N_28263,N_27805,N_27811);
and U28264 (N_28264,N_27560,N_27223);
or U28265 (N_28265,N_26276,N_26580);
and U28266 (N_28266,N_26719,N_26573);
nor U28267 (N_28267,N_26528,N_27960);
nor U28268 (N_28268,N_27568,N_27703);
nor U28269 (N_28269,N_27173,N_26207);
or U28270 (N_28270,N_26971,N_26586);
nor U28271 (N_28271,N_26479,N_27980);
nor U28272 (N_28272,N_26493,N_26168);
xor U28273 (N_28273,N_27012,N_27320);
nand U28274 (N_28274,N_26716,N_26073);
xnor U28275 (N_28275,N_27453,N_26776);
nor U28276 (N_28276,N_27494,N_27697);
or U28277 (N_28277,N_27870,N_27098);
xnor U28278 (N_28278,N_26474,N_27305);
and U28279 (N_28279,N_26097,N_27624);
or U28280 (N_28280,N_26069,N_26558);
or U28281 (N_28281,N_27121,N_27150);
and U28282 (N_28282,N_27198,N_26223);
nor U28283 (N_28283,N_26455,N_27278);
nor U28284 (N_28284,N_27025,N_27844);
and U28285 (N_28285,N_27186,N_26400);
xnor U28286 (N_28286,N_26452,N_26826);
and U28287 (N_28287,N_26485,N_26372);
nand U28288 (N_28288,N_26507,N_27579);
nor U28289 (N_28289,N_26310,N_26422);
nor U28290 (N_28290,N_27407,N_26029);
xnor U28291 (N_28291,N_27061,N_27504);
and U28292 (N_28292,N_26554,N_26129);
and U28293 (N_28293,N_27621,N_26763);
and U28294 (N_28294,N_27466,N_26030);
nand U28295 (N_28295,N_26561,N_27215);
nand U28296 (N_28296,N_27454,N_27741);
nand U28297 (N_28297,N_27495,N_26853);
xnor U28298 (N_28298,N_27071,N_26880);
or U28299 (N_28299,N_26035,N_26529);
nor U28300 (N_28300,N_26858,N_27747);
xor U28301 (N_28301,N_26712,N_27581);
and U28302 (N_28302,N_26599,N_26306);
and U28303 (N_28303,N_26522,N_27716);
nand U28304 (N_28304,N_26389,N_26054);
or U28305 (N_28305,N_27123,N_26122);
nand U28306 (N_28306,N_27654,N_27195);
nor U28307 (N_28307,N_26544,N_26854);
and U28308 (N_28308,N_26915,N_26940);
or U28309 (N_28309,N_27968,N_26829);
nor U28310 (N_28310,N_26157,N_27761);
nor U28311 (N_28311,N_26796,N_26709);
or U28312 (N_28312,N_26088,N_26234);
and U28313 (N_28313,N_27626,N_26779);
or U28314 (N_28314,N_26315,N_26192);
and U28315 (N_28315,N_26244,N_26067);
nand U28316 (N_28316,N_26848,N_26335);
or U28317 (N_28317,N_27104,N_27550);
nor U28318 (N_28318,N_26331,N_26481);
and U28319 (N_28319,N_26120,N_26837);
or U28320 (N_28320,N_27271,N_27675);
or U28321 (N_28321,N_27356,N_27346);
and U28322 (N_28322,N_26396,N_26028);
or U28323 (N_28323,N_27881,N_26304);
and U28324 (N_28324,N_27157,N_27561);
nor U28325 (N_28325,N_27463,N_26782);
nor U28326 (N_28326,N_27974,N_26446);
nor U28327 (N_28327,N_27800,N_26089);
xor U28328 (N_28328,N_27913,N_26235);
or U28329 (N_28329,N_27687,N_27221);
xnor U28330 (N_28330,N_27825,N_27849);
nor U28331 (N_28331,N_27963,N_27997);
nor U28332 (N_28332,N_26928,N_26868);
nor U28333 (N_28333,N_27552,N_27564);
or U28334 (N_28334,N_27291,N_27847);
nor U28335 (N_28335,N_27402,N_27998);
and U28336 (N_28336,N_26885,N_26575);
and U28337 (N_28337,N_27982,N_27729);
xnor U28338 (N_28338,N_27174,N_26392);
xor U28339 (N_28339,N_27756,N_27514);
or U28340 (N_28340,N_27109,N_27634);
and U28341 (N_28341,N_26159,N_26070);
or U28342 (N_28342,N_26875,N_26194);
nand U28343 (N_28343,N_27160,N_27425);
nand U28344 (N_28344,N_26923,N_26741);
nand U28345 (N_28345,N_26930,N_27695);
nor U28346 (N_28346,N_27768,N_26098);
or U28347 (N_28347,N_26753,N_27821);
and U28348 (N_28348,N_27452,N_26238);
or U28349 (N_28349,N_26533,N_26726);
xnor U28350 (N_28350,N_26082,N_26515);
xor U28351 (N_28351,N_27858,N_26173);
or U28352 (N_28352,N_26831,N_26071);
nand U28353 (N_28353,N_26806,N_26212);
nand U28354 (N_28354,N_26216,N_27456);
nand U28355 (N_28355,N_26172,N_27011);
nor U28356 (N_28356,N_27298,N_27757);
or U28357 (N_28357,N_27092,N_26370);
nor U28358 (N_28358,N_27465,N_26892);
nand U28359 (N_28359,N_26204,N_27114);
or U28360 (N_28360,N_26232,N_27597);
nand U28361 (N_28361,N_27677,N_27584);
nand U28362 (N_28362,N_26432,N_27547);
xnor U28363 (N_28363,N_26055,N_27395);
or U28364 (N_28364,N_26041,N_27854);
and U28365 (N_28365,N_26982,N_27604);
and U28366 (N_28366,N_26840,N_26815);
and U28367 (N_28367,N_27585,N_27266);
xnor U28368 (N_28368,N_26912,N_26957);
or U28369 (N_28369,N_27609,N_27835);
nand U28370 (N_28370,N_27227,N_26773);
xor U28371 (N_28371,N_27498,N_26450);
nand U28372 (N_28372,N_26005,N_26994);
or U28373 (N_28373,N_26860,N_27152);
or U28374 (N_28374,N_26634,N_27943);
nor U28375 (N_28375,N_27257,N_27672);
nand U28376 (N_28376,N_27957,N_26894);
xor U28377 (N_28377,N_27706,N_27975);
and U28378 (N_28378,N_27249,N_26427);
or U28379 (N_28379,N_26568,N_27393);
nor U28380 (N_28380,N_27387,N_27357);
or U28381 (N_28381,N_27802,N_26792);
and U28382 (N_28382,N_26360,N_26431);
xnor U28383 (N_28383,N_27330,N_26391);
or U28384 (N_28384,N_27941,N_26660);
xnor U28385 (N_28385,N_26873,N_27801);
and U28386 (N_28386,N_27210,N_26824);
nor U28387 (N_28387,N_27349,N_26072);
xnor U28388 (N_28388,N_27342,N_26635);
or U28389 (N_28389,N_26924,N_26085);
xor U28390 (N_28390,N_26995,N_26666);
and U28391 (N_28391,N_26877,N_26985);
xnor U28392 (N_28392,N_26349,N_26620);
nand U28393 (N_28393,N_26605,N_26034);
xnor U28394 (N_28394,N_26313,N_26749);
and U28395 (N_28395,N_26388,N_26468);
xor U28396 (N_28396,N_26584,N_26033);
and U28397 (N_28397,N_26477,N_26043);
xnor U28398 (N_28398,N_27462,N_26294);
or U28399 (N_28399,N_27773,N_27623);
nand U28400 (N_28400,N_27611,N_26539);
nor U28401 (N_28401,N_27708,N_26287);
and U28402 (N_28402,N_27073,N_26516);
xnor U28403 (N_28403,N_26855,N_27268);
nor U28404 (N_28404,N_27335,N_27614);
or U28405 (N_28405,N_27277,N_27345);
nand U28406 (N_28406,N_26259,N_27162);
nand U28407 (N_28407,N_26990,N_27343);
or U28408 (N_28408,N_27334,N_27945);
xor U28409 (N_28409,N_27715,N_26221);
nor U28410 (N_28410,N_27643,N_27212);
xor U28411 (N_28411,N_26975,N_26401);
or U28412 (N_28412,N_26137,N_27803);
and U28413 (N_28413,N_27410,N_26333);
or U28414 (N_28414,N_27833,N_26366);
xor U28415 (N_28415,N_26453,N_27222);
xnor U28416 (N_28416,N_26500,N_26787);
and U28417 (N_28417,N_27810,N_26320);
nor U28418 (N_28418,N_27513,N_26624);
nand U28419 (N_28419,N_27288,N_26136);
nand U28420 (N_28420,N_27048,N_27206);
xnor U28421 (N_28421,N_27254,N_26750);
and U28422 (N_28422,N_27189,N_27164);
nand U28423 (N_28423,N_27304,N_27190);
or U28424 (N_28424,N_26711,N_26564);
and U28425 (N_28425,N_27932,N_26710);
nor U28426 (N_28426,N_27264,N_27744);
nor U28427 (N_28427,N_26821,N_26270);
or U28428 (N_28428,N_26260,N_27445);
xnor U28429 (N_28429,N_26999,N_27156);
nand U28430 (N_28430,N_26000,N_27193);
nor U28431 (N_28431,N_27929,N_26152);
nor U28432 (N_28432,N_27765,N_27170);
or U28433 (N_28433,N_27521,N_26058);
nand U28434 (N_28434,N_27208,N_27594);
xor U28435 (N_28435,N_27923,N_27520);
nand U28436 (N_28436,N_26549,N_27241);
or U28437 (N_28437,N_26051,N_27289);
or U28438 (N_28438,N_27586,N_26390);
nor U28439 (N_28439,N_27066,N_26663);
and U28440 (N_28440,N_27364,N_26715);
or U28441 (N_28441,N_27723,N_26308);
and U28442 (N_28442,N_27397,N_27269);
or U28443 (N_28443,N_26284,N_27935);
nand U28444 (N_28444,N_27355,N_26492);
nor U28445 (N_28445,N_26449,N_27489);
and U28446 (N_28446,N_27163,N_27147);
or U28447 (N_28447,N_26888,N_27583);
nor U28448 (N_28448,N_27122,N_26649);
xnor U28449 (N_28449,N_26105,N_26944);
or U28450 (N_28450,N_26943,N_27250);
nand U28451 (N_28451,N_26302,N_26256);
or U28452 (N_28452,N_26743,N_27641);
xor U28453 (N_28453,N_26647,N_27430);
nor U28454 (N_28454,N_27515,N_26764);
xnor U28455 (N_28455,N_26095,N_26112);
and U28456 (N_28456,N_26502,N_27046);
nand U28457 (N_28457,N_26077,N_27444);
nor U28458 (N_28458,N_27545,N_26595);
and U28459 (N_28459,N_26380,N_26508);
or U28460 (N_28460,N_27484,N_26126);
nand U28461 (N_28461,N_26744,N_26007);
nor U28462 (N_28462,N_26038,N_26478);
nor U28463 (N_28463,N_26588,N_27556);
or U28464 (N_28464,N_26747,N_26140);
xnor U28465 (N_28465,N_26611,N_27947);
and U28466 (N_28466,N_27888,N_26993);
nand U28467 (N_28467,N_26026,N_26298);
nor U28468 (N_28468,N_27168,N_27331);
or U28469 (N_28469,N_26061,N_26020);
xnor U28470 (N_28470,N_26984,N_27293);
nor U28471 (N_28471,N_26633,N_26503);
nor U28472 (N_28472,N_26988,N_26781);
nand U28473 (N_28473,N_27908,N_26394);
and U28474 (N_28474,N_26910,N_26180);
nand U28475 (N_28475,N_26760,N_26683);
nor U28476 (N_28476,N_27738,N_27775);
nand U28477 (N_28477,N_27549,N_26630);
or U28478 (N_28478,N_27693,N_26312);
and U28479 (N_28479,N_26638,N_26209);
nor U28480 (N_28480,N_26882,N_26547);
xnor U28481 (N_28481,N_26032,N_27853);
and U28482 (N_28482,N_27060,N_26772);
xnor U28483 (N_28483,N_26415,N_27408);
or U28484 (N_28484,N_26667,N_26846);
nor U28485 (N_28485,N_26104,N_26931);
xnor U28486 (N_28486,N_27372,N_27479);
and U28487 (N_28487,N_26087,N_27317);
xnor U28488 (N_28488,N_26003,N_27796);
and U28489 (N_28489,N_27841,N_27120);
nand U28490 (N_28490,N_26206,N_26780);
xor U28491 (N_28491,N_27378,N_26151);
nand U28492 (N_28492,N_27177,N_26619);
or U28493 (N_28493,N_27905,N_26607);
and U28494 (N_28494,N_27743,N_26545);
nand U28495 (N_28495,N_27085,N_27928);
and U28496 (N_28496,N_27784,N_27660);
nor U28497 (N_28497,N_27369,N_27575);
and U28498 (N_28498,N_27418,N_27668);
nand U28499 (N_28499,N_27789,N_26040);
nand U28500 (N_28500,N_26266,N_26115);
and U28501 (N_28501,N_27488,N_26227);
nand U28502 (N_28502,N_26079,N_27218);
xnor U28503 (N_28503,N_27176,N_27722);
nand U28504 (N_28504,N_27083,N_26992);
xor U28505 (N_28505,N_27350,N_26687);
nor U28506 (N_28506,N_27724,N_26484);
nand U28507 (N_28507,N_27685,N_26267);
nor U28508 (N_28508,N_26224,N_26514);
and U28509 (N_28509,N_27016,N_26282);
xor U28510 (N_28510,N_26680,N_27119);
nand U28511 (N_28511,N_26257,N_26210);
xnor U28512 (N_28512,N_26830,N_26230);
and U28513 (N_28513,N_26374,N_26813);
nor U28514 (N_28514,N_27084,N_27539);
or U28515 (N_28515,N_26521,N_27203);
nor U28516 (N_28516,N_27267,N_26358);
nand U28517 (N_28517,N_26240,N_27509);
xnor U28518 (N_28518,N_26386,N_27735);
xnor U28519 (N_28519,N_27588,N_27619);
and U28520 (N_28520,N_26280,N_27548);
nor U28521 (N_28521,N_27558,N_26417);
nor U28522 (N_28522,N_27486,N_26361);
and U28523 (N_28523,N_27996,N_26214);
nor U28524 (N_28524,N_26793,N_27651);
xor U28525 (N_28525,N_27125,N_27993);
xor U28526 (N_28526,N_26397,N_27306);
nand U28527 (N_28527,N_27235,N_26444);
xor U28528 (N_28528,N_27468,N_26548);
nand U28529 (N_28529,N_27000,N_27129);
nand U28530 (N_28530,N_26362,N_26327);
and U28531 (N_28531,N_27599,N_27664);
nand U28532 (N_28532,N_26721,N_27699);
xnor U28533 (N_28533,N_27557,N_27014);
nand U28534 (N_28534,N_26914,N_26066);
and U28535 (N_28535,N_26460,N_26585);
and U28536 (N_28536,N_26149,N_27131);
xor U28537 (N_28537,N_26044,N_27860);
nand U28538 (N_28538,N_27263,N_27031);
nor U28539 (N_28539,N_27392,N_27483);
or U28540 (N_28540,N_27044,N_26671);
xor U28541 (N_28541,N_27793,N_27646);
nor U28542 (N_28542,N_27684,N_26895);
and U28543 (N_28543,N_27180,N_26769);
xnor U28544 (N_28544,N_27704,N_26334);
or U28545 (N_28545,N_27880,N_27771);
or U28546 (N_28546,N_26890,N_27727);
and U28547 (N_28547,N_26426,N_26790);
nor U28548 (N_28548,N_26756,N_26704);
xor U28549 (N_28549,N_27493,N_26523);
and U28550 (N_28550,N_27382,N_26001);
or U28551 (N_28551,N_26876,N_27606);
and U28552 (N_28552,N_26458,N_26617);
xor U28553 (N_28553,N_27373,N_26254);
nand U28554 (N_28554,N_27354,N_27219);
nand U28555 (N_28555,N_26567,N_27962);
nor U28556 (N_28556,N_26359,N_26111);
xnor U28557 (N_28557,N_27067,N_27754);
xnor U28558 (N_28558,N_26363,N_26196);
xnor U28559 (N_28559,N_26864,N_26559);
and U28560 (N_28560,N_27852,N_27917);
and U28561 (N_28561,N_26113,N_27258);
nand U28562 (N_28562,N_26008,N_26255);
or U28563 (N_28563,N_26531,N_26324);
xnor U28564 (N_28564,N_26425,N_26978);
nor U28565 (N_28565,N_27900,N_27846);
or U28566 (N_28566,N_26654,N_27197);
or U28567 (N_28567,N_26518,N_27953);
nand U28568 (N_28568,N_27200,N_27144);
and U28569 (N_28569,N_26511,N_27246);
or U28570 (N_28570,N_26832,N_26176);
and U28571 (N_28571,N_27700,N_27406);
and U28572 (N_28572,N_26251,N_26608);
and U28573 (N_28573,N_26543,N_26341);
nand U28574 (N_28574,N_26319,N_27285);
nand U28575 (N_28575,N_26084,N_27663);
and U28576 (N_28576,N_27839,N_27613);
and U28577 (N_28577,N_27898,N_26643);
or U28578 (N_28578,N_26786,N_26706);
or U28579 (N_28579,N_27101,N_26534);
nor U28580 (N_28580,N_26884,N_27692);
and U28581 (N_28581,N_27702,N_27954);
or U28582 (N_28582,N_27755,N_27295);
nand U28583 (N_28583,N_26476,N_27887);
nand U28584 (N_28584,N_27008,N_26470);
and U28585 (N_28585,N_26762,N_26843);
and U28586 (N_28586,N_27216,N_26184);
or U28587 (N_28587,N_26307,N_27497);
and U28588 (N_28588,N_27837,N_26213);
nor U28589 (N_28589,N_27813,N_27912);
or U28590 (N_28590,N_26774,N_26794);
nor U28591 (N_28591,N_27299,N_26968);
xor U28592 (N_28592,N_27002,N_26146);
nor U28593 (N_28593,N_27855,N_27786);
nand U28594 (N_28594,N_27949,N_27351);
and U28595 (N_28595,N_26665,N_26939);
nor U28596 (N_28596,N_27302,N_27502);
xnor U28597 (N_28597,N_27234,N_26247);
nor U28598 (N_28598,N_26059,N_26258);
or U28599 (N_28599,N_26365,N_26748);
nor U28600 (N_28600,N_26552,N_27321);
nor U28601 (N_28601,N_27196,N_27555);
nand U28602 (N_28602,N_26408,N_27907);
nand U28603 (N_28603,N_27726,N_27033);
xnor U28604 (N_28604,N_26013,N_27896);
xnor U28605 (N_28605,N_27915,N_26628);
and U28606 (N_28606,N_26261,N_27388);
nor U28607 (N_28607,N_27911,N_27916);
and U28608 (N_28608,N_27404,N_26937);
or U28609 (N_28609,N_26316,N_27580);
nand U28610 (N_28610,N_26927,N_26661);
xor U28611 (N_28611,N_26582,N_27746);
or U28612 (N_28612,N_26268,N_26099);
nand U28613 (N_28613,N_26293,N_26179);
nand U28614 (N_28614,N_26714,N_27779);
xor U28615 (N_28615,N_26046,N_26765);
or U28616 (N_28616,N_27353,N_27361);
nand U28617 (N_28617,N_27472,N_27139);
and U28618 (N_28618,N_27028,N_26562);
or U28619 (N_28619,N_27094,N_27178);
nor U28620 (N_28620,N_27518,N_27282);
or U28621 (N_28621,N_27021,N_26497);
xor U28622 (N_28622,N_26339,N_26606);
xnor U28623 (N_28623,N_27559,N_27574);
and U28624 (N_28624,N_26006,N_27644);
xor U28625 (N_28625,N_26023,N_27652);
and U28626 (N_28626,N_26018,N_27795);
xor U28627 (N_28627,N_26336,N_27942);
nand U28628 (N_28628,N_26670,N_27142);
and U28629 (N_28629,N_26190,N_27582);
or U28630 (N_28630,N_26128,N_26382);
nand U28631 (N_28631,N_26075,N_27464);
nor U28632 (N_28632,N_26618,N_26004);
and U28633 (N_28633,N_26669,N_27429);
nand U28634 (N_28634,N_27748,N_26229);
xor U28635 (N_28635,N_27937,N_27925);
and U28636 (N_28636,N_26997,N_27088);
and U28637 (N_28637,N_26471,N_26462);
and U28638 (N_28638,N_27782,N_26483);
nor U28639 (N_28639,N_26911,N_27995);
xnor U28640 (N_28640,N_26125,N_26811);
nand U28641 (N_28641,N_27959,N_26171);
xor U28642 (N_28642,N_27460,N_26642);
nand U28643 (N_28643,N_26249,N_26745);
nor U28644 (N_28644,N_27778,N_27966);
or U28645 (N_28645,N_26784,N_26411);
nor U28646 (N_28646,N_27411,N_26285);
or U28647 (N_28647,N_27035,N_27972);
nor U28648 (N_28648,N_26814,N_26560);
nand U28649 (N_28649,N_27253,N_27750);
nor U28650 (N_28650,N_27532,N_27840);
nand U28651 (N_28651,N_27759,N_26998);
nand U28652 (N_28652,N_26127,N_27478);
or U28653 (N_28653,N_26286,N_26659);
and U28654 (N_28654,N_27589,N_27205);
nor U28655 (N_28655,N_26012,N_27475);
xnor U28656 (N_28656,N_27602,N_27090);
xnor U28657 (N_28657,N_27787,N_27265);
nand U28658 (N_28658,N_27885,N_26612);
nand U28659 (N_28659,N_27820,N_27252);
xor U28660 (N_28660,N_26488,N_27667);
nor U28661 (N_28661,N_27015,N_26385);
or U28662 (N_28662,N_26342,N_27211);
nand U28663 (N_28663,N_27785,N_27199);
or U28664 (N_28664,N_27823,N_26613);
or U28665 (N_28665,N_26291,N_26439);
xor U28666 (N_28666,N_26693,N_26655);
xnor U28667 (N_28667,N_26237,N_26424);
and U28668 (N_28668,N_26972,N_27500);
xnor U28669 (N_28669,N_26520,N_27287);
and U28670 (N_28670,N_26434,N_26570);
nor U28671 (N_28671,N_27363,N_26788);
nand U28672 (N_28672,N_27590,N_26974);
and U28673 (N_28673,N_27442,N_27510);
and U28674 (N_28674,N_26203,N_27633);
xor U28675 (N_28675,N_27740,N_27100);
or U28676 (N_28676,N_26490,N_27043);
and U28677 (N_28677,N_27165,N_26118);
nor U28678 (N_28678,N_27542,N_26640);
nand U28679 (N_28679,N_26834,N_27984);
or U28680 (N_28680,N_27688,N_27848);
nand U28681 (N_28681,N_26371,N_27620);
nand U28682 (N_28682,N_27691,N_26862);
nand U28683 (N_28683,N_26791,N_26870);
and U28684 (N_28684,N_27886,N_27099);
or U28685 (N_28685,N_26506,N_27674);
or U28686 (N_28686,N_27137,N_26836);
or U28687 (N_28687,N_26404,N_26325);
nor U28688 (N_28688,N_26217,N_26842);
nand U28689 (N_28689,N_26903,N_26810);
and U28690 (N_28690,N_27422,N_26486);
xnor U28691 (N_28691,N_27512,N_27689);
nand U28692 (N_28692,N_27576,N_27739);
nand U28693 (N_28693,N_27181,N_27481);
nand U28694 (N_28694,N_27592,N_27325);
or U28695 (N_28695,N_27213,N_27275);
nor U28696 (N_28696,N_27524,N_27927);
nor U28697 (N_28697,N_26403,N_26037);
or U28698 (N_28698,N_26725,N_27172);
and U28699 (N_28699,N_26211,N_27632);
and U28700 (N_28700,N_27292,N_26947);
nand U28701 (N_28701,N_26622,N_26290);
nand U28702 (N_28702,N_26536,N_27041);
or U28703 (N_28703,N_27903,N_27529);
and U28704 (N_28704,N_27806,N_27653);
or U28705 (N_28705,N_26438,N_26941);
or U28706 (N_28706,N_26373,N_27029);
nor U28707 (N_28707,N_26959,N_26981);
xnor U28708 (N_28708,N_26701,N_26819);
and U28709 (N_28709,N_26353,N_26969);
nand U28710 (N_28710,N_27089,N_27419);
nand U28711 (N_28711,N_27435,N_27958);
nor U28712 (N_28712,N_26828,N_26279);
nand U28713 (N_28713,N_26899,N_26657);
or U28714 (N_28714,N_27622,N_26191);
xnor U28715 (N_28715,N_26976,N_27030);
and U28716 (N_28716,N_27143,N_26025);
xor U28717 (N_28717,N_27573,N_27111);
nor U28718 (N_28718,N_27179,N_26387);
or U28719 (N_28719,N_27899,N_27760);
nand U28720 (N_28720,N_27117,N_26277);
nand U28721 (N_28721,N_26347,N_27107);
nand U28722 (N_28722,N_26395,N_26393);
nor U28723 (N_28723,N_26598,N_27617);
xor U28724 (N_28724,N_27618,N_27323);
nand U28725 (N_28725,N_27081,N_27338);
or U28726 (N_28726,N_26960,N_27767);
xor U28727 (N_28727,N_27068,N_26581);
xor U28728 (N_28728,N_27010,N_26675);
or U28729 (N_28729,N_26182,N_27451);
and U28730 (N_28730,N_27830,N_27242);
or U28731 (N_28731,N_26625,N_27868);
and U28732 (N_28732,N_27140,N_27507);
and U28733 (N_28733,N_27777,N_27918);
or U28734 (N_28734,N_27311,N_27401);
xnor U28735 (N_28735,N_26123,N_26664);
nor U28736 (N_28736,N_27236,N_27690);
nand U28737 (N_28737,N_27233,N_27417);
and U28738 (N_28738,N_26703,N_27901);
nor U28739 (N_28739,N_27091,N_26027);
nor U28740 (N_28740,N_26754,N_26730);
xnor U28741 (N_28741,N_26504,N_27413);
nand U28742 (N_28742,N_26466,N_26354);
and U28743 (N_28743,N_26801,N_27471);
nand U28744 (N_28744,N_27814,N_27914);
nand U28745 (N_28745,N_26996,N_26463);
nand U28746 (N_28746,N_27491,N_27894);
nor U28747 (N_28747,N_26579,N_27192);
or U28748 (N_28748,N_26789,N_26063);
nor U28749 (N_28749,N_27809,N_27290);
nand U28750 (N_28750,N_26162,N_26117);
nor U28751 (N_28751,N_27459,N_26252);
and U28752 (N_28752,N_27256,N_27096);
nor U28753 (N_28753,N_26979,N_26767);
or U28754 (N_28754,N_27294,N_26768);
or U28755 (N_28755,N_27926,N_27850);
nor U28756 (N_28756,N_27713,N_26494);
nand U28757 (N_28757,N_27701,N_26648);
or U28758 (N_28758,N_27530,N_27365);
nor U28759 (N_28759,N_27709,N_27384);
and U28760 (N_28760,N_26174,N_27838);
nand U28761 (N_28761,N_27780,N_27344);
and U28762 (N_28762,N_26909,N_27013);
and U28763 (N_28763,N_27666,N_27842);
nand U28764 (N_28764,N_26114,N_27822);
and U28765 (N_28765,N_27829,N_27072);
xnor U28766 (N_28766,N_27994,N_27673);
nand U28767 (N_28767,N_26384,N_27836);
nor U28768 (N_28768,N_26448,N_26269);
nand U28769 (N_28769,N_27503,N_26505);
and U28770 (N_28770,N_27188,N_27676);
xnor U28771 (N_28771,N_26907,N_27776);
nor U28772 (N_28772,N_26797,N_26248);
or U28773 (N_28773,N_27379,N_27359);
or U28774 (N_28774,N_27523,N_26355);
nand U28775 (N_28775,N_26817,N_27055);
nor U28776 (N_28776,N_26954,N_26953);
or U28777 (N_28777,N_27169,N_26475);
and U28778 (N_28778,N_26989,N_27978);
and U28779 (N_28779,N_27374,N_26156);
xnor U28780 (N_28780,N_26541,N_27247);
nor U28781 (N_28781,N_27207,N_27336);
and U28782 (N_28782,N_26592,N_27003);
xnor U28783 (N_28783,N_26869,N_26274);
nand U28784 (N_28784,N_26090,N_27039);
xor U28785 (N_28785,N_27920,N_27064);
xor U28786 (N_28786,N_26435,N_27638);
nand U28787 (N_28787,N_27772,N_27281);
nand U28788 (N_28788,N_26134,N_26677);
and U28789 (N_28789,N_27537,N_27657);
or U28790 (N_28790,N_27280,N_26551);
or U28791 (N_28791,N_26601,N_27683);
and U28792 (N_28792,N_26844,N_27519);
xnor U28793 (N_28793,N_27020,N_27436);
nand U28794 (N_28794,N_26867,N_26955);
nand U28795 (N_28795,N_27228,N_26167);
and U28796 (N_28796,N_26464,N_26135);
xor U28797 (N_28797,N_27381,N_26639);
nand U28798 (N_28798,N_26938,N_26751);
and U28799 (N_28799,N_26501,N_26732);
nor U28800 (N_28800,N_26878,N_27182);
and U28801 (N_28801,N_26378,N_27127);
and U28802 (N_28802,N_26557,N_26835);
and U28803 (N_28803,N_27284,N_27309);
and U28804 (N_28804,N_27112,N_26816);
xor U28805 (N_28805,N_27717,N_26379);
or U28806 (N_28806,N_26321,N_26777);
nor U28807 (N_28807,N_27971,N_27541);
and U28808 (N_28808,N_27310,N_26731);
and U28809 (N_28809,N_27232,N_26681);
or U28810 (N_28810,N_26060,N_27368);
or U28811 (N_28811,N_27079,N_26626);
and U28812 (N_28812,N_27535,N_27158);
or U28813 (N_28813,N_26143,N_27051);
nor U28814 (N_28814,N_26646,N_27857);
xnor U28815 (N_28815,N_27909,N_26823);
nor U28816 (N_28816,N_27229,N_26919);
and U28817 (N_28817,N_27214,N_26920);
xnor U28818 (N_28818,N_26419,N_26775);
xnor U28819 (N_28819,N_26219,N_27808);
xnor U28820 (N_28820,N_27711,N_27631);
and U28821 (N_28821,N_27341,N_27473);
nand U28822 (N_28822,N_26621,N_26119);
nor U28823 (N_28823,N_27461,N_26929);
xor U28824 (N_28824,N_27774,N_26301);
nor U28825 (N_28825,N_27924,N_26170);
xnor U28826 (N_28826,N_27492,N_27610);
nor U28827 (N_28827,N_26849,N_26803);
nor U28828 (N_28828,N_27625,N_27669);
or U28829 (N_28829,N_26239,N_27869);
or U28830 (N_28830,N_26512,N_26636);
or U28831 (N_28831,N_27102,N_26653);
and U28832 (N_28832,N_26571,N_27696);
and U28833 (N_28833,N_27187,N_26700);
and U28834 (N_28834,N_27511,N_26245);
xnor U28835 (N_28835,N_27134,N_26116);
nor U28836 (N_28836,N_27130,N_26759);
and U28837 (N_28837,N_27872,N_27022);
xor U28838 (N_28838,N_27103,N_26193);
xor U28839 (N_28839,N_27070,N_26340);
nand U28840 (N_28840,N_26717,N_26802);
and U28841 (N_28841,N_27819,N_27783);
xnor U28842 (N_28842,N_27615,N_27426);
xnor U28843 (N_28843,N_27224,N_26986);
and U28844 (N_28844,N_26311,N_26866);
and U28845 (N_28845,N_26897,N_27126);
and U28846 (N_28846,N_26952,N_26300);
xor U28847 (N_28847,N_26163,N_27616);
or U28848 (N_28848,N_26141,N_27734);
and U28849 (N_28849,N_26155,N_26891);
and U28850 (N_28850,N_27154,N_27629);
and U28851 (N_28851,N_26688,N_27902);
nand U28852 (N_28852,N_26513,N_26010);
or U28853 (N_28853,N_26451,N_26684);
nand U28854 (N_28854,N_27272,N_26350);
and U28855 (N_28855,N_27171,N_27948);
nor U28856 (N_28856,N_26946,N_27230);
nor U28857 (N_28857,N_26472,N_27650);
xnor U28858 (N_28858,N_27095,N_27259);
and U28859 (N_28859,N_27420,N_26550);
nor U28860 (N_28860,N_26158,N_26740);
xnor U28861 (N_28861,N_27956,N_27571);
and U28862 (N_28862,N_27261,N_27428);
and U28863 (N_28863,N_27017,N_27409);
nor U28864 (N_28864,N_27412,N_26945);
nand U28865 (N_28865,N_26473,N_26263);
or U28866 (N_28866,N_27961,N_27546);
and U28867 (N_28867,N_26337,N_26132);
nand U28868 (N_28868,N_26851,N_27148);
or U28869 (N_28869,N_26566,N_26902);
nor U28870 (N_28870,N_26175,N_27097);
xor U28871 (N_28871,N_26039,N_26674);
xnor U28872 (N_28872,N_26154,N_27040);
nor U28873 (N_28873,N_26852,N_27065);
nor U28874 (N_28874,N_26728,N_27005);
or U28875 (N_28875,N_26317,N_26676);
and U28876 (N_28876,N_27348,N_27608);
and U28877 (N_28877,N_26243,N_26856);
nand U28878 (N_28878,N_27866,N_26637);
nor U28879 (N_28879,N_26246,N_27940);
or U28880 (N_28880,N_27578,N_26343);
and U28881 (N_28881,N_27714,N_27245);
xor U28882 (N_28882,N_27517,N_27832);
and U28883 (N_28883,N_27138,N_26746);
xnor U28884 (N_28884,N_27988,N_27766);
nand U28885 (N_28885,N_27301,N_26656);
or U28886 (N_28886,N_27118,N_26783);
nand U28887 (N_28887,N_26169,N_27052);
xor U28888 (N_28888,N_26896,N_27054);
xnor U28889 (N_28889,N_26537,N_26047);
nand U28890 (N_28890,N_26181,N_26131);
nor U28891 (N_28891,N_27308,N_26202);
nor U28892 (N_28892,N_27867,N_26338);
xor U28893 (N_28893,N_27788,N_27487);
nand U28894 (N_28894,N_26977,N_26303);
or U28895 (N_28895,N_26689,N_26800);
and U28896 (N_28896,N_26948,N_26734);
and U28897 (N_28897,N_27108,N_26785);
nor U28898 (N_28898,N_27587,N_27389);
and U28899 (N_28899,N_26838,N_27080);
or U28900 (N_28900,N_26016,N_26572);
xnor U28901 (N_28901,N_27415,N_26583);
and U28902 (N_28902,N_27851,N_27026);
nand U28903 (N_28903,N_26461,N_27480);
or U28904 (N_28904,N_27790,N_27598);
xnor U28905 (N_28905,N_26253,N_26093);
nor U28906 (N_28906,N_26857,N_27038);
or U28907 (N_28907,N_26705,N_27906);
and U28908 (N_28908,N_26822,N_27770);
nor U28909 (N_28909,N_27647,N_26807);
and U28910 (N_28910,N_26405,N_27596);
nand U28911 (N_28911,N_26738,N_26942);
nand U28912 (N_28912,N_27845,N_26145);
xnor U28913 (N_28913,N_26863,N_27799);
and U28914 (N_28914,N_26917,N_26328);
xnor U28915 (N_28915,N_26694,N_27884);
and U28916 (N_28916,N_27733,N_26443);
or U28917 (N_28917,N_26587,N_26297);
nor U28918 (N_28918,N_26402,N_27050);
nand U28919 (N_28919,N_27919,N_27969);
or U28920 (N_28920,N_27985,N_27680);
and U28921 (N_28921,N_26698,N_27921);
xnor U28922 (N_28922,N_26102,N_27979);
nand U28923 (N_28923,N_26133,N_26189);
xor U28924 (N_28924,N_26542,N_27642);
xor U28925 (N_28925,N_27220,N_27316);
and U28926 (N_28926,N_27720,N_27394);
xor U28927 (N_28927,N_27763,N_26031);
or U28928 (N_28928,N_27525,N_27977);
or U28929 (N_28929,N_27377,N_27694);
nand U28930 (N_28930,N_27864,N_26658);
nor U28931 (N_28931,N_27983,N_27607);
or U28932 (N_28932,N_26108,N_26650);
nand U28933 (N_28933,N_27648,N_26036);
and U28934 (N_28934,N_26589,N_27791);
and U28935 (N_28935,N_26886,N_26447);
xor U28936 (N_28936,N_27427,N_27159);
and U28937 (N_28937,N_27681,N_27570);
nand U28938 (N_28938,N_26691,N_26139);
and U28939 (N_28939,N_26283,N_27612);
and U28940 (N_28940,N_26925,N_26766);
nor U28941 (N_28941,N_26205,N_27371);
xor U28942 (N_28942,N_26109,N_26591);
or U28943 (N_28943,N_27053,N_27136);
nand U28944 (N_28944,N_26124,N_27732);
nor U28945 (N_28945,N_26049,N_26798);
or U28946 (N_28946,N_27209,N_27816);
nand U28947 (N_28947,N_26871,N_27758);
or U28948 (N_28948,N_26859,N_26014);
and U28949 (N_28949,N_26160,N_26932);
nor U28950 (N_28950,N_27106,N_27286);
or U28951 (N_28951,N_26934,N_26200);
nor U28952 (N_28952,N_26881,N_27992);
nor U28953 (N_28953,N_26662,N_26110);
or U28954 (N_28954,N_27873,N_26757);
or U28955 (N_28955,N_26906,N_26121);
xnor U28956 (N_28956,N_26673,N_27009);
xor U28957 (N_28957,N_27324,N_27006);
nor U28958 (N_28958,N_26973,N_27730);
or U28959 (N_28959,N_27225,N_26078);
or U28960 (N_28960,N_26048,N_26351);
or U28961 (N_28961,N_26699,N_27399);
or U28962 (N_28962,N_27964,N_27731);
nor U28963 (N_28963,N_27161,N_26565);
nand U28964 (N_28964,N_27649,N_27707);
nand U28965 (N_28965,N_27991,N_26936);
nand U28966 (N_28966,N_26272,N_26965);
nand U28967 (N_28967,N_26220,N_27116);
xnor U28968 (N_28968,N_26414,N_26833);
and U28969 (N_28969,N_27360,N_26887);
xor U28970 (N_28970,N_26428,N_27312);
or U28971 (N_28971,N_27764,N_27448);
nand U28972 (N_28972,N_27243,N_26956);
xnor U28973 (N_28973,N_27457,N_27798);
nand U28974 (N_28974,N_26381,N_27414);
nor U28975 (N_28975,N_26445,N_26278);
and U28976 (N_28976,N_26951,N_27078);
nor U28977 (N_28977,N_26457,N_26423);
nor U28978 (N_28978,N_26901,N_26416);
or U28979 (N_28979,N_27086,N_26812);
and U28980 (N_28980,N_26991,N_26062);
nand U28981 (N_28981,N_26024,N_27201);
nand U28982 (N_28982,N_27826,N_26602);
nand U28983 (N_28983,N_26398,N_27380);
xor U28984 (N_28984,N_27950,N_27976);
nand U28985 (N_28985,N_27904,N_26696);
nor U28986 (N_28986,N_27204,N_27433);
xor U28987 (N_28987,N_27934,N_26096);
nand U28988 (N_28988,N_27300,N_27307);
or U28989 (N_28989,N_27175,N_27482);
nor U28990 (N_28990,N_26538,N_26348);
xnor U28991 (N_28991,N_26410,N_27337);
xnor U28992 (N_28992,N_26299,N_27202);
xnor U28993 (N_28993,N_27637,N_26399);
xnor U28994 (N_28994,N_26065,N_26517);
xor U28995 (N_28995,N_27536,N_27725);
and U28996 (N_28996,N_26345,N_27467);
or U28997 (N_28997,N_26627,N_26949);
xor U28998 (N_28998,N_26546,N_26809);
or U28999 (N_28999,N_26441,N_27721);
nand U29000 (N_29000,N_27450,N_27514);
nor U29001 (N_29001,N_26444,N_26641);
or U29002 (N_29002,N_26641,N_26721);
and U29003 (N_29003,N_27182,N_26098);
and U29004 (N_29004,N_27581,N_26480);
nand U29005 (N_29005,N_26857,N_26209);
nor U29006 (N_29006,N_26272,N_27607);
xnor U29007 (N_29007,N_27706,N_26553);
or U29008 (N_29008,N_26812,N_26435);
xnor U29009 (N_29009,N_26624,N_27009);
xnor U29010 (N_29010,N_27401,N_27895);
and U29011 (N_29011,N_26857,N_26501);
nand U29012 (N_29012,N_26088,N_27083);
nand U29013 (N_29013,N_27215,N_27068);
nor U29014 (N_29014,N_26333,N_27644);
or U29015 (N_29015,N_26174,N_26692);
nand U29016 (N_29016,N_26238,N_26959);
or U29017 (N_29017,N_27855,N_26784);
nor U29018 (N_29018,N_27828,N_27931);
nand U29019 (N_29019,N_27468,N_26905);
nor U29020 (N_29020,N_27586,N_27811);
xnor U29021 (N_29021,N_27274,N_27791);
and U29022 (N_29022,N_26596,N_27878);
xor U29023 (N_29023,N_27706,N_27724);
or U29024 (N_29024,N_26493,N_26926);
or U29025 (N_29025,N_26301,N_27106);
or U29026 (N_29026,N_26581,N_27430);
xor U29027 (N_29027,N_27836,N_26962);
and U29028 (N_29028,N_26170,N_27993);
nor U29029 (N_29029,N_26211,N_27465);
or U29030 (N_29030,N_27996,N_27093);
nand U29031 (N_29031,N_27315,N_27655);
nand U29032 (N_29032,N_27068,N_26100);
nor U29033 (N_29033,N_27716,N_26859);
or U29034 (N_29034,N_27661,N_26811);
xnor U29035 (N_29035,N_27827,N_26769);
xor U29036 (N_29036,N_26409,N_26936);
and U29037 (N_29037,N_27745,N_26991);
and U29038 (N_29038,N_26993,N_27705);
nand U29039 (N_29039,N_26712,N_26659);
and U29040 (N_29040,N_27803,N_27684);
nor U29041 (N_29041,N_26531,N_26487);
xnor U29042 (N_29042,N_27937,N_27226);
nand U29043 (N_29043,N_26373,N_27987);
and U29044 (N_29044,N_27022,N_26818);
nor U29045 (N_29045,N_27835,N_27559);
or U29046 (N_29046,N_26404,N_27316);
or U29047 (N_29047,N_26716,N_26705);
nand U29048 (N_29048,N_26415,N_27424);
nand U29049 (N_29049,N_27749,N_27992);
or U29050 (N_29050,N_26702,N_27513);
xor U29051 (N_29051,N_26120,N_27918);
nor U29052 (N_29052,N_26908,N_26020);
and U29053 (N_29053,N_27875,N_26226);
xnor U29054 (N_29054,N_26588,N_26297);
or U29055 (N_29055,N_27251,N_27427);
nand U29056 (N_29056,N_26111,N_27533);
and U29057 (N_29057,N_26623,N_26944);
or U29058 (N_29058,N_27323,N_27970);
xor U29059 (N_29059,N_26316,N_27646);
and U29060 (N_29060,N_27571,N_27061);
nand U29061 (N_29061,N_26220,N_27820);
nand U29062 (N_29062,N_27035,N_26693);
nor U29063 (N_29063,N_27418,N_27881);
nor U29064 (N_29064,N_27252,N_27744);
nand U29065 (N_29065,N_27953,N_27743);
or U29066 (N_29066,N_26334,N_26923);
or U29067 (N_29067,N_26370,N_26954);
nand U29068 (N_29068,N_27557,N_26216);
nand U29069 (N_29069,N_26073,N_26456);
and U29070 (N_29070,N_27902,N_26631);
xor U29071 (N_29071,N_26699,N_27912);
xor U29072 (N_29072,N_27298,N_27260);
nand U29073 (N_29073,N_26244,N_27624);
or U29074 (N_29074,N_26290,N_26695);
and U29075 (N_29075,N_27432,N_26368);
nand U29076 (N_29076,N_27518,N_27124);
nor U29077 (N_29077,N_26715,N_26585);
or U29078 (N_29078,N_26362,N_26851);
nand U29079 (N_29079,N_26419,N_26572);
and U29080 (N_29080,N_26030,N_26321);
and U29081 (N_29081,N_27617,N_27220);
nor U29082 (N_29082,N_27022,N_27611);
xor U29083 (N_29083,N_26211,N_26045);
nor U29084 (N_29084,N_27691,N_26757);
or U29085 (N_29085,N_26639,N_26660);
nand U29086 (N_29086,N_26507,N_26150);
and U29087 (N_29087,N_27000,N_27896);
and U29088 (N_29088,N_27227,N_26859);
nand U29089 (N_29089,N_27027,N_27456);
and U29090 (N_29090,N_26621,N_27303);
nand U29091 (N_29091,N_27867,N_26498);
xnor U29092 (N_29092,N_27175,N_26273);
xor U29093 (N_29093,N_27609,N_27205);
or U29094 (N_29094,N_26228,N_27495);
or U29095 (N_29095,N_26263,N_27404);
xnor U29096 (N_29096,N_26436,N_26967);
nand U29097 (N_29097,N_27713,N_27977);
or U29098 (N_29098,N_27964,N_26383);
or U29099 (N_29099,N_26033,N_26421);
xnor U29100 (N_29100,N_27304,N_26556);
nand U29101 (N_29101,N_26009,N_27787);
or U29102 (N_29102,N_27710,N_26231);
and U29103 (N_29103,N_27264,N_27785);
xnor U29104 (N_29104,N_27564,N_26773);
nor U29105 (N_29105,N_26480,N_27499);
or U29106 (N_29106,N_27567,N_26439);
nand U29107 (N_29107,N_26950,N_26471);
or U29108 (N_29108,N_27694,N_26588);
nand U29109 (N_29109,N_26633,N_27538);
or U29110 (N_29110,N_26922,N_27292);
nand U29111 (N_29111,N_27809,N_26431);
and U29112 (N_29112,N_27606,N_27134);
xor U29113 (N_29113,N_26886,N_27673);
and U29114 (N_29114,N_27087,N_26430);
xor U29115 (N_29115,N_27357,N_27851);
nand U29116 (N_29116,N_26178,N_26827);
or U29117 (N_29117,N_26896,N_27495);
xnor U29118 (N_29118,N_27483,N_27439);
nand U29119 (N_29119,N_27119,N_26084);
and U29120 (N_29120,N_26192,N_27321);
or U29121 (N_29121,N_26421,N_27037);
nand U29122 (N_29122,N_26102,N_26862);
nor U29123 (N_29123,N_26767,N_27028);
xor U29124 (N_29124,N_27954,N_27286);
and U29125 (N_29125,N_26494,N_27975);
and U29126 (N_29126,N_27218,N_26043);
xnor U29127 (N_29127,N_26139,N_27286);
nand U29128 (N_29128,N_26093,N_26305);
xnor U29129 (N_29129,N_26706,N_26306);
nor U29130 (N_29130,N_27012,N_26602);
xor U29131 (N_29131,N_26676,N_27062);
nor U29132 (N_29132,N_26968,N_26738);
nor U29133 (N_29133,N_27091,N_26770);
and U29134 (N_29134,N_26740,N_27382);
xor U29135 (N_29135,N_26441,N_27993);
nand U29136 (N_29136,N_27989,N_26320);
nor U29137 (N_29137,N_27837,N_26959);
xor U29138 (N_29138,N_27642,N_26163);
or U29139 (N_29139,N_27791,N_26924);
nand U29140 (N_29140,N_27140,N_27993);
and U29141 (N_29141,N_27372,N_27738);
or U29142 (N_29142,N_27530,N_27140);
or U29143 (N_29143,N_27866,N_27844);
nand U29144 (N_29144,N_26412,N_27089);
or U29145 (N_29145,N_27928,N_26435);
and U29146 (N_29146,N_26293,N_27265);
or U29147 (N_29147,N_26478,N_26460);
or U29148 (N_29148,N_26768,N_26247);
nand U29149 (N_29149,N_27693,N_26899);
nand U29150 (N_29150,N_26484,N_26979);
or U29151 (N_29151,N_27299,N_27455);
nand U29152 (N_29152,N_26348,N_27215);
xor U29153 (N_29153,N_26658,N_27381);
xnor U29154 (N_29154,N_26835,N_27697);
and U29155 (N_29155,N_26163,N_26840);
or U29156 (N_29156,N_27316,N_26723);
xnor U29157 (N_29157,N_26247,N_26061);
xnor U29158 (N_29158,N_26815,N_26803);
or U29159 (N_29159,N_27152,N_27738);
or U29160 (N_29160,N_27199,N_26909);
nor U29161 (N_29161,N_27387,N_27272);
and U29162 (N_29162,N_26620,N_26903);
nor U29163 (N_29163,N_27487,N_27221);
or U29164 (N_29164,N_26387,N_27842);
nand U29165 (N_29165,N_26732,N_27855);
xnor U29166 (N_29166,N_27626,N_26878);
or U29167 (N_29167,N_27096,N_27517);
xnor U29168 (N_29168,N_27905,N_27926);
nor U29169 (N_29169,N_26778,N_26508);
nand U29170 (N_29170,N_27222,N_26996);
nor U29171 (N_29171,N_27130,N_26069);
nor U29172 (N_29172,N_26464,N_26327);
nor U29173 (N_29173,N_26593,N_27342);
or U29174 (N_29174,N_27696,N_27568);
xnor U29175 (N_29175,N_26956,N_27735);
and U29176 (N_29176,N_27889,N_27704);
and U29177 (N_29177,N_27469,N_26363);
nand U29178 (N_29178,N_26071,N_26844);
nor U29179 (N_29179,N_26590,N_26926);
and U29180 (N_29180,N_26983,N_27044);
nor U29181 (N_29181,N_26247,N_27799);
nand U29182 (N_29182,N_26312,N_27525);
or U29183 (N_29183,N_26937,N_27550);
nor U29184 (N_29184,N_26867,N_27170);
nor U29185 (N_29185,N_27155,N_27529);
xnor U29186 (N_29186,N_27738,N_26019);
xnor U29187 (N_29187,N_27065,N_27224);
and U29188 (N_29188,N_26346,N_27233);
and U29189 (N_29189,N_26860,N_26040);
or U29190 (N_29190,N_26463,N_26178);
nor U29191 (N_29191,N_26703,N_27012);
xor U29192 (N_29192,N_27906,N_26961);
or U29193 (N_29193,N_26264,N_26437);
or U29194 (N_29194,N_26008,N_27804);
nand U29195 (N_29195,N_26117,N_27668);
or U29196 (N_29196,N_26660,N_26638);
and U29197 (N_29197,N_26568,N_27958);
or U29198 (N_29198,N_26054,N_26696);
and U29199 (N_29199,N_27913,N_26917);
nand U29200 (N_29200,N_27919,N_26144);
xor U29201 (N_29201,N_26969,N_27229);
xnor U29202 (N_29202,N_27851,N_27207);
nand U29203 (N_29203,N_26255,N_27763);
xnor U29204 (N_29204,N_27229,N_26124);
or U29205 (N_29205,N_27266,N_26599);
or U29206 (N_29206,N_26291,N_27224);
nor U29207 (N_29207,N_27372,N_26380);
and U29208 (N_29208,N_26092,N_26945);
and U29209 (N_29209,N_26605,N_26528);
or U29210 (N_29210,N_26049,N_27807);
nor U29211 (N_29211,N_26123,N_26111);
nand U29212 (N_29212,N_26145,N_26605);
or U29213 (N_29213,N_27712,N_26803);
nor U29214 (N_29214,N_27126,N_26726);
nand U29215 (N_29215,N_27512,N_26909);
nor U29216 (N_29216,N_26699,N_26070);
nor U29217 (N_29217,N_27632,N_27565);
and U29218 (N_29218,N_27410,N_27800);
nand U29219 (N_29219,N_27087,N_27225);
nor U29220 (N_29220,N_27613,N_26022);
or U29221 (N_29221,N_27275,N_26391);
nand U29222 (N_29222,N_27568,N_27250);
nand U29223 (N_29223,N_27412,N_27853);
or U29224 (N_29224,N_26011,N_26128);
xor U29225 (N_29225,N_27695,N_26446);
nor U29226 (N_29226,N_27500,N_27958);
and U29227 (N_29227,N_26256,N_27059);
and U29228 (N_29228,N_26101,N_26792);
and U29229 (N_29229,N_27485,N_26244);
and U29230 (N_29230,N_26407,N_27710);
nor U29231 (N_29231,N_27739,N_27131);
and U29232 (N_29232,N_26289,N_27512);
nand U29233 (N_29233,N_27967,N_27826);
xor U29234 (N_29234,N_26187,N_27913);
nand U29235 (N_29235,N_26977,N_26133);
or U29236 (N_29236,N_26190,N_26222);
or U29237 (N_29237,N_27565,N_26305);
xnor U29238 (N_29238,N_26242,N_26118);
or U29239 (N_29239,N_26852,N_26315);
or U29240 (N_29240,N_27633,N_26370);
xor U29241 (N_29241,N_27644,N_26447);
and U29242 (N_29242,N_27220,N_26395);
or U29243 (N_29243,N_27383,N_26152);
or U29244 (N_29244,N_27835,N_27479);
nor U29245 (N_29245,N_27336,N_26493);
nand U29246 (N_29246,N_26403,N_26286);
or U29247 (N_29247,N_27843,N_26878);
and U29248 (N_29248,N_27179,N_26639);
and U29249 (N_29249,N_27125,N_27461);
and U29250 (N_29250,N_27429,N_26578);
or U29251 (N_29251,N_26100,N_26615);
nor U29252 (N_29252,N_26555,N_26224);
xnor U29253 (N_29253,N_26618,N_27219);
nand U29254 (N_29254,N_26397,N_26941);
nand U29255 (N_29255,N_27687,N_27727);
and U29256 (N_29256,N_27610,N_27434);
nand U29257 (N_29257,N_26268,N_27769);
xor U29258 (N_29258,N_27712,N_26619);
and U29259 (N_29259,N_27282,N_27432);
nand U29260 (N_29260,N_26695,N_27062);
xnor U29261 (N_29261,N_27340,N_27465);
nor U29262 (N_29262,N_27369,N_26014);
xnor U29263 (N_29263,N_27978,N_27679);
xor U29264 (N_29264,N_26823,N_26310);
and U29265 (N_29265,N_26467,N_27867);
nor U29266 (N_29266,N_26435,N_26843);
nand U29267 (N_29267,N_27819,N_26057);
xnor U29268 (N_29268,N_26759,N_26415);
or U29269 (N_29269,N_27284,N_26243);
xnor U29270 (N_29270,N_27241,N_26651);
xnor U29271 (N_29271,N_26091,N_27799);
nand U29272 (N_29272,N_26264,N_27100);
nor U29273 (N_29273,N_27573,N_26156);
and U29274 (N_29274,N_27318,N_27171);
nor U29275 (N_29275,N_27463,N_26258);
xnor U29276 (N_29276,N_26176,N_27233);
and U29277 (N_29277,N_27069,N_27187);
nor U29278 (N_29278,N_26870,N_26675);
xnor U29279 (N_29279,N_27522,N_27887);
xor U29280 (N_29280,N_26848,N_26911);
xor U29281 (N_29281,N_27428,N_27245);
nand U29282 (N_29282,N_27776,N_27810);
xnor U29283 (N_29283,N_26743,N_27670);
or U29284 (N_29284,N_27078,N_26772);
nor U29285 (N_29285,N_26013,N_26594);
or U29286 (N_29286,N_27149,N_26086);
nor U29287 (N_29287,N_27748,N_26452);
and U29288 (N_29288,N_27280,N_26894);
nand U29289 (N_29289,N_27532,N_27054);
and U29290 (N_29290,N_26108,N_26492);
xor U29291 (N_29291,N_26804,N_27975);
nor U29292 (N_29292,N_26889,N_27430);
and U29293 (N_29293,N_27647,N_27572);
nor U29294 (N_29294,N_26909,N_27043);
nor U29295 (N_29295,N_26813,N_26193);
and U29296 (N_29296,N_26373,N_27811);
or U29297 (N_29297,N_26161,N_26723);
xnor U29298 (N_29298,N_26120,N_27694);
nand U29299 (N_29299,N_27590,N_26097);
and U29300 (N_29300,N_27117,N_27760);
xor U29301 (N_29301,N_26897,N_26951);
and U29302 (N_29302,N_26264,N_27284);
and U29303 (N_29303,N_27593,N_27693);
nor U29304 (N_29304,N_27774,N_26520);
xnor U29305 (N_29305,N_27390,N_27927);
xnor U29306 (N_29306,N_27624,N_26580);
nand U29307 (N_29307,N_26371,N_26741);
nand U29308 (N_29308,N_27607,N_27688);
nand U29309 (N_29309,N_27208,N_26612);
nand U29310 (N_29310,N_26699,N_26769);
and U29311 (N_29311,N_27457,N_27359);
nor U29312 (N_29312,N_26788,N_27177);
nor U29313 (N_29313,N_26585,N_26919);
nor U29314 (N_29314,N_26950,N_27645);
xor U29315 (N_29315,N_27253,N_27167);
and U29316 (N_29316,N_27128,N_27409);
xnor U29317 (N_29317,N_27339,N_26348);
and U29318 (N_29318,N_27082,N_27364);
or U29319 (N_29319,N_26467,N_26838);
nand U29320 (N_29320,N_27116,N_27019);
and U29321 (N_29321,N_26077,N_27244);
or U29322 (N_29322,N_26688,N_26999);
or U29323 (N_29323,N_27045,N_26057);
nor U29324 (N_29324,N_26890,N_27753);
xnor U29325 (N_29325,N_26877,N_26379);
xnor U29326 (N_29326,N_27952,N_26425);
and U29327 (N_29327,N_26583,N_27593);
and U29328 (N_29328,N_26381,N_26052);
or U29329 (N_29329,N_26205,N_26498);
nor U29330 (N_29330,N_26646,N_26732);
xor U29331 (N_29331,N_26569,N_27350);
and U29332 (N_29332,N_26997,N_26718);
nand U29333 (N_29333,N_27180,N_26223);
nor U29334 (N_29334,N_27241,N_27826);
nand U29335 (N_29335,N_26548,N_26774);
or U29336 (N_29336,N_26788,N_27258);
nand U29337 (N_29337,N_26503,N_26519);
nor U29338 (N_29338,N_27066,N_26124);
and U29339 (N_29339,N_27081,N_26186);
nor U29340 (N_29340,N_26308,N_27815);
or U29341 (N_29341,N_27677,N_27993);
or U29342 (N_29342,N_26906,N_26180);
and U29343 (N_29343,N_27769,N_27899);
or U29344 (N_29344,N_26423,N_27848);
nor U29345 (N_29345,N_27273,N_27363);
nand U29346 (N_29346,N_26216,N_27416);
xnor U29347 (N_29347,N_27861,N_26487);
nand U29348 (N_29348,N_27293,N_26416);
xnor U29349 (N_29349,N_27321,N_26244);
xor U29350 (N_29350,N_27859,N_26298);
or U29351 (N_29351,N_27872,N_26762);
and U29352 (N_29352,N_26394,N_26953);
nor U29353 (N_29353,N_26494,N_27504);
xnor U29354 (N_29354,N_26973,N_27312);
and U29355 (N_29355,N_27558,N_26575);
nand U29356 (N_29356,N_27183,N_27001);
and U29357 (N_29357,N_26495,N_27230);
nor U29358 (N_29358,N_27939,N_27445);
or U29359 (N_29359,N_27245,N_26008);
or U29360 (N_29360,N_26143,N_26333);
or U29361 (N_29361,N_26283,N_26535);
nor U29362 (N_29362,N_27430,N_27168);
nand U29363 (N_29363,N_27756,N_26007);
or U29364 (N_29364,N_26641,N_27172);
nand U29365 (N_29365,N_26200,N_27762);
xor U29366 (N_29366,N_26207,N_26296);
or U29367 (N_29367,N_26672,N_27455);
xnor U29368 (N_29368,N_27442,N_27007);
nand U29369 (N_29369,N_27404,N_27004);
nor U29370 (N_29370,N_26403,N_27212);
xor U29371 (N_29371,N_26045,N_27152);
and U29372 (N_29372,N_27661,N_27554);
and U29373 (N_29373,N_26495,N_26733);
and U29374 (N_29374,N_26502,N_27439);
or U29375 (N_29375,N_26796,N_26584);
nor U29376 (N_29376,N_26474,N_27639);
nor U29377 (N_29377,N_27301,N_27819);
nor U29378 (N_29378,N_26020,N_26717);
or U29379 (N_29379,N_26334,N_27894);
xor U29380 (N_29380,N_26971,N_26220);
or U29381 (N_29381,N_26509,N_26436);
and U29382 (N_29382,N_26370,N_27487);
or U29383 (N_29383,N_26675,N_27564);
or U29384 (N_29384,N_26660,N_26161);
or U29385 (N_29385,N_26842,N_26146);
xor U29386 (N_29386,N_26619,N_26652);
nand U29387 (N_29387,N_26386,N_27741);
and U29388 (N_29388,N_27662,N_27409);
and U29389 (N_29389,N_27833,N_26576);
nor U29390 (N_29390,N_27743,N_27849);
nand U29391 (N_29391,N_27487,N_27813);
and U29392 (N_29392,N_27278,N_26440);
or U29393 (N_29393,N_27404,N_26465);
or U29394 (N_29394,N_27311,N_26554);
nor U29395 (N_29395,N_26563,N_26341);
nand U29396 (N_29396,N_26113,N_27125);
or U29397 (N_29397,N_26033,N_27004);
and U29398 (N_29398,N_26033,N_27264);
nand U29399 (N_29399,N_27490,N_26492);
xor U29400 (N_29400,N_26224,N_27244);
xnor U29401 (N_29401,N_26631,N_26594);
or U29402 (N_29402,N_26547,N_27859);
xor U29403 (N_29403,N_26422,N_27409);
and U29404 (N_29404,N_27250,N_26292);
nor U29405 (N_29405,N_27312,N_26535);
nand U29406 (N_29406,N_27491,N_26732);
and U29407 (N_29407,N_27709,N_26271);
or U29408 (N_29408,N_27461,N_26566);
nor U29409 (N_29409,N_26482,N_27863);
and U29410 (N_29410,N_27941,N_26937);
nand U29411 (N_29411,N_27400,N_27010);
nand U29412 (N_29412,N_26567,N_26593);
nor U29413 (N_29413,N_26988,N_27810);
and U29414 (N_29414,N_26554,N_27625);
nand U29415 (N_29415,N_27296,N_27497);
nor U29416 (N_29416,N_27922,N_27304);
xnor U29417 (N_29417,N_27750,N_27393);
xor U29418 (N_29418,N_26538,N_26148);
xnor U29419 (N_29419,N_27518,N_27110);
nand U29420 (N_29420,N_26904,N_27753);
nand U29421 (N_29421,N_27505,N_27405);
nor U29422 (N_29422,N_27001,N_26228);
nand U29423 (N_29423,N_26236,N_26460);
nor U29424 (N_29424,N_26988,N_26252);
xnor U29425 (N_29425,N_26604,N_27124);
nor U29426 (N_29426,N_26722,N_27146);
nor U29427 (N_29427,N_27173,N_26022);
xnor U29428 (N_29428,N_26378,N_27387);
xnor U29429 (N_29429,N_26674,N_26211);
or U29430 (N_29430,N_27276,N_27513);
or U29431 (N_29431,N_26309,N_27996);
xnor U29432 (N_29432,N_26993,N_27588);
nand U29433 (N_29433,N_27767,N_27025);
nand U29434 (N_29434,N_27953,N_27322);
nor U29435 (N_29435,N_26123,N_26845);
and U29436 (N_29436,N_27964,N_26266);
or U29437 (N_29437,N_26717,N_27780);
nand U29438 (N_29438,N_26225,N_27632);
nand U29439 (N_29439,N_27623,N_26543);
and U29440 (N_29440,N_27461,N_26127);
and U29441 (N_29441,N_27011,N_26121);
nand U29442 (N_29442,N_26666,N_26390);
xnor U29443 (N_29443,N_26956,N_26108);
nor U29444 (N_29444,N_27724,N_26207);
or U29445 (N_29445,N_26138,N_27083);
and U29446 (N_29446,N_27766,N_26312);
xor U29447 (N_29447,N_26779,N_26613);
nor U29448 (N_29448,N_27831,N_26296);
nand U29449 (N_29449,N_26799,N_26737);
or U29450 (N_29450,N_26424,N_26869);
nand U29451 (N_29451,N_27982,N_27692);
xor U29452 (N_29452,N_26532,N_26803);
and U29453 (N_29453,N_27519,N_26450);
nor U29454 (N_29454,N_26431,N_27824);
nand U29455 (N_29455,N_27975,N_26369);
and U29456 (N_29456,N_26497,N_26534);
nand U29457 (N_29457,N_27648,N_27583);
and U29458 (N_29458,N_27257,N_27707);
or U29459 (N_29459,N_26354,N_26491);
or U29460 (N_29460,N_26727,N_27098);
and U29461 (N_29461,N_27838,N_26597);
and U29462 (N_29462,N_27727,N_26571);
or U29463 (N_29463,N_26150,N_26992);
nand U29464 (N_29464,N_26048,N_27057);
or U29465 (N_29465,N_27892,N_26777);
nor U29466 (N_29466,N_26706,N_27987);
nand U29467 (N_29467,N_26800,N_26325);
or U29468 (N_29468,N_26479,N_26235);
or U29469 (N_29469,N_26306,N_27542);
nor U29470 (N_29470,N_26479,N_26025);
nand U29471 (N_29471,N_27508,N_26320);
nand U29472 (N_29472,N_26917,N_26911);
nor U29473 (N_29473,N_26553,N_27169);
nand U29474 (N_29474,N_27139,N_26625);
nand U29475 (N_29475,N_27575,N_27219);
and U29476 (N_29476,N_26307,N_26234);
nand U29477 (N_29477,N_27998,N_27551);
or U29478 (N_29478,N_26398,N_27905);
nor U29479 (N_29479,N_27617,N_26823);
nand U29480 (N_29480,N_26546,N_26877);
nand U29481 (N_29481,N_27083,N_26517);
or U29482 (N_29482,N_26048,N_26982);
or U29483 (N_29483,N_26457,N_26239);
nor U29484 (N_29484,N_27186,N_26390);
nand U29485 (N_29485,N_27649,N_27645);
or U29486 (N_29486,N_27794,N_26377);
and U29487 (N_29487,N_26668,N_26535);
xnor U29488 (N_29488,N_26917,N_26118);
xor U29489 (N_29489,N_27525,N_26588);
and U29490 (N_29490,N_27008,N_26624);
or U29491 (N_29491,N_26022,N_27747);
or U29492 (N_29492,N_26183,N_27063);
nand U29493 (N_29493,N_27919,N_26528);
nand U29494 (N_29494,N_27079,N_26394);
nor U29495 (N_29495,N_27057,N_27717);
xnor U29496 (N_29496,N_27581,N_27472);
and U29497 (N_29497,N_27336,N_26149);
and U29498 (N_29498,N_26104,N_26903);
xnor U29499 (N_29499,N_27226,N_27006);
or U29500 (N_29500,N_26747,N_27204);
or U29501 (N_29501,N_26043,N_27470);
or U29502 (N_29502,N_26156,N_26795);
or U29503 (N_29503,N_26461,N_26308);
nor U29504 (N_29504,N_26990,N_26333);
nand U29505 (N_29505,N_26287,N_26779);
nand U29506 (N_29506,N_26467,N_26514);
or U29507 (N_29507,N_26112,N_26467);
nor U29508 (N_29508,N_26182,N_26684);
and U29509 (N_29509,N_27401,N_27398);
nor U29510 (N_29510,N_27922,N_27256);
xnor U29511 (N_29511,N_26359,N_27054);
and U29512 (N_29512,N_27205,N_27147);
xnor U29513 (N_29513,N_26927,N_27682);
nor U29514 (N_29514,N_26284,N_26173);
or U29515 (N_29515,N_26148,N_27365);
and U29516 (N_29516,N_27346,N_26767);
and U29517 (N_29517,N_26219,N_26792);
and U29518 (N_29518,N_26202,N_26210);
xnor U29519 (N_29519,N_27685,N_27235);
or U29520 (N_29520,N_26770,N_27952);
nor U29521 (N_29521,N_26080,N_26553);
nand U29522 (N_29522,N_27954,N_26905);
nor U29523 (N_29523,N_27058,N_26844);
xor U29524 (N_29524,N_27409,N_27881);
nor U29525 (N_29525,N_27566,N_26887);
or U29526 (N_29526,N_27353,N_26097);
xnor U29527 (N_29527,N_26542,N_27643);
and U29528 (N_29528,N_26881,N_27617);
nor U29529 (N_29529,N_27474,N_27471);
nor U29530 (N_29530,N_27685,N_26992);
and U29531 (N_29531,N_26599,N_26514);
xnor U29532 (N_29532,N_27042,N_26694);
or U29533 (N_29533,N_26580,N_26512);
nor U29534 (N_29534,N_27986,N_27029);
nor U29535 (N_29535,N_26418,N_27948);
xnor U29536 (N_29536,N_26762,N_26958);
nand U29537 (N_29537,N_27215,N_26918);
and U29538 (N_29538,N_27145,N_26823);
nor U29539 (N_29539,N_26362,N_27362);
xnor U29540 (N_29540,N_27389,N_26541);
nor U29541 (N_29541,N_26968,N_26248);
nor U29542 (N_29542,N_27057,N_26619);
xor U29543 (N_29543,N_26554,N_27037);
nor U29544 (N_29544,N_26104,N_27875);
nor U29545 (N_29545,N_26952,N_26939);
or U29546 (N_29546,N_26354,N_27399);
nor U29547 (N_29547,N_26248,N_26950);
nand U29548 (N_29548,N_27443,N_26626);
nor U29549 (N_29549,N_27972,N_26731);
or U29550 (N_29550,N_26365,N_26144);
nand U29551 (N_29551,N_27863,N_26210);
nor U29552 (N_29552,N_26212,N_26913);
nand U29553 (N_29553,N_27210,N_27845);
nand U29554 (N_29554,N_26962,N_26022);
nor U29555 (N_29555,N_27333,N_27399);
or U29556 (N_29556,N_27921,N_26080);
nor U29557 (N_29557,N_27191,N_26479);
nor U29558 (N_29558,N_27631,N_26473);
or U29559 (N_29559,N_27517,N_27717);
nor U29560 (N_29560,N_26999,N_27813);
or U29561 (N_29561,N_27972,N_26554);
or U29562 (N_29562,N_26092,N_27179);
nor U29563 (N_29563,N_27796,N_26031);
nor U29564 (N_29564,N_27539,N_26335);
xor U29565 (N_29565,N_27694,N_26690);
nor U29566 (N_29566,N_27635,N_26798);
nor U29567 (N_29567,N_27206,N_27185);
nor U29568 (N_29568,N_26584,N_26735);
xnor U29569 (N_29569,N_26114,N_26014);
and U29570 (N_29570,N_26543,N_26350);
nand U29571 (N_29571,N_26776,N_27255);
or U29572 (N_29572,N_26375,N_26545);
xor U29573 (N_29573,N_27198,N_27781);
nor U29574 (N_29574,N_26484,N_27457);
or U29575 (N_29575,N_27119,N_27981);
and U29576 (N_29576,N_26604,N_26554);
or U29577 (N_29577,N_26258,N_27099);
or U29578 (N_29578,N_27109,N_26442);
nand U29579 (N_29579,N_27303,N_27771);
and U29580 (N_29580,N_27101,N_27085);
nand U29581 (N_29581,N_26574,N_26998);
and U29582 (N_29582,N_26805,N_27127);
nor U29583 (N_29583,N_27590,N_26683);
nor U29584 (N_29584,N_27531,N_26686);
or U29585 (N_29585,N_27442,N_27359);
or U29586 (N_29586,N_27688,N_27933);
nand U29587 (N_29587,N_26715,N_26311);
xor U29588 (N_29588,N_27231,N_27662);
nand U29589 (N_29589,N_27922,N_27402);
or U29590 (N_29590,N_26651,N_27594);
or U29591 (N_29591,N_26081,N_27375);
nand U29592 (N_29592,N_26103,N_27587);
nor U29593 (N_29593,N_27825,N_27387);
nand U29594 (N_29594,N_27794,N_27204);
or U29595 (N_29595,N_27388,N_27123);
nor U29596 (N_29596,N_27486,N_27205);
nand U29597 (N_29597,N_26817,N_26144);
or U29598 (N_29598,N_26939,N_26692);
xnor U29599 (N_29599,N_27029,N_26719);
and U29600 (N_29600,N_27389,N_27192);
nor U29601 (N_29601,N_27777,N_26422);
nand U29602 (N_29602,N_26165,N_26328);
nand U29603 (N_29603,N_27342,N_26102);
or U29604 (N_29604,N_26099,N_27886);
or U29605 (N_29605,N_26968,N_27680);
and U29606 (N_29606,N_27768,N_27257);
and U29607 (N_29607,N_27046,N_26995);
xor U29608 (N_29608,N_27797,N_27753);
nor U29609 (N_29609,N_26913,N_26078);
xor U29610 (N_29610,N_26012,N_27165);
and U29611 (N_29611,N_26863,N_27480);
nor U29612 (N_29612,N_27166,N_27221);
nor U29613 (N_29613,N_26811,N_27942);
xnor U29614 (N_29614,N_26900,N_27185);
nand U29615 (N_29615,N_27453,N_26027);
xor U29616 (N_29616,N_27091,N_27338);
or U29617 (N_29617,N_26852,N_27242);
and U29618 (N_29618,N_27333,N_27547);
or U29619 (N_29619,N_26235,N_27560);
nor U29620 (N_29620,N_26991,N_27613);
or U29621 (N_29621,N_26555,N_27854);
xor U29622 (N_29622,N_26629,N_27564);
xor U29623 (N_29623,N_26903,N_27965);
nor U29624 (N_29624,N_26645,N_26226);
nor U29625 (N_29625,N_27909,N_27688);
nand U29626 (N_29626,N_26099,N_27671);
nor U29627 (N_29627,N_26133,N_27526);
nor U29628 (N_29628,N_27843,N_26975);
and U29629 (N_29629,N_27557,N_26134);
nor U29630 (N_29630,N_27047,N_26053);
nor U29631 (N_29631,N_27683,N_26912);
xor U29632 (N_29632,N_26065,N_26324);
nor U29633 (N_29633,N_27237,N_27985);
xnor U29634 (N_29634,N_26179,N_26904);
or U29635 (N_29635,N_26570,N_26543);
nor U29636 (N_29636,N_27163,N_27081);
nand U29637 (N_29637,N_27311,N_27321);
xor U29638 (N_29638,N_27436,N_26310);
or U29639 (N_29639,N_27631,N_27017);
or U29640 (N_29640,N_26159,N_27745);
and U29641 (N_29641,N_27251,N_27993);
nand U29642 (N_29642,N_27251,N_26486);
nand U29643 (N_29643,N_26952,N_26742);
and U29644 (N_29644,N_27297,N_26229);
and U29645 (N_29645,N_26527,N_27089);
nor U29646 (N_29646,N_27827,N_27465);
or U29647 (N_29647,N_26579,N_26623);
or U29648 (N_29648,N_27885,N_27451);
xnor U29649 (N_29649,N_27049,N_27354);
xnor U29650 (N_29650,N_27533,N_27365);
nand U29651 (N_29651,N_27956,N_26564);
nand U29652 (N_29652,N_27370,N_26352);
xor U29653 (N_29653,N_27588,N_27546);
or U29654 (N_29654,N_27528,N_26231);
nor U29655 (N_29655,N_26895,N_26935);
or U29656 (N_29656,N_27781,N_26579);
xnor U29657 (N_29657,N_26527,N_26097);
nand U29658 (N_29658,N_27456,N_26034);
nor U29659 (N_29659,N_26338,N_26484);
or U29660 (N_29660,N_26310,N_26804);
and U29661 (N_29661,N_27060,N_27022);
and U29662 (N_29662,N_27011,N_26456);
xnor U29663 (N_29663,N_27323,N_27553);
or U29664 (N_29664,N_26552,N_27020);
nor U29665 (N_29665,N_27030,N_27587);
and U29666 (N_29666,N_27132,N_26694);
xor U29667 (N_29667,N_26763,N_26056);
xor U29668 (N_29668,N_26729,N_27663);
nor U29669 (N_29669,N_27177,N_26981);
xnor U29670 (N_29670,N_26244,N_27856);
nand U29671 (N_29671,N_26869,N_26506);
nand U29672 (N_29672,N_27794,N_26755);
nor U29673 (N_29673,N_27524,N_26400);
or U29674 (N_29674,N_26555,N_26674);
xor U29675 (N_29675,N_26305,N_26952);
xor U29676 (N_29676,N_26032,N_27198);
xnor U29677 (N_29677,N_26656,N_26406);
xor U29678 (N_29678,N_27512,N_27303);
xnor U29679 (N_29679,N_26803,N_26497);
or U29680 (N_29680,N_26862,N_27936);
and U29681 (N_29681,N_26905,N_27048);
nor U29682 (N_29682,N_27540,N_27869);
nand U29683 (N_29683,N_27533,N_27654);
xor U29684 (N_29684,N_26317,N_27033);
nand U29685 (N_29685,N_26931,N_26146);
and U29686 (N_29686,N_26984,N_27943);
and U29687 (N_29687,N_27413,N_26029);
nor U29688 (N_29688,N_27475,N_27673);
or U29689 (N_29689,N_26954,N_27396);
nand U29690 (N_29690,N_27507,N_26375);
or U29691 (N_29691,N_27235,N_27120);
and U29692 (N_29692,N_26008,N_26227);
and U29693 (N_29693,N_27231,N_27270);
xor U29694 (N_29694,N_27545,N_27992);
nand U29695 (N_29695,N_27693,N_26220);
nand U29696 (N_29696,N_27808,N_27888);
nand U29697 (N_29697,N_27004,N_27351);
nand U29698 (N_29698,N_26280,N_27352);
nand U29699 (N_29699,N_27674,N_27817);
nand U29700 (N_29700,N_27916,N_27149);
nor U29701 (N_29701,N_26094,N_26233);
xnor U29702 (N_29702,N_26967,N_27347);
and U29703 (N_29703,N_26394,N_27476);
nand U29704 (N_29704,N_26982,N_27968);
nor U29705 (N_29705,N_26024,N_26265);
nand U29706 (N_29706,N_26727,N_27340);
xnor U29707 (N_29707,N_27458,N_26261);
or U29708 (N_29708,N_27841,N_26454);
xor U29709 (N_29709,N_26136,N_26455);
or U29710 (N_29710,N_26272,N_26868);
xnor U29711 (N_29711,N_26282,N_26671);
xor U29712 (N_29712,N_27103,N_27935);
or U29713 (N_29713,N_27020,N_27967);
and U29714 (N_29714,N_26928,N_27521);
and U29715 (N_29715,N_27349,N_26077);
or U29716 (N_29716,N_26566,N_27326);
and U29717 (N_29717,N_26281,N_27071);
nor U29718 (N_29718,N_27965,N_26917);
xnor U29719 (N_29719,N_27840,N_26160);
nand U29720 (N_29720,N_26479,N_26113);
or U29721 (N_29721,N_27310,N_26467);
and U29722 (N_29722,N_27345,N_26257);
and U29723 (N_29723,N_26454,N_27311);
or U29724 (N_29724,N_26086,N_27198);
xor U29725 (N_29725,N_26813,N_26996);
nor U29726 (N_29726,N_27389,N_27296);
or U29727 (N_29727,N_26807,N_27157);
xnor U29728 (N_29728,N_26796,N_27187);
nand U29729 (N_29729,N_27822,N_27105);
nor U29730 (N_29730,N_26804,N_27735);
nand U29731 (N_29731,N_26836,N_27668);
and U29732 (N_29732,N_26248,N_27011);
or U29733 (N_29733,N_26907,N_26792);
nor U29734 (N_29734,N_27787,N_27395);
nand U29735 (N_29735,N_27444,N_27841);
or U29736 (N_29736,N_27225,N_26974);
nand U29737 (N_29737,N_26755,N_27999);
xor U29738 (N_29738,N_27850,N_27361);
or U29739 (N_29739,N_27428,N_27445);
nand U29740 (N_29740,N_27092,N_27425);
nor U29741 (N_29741,N_27103,N_26884);
nor U29742 (N_29742,N_26237,N_27033);
or U29743 (N_29743,N_27573,N_26194);
xnor U29744 (N_29744,N_26348,N_27655);
nand U29745 (N_29745,N_27526,N_26737);
xnor U29746 (N_29746,N_26273,N_27270);
or U29747 (N_29747,N_26834,N_26714);
nor U29748 (N_29748,N_27469,N_26528);
nand U29749 (N_29749,N_27755,N_26422);
nor U29750 (N_29750,N_27010,N_27218);
nand U29751 (N_29751,N_27932,N_27757);
or U29752 (N_29752,N_26261,N_27022);
or U29753 (N_29753,N_27784,N_26347);
nor U29754 (N_29754,N_27460,N_27316);
and U29755 (N_29755,N_27469,N_26587);
xnor U29756 (N_29756,N_26788,N_27257);
nor U29757 (N_29757,N_27275,N_26018);
nand U29758 (N_29758,N_26296,N_26848);
nand U29759 (N_29759,N_27201,N_27132);
or U29760 (N_29760,N_26598,N_26565);
xnor U29761 (N_29761,N_27808,N_27568);
nand U29762 (N_29762,N_26547,N_27381);
nand U29763 (N_29763,N_26641,N_27678);
nand U29764 (N_29764,N_26254,N_26917);
xnor U29765 (N_29765,N_26142,N_27064);
and U29766 (N_29766,N_26809,N_27792);
or U29767 (N_29767,N_26925,N_26733);
nand U29768 (N_29768,N_27744,N_26342);
or U29769 (N_29769,N_27410,N_27003);
xnor U29770 (N_29770,N_27228,N_26776);
nor U29771 (N_29771,N_27502,N_26913);
nand U29772 (N_29772,N_27601,N_27771);
and U29773 (N_29773,N_27607,N_26903);
nor U29774 (N_29774,N_27509,N_26383);
nor U29775 (N_29775,N_26498,N_26424);
nor U29776 (N_29776,N_26563,N_26342);
xnor U29777 (N_29777,N_26776,N_26312);
nand U29778 (N_29778,N_26192,N_27372);
nand U29779 (N_29779,N_26610,N_27429);
and U29780 (N_29780,N_26379,N_26223);
and U29781 (N_29781,N_27458,N_27446);
xor U29782 (N_29782,N_27452,N_26581);
nand U29783 (N_29783,N_27548,N_26457);
or U29784 (N_29784,N_27763,N_27910);
and U29785 (N_29785,N_27461,N_26434);
nor U29786 (N_29786,N_27774,N_27750);
nor U29787 (N_29787,N_27558,N_27658);
or U29788 (N_29788,N_26689,N_26764);
nor U29789 (N_29789,N_26087,N_27287);
or U29790 (N_29790,N_27486,N_27556);
xor U29791 (N_29791,N_27818,N_27544);
and U29792 (N_29792,N_27632,N_27201);
xor U29793 (N_29793,N_26266,N_26514);
and U29794 (N_29794,N_27760,N_26799);
xor U29795 (N_29795,N_26563,N_27681);
nor U29796 (N_29796,N_27536,N_27136);
and U29797 (N_29797,N_27968,N_26090);
or U29798 (N_29798,N_27802,N_27575);
or U29799 (N_29799,N_27085,N_27095);
nand U29800 (N_29800,N_27638,N_27568);
and U29801 (N_29801,N_27995,N_27960);
and U29802 (N_29802,N_27786,N_27634);
and U29803 (N_29803,N_26795,N_26084);
and U29804 (N_29804,N_27864,N_26134);
xor U29805 (N_29805,N_26743,N_27543);
xor U29806 (N_29806,N_26518,N_27869);
xor U29807 (N_29807,N_26219,N_26175);
and U29808 (N_29808,N_27092,N_27006);
xor U29809 (N_29809,N_27337,N_27367);
and U29810 (N_29810,N_26293,N_27600);
and U29811 (N_29811,N_26249,N_26530);
and U29812 (N_29812,N_27549,N_27907);
nor U29813 (N_29813,N_26487,N_27100);
nor U29814 (N_29814,N_26166,N_26669);
nor U29815 (N_29815,N_27385,N_26469);
nor U29816 (N_29816,N_27459,N_27892);
nand U29817 (N_29817,N_27076,N_27995);
nor U29818 (N_29818,N_27487,N_27870);
nor U29819 (N_29819,N_26251,N_26365);
or U29820 (N_29820,N_27335,N_27264);
or U29821 (N_29821,N_26452,N_26082);
nand U29822 (N_29822,N_27435,N_26427);
xor U29823 (N_29823,N_26976,N_27247);
nand U29824 (N_29824,N_27137,N_26702);
nor U29825 (N_29825,N_27463,N_26055);
nand U29826 (N_29826,N_27164,N_26068);
and U29827 (N_29827,N_27412,N_27553);
and U29828 (N_29828,N_27916,N_27497);
nor U29829 (N_29829,N_27322,N_26048);
nor U29830 (N_29830,N_26612,N_27206);
nor U29831 (N_29831,N_27758,N_26987);
xor U29832 (N_29832,N_26324,N_27564);
nand U29833 (N_29833,N_27956,N_27346);
or U29834 (N_29834,N_26381,N_27773);
and U29835 (N_29835,N_26147,N_26588);
and U29836 (N_29836,N_27699,N_26910);
or U29837 (N_29837,N_26565,N_26514);
nor U29838 (N_29838,N_26649,N_26060);
xnor U29839 (N_29839,N_27864,N_26199);
xor U29840 (N_29840,N_26241,N_26006);
nor U29841 (N_29841,N_27439,N_27976);
xor U29842 (N_29842,N_27770,N_26494);
or U29843 (N_29843,N_27664,N_26296);
nand U29844 (N_29844,N_26382,N_26142);
or U29845 (N_29845,N_27443,N_26445);
xnor U29846 (N_29846,N_27104,N_27025);
nand U29847 (N_29847,N_26878,N_27672);
nand U29848 (N_29848,N_27623,N_27580);
nand U29849 (N_29849,N_27320,N_26343);
nor U29850 (N_29850,N_27358,N_27550);
nand U29851 (N_29851,N_27791,N_26389);
nor U29852 (N_29852,N_27119,N_26604);
xnor U29853 (N_29853,N_27162,N_26384);
nand U29854 (N_29854,N_27505,N_26311);
nor U29855 (N_29855,N_27217,N_27048);
and U29856 (N_29856,N_27600,N_26106);
nor U29857 (N_29857,N_26091,N_27542);
nand U29858 (N_29858,N_26311,N_27788);
and U29859 (N_29859,N_27015,N_26827);
or U29860 (N_29860,N_26390,N_26435);
nor U29861 (N_29861,N_26067,N_27187);
nand U29862 (N_29862,N_26321,N_27730);
and U29863 (N_29863,N_27835,N_26604);
or U29864 (N_29864,N_26382,N_27193);
and U29865 (N_29865,N_27777,N_27469);
or U29866 (N_29866,N_27141,N_27390);
and U29867 (N_29867,N_27380,N_26411);
and U29868 (N_29868,N_27658,N_26593);
and U29869 (N_29869,N_27056,N_27154);
xnor U29870 (N_29870,N_27223,N_27719);
nand U29871 (N_29871,N_27815,N_26023);
xnor U29872 (N_29872,N_26777,N_27937);
or U29873 (N_29873,N_27108,N_27142);
nor U29874 (N_29874,N_26396,N_26167);
nand U29875 (N_29875,N_27761,N_26530);
nand U29876 (N_29876,N_26229,N_27272);
nor U29877 (N_29877,N_26712,N_26076);
and U29878 (N_29878,N_26056,N_26091);
nor U29879 (N_29879,N_26955,N_27872);
and U29880 (N_29880,N_27891,N_27389);
nor U29881 (N_29881,N_26066,N_26105);
nand U29882 (N_29882,N_26782,N_27126);
nor U29883 (N_29883,N_26006,N_27659);
and U29884 (N_29884,N_26068,N_26257);
or U29885 (N_29885,N_26212,N_26040);
or U29886 (N_29886,N_27826,N_26244);
and U29887 (N_29887,N_26006,N_26852);
nor U29888 (N_29888,N_26856,N_26657);
or U29889 (N_29889,N_26314,N_26030);
nor U29890 (N_29890,N_26232,N_26914);
or U29891 (N_29891,N_26649,N_27602);
nand U29892 (N_29892,N_26897,N_27815);
or U29893 (N_29893,N_27074,N_26518);
xor U29894 (N_29894,N_27549,N_27792);
and U29895 (N_29895,N_27482,N_26014);
or U29896 (N_29896,N_26935,N_27648);
nand U29897 (N_29897,N_27835,N_27209);
or U29898 (N_29898,N_27042,N_27808);
and U29899 (N_29899,N_27922,N_26374);
or U29900 (N_29900,N_27684,N_26991);
nand U29901 (N_29901,N_27925,N_27796);
or U29902 (N_29902,N_26512,N_26459);
xor U29903 (N_29903,N_26912,N_26055);
nor U29904 (N_29904,N_26158,N_27517);
nand U29905 (N_29905,N_26194,N_26753);
nand U29906 (N_29906,N_26457,N_26011);
nor U29907 (N_29907,N_26987,N_26474);
xnor U29908 (N_29908,N_27819,N_26375);
nand U29909 (N_29909,N_27298,N_26868);
and U29910 (N_29910,N_27683,N_27410);
nor U29911 (N_29911,N_27838,N_27321);
nor U29912 (N_29912,N_27919,N_26427);
and U29913 (N_29913,N_27876,N_27167);
nor U29914 (N_29914,N_27056,N_27611);
xnor U29915 (N_29915,N_27810,N_27249);
nor U29916 (N_29916,N_26197,N_27249);
xor U29917 (N_29917,N_27475,N_27704);
and U29918 (N_29918,N_26346,N_26213);
nand U29919 (N_29919,N_27344,N_26047);
and U29920 (N_29920,N_27585,N_27320);
nor U29921 (N_29921,N_26920,N_26581);
nand U29922 (N_29922,N_26825,N_26447);
nor U29923 (N_29923,N_26558,N_27163);
nor U29924 (N_29924,N_26604,N_26504);
and U29925 (N_29925,N_27688,N_27456);
or U29926 (N_29926,N_27766,N_27626);
nor U29927 (N_29927,N_26931,N_26278);
nand U29928 (N_29928,N_27003,N_26438);
nor U29929 (N_29929,N_27579,N_27615);
or U29930 (N_29930,N_27762,N_27175);
or U29931 (N_29931,N_26688,N_26514);
nand U29932 (N_29932,N_27887,N_26239);
xnor U29933 (N_29933,N_26320,N_27261);
xor U29934 (N_29934,N_27056,N_26148);
or U29935 (N_29935,N_27757,N_27940);
nand U29936 (N_29936,N_26879,N_27196);
xnor U29937 (N_29937,N_26098,N_26134);
xnor U29938 (N_29938,N_26847,N_26772);
xor U29939 (N_29939,N_26164,N_27473);
nor U29940 (N_29940,N_27995,N_27991);
or U29941 (N_29941,N_27269,N_26796);
nand U29942 (N_29942,N_26932,N_26269);
nand U29943 (N_29943,N_27975,N_26852);
nor U29944 (N_29944,N_26714,N_26985);
xor U29945 (N_29945,N_27604,N_27098);
xor U29946 (N_29946,N_27632,N_26636);
or U29947 (N_29947,N_27300,N_26459);
nor U29948 (N_29948,N_26418,N_26986);
nand U29949 (N_29949,N_26711,N_26780);
or U29950 (N_29950,N_27226,N_27806);
xor U29951 (N_29951,N_26227,N_26796);
and U29952 (N_29952,N_27880,N_26315);
xnor U29953 (N_29953,N_26644,N_26346);
or U29954 (N_29954,N_26223,N_26279);
or U29955 (N_29955,N_26183,N_27829);
or U29956 (N_29956,N_27830,N_27511);
and U29957 (N_29957,N_27979,N_26148);
and U29958 (N_29958,N_27535,N_27659);
nand U29959 (N_29959,N_26070,N_26298);
and U29960 (N_29960,N_26088,N_26844);
nor U29961 (N_29961,N_26044,N_26840);
and U29962 (N_29962,N_27733,N_26317);
xor U29963 (N_29963,N_27299,N_27054);
and U29964 (N_29964,N_27667,N_26101);
and U29965 (N_29965,N_26151,N_26126);
nor U29966 (N_29966,N_26261,N_27754);
xnor U29967 (N_29967,N_27084,N_27767);
nor U29968 (N_29968,N_26202,N_27034);
or U29969 (N_29969,N_27105,N_26728);
nand U29970 (N_29970,N_26393,N_26161);
or U29971 (N_29971,N_27279,N_26238);
or U29972 (N_29972,N_27223,N_27198);
or U29973 (N_29973,N_27347,N_26617);
xor U29974 (N_29974,N_26233,N_27107);
and U29975 (N_29975,N_27416,N_26979);
or U29976 (N_29976,N_27035,N_26127);
xor U29977 (N_29977,N_26733,N_26778);
and U29978 (N_29978,N_26875,N_27057);
and U29979 (N_29979,N_26938,N_27621);
nand U29980 (N_29980,N_27593,N_26934);
nand U29981 (N_29981,N_26157,N_26491);
nand U29982 (N_29982,N_26355,N_27159);
and U29983 (N_29983,N_27860,N_27494);
xnor U29984 (N_29984,N_26677,N_27723);
or U29985 (N_29985,N_26824,N_26346);
and U29986 (N_29986,N_27712,N_26228);
nand U29987 (N_29987,N_27223,N_26071);
or U29988 (N_29988,N_26887,N_27201);
xor U29989 (N_29989,N_27962,N_26707);
nand U29990 (N_29990,N_26958,N_27040);
nand U29991 (N_29991,N_26722,N_26650);
nor U29992 (N_29992,N_27569,N_26997);
and U29993 (N_29993,N_26089,N_27962);
nand U29994 (N_29994,N_26482,N_27484);
nor U29995 (N_29995,N_27500,N_26346);
or U29996 (N_29996,N_27810,N_26439);
or U29997 (N_29997,N_27353,N_27964);
or U29998 (N_29998,N_27707,N_26827);
and U29999 (N_29999,N_27588,N_27879);
xor U30000 (N_30000,N_28135,N_28825);
or U30001 (N_30001,N_29969,N_29542);
nor U30002 (N_30002,N_28468,N_28762);
nand U30003 (N_30003,N_29663,N_29816);
nand U30004 (N_30004,N_28738,N_28037);
xnor U30005 (N_30005,N_29831,N_29734);
nor U30006 (N_30006,N_28808,N_29789);
nor U30007 (N_30007,N_28000,N_29437);
nor U30008 (N_30008,N_28906,N_29088);
xor U30009 (N_30009,N_29333,N_29533);
xnor U30010 (N_30010,N_29003,N_28731);
xnor U30011 (N_30011,N_28050,N_28043);
nor U30012 (N_30012,N_29595,N_29892);
or U30013 (N_30013,N_29729,N_28301);
nor U30014 (N_30014,N_28939,N_28042);
and U30015 (N_30015,N_29900,N_29047);
and U30016 (N_30016,N_29091,N_28976);
xnor U30017 (N_30017,N_28572,N_28790);
or U30018 (N_30018,N_28706,N_28845);
nand U30019 (N_30019,N_29021,N_29246);
or U30020 (N_30020,N_28036,N_29097);
and U30021 (N_30021,N_29929,N_29353);
or U30022 (N_30022,N_29356,N_29588);
xnor U30023 (N_30023,N_28151,N_28996);
xnor U30024 (N_30024,N_29584,N_28127);
nand U30025 (N_30025,N_29976,N_29611);
or U30026 (N_30026,N_29064,N_28575);
nor U30027 (N_30027,N_28262,N_28697);
or U30028 (N_30028,N_28792,N_29369);
or U30029 (N_30029,N_28723,N_29518);
nand U30030 (N_30030,N_28476,N_29860);
nand U30031 (N_30031,N_28435,N_29251);
nor U30032 (N_30032,N_28561,N_29308);
or U30033 (N_30033,N_28531,N_29548);
xor U30034 (N_30034,N_29701,N_28394);
nor U30035 (N_30035,N_29494,N_29104);
or U30036 (N_30036,N_28388,N_29079);
xor U30037 (N_30037,N_28479,N_28728);
nand U30038 (N_30038,N_28876,N_29309);
xor U30039 (N_30039,N_29297,N_28196);
nor U30040 (N_30040,N_28497,N_29268);
nor U30041 (N_30041,N_29972,N_29373);
nor U30042 (N_30042,N_29001,N_28460);
or U30043 (N_30043,N_28713,N_29241);
xnor U30044 (N_30044,N_29887,N_29193);
or U30045 (N_30045,N_29582,N_28039);
and U30046 (N_30046,N_29429,N_28611);
nor U30047 (N_30047,N_29675,N_28137);
nand U30048 (N_30048,N_28250,N_28844);
nor U30049 (N_30049,N_28401,N_28954);
or U30050 (N_30050,N_29067,N_29525);
nor U30051 (N_30051,N_28699,N_28072);
nor U30052 (N_30052,N_28437,N_28383);
or U30053 (N_30053,N_29866,N_28364);
nor U30054 (N_30054,N_28970,N_29726);
and U30055 (N_30055,N_29817,N_28889);
or U30056 (N_30056,N_28756,N_29819);
and U30057 (N_30057,N_28136,N_29211);
nand U30058 (N_30058,N_28170,N_29813);
nand U30059 (N_30059,N_29412,N_29823);
xnor U30060 (N_30060,N_29747,N_28812);
nor U30061 (N_30061,N_29068,N_29247);
xnor U30062 (N_30062,N_28667,N_29295);
or U30063 (N_30063,N_28570,N_29253);
xor U30064 (N_30064,N_28701,N_29826);
or U30065 (N_30065,N_29464,N_29618);
nor U30066 (N_30066,N_28244,N_28436);
xor U30067 (N_30067,N_29000,N_29706);
nor U30068 (N_30068,N_28556,N_28909);
and U30069 (N_30069,N_29818,N_29554);
xor U30070 (N_30070,N_28576,N_29366);
and U30071 (N_30071,N_29620,N_29481);
nand U30072 (N_30072,N_28323,N_28004);
and U30073 (N_30073,N_28217,N_28178);
xor U30074 (N_30074,N_29472,N_28732);
nand U30075 (N_30075,N_29009,N_28271);
xor U30076 (N_30076,N_29199,N_28514);
and U30077 (N_30077,N_28222,N_29705);
and U30078 (N_30078,N_28141,N_29514);
nand U30079 (N_30079,N_28492,N_29797);
or U30080 (N_30080,N_28333,N_28986);
and U30081 (N_30081,N_29229,N_29863);
nor U30082 (N_30082,N_29617,N_28863);
nand U30083 (N_30083,N_29640,N_29678);
or U30084 (N_30084,N_28221,N_29111);
nand U30085 (N_30085,N_29650,N_29249);
xor U30086 (N_30086,N_28098,N_28409);
nand U30087 (N_30087,N_29228,N_29758);
or U30088 (N_30088,N_29551,N_28983);
and U30089 (N_30089,N_28289,N_28320);
nand U30090 (N_30090,N_28950,N_28851);
nand U30091 (N_30091,N_29383,N_28559);
xor U30092 (N_30092,N_28107,N_28972);
xnor U30093 (N_30093,N_29793,N_29530);
or U30094 (N_30094,N_29184,N_28060);
or U30095 (N_30095,N_29360,N_29165);
nand U30096 (N_30096,N_28375,N_28524);
nand U30097 (N_30097,N_29547,N_29778);
and U30098 (N_30098,N_29833,N_29851);
and U30099 (N_30099,N_29973,N_28140);
nor U30100 (N_30100,N_28429,N_28430);
or U30101 (N_30101,N_29766,N_28526);
xor U30102 (N_30102,N_28233,N_28786);
nand U30103 (N_30103,N_29460,N_29508);
or U30104 (N_30104,N_28758,N_28617);
xor U30105 (N_30105,N_28980,N_28771);
and U30106 (N_30106,N_28454,N_29462);
nand U30107 (N_30107,N_28515,N_28405);
nand U30108 (N_30108,N_29754,N_29779);
or U30109 (N_30109,N_28630,N_29132);
and U30110 (N_30110,N_28999,N_29915);
xor U30111 (N_30111,N_29441,N_29343);
or U30112 (N_30112,N_28255,N_29536);
and U30113 (N_30113,N_28188,N_29970);
xor U30114 (N_30114,N_28900,N_28563);
nand U30115 (N_30115,N_28940,N_29114);
or U30116 (N_30116,N_28836,N_28849);
xor U30117 (N_30117,N_28331,N_28292);
or U30118 (N_30118,N_29160,N_29210);
nand U30119 (N_30119,N_28165,N_28560);
xor U30120 (N_30120,N_29157,N_29265);
or U30121 (N_30121,N_28294,N_28604);
xor U30122 (N_30122,N_29733,N_29313);
nor U30123 (N_30123,N_28215,N_28833);
nor U30124 (N_30124,N_28595,N_28607);
nand U30125 (N_30125,N_28696,N_29528);
nand U30126 (N_30126,N_29662,N_28206);
or U30127 (N_30127,N_29304,N_29188);
nand U30128 (N_30128,N_29987,N_28658);
and U30129 (N_30129,N_28312,N_29834);
nand U30130 (N_30130,N_28382,N_28615);
nand U30131 (N_30131,N_29093,N_29478);
xnor U30132 (N_30132,N_28419,N_28627);
nand U30133 (N_30133,N_29459,N_29415);
xor U30134 (N_30134,N_28266,N_29155);
nor U30135 (N_30135,N_28772,N_29034);
nand U30136 (N_30136,N_28788,N_28660);
and U30137 (N_30137,N_28315,N_28452);
nor U30138 (N_30138,N_28358,N_28190);
and U30139 (N_30139,N_28534,N_28548);
nor U30140 (N_30140,N_28525,N_28003);
or U30141 (N_30141,N_29107,N_28528);
nand U30142 (N_30142,N_28277,N_29074);
xor U30143 (N_30143,N_29896,N_29127);
and U30144 (N_30144,N_28730,N_29612);
nand U30145 (N_30145,N_28057,N_29116);
nor U30146 (N_30146,N_28441,N_28782);
nor U30147 (N_30147,N_28979,N_29479);
xnor U30148 (N_30148,N_28487,N_29868);
nand U30149 (N_30149,N_28432,N_28574);
nor U30150 (N_30150,N_28086,N_28481);
nor U30151 (N_30151,N_29142,N_29041);
nor U30152 (N_30152,N_29982,N_28894);
or U30153 (N_30153,N_28353,N_29578);
nor U30154 (N_30154,N_29967,N_28915);
nand U30155 (N_30155,N_28582,N_29538);
and U30156 (N_30156,N_29621,N_28332);
nor U30157 (N_30157,N_29714,N_29349);
nand U30158 (N_30158,N_29002,N_29205);
or U30159 (N_30159,N_29845,N_28775);
nand U30160 (N_30160,N_29657,N_28577);
or U30161 (N_30161,N_29431,N_29444);
nand U30162 (N_30162,N_28020,N_28944);
nand U30163 (N_30163,N_28112,N_29791);
nor U30164 (N_30164,N_28819,N_29432);
xnor U30165 (N_30165,N_28977,N_28109);
or U30166 (N_30166,N_28070,N_28916);
nor U30167 (N_30167,N_29944,N_29109);
xnor U30168 (N_30168,N_29893,N_28108);
and U30169 (N_30169,N_28032,N_29317);
or U30170 (N_30170,N_28523,N_28789);
xor U30171 (N_30171,N_29261,N_28583);
and U30172 (N_30172,N_28114,N_28911);
nor U30173 (N_30173,N_29568,N_28091);
or U30174 (N_30174,N_29121,N_28877);
nand U30175 (N_30175,N_29722,N_28022);
or U30176 (N_30176,N_28761,N_28488);
nor U30177 (N_30177,N_28268,N_28500);
xor U30178 (N_30178,N_28148,N_28647);
nor U30179 (N_30179,N_29052,N_29457);
nor U30180 (N_30180,N_29832,N_28182);
or U30181 (N_30181,N_29335,N_28021);
nand U30182 (N_30182,N_29581,N_28903);
xor U30183 (N_30183,N_28156,N_29045);
or U30184 (N_30184,N_28638,N_29553);
nor U30185 (N_30185,N_29785,N_29103);
or U30186 (N_30186,N_28711,N_28748);
nor U30187 (N_30187,N_29753,N_28425);
nor U30188 (N_30188,N_29144,N_28663);
xnor U30189 (N_30189,N_29952,N_29909);
xor U30190 (N_30190,N_28550,N_28882);
xor U30191 (N_30191,N_28062,N_29783);
nor U30192 (N_30192,N_28123,N_29661);
nor U30193 (N_30193,N_28593,N_28739);
xnor U30194 (N_30194,N_28517,N_29639);
nand U30195 (N_30195,N_28279,N_28662);
or U30196 (N_30196,N_29985,N_29348);
and U30197 (N_30197,N_29852,N_28875);
nor U30198 (N_30198,N_29961,N_28442);
nand U30199 (N_30199,N_29713,N_28200);
or U30200 (N_30200,N_28824,N_29280);
or U30201 (N_30201,N_29135,N_28404);
and U30202 (N_30202,N_28989,N_29399);
xnor U30203 (N_30203,N_28703,N_28120);
nand U30204 (N_30204,N_29314,N_29943);
nor U30205 (N_30205,N_28951,N_29438);
or U30206 (N_30206,N_28619,N_28634);
nand U30207 (N_30207,N_29959,N_28931);
nor U30208 (N_30208,N_29040,N_29587);
nand U30209 (N_30209,N_29322,N_28334);
nand U30210 (N_30210,N_29759,N_29435);
or U30211 (N_30211,N_29699,N_29709);
nand U30212 (N_30212,N_29926,N_28205);
nand U30213 (N_30213,N_29539,N_28313);
nand U30214 (N_30214,N_28859,N_28229);
xor U30215 (N_30215,N_28439,N_28541);
xnor U30216 (N_30216,N_29798,N_29393);
nand U30217 (N_30217,N_28457,N_28890);
nor U30218 (N_30218,N_29505,N_28985);
nand U30219 (N_30219,N_29487,N_29396);
nor U30220 (N_30220,N_28848,N_29351);
and U30221 (N_30221,N_29978,N_28935);
or U30222 (N_30222,N_29767,N_29048);
nor U30223 (N_30223,N_29061,N_29183);
and U30224 (N_30224,N_29167,N_28483);
xor U30225 (N_30225,N_28818,N_28930);
nand U30226 (N_30226,N_28672,N_29880);
xor U30227 (N_30227,N_29381,N_28892);
or U30228 (N_30228,N_28866,N_29019);
or U30229 (N_30229,N_29574,N_29993);
xor U30230 (N_30230,N_28132,N_28183);
xnor U30231 (N_30231,N_28234,N_28506);
nor U30232 (N_30232,N_29565,N_29989);
and U30233 (N_30233,N_29654,N_28090);
and U30234 (N_30234,N_28318,N_28321);
or U30235 (N_30235,N_29932,N_28444);
nor U30236 (N_30236,N_29287,N_28549);
xor U30237 (N_30237,N_29524,N_28805);
xor U30238 (N_30238,N_28379,N_28048);
nor U30239 (N_30239,N_29147,N_28800);
and U30240 (N_30240,N_29452,N_28092);
nor U30241 (N_30241,N_29060,N_28041);
xnor U30242 (N_30242,N_28263,N_29179);
nand U30243 (N_30243,N_28324,N_29476);
or U30244 (N_30244,N_28464,N_29468);
nand U30245 (N_30245,N_28811,N_29303);
nor U30246 (N_30246,N_28657,N_29728);
and U30247 (N_30247,N_29497,N_29750);
or U30248 (N_30248,N_28180,N_29503);
or U30249 (N_30249,N_28414,N_29471);
and U30250 (N_30250,N_29599,N_28480);
or U30251 (N_30251,N_29672,N_29787);
xor U30252 (N_30252,N_28714,N_29695);
or U30253 (N_30253,N_28609,N_29903);
nand U30254 (N_30254,N_28540,N_29928);
nor U30255 (N_30255,N_28769,N_28678);
or U30256 (N_30256,N_29202,N_29004);
nand U30257 (N_30257,N_29800,N_29828);
nand U30258 (N_30258,N_28498,N_28538);
or U30259 (N_30259,N_29844,N_29178);
and U30260 (N_30260,N_28878,N_28766);
or U30261 (N_30261,N_29875,N_28695);
nand U30262 (N_30262,N_29286,N_28285);
and U30263 (N_30263,N_29367,N_29421);
or U30264 (N_30264,N_28264,N_29024);
or U30265 (N_30265,N_29240,N_29516);
nand U30266 (N_30266,N_29693,N_29365);
and U30267 (N_30267,N_29401,N_29564);
xnor U30268 (N_30268,N_28343,N_29613);
and U30269 (N_30269,N_28934,N_29513);
nor U30270 (N_30270,N_29424,N_28505);
nor U30271 (N_30271,N_28445,N_29090);
nand U30272 (N_30272,N_29131,N_28208);
xnor U30273 (N_30273,N_28623,N_28291);
nand U30274 (N_30274,N_28671,N_28161);
nor U30275 (N_30275,N_29520,N_28040);
xnor U30276 (N_30276,N_28997,N_28245);
and U30277 (N_30277,N_29310,N_29260);
nand U30278 (N_30278,N_29129,N_28650);
and U30279 (N_30279,N_28385,N_29329);
xor U30280 (N_30280,N_28850,N_29942);
or U30281 (N_30281,N_28616,N_29688);
nor U30282 (N_30282,N_28910,N_29814);
xor U30283 (N_30283,N_29130,N_28880);
or U30284 (N_30284,N_28362,N_28661);
and U30285 (N_30285,N_29630,N_28629);
nand U30286 (N_30286,N_28261,N_28296);
nand U30287 (N_30287,N_29106,N_29252);
or U30288 (N_30288,N_29710,N_29277);
nand U30289 (N_30289,N_28557,N_28917);
nand U30290 (N_30290,N_28924,N_29032);
nand U30291 (N_30291,N_28297,N_29300);
nor U30292 (N_30292,N_29406,N_29043);
xor U30293 (N_30293,N_28053,N_28644);
nand U30294 (N_30294,N_28547,N_29737);
and U30295 (N_30295,N_28104,N_28026);
or U30296 (N_30296,N_28093,N_28155);
xor U30297 (N_30297,N_29124,N_29938);
or U30298 (N_30298,N_29874,N_28945);
nor U30299 (N_30299,N_29491,N_28648);
nor U30300 (N_30300,N_29180,N_29891);
and U30301 (N_30301,N_29752,N_29363);
or U30302 (N_30302,N_28864,N_29133);
and U30303 (N_30303,N_29123,N_28729);
nand U30304 (N_30304,N_29203,N_28814);
nor U30305 (N_30305,N_28520,N_29311);
and U30306 (N_30306,N_29307,N_29148);
or U30307 (N_30307,N_29143,N_29719);
nor U30308 (N_30308,N_28248,N_29974);
and U30309 (N_30309,N_29625,N_29404);
xnor U30310 (N_30310,N_29770,N_29259);
nand U30311 (N_30311,N_29506,N_28794);
xor U30312 (N_30312,N_28288,N_28928);
nand U30313 (N_30313,N_28975,N_28219);
xnor U30314 (N_30314,N_29062,N_28791);
nor U30315 (N_30315,N_28254,N_29628);
nor U30316 (N_30316,N_28386,N_28339);
xnor U30317 (N_30317,N_28453,N_29145);
nand U30318 (N_30318,N_28393,N_29339);
nand U30319 (N_30319,N_28100,N_29677);
nor U30320 (N_30320,N_29664,N_28283);
nor U30321 (N_30321,N_28016,N_28943);
or U30322 (N_30322,N_28501,N_28069);
or U30323 (N_30323,N_28533,N_28965);
or U30324 (N_30324,N_29741,N_28166);
nor U30325 (N_30325,N_28688,N_28816);
or U30326 (N_30326,N_29897,N_28482);
and U30327 (N_30327,N_28763,N_29039);
nor U30328 (N_30328,N_28002,N_29667);
nand U30329 (N_30329,N_29856,N_29603);
nor U30330 (N_30330,N_29805,N_28591);
nand U30331 (N_30331,N_29126,N_28067);
and U30332 (N_30332,N_28636,N_28061);
xor U30333 (N_30333,N_28753,N_28223);
xor U30334 (N_30334,N_28680,N_29683);
and U30335 (N_30335,N_28073,N_29331);
nand U30336 (N_30336,N_29291,N_28126);
and U30337 (N_30337,N_28959,N_29388);
nand U30338 (N_30338,N_29531,N_28612);
nand U30339 (N_30339,N_28396,N_29271);
nand U30340 (N_30340,N_28105,N_28011);
nor U30341 (N_30341,N_28051,N_29669);
and U30342 (N_30342,N_29274,N_29724);
nor U30343 (N_30343,N_29453,N_28172);
or U30344 (N_30344,N_29712,N_29500);
and U30345 (N_30345,N_29950,N_28010);
xor U30346 (N_30346,N_29872,N_29011);
nor U30347 (N_30347,N_29092,N_29390);
xnor U30348 (N_30348,N_29725,N_29195);
nand U30349 (N_30349,N_29792,N_29532);
and U30350 (N_30350,N_28955,N_29031);
xor U30351 (N_30351,N_28743,N_29208);
and U30352 (N_30352,N_28345,N_28806);
nor U30353 (N_30353,N_29507,N_28082);
and U30354 (N_30354,N_29445,N_28922);
or U30355 (N_30355,N_29643,N_29594);
xor U30356 (N_30356,N_28799,N_29642);
nand U30357 (N_30357,N_28737,N_29134);
nor U30358 (N_30358,N_29219,N_28717);
and U30359 (N_30359,N_28191,N_28220);
xnor U30360 (N_30360,N_29495,N_29761);
xnor U30361 (N_30361,N_28031,N_28046);
nand U30362 (N_30362,N_28326,N_28484);
and U30363 (N_30363,N_28101,N_29477);
and U30364 (N_30364,N_29344,N_29008);
nand U30365 (N_30365,N_28529,N_29250);
nor U30366 (N_30366,N_28478,N_28840);
nor U30367 (N_30367,N_29924,N_29358);
or U30368 (N_30368,N_28342,N_29112);
and U30369 (N_30369,N_28238,N_28752);
xor U30370 (N_30370,N_28237,N_28747);
xnor U30371 (N_30371,N_28586,N_28189);
nand U30372 (N_30372,N_29440,N_29673);
or U30373 (N_30373,N_28974,N_29150);
and U30374 (N_30374,N_29325,N_28578);
nand U30375 (N_30375,N_29086,N_28162);
nand U30376 (N_30376,N_28597,N_28727);
xor U30377 (N_30377,N_28804,N_29244);
nor U30378 (N_30378,N_29912,N_29028);
nor U30379 (N_30379,N_29336,N_29474);
nand U30380 (N_30380,N_28870,N_29151);
xor U30381 (N_30381,N_29023,N_29540);
nor U30382 (N_30382,N_28272,N_29634);
nor U30383 (N_30383,N_28443,N_28054);
xor U30384 (N_30384,N_29402,N_29117);
and U30385 (N_30385,N_28646,N_28639);
xor U30386 (N_30386,N_29806,N_28914);
or U30387 (N_30387,N_28477,N_28322);
and U30388 (N_30388,N_28742,N_29602);
and U30389 (N_30389,N_28253,N_28145);
nand U30390 (N_30390,N_29649,N_29377);
and U30391 (N_30391,N_28749,N_28169);
nand U30392 (N_30392,N_28904,N_29095);
nand U30393 (N_30393,N_28372,N_28265);
xnor U30394 (N_30394,N_29347,N_28925);
nor U30395 (N_30395,N_29227,N_29659);
or U30396 (N_30396,N_29871,N_28902);
xnor U30397 (N_30397,N_29201,N_28079);
and U30398 (N_30398,N_28417,N_29839);
or U30399 (N_30399,N_29955,N_29689);
nor U30400 (N_30400,N_28198,N_28088);
nand U30401 (N_30401,N_28679,N_28508);
and U30402 (N_30402,N_28495,N_29881);
nand U30403 (N_30403,N_29768,N_29991);
or U30404 (N_30404,N_29939,N_29038);
or U30405 (N_30405,N_28767,N_28179);
xnor U30406 (N_30406,N_29030,N_28868);
and U30407 (N_30407,N_28821,N_28670);
xnor U30408 (N_30408,N_29555,N_28510);
nor U30409 (N_30409,N_28489,N_28361);
nor U30410 (N_30410,N_28602,N_29204);
nor U30411 (N_30411,N_28837,N_28905);
or U30412 (N_30412,N_28350,N_29980);
xor U30413 (N_30413,N_29425,N_29315);
xor U30414 (N_30414,N_28034,N_29416);
nand U30415 (N_30415,N_28736,N_28280);
xor U30416 (N_30416,N_28891,N_29511);
or U30417 (N_30417,N_28075,N_28869);
or U30418 (N_30418,N_29808,N_29215);
and U30419 (N_30419,N_29906,N_28349);
xnor U30420 (N_30420,N_28408,N_28142);
nand U30421 (N_30421,N_29931,N_29306);
or U30422 (N_30422,N_28527,N_28551);
and U30423 (N_30423,N_29189,N_28860);
or U30424 (N_30424,N_28596,N_28111);
nor U30425 (N_30425,N_29849,N_28337);
nor U30426 (N_30426,N_29563,N_28449);
xor U30427 (N_30427,N_29138,N_29707);
and U30428 (N_30428,N_28485,N_29862);
nand U30429 (N_30429,N_28684,N_29380);
or U30430 (N_30430,N_29697,N_28210);
or U30431 (N_30431,N_29036,N_28635);
or U30432 (N_30432,N_29262,N_29746);
or U30433 (N_30433,N_28676,N_29898);
nor U30434 (N_30434,N_29301,N_28949);
nand U30435 (N_30435,N_28918,N_29458);
nor U30436 (N_30436,N_28553,N_28017);
nor U30437 (N_30437,N_28018,N_28403);
or U30438 (N_30438,N_29499,N_28038);
or U30439 (N_30439,N_28700,N_28565);
xor U30440 (N_30440,N_29063,N_28793);
or U30441 (N_30441,N_29788,N_29690);
nor U30442 (N_30442,N_28956,N_28094);
and U30443 (N_30443,N_28099,N_29171);
or U30444 (N_30444,N_29796,N_28608);
nor U30445 (N_30445,N_29484,N_28276);
or U30446 (N_30446,N_29560,N_29933);
or U30447 (N_30447,N_29051,N_28991);
xor U30448 (N_30448,N_29914,N_29586);
xor U30449 (N_30449,N_29146,N_29279);
nor U30450 (N_30450,N_28692,N_28998);
xnor U30451 (N_30451,N_28458,N_29427);
or U30452 (N_30452,N_29159,N_29368);
xor U30453 (N_30453,N_28751,N_29609);
nand U30454 (N_30454,N_29886,N_29098);
xnor U30455 (N_30455,N_28144,N_28197);
nor U30456 (N_30456,N_29527,N_28465);
xnor U30457 (N_30457,N_29233,N_29526);
nand U30458 (N_30458,N_28058,N_29988);
xnor U30459 (N_30459,N_29883,N_29825);
and U30460 (N_30460,N_28774,N_28886);
nand U30461 (N_30461,N_28704,N_29781);
xnor U30462 (N_30462,N_28542,N_29237);
nor U30463 (N_30463,N_29815,N_29632);
and U30464 (N_30464,N_28118,N_28216);
nor U30465 (N_30465,N_28456,N_29018);
nand U30466 (N_30466,N_28269,N_29771);
nand U30467 (N_30467,N_28502,N_29731);
nor U30468 (N_30468,N_28371,N_29601);
and U30469 (N_30469,N_29120,N_29850);
or U30470 (N_30470,N_29730,N_28948);
nand U30471 (N_30471,N_28537,N_29854);
nor U30472 (N_30472,N_28626,N_29890);
or U30473 (N_30473,N_28392,N_28171);
xor U30474 (N_30474,N_29057,N_29055);
nand U30475 (N_30475,N_28947,N_29073);
or U30476 (N_30476,N_29723,N_28116);
xor U30477 (N_30477,N_29164,N_29760);
nor U30478 (N_30478,N_28938,N_29836);
or U30479 (N_30479,N_29122,N_29812);
nand U30480 (N_30480,N_29273,N_28256);
or U30481 (N_30481,N_29082,N_28400);
or U30482 (N_30482,N_29266,N_29575);
or U30483 (N_30483,N_29359,N_29512);
and U30484 (N_30484,N_28781,N_29059);
or U30485 (N_30485,N_28096,N_29894);
and U30486 (N_30486,N_29930,N_28828);
or U30487 (N_30487,N_29469,N_29345);
nand U30488 (N_30488,N_28843,N_29293);
xor U30489 (N_30489,N_28852,N_29908);
nor U30490 (N_30490,N_28211,N_28839);
nand U30491 (N_30491,N_28830,N_28427);
xor U30492 (N_30492,N_29434,N_28275);
xor U30493 (N_30493,N_28967,N_28387);
or U30494 (N_30494,N_28490,N_28901);
nand U30495 (N_30495,N_29409,N_28601);
or U30496 (N_30496,N_29680,N_28600);
nor U30497 (N_30497,N_29362,N_28076);
xor U30498 (N_30498,N_29700,N_28919);
xnor U30499 (N_30499,N_29224,N_29614);
xnor U30500 (N_30500,N_29414,N_28095);
or U30501 (N_30501,N_28055,N_28598);
nand U30502 (N_30502,N_28606,N_28327);
and U30503 (N_30503,N_28785,N_29966);
xnor U30504 (N_30504,N_29696,N_28491);
nand U30505 (N_30505,N_28426,N_28305);
or U30506 (N_30506,N_29181,N_29997);
and U30507 (N_30507,N_28235,N_28573);
and U30508 (N_30508,N_29113,N_28984);
or U30509 (N_30509,N_29960,N_28066);
or U30510 (N_30510,N_28757,N_28359);
or U30511 (N_30511,N_28357,N_28065);
nor U30512 (N_30512,N_29156,N_29276);
xor U30513 (N_30513,N_28666,N_28252);
nor U30514 (N_30514,N_28153,N_28963);
nand U30515 (N_30515,N_29275,N_29557);
nor U30516 (N_30516,N_29270,N_28314);
and U30517 (N_30517,N_28173,N_29426);
or U30518 (N_30518,N_29666,N_29708);
nand U30519 (N_30519,N_29190,N_28539);
or U30520 (N_30520,N_29014,N_29676);
or U30521 (N_30521,N_29604,N_29196);
nand U30522 (N_30522,N_28351,N_29254);
nor U30523 (N_30523,N_29902,N_28071);
and U30524 (N_30524,N_28415,N_28689);
and U30525 (N_30525,N_28873,N_29990);
nor U30526 (N_30526,N_29537,N_28440);
nor U30527 (N_30527,N_29589,N_28926);
nand U30528 (N_30528,N_29174,N_28341);
or U30529 (N_30529,N_28360,N_28290);
and U30530 (N_30530,N_29436,N_28854);
nand U30531 (N_30531,N_29005,N_29278);
and U30532 (N_30532,N_29840,N_29069);
xnor U30533 (N_30533,N_29879,N_29027);
nor U30534 (N_30534,N_29361,N_29646);
nor U30535 (N_30535,N_28923,N_29411);
xor U30536 (N_30536,N_28078,N_28446);
or U30537 (N_30537,N_29099,N_29364);
nand U30538 (N_30538,N_28961,N_28257);
nand U30539 (N_30539,N_29139,N_29670);
nand U30540 (N_30540,N_28705,N_29718);
xnor U30541 (N_30541,N_29428,N_29544);
nor U30542 (N_30542,N_28555,N_28605);
or U30543 (N_30543,N_28397,N_28081);
and U30544 (N_30544,N_29408,N_29608);
or U30545 (N_30545,N_29681,N_28740);
or U30546 (N_30546,N_29992,N_28656);
and U30547 (N_30547,N_29848,N_28942);
or U30548 (N_30548,N_28579,N_28434);
and U30549 (N_30549,N_29161,N_29166);
nor U30550 (N_30550,N_28669,N_28047);
or U30551 (N_30551,N_28585,N_28494);
or U30552 (N_30552,N_29627,N_29936);
nor U30553 (N_30553,N_28175,N_29651);
nor U30554 (N_30554,N_28817,N_28325);
xor U30555 (N_30555,N_29698,N_29635);
nand U30556 (N_30556,N_29025,N_29316);
and U30557 (N_30557,N_29801,N_28499);
nand U30558 (N_30558,N_29644,N_29763);
nand U30559 (N_30559,N_28131,N_28893);
nor U30560 (N_30560,N_29945,N_28815);
and U30561 (N_30561,N_29328,N_28512);
and U30562 (N_30562,N_29837,N_29515);
nand U30563 (N_30563,N_28776,N_28129);
nand U30564 (N_30564,N_29288,N_29764);
and U30565 (N_30565,N_28193,N_28779);
and U30566 (N_30566,N_29149,N_28455);
nor U30567 (N_30567,N_28496,N_28157);
nand U30568 (N_30568,N_28770,N_29501);
nor U30569 (N_30569,N_28795,N_29720);
nand U30570 (N_30570,N_28281,N_28374);
and U30571 (N_30571,N_29182,N_29289);
and U30572 (N_30572,N_28725,N_28063);
nor U30573 (N_30573,N_29577,N_28895);
or U30574 (N_30574,N_29403,N_29294);
and U30575 (N_30575,N_28160,N_28568);
and U30576 (N_30576,N_29566,N_29389);
nand U30577 (N_30577,N_29355,N_28421);
xnor U30578 (N_30578,N_29692,N_29986);
xnor U30579 (N_30579,N_28710,N_29543);
nand U30580 (N_30580,N_28012,N_28412);
or U30581 (N_30581,N_29169,N_29264);
nand U30582 (N_30582,N_29226,N_28543);
and U30583 (N_30583,N_29492,N_29841);
or U30584 (N_30584,N_29964,N_29979);
xor U30585 (N_30585,N_28231,N_29026);
nand U30586 (N_30586,N_28773,N_28686);
xor U30587 (N_30587,N_28832,N_28898);
or U30588 (N_30588,N_28355,N_29077);
and U30589 (N_30589,N_28293,N_28665);
nor U30590 (N_30590,N_29765,N_28259);
or U30591 (N_30591,N_28513,N_29999);
nand U30592 (N_30592,N_29864,N_28855);
nor U30593 (N_30593,N_29509,N_29214);
xnor U30594 (N_30594,N_29922,N_28424);
and U30595 (N_30595,N_28777,N_28995);
xor U30596 (N_30596,N_28518,N_29222);
xnor U30597 (N_30597,N_29829,N_29070);
or U30598 (N_30598,N_29447,N_28150);
xnor U30599 (N_30599,N_28764,N_28367);
and U30600 (N_30600,N_29318,N_28273);
or U30601 (N_30601,N_28304,N_28532);
and U30602 (N_30602,N_28625,N_29656);
or U30603 (N_30603,N_29257,N_28428);
nor U30604 (N_30604,N_29154,N_29177);
or U30605 (N_30605,N_29242,N_28797);
nor U30606 (N_30606,N_29175,N_29158);
nor U30607 (N_30607,N_28655,N_29739);
or U30608 (N_30608,N_29094,N_29596);
and U30609 (N_30609,N_28473,N_29743);
and U30610 (N_30610,N_28251,N_29305);
nand U30611 (N_30611,N_29616,N_28971);
nor U30612 (N_30612,N_28340,N_28719);
or U30613 (N_30613,N_28621,N_28295);
and U30614 (N_30614,N_29152,N_29885);
nand U30615 (N_30615,N_29320,N_28896);
nand U30616 (N_30616,N_28994,N_28202);
nor U30617 (N_30617,N_29053,N_28783);
and U30618 (N_30618,N_28829,N_29975);
and U30619 (N_30619,N_29085,N_29755);
nand U30620 (N_30620,N_29878,N_29080);
nor U30621 (N_30621,N_28227,N_29916);
nand U30622 (N_30622,N_28284,N_29827);
or U30623 (N_30623,N_29535,N_29102);
nor U30624 (N_30624,N_29716,N_28168);
nand U30625 (N_30625,N_28668,N_29888);
nand U30626 (N_30626,N_28306,N_29773);
nor U30627 (N_30627,N_28702,N_28637);
nor U30628 (N_30628,N_28356,N_29065);
nor U30629 (N_30629,N_28187,N_28459);
xnor U30630 (N_30630,N_28319,N_28122);
xor U30631 (N_30631,N_29327,N_29482);
or U30632 (N_30632,N_29615,N_28005);
nor U30633 (N_30633,N_29977,N_29619);
and U30634 (N_30634,N_28897,N_29470);
and U30635 (N_30635,N_28064,N_29572);
nor U30636 (N_30636,N_28810,N_28675);
nor U30637 (N_30637,N_28049,N_29037);
or U30638 (N_30638,N_29686,N_29346);
nand U30639 (N_30639,N_29108,N_28236);
nand U30640 (N_30640,N_29641,N_28564);
or U30641 (N_30641,N_29963,N_29799);
xnor U30642 (N_30642,N_28335,N_29400);
xor U30643 (N_30643,N_28807,N_28014);
or U30644 (N_30644,N_28282,N_28370);
nand U30645 (N_30645,N_28103,N_28708);
nor U30646 (N_30646,N_29296,N_29467);
xor U30647 (N_30647,N_29269,N_29727);
xor U30648 (N_30648,N_29721,N_28690);
xor U30649 (N_30649,N_28872,N_28645);
xnor U30650 (N_30650,N_29081,N_29326);
xor U30651 (N_30651,N_29475,N_28589);
nand U30652 (N_30652,N_28214,N_29292);
and U30653 (N_30653,N_29096,N_28467);
nor U30654 (N_30654,N_28937,N_29671);
and U30655 (N_30655,N_28311,N_28423);
or U30656 (N_30656,N_29679,N_29386);
nand U30657 (N_30657,N_29258,N_29655);
or U30658 (N_30658,N_29209,N_28199);
xor U30659 (N_30659,N_28402,N_28212);
nand U30660 (N_30660,N_28603,N_28287);
nor U30661 (N_30661,N_29486,N_29330);
or U30662 (N_30662,N_29443,N_29420);
xnor U30663 (N_30663,N_29576,N_29374);
xor U30664 (N_30664,N_28336,N_28399);
xnor U30665 (N_30665,N_29927,N_28438);
nor U30666 (N_30666,N_29044,N_29772);
or U30667 (N_30667,N_28194,N_28885);
nand U30668 (N_30668,N_28209,N_28420);
nor U30669 (N_30669,N_29607,N_29033);
xor U30670 (N_30670,N_29633,N_28085);
and U30671 (N_30671,N_28469,N_29186);
nand U30672 (N_30672,N_28726,N_28957);
or U30673 (N_30673,N_29957,N_29593);
and U30674 (N_30674,N_28028,N_28990);
xnor U30675 (N_30675,N_28641,N_29523);
xnor U30676 (N_30676,N_28147,N_29946);
nor U30677 (N_30677,N_28569,N_29418);
xnor U30678 (N_30678,N_29485,N_29089);
nand U30679 (N_30679,N_29996,N_28698);
xnor U30680 (N_30680,N_29809,N_28247);
xnor U30681 (N_30681,N_29455,N_29504);
nor U30682 (N_30682,N_28056,N_29197);
and U30683 (N_30683,N_29674,N_29769);
nor U30684 (N_30684,N_29206,N_28226);
and U30685 (N_30685,N_28115,N_28174);
nor U30686 (N_30686,N_28267,N_29790);
nor U30687 (N_30687,N_28516,N_29125);
xnor U30688 (N_30688,N_29913,N_29128);
nor U30689 (N_30689,N_28035,N_29391);
or U30690 (N_30690,N_28470,N_29172);
or U30691 (N_30691,N_29101,N_29647);
or U30692 (N_30692,N_28992,N_28674);
or U30693 (N_30693,N_28106,N_28128);
xor U30694 (N_30694,N_28378,N_28395);
nor U30695 (N_30695,N_29953,N_29751);
nor U30696 (N_30696,N_28535,N_28338);
or U30697 (N_30697,N_28373,N_29382);
nor U30698 (N_30698,N_29591,N_28536);
xnor U30699 (N_30699,N_28827,N_28587);
xnor U30700 (N_30700,N_28389,N_29776);
and U30701 (N_30701,N_29561,N_29556);
nand U30702 (N_30702,N_29216,N_28908);
and U30703 (N_30703,N_28029,N_28328);
and U30704 (N_30704,N_28347,N_29660);
or U30705 (N_30705,N_29921,N_29087);
xnor U30706 (N_30706,N_29058,N_28960);
and U30707 (N_30707,N_29022,N_29493);
and U30708 (N_30708,N_28249,N_29387);
or U30709 (N_30709,N_29652,N_29853);
nand U30710 (N_30710,N_29958,N_29835);
xnor U30711 (N_30711,N_29029,N_28113);
and U30712 (N_30712,N_29357,N_28232);
nor U30713 (N_30713,N_29665,N_28087);
or U30714 (N_30714,N_28952,N_28316);
or U30715 (N_30715,N_28080,N_28682);
and U30716 (N_30716,N_29867,N_29567);
or U30717 (N_30717,N_29413,N_29217);
xnor U30718 (N_30718,N_29579,N_28610);
nor U30719 (N_30719,N_28344,N_29046);
nand U30720 (N_30720,N_29466,N_29610);
nor U30721 (N_30721,N_28463,N_28493);
nor U30722 (N_30722,N_28580,N_28545);
nand U30723 (N_30723,N_28009,N_29745);
and U30724 (N_30724,N_29857,N_28329);
nor U30725 (N_30725,N_29020,N_29934);
nor U30726 (N_30726,N_29223,N_29645);
and U30727 (N_30727,N_29598,N_28907);
xnor U30728 (N_30728,N_28391,N_28376);
or U30729 (N_30729,N_29496,N_29372);
xor U30730 (N_30730,N_29744,N_28899);
nor U30731 (N_30731,N_28228,N_29448);
nor U30732 (N_30732,N_28881,N_28258);
nor U30733 (N_30733,N_29248,N_28681);
nand U30734 (N_30734,N_29901,N_29465);
nor U30735 (N_30735,N_29042,N_28631);
xor U30736 (N_30736,N_29385,N_29983);
or U30737 (N_30737,N_28407,N_28008);
and U30738 (N_30738,N_29267,N_28133);
and U30739 (N_30739,N_28317,N_29918);
nor U30740 (N_30740,N_29323,N_29238);
nor U30741 (N_30741,N_28240,N_29105);
and U30742 (N_30742,N_29738,N_29821);
and U30743 (N_30743,N_29510,N_28745);
nand U30744 (N_30744,N_29352,N_29430);
nor U30745 (N_30745,N_28823,N_28862);
nand U30746 (N_30746,N_28023,N_28059);
xor U30747 (N_30747,N_28632,N_29321);
nor U30748 (N_30748,N_29956,N_29334);
nor U30749 (N_30749,N_28687,N_29332);
nand U30750 (N_30750,N_28422,N_29749);
nand U30751 (N_30751,N_29354,N_29417);
nor U30752 (N_30752,N_28368,N_28718);
nand U30753 (N_30753,N_29012,N_28117);
xnor U30754 (N_30754,N_29239,N_29842);
nor U30755 (N_30755,N_29925,N_28754);
or U30756 (N_30756,N_29376,N_29636);
or U30757 (N_30757,N_29370,N_28504);
nand U30758 (N_30758,N_28068,N_29256);
nand U30759 (N_30759,N_28953,N_29522);
and U30760 (N_30760,N_28089,N_28857);
or U30761 (N_30761,N_29422,N_29232);
and U30762 (N_30762,N_29449,N_29245);
xor U30763 (N_30763,N_28309,N_29200);
or U30764 (N_30764,N_29810,N_28649);
xor U30765 (N_30765,N_29995,N_29748);
and U30766 (N_30766,N_29637,N_29552);
xnor U30767 (N_30767,N_29302,N_28588);
xor U30768 (N_30768,N_28787,N_28933);
or U30769 (N_30769,N_29895,N_29049);
and U30770 (N_30770,N_29371,N_28471);
and U30771 (N_30771,N_29843,N_29450);
nor U30772 (N_30772,N_28778,N_29782);
or U30773 (N_30773,N_28653,N_28030);
xor U30774 (N_30774,N_29006,N_28741);
xor U30775 (N_30775,N_28988,N_29717);
nand U30776 (N_30776,N_28820,N_28007);
nand U30777 (N_30777,N_28716,N_28413);
or U30778 (N_30778,N_28720,N_28398);
or U30779 (N_30779,N_29488,N_29948);
nor U30780 (N_30780,N_28348,N_29998);
and U30781 (N_30781,N_28768,N_29115);
or U30782 (N_30782,N_28640,N_29629);
or U30783 (N_30783,N_28780,N_29631);
nor U30784 (N_30784,N_28243,N_28390);
nor U30785 (N_30785,N_28164,N_28149);
nand U30786 (N_30786,N_29384,N_28826);
nor U30787 (N_30787,N_28552,N_29971);
nand U30788 (N_30788,N_28260,N_29176);
nand U30789 (N_30789,N_29736,N_28097);
or U30790 (N_30790,N_29703,N_29225);
nor U30791 (N_30791,N_28006,N_28867);
and U30792 (N_30792,N_29937,N_28299);
or U30793 (N_30793,N_29559,N_29859);
nor U30794 (N_30794,N_29838,N_29694);
and U30795 (N_30795,N_29198,N_29899);
xnor U30796 (N_30796,N_29541,N_29140);
nor U30797 (N_30797,N_28303,N_29811);
or U30798 (N_30798,N_28978,N_28074);
and U30799 (N_30799,N_29580,N_28013);
nand U30800 (N_30800,N_28363,N_29994);
nand U30801 (N_30801,N_28384,N_28599);
or U30802 (N_30802,N_29756,N_28507);
nand U30803 (N_30803,N_29606,N_29935);
xor U30804 (N_30804,N_29889,N_29017);
and U30805 (N_30805,N_28330,N_29534);
xor U30806 (N_30806,N_29923,N_28856);
nand U30807 (N_30807,N_29907,N_28888);
or U30808 (N_30808,N_29949,N_29740);
nor U30809 (N_30809,N_28519,N_29281);
nand U30810 (N_30810,N_29110,N_29118);
or U30811 (N_30811,N_29910,N_29337);
nand U30812 (N_30812,N_28346,N_29622);
nor U30813 (N_30813,N_29570,N_28246);
xnor U30814 (N_30814,N_28654,N_28558);
nand U30815 (N_30815,N_29319,N_29423);
nor U30816 (N_30816,N_29185,N_29072);
or U30817 (N_30817,N_29545,N_28033);
xnor U30818 (N_30818,N_28913,N_28380);
and U30819 (N_30819,N_28750,N_28146);
xnor U30820 (N_30820,N_28592,N_29962);
nand U30821 (N_30821,N_29170,N_28377);
and U30822 (N_30822,N_29076,N_28835);
xor U30823 (N_30823,N_28461,N_28186);
xor U30824 (N_30824,N_29340,N_29299);
or U30825 (N_30825,N_29213,N_29083);
xnor U30826 (N_30826,N_29653,N_29571);
nor U30827 (N_30827,N_29624,N_28143);
nand U30828 (N_30828,N_29638,N_29905);
and U30829 (N_30829,N_29786,N_28241);
nand U30830 (N_30830,N_28683,N_28941);
or U30831 (N_30831,N_29312,N_28920);
nor U30832 (N_30832,N_28929,N_28746);
xnor U30833 (N_30833,N_28652,N_28130);
nor U30834 (N_30834,N_29762,N_28110);
or U30835 (N_30835,N_29480,N_29807);
xnor U30836 (N_30836,N_28879,N_28474);
or U30837 (N_30837,N_29473,N_29015);
xnor U30838 (N_30838,N_28546,N_29071);
or U30839 (N_30839,N_29035,N_29168);
nor U30840 (N_30840,N_29446,N_28853);
xnor U30841 (N_30841,N_29236,N_29784);
and U30842 (N_30842,N_29298,N_28121);
nand U30843 (N_30843,N_28759,N_28628);
or U30844 (N_30844,N_28958,N_28416);
xnor U30845 (N_30845,N_29585,N_29917);
xnor U30846 (N_30846,N_28677,N_29078);
xor U30847 (N_30847,N_29136,N_28204);
or U30848 (N_30848,N_29846,N_29884);
nor U30849 (N_30849,N_29137,N_28352);
and U30850 (N_30850,N_28659,N_29691);
nand U30851 (N_30851,N_28024,N_29489);
nor U30852 (N_30852,N_29283,N_28842);
nand U30853 (N_30853,N_29173,N_28847);
or U30854 (N_30854,N_28381,N_28973);
xor U30855 (N_30855,N_28685,N_29830);
and U30856 (N_30856,N_29338,N_28167);
or U30857 (N_30857,N_29824,N_28693);
nand U30858 (N_30858,N_29940,N_28722);
or U30859 (N_30859,N_29231,N_28184);
nor U30860 (N_30860,N_28964,N_28993);
and U30861 (N_30861,N_28192,N_28447);
xor U30862 (N_30862,N_28270,N_29284);
xnor U30863 (N_30863,N_28642,N_29218);
or U30864 (N_30864,N_28019,N_29941);
or U30865 (N_30865,N_29775,N_29419);
and U30866 (N_30866,N_29324,N_28673);
xnor U30867 (N_30867,N_29658,N_29375);
or U30868 (N_30868,N_28822,N_29290);
nor U30869 (N_30869,N_28755,N_28522);
or U30870 (N_30870,N_29820,N_29263);
nor U30871 (N_30871,N_28084,N_29084);
and U30872 (N_30872,N_29873,N_28274);
nand U30873 (N_30873,N_29558,N_28181);
nand U30874 (N_30874,N_29395,N_29398);
nor U30875 (N_30875,N_29066,N_29794);
nor U30876 (N_30876,N_28448,N_28077);
and U30877 (N_30877,N_28946,N_29461);
or U30878 (N_30878,N_28286,N_29243);
and U30879 (N_30879,N_29162,N_29141);
nor U30880 (N_30880,N_29735,N_28462);
nor U30881 (N_30881,N_29919,N_29802);
nand U30882 (N_30882,N_29454,N_28784);
or U30883 (N_30883,N_28721,N_29405);
or U30884 (N_30884,N_29230,N_28567);
nand U30885 (N_30885,N_28643,N_29965);
xnor U30886 (N_30886,N_28195,N_28521);
and U30887 (N_30887,N_28966,N_28154);
xnor U30888 (N_30888,N_29234,N_28025);
and U30889 (N_30889,N_29904,N_29056);
or U30890 (N_30890,N_28302,N_29855);
xnor U30891 (N_30891,N_28431,N_28451);
nor U30892 (N_30892,N_28861,N_29573);
and U30893 (N_30893,N_29187,N_28213);
nand U30894 (N_30894,N_28724,N_28594);
nor U30895 (N_30895,N_28102,N_29847);
nor U30896 (N_30896,N_28912,N_29715);
nand U30897 (N_30897,N_28932,N_29451);
and U30898 (N_30898,N_28163,N_28239);
and U30899 (N_30899,N_29704,N_28813);
xnor U30900 (N_30900,N_29968,N_28139);
and U30901 (N_30901,N_29682,N_28571);
and U30902 (N_30902,N_28410,N_29163);
xnor U30903 (N_30903,N_29803,N_28831);
or U30904 (N_30904,N_29075,N_28927);
nand U30905 (N_30905,N_28874,N_28433);
and U30906 (N_30906,N_28159,N_28158);
xor U30907 (N_30907,N_28176,N_28177);
or U30908 (N_30908,N_28733,N_29378);
nand U30909 (N_30909,N_29207,N_29191);
and U30910 (N_30910,N_29954,N_29648);
or U30911 (N_30911,N_28503,N_28230);
xor U30912 (N_30912,N_28887,N_28613);
xnor U30913 (N_30913,N_28562,N_29410);
or U30914 (N_30914,N_28218,N_28801);
xnor U30915 (N_30915,N_29549,N_28203);
nor U30916 (N_30916,N_29498,N_29920);
and U30917 (N_30917,N_28124,N_28622);
nand U30918 (N_30918,N_28152,N_28566);
xor U30919 (N_30919,N_29192,N_28841);
xor U30920 (N_30920,N_29490,N_29822);
nand U30921 (N_30921,N_28486,N_29861);
and U30922 (N_30922,N_28802,N_28366);
or U30923 (N_30923,N_29984,N_29702);
nand U30924 (N_30924,N_29780,N_28590);
or U30925 (N_30925,N_29684,N_29016);
nor U30926 (N_30926,N_29463,N_28001);
nor U30927 (N_30927,N_28418,N_29583);
or U30928 (N_30928,N_28224,N_29255);
nor U30929 (N_30929,N_29777,N_28369);
nor U30930 (N_30930,N_29742,N_29282);
or U30931 (N_30931,N_28406,N_29562);
nand U30932 (N_30932,N_29605,N_29119);
and U30933 (N_30933,N_28624,N_28936);
xnor U30934 (N_30934,N_28278,N_28044);
or U30935 (N_30935,N_29858,N_29711);
and U30936 (N_30936,N_29981,N_29342);
and U30937 (N_30937,N_28475,N_28962);
xnor U30938 (N_30938,N_29951,N_29100);
xor U30939 (N_30939,N_28633,N_28838);
xnor U30940 (N_30940,N_29877,N_28185);
xnor U30941 (N_30941,N_28310,N_28554);
and U30942 (N_30942,N_28450,N_28987);
nor U30943 (N_30943,N_28225,N_28981);
and U30944 (N_30944,N_29732,N_29379);
nand U30945 (N_30945,N_28735,N_28472);
nand U30946 (N_30946,N_28411,N_29341);
nand U30947 (N_30947,N_29626,N_29013);
or U30948 (N_30948,N_28620,N_29911);
nor U30949 (N_30949,N_28760,N_28765);
xor U30950 (N_30950,N_28581,N_29050);
xnor U30951 (N_30951,N_28300,N_28618);
nand U30952 (N_30952,N_28709,N_28530);
nor U30953 (N_30953,N_28707,N_29456);
nor U30954 (N_30954,N_29221,N_29433);
and U30955 (N_30955,N_29442,N_29350);
or U30956 (N_30956,N_28734,N_29623);
nand U30957 (N_30957,N_28803,N_29869);
nand U30958 (N_30958,N_28511,N_29590);
and U30959 (N_30959,N_28134,N_28809);
xor U30960 (N_30960,N_28298,N_29597);
nor U30961 (N_30961,N_29397,N_28083);
nor U30962 (N_30962,N_28712,N_28871);
nand U30963 (N_30963,N_28834,N_28052);
xor U30964 (N_30964,N_29685,N_28307);
xnor U30965 (N_30965,N_28651,N_28798);
or U30966 (N_30966,N_29212,N_29235);
or U30967 (N_30967,N_28715,N_29394);
and U30968 (N_30968,N_28365,N_29483);
xnor U30969 (N_30969,N_28969,N_28883);
xor U30970 (N_30970,N_28138,N_28694);
nand U30971 (N_30971,N_28865,N_28027);
or U30972 (N_30972,N_28744,N_29870);
nand U30973 (N_30973,N_28466,N_28509);
nand U30974 (N_30974,N_29517,N_29550);
nand U30975 (N_30975,N_29007,N_29392);
xor U30976 (N_30976,N_29865,N_29272);
or U30977 (N_30977,N_29876,N_28691);
nand U30978 (N_30978,N_28884,N_28354);
xor U30979 (N_30979,N_29153,N_28968);
xor U30980 (N_30980,N_29194,N_28125);
and U30981 (N_30981,N_29529,N_29220);
xor U30982 (N_30982,N_29569,N_28544);
or U30983 (N_30983,N_29668,N_28207);
xnor U30984 (N_30984,N_28664,N_29502);
nor U30985 (N_30985,N_29546,N_29407);
and U30986 (N_30986,N_28584,N_29285);
or U30987 (N_30987,N_29795,N_29592);
xnor U30988 (N_30988,N_29882,N_28201);
or U30989 (N_30989,N_28921,N_28614);
nor U30990 (N_30990,N_28846,N_28858);
and U30991 (N_30991,N_29439,N_29519);
xor U30992 (N_30992,N_29947,N_29010);
nand U30993 (N_30993,N_29757,N_29521);
or U30994 (N_30994,N_29600,N_28015);
and U30995 (N_30995,N_28045,N_29054);
or U30996 (N_30996,N_29804,N_28242);
nor U30997 (N_30997,N_28308,N_28982);
nor U30998 (N_30998,N_28796,N_29774);
nand U30999 (N_30999,N_28119,N_29687);
xnor U31000 (N_31000,N_28845,N_29698);
or U31001 (N_31001,N_28258,N_28761);
or U31002 (N_31002,N_29868,N_28459);
xnor U31003 (N_31003,N_28206,N_28693);
xnor U31004 (N_31004,N_28488,N_29634);
nor U31005 (N_31005,N_28071,N_29042);
xnor U31006 (N_31006,N_28715,N_29959);
or U31007 (N_31007,N_29033,N_28004);
xnor U31008 (N_31008,N_28614,N_29293);
nand U31009 (N_31009,N_29539,N_29647);
or U31010 (N_31010,N_28546,N_28702);
or U31011 (N_31011,N_28725,N_29743);
or U31012 (N_31012,N_29534,N_28397);
xor U31013 (N_31013,N_28814,N_28472);
nand U31014 (N_31014,N_29387,N_29748);
and U31015 (N_31015,N_28594,N_28926);
and U31016 (N_31016,N_29171,N_29317);
nand U31017 (N_31017,N_28589,N_29182);
or U31018 (N_31018,N_28009,N_28860);
nor U31019 (N_31019,N_28942,N_28440);
nand U31020 (N_31020,N_29942,N_28495);
xnor U31021 (N_31021,N_28475,N_29284);
nand U31022 (N_31022,N_28192,N_29521);
nor U31023 (N_31023,N_28535,N_28009);
or U31024 (N_31024,N_29645,N_29743);
nand U31025 (N_31025,N_28110,N_29892);
and U31026 (N_31026,N_28344,N_29804);
and U31027 (N_31027,N_28825,N_29016);
nor U31028 (N_31028,N_28363,N_28156);
or U31029 (N_31029,N_28697,N_28731);
or U31030 (N_31030,N_28264,N_28768);
or U31031 (N_31031,N_29132,N_28180);
nor U31032 (N_31032,N_28607,N_28671);
nand U31033 (N_31033,N_28384,N_29100);
xnor U31034 (N_31034,N_28166,N_28609);
nand U31035 (N_31035,N_29887,N_29129);
or U31036 (N_31036,N_29804,N_29403);
and U31037 (N_31037,N_28371,N_29605);
nand U31038 (N_31038,N_28680,N_29476);
nand U31039 (N_31039,N_28886,N_28821);
and U31040 (N_31040,N_29497,N_29694);
xnor U31041 (N_31041,N_28314,N_29335);
nand U31042 (N_31042,N_29134,N_29021);
xor U31043 (N_31043,N_28938,N_29275);
nand U31044 (N_31044,N_28777,N_29125);
nor U31045 (N_31045,N_28414,N_29348);
nor U31046 (N_31046,N_29585,N_28630);
or U31047 (N_31047,N_28601,N_29989);
xor U31048 (N_31048,N_29263,N_29374);
or U31049 (N_31049,N_28757,N_28692);
and U31050 (N_31050,N_29199,N_29720);
nor U31051 (N_31051,N_28025,N_28017);
or U31052 (N_31052,N_28678,N_28533);
nor U31053 (N_31053,N_29781,N_29954);
nor U31054 (N_31054,N_28032,N_29235);
nand U31055 (N_31055,N_29916,N_28675);
nor U31056 (N_31056,N_28255,N_29382);
nand U31057 (N_31057,N_28689,N_28584);
nand U31058 (N_31058,N_29726,N_28456);
nor U31059 (N_31059,N_29927,N_28621);
xor U31060 (N_31060,N_29115,N_28284);
nor U31061 (N_31061,N_29494,N_29462);
and U31062 (N_31062,N_28450,N_29917);
or U31063 (N_31063,N_28418,N_28271);
xnor U31064 (N_31064,N_28442,N_28365);
nor U31065 (N_31065,N_28880,N_28845);
and U31066 (N_31066,N_28822,N_29075);
nor U31067 (N_31067,N_28466,N_28781);
nand U31068 (N_31068,N_28332,N_29123);
nor U31069 (N_31069,N_29621,N_29488);
nand U31070 (N_31070,N_28546,N_28970);
and U31071 (N_31071,N_29144,N_28743);
or U31072 (N_31072,N_28678,N_28218);
xor U31073 (N_31073,N_29861,N_29792);
or U31074 (N_31074,N_29303,N_29592);
nor U31075 (N_31075,N_29503,N_28136);
xor U31076 (N_31076,N_29203,N_28125);
xor U31077 (N_31077,N_29815,N_29291);
and U31078 (N_31078,N_29372,N_28241);
nor U31079 (N_31079,N_29784,N_28957);
nand U31080 (N_31080,N_28633,N_28398);
and U31081 (N_31081,N_29614,N_28743);
and U31082 (N_31082,N_29613,N_28852);
or U31083 (N_31083,N_29591,N_28677);
or U31084 (N_31084,N_29354,N_28041);
or U31085 (N_31085,N_28659,N_29641);
xnor U31086 (N_31086,N_29610,N_28774);
nand U31087 (N_31087,N_28418,N_28475);
nor U31088 (N_31088,N_29788,N_28974);
nor U31089 (N_31089,N_28402,N_29189);
xor U31090 (N_31090,N_29616,N_28696);
xnor U31091 (N_31091,N_29762,N_29757);
and U31092 (N_31092,N_28814,N_29890);
and U31093 (N_31093,N_28306,N_29876);
or U31094 (N_31094,N_28983,N_28823);
or U31095 (N_31095,N_29419,N_29149);
xor U31096 (N_31096,N_29484,N_28155);
or U31097 (N_31097,N_29818,N_29770);
and U31098 (N_31098,N_28758,N_29424);
or U31099 (N_31099,N_29863,N_29474);
xnor U31100 (N_31100,N_29141,N_29308);
and U31101 (N_31101,N_29504,N_29060);
xnor U31102 (N_31102,N_28396,N_28074);
or U31103 (N_31103,N_29078,N_29881);
xnor U31104 (N_31104,N_28559,N_28604);
nor U31105 (N_31105,N_28985,N_29202);
nand U31106 (N_31106,N_28809,N_29853);
xor U31107 (N_31107,N_29648,N_28930);
or U31108 (N_31108,N_29544,N_29399);
nor U31109 (N_31109,N_28277,N_28268);
and U31110 (N_31110,N_28529,N_29145);
and U31111 (N_31111,N_29657,N_29483);
and U31112 (N_31112,N_28895,N_29006);
or U31113 (N_31113,N_29631,N_28822);
nand U31114 (N_31114,N_28178,N_28593);
or U31115 (N_31115,N_28464,N_28244);
nor U31116 (N_31116,N_29080,N_29296);
xor U31117 (N_31117,N_29165,N_29306);
or U31118 (N_31118,N_28617,N_29864);
and U31119 (N_31119,N_29247,N_28341);
and U31120 (N_31120,N_29501,N_29222);
nand U31121 (N_31121,N_29695,N_28032);
and U31122 (N_31122,N_29846,N_28626);
or U31123 (N_31123,N_28869,N_29696);
xnor U31124 (N_31124,N_28930,N_29128);
xnor U31125 (N_31125,N_29747,N_28700);
xnor U31126 (N_31126,N_29585,N_29492);
and U31127 (N_31127,N_29728,N_28386);
xor U31128 (N_31128,N_29545,N_29006);
nand U31129 (N_31129,N_28432,N_29114);
or U31130 (N_31130,N_28122,N_28078);
nor U31131 (N_31131,N_29878,N_28325);
xnor U31132 (N_31132,N_29679,N_28409);
nor U31133 (N_31133,N_29068,N_29796);
nor U31134 (N_31134,N_28576,N_28597);
or U31135 (N_31135,N_29463,N_28841);
and U31136 (N_31136,N_28690,N_29567);
nand U31137 (N_31137,N_29424,N_28604);
xor U31138 (N_31138,N_28932,N_28563);
and U31139 (N_31139,N_29751,N_29635);
xor U31140 (N_31140,N_29983,N_29855);
or U31141 (N_31141,N_28990,N_28458);
xnor U31142 (N_31142,N_29665,N_29396);
and U31143 (N_31143,N_29668,N_28154);
or U31144 (N_31144,N_29548,N_28771);
and U31145 (N_31145,N_28714,N_28709);
xor U31146 (N_31146,N_28989,N_28498);
or U31147 (N_31147,N_28666,N_29595);
nand U31148 (N_31148,N_29520,N_29920);
or U31149 (N_31149,N_28736,N_28285);
or U31150 (N_31150,N_29185,N_29028);
nor U31151 (N_31151,N_28562,N_29099);
xnor U31152 (N_31152,N_28207,N_29748);
nor U31153 (N_31153,N_29571,N_29033);
nand U31154 (N_31154,N_29111,N_28728);
or U31155 (N_31155,N_29426,N_29755);
xor U31156 (N_31156,N_28739,N_28676);
or U31157 (N_31157,N_29057,N_29106);
xor U31158 (N_31158,N_29002,N_28227);
nand U31159 (N_31159,N_29420,N_28224);
xor U31160 (N_31160,N_29280,N_29768);
nand U31161 (N_31161,N_29396,N_28367);
nor U31162 (N_31162,N_29714,N_28281);
and U31163 (N_31163,N_28876,N_29334);
or U31164 (N_31164,N_28183,N_28643);
nor U31165 (N_31165,N_28057,N_29545);
or U31166 (N_31166,N_29330,N_28069);
or U31167 (N_31167,N_29248,N_28797);
or U31168 (N_31168,N_28130,N_28945);
and U31169 (N_31169,N_29512,N_28372);
nor U31170 (N_31170,N_29864,N_28531);
or U31171 (N_31171,N_29464,N_29276);
xor U31172 (N_31172,N_28974,N_28529);
and U31173 (N_31173,N_28821,N_29099);
or U31174 (N_31174,N_29980,N_28496);
xor U31175 (N_31175,N_29721,N_28631);
or U31176 (N_31176,N_28206,N_29167);
xor U31177 (N_31177,N_28445,N_28684);
nand U31178 (N_31178,N_29571,N_29816);
nand U31179 (N_31179,N_29054,N_29485);
and U31180 (N_31180,N_28299,N_28185);
nor U31181 (N_31181,N_29750,N_29049);
nand U31182 (N_31182,N_28404,N_29533);
xor U31183 (N_31183,N_28211,N_28931);
xnor U31184 (N_31184,N_29070,N_28059);
xor U31185 (N_31185,N_29060,N_28354);
nor U31186 (N_31186,N_28592,N_28887);
and U31187 (N_31187,N_28251,N_28293);
nand U31188 (N_31188,N_28227,N_29413);
xor U31189 (N_31189,N_29672,N_28712);
xnor U31190 (N_31190,N_29182,N_28192);
or U31191 (N_31191,N_29696,N_29672);
xnor U31192 (N_31192,N_29063,N_29712);
xor U31193 (N_31193,N_28344,N_29591);
xor U31194 (N_31194,N_29174,N_28840);
and U31195 (N_31195,N_29319,N_29438);
xor U31196 (N_31196,N_28797,N_28558);
xnor U31197 (N_31197,N_29942,N_29188);
and U31198 (N_31198,N_29371,N_28940);
xor U31199 (N_31199,N_29418,N_29844);
xnor U31200 (N_31200,N_28738,N_29724);
nand U31201 (N_31201,N_28651,N_28040);
or U31202 (N_31202,N_29952,N_29770);
and U31203 (N_31203,N_28231,N_29100);
xor U31204 (N_31204,N_28902,N_29197);
or U31205 (N_31205,N_29999,N_28706);
nand U31206 (N_31206,N_29523,N_29512);
nand U31207 (N_31207,N_28579,N_28945);
or U31208 (N_31208,N_29124,N_29528);
xor U31209 (N_31209,N_29984,N_28101);
xor U31210 (N_31210,N_28038,N_28821);
nand U31211 (N_31211,N_29116,N_29478);
or U31212 (N_31212,N_28628,N_28321);
xor U31213 (N_31213,N_28082,N_28529);
xnor U31214 (N_31214,N_28424,N_28459);
and U31215 (N_31215,N_29937,N_29867);
nor U31216 (N_31216,N_29394,N_28086);
xor U31217 (N_31217,N_29700,N_28235);
and U31218 (N_31218,N_29782,N_29451);
and U31219 (N_31219,N_28370,N_28421);
nand U31220 (N_31220,N_29371,N_28043);
or U31221 (N_31221,N_29945,N_29126);
or U31222 (N_31222,N_29362,N_28461);
xnor U31223 (N_31223,N_28290,N_28919);
xnor U31224 (N_31224,N_29782,N_28072);
nor U31225 (N_31225,N_28016,N_28326);
nor U31226 (N_31226,N_28151,N_28554);
nor U31227 (N_31227,N_28553,N_29980);
nand U31228 (N_31228,N_28440,N_28249);
nand U31229 (N_31229,N_29500,N_29629);
and U31230 (N_31230,N_29495,N_28602);
nor U31231 (N_31231,N_29936,N_28492);
and U31232 (N_31232,N_29670,N_29464);
nor U31233 (N_31233,N_28959,N_28859);
or U31234 (N_31234,N_28936,N_29842);
and U31235 (N_31235,N_28543,N_28024);
nor U31236 (N_31236,N_28606,N_28265);
xnor U31237 (N_31237,N_28486,N_29113);
and U31238 (N_31238,N_28281,N_29150);
nand U31239 (N_31239,N_28504,N_29606);
xor U31240 (N_31240,N_29474,N_29141);
nor U31241 (N_31241,N_28394,N_29776);
xnor U31242 (N_31242,N_29123,N_28327);
xnor U31243 (N_31243,N_29379,N_29920);
xnor U31244 (N_31244,N_28445,N_29699);
and U31245 (N_31245,N_29070,N_28880);
xnor U31246 (N_31246,N_28914,N_28457);
xor U31247 (N_31247,N_29221,N_28222);
or U31248 (N_31248,N_28682,N_28120);
xor U31249 (N_31249,N_29326,N_28590);
or U31250 (N_31250,N_28007,N_28922);
and U31251 (N_31251,N_28913,N_29376);
nand U31252 (N_31252,N_28451,N_28120);
and U31253 (N_31253,N_28018,N_28613);
or U31254 (N_31254,N_29957,N_29444);
xnor U31255 (N_31255,N_29756,N_29732);
nor U31256 (N_31256,N_28722,N_29516);
or U31257 (N_31257,N_29542,N_28443);
and U31258 (N_31258,N_29054,N_29493);
nor U31259 (N_31259,N_29833,N_28501);
nand U31260 (N_31260,N_28914,N_29551);
or U31261 (N_31261,N_28906,N_28087);
and U31262 (N_31262,N_29129,N_29509);
nand U31263 (N_31263,N_28451,N_29101);
xor U31264 (N_31264,N_28740,N_29273);
and U31265 (N_31265,N_29558,N_28503);
and U31266 (N_31266,N_29293,N_28509);
xor U31267 (N_31267,N_29608,N_28679);
and U31268 (N_31268,N_28482,N_29809);
and U31269 (N_31269,N_28903,N_29485);
or U31270 (N_31270,N_28285,N_28492);
xor U31271 (N_31271,N_29628,N_29899);
nand U31272 (N_31272,N_29561,N_28624);
or U31273 (N_31273,N_28071,N_29223);
nand U31274 (N_31274,N_29254,N_29983);
xor U31275 (N_31275,N_29770,N_28512);
and U31276 (N_31276,N_28330,N_28528);
and U31277 (N_31277,N_28887,N_28609);
nand U31278 (N_31278,N_28643,N_28751);
or U31279 (N_31279,N_28829,N_28385);
or U31280 (N_31280,N_28359,N_28187);
or U31281 (N_31281,N_28622,N_29580);
or U31282 (N_31282,N_28234,N_29155);
nor U31283 (N_31283,N_29509,N_28238);
nor U31284 (N_31284,N_29528,N_28342);
xor U31285 (N_31285,N_29882,N_29477);
nor U31286 (N_31286,N_28731,N_29179);
nand U31287 (N_31287,N_29058,N_28245);
xor U31288 (N_31288,N_29801,N_29411);
and U31289 (N_31289,N_29875,N_28996);
nor U31290 (N_31290,N_29408,N_28479);
nor U31291 (N_31291,N_29184,N_29634);
nand U31292 (N_31292,N_28208,N_29666);
and U31293 (N_31293,N_29423,N_29646);
nand U31294 (N_31294,N_28421,N_28827);
and U31295 (N_31295,N_29828,N_28925);
nand U31296 (N_31296,N_28037,N_28631);
xnor U31297 (N_31297,N_29614,N_29182);
nand U31298 (N_31298,N_29561,N_29272);
or U31299 (N_31299,N_29118,N_29488);
xnor U31300 (N_31300,N_29084,N_28717);
or U31301 (N_31301,N_28587,N_28523);
and U31302 (N_31302,N_28891,N_29463);
or U31303 (N_31303,N_29127,N_28762);
nand U31304 (N_31304,N_29802,N_28588);
and U31305 (N_31305,N_28065,N_28240);
nor U31306 (N_31306,N_28943,N_28939);
and U31307 (N_31307,N_29581,N_28613);
nand U31308 (N_31308,N_28028,N_29368);
and U31309 (N_31309,N_29305,N_28032);
xnor U31310 (N_31310,N_28592,N_29318);
nand U31311 (N_31311,N_29682,N_28242);
nor U31312 (N_31312,N_28099,N_28567);
nand U31313 (N_31313,N_29687,N_29124);
nand U31314 (N_31314,N_29054,N_28980);
or U31315 (N_31315,N_29609,N_28930);
or U31316 (N_31316,N_29139,N_29760);
xor U31317 (N_31317,N_28772,N_28704);
and U31318 (N_31318,N_28219,N_29861);
nand U31319 (N_31319,N_29514,N_28182);
xnor U31320 (N_31320,N_28777,N_28012);
xnor U31321 (N_31321,N_29519,N_29669);
nand U31322 (N_31322,N_28156,N_28878);
or U31323 (N_31323,N_28407,N_29097);
nand U31324 (N_31324,N_28273,N_29453);
and U31325 (N_31325,N_28592,N_29184);
xnor U31326 (N_31326,N_29517,N_28374);
nand U31327 (N_31327,N_28066,N_29011);
nor U31328 (N_31328,N_28601,N_29153);
or U31329 (N_31329,N_29862,N_29681);
xnor U31330 (N_31330,N_29752,N_28317);
nor U31331 (N_31331,N_29302,N_29558);
xnor U31332 (N_31332,N_28675,N_28453);
or U31333 (N_31333,N_28931,N_28237);
and U31334 (N_31334,N_29113,N_28273);
nand U31335 (N_31335,N_29956,N_28880);
xnor U31336 (N_31336,N_29383,N_28616);
or U31337 (N_31337,N_29203,N_29128);
xor U31338 (N_31338,N_28374,N_29212);
nand U31339 (N_31339,N_28717,N_28289);
and U31340 (N_31340,N_29168,N_29350);
xnor U31341 (N_31341,N_28181,N_28415);
xnor U31342 (N_31342,N_29568,N_28601);
nand U31343 (N_31343,N_28393,N_29013);
or U31344 (N_31344,N_28014,N_29241);
or U31345 (N_31345,N_29661,N_29128);
and U31346 (N_31346,N_28106,N_28304);
xnor U31347 (N_31347,N_29900,N_28737);
nand U31348 (N_31348,N_28730,N_29042);
xor U31349 (N_31349,N_29359,N_29302);
xnor U31350 (N_31350,N_29031,N_28593);
and U31351 (N_31351,N_29280,N_28053);
or U31352 (N_31352,N_29700,N_29175);
nand U31353 (N_31353,N_29672,N_28833);
nor U31354 (N_31354,N_29930,N_29079);
and U31355 (N_31355,N_29492,N_29969);
xnor U31356 (N_31356,N_28362,N_29196);
nand U31357 (N_31357,N_29555,N_28831);
and U31358 (N_31358,N_28987,N_28728);
and U31359 (N_31359,N_29821,N_28682);
nand U31360 (N_31360,N_29352,N_29703);
or U31361 (N_31361,N_29614,N_28676);
nand U31362 (N_31362,N_29145,N_28144);
nand U31363 (N_31363,N_28434,N_28501);
and U31364 (N_31364,N_29749,N_28512);
and U31365 (N_31365,N_28923,N_28688);
nor U31366 (N_31366,N_28695,N_28861);
and U31367 (N_31367,N_29107,N_28771);
nor U31368 (N_31368,N_29006,N_28715);
nor U31369 (N_31369,N_29942,N_28615);
nand U31370 (N_31370,N_29944,N_29841);
and U31371 (N_31371,N_29014,N_28256);
or U31372 (N_31372,N_28118,N_28772);
xor U31373 (N_31373,N_29566,N_28762);
and U31374 (N_31374,N_28233,N_28599);
nor U31375 (N_31375,N_28430,N_28645);
nor U31376 (N_31376,N_29370,N_28354);
xnor U31377 (N_31377,N_29145,N_28394);
xnor U31378 (N_31378,N_29790,N_28350);
nand U31379 (N_31379,N_28128,N_29156);
nor U31380 (N_31380,N_28248,N_29261);
xnor U31381 (N_31381,N_28613,N_28578);
nand U31382 (N_31382,N_28419,N_29448);
xor U31383 (N_31383,N_28954,N_29394);
xor U31384 (N_31384,N_29771,N_29199);
and U31385 (N_31385,N_28984,N_28134);
nor U31386 (N_31386,N_29056,N_29110);
nand U31387 (N_31387,N_28661,N_28874);
xnor U31388 (N_31388,N_29060,N_28783);
and U31389 (N_31389,N_28734,N_28859);
and U31390 (N_31390,N_28772,N_29537);
xnor U31391 (N_31391,N_28099,N_28883);
xnor U31392 (N_31392,N_29912,N_29361);
and U31393 (N_31393,N_28975,N_28810);
nor U31394 (N_31394,N_29070,N_29403);
and U31395 (N_31395,N_28694,N_28791);
nor U31396 (N_31396,N_28478,N_28356);
xnor U31397 (N_31397,N_29007,N_29696);
nand U31398 (N_31398,N_28731,N_28764);
nand U31399 (N_31399,N_29271,N_28648);
nor U31400 (N_31400,N_29077,N_29577);
nand U31401 (N_31401,N_29437,N_28075);
xor U31402 (N_31402,N_28811,N_29701);
and U31403 (N_31403,N_29897,N_29782);
nor U31404 (N_31404,N_29119,N_29658);
xnor U31405 (N_31405,N_28338,N_29737);
and U31406 (N_31406,N_29060,N_28848);
nand U31407 (N_31407,N_29507,N_29301);
xnor U31408 (N_31408,N_29727,N_29286);
or U31409 (N_31409,N_28236,N_29325);
nand U31410 (N_31410,N_28809,N_28419);
nor U31411 (N_31411,N_28908,N_29960);
xnor U31412 (N_31412,N_29396,N_29109);
or U31413 (N_31413,N_29253,N_29488);
nand U31414 (N_31414,N_29325,N_28492);
nand U31415 (N_31415,N_28801,N_29529);
nand U31416 (N_31416,N_28644,N_29332);
or U31417 (N_31417,N_28392,N_28554);
nor U31418 (N_31418,N_29475,N_28022);
xor U31419 (N_31419,N_28967,N_29232);
or U31420 (N_31420,N_29341,N_28415);
and U31421 (N_31421,N_29942,N_28231);
xor U31422 (N_31422,N_29216,N_29964);
and U31423 (N_31423,N_28119,N_28068);
xnor U31424 (N_31424,N_29690,N_29719);
nor U31425 (N_31425,N_29182,N_28886);
xnor U31426 (N_31426,N_29970,N_29176);
or U31427 (N_31427,N_29364,N_28621);
or U31428 (N_31428,N_29423,N_29499);
or U31429 (N_31429,N_28917,N_29599);
nand U31430 (N_31430,N_28965,N_28081);
and U31431 (N_31431,N_29321,N_29326);
xnor U31432 (N_31432,N_29411,N_29223);
nand U31433 (N_31433,N_28726,N_29564);
nor U31434 (N_31434,N_29800,N_28253);
nor U31435 (N_31435,N_29839,N_28311);
nor U31436 (N_31436,N_29925,N_29701);
and U31437 (N_31437,N_29200,N_28238);
xnor U31438 (N_31438,N_29312,N_29687);
xor U31439 (N_31439,N_29796,N_28977);
and U31440 (N_31440,N_28534,N_29830);
nor U31441 (N_31441,N_29068,N_29069);
xnor U31442 (N_31442,N_28379,N_28891);
xnor U31443 (N_31443,N_29921,N_28606);
and U31444 (N_31444,N_28710,N_28057);
nor U31445 (N_31445,N_28360,N_28313);
nor U31446 (N_31446,N_28270,N_28546);
or U31447 (N_31447,N_28669,N_28798);
nor U31448 (N_31448,N_28012,N_28156);
and U31449 (N_31449,N_28333,N_29789);
xor U31450 (N_31450,N_28099,N_29083);
and U31451 (N_31451,N_28162,N_28963);
and U31452 (N_31452,N_28321,N_29133);
or U31453 (N_31453,N_28888,N_28978);
nand U31454 (N_31454,N_28071,N_28684);
nor U31455 (N_31455,N_29630,N_29715);
or U31456 (N_31456,N_29756,N_28792);
nor U31457 (N_31457,N_29960,N_29050);
nand U31458 (N_31458,N_29444,N_28215);
and U31459 (N_31459,N_28007,N_28957);
nand U31460 (N_31460,N_29991,N_29356);
nor U31461 (N_31461,N_28812,N_29327);
and U31462 (N_31462,N_29970,N_29347);
xnor U31463 (N_31463,N_28776,N_28162);
and U31464 (N_31464,N_29940,N_29888);
nor U31465 (N_31465,N_28327,N_29855);
nand U31466 (N_31466,N_28348,N_28336);
and U31467 (N_31467,N_29327,N_29415);
and U31468 (N_31468,N_29807,N_28084);
and U31469 (N_31469,N_28871,N_28099);
xnor U31470 (N_31470,N_28405,N_29675);
xor U31471 (N_31471,N_29589,N_28973);
nand U31472 (N_31472,N_29867,N_28562);
nand U31473 (N_31473,N_29833,N_28896);
or U31474 (N_31474,N_29713,N_28899);
or U31475 (N_31475,N_29823,N_28451);
or U31476 (N_31476,N_29239,N_29843);
or U31477 (N_31477,N_28890,N_28896);
nor U31478 (N_31478,N_29514,N_29633);
or U31479 (N_31479,N_29561,N_28055);
nor U31480 (N_31480,N_28312,N_28115);
xnor U31481 (N_31481,N_28158,N_28357);
nor U31482 (N_31482,N_29965,N_29322);
or U31483 (N_31483,N_29444,N_28710);
or U31484 (N_31484,N_29274,N_29155);
or U31485 (N_31485,N_29963,N_28709);
nor U31486 (N_31486,N_28682,N_29003);
xnor U31487 (N_31487,N_28962,N_28629);
and U31488 (N_31488,N_29044,N_28653);
and U31489 (N_31489,N_29213,N_29028);
nand U31490 (N_31490,N_28088,N_28071);
nor U31491 (N_31491,N_28024,N_28944);
xor U31492 (N_31492,N_28198,N_29481);
xnor U31493 (N_31493,N_29764,N_28669);
and U31494 (N_31494,N_29715,N_29323);
or U31495 (N_31495,N_29923,N_28411);
or U31496 (N_31496,N_28735,N_29172);
nor U31497 (N_31497,N_28738,N_28759);
xnor U31498 (N_31498,N_29559,N_28382);
and U31499 (N_31499,N_28961,N_28900);
or U31500 (N_31500,N_28354,N_28454);
or U31501 (N_31501,N_28421,N_28826);
or U31502 (N_31502,N_29867,N_28396);
xnor U31503 (N_31503,N_28620,N_28107);
or U31504 (N_31504,N_29278,N_28384);
nand U31505 (N_31505,N_28700,N_29478);
and U31506 (N_31506,N_28427,N_28411);
nor U31507 (N_31507,N_28698,N_28820);
xnor U31508 (N_31508,N_29394,N_29609);
nor U31509 (N_31509,N_29493,N_29782);
nor U31510 (N_31510,N_28625,N_28147);
nor U31511 (N_31511,N_28874,N_28720);
xor U31512 (N_31512,N_28960,N_28117);
nand U31513 (N_31513,N_28122,N_29984);
nor U31514 (N_31514,N_29854,N_28627);
and U31515 (N_31515,N_28209,N_29402);
xnor U31516 (N_31516,N_29826,N_28186);
nor U31517 (N_31517,N_28341,N_29884);
or U31518 (N_31518,N_28891,N_29889);
nor U31519 (N_31519,N_28389,N_29349);
xor U31520 (N_31520,N_29859,N_29982);
nor U31521 (N_31521,N_29850,N_29609);
nor U31522 (N_31522,N_29405,N_29463);
or U31523 (N_31523,N_29211,N_28949);
nand U31524 (N_31524,N_28778,N_29650);
nand U31525 (N_31525,N_29195,N_28594);
nor U31526 (N_31526,N_28774,N_28646);
nand U31527 (N_31527,N_28604,N_29774);
or U31528 (N_31528,N_28102,N_29769);
xor U31529 (N_31529,N_28676,N_28971);
or U31530 (N_31530,N_28495,N_29403);
nand U31531 (N_31531,N_28901,N_28596);
xor U31532 (N_31532,N_28352,N_28204);
nor U31533 (N_31533,N_28217,N_28766);
nand U31534 (N_31534,N_29234,N_29427);
nand U31535 (N_31535,N_28924,N_28471);
and U31536 (N_31536,N_29978,N_28387);
nor U31537 (N_31537,N_28561,N_28779);
or U31538 (N_31538,N_28069,N_29092);
nor U31539 (N_31539,N_29831,N_29925);
and U31540 (N_31540,N_28000,N_29159);
xnor U31541 (N_31541,N_28944,N_28541);
nor U31542 (N_31542,N_28160,N_28177);
or U31543 (N_31543,N_29424,N_28105);
xor U31544 (N_31544,N_28851,N_28032);
xor U31545 (N_31545,N_28452,N_29473);
nand U31546 (N_31546,N_28912,N_28586);
nor U31547 (N_31547,N_29955,N_28816);
xnor U31548 (N_31548,N_28580,N_28789);
or U31549 (N_31549,N_28831,N_29009);
and U31550 (N_31550,N_29147,N_29415);
and U31551 (N_31551,N_28152,N_28563);
xor U31552 (N_31552,N_28376,N_28909);
nand U31553 (N_31553,N_28385,N_28625);
nand U31554 (N_31554,N_29058,N_29782);
nor U31555 (N_31555,N_29990,N_28646);
and U31556 (N_31556,N_28494,N_28246);
nand U31557 (N_31557,N_29763,N_28695);
nand U31558 (N_31558,N_29595,N_28492);
nor U31559 (N_31559,N_28964,N_29649);
nand U31560 (N_31560,N_29178,N_28626);
xor U31561 (N_31561,N_28887,N_28208);
and U31562 (N_31562,N_29644,N_28143);
nor U31563 (N_31563,N_28210,N_29849);
or U31564 (N_31564,N_28698,N_29987);
or U31565 (N_31565,N_28017,N_28396);
and U31566 (N_31566,N_28975,N_28960);
nand U31567 (N_31567,N_28282,N_29633);
or U31568 (N_31568,N_28372,N_29414);
and U31569 (N_31569,N_28754,N_29474);
nor U31570 (N_31570,N_29776,N_28116);
nor U31571 (N_31571,N_29298,N_28623);
and U31572 (N_31572,N_29099,N_29193);
nor U31573 (N_31573,N_29559,N_28010);
nand U31574 (N_31574,N_28691,N_29689);
or U31575 (N_31575,N_29504,N_29156);
xnor U31576 (N_31576,N_29817,N_29900);
nand U31577 (N_31577,N_28329,N_28752);
xor U31578 (N_31578,N_28388,N_28742);
and U31579 (N_31579,N_28670,N_29713);
nor U31580 (N_31580,N_28120,N_29264);
or U31581 (N_31581,N_29920,N_29094);
and U31582 (N_31582,N_29122,N_29566);
or U31583 (N_31583,N_29988,N_28024);
nor U31584 (N_31584,N_29499,N_29743);
or U31585 (N_31585,N_29576,N_29103);
xor U31586 (N_31586,N_28843,N_29697);
and U31587 (N_31587,N_29809,N_28256);
and U31588 (N_31588,N_28331,N_29513);
and U31589 (N_31589,N_28834,N_28846);
and U31590 (N_31590,N_28709,N_28256);
and U31591 (N_31591,N_28569,N_28771);
xor U31592 (N_31592,N_28295,N_29713);
nand U31593 (N_31593,N_29215,N_29970);
nand U31594 (N_31594,N_28785,N_28775);
or U31595 (N_31595,N_29228,N_28875);
nor U31596 (N_31596,N_28421,N_29424);
and U31597 (N_31597,N_28544,N_29829);
xnor U31598 (N_31598,N_29203,N_29347);
nor U31599 (N_31599,N_28389,N_28694);
nor U31600 (N_31600,N_29490,N_29443);
nor U31601 (N_31601,N_29395,N_28300);
or U31602 (N_31602,N_28817,N_28968);
or U31603 (N_31603,N_29768,N_29981);
nor U31604 (N_31604,N_28668,N_28600);
or U31605 (N_31605,N_28709,N_29970);
nor U31606 (N_31606,N_28396,N_29661);
xnor U31607 (N_31607,N_29298,N_28562);
nand U31608 (N_31608,N_28598,N_29100);
and U31609 (N_31609,N_29513,N_28614);
or U31610 (N_31610,N_29281,N_28284);
nand U31611 (N_31611,N_29627,N_29392);
nand U31612 (N_31612,N_28643,N_28717);
nor U31613 (N_31613,N_29438,N_28961);
nand U31614 (N_31614,N_29986,N_28132);
and U31615 (N_31615,N_29645,N_28147);
or U31616 (N_31616,N_29786,N_29289);
and U31617 (N_31617,N_29423,N_29824);
nand U31618 (N_31618,N_29964,N_28387);
and U31619 (N_31619,N_28709,N_28460);
nand U31620 (N_31620,N_29893,N_29451);
nor U31621 (N_31621,N_29016,N_28288);
nand U31622 (N_31622,N_28876,N_28517);
and U31623 (N_31623,N_28905,N_29662);
and U31624 (N_31624,N_28451,N_28902);
nand U31625 (N_31625,N_29166,N_29097);
or U31626 (N_31626,N_29070,N_28990);
or U31627 (N_31627,N_28181,N_29827);
and U31628 (N_31628,N_28944,N_29646);
or U31629 (N_31629,N_29858,N_28632);
nand U31630 (N_31630,N_29149,N_29644);
nand U31631 (N_31631,N_28674,N_29042);
nand U31632 (N_31632,N_29979,N_28379);
xor U31633 (N_31633,N_28633,N_28618);
nor U31634 (N_31634,N_29963,N_28317);
nand U31635 (N_31635,N_29659,N_28538);
xor U31636 (N_31636,N_29036,N_28648);
or U31637 (N_31637,N_29331,N_29441);
or U31638 (N_31638,N_28492,N_29944);
nor U31639 (N_31639,N_29160,N_28034);
xnor U31640 (N_31640,N_29594,N_28857);
nand U31641 (N_31641,N_28714,N_29201);
nor U31642 (N_31642,N_28553,N_29638);
or U31643 (N_31643,N_29499,N_28965);
or U31644 (N_31644,N_28330,N_28435);
nor U31645 (N_31645,N_28174,N_29789);
and U31646 (N_31646,N_29131,N_29183);
and U31647 (N_31647,N_29388,N_28016);
or U31648 (N_31648,N_28244,N_28634);
nand U31649 (N_31649,N_28928,N_28634);
or U31650 (N_31650,N_28008,N_28395);
nand U31651 (N_31651,N_28388,N_28282);
and U31652 (N_31652,N_29744,N_28263);
and U31653 (N_31653,N_29810,N_28284);
xor U31654 (N_31654,N_29380,N_29587);
or U31655 (N_31655,N_28039,N_29728);
nand U31656 (N_31656,N_28121,N_28188);
nand U31657 (N_31657,N_29397,N_29956);
nor U31658 (N_31658,N_28333,N_28526);
nand U31659 (N_31659,N_28853,N_28428);
and U31660 (N_31660,N_29414,N_29208);
or U31661 (N_31661,N_28833,N_29357);
xnor U31662 (N_31662,N_28986,N_28805);
and U31663 (N_31663,N_28598,N_29200);
nor U31664 (N_31664,N_28186,N_28583);
or U31665 (N_31665,N_29232,N_28497);
nor U31666 (N_31666,N_28770,N_29598);
or U31667 (N_31667,N_29843,N_28876);
nand U31668 (N_31668,N_29515,N_28650);
xor U31669 (N_31669,N_28884,N_29600);
xnor U31670 (N_31670,N_29764,N_29448);
and U31671 (N_31671,N_29077,N_29171);
nand U31672 (N_31672,N_29503,N_28256);
nor U31673 (N_31673,N_29817,N_28749);
nand U31674 (N_31674,N_29655,N_28552);
nand U31675 (N_31675,N_28885,N_28468);
and U31676 (N_31676,N_28312,N_29317);
xnor U31677 (N_31677,N_28383,N_29763);
and U31678 (N_31678,N_28710,N_28284);
nor U31679 (N_31679,N_28823,N_28727);
xnor U31680 (N_31680,N_29389,N_29310);
nand U31681 (N_31681,N_28020,N_29496);
nor U31682 (N_31682,N_29637,N_28352);
nor U31683 (N_31683,N_29263,N_28619);
or U31684 (N_31684,N_29872,N_28721);
xor U31685 (N_31685,N_28053,N_29297);
nor U31686 (N_31686,N_28914,N_28283);
or U31687 (N_31687,N_28499,N_29576);
or U31688 (N_31688,N_28294,N_28105);
nand U31689 (N_31689,N_29931,N_29007);
or U31690 (N_31690,N_28213,N_28281);
nor U31691 (N_31691,N_28198,N_28901);
nor U31692 (N_31692,N_28700,N_28502);
xnor U31693 (N_31693,N_29648,N_28600);
or U31694 (N_31694,N_28844,N_29658);
nor U31695 (N_31695,N_29710,N_28301);
or U31696 (N_31696,N_29689,N_28879);
and U31697 (N_31697,N_28556,N_28360);
or U31698 (N_31698,N_28791,N_28956);
nor U31699 (N_31699,N_29516,N_28701);
nor U31700 (N_31700,N_29460,N_29261);
xnor U31701 (N_31701,N_29863,N_28778);
and U31702 (N_31702,N_29909,N_29949);
and U31703 (N_31703,N_28312,N_29921);
nor U31704 (N_31704,N_28502,N_29858);
xor U31705 (N_31705,N_28826,N_29860);
or U31706 (N_31706,N_28802,N_29258);
and U31707 (N_31707,N_28073,N_28832);
nor U31708 (N_31708,N_28559,N_28804);
or U31709 (N_31709,N_28984,N_29290);
and U31710 (N_31710,N_28396,N_29065);
xor U31711 (N_31711,N_28413,N_28326);
nand U31712 (N_31712,N_29940,N_28443);
xor U31713 (N_31713,N_29050,N_28441);
and U31714 (N_31714,N_28307,N_28399);
nand U31715 (N_31715,N_28344,N_28007);
nor U31716 (N_31716,N_29436,N_29171);
and U31717 (N_31717,N_28906,N_29312);
nand U31718 (N_31718,N_28851,N_29138);
xor U31719 (N_31719,N_28182,N_28812);
and U31720 (N_31720,N_29696,N_28820);
or U31721 (N_31721,N_28444,N_28518);
nand U31722 (N_31722,N_28048,N_28725);
xor U31723 (N_31723,N_28152,N_29198);
nand U31724 (N_31724,N_28899,N_28054);
and U31725 (N_31725,N_28723,N_29175);
and U31726 (N_31726,N_29544,N_29221);
and U31727 (N_31727,N_29078,N_28109);
nor U31728 (N_31728,N_28092,N_29544);
and U31729 (N_31729,N_28399,N_28637);
nand U31730 (N_31730,N_28460,N_29305);
or U31731 (N_31731,N_29191,N_29360);
nand U31732 (N_31732,N_29126,N_28608);
nor U31733 (N_31733,N_29194,N_29580);
and U31734 (N_31734,N_29679,N_28117);
nand U31735 (N_31735,N_28713,N_29315);
xnor U31736 (N_31736,N_29316,N_28344);
and U31737 (N_31737,N_29845,N_29617);
and U31738 (N_31738,N_28808,N_28265);
or U31739 (N_31739,N_28008,N_28758);
xnor U31740 (N_31740,N_28396,N_29293);
nand U31741 (N_31741,N_29789,N_28599);
or U31742 (N_31742,N_28730,N_28835);
nor U31743 (N_31743,N_28651,N_28497);
and U31744 (N_31744,N_29431,N_28427);
nand U31745 (N_31745,N_28283,N_29836);
nor U31746 (N_31746,N_28853,N_29619);
and U31747 (N_31747,N_28612,N_28958);
and U31748 (N_31748,N_29520,N_28097);
or U31749 (N_31749,N_28080,N_29339);
or U31750 (N_31750,N_29271,N_28807);
or U31751 (N_31751,N_28255,N_28449);
xor U31752 (N_31752,N_29203,N_28896);
nor U31753 (N_31753,N_29196,N_29950);
nor U31754 (N_31754,N_29550,N_28562);
nor U31755 (N_31755,N_28423,N_29550);
nor U31756 (N_31756,N_29137,N_28125);
xnor U31757 (N_31757,N_28066,N_29327);
xor U31758 (N_31758,N_28416,N_28128);
and U31759 (N_31759,N_28552,N_29769);
xnor U31760 (N_31760,N_29360,N_28521);
and U31761 (N_31761,N_28899,N_29833);
and U31762 (N_31762,N_28044,N_29399);
nand U31763 (N_31763,N_28662,N_29212);
nor U31764 (N_31764,N_28804,N_28896);
or U31765 (N_31765,N_29051,N_28821);
xnor U31766 (N_31766,N_29514,N_28475);
and U31767 (N_31767,N_28350,N_28643);
nand U31768 (N_31768,N_29018,N_28386);
xor U31769 (N_31769,N_28658,N_28386);
or U31770 (N_31770,N_28059,N_28167);
nand U31771 (N_31771,N_28870,N_28609);
nand U31772 (N_31772,N_29423,N_29292);
or U31773 (N_31773,N_29189,N_28113);
or U31774 (N_31774,N_29313,N_28546);
and U31775 (N_31775,N_28032,N_29411);
xnor U31776 (N_31776,N_28680,N_28247);
and U31777 (N_31777,N_28922,N_28510);
xnor U31778 (N_31778,N_29080,N_29092);
and U31779 (N_31779,N_28897,N_28396);
and U31780 (N_31780,N_28829,N_29571);
and U31781 (N_31781,N_29444,N_28259);
and U31782 (N_31782,N_28220,N_29289);
nand U31783 (N_31783,N_29658,N_28853);
nand U31784 (N_31784,N_28203,N_28082);
xnor U31785 (N_31785,N_29309,N_28717);
or U31786 (N_31786,N_29311,N_29156);
and U31787 (N_31787,N_28243,N_29107);
xnor U31788 (N_31788,N_29293,N_28438);
nor U31789 (N_31789,N_29961,N_29295);
and U31790 (N_31790,N_28428,N_28371);
and U31791 (N_31791,N_29775,N_28571);
nor U31792 (N_31792,N_28629,N_29816);
and U31793 (N_31793,N_28482,N_29263);
and U31794 (N_31794,N_28323,N_29691);
or U31795 (N_31795,N_28144,N_28696);
xor U31796 (N_31796,N_28831,N_29753);
or U31797 (N_31797,N_28482,N_28334);
and U31798 (N_31798,N_29990,N_29256);
and U31799 (N_31799,N_28205,N_29506);
and U31800 (N_31800,N_28319,N_29285);
and U31801 (N_31801,N_28132,N_28012);
nor U31802 (N_31802,N_29131,N_28627);
and U31803 (N_31803,N_29046,N_29898);
nand U31804 (N_31804,N_28231,N_29747);
and U31805 (N_31805,N_29634,N_28695);
xnor U31806 (N_31806,N_28067,N_29497);
nand U31807 (N_31807,N_28873,N_28890);
nand U31808 (N_31808,N_28038,N_28587);
nand U31809 (N_31809,N_29069,N_29235);
or U31810 (N_31810,N_29912,N_28649);
nor U31811 (N_31811,N_28357,N_28876);
nor U31812 (N_31812,N_29704,N_28961);
nand U31813 (N_31813,N_28604,N_28420);
nor U31814 (N_31814,N_29700,N_28870);
or U31815 (N_31815,N_29287,N_29550);
nand U31816 (N_31816,N_28180,N_28850);
nand U31817 (N_31817,N_28546,N_29899);
nand U31818 (N_31818,N_28460,N_28235);
nor U31819 (N_31819,N_28286,N_29703);
and U31820 (N_31820,N_28840,N_28857);
or U31821 (N_31821,N_28590,N_28836);
and U31822 (N_31822,N_28280,N_28908);
nand U31823 (N_31823,N_29845,N_29145);
and U31824 (N_31824,N_29825,N_28438);
nand U31825 (N_31825,N_29366,N_29621);
nand U31826 (N_31826,N_29625,N_29089);
and U31827 (N_31827,N_29872,N_29524);
xnor U31828 (N_31828,N_29873,N_29952);
nand U31829 (N_31829,N_28984,N_29533);
nand U31830 (N_31830,N_28487,N_28250);
and U31831 (N_31831,N_29098,N_29454);
xor U31832 (N_31832,N_28712,N_28861);
xnor U31833 (N_31833,N_29196,N_28282);
nand U31834 (N_31834,N_29664,N_28724);
nor U31835 (N_31835,N_29310,N_29726);
or U31836 (N_31836,N_29525,N_28193);
nor U31837 (N_31837,N_29311,N_28908);
nand U31838 (N_31838,N_29492,N_28418);
and U31839 (N_31839,N_29691,N_29510);
or U31840 (N_31840,N_29453,N_28764);
xnor U31841 (N_31841,N_29479,N_29729);
nand U31842 (N_31842,N_29547,N_29635);
or U31843 (N_31843,N_29538,N_29461);
and U31844 (N_31844,N_28588,N_28675);
nand U31845 (N_31845,N_29467,N_29721);
nor U31846 (N_31846,N_28099,N_28683);
nand U31847 (N_31847,N_29160,N_29955);
and U31848 (N_31848,N_29003,N_29373);
and U31849 (N_31849,N_29310,N_29702);
nand U31850 (N_31850,N_29966,N_28742);
nor U31851 (N_31851,N_28074,N_29665);
xnor U31852 (N_31852,N_29377,N_28882);
and U31853 (N_31853,N_28788,N_29703);
or U31854 (N_31854,N_29344,N_28742);
nor U31855 (N_31855,N_29271,N_29363);
nand U31856 (N_31856,N_28907,N_28138);
nor U31857 (N_31857,N_28207,N_29484);
xnor U31858 (N_31858,N_29847,N_28540);
xor U31859 (N_31859,N_28857,N_29252);
nor U31860 (N_31860,N_28861,N_28336);
xor U31861 (N_31861,N_28900,N_29696);
xnor U31862 (N_31862,N_29754,N_28718);
nor U31863 (N_31863,N_29608,N_29538);
nor U31864 (N_31864,N_29208,N_28157);
nand U31865 (N_31865,N_28055,N_29597);
nand U31866 (N_31866,N_28667,N_29671);
or U31867 (N_31867,N_28155,N_29897);
or U31868 (N_31868,N_29033,N_28135);
nand U31869 (N_31869,N_28485,N_29887);
xnor U31870 (N_31870,N_28857,N_29027);
or U31871 (N_31871,N_29489,N_29654);
or U31872 (N_31872,N_28439,N_29266);
nor U31873 (N_31873,N_28685,N_29034);
xor U31874 (N_31874,N_29391,N_29362);
or U31875 (N_31875,N_28489,N_29088);
and U31876 (N_31876,N_28070,N_28008);
and U31877 (N_31877,N_28204,N_29436);
xor U31878 (N_31878,N_28969,N_28505);
xor U31879 (N_31879,N_29608,N_29533);
or U31880 (N_31880,N_29328,N_28449);
nand U31881 (N_31881,N_29076,N_28774);
nand U31882 (N_31882,N_28464,N_29913);
xor U31883 (N_31883,N_29787,N_29134);
nor U31884 (N_31884,N_29371,N_29921);
nand U31885 (N_31885,N_28315,N_29813);
xor U31886 (N_31886,N_28823,N_28336);
xnor U31887 (N_31887,N_29893,N_29087);
nor U31888 (N_31888,N_28389,N_29272);
xnor U31889 (N_31889,N_29597,N_29060);
xnor U31890 (N_31890,N_29720,N_29717);
nor U31891 (N_31891,N_28397,N_28190);
xor U31892 (N_31892,N_29967,N_29691);
and U31893 (N_31893,N_28807,N_29654);
xor U31894 (N_31894,N_29222,N_28104);
xor U31895 (N_31895,N_28576,N_28162);
or U31896 (N_31896,N_28768,N_29969);
nor U31897 (N_31897,N_29813,N_28330);
nand U31898 (N_31898,N_29029,N_29313);
nand U31899 (N_31899,N_29220,N_28915);
nor U31900 (N_31900,N_29054,N_29909);
and U31901 (N_31901,N_29095,N_29140);
xnor U31902 (N_31902,N_29722,N_28591);
nand U31903 (N_31903,N_28020,N_28353);
and U31904 (N_31904,N_28316,N_28381);
or U31905 (N_31905,N_28666,N_28036);
and U31906 (N_31906,N_28753,N_29255);
and U31907 (N_31907,N_29857,N_29346);
nand U31908 (N_31908,N_28210,N_29819);
nor U31909 (N_31909,N_29731,N_29143);
and U31910 (N_31910,N_29976,N_29616);
nor U31911 (N_31911,N_29142,N_29617);
nor U31912 (N_31912,N_28839,N_28243);
nor U31913 (N_31913,N_29898,N_28997);
xor U31914 (N_31914,N_29718,N_28046);
or U31915 (N_31915,N_29792,N_29554);
and U31916 (N_31916,N_29373,N_28066);
xnor U31917 (N_31917,N_29989,N_29194);
and U31918 (N_31918,N_28631,N_29064);
xnor U31919 (N_31919,N_29919,N_28612);
xnor U31920 (N_31920,N_28610,N_29572);
or U31921 (N_31921,N_29007,N_28302);
nand U31922 (N_31922,N_29453,N_29462);
nor U31923 (N_31923,N_28350,N_28440);
nand U31924 (N_31924,N_28066,N_29446);
nor U31925 (N_31925,N_28752,N_28458);
or U31926 (N_31926,N_28985,N_28877);
or U31927 (N_31927,N_28643,N_28446);
nand U31928 (N_31928,N_29952,N_28524);
and U31929 (N_31929,N_28815,N_29509);
and U31930 (N_31930,N_29076,N_29984);
and U31931 (N_31931,N_29616,N_28451);
xnor U31932 (N_31932,N_28240,N_29304);
or U31933 (N_31933,N_29202,N_29585);
nor U31934 (N_31934,N_28606,N_29955);
xnor U31935 (N_31935,N_28997,N_29985);
nand U31936 (N_31936,N_29099,N_29974);
or U31937 (N_31937,N_29587,N_29090);
nand U31938 (N_31938,N_28761,N_29096);
xor U31939 (N_31939,N_29480,N_28245);
and U31940 (N_31940,N_29435,N_28578);
or U31941 (N_31941,N_29020,N_29284);
nand U31942 (N_31942,N_28112,N_28275);
and U31943 (N_31943,N_28359,N_29468);
nand U31944 (N_31944,N_29030,N_28557);
or U31945 (N_31945,N_28761,N_29552);
or U31946 (N_31946,N_29721,N_28780);
and U31947 (N_31947,N_29878,N_28978);
or U31948 (N_31948,N_28950,N_28962);
or U31949 (N_31949,N_28084,N_29559);
or U31950 (N_31950,N_29858,N_28446);
nand U31951 (N_31951,N_29525,N_28537);
nor U31952 (N_31952,N_28229,N_29344);
nand U31953 (N_31953,N_28334,N_28978);
or U31954 (N_31954,N_29805,N_29954);
xor U31955 (N_31955,N_29942,N_29808);
nand U31956 (N_31956,N_28474,N_28293);
xnor U31957 (N_31957,N_28783,N_29713);
and U31958 (N_31958,N_29372,N_28825);
or U31959 (N_31959,N_29939,N_29620);
or U31960 (N_31960,N_28624,N_28826);
xor U31961 (N_31961,N_29125,N_29991);
nand U31962 (N_31962,N_29985,N_29717);
xnor U31963 (N_31963,N_29452,N_28193);
and U31964 (N_31964,N_29569,N_28757);
nand U31965 (N_31965,N_28313,N_29136);
nor U31966 (N_31966,N_29393,N_28121);
xor U31967 (N_31967,N_28376,N_28213);
and U31968 (N_31968,N_28361,N_28071);
nand U31969 (N_31969,N_28325,N_29844);
nand U31970 (N_31970,N_29921,N_28253);
nand U31971 (N_31971,N_28892,N_29083);
and U31972 (N_31972,N_28542,N_29794);
or U31973 (N_31973,N_29355,N_29327);
and U31974 (N_31974,N_29011,N_29292);
xnor U31975 (N_31975,N_28328,N_29125);
nor U31976 (N_31976,N_28345,N_29511);
and U31977 (N_31977,N_28861,N_29376);
and U31978 (N_31978,N_28453,N_29032);
nor U31979 (N_31979,N_28781,N_29968);
and U31980 (N_31980,N_29569,N_29914);
nor U31981 (N_31981,N_28490,N_29178);
xnor U31982 (N_31982,N_28035,N_29950);
nand U31983 (N_31983,N_28972,N_29232);
nor U31984 (N_31984,N_28763,N_29112);
xnor U31985 (N_31985,N_29251,N_28136);
xnor U31986 (N_31986,N_29230,N_28164);
nand U31987 (N_31987,N_29764,N_28733);
xor U31988 (N_31988,N_29705,N_28565);
and U31989 (N_31989,N_28833,N_28852);
or U31990 (N_31990,N_29267,N_29543);
and U31991 (N_31991,N_28540,N_29688);
nor U31992 (N_31992,N_29299,N_29792);
or U31993 (N_31993,N_28554,N_28520);
nor U31994 (N_31994,N_28739,N_28955);
or U31995 (N_31995,N_29031,N_28866);
nand U31996 (N_31996,N_29142,N_29134);
nand U31997 (N_31997,N_29576,N_28042);
and U31998 (N_31998,N_28740,N_29058);
xor U31999 (N_31999,N_29880,N_28282);
xnor U32000 (N_32000,N_30882,N_30852);
and U32001 (N_32001,N_31788,N_30503);
xor U32002 (N_32002,N_30556,N_30025);
xor U32003 (N_32003,N_31947,N_31769);
or U32004 (N_32004,N_30703,N_31503);
nand U32005 (N_32005,N_31349,N_30416);
nand U32006 (N_32006,N_31814,N_30599);
nor U32007 (N_32007,N_30821,N_31168);
or U32008 (N_32008,N_30762,N_31583);
or U32009 (N_32009,N_30245,N_31823);
xor U32010 (N_32010,N_30452,N_31596);
or U32011 (N_32011,N_30621,N_31079);
xnor U32012 (N_32012,N_30458,N_31341);
nor U32013 (N_32013,N_30966,N_31157);
and U32014 (N_32014,N_30205,N_30941);
and U32015 (N_32015,N_31226,N_30402);
xnor U32016 (N_32016,N_31254,N_31830);
nand U32017 (N_32017,N_30430,N_31277);
and U32018 (N_32018,N_31003,N_31749);
xnor U32019 (N_32019,N_30020,N_31574);
and U32020 (N_32020,N_30252,N_31203);
xor U32021 (N_32021,N_30925,N_31722);
xnor U32022 (N_32022,N_30275,N_30758);
nand U32023 (N_32023,N_31452,N_31494);
and U32024 (N_32024,N_31888,N_30360);
or U32025 (N_32025,N_31819,N_31197);
nor U32026 (N_32026,N_31031,N_31979);
nor U32027 (N_32027,N_31694,N_31380);
nand U32028 (N_32028,N_31971,N_30604);
nor U32029 (N_32029,N_31133,N_30667);
nand U32030 (N_32030,N_31711,N_31478);
nor U32031 (N_32031,N_30792,N_31643);
nand U32032 (N_32032,N_30432,N_31018);
nand U32033 (N_32033,N_30435,N_31198);
nand U32034 (N_32034,N_30346,N_30746);
xor U32035 (N_32035,N_31850,N_31662);
nand U32036 (N_32036,N_30831,N_31153);
or U32037 (N_32037,N_30104,N_31060);
nand U32038 (N_32038,N_31042,N_30612);
nor U32039 (N_32039,N_30166,N_30548);
nand U32040 (N_32040,N_31086,N_31732);
xor U32041 (N_32041,N_31316,N_30763);
nand U32042 (N_32042,N_31860,N_31354);
xnor U32043 (N_32043,N_31172,N_30456);
xnor U32044 (N_32044,N_30133,N_31450);
xor U32045 (N_32045,N_31324,N_30158);
nand U32046 (N_32046,N_31024,N_31783);
xnor U32047 (N_32047,N_31631,N_30135);
or U32048 (N_32048,N_31713,N_30847);
or U32049 (N_32049,N_30980,N_30915);
nor U32050 (N_32050,N_31963,N_30454);
or U32051 (N_32051,N_30640,N_31136);
xor U32052 (N_32052,N_30944,N_30487);
nand U32053 (N_32053,N_30871,N_30991);
nor U32054 (N_32054,N_30415,N_31671);
nand U32055 (N_32055,N_31855,N_30839);
and U32056 (N_32056,N_31960,N_30339);
xor U32057 (N_32057,N_31539,N_30564);
xor U32058 (N_32058,N_30325,N_31233);
and U32059 (N_32059,N_30068,N_31798);
or U32060 (N_32060,N_30560,N_30884);
nor U32061 (N_32061,N_30835,N_31650);
xor U32062 (N_32062,N_30265,N_31497);
nor U32063 (N_32063,N_30397,N_31999);
nand U32064 (N_32064,N_30668,N_31384);
nor U32065 (N_32065,N_31106,N_30192);
nand U32066 (N_32066,N_30094,N_31771);
or U32067 (N_32067,N_30529,N_30506);
nand U32068 (N_32068,N_31074,N_31718);
and U32069 (N_32069,N_31289,N_31614);
nand U32070 (N_32070,N_31842,N_31400);
or U32071 (N_32071,N_31177,N_31518);
and U32072 (N_32072,N_31087,N_31459);
nor U32073 (N_32073,N_30127,N_30679);
nor U32074 (N_32074,N_31707,N_31760);
nor U32075 (N_32075,N_31209,N_30664);
xor U32076 (N_32076,N_31689,N_31190);
or U32077 (N_32077,N_30954,N_30536);
or U32078 (N_32078,N_31591,N_31890);
xor U32079 (N_32079,N_31602,N_31525);
nand U32080 (N_32080,N_30008,N_31049);
or U32081 (N_32081,N_30616,N_31192);
and U32082 (N_32082,N_31682,N_31223);
nor U32083 (N_32083,N_31791,N_30311);
nor U32084 (N_32084,N_31430,N_31826);
and U32085 (N_32085,N_31986,N_31550);
nor U32086 (N_32086,N_30894,N_31144);
xnor U32087 (N_32087,N_31010,N_30651);
and U32088 (N_32088,N_31683,N_30421);
xnor U32089 (N_32089,N_31364,N_30708);
xor U32090 (N_32090,N_31931,N_30394);
nor U32091 (N_32091,N_30748,N_31693);
or U32092 (N_32092,N_30910,N_31121);
or U32093 (N_32093,N_30331,N_31975);
or U32094 (N_32094,N_30182,N_31978);
nand U32095 (N_32095,N_31323,N_31204);
xnor U32096 (N_32096,N_30371,N_31340);
nand U32097 (N_32097,N_31005,N_30555);
nor U32098 (N_32098,N_31951,N_30934);
xor U32099 (N_32099,N_30255,N_31943);
xnor U32100 (N_32100,N_30964,N_31734);
xnor U32101 (N_32101,N_30507,N_30856);
nor U32102 (N_32102,N_31259,N_30030);
nor U32103 (N_32103,N_31758,N_31556);
xnor U32104 (N_32104,N_30544,N_31363);
nor U32105 (N_32105,N_30519,N_31582);
nand U32106 (N_32106,N_31044,N_31577);
nor U32107 (N_32107,N_31280,N_31426);
nor U32108 (N_32108,N_30411,N_30408);
nand U32109 (N_32109,N_30515,N_30911);
and U32110 (N_32110,N_31211,N_31174);
and U32111 (N_32111,N_30033,N_31627);
and U32112 (N_32112,N_31716,N_30422);
nand U32113 (N_32113,N_30726,N_31269);
or U32114 (N_32114,N_30368,N_30801);
or U32115 (N_32115,N_31398,N_30681);
or U32116 (N_32116,N_30053,N_30330);
nand U32117 (N_32117,N_31064,N_31606);
xnor U32118 (N_32118,N_30419,N_31976);
or U32119 (N_32119,N_30052,N_31942);
and U32120 (N_32120,N_31187,N_31275);
nor U32121 (N_32121,N_31628,N_31148);
and U32122 (N_32122,N_31498,N_31592);
and U32123 (N_32123,N_31970,N_30671);
or U32124 (N_32124,N_31433,N_30957);
nor U32125 (N_32125,N_30753,N_30993);
and U32126 (N_32126,N_31102,N_31792);
nor U32127 (N_32127,N_30550,N_31623);
xor U32128 (N_32128,N_30736,N_31502);
or U32129 (N_32129,N_30822,N_31131);
nand U32130 (N_32130,N_31481,N_30573);
or U32131 (N_32131,N_30404,N_31376);
nand U32132 (N_32132,N_31762,N_30596);
nand U32133 (N_32133,N_31117,N_31572);
nand U32134 (N_32134,N_31950,N_30752);
or U32135 (N_32135,N_30782,N_30140);
and U32136 (N_32136,N_31569,N_31507);
nor U32137 (N_32137,N_31167,N_30409);
nor U32138 (N_32138,N_31446,N_30778);
xnor U32139 (N_32139,N_31506,N_30885);
nand U32140 (N_32140,N_31490,N_30049);
nor U32141 (N_32141,N_31253,N_31917);
or U32142 (N_32142,N_31270,N_31404);
nand U32143 (N_32143,N_30018,N_30460);
and U32144 (N_32144,N_31441,N_30994);
nor U32145 (N_32145,N_30222,N_30563);
nor U32146 (N_32146,N_30069,N_31797);
or U32147 (N_32147,N_31753,N_30654);
or U32148 (N_32148,N_30465,N_30321);
nor U32149 (N_32149,N_30179,N_31138);
and U32150 (N_32150,N_30355,N_30986);
and U32151 (N_32151,N_30526,N_31879);
or U32152 (N_32152,N_30656,N_31368);
nor U32153 (N_32153,N_31006,N_30308);
nor U32154 (N_32154,N_30795,N_30844);
nand U32155 (N_32155,N_30716,N_30825);
nor U32156 (N_32156,N_31093,N_31073);
or U32157 (N_32157,N_31048,N_30082);
xor U32158 (N_32158,N_31822,N_31229);
xor U32159 (N_32159,N_31900,N_31742);
nand U32160 (N_32160,N_31526,N_31184);
nor U32161 (N_32161,N_30388,N_30491);
nand U32162 (N_32162,N_30619,N_31670);
and U32163 (N_32163,N_30953,N_31181);
nor U32164 (N_32164,N_31059,N_31756);
nand U32165 (N_32165,N_30974,N_31486);
or U32166 (N_32166,N_31660,N_31540);
or U32167 (N_32167,N_30976,N_30171);
nor U32168 (N_32168,N_31081,N_30072);
or U32169 (N_32169,N_30783,N_30260);
or U32170 (N_32170,N_30400,N_31183);
or U32171 (N_32171,N_30862,N_31436);
xor U32172 (N_32172,N_30985,N_30493);
nand U32173 (N_32173,N_31315,N_31821);
and U32174 (N_32174,N_30023,N_31968);
nor U32175 (N_32175,N_31206,N_30376);
nor U32176 (N_32176,N_31479,N_31065);
and U32177 (N_32177,N_30223,N_31448);
xnor U32178 (N_32178,N_30733,N_31794);
nand U32179 (N_32179,N_31688,N_30144);
xnor U32180 (N_32180,N_30786,N_31719);
or U32181 (N_32181,N_31695,N_31043);
or U32182 (N_32182,N_30730,N_30863);
nor U32183 (N_32183,N_31657,N_31553);
or U32184 (N_32184,N_30276,N_31317);
nor U32185 (N_32185,N_30324,N_30424);
nor U32186 (N_32186,N_30605,N_31300);
nand U32187 (N_32187,N_31234,N_30901);
nand U32188 (N_32188,N_31487,N_31112);
and U32189 (N_32189,N_30684,N_30745);
xor U32190 (N_32190,N_30955,N_30567);
nand U32191 (N_32191,N_31263,N_30113);
and U32192 (N_32192,N_31748,N_31170);
or U32193 (N_32193,N_31122,N_30216);
and U32194 (N_32194,N_31562,N_31098);
and U32195 (N_32195,N_30129,N_30879);
or U32196 (N_32196,N_30317,N_31374);
nor U32197 (N_32197,N_30921,N_30010);
and U32198 (N_32198,N_30765,N_30546);
nor U32199 (N_32199,N_31777,N_31243);
and U32200 (N_32200,N_30772,N_30288);
or U32201 (N_32201,N_30187,N_31213);
and U32202 (N_32202,N_31913,N_30774);
xor U32203 (N_32203,N_31790,N_31033);
nor U32204 (N_32204,N_30836,N_31366);
or U32205 (N_32205,N_30717,N_31731);
or U32206 (N_32206,N_31442,N_30084);
nor U32207 (N_32207,N_31451,N_31130);
or U32208 (N_32208,N_31186,N_30157);
and U32209 (N_32209,N_31840,N_31035);
nand U32210 (N_32210,N_31207,N_30039);
xnor U32211 (N_32211,N_30741,N_30568);
nand U32212 (N_32212,N_31573,N_31952);
and U32213 (N_32213,N_30429,N_30273);
and U32214 (N_32214,N_30942,N_31641);
or U32215 (N_32215,N_31500,N_30749);
nor U32216 (N_32216,N_30309,N_30410);
xor U32217 (N_32217,N_30969,N_30649);
xor U32218 (N_32218,N_30480,N_31558);
or U32219 (N_32219,N_31360,N_30470);
or U32220 (N_32220,N_30302,N_31397);
and U32221 (N_32221,N_31899,N_31767);
or U32222 (N_32222,N_31648,N_31140);
or U32223 (N_32223,N_30575,N_31861);
nor U32224 (N_32224,N_31754,N_30789);
or U32225 (N_32225,N_31841,N_31954);
nor U32226 (N_32226,N_30472,N_30982);
nand U32227 (N_32227,N_30665,N_30221);
xnor U32228 (N_32228,N_30202,N_30439);
or U32229 (N_32229,N_30074,N_30455);
or U32230 (N_32230,N_30562,N_31402);
nor U32231 (N_32231,N_30577,N_30532);
xnor U32232 (N_32232,N_31630,N_30414);
or U32233 (N_32233,N_31563,N_30670);
nand U32234 (N_32234,N_31661,N_31414);
xor U32235 (N_32235,N_31394,N_30070);
and U32236 (N_32236,N_31845,N_30678);
and U32237 (N_32237,N_30357,N_30866);
nand U32238 (N_32238,N_31178,N_31428);
nor U32239 (N_32239,N_30636,N_30370);
nor U32240 (N_32240,N_30254,N_30057);
nand U32241 (N_32241,N_31373,N_31745);
xnor U32242 (N_32242,N_31029,N_31825);
and U32243 (N_32243,N_30677,N_31405);
and U32244 (N_32244,N_31217,N_30541);
xnor U32245 (N_32245,N_31482,N_31417);
nor U32246 (N_32246,N_30248,N_31094);
nand U32247 (N_32247,N_31761,N_31709);
nand U32248 (N_32248,N_31145,N_31396);
nor U32249 (N_32249,N_31313,N_30860);
xor U32250 (N_32250,N_31907,N_31422);
xor U32251 (N_32251,N_31835,N_31246);
nand U32252 (N_32252,N_31240,N_31389);
nand U32253 (N_32253,N_30501,N_31371);
nor U32254 (N_32254,N_30201,N_30586);
or U32255 (N_32255,N_31938,N_30600);
nor U32256 (N_32256,N_31132,N_31222);
and U32257 (N_32257,N_30285,N_31116);
nand U32258 (N_32258,N_30294,N_31342);
nand U32259 (N_32259,N_30119,N_30055);
xnor U32260 (N_32260,N_31001,N_31714);
and U32261 (N_32261,N_30322,N_31423);
nor U32262 (N_32262,N_31723,N_30891);
nor U32263 (N_32263,N_31291,N_30431);
and U32264 (N_32264,N_31629,N_30781);
nor U32265 (N_32265,N_30706,N_31485);
and U32266 (N_32266,N_31166,N_30939);
xor U32267 (N_32267,N_30881,N_30261);
nor U32268 (N_32268,N_30642,N_30184);
nand U32269 (N_32269,N_31169,N_31182);
xnor U32270 (N_32270,N_30130,N_30534);
nor U32271 (N_32271,N_30992,N_31815);
nor U32272 (N_32272,N_30334,N_31311);
and U32273 (N_32273,N_30219,N_31336);
and U32274 (N_32274,N_31864,N_31058);
and U32275 (N_32275,N_30851,N_30947);
or U32276 (N_32276,N_31961,N_31295);
and U32277 (N_32277,N_30352,N_30466);
nand U32278 (N_32278,N_31128,N_30138);
nor U32279 (N_32279,N_31196,N_30029);
xor U32280 (N_32280,N_30510,N_30811);
nor U32281 (N_32281,N_31070,N_31915);
nand U32282 (N_32282,N_30843,N_31524);
xnor U32283 (N_32283,N_31296,N_30554);
xor U32284 (N_32284,N_30676,N_30436);
and U32285 (N_32285,N_31989,N_30278);
and U32286 (N_32286,N_31047,N_30858);
or U32287 (N_32287,N_31504,N_30806);
and U32288 (N_32288,N_30926,N_30191);
nor U32289 (N_32289,N_31877,N_30481);
xnor U32290 (N_32290,N_30511,N_31036);
nor U32291 (N_32291,N_30613,N_30213);
and U32292 (N_32292,N_31472,N_30837);
nand U32293 (N_32293,N_30732,N_31322);
nand U32294 (N_32294,N_30167,N_31774);
nand U32295 (N_32295,N_31530,N_30034);
nand U32296 (N_32296,N_31611,N_30338);
or U32297 (N_32297,N_30373,N_30079);
xnor U32298 (N_32298,N_31383,N_31655);
or U32299 (N_32299,N_30141,N_31355);
or U32300 (N_32300,N_31514,N_31063);
nor U32301 (N_32301,N_31164,N_30405);
and U32302 (N_32302,N_31692,N_30485);
nor U32303 (N_32303,N_31729,N_31773);
nor U32304 (N_32304,N_31370,N_31956);
nor U32305 (N_32305,N_30139,N_30464);
and U32306 (N_32306,N_31759,N_30151);
and U32307 (N_32307,N_31772,N_31066);
and U32308 (N_32308,N_30146,N_30614);
and U32309 (N_32309,N_30242,N_30241);
nand U32310 (N_32310,N_30272,N_30282);
xnor U32311 (N_32311,N_30794,N_31235);
nand U32312 (N_32312,N_31257,N_31134);
xor U32313 (N_32313,N_31244,N_31546);
or U32314 (N_32314,N_30112,N_31410);
xor U32315 (N_32315,N_30697,N_31896);
nor U32316 (N_32316,N_31785,N_30785);
xor U32317 (N_32317,N_30583,N_31260);
and U32318 (N_32318,N_30951,N_30022);
and U32319 (N_32319,N_30027,N_30335);
xor U32320 (N_32320,N_31706,N_31740);
nor U32321 (N_32321,N_31320,N_30854);
nand U32322 (N_32322,N_30313,N_30528);
or U32323 (N_32323,N_30423,N_31118);
nand U32324 (N_32324,N_30395,N_31529);
nand U32325 (N_32325,N_31028,N_31054);
or U32326 (N_32326,N_31510,N_31496);
nand U32327 (N_32327,N_31571,N_31467);
or U32328 (N_32328,N_31113,N_31843);
and U32329 (N_32329,N_30631,N_30489);
nand U32330 (N_32330,N_31356,N_30912);
nand U32331 (N_32331,N_31610,N_31050);
nand U32332 (N_32332,N_31266,N_31594);
nand U32333 (N_32333,N_30087,N_31541);
and U32334 (N_32334,N_30592,N_31549);
and U32335 (N_32335,N_30900,N_30253);
or U32336 (N_32336,N_30212,N_31664);
or U32337 (N_32337,N_30152,N_30938);
nor U32338 (N_32338,N_30551,N_30341);
and U32339 (N_32339,N_31807,N_30374);
nand U32340 (N_32340,N_30169,N_31836);
nor U32341 (N_32341,N_31221,N_31666);
nor U32342 (N_32342,N_30380,N_30078);
nand U32343 (N_32343,N_30204,N_30249);
nor U32344 (N_32344,N_31232,N_30919);
nand U32345 (N_32345,N_30597,N_30005);
nor U32346 (N_32346,N_31161,N_31250);
nor U32347 (N_32347,N_30952,N_31651);
nor U32348 (N_32348,N_31897,N_30977);
nand U32349 (N_32349,N_31421,N_31002);
nor U32350 (N_32350,N_30398,N_31511);
nand U32351 (N_32351,N_31957,N_30658);
nor U32352 (N_32352,N_31332,N_30093);
and U32353 (N_32353,N_30271,N_30088);
nand U32354 (N_32354,N_30494,N_31016);
and U32355 (N_32355,N_30496,N_30476);
nor U32356 (N_32356,N_31810,N_30530);
nand U32357 (N_32357,N_31616,N_30516);
nor U32358 (N_32358,N_30342,N_30343);
nor U32359 (N_32359,N_30156,N_31365);
or U32360 (N_32360,N_31447,N_30561);
or U32361 (N_32361,N_31634,N_31534);
xor U32362 (N_32362,N_31252,N_30890);
or U32363 (N_32363,N_30389,N_30707);
xnor U32364 (N_32364,N_31012,N_30788);
and U32365 (N_32365,N_30488,N_31267);
nand U32366 (N_32366,N_31918,N_31652);
and U32367 (N_32367,N_31939,N_30666);
and U32368 (N_32368,N_31101,N_30645);
nor U32369 (N_32369,N_30114,N_31361);
and U32370 (N_32370,N_31875,N_30206);
nand U32371 (N_32371,N_30727,N_30186);
or U32372 (N_32372,N_30236,N_31928);
xnor U32373 (N_32373,N_30943,N_30462);
nand U32374 (N_32374,N_30401,N_30594);
xnor U32375 (N_32375,N_30286,N_31282);
xnor U32376 (N_32376,N_30417,N_30060);
xor U32377 (N_32377,N_31744,N_30289);
nand U32378 (N_32378,N_31292,N_30999);
nand U32379 (N_32379,N_30539,N_30483);
nor U32380 (N_32380,N_30566,N_31808);
nor U32381 (N_32381,N_30165,N_31559);
or U32382 (N_32382,N_30369,N_31837);
and U32383 (N_32383,N_31026,N_30359);
nand U32384 (N_32384,N_31165,N_30310);
nand U32385 (N_32385,N_30433,N_30207);
and U32386 (N_32386,N_30305,N_31399);
and U32387 (N_32387,N_31480,N_30634);
xnor U32388 (N_32388,N_30683,N_30533);
xnor U32389 (N_32389,N_30092,N_31930);
nor U32390 (N_32390,N_30589,N_31799);
nand U32391 (N_32391,N_30715,N_31598);
nand U32392 (N_32392,N_31523,N_31565);
nand U32393 (N_32393,N_30438,N_31215);
xnor U32394 (N_32394,N_30413,N_31801);
or U32395 (N_32395,N_31308,N_31816);
and U32396 (N_32396,N_31199,N_31870);
xor U32397 (N_32397,N_31675,N_30117);
nand U32398 (N_32398,N_30484,N_30633);
nand U32399 (N_32399,N_31887,N_31279);
nor U32400 (N_32400,N_30812,N_31589);
or U32401 (N_32401,N_30163,N_31492);
nor U32402 (N_32402,N_30280,N_30292);
and U32403 (N_32403,N_30978,N_30047);
xor U32404 (N_32404,N_31395,N_31307);
and U32405 (N_32405,N_30428,N_30231);
and U32406 (N_32406,N_31601,N_31544);
nor U32407 (N_32407,N_30065,N_30434);
nand U32408 (N_32408,N_31528,N_31429);
and U32409 (N_32409,N_31443,N_31561);
xor U32410 (N_32410,N_31672,N_30062);
nand U32411 (N_32411,N_31352,N_31985);
nor U32412 (N_32412,N_31889,N_31653);
and U32413 (N_32413,N_31137,N_31019);
xnor U32414 (N_32414,N_31784,N_31152);
xnor U32415 (N_32415,N_30688,N_31377);
xor U32416 (N_32416,N_30520,N_30391);
nand U32417 (N_32417,N_30868,N_31100);
nand U32418 (N_32418,N_31697,N_30106);
xor U32419 (N_32419,N_31893,N_30922);
nand U32420 (N_32420,N_31237,N_31249);
xnor U32421 (N_32421,N_31193,N_31965);
and U32422 (N_32422,N_30987,N_30759);
nor U32423 (N_32423,N_30815,N_31242);
or U32424 (N_32424,N_31704,N_30933);
and U32425 (N_32425,N_30449,N_30899);
nor U32426 (N_32426,N_30518,N_31413);
nand U32427 (N_32427,N_30035,N_30102);
and U32428 (N_32428,N_31271,N_30362);
nand U32429 (N_32429,N_30793,N_31621);
xor U32430 (N_32430,N_31255,N_30486);
xor U32431 (N_32431,N_31495,N_31105);
and U32432 (N_32432,N_31474,N_31025);
or U32433 (N_32433,N_31185,N_31743);
nor U32434 (N_32434,N_31046,N_30864);
or U32435 (N_32435,N_30784,N_30845);
or U32436 (N_32436,N_30979,N_30447);
or U32437 (N_32437,N_30962,N_30602);
or U32438 (N_32438,N_31306,N_31516);
nor U32439 (N_32439,N_30199,N_30258);
nand U32440 (N_32440,N_31123,N_30063);
and U32441 (N_32441,N_31096,N_30637);
nand U32442 (N_32442,N_30181,N_30209);
nand U32443 (N_32443,N_31171,N_30737);
nor U32444 (N_32444,N_30300,N_31998);
and U32445 (N_32445,N_31427,N_30657);
nor U32446 (N_32446,N_30083,N_31470);
nand U32447 (N_32447,N_31241,N_30103);
nand U32448 (N_32448,N_31339,N_30024);
xor U32449 (N_32449,N_30552,N_31624);
nand U32450 (N_32450,N_30842,N_31868);
nand U32451 (N_32451,N_31484,N_30755);
nor U32452 (N_32452,N_30513,N_31593);
nor U32453 (N_32453,N_30580,N_30080);
and U32454 (N_32454,N_30482,N_30861);
xor U32455 (N_32455,N_30215,N_30149);
nand U32456 (N_32456,N_30044,N_30578);
nor U32457 (N_32457,N_30887,N_31779);
or U32458 (N_32458,N_31604,N_30663);
nand U32459 (N_32459,N_30874,N_31146);
nand U32460 (N_32460,N_30195,N_30509);
xnor U32461 (N_32461,N_30468,N_31778);
nand U32462 (N_32462,N_30673,N_31995);
or U32463 (N_32463,N_31800,N_30913);
nand U32464 (N_32464,N_30796,N_31834);
nor U32465 (N_32465,N_31375,N_30332);
and U32466 (N_32466,N_31647,N_31258);
nor U32467 (N_32467,N_30905,N_31590);
or U32468 (N_32468,N_31678,N_30963);
and U32469 (N_32469,N_31392,N_30872);
xnor U32470 (N_32470,N_30607,N_31964);
nor U32471 (N_32471,N_30995,N_30091);
nor U32472 (N_32472,N_30984,N_30527);
and U32473 (N_32473,N_31449,N_30230);
xnor U32474 (N_32474,N_30584,N_31393);
or U32475 (N_32475,N_31977,N_31796);
nor U32476 (N_32476,N_31149,N_30393);
and U32477 (N_32477,N_30407,N_30326);
nand U32478 (N_32478,N_30495,N_31805);
xnor U32479 (N_32479,N_31469,N_30504);
xnor U32480 (N_32480,N_30451,N_31780);
xor U32481 (N_32481,N_31139,N_31056);
or U32482 (N_32482,N_31728,N_30295);
or U32483 (N_32483,N_30647,N_31912);
or U32484 (N_32484,N_30479,N_30086);
nand U32485 (N_32485,N_31923,N_30121);
nor U32486 (N_32486,N_31343,N_30379);
xnor U32487 (N_32487,N_30319,N_30768);
xor U32488 (N_32488,N_30877,N_30779);
and U32489 (N_32489,N_30775,N_31605);
nand U32490 (N_32490,N_31595,N_31162);
and U32491 (N_32491,N_30643,N_31188);
or U32492 (N_32492,N_30134,N_31214);
nand U32493 (N_32493,N_31656,N_31537);
and U32494 (N_32494,N_30274,N_31444);
or U32495 (N_32495,N_31633,N_31545);
or U32496 (N_32496,N_31435,N_31344);
nand U32497 (N_32497,N_30712,N_30269);
xor U32498 (N_32498,N_30128,N_30075);
nand U32499 (N_32499,N_30787,N_31878);
or U32500 (N_32500,N_31386,N_31304);
nor U32501 (N_32501,N_31717,N_30257);
nor U32502 (N_32502,N_31649,N_30126);
and U32503 (N_32503,N_31247,N_31351);
nor U32504 (N_32504,N_30998,N_31501);
or U32505 (N_32505,N_31180,N_30603);
or U32506 (N_32506,N_31937,N_31261);
xnor U32507 (N_32507,N_30961,N_30971);
nand U32508 (N_32508,N_30467,N_30610);
nor U32509 (N_32509,N_31156,N_31416);
or U32510 (N_32510,N_31959,N_31076);
and U32511 (N_32511,N_31894,N_31319);
nor U32512 (N_32512,N_31852,N_30967);
and U32513 (N_32513,N_31119,N_31030);
and U32514 (N_32514,N_30970,N_30808);
and U32515 (N_32515,N_31358,N_31551);
nand U32516 (N_32516,N_30316,N_31891);
nor U32517 (N_32517,N_30200,N_31936);
or U32518 (N_32518,N_31752,N_30143);
or U32519 (N_32519,N_30829,N_31775);
or U32520 (N_32520,N_31575,N_31160);
nor U32521 (N_32521,N_31173,N_31293);
and U32522 (N_32522,N_30392,N_31827);
or U32523 (N_32523,N_30366,N_31473);
xnor U32524 (N_32524,N_30813,N_30363);
nor U32525 (N_32525,N_30728,N_30735);
xor U32526 (N_32526,N_31390,N_30791);
or U32527 (N_32527,N_31806,N_31265);
or U32528 (N_32528,N_31191,N_31934);
nand U32529 (N_32529,N_31346,N_30002);
nor U32530 (N_32530,N_30512,N_30721);
and U32531 (N_32531,N_30256,N_30659);
nand U32532 (N_32532,N_31969,N_30849);
or U32533 (N_32533,N_30635,N_31445);
nor U32534 (N_32534,N_30240,N_30233);
nor U32535 (N_32535,N_31669,N_30918);
nand U32536 (N_32536,N_31381,N_31910);
nand U32537 (N_32537,N_30814,N_30522);
and U32538 (N_32538,N_31768,N_31077);
and U32539 (N_32539,N_31051,N_30723);
xnor U32540 (N_32540,N_31699,N_30007);
nand U32541 (N_32541,N_30959,N_30797);
and U32542 (N_32542,N_31285,N_30972);
nor U32543 (N_32543,N_30382,N_30095);
xor U32544 (N_32544,N_31378,N_31955);
xnor U32545 (N_32545,N_31512,N_30159);
xnor U32546 (N_32546,N_31236,N_30595);
xnor U32547 (N_32547,N_30026,N_30805);
nor U32548 (N_32548,N_30638,N_31585);
xor U32549 (N_32549,N_30243,N_30323);
and U32550 (N_32550,N_31200,N_30471);
nor U32551 (N_32551,N_31944,N_30361);
nor U32552 (N_32552,N_31264,N_31491);
or U32553 (N_32553,N_30137,N_31158);
nand U32554 (N_32554,N_31880,N_30945);
or U32555 (N_32555,N_31881,N_30770);
nand U32556 (N_32556,N_30936,N_30639);
nor U32557 (N_32557,N_31301,N_31513);
and U32558 (N_32558,N_30824,N_30081);
xor U32559 (N_32559,N_30232,N_30210);
xnor U32560 (N_32560,N_31219,N_30704);
and U32561 (N_32561,N_31552,N_30826);
or U32562 (N_32562,N_30660,N_30356);
or U32563 (N_32563,N_31700,N_30958);
and U32564 (N_32564,N_30315,N_30698);
xor U32565 (N_32565,N_31517,N_30694);
and U32566 (N_32566,N_30214,N_30329);
xor U32567 (N_32567,N_31576,N_31089);
and U32568 (N_32568,N_30646,N_30228);
and U32569 (N_32569,N_31638,N_30830);
nand U32570 (N_32570,N_31456,N_31251);
nand U32571 (N_32571,N_31091,N_30440);
or U32572 (N_32572,N_31129,N_31176);
nor U32573 (N_32573,N_30540,N_31432);
or U32574 (N_32574,N_31690,N_30443);
and U32575 (N_32575,N_30096,N_31984);
nor U32576 (N_32576,N_31736,N_30608);
xnor U32577 (N_32577,N_31273,N_31208);
and U32578 (N_32578,N_30234,N_31982);
nor U32579 (N_32579,N_30478,N_30101);
nand U32580 (N_32580,N_30148,N_30892);
or U32581 (N_32581,N_31276,N_30524);
nor U32582 (N_32582,N_31220,N_30390);
nor U32583 (N_32583,N_31795,N_30185);
or U32584 (N_32584,N_30372,N_30558);
nor U32585 (N_32585,N_31674,N_31231);
nand U32586 (N_32586,N_30312,N_31739);
nor U32587 (N_32587,N_30406,N_30574);
or U32588 (N_32588,N_30724,N_30615);
and U32589 (N_32589,N_31751,N_30263);
nor U32590 (N_32590,N_30132,N_30692);
nand U32591 (N_32591,N_30820,N_30729);
and U32592 (N_32592,N_31838,N_30767);
or U32593 (N_32593,N_31636,N_30535);
xor U32594 (N_32594,N_30816,N_30537);
or U32595 (N_32595,N_31321,N_31538);
and U32596 (N_32596,N_31439,N_30620);
or U32597 (N_32597,N_31882,N_31766);
or U32598 (N_32598,N_31786,N_30923);
and U32599 (N_32599,N_30354,N_30189);
xor U32600 (N_32600,N_30622,N_31110);
nand U32601 (N_32601,N_30525,N_31345);
xnor U32602 (N_32602,N_31202,N_31262);
xnor U32603 (N_32603,N_30367,N_31283);
nand U32604 (N_32604,N_30543,N_30203);
and U32605 (N_32605,N_31347,N_30691);
or U32606 (N_32606,N_31817,N_30585);
nand U32607 (N_32607,N_30107,N_30016);
nor U32608 (N_32608,N_31587,N_30246);
xnor U32609 (N_32609,N_31924,N_30009);
nand U32610 (N_32610,N_31353,N_31922);
xnor U32611 (N_32611,N_30054,N_30279);
and U32612 (N_32612,N_31205,N_30873);
nor U32613 (N_32613,N_31412,N_31691);
nand U32614 (N_32614,N_30928,N_31632);
nor U32615 (N_32615,N_30799,N_30076);
or U32616 (N_32616,N_30445,N_30840);
nand U32617 (N_32617,N_31256,N_30895);
xnor U32618 (N_32618,N_31369,N_31107);
nand U32619 (N_32619,N_31584,N_31946);
nand U32620 (N_32620,N_30155,N_31078);
nand U32621 (N_32621,N_30711,N_30211);
or U32622 (N_32622,N_30333,N_31420);
xnor U32623 (N_32623,N_31382,N_31581);
nor U32624 (N_32624,N_31726,N_31379);
or U32625 (N_32625,N_31477,N_31023);
and U32626 (N_32626,N_31958,N_31904);
nand U32627 (N_32627,N_30798,N_30238);
nand U32628 (N_32628,N_30160,N_31425);
or U32629 (N_32629,N_31475,N_31673);
xnor U32630 (N_32630,N_31919,N_31962);
nor U32631 (N_32631,N_30932,N_30930);
nand U32632 (N_32632,N_30229,N_30108);
or U32633 (N_32633,N_31828,N_31418);
and U32634 (N_32634,N_31844,N_31637);
and U32635 (N_32635,N_30046,N_30517);
or U32636 (N_32636,N_30857,N_30718);
xnor U32637 (N_32637,N_30304,N_31809);
or U32638 (N_32638,N_30105,N_31599);
xor U32639 (N_32639,N_30375,N_30041);
and U32640 (N_32640,N_31294,N_31095);
nand U32641 (N_32641,N_30350,N_30846);
nand U32642 (N_32642,N_30178,N_30153);
nand U32643 (N_32643,N_30738,N_30713);
or U32644 (N_32644,N_30296,N_30077);
nand U32645 (N_32645,N_30177,N_30848);
or U32646 (N_32646,N_30760,N_31189);
and U32647 (N_32647,N_31940,N_30579);
or U32648 (N_32648,N_31987,N_30508);
or U32649 (N_32649,N_31884,N_30345);
nor U32650 (N_32650,N_30118,N_31741);
nor U32651 (N_32651,N_30174,N_31859);
or U32652 (N_32652,N_30297,N_31724);
nor U32653 (N_32653,N_30031,N_31941);
nor U32654 (N_32654,N_30514,N_30699);
and U32655 (N_32655,N_31287,N_30769);
or U32656 (N_32656,N_31508,N_31612);
and U32657 (N_32657,N_31831,N_31034);
or U32658 (N_32658,N_30675,N_30291);
or U32659 (N_32659,N_31914,N_30880);
nand U32660 (N_32660,N_31458,N_30687);
nor U32661 (N_32661,N_31083,N_30853);
and U32662 (N_32662,N_31454,N_30731);
nor U32663 (N_32663,N_31125,N_31298);
or U32664 (N_32664,N_31097,N_30757);
xor U32665 (N_32665,N_30931,N_30626);
nand U32666 (N_32666,N_30115,N_31853);
xnor U32667 (N_32667,N_30804,N_30935);
xnor U32668 (N_32668,N_30810,N_30701);
nor U32669 (N_32669,N_31902,N_30003);
nand U32670 (N_32670,N_31974,N_30498);
nor U32671 (N_32671,N_30384,N_30098);
nand U32672 (N_32672,N_31464,N_31566);
or U32673 (N_32673,N_30420,N_31225);
nor U32674 (N_32674,N_30006,N_30122);
nor U32675 (N_32675,N_31437,N_30818);
and U32676 (N_32676,N_31092,N_31069);
nand U32677 (N_32677,N_30617,N_30038);
or U32678 (N_32678,N_30164,N_31812);
or U32679 (N_32679,N_31461,N_31216);
nand U32680 (N_32680,N_31111,N_30015);
xnor U32681 (N_32681,N_31725,N_30225);
or U32682 (N_32682,N_30441,N_31681);
and U32683 (N_32683,N_31953,N_30802);
and U32684 (N_32684,N_30632,N_30696);
or U32685 (N_32685,N_31658,N_31548);
and U32686 (N_32686,N_30623,N_31607);
xnor U32687 (N_32687,N_30224,N_31687);
nand U32688 (N_32688,N_30004,N_31613);
and U32689 (N_32689,N_30461,N_30593);
nand U32690 (N_32690,N_31750,N_31820);
xor U32691 (N_32691,N_30097,N_30183);
nor U32692 (N_32692,N_31804,N_31932);
xnor U32693 (N_32693,N_31802,N_31391);
nand U32694 (N_32694,N_30120,N_31608);
xnor U32695 (N_32695,N_30771,N_30043);
nand U32696 (N_32696,N_31310,N_30172);
nand U32697 (N_32697,N_31085,N_31325);
or U32698 (N_32698,N_31115,N_31908);
nor U32699 (N_32699,N_31288,N_30627);
or U32700 (N_32700,N_31972,N_30908);
or U32701 (N_32701,N_31588,N_31869);
nand U32702 (N_32702,N_31127,N_31305);
xnor U32703 (N_32703,N_30180,N_31945);
and U32704 (N_32704,N_30661,N_31715);
xnor U32705 (N_32705,N_31175,N_30017);
and U32706 (N_32706,N_31597,N_31570);
nand U32707 (N_32707,N_30850,N_30142);
xor U32708 (N_32708,N_30100,N_30381);
xnor U32709 (N_32709,N_30340,N_30001);
and U32710 (N_32710,N_31372,N_30299);
nor U32711 (N_32711,N_30014,N_30989);
nor U32712 (N_32712,N_31871,N_31885);
nand U32713 (N_32713,N_30569,N_31679);
xor U32714 (N_32714,N_30505,N_30690);
or U32715 (N_32715,N_31415,N_30277);
and U32716 (N_32716,N_30841,N_31278);
nor U32717 (N_32717,N_31407,N_31644);
and U32718 (N_32718,N_30012,N_30587);
xor U32719 (N_32719,N_31212,N_31350);
xor U32720 (N_32720,N_30448,N_30809);
nor U32721 (N_32721,N_30064,N_30920);
nor U32722 (N_32722,N_30196,N_31920);
xor U32723 (N_32723,N_31067,N_31303);
xor U32724 (N_32724,N_30739,N_31927);
xor U32725 (N_32725,N_30990,N_31032);
and U32726 (N_32726,N_31684,N_31993);
nor U32727 (N_32727,N_31948,N_31424);
xor U32728 (N_32728,N_31685,N_31334);
nand U32729 (N_32729,N_31793,N_31921);
and U32730 (N_32730,N_31522,N_31411);
or U32731 (N_32731,N_30193,N_31515);
and U32732 (N_32732,N_30823,N_30327);
nor U32733 (N_32733,N_30902,N_31014);
xor U32734 (N_32734,N_31535,N_30754);
and U32735 (N_32735,N_30442,N_30089);
or U32736 (N_32736,N_31135,N_31701);
xor U32737 (N_32737,N_31385,N_31727);
and U32738 (N_32738,N_31519,N_30244);
nand U32739 (N_32739,N_30194,N_31052);
xnor U32740 (N_32740,N_30336,N_30217);
nand U32741 (N_32741,N_30349,N_31776);
xnor U32742 (N_32742,N_30878,N_31895);
nor U32743 (N_32743,N_31702,N_31737);
or U32744 (N_32744,N_30669,N_30283);
xnor U32745 (N_32745,N_31057,N_30028);
xor U32746 (N_32746,N_31109,N_31357);
nor U32747 (N_32747,N_30766,N_31521);
and U32748 (N_32748,N_31218,N_31274);
nor U32749 (N_32749,N_30109,N_30353);
and U32750 (N_32750,N_30720,N_30268);
xor U32751 (N_32751,N_31120,N_30648);
and U32752 (N_32752,N_30710,N_31824);
nor U32753 (N_32753,N_30124,N_30226);
nor U32754 (N_32754,N_31419,N_30358);
nand U32755 (N_32755,N_30307,N_31618);
nand U32756 (N_32756,N_31720,N_30705);
nand U32757 (N_32757,N_30110,N_31460);
nand U32758 (N_32758,N_31154,N_31874);
nor U32759 (N_32759,N_31290,N_30262);
nand U32760 (N_32760,N_30364,N_30652);
nor U32761 (N_32761,N_30290,N_31532);
xor U32762 (N_32762,N_30565,N_31126);
or U32763 (N_32763,N_30903,N_31075);
nor U32764 (N_32764,N_31557,N_31996);
xor U32765 (N_32765,N_30819,N_30618);
xor U32766 (N_32766,N_31872,N_30067);
or U32767 (N_32767,N_31143,N_30950);
nor U32768 (N_32768,N_31045,N_30190);
or U32769 (N_32769,N_31108,N_31483);
and U32770 (N_32770,N_31698,N_30387);
xnor U32771 (N_32771,N_30073,N_31916);
and U32772 (N_32772,N_30168,N_30473);
or U32773 (N_32773,N_30725,N_30598);
nand U32774 (N_32774,N_30924,N_30807);
or U32775 (N_32775,N_31040,N_31705);
nor U32776 (N_32776,N_30344,N_31883);
or U32777 (N_32777,N_30538,N_30188);
nand U32778 (N_32778,N_30475,N_30116);
nor U32779 (N_32779,N_31312,N_30997);
or U32780 (N_32780,N_31625,N_30056);
and U32781 (N_32781,N_30686,N_30418);
and U32782 (N_32782,N_31068,N_31348);
or U32783 (N_32783,N_31639,N_31925);
nand U32784 (N_32784,N_30446,N_30303);
or U32785 (N_32785,N_31663,N_31359);
xor U32786 (N_32786,N_31854,N_30611);
nor U32787 (N_32787,N_31642,N_30996);
nor U32788 (N_32788,N_31533,N_31622);
or U32789 (N_32789,N_30111,N_31781);
nor U32790 (N_32790,N_30497,N_30499);
nor U32791 (N_32791,N_31848,N_30251);
and U32792 (N_32792,N_30450,N_31489);
nand U32793 (N_32793,N_31531,N_31009);
nand U32794 (N_32794,N_31926,N_30125);
and U32795 (N_32795,N_30218,N_30937);
nor U32796 (N_32796,N_31646,N_30680);
or U32797 (N_32797,N_30173,N_30061);
nor U32798 (N_32798,N_30385,N_31462);
nor U32799 (N_32799,N_30457,N_31905);
xor U32800 (N_32800,N_31327,N_31022);
and U32801 (N_32801,N_31409,N_31017);
xnor U32802 (N_32802,N_31163,N_31388);
or U32803 (N_32803,N_31782,N_30170);
nand U32804 (N_32804,N_31763,N_31721);
nor U32805 (N_32805,N_30719,N_30888);
nor U32806 (N_32806,N_31457,N_30301);
xor U32807 (N_32807,N_30247,N_30883);
and U32808 (N_32808,N_30293,N_30742);
or U32809 (N_32809,N_31335,N_30549);
and U32810 (N_32810,N_30284,N_30949);
nand U32811 (N_32811,N_30444,N_31151);
or U32812 (N_32812,N_31194,N_31248);
nand U32813 (N_32813,N_30744,N_31832);
nand U32814 (N_32814,N_30761,N_31013);
and U32815 (N_32815,N_31567,N_30314);
and U32816 (N_32816,N_31284,N_30625);
nor U32817 (N_32817,N_31866,N_31281);
nor U32818 (N_32818,N_31080,N_30973);
nor U32819 (N_32819,N_31586,N_31757);
or U32820 (N_32820,N_30695,N_30751);
xor U32821 (N_32821,N_31626,N_30557);
or U32822 (N_32822,N_31686,N_31764);
nor U32823 (N_32823,N_30777,N_30689);
or U32824 (N_32824,N_31387,N_31000);
and U32825 (N_32825,N_31326,N_31210);
nor U32826 (N_32826,N_31141,N_30136);
xnor U32827 (N_32827,N_30628,N_30629);
nor U32828 (N_32828,N_31813,N_30469);
or U32829 (N_32829,N_30175,N_31493);
and U32830 (N_32830,N_30896,N_30351);
xnor U32831 (N_32831,N_30581,N_30281);
nor U32832 (N_32832,N_31084,N_31455);
nand U32833 (N_32833,N_31527,N_30960);
nand U32834 (N_32834,N_31227,N_31856);
or U32835 (N_32835,N_30773,N_31667);
and U32836 (N_32836,N_31331,N_30239);
or U32837 (N_32837,N_30237,N_30828);
xor U32838 (N_32838,N_30197,N_30590);
or U32839 (N_32839,N_30834,N_31554);
nand U32840 (N_32840,N_31755,N_31839);
and U32841 (N_32841,N_30653,N_30624);
xnor U32842 (N_32842,N_31909,N_30838);
xnor U32843 (N_32843,N_30147,N_31179);
nand U32844 (N_32844,N_31747,N_31677);
nand U32845 (N_32845,N_31408,N_30474);
nand U32846 (N_32846,N_30662,N_31992);
nor U32847 (N_32847,N_30347,N_31547);
and U32848 (N_32848,N_31730,N_31297);
nand U32849 (N_32849,N_30946,N_31509);
nand U32850 (N_32850,N_31367,N_30609);
nor U32851 (N_32851,N_30641,N_30907);
nor U32852 (N_32852,N_30250,N_31994);
or U32853 (N_32853,N_31617,N_30383);
xnor U32854 (N_32854,N_31239,N_30021);
and U32855 (N_32855,N_30396,N_31061);
nor U32856 (N_32856,N_31579,N_30803);
xnor U32857 (N_32857,N_31933,N_31072);
nand U32858 (N_32858,N_31555,N_30571);
nand U32859 (N_32859,N_30287,N_30644);
or U32860 (N_32860,N_31988,N_31708);
and U32861 (N_32861,N_31789,N_31468);
nor U32862 (N_32862,N_30914,N_31973);
and U32863 (N_32863,N_30492,N_31245);
nor U32864 (N_32864,N_30790,N_30013);
or U32865 (N_32865,N_31803,N_31338);
or U32866 (N_32866,N_31471,N_30780);
and U32867 (N_32867,N_30545,N_30176);
xnor U32868 (N_32868,N_31733,N_30521);
nor U32869 (N_32869,N_31007,N_30800);
and U32870 (N_32870,N_30090,N_30909);
nor U32871 (N_32871,N_31155,N_30734);
and U32872 (N_32872,N_30572,N_31849);
and U32873 (N_32873,N_31015,N_30601);
nand U32874 (N_32874,N_31224,N_30477);
nand U32875 (N_32875,N_31847,N_30855);
nor U32876 (N_32876,N_31765,N_31465);
xnor U32877 (N_32877,N_30059,N_31746);
nand U32878 (N_32878,N_31990,N_31147);
and U32879 (N_32879,N_31505,N_30553);
xor U32880 (N_32880,N_30682,N_31903);
and U32881 (N_32881,N_31665,N_31929);
xor U32882 (N_32882,N_30198,N_31703);
and U32883 (N_32883,N_30045,N_31272);
nand U32884 (N_32884,N_30859,N_31337);
nand U32885 (N_32885,N_31071,N_31654);
nand U32886 (N_32886,N_30019,N_30542);
nor U32887 (N_32887,N_30399,N_30320);
nand U32888 (N_32888,N_31892,N_31615);
nand U32889 (N_32889,N_30298,N_31833);
nor U32890 (N_32890,N_30886,N_31406);
nand U32891 (N_32891,N_30099,N_31735);
nor U32892 (N_32892,N_31863,N_31268);
or U32893 (N_32893,N_31580,N_30412);
and U32894 (N_32894,N_31088,N_30655);
xor U32895 (N_32895,N_30975,N_31603);
or U32896 (N_32896,N_30502,N_30722);
nand U32897 (N_32897,N_30865,N_31099);
nor U32898 (N_32898,N_31645,N_31811);
nand U32899 (N_32899,N_30071,N_31403);
nor U32900 (N_32900,N_30032,N_31668);
or U32901 (N_32901,N_30208,N_30306);
and U32902 (N_32902,N_31027,N_30740);
and U32903 (N_32903,N_31062,N_31228);
or U32904 (N_32904,N_31710,N_30437);
xnor U32905 (N_32905,N_30048,N_31935);
and U32906 (N_32906,N_31476,N_30948);
xor U32907 (N_32907,N_31401,N_31037);
nand U32908 (N_32908,N_30968,N_30630);
and U32909 (N_32909,N_31543,N_30051);
nand U32910 (N_32910,N_31867,N_31857);
or U32911 (N_32911,N_30259,N_30869);
xor U32912 (N_32912,N_30916,N_31635);
nand U32913 (N_32913,N_30876,N_31333);
nand U32914 (N_32914,N_31851,N_30145);
nand U32915 (N_32915,N_30827,N_30956);
xnor U32916 (N_32916,N_30893,N_30150);
or U32917 (N_32917,N_31873,N_31640);
xnor U32918 (N_32918,N_30426,N_31680);
xor U32919 (N_32919,N_30161,N_30378);
nand U32920 (N_32920,N_31434,N_31600);
and U32921 (N_32921,N_30264,N_31949);
or U32922 (N_32922,N_31787,N_31906);
nor U32923 (N_32923,N_30570,N_30817);
and U32924 (N_32924,N_30040,N_31865);
nor U32925 (N_32925,N_31738,N_31004);
or U32926 (N_32926,N_31362,N_31440);
nand U32927 (N_32927,N_31659,N_31981);
xor U32928 (N_32928,N_31676,N_30672);
and U32929 (N_32929,N_31983,N_30050);
nor U32930 (N_32930,N_30042,N_30743);
xnor U32931 (N_32931,N_30220,N_30983);
and U32932 (N_32932,N_30776,N_30693);
nand U32933 (N_32933,N_30162,N_30227);
nor U32934 (N_32934,N_31159,N_30348);
nand U32935 (N_32935,N_30833,N_31082);
xor U32936 (N_32936,N_30588,N_30940);
nand U32937 (N_32937,N_31053,N_30085);
nor U32938 (N_32938,N_31520,N_31114);
nor U32939 (N_32939,N_31980,N_30318);
xor U32940 (N_32940,N_30929,N_30523);
nor U32941 (N_32941,N_31103,N_30459);
xnor U32942 (N_32942,N_31568,N_30832);
nand U32943 (N_32943,N_30386,N_31829);
and U32944 (N_32944,N_31318,N_30764);
xnor U32945 (N_32945,N_31463,N_31142);
nor U32946 (N_32946,N_30650,N_30709);
or U32947 (N_32947,N_31564,N_31846);
xor U32948 (N_32948,N_30685,N_30403);
nor U32949 (N_32949,N_30427,N_31858);
and U32950 (N_32950,N_31911,N_30058);
nor U32951 (N_32951,N_30365,N_31328);
and U32952 (N_32952,N_30867,N_31195);
xor U32953 (N_32953,N_30889,N_30011);
xor U32954 (N_32954,N_30700,N_30463);
nor U32955 (N_32955,N_30927,N_31038);
and U32956 (N_32956,N_31039,N_30904);
nor U32957 (N_32957,N_30066,N_30870);
nor U32958 (N_32958,N_30154,N_31329);
or U32959 (N_32959,N_30750,N_31619);
and U32960 (N_32960,N_31230,N_30267);
and U32961 (N_32961,N_31536,N_31008);
xor U32962 (N_32962,N_30453,N_30965);
or U32963 (N_32963,N_30235,N_30906);
nand U32964 (N_32964,N_31090,N_30981);
nand U32965 (N_32965,N_31299,N_31609);
or U32966 (N_32966,N_31309,N_30490);
or U32967 (N_32967,N_30576,N_30036);
and U32968 (N_32968,N_30131,N_30337);
and U32969 (N_32969,N_31967,N_30328);
xnor U32970 (N_32970,N_31011,N_30425);
or U32971 (N_32971,N_30702,N_30897);
xor U32972 (N_32972,N_31818,N_31021);
xor U32973 (N_32973,N_31560,N_31966);
or U32974 (N_32974,N_30037,N_31898);
or U32975 (N_32975,N_30547,N_30756);
or U32976 (N_32976,N_31438,N_31041);
nand U32977 (N_32977,N_30123,N_30266);
nand U32978 (N_32978,N_31578,N_30531);
nor U32979 (N_32979,N_30000,N_31201);
nand U32980 (N_32980,N_30988,N_30714);
and U32981 (N_32981,N_31238,N_30875);
xor U32982 (N_32982,N_31488,N_31997);
xor U32983 (N_32983,N_30606,N_31886);
xnor U32984 (N_32984,N_30674,N_31712);
nand U32985 (N_32985,N_31620,N_31901);
nor U32986 (N_32986,N_31150,N_30377);
and U32987 (N_32987,N_30747,N_31696);
and U32988 (N_32988,N_30270,N_31499);
nor U32989 (N_32989,N_31862,N_31314);
and U32990 (N_32990,N_30898,N_31055);
nor U32991 (N_32991,N_30582,N_31431);
nor U32992 (N_32992,N_31466,N_31876);
or U32993 (N_32993,N_31104,N_30559);
or U32994 (N_32994,N_31124,N_31302);
and U32995 (N_32995,N_31330,N_30500);
nor U32996 (N_32996,N_30917,N_31770);
nand U32997 (N_32997,N_31286,N_31020);
or U32998 (N_32998,N_30591,N_31453);
and U32999 (N_32999,N_31542,N_31991);
and U33000 (N_33000,N_30521,N_30984);
nand U33001 (N_33001,N_30479,N_31712);
xnor U33002 (N_33002,N_30019,N_30165);
nand U33003 (N_33003,N_31787,N_31410);
nor U33004 (N_33004,N_31127,N_30696);
and U33005 (N_33005,N_30826,N_30697);
xnor U33006 (N_33006,N_30865,N_30205);
nor U33007 (N_33007,N_30418,N_31777);
xor U33008 (N_33008,N_31069,N_31766);
and U33009 (N_33009,N_30539,N_30172);
nor U33010 (N_33010,N_30408,N_31108);
nor U33011 (N_33011,N_31908,N_31403);
and U33012 (N_33012,N_30223,N_31010);
nand U33013 (N_33013,N_31158,N_31664);
nor U33014 (N_33014,N_31045,N_30798);
and U33015 (N_33015,N_30460,N_30247);
or U33016 (N_33016,N_30620,N_31901);
nor U33017 (N_33017,N_30821,N_30927);
nor U33018 (N_33018,N_31175,N_30422);
and U33019 (N_33019,N_31943,N_30106);
or U33020 (N_33020,N_31717,N_31857);
or U33021 (N_33021,N_30707,N_30498);
or U33022 (N_33022,N_31349,N_30444);
nand U33023 (N_33023,N_30321,N_31687);
xor U33024 (N_33024,N_30413,N_31083);
nand U33025 (N_33025,N_31884,N_30889);
and U33026 (N_33026,N_30553,N_31971);
and U33027 (N_33027,N_31851,N_31339);
nand U33028 (N_33028,N_30223,N_31242);
nand U33029 (N_33029,N_31470,N_30364);
nor U33030 (N_33030,N_31859,N_31762);
or U33031 (N_33031,N_31009,N_31219);
nand U33032 (N_33032,N_30972,N_30748);
nand U33033 (N_33033,N_31122,N_30107);
xnor U33034 (N_33034,N_31178,N_30960);
and U33035 (N_33035,N_30031,N_31989);
nor U33036 (N_33036,N_30867,N_31861);
nor U33037 (N_33037,N_30716,N_31149);
nor U33038 (N_33038,N_30546,N_31288);
and U33039 (N_33039,N_31977,N_30755);
or U33040 (N_33040,N_30253,N_30762);
and U33041 (N_33041,N_30686,N_31490);
and U33042 (N_33042,N_31132,N_30088);
xnor U33043 (N_33043,N_31323,N_31889);
xnor U33044 (N_33044,N_30511,N_30535);
and U33045 (N_33045,N_30398,N_30833);
nand U33046 (N_33046,N_31553,N_30830);
nor U33047 (N_33047,N_30427,N_30626);
nor U33048 (N_33048,N_30093,N_30943);
nor U33049 (N_33049,N_30549,N_30889);
nor U33050 (N_33050,N_31945,N_31856);
xor U33051 (N_33051,N_31065,N_31763);
or U33052 (N_33052,N_30304,N_30648);
nor U33053 (N_33053,N_31188,N_30135);
nor U33054 (N_33054,N_31393,N_31108);
xnor U33055 (N_33055,N_30553,N_31452);
xnor U33056 (N_33056,N_31753,N_30785);
nor U33057 (N_33057,N_30102,N_31517);
nor U33058 (N_33058,N_31470,N_30487);
nand U33059 (N_33059,N_30804,N_31354);
xor U33060 (N_33060,N_31304,N_30422);
and U33061 (N_33061,N_30518,N_31313);
or U33062 (N_33062,N_30125,N_31399);
nand U33063 (N_33063,N_30253,N_31016);
or U33064 (N_33064,N_31501,N_31854);
nor U33065 (N_33065,N_30879,N_30336);
or U33066 (N_33066,N_31021,N_31506);
nand U33067 (N_33067,N_31202,N_30641);
xnor U33068 (N_33068,N_30027,N_31863);
nand U33069 (N_33069,N_31585,N_31860);
nand U33070 (N_33070,N_31223,N_31521);
nor U33071 (N_33071,N_31352,N_31777);
xnor U33072 (N_33072,N_31846,N_30984);
or U33073 (N_33073,N_31620,N_31516);
nor U33074 (N_33074,N_30583,N_30178);
and U33075 (N_33075,N_31144,N_30259);
xnor U33076 (N_33076,N_31029,N_31437);
xor U33077 (N_33077,N_31084,N_31019);
nand U33078 (N_33078,N_31349,N_31385);
xnor U33079 (N_33079,N_30166,N_30177);
nor U33080 (N_33080,N_31772,N_30567);
and U33081 (N_33081,N_31207,N_31699);
xor U33082 (N_33082,N_30415,N_31485);
and U33083 (N_33083,N_30800,N_30388);
and U33084 (N_33084,N_30504,N_31162);
xor U33085 (N_33085,N_31159,N_31575);
xnor U33086 (N_33086,N_30851,N_31846);
and U33087 (N_33087,N_30097,N_30985);
nor U33088 (N_33088,N_30672,N_30915);
and U33089 (N_33089,N_31672,N_30668);
nor U33090 (N_33090,N_31455,N_30781);
xnor U33091 (N_33091,N_30173,N_31214);
nand U33092 (N_33092,N_30230,N_31803);
nand U33093 (N_33093,N_31262,N_31956);
xor U33094 (N_33094,N_31805,N_30701);
nand U33095 (N_33095,N_31285,N_31627);
nand U33096 (N_33096,N_30045,N_30224);
or U33097 (N_33097,N_30438,N_30558);
xnor U33098 (N_33098,N_30104,N_30134);
and U33099 (N_33099,N_31758,N_30910);
nor U33100 (N_33100,N_30957,N_30780);
and U33101 (N_33101,N_31157,N_31876);
nand U33102 (N_33102,N_30988,N_31565);
xnor U33103 (N_33103,N_31531,N_30817);
nand U33104 (N_33104,N_30312,N_31098);
nor U33105 (N_33105,N_31717,N_30470);
xor U33106 (N_33106,N_31109,N_30938);
and U33107 (N_33107,N_31042,N_30811);
nand U33108 (N_33108,N_30920,N_31647);
or U33109 (N_33109,N_30730,N_30361);
nor U33110 (N_33110,N_31868,N_31876);
and U33111 (N_33111,N_30838,N_30549);
and U33112 (N_33112,N_30549,N_30087);
and U33113 (N_33113,N_31382,N_31116);
and U33114 (N_33114,N_30053,N_30373);
nand U33115 (N_33115,N_30464,N_30267);
or U33116 (N_33116,N_30683,N_31077);
xnor U33117 (N_33117,N_31182,N_31633);
or U33118 (N_33118,N_31558,N_31578);
nand U33119 (N_33119,N_30181,N_30736);
and U33120 (N_33120,N_30156,N_30123);
nand U33121 (N_33121,N_30788,N_31357);
nor U33122 (N_33122,N_30255,N_31025);
and U33123 (N_33123,N_31469,N_30814);
nand U33124 (N_33124,N_31889,N_31308);
nor U33125 (N_33125,N_31305,N_30798);
xor U33126 (N_33126,N_30678,N_31685);
xnor U33127 (N_33127,N_30951,N_31417);
xnor U33128 (N_33128,N_30554,N_30696);
xor U33129 (N_33129,N_31561,N_30289);
nand U33130 (N_33130,N_31107,N_31890);
nor U33131 (N_33131,N_30491,N_30615);
and U33132 (N_33132,N_30928,N_30775);
nand U33133 (N_33133,N_30280,N_30124);
and U33134 (N_33134,N_31284,N_30959);
xor U33135 (N_33135,N_31344,N_30794);
nor U33136 (N_33136,N_30364,N_31353);
or U33137 (N_33137,N_30369,N_31190);
xnor U33138 (N_33138,N_30841,N_31494);
nand U33139 (N_33139,N_31667,N_30230);
or U33140 (N_33140,N_31334,N_31489);
and U33141 (N_33141,N_30911,N_30540);
nor U33142 (N_33142,N_31382,N_30721);
and U33143 (N_33143,N_30131,N_30818);
xor U33144 (N_33144,N_31436,N_31432);
nand U33145 (N_33145,N_31979,N_31863);
or U33146 (N_33146,N_31977,N_31031);
nor U33147 (N_33147,N_31958,N_31585);
or U33148 (N_33148,N_31682,N_31450);
and U33149 (N_33149,N_30169,N_31899);
xor U33150 (N_33150,N_31725,N_31474);
xor U33151 (N_33151,N_30546,N_31910);
xor U33152 (N_33152,N_30547,N_31265);
and U33153 (N_33153,N_30364,N_31201);
nand U33154 (N_33154,N_31219,N_30146);
nor U33155 (N_33155,N_30929,N_31665);
or U33156 (N_33156,N_30980,N_30278);
and U33157 (N_33157,N_30033,N_31684);
and U33158 (N_33158,N_30961,N_30357);
and U33159 (N_33159,N_30764,N_30828);
or U33160 (N_33160,N_31751,N_30260);
nand U33161 (N_33161,N_31923,N_31444);
nand U33162 (N_33162,N_31030,N_31831);
nand U33163 (N_33163,N_31111,N_31753);
or U33164 (N_33164,N_30126,N_31475);
nand U33165 (N_33165,N_31966,N_30298);
nand U33166 (N_33166,N_30050,N_30956);
nand U33167 (N_33167,N_31207,N_31742);
nand U33168 (N_33168,N_30474,N_31773);
xor U33169 (N_33169,N_31075,N_30554);
and U33170 (N_33170,N_30815,N_31906);
nor U33171 (N_33171,N_30116,N_31416);
nand U33172 (N_33172,N_31299,N_30144);
nand U33173 (N_33173,N_31602,N_30822);
or U33174 (N_33174,N_31457,N_30038);
nor U33175 (N_33175,N_31218,N_30220);
nand U33176 (N_33176,N_31782,N_31644);
nor U33177 (N_33177,N_30175,N_30802);
or U33178 (N_33178,N_31928,N_30779);
or U33179 (N_33179,N_30274,N_30439);
xor U33180 (N_33180,N_30087,N_30534);
xnor U33181 (N_33181,N_30734,N_30966);
or U33182 (N_33182,N_31482,N_30341);
nor U33183 (N_33183,N_31201,N_31789);
and U33184 (N_33184,N_31329,N_30832);
nand U33185 (N_33185,N_31785,N_30284);
or U33186 (N_33186,N_31761,N_30098);
and U33187 (N_33187,N_30584,N_31511);
nor U33188 (N_33188,N_31993,N_30604);
and U33189 (N_33189,N_30144,N_30407);
xor U33190 (N_33190,N_31135,N_31113);
and U33191 (N_33191,N_31345,N_30964);
xnor U33192 (N_33192,N_31283,N_31162);
xnor U33193 (N_33193,N_30363,N_31292);
nor U33194 (N_33194,N_30237,N_30840);
or U33195 (N_33195,N_31415,N_31093);
or U33196 (N_33196,N_31730,N_31152);
xnor U33197 (N_33197,N_30184,N_31898);
nor U33198 (N_33198,N_30568,N_30365);
and U33199 (N_33199,N_31819,N_31824);
nand U33200 (N_33200,N_31406,N_30681);
or U33201 (N_33201,N_30411,N_30794);
and U33202 (N_33202,N_31918,N_30806);
and U33203 (N_33203,N_30595,N_31383);
and U33204 (N_33204,N_30827,N_31680);
and U33205 (N_33205,N_31004,N_30176);
xnor U33206 (N_33206,N_31761,N_31275);
xor U33207 (N_33207,N_31963,N_30711);
or U33208 (N_33208,N_30040,N_31041);
or U33209 (N_33209,N_31695,N_31124);
xnor U33210 (N_33210,N_30824,N_31205);
xnor U33211 (N_33211,N_30350,N_30106);
xnor U33212 (N_33212,N_30173,N_31140);
xnor U33213 (N_33213,N_30983,N_31170);
or U33214 (N_33214,N_30682,N_30990);
and U33215 (N_33215,N_31365,N_31070);
xnor U33216 (N_33216,N_31346,N_31796);
nand U33217 (N_33217,N_30338,N_30258);
and U33218 (N_33218,N_31085,N_30700);
or U33219 (N_33219,N_31798,N_31642);
xnor U33220 (N_33220,N_31439,N_31570);
nor U33221 (N_33221,N_30021,N_31446);
and U33222 (N_33222,N_30008,N_31194);
or U33223 (N_33223,N_31640,N_30896);
xor U33224 (N_33224,N_31992,N_30197);
or U33225 (N_33225,N_31230,N_30214);
and U33226 (N_33226,N_31774,N_31176);
nor U33227 (N_33227,N_30200,N_30566);
nor U33228 (N_33228,N_31167,N_31702);
nand U33229 (N_33229,N_31000,N_31995);
nand U33230 (N_33230,N_30498,N_31700);
or U33231 (N_33231,N_31216,N_31147);
or U33232 (N_33232,N_30545,N_30790);
xor U33233 (N_33233,N_31945,N_31019);
nor U33234 (N_33234,N_31279,N_31482);
and U33235 (N_33235,N_31056,N_30427);
nand U33236 (N_33236,N_30654,N_30269);
xnor U33237 (N_33237,N_31621,N_31281);
or U33238 (N_33238,N_30711,N_30251);
xnor U33239 (N_33239,N_30397,N_30701);
nand U33240 (N_33240,N_30632,N_31662);
nor U33241 (N_33241,N_30032,N_30854);
xor U33242 (N_33242,N_31212,N_31282);
nand U33243 (N_33243,N_30980,N_31809);
or U33244 (N_33244,N_31720,N_30848);
and U33245 (N_33245,N_30074,N_31168);
nor U33246 (N_33246,N_31312,N_30767);
and U33247 (N_33247,N_30218,N_30821);
xor U33248 (N_33248,N_31201,N_31718);
nor U33249 (N_33249,N_30889,N_31625);
or U33250 (N_33250,N_30540,N_30471);
xor U33251 (N_33251,N_30373,N_30094);
xor U33252 (N_33252,N_30400,N_31449);
xnor U33253 (N_33253,N_30777,N_30019);
nand U33254 (N_33254,N_30364,N_30980);
or U33255 (N_33255,N_30850,N_31331);
xor U33256 (N_33256,N_30977,N_30639);
nand U33257 (N_33257,N_30959,N_30112);
nand U33258 (N_33258,N_31661,N_30362);
or U33259 (N_33259,N_31519,N_31264);
and U33260 (N_33260,N_31684,N_30599);
and U33261 (N_33261,N_30641,N_31512);
xor U33262 (N_33262,N_30095,N_31162);
and U33263 (N_33263,N_30657,N_30479);
xor U33264 (N_33264,N_30167,N_31390);
or U33265 (N_33265,N_30360,N_30914);
or U33266 (N_33266,N_31130,N_30457);
or U33267 (N_33267,N_31813,N_30370);
xnor U33268 (N_33268,N_31296,N_30609);
and U33269 (N_33269,N_30179,N_30670);
xnor U33270 (N_33270,N_31429,N_31250);
and U33271 (N_33271,N_31867,N_31825);
or U33272 (N_33272,N_30183,N_30280);
nand U33273 (N_33273,N_30554,N_31616);
nor U33274 (N_33274,N_30244,N_30278);
nor U33275 (N_33275,N_30094,N_31677);
xor U33276 (N_33276,N_31243,N_30906);
or U33277 (N_33277,N_30795,N_30829);
nand U33278 (N_33278,N_31524,N_31556);
or U33279 (N_33279,N_31224,N_31225);
and U33280 (N_33280,N_30916,N_31959);
and U33281 (N_33281,N_30284,N_30905);
or U33282 (N_33282,N_31965,N_31227);
xnor U33283 (N_33283,N_30159,N_30096);
nand U33284 (N_33284,N_30695,N_30812);
nand U33285 (N_33285,N_30664,N_30240);
nor U33286 (N_33286,N_30709,N_31129);
and U33287 (N_33287,N_31366,N_30503);
nand U33288 (N_33288,N_31576,N_31112);
or U33289 (N_33289,N_31610,N_31997);
or U33290 (N_33290,N_30515,N_30546);
or U33291 (N_33291,N_30398,N_30181);
xnor U33292 (N_33292,N_30447,N_30458);
nand U33293 (N_33293,N_30256,N_30567);
and U33294 (N_33294,N_31253,N_31913);
or U33295 (N_33295,N_31209,N_30983);
nor U33296 (N_33296,N_31991,N_30123);
or U33297 (N_33297,N_30915,N_31732);
nor U33298 (N_33298,N_31163,N_31008);
and U33299 (N_33299,N_31942,N_30372);
xor U33300 (N_33300,N_30279,N_31272);
nand U33301 (N_33301,N_31160,N_30065);
nor U33302 (N_33302,N_31674,N_30958);
nand U33303 (N_33303,N_30429,N_30415);
and U33304 (N_33304,N_31039,N_31236);
or U33305 (N_33305,N_30310,N_31263);
xor U33306 (N_33306,N_31997,N_31053);
nor U33307 (N_33307,N_30065,N_31222);
nand U33308 (N_33308,N_31515,N_31300);
and U33309 (N_33309,N_31381,N_30261);
or U33310 (N_33310,N_30989,N_30406);
nand U33311 (N_33311,N_31849,N_31372);
xnor U33312 (N_33312,N_30700,N_31290);
and U33313 (N_33313,N_30381,N_30592);
xnor U33314 (N_33314,N_30572,N_30478);
xor U33315 (N_33315,N_30059,N_30764);
and U33316 (N_33316,N_30244,N_30491);
nor U33317 (N_33317,N_30362,N_31084);
nand U33318 (N_33318,N_30422,N_31470);
nand U33319 (N_33319,N_30229,N_30246);
and U33320 (N_33320,N_31416,N_31172);
and U33321 (N_33321,N_31955,N_30718);
nor U33322 (N_33322,N_30083,N_30249);
nor U33323 (N_33323,N_31711,N_30360);
nor U33324 (N_33324,N_31715,N_30442);
xor U33325 (N_33325,N_30851,N_31474);
and U33326 (N_33326,N_30084,N_31598);
nor U33327 (N_33327,N_31161,N_31173);
or U33328 (N_33328,N_30687,N_30587);
nor U33329 (N_33329,N_30043,N_31948);
nor U33330 (N_33330,N_31167,N_31166);
nand U33331 (N_33331,N_30027,N_31547);
xor U33332 (N_33332,N_30054,N_31505);
or U33333 (N_33333,N_31848,N_31023);
xnor U33334 (N_33334,N_30782,N_31054);
nand U33335 (N_33335,N_31026,N_30813);
xnor U33336 (N_33336,N_31797,N_31720);
nor U33337 (N_33337,N_31600,N_30115);
nand U33338 (N_33338,N_30248,N_31676);
nand U33339 (N_33339,N_30318,N_31865);
or U33340 (N_33340,N_31850,N_30760);
or U33341 (N_33341,N_30362,N_31721);
and U33342 (N_33342,N_30846,N_31179);
xnor U33343 (N_33343,N_30884,N_31999);
and U33344 (N_33344,N_30152,N_30479);
xor U33345 (N_33345,N_31806,N_31898);
and U33346 (N_33346,N_31904,N_31791);
or U33347 (N_33347,N_31019,N_30289);
and U33348 (N_33348,N_31642,N_30972);
nand U33349 (N_33349,N_31466,N_30541);
nor U33350 (N_33350,N_30891,N_31470);
nor U33351 (N_33351,N_30238,N_31965);
and U33352 (N_33352,N_31081,N_31763);
or U33353 (N_33353,N_30232,N_31007);
or U33354 (N_33354,N_30845,N_30997);
xor U33355 (N_33355,N_31761,N_31548);
and U33356 (N_33356,N_31598,N_30492);
nand U33357 (N_33357,N_30092,N_30604);
or U33358 (N_33358,N_30891,N_31087);
and U33359 (N_33359,N_30925,N_30088);
and U33360 (N_33360,N_30946,N_30455);
xor U33361 (N_33361,N_31002,N_31007);
nor U33362 (N_33362,N_30982,N_30995);
nand U33363 (N_33363,N_31812,N_30090);
xnor U33364 (N_33364,N_30470,N_30926);
xnor U33365 (N_33365,N_31239,N_31005);
or U33366 (N_33366,N_31967,N_31147);
nor U33367 (N_33367,N_30895,N_31477);
xor U33368 (N_33368,N_31178,N_31438);
nand U33369 (N_33369,N_30254,N_30517);
nor U33370 (N_33370,N_30843,N_31389);
or U33371 (N_33371,N_30428,N_30185);
nor U33372 (N_33372,N_30108,N_30521);
nor U33373 (N_33373,N_30404,N_31188);
and U33374 (N_33374,N_31587,N_31578);
or U33375 (N_33375,N_30434,N_30258);
or U33376 (N_33376,N_30414,N_30400);
nor U33377 (N_33377,N_31936,N_30218);
nand U33378 (N_33378,N_31061,N_31636);
or U33379 (N_33379,N_31449,N_30764);
and U33380 (N_33380,N_30412,N_30798);
xnor U33381 (N_33381,N_31907,N_30430);
or U33382 (N_33382,N_31376,N_31751);
or U33383 (N_33383,N_30890,N_31071);
nand U33384 (N_33384,N_31046,N_31600);
and U33385 (N_33385,N_30633,N_31643);
xnor U33386 (N_33386,N_31949,N_31231);
nor U33387 (N_33387,N_30383,N_31800);
nor U33388 (N_33388,N_30936,N_31347);
and U33389 (N_33389,N_30949,N_30043);
xor U33390 (N_33390,N_30285,N_30794);
or U33391 (N_33391,N_31307,N_30956);
nand U33392 (N_33392,N_31901,N_31205);
nor U33393 (N_33393,N_31939,N_31396);
xnor U33394 (N_33394,N_31310,N_31802);
nor U33395 (N_33395,N_31313,N_30850);
or U33396 (N_33396,N_31588,N_31564);
nor U33397 (N_33397,N_30432,N_30861);
nand U33398 (N_33398,N_31978,N_31351);
xor U33399 (N_33399,N_31934,N_31099);
nor U33400 (N_33400,N_31960,N_31088);
or U33401 (N_33401,N_31004,N_30501);
nor U33402 (N_33402,N_31832,N_30523);
or U33403 (N_33403,N_31232,N_31609);
or U33404 (N_33404,N_31438,N_31890);
and U33405 (N_33405,N_30428,N_30402);
nor U33406 (N_33406,N_31657,N_30659);
nor U33407 (N_33407,N_30792,N_31368);
xor U33408 (N_33408,N_30124,N_30382);
or U33409 (N_33409,N_31387,N_30093);
or U33410 (N_33410,N_31586,N_30181);
or U33411 (N_33411,N_30136,N_31859);
xnor U33412 (N_33412,N_31781,N_30907);
or U33413 (N_33413,N_30636,N_30138);
nand U33414 (N_33414,N_30337,N_30300);
nor U33415 (N_33415,N_30270,N_31830);
nor U33416 (N_33416,N_30055,N_31448);
and U33417 (N_33417,N_30115,N_30275);
and U33418 (N_33418,N_30658,N_31740);
or U33419 (N_33419,N_30785,N_31842);
and U33420 (N_33420,N_31193,N_31448);
and U33421 (N_33421,N_30781,N_31754);
or U33422 (N_33422,N_30974,N_30403);
or U33423 (N_33423,N_30056,N_30273);
nor U33424 (N_33424,N_31232,N_31803);
xor U33425 (N_33425,N_30657,N_31627);
or U33426 (N_33426,N_30322,N_31394);
or U33427 (N_33427,N_30843,N_30359);
or U33428 (N_33428,N_30158,N_31739);
and U33429 (N_33429,N_30166,N_30508);
nor U33430 (N_33430,N_31733,N_31734);
and U33431 (N_33431,N_31136,N_31441);
nand U33432 (N_33432,N_31605,N_31854);
or U33433 (N_33433,N_31277,N_30229);
or U33434 (N_33434,N_30700,N_31146);
nor U33435 (N_33435,N_30150,N_30671);
xnor U33436 (N_33436,N_31565,N_31409);
nand U33437 (N_33437,N_31382,N_30643);
nor U33438 (N_33438,N_31721,N_30774);
or U33439 (N_33439,N_31200,N_31770);
nor U33440 (N_33440,N_30891,N_30450);
or U33441 (N_33441,N_30522,N_31668);
nand U33442 (N_33442,N_31587,N_30934);
nor U33443 (N_33443,N_31471,N_31376);
and U33444 (N_33444,N_31766,N_31676);
xnor U33445 (N_33445,N_31970,N_30938);
and U33446 (N_33446,N_31698,N_31439);
nand U33447 (N_33447,N_31242,N_30655);
nand U33448 (N_33448,N_30314,N_30993);
or U33449 (N_33449,N_30091,N_31839);
and U33450 (N_33450,N_31930,N_31862);
nor U33451 (N_33451,N_30567,N_31667);
xnor U33452 (N_33452,N_30398,N_31658);
nand U33453 (N_33453,N_30407,N_31053);
nor U33454 (N_33454,N_30940,N_31759);
xor U33455 (N_33455,N_31286,N_30484);
or U33456 (N_33456,N_30972,N_31933);
xor U33457 (N_33457,N_31429,N_31576);
nor U33458 (N_33458,N_31343,N_31998);
xnor U33459 (N_33459,N_31573,N_31232);
nand U33460 (N_33460,N_31883,N_30817);
or U33461 (N_33461,N_30478,N_30710);
and U33462 (N_33462,N_30003,N_30060);
and U33463 (N_33463,N_31099,N_31015);
or U33464 (N_33464,N_31025,N_30404);
nor U33465 (N_33465,N_30644,N_30221);
nand U33466 (N_33466,N_30755,N_30813);
or U33467 (N_33467,N_30388,N_30074);
nand U33468 (N_33468,N_31354,N_31806);
and U33469 (N_33469,N_31021,N_30912);
nor U33470 (N_33470,N_30668,N_31858);
and U33471 (N_33471,N_30277,N_31109);
nor U33472 (N_33472,N_30793,N_30523);
or U33473 (N_33473,N_31023,N_31499);
and U33474 (N_33474,N_31654,N_31624);
nand U33475 (N_33475,N_31144,N_31821);
nor U33476 (N_33476,N_31018,N_31552);
or U33477 (N_33477,N_31239,N_31695);
and U33478 (N_33478,N_31586,N_31786);
xnor U33479 (N_33479,N_31173,N_31772);
and U33480 (N_33480,N_31832,N_31811);
nor U33481 (N_33481,N_31220,N_30773);
nand U33482 (N_33482,N_30877,N_30684);
and U33483 (N_33483,N_31690,N_30476);
nand U33484 (N_33484,N_31099,N_31393);
or U33485 (N_33485,N_31629,N_31454);
or U33486 (N_33486,N_30271,N_31322);
and U33487 (N_33487,N_30190,N_30587);
nand U33488 (N_33488,N_31963,N_31952);
and U33489 (N_33489,N_30882,N_30848);
and U33490 (N_33490,N_30409,N_31318);
and U33491 (N_33491,N_31483,N_31429);
or U33492 (N_33492,N_31712,N_31358);
or U33493 (N_33493,N_31595,N_30805);
xor U33494 (N_33494,N_30067,N_30037);
or U33495 (N_33495,N_31858,N_30988);
nor U33496 (N_33496,N_31717,N_31939);
and U33497 (N_33497,N_30925,N_30033);
and U33498 (N_33498,N_31965,N_31239);
nor U33499 (N_33499,N_31332,N_31860);
nand U33500 (N_33500,N_31683,N_30938);
xor U33501 (N_33501,N_30561,N_31212);
and U33502 (N_33502,N_30485,N_30870);
or U33503 (N_33503,N_30416,N_31499);
and U33504 (N_33504,N_31726,N_30129);
xnor U33505 (N_33505,N_31160,N_30430);
nand U33506 (N_33506,N_30423,N_31201);
and U33507 (N_33507,N_31361,N_31206);
nor U33508 (N_33508,N_31418,N_31875);
or U33509 (N_33509,N_31685,N_30949);
or U33510 (N_33510,N_31941,N_31333);
or U33511 (N_33511,N_30466,N_31354);
nor U33512 (N_33512,N_30652,N_30962);
xor U33513 (N_33513,N_31651,N_31649);
xnor U33514 (N_33514,N_30125,N_30103);
xnor U33515 (N_33515,N_30350,N_31162);
xor U33516 (N_33516,N_31993,N_31456);
nand U33517 (N_33517,N_30796,N_30584);
nor U33518 (N_33518,N_31674,N_31404);
xor U33519 (N_33519,N_31196,N_30774);
nand U33520 (N_33520,N_30574,N_30372);
nor U33521 (N_33521,N_31633,N_31409);
nand U33522 (N_33522,N_30013,N_30505);
and U33523 (N_33523,N_31666,N_30144);
and U33524 (N_33524,N_31704,N_31834);
or U33525 (N_33525,N_30195,N_31972);
xor U33526 (N_33526,N_31931,N_30972);
or U33527 (N_33527,N_30332,N_30564);
nor U33528 (N_33528,N_30627,N_30874);
or U33529 (N_33529,N_30946,N_31413);
nand U33530 (N_33530,N_30816,N_30350);
and U33531 (N_33531,N_31883,N_31921);
and U33532 (N_33532,N_30466,N_31522);
or U33533 (N_33533,N_30083,N_30824);
and U33534 (N_33534,N_30712,N_31197);
nor U33535 (N_33535,N_31813,N_31386);
nand U33536 (N_33536,N_30284,N_31914);
nand U33537 (N_33537,N_30844,N_30722);
xor U33538 (N_33538,N_30571,N_31444);
xor U33539 (N_33539,N_30015,N_31134);
xnor U33540 (N_33540,N_31240,N_30152);
and U33541 (N_33541,N_30832,N_30543);
xnor U33542 (N_33542,N_31464,N_31727);
or U33543 (N_33543,N_30217,N_30603);
and U33544 (N_33544,N_30974,N_31477);
nor U33545 (N_33545,N_31323,N_31829);
and U33546 (N_33546,N_31727,N_30328);
nor U33547 (N_33547,N_31166,N_31312);
nor U33548 (N_33548,N_31908,N_31558);
nand U33549 (N_33549,N_30574,N_30867);
nand U33550 (N_33550,N_30935,N_30584);
or U33551 (N_33551,N_30021,N_30353);
nand U33552 (N_33552,N_30804,N_30225);
and U33553 (N_33553,N_31392,N_30039);
xnor U33554 (N_33554,N_31417,N_30870);
and U33555 (N_33555,N_30804,N_30476);
nand U33556 (N_33556,N_31803,N_30720);
and U33557 (N_33557,N_31899,N_31608);
nand U33558 (N_33558,N_30850,N_31989);
xor U33559 (N_33559,N_31238,N_31434);
nor U33560 (N_33560,N_31839,N_30066);
nand U33561 (N_33561,N_30027,N_31536);
nor U33562 (N_33562,N_30284,N_31382);
xor U33563 (N_33563,N_30472,N_31639);
nand U33564 (N_33564,N_30392,N_30756);
nor U33565 (N_33565,N_30658,N_31288);
nand U33566 (N_33566,N_30814,N_30005);
nor U33567 (N_33567,N_30229,N_31137);
or U33568 (N_33568,N_31041,N_31203);
nor U33569 (N_33569,N_30294,N_30404);
or U33570 (N_33570,N_30342,N_30009);
xor U33571 (N_33571,N_30578,N_31302);
nand U33572 (N_33572,N_31941,N_30012);
and U33573 (N_33573,N_31452,N_30741);
xor U33574 (N_33574,N_30345,N_30272);
and U33575 (N_33575,N_31146,N_30894);
and U33576 (N_33576,N_31248,N_30401);
xnor U33577 (N_33577,N_31811,N_30712);
or U33578 (N_33578,N_31784,N_30841);
and U33579 (N_33579,N_30023,N_30176);
xnor U33580 (N_33580,N_30235,N_30309);
nor U33581 (N_33581,N_30609,N_30009);
xor U33582 (N_33582,N_31042,N_30686);
xnor U33583 (N_33583,N_31542,N_30108);
and U33584 (N_33584,N_31664,N_31246);
nand U33585 (N_33585,N_31622,N_30855);
and U33586 (N_33586,N_31500,N_31514);
nand U33587 (N_33587,N_31407,N_30795);
xor U33588 (N_33588,N_31695,N_31450);
nor U33589 (N_33589,N_31021,N_31691);
nand U33590 (N_33590,N_30358,N_31788);
or U33591 (N_33591,N_30085,N_30922);
xor U33592 (N_33592,N_31767,N_30504);
nor U33593 (N_33593,N_30181,N_30515);
nor U33594 (N_33594,N_31851,N_30231);
and U33595 (N_33595,N_31860,N_31740);
and U33596 (N_33596,N_31862,N_30925);
xnor U33597 (N_33597,N_31112,N_31443);
nand U33598 (N_33598,N_30955,N_30144);
nor U33599 (N_33599,N_30316,N_31305);
and U33600 (N_33600,N_30505,N_31829);
xor U33601 (N_33601,N_31524,N_30388);
nor U33602 (N_33602,N_31160,N_30887);
nor U33603 (N_33603,N_31201,N_31144);
xnor U33604 (N_33604,N_31418,N_31309);
xnor U33605 (N_33605,N_31077,N_30915);
xnor U33606 (N_33606,N_30011,N_30648);
or U33607 (N_33607,N_31776,N_31766);
nor U33608 (N_33608,N_30191,N_31729);
nand U33609 (N_33609,N_30628,N_31650);
nand U33610 (N_33610,N_31382,N_30314);
and U33611 (N_33611,N_30733,N_30896);
or U33612 (N_33612,N_31148,N_31366);
or U33613 (N_33613,N_31528,N_31763);
and U33614 (N_33614,N_30034,N_30630);
nand U33615 (N_33615,N_30429,N_30546);
or U33616 (N_33616,N_30850,N_30914);
xnor U33617 (N_33617,N_31525,N_31379);
and U33618 (N_33618,N_30854,N_30595);
and U33619 (N_33619,N_31795,N_30069);
nand U33620 (N_33620,N_31408,N_31793);
or U33621 (N_33621,N_31359,N_31341);
and U33622 (N_33622,N_31742,N_30520);
or U33623 (N_33623,N_31956,N_30653);
nor U33624 (N_33624,N_31524,N_30780);
and U33625 (N_33625,N_31300,N_30251);
nand U33626 (N_33626,N_31080,N_31204);
nand U33627 (N_33627,N_30537,N_30191);
and U33628 (N_33628,N_31604,N_30420);
nor U33629 (N_33629,N_30313,N_31830);
nor U33630 (N_33630,N_31669,N_30030);
and U33631 (N_33631,N_31612,N_30017);
nand U33632 (N_33632,N_30493,N_30258);
nor U33633 (N_33633,N_30807,N_30392);
xnor U33634 (N_33634,N_30303,N_31107);
xnor U33635 (N_33635,N_31477,N_30621);
and U33636 (N_33636,N_31226,N_30808);
xnor U33637 (N_33637,N_31990,N_31915);
and U33638 (N_33638,N_30740,N_30365);
or U33639 (N_33639,N_31002,N_31371);
xnor U33640 (N_33640,N_30279,N_31213);
xnor U33641 (N_33641,N_30312,N_31301);
and U33642 (N_33642,N_31994,N_30961);
nor U33643 (N_33643,N_31186,N_30241);
and U33644 (N_33644,N_30158,N_31968);
nor U33645 (N_33645,N_31538,N_31703);
nand U33646 (N_33646,N_31545,N_31517);
xnor U33647 (N_33647,N_30694,N_31475);
or U33648 (N_33648,N_31266,N_31883);
nor U33649 (N_33649,N_31970,N_30904);
nand U33650 (N_33650,N_30312,N_30391);
and U33651 (N_33651,N_30793,N_30096);
nor U33652 (N_33652,N_31284,N_30012);
or U33653 (N_33653,N_31283,N_31727);
or U33654 (N_33654,N_30612,N_31877);
nand U33655 (N_33655,N_31522,N_30681);
nand U33656 (N_33656,N_30104,N_31810);
nor U33657 (N_33657,N_31248,N_30167);
or U33658 (N_33658,N_31188,N_30137);
xnor U33659 (N_33659,N_30325,N_30941);
and U33660 (N_33660,N_31888,N_30189);
nand U33661 (N_33661,N_31768,N_31827);
or U33662 (N_33662,N_31642,N_31317);
xnor U33663 (N_33663,N_30782,N_30573);
nor U33664 (N_33664,N_31950,N_30029);
nor U33665 (N_33665,N_30270,N_30532);
nand U33666 (N_33666,N_30863,N_30234);
xor U33667 (N_33667,N_31476,N_30504);
nand U33668 (N_33668,N_31943,N_31850);
and U33669 (N_33669,N_30548,N_31768);
nor U33670 (N_33670,N_31538,N_30863);
xor U33671 (N_33671,N_31357,N_30820);
and U33672 (N_33672,N_30477,N_31969);
nand U33673 (N_33673,N_31664,N_31641);
nand U33674 (N_33674,N_30536,N_30373);
xor U33675 (N_33675,N_30358,N_30474);
and U33676 (N_33676,N_30192,N_31446);
and U33677 (N_33677,N_30668,N_31616);
nor U33678 (N_33678,N_30155,N_31722);
xnor U33679 (N_33679,N_30510,N_31625);
or U33680 (N_33680,N_30658,N_30152);
or U33681 (N_33681,N_30807,N_31668);
nor U33682 (N_33682,N_31555,N_30694);
xnor U33683 (N_33683,N_31191,N_31858);
xor U33684 (N_33684,N_31341,N_31571);
nand U33685 (N_33685,N_31818,N_31860);
and U33686 (N_33686,N_30760,N_31202);
nor U33687 (N_33687,N_30917,N_31642);
nand U33688 (N_33688,N_31231,N_31309);
nand U33689 (N_33689,N_30669,N_30339);
xnor U33690 (N_33690,N_30415,N_30109);
or U33691 (N_33691,N_30879,N_31370);
xnor U33692 (N_33692,N_31471,N_30984);
and U33693 (N_33693,N_31887,N_30677);
nand U33694 (N_33694,N_31418,N_30038);
xnor U33695 (N_33695,N_30660,N_30599);
xor U33696 (N_33696,N_30893,N_31589);
nor U33697 (N_33697,N_30051,N_30956);
or U33698 (N_33698,N_31523,N_30649);
nor U33699 (N_33699,N_31079,N_31204);
xnor U33700 (N_33700,N_31497,N_31566);
and U33701 (N_33701,N_30331,N_31263);
nor U33702 (N_33702,N_30552,N_31007);
and U33703 (N_33703,N_30201,N_30727);
nor U33704 (N_33704,N_30137,N_30709);
nor U33705 (N_33705,N_30655,N_31253);
nand U33706 (N_33706,N_30126,N_31856);
or U33707 (N_33707,N_30180,N_31019);
xnor U33708 (N_33708,N_31481,N_31636);
or U33709 (N_33709,N_30080,N_30369);
nand U33710 (N_33710,N_30319,N_31211);
and U33711 (N_33711,N_31994,N_30432);
or U33712 (N_33712,N_31137,N_30153);
nor U33713 (N_33713,N_30243,N_30846);
xnor U33714 (N_33714,N_30507,N_30097);
xnor U33715 (N_33715,N_31715,N_30884);
xnor U33716 (N_33716,N_31868,N_31481);
nand U33717 (N_33717,N_31678,N_31758);
nor U33718 (N_33718,N_31113,N_31107);
nor U33719 (N_33719,N_31136,N_31529);
nand U33720 (N_33720,N_31830,N_31703);
xor U33721 (N_33721,N_30242,N_31027);
nor U33722 (N_33722,N_31969,N_31454);
or U33723 (N_33723,N_31179,N_30196);
or U33724 (N_33724,N_31045,N_30353);
or U33725 (N_33725,N_31438,N_31982);
nand U33726 (N_33726,N_31148,N_31283);
and U33727 (N_33727,N_30487,N_30550);
or U33728 (N_33728,N_30976,N_30890);
or U33729 (N_33729,N_30679,N_30459);
or U33730 (N_33730,N_30807,N_31407);
and U33731 (N_33731,N_31615,N_31873);
xor U33732 (N_33732,N_31767,N_30147);
nand U33733 (N_33733,N_31222,N_30572);
xor U33734 (N_33734,N_31454,N_30415);
and U33735 (N_33735,N_31433,N_30347);
or U33736 (N_33736,N_31682,N_30191);
and U33737 (N_33737,N_30769,N_30764);
xnor U33738 (N_33738,N_30539,N_30274);
nor U33739 (N_33739,N_31024,N_31910);
nand U33740 (N_33740,N_31196,N_31824);
or U33741 (N_33741,N_31412,N_31335);
nor U33742 (N_33742,N_30214,N_30488);
nand U33743 (N_33743,N_31269,N_30229);
or U33744 (N_33744,N_31862,N_30125);
xnor U33745 (N_33745,N_31755,N_31783);
nand U33746 (N_33746,N_30231,N_30616);
nor U33747 (N_33747,N_30832,N_30532);
and U33748 (N_33748,N_30916,N_30213);
or U33749 (N_33749,N_30560,N_30612);
xor U33750 (N_33750,N_30625,N_30596);
nor U33751 (N_33751,N_30463,N_31356);
nor U33752 (N_33752,N_31673,N_31328);
or U33753 (N_33753,N_31802,N_31252);
xor U33754 (N_33754,N_30787,N_30573);
or U33755 (N_33755,N_30154,N_31912);
xnor U33756 (N_33756,N_31970,N_31962);
xor U33757 (N_33757,N_31315,N_30814);
or U33758 (N_33758,N_31416,N_30965);
or U33759 (N_33759,N_31520,N_30230);
xor U33760 (N_33760,N_31643,N_31268);
xor U33761 (N_33761,N_30338,N_31231);
nor U33762 (N_33762,N_30728,N_30802);
or U33763 (N_33763,N_31018,N_31945);
xnor U33764 (N_33764,N_31374,N_30441);
and U33765 (N_33765,N_30953,N_31919);
nor U33766 (N_33766,N_30681,N_30084);
and U33767 (N_33767,N_30031,N_31950);
nor U33768 (N_33768,N_30835,N_30302);
nand U33769 (N_33769,N_30749,N_30975);
xor U33770 (N_33770,N_30817,N_31911);
or U33771 (N_33771,N_31161,N_30883);
xnor U33772 (N_33772,N_31419,N_31896);
and U33773 (N_33773,N_31279,N_30318);
xor U33774 (N_33774,N_31546,N_31533);
or U33775 (N_33775,N_31075,N_31497);
xor U33776 (N_33776,N_31284,N_30915);
or U33777 (N_33777,N_30199,N_30361);
and U33778 (N_33778,N_30469,N_30438);
and U33779 (N_33779,N_30568,N_30293);
xor U33780 (N_33780,N_30437,N_31803);
nand U33781 (N_33781,N_31024,N_30756);
nor U33782 (N_33782,N_30509,N_30514);
and U33783 (N_33783,N_31761,N_31511);
nor U33784 (N_33784,N_31421,N_30116);
nor U33785 (N_33785,N_31359,N_31038);
nand U33786 (N_33786,N_31630,N_31344);
nor U33787 (N_33787,N_30255,N_31227);
and U33788 (N_33788,N_31155,N_30022);
and U33789 (N_33789,N_30397,N_30832);
nand U33790 (N_33790,N_30522,N_31199);
nand U33791 (N_33791,N_30980,N_30457);
xnor U33792 (N_33792,N_31814,N_31271);
nor U33793 (N_33793,N_31675,N_30236);
nand U33794 (N_33794,N_31491,N_30700);
and U33795 (N_33795,N_30700,N_31528);
nand U33796 (N_33796,N_31586,N_31144);
nand U33797 (N_33797,N_30243,N_30406);
or U33798 (N_33798,N_31555,N_31922);
nand U33799 (N_33799,N_30440,N_30365);
or U33800 (N_33800,N_30439,N_30945);
and U33801 (N_33801,N_31207,N_30093);
xor U33802 (N_33802,N_30116,N_30675);
nor U33803 (N_33803,N_30505,N_31588);
or U33804 (N_33804,N_31744,N_30630);
nand U33805 (N_33805,N_30662,N_31780);
or U33806 (N_33806,N_30669,N_31569);
and U33807 (N_33807,N_31873,N_30032);
and U33808 (N_33808,N_31728,N_31945);
nand U33809 (N_33809,N_30134,N_31302);
or U33810 (N_33810,N_31125,N_31396);
nor U33811 (N_33811,N_30920,N_31231);
nand U33812 (N_33812,N_30556,N_30760);
or U33813 (N_33813,N_31856,N_31917);
xor U33814 (N_33814,N_30079,N_30932);
xor U33815 (N_33815,N_30789,N_30917);
xor U33816 (N_33816,N_31597,N_30634);
nand U33817 (N_33817,N_31708,N_30895);
and U33818 (N_33818,N_31424,N_30054);
nor U33819 (N_33819,N_31849,N_31827);
xnor U33820 (N_33820,N_31277,N_31761);
and U33821 (N_33821,N_31565,N_30433);
and U33822 (N_33822,N_31602,N_31964);
nor U33823 (N_33823,N_30083,N_31136);
nor U33824 (N_33824,N_31329,N_31548);
xor U33825 (N_33825,N_31280,N_31942);
xor U33826 (N_33826,N_30593,N_31121);
xnor U33827 (N_33827,N_31942,N_31425);
or U33828 (N_33828,N_30493,N_30201);
nand U33829 (N_33829,N_31486,N_30792);
and U33830 (N_33830,N_31616,N_30088);
xnor U33831 (N_33831,N_31164,N_30465);
nor U33832 (N_33832,N_30625,N_31649);
nand U33833 (N_33833,N_31359,N_31180);
and U33834 (N_33834,N_30071,N_30760);
xnor U33835 (N_33835,N_30534,N_31796);
nor U33836 (N_33836,N_30603,N_30508);
nor U33837 (N_33837,N_31892,N_31906);
xor U33838 (N_33838,N_31729,N_30986);
nor U33839 (N_33839,N_30580,N_30019);
xor U33840 (N_33840,N_30438,N_31194);
nand U33841 (N_33841,N_31505,N_31863);
nor U33842 (N_33842,N_30071,N_30811);
and U33843 (N_33843,N_31936,N_31343);
and U33844 (N_33844,N_30078,N_31883);
xnor U33845 (N_33845,N_31335,N_30631);
nand U33846 (N_33846,N_31383,N_30833);
xor U33847 (N_33847,N_31173,N_31454);
and U33848 (N_33848,N_31913,N_30882);
nor U33849 (N_33849,N_31392,N_31264);
or U33850 (N_33850,N_31948,N_30919);
xor U33851 (N_33851,N_31151,N_31793);
nand U33852 (N_33852,N_31266,N_31732);
nand U33853 (N_33853,N_31070,N_30035);
nor U33854 (N_33854,N_31013,N_31357);
nor U33855 (N_33855,N_30070,N_31007);
xnor U33856 (N_33856,N_31375,N_30773);
and U33857 (N_33857,N_31326,N_31422);
nand U33858 (N_33858,N_31218,N_31515);
nor U33859 (N_33859,N_30507,N_30476);
xnor U33860 (N_33860,N_31981,N_31968);
nand U33861 (N_33861,N_30019,N_31906);
nor U33862 (N_33862,N_30758,N_30450);
nor U33863 (N_33863,N_31011,N_31706);
xnor U33864 (N_33864,N_30889,N_31788);
or U33865 (N_33865,N_31072,N_31375);
xnor U33866 (N_33866,N_30331,N_31243);
xor U33867 (N_33867,N_31637,N_31581);
nor U33868 (N_33868,N_31329,N_30583);
or U33869 (N_33869,N_31580,N_31669);
xnor U33870 (N_33870,N_30994,N_30152);
or U33871 (N_33871,N_31115,N_30051);
nor U33872 (N_33872,N_30489,N_31536);
nand U33873 (N_33873,N_30166,N_31572);
nor U33874 (N_33874,N_30598,N_31095);
and U33875 (N_33875,N_31085,N_31224);
nand U33876 (N_33876,N_31905,N_30390);
and U33877 (N_33877,N_31256,N_30389);
nand U33878 (N_33878,N_31531,N_31880);
nand U33879 (N_33879,N_30532,N_30484);
and U33880 (N_33880,N_30220,N_30707);
nand U33881 (N_33881,N_30010,N_31364);
and U33882 (N_33882,N_31554,N_30453);
nor U33883 (N_33883,N_30008,N_30170);
and U33884 (N_33884,N_30751,N_30792);
or U33885 (N_33885,N_31406,N_31317);
nand U33886 (N_33886,N_31689,N_31990);
or U33887 (N_33887,N_31313,N_31081);
xnor U33888 (N_33888,N_31600,N_31378);
and U33889 (N_33889,N_30394,N_30483);
nor U33890 (N_33890,N_31946,N_31319);
and U33891 (N_33891,N_30959,N_30913);
nand U33892 (N_33892,N_31537,N_31629);
and U33893 (N_33893,N_30343,N_31845);
and U33894 (N_33894,N_31230,N_31216);
nand U33895 (N_33895,N_30034,N_30187);
xor U33896 (N_33896,N_30075,N_31013);
nor U33897 (N_33897,N_30021,N_31035);
nor U33898 (N_33898,N_31117,N_30359);
nor U33899 (N_33899,N_30734,N_31568);
xnor U33900 (N_33900,N_30897,N_30103);
and U33901 (N_33901,N_30015,N_31115);
nand U33902 (N_33902,N_31501,N_31889);
nor U33903 (N_33903,N_31193,N_31720);
and U33904 (N_33904,N_31026,N_30154);
nand U33905 (N_33905,N_30044,N_30308);
and U33906 (N_33906,N_30426,N_31572);
nand U33907 (N_33907,N_31263,N_30641);
and U33908 (N_33908,N_30732,N_31783);
and U33909 (N_33909,N_31313,N_31117);
xnor U33910 (N_33910,N_30155,N_30486);
or U33911 (N_33911,N_31123,N_30010);
nor U33912 (N_33912,N_31181,N_30692);
xnor U33913 (N_33913,N_30291,N_30185);
nor U33914 (N_33914,N_30643,N_30913);
nor U33915 (N_33915,N_30652,N_30775);
and U33916 (N_33916,N_31520,N_30287);
or U33917 (N_33917,N_31157,N_30370);
and U33918 (N_33918,N_31259,N_30027);
or U33919 (N_33919,N_31144,N_31264);
nor U33920 (N_33920,N_31101,N_30716);
or U33921 (N_33921,N_31193,N_30266);
xnor U33922 (N_33922,N_30728,N_31425);
nor U33923 (N_33923,N_30891,N_31541);
or U33924 (N_33924,N_31813,N_31891);
xor U33925 (N_33925,N_30912,N_30097);
or U33926 (N_33926,N_31042,N_30943);
nor U33927 (N_33927,N_31523,N_31039);
xnor U33928 (N_33928,N_30560,N_31782);
nand U33929 (N_33929,N_30830,N_30697);
or U33930 (N_33930,N_30756,N_30940);
and U33931 (N_33931,N_31712,N_31837);
or U33932 (N_33932,N_31896,N_30626);
and U33933 (N_33933,N_31296,N_30396);
or U33934 (N_33934,N_30065,N_31131);
and U33935 (N_33935,N_31975,N_31044);
xnor U33936 (N_33936,N_30640,N_31884);
or U33937 (N_33937,N_31899,N_30711);
nand U33938 (N_33938,N_31488,N_31378);
nor U33939 (N_33939,N_31207,N_30591);
xnor U33940 (N_33940,N_31776,N_30015);
nand U33941 (N_33941,N_31158,N_31347);
nand U33942 (N_33942,N_31607,N_31667);
and U33943 (N_33943,N_30450,N_31996);
and U33944 (N_33944,N_31536,N_31961);
nand U33945 (N_33945,N_31501,N_31193);
or U33946 (N_33946,N_31455,N_31783);
and U33947 (N_33947,N_31852,N_31956);
or U33948 (N_33948,N_31534,N_31132);
xnor U33949 (N_33949,N_30796,N_30162);
and U33950 (N_33950,N_30343,N_30309);
or U33951 (N_33951,N_31052,N_31332);
or U33952 (N_33952,N_30801,N_30189);
xnor U33953 (N_33953,N_30405,N_30737);
or U33954 (N_33954,N_30688,N_30932);
nor U33955 (N_33955,N_31506,N_30368);
or U33956 (N_33956,N_31377,N_31168);
nor U33957 (N_33957,N_30629,N_31340);
or U33958 (N_33958,N_30956,N_31207);
nand U33959 (N_33959,N_31055,N_31661);
nand U33960 (N_33960,N_31896,N_30650);
and U33961 (N_33961,N_31411,N_31549);
xnor U33962 (N_33962,N_31978,N_31080);
nand U33963 (N_33963,N_30027,N_31190);
nand U33964 (N_33964,N_30545,N_31138);
or U33965 (N_33965,N_30148,N_30513);
and U33966 (N_33966,N_31025,N_30448);
nor U33967 (N_33967,N_31731,N_31403);
nand U33968 (N_33968,N_31499,N_30568);
and U33969 (N_33969,N_31712,N_31324);
nand U33970 (N_33970,N_31651,N_31429);
nor U33971 (N_33971,N_31232,N_30030);
xnor U33972 (N_33972,N_30713,N_30192);
or U33973 (N_33973,N_31760,N_30530);
xnor U33974 (N_33974,N_31779,N_31480);
and U33975 (N_33975,N_31558,N_31495);
and U33976 (N_33976,N_30466,N_31214);
nand U33977 (N_33977,N_31227,N_31683);
or U33978 (N_33978,N_30784,N_30157);
xnor U33979 (N_33979,N_30925,N_30220);
or U33980 (N_33980,N_30148,N_30941);
nand U33981 (N_33981,N_31187,N_30447);
nand U33982 (N_33982,N_31601,N_31066);
or U33983 (N_33983,N_31744,N_31342);
xor U33984 (N_33984,N_31215,N_30403);
nand U33985 (N_33985,N_30173,N_31469);
nor U33986 (N_33986,N_31851,N_30770);
or U33987 (N_33987,N_31164,N_30935);
and U33988 (N_33988,N_30559,N_30168);
and U33989 (N_33989,N_31304,N_31190);
xnor U33990 (N_33990,N_31430,N_31290);
nand U33991 (N_33991,N_31704,N_31930);
nor U33992 (N_33992,N_30195,N_31441);
nand U33993 (N_33993,N_31449,N_31849);
or U33994 (N_33994,N_30281,N_30866);
xor U33995 (N_33995,N_31825,N_30878);
nand U33996 (N_33996,N_31324,N_30883);
nand U33997 (N_33997,N_30483,N_31269);
or U33998 (N_33998,N_30459,N_31493);
nor U33999 (N_33999,N_30043,N_30069);
and U34000 (N_34000,N_33408,N_32766);
nand U34001 (N_34001,N_32627,N_33739);
nand U34002 (N_34002,N_32964,N_33835);
and U34003 (N_34003,N_33565,N_33079);
and U34004 (N_34004,N_32296,N_32815);
and U34005 (N_34005,N_33412,N_32406);
nand U34006 (N_34006,N_32929,N_33826);
and U34007 (N_34007,N_32449,N_32615);
nand U34008 (N_34008,N_33955,N_32765);
nand U34009 (N_34009,N_32890,N_32813);
or U34010 (N_34010,N_33753,N_33794);
or U34011 (N_34011,N_33454,N_33623);
xor U34012 (N_34012,N_32421,N_33076);
and U34013 (N_34013,N_33866,N_33629);
and U34014 (N_34014,N_33677,N_33364);
xor U34015 (N_34015,N_33429,N_33875);
nand U34016 (N_34016,N_33821,N_32703);
nor U34017 (N_34017,N_33208,N_32363);
nor U34018 (N_34018,N_33437,N_33746);
xnor U34019 (N_34019,N_33928,N_32188);
and U34020 (N_34020,N_33799,N_32844);
xnor U34021 (N_34021,N_32286,N_33180);
xnor U34022 (N_34022,N_33787,N_32169);
nand U34023 (N_34023,N_33413,N_32837);
nor U34024 (N_34024,N_32331,N_32553);
or U34025 (N_34025,N_33020,N_33756);
and U34026 (N_34026,N_33555,N_33811);
nand U34027 (N_34027,N_33196,N_32109);
and U34028 (N_34028,N_33450,N_33231);
xnor U34029 (N_34029,N_33944,N_33065);
and U34030 (N_34030,N_33315,N_33127);
nand U34031 (N_34031,N_32757,N_33625);
or U34032 (N_34032,N_32616,N_32751);
and U34033 (N_34033,N_32504,N_33317);
nor U34034 (N_34034,N_32263,N_33604);
nor U34035 (N_34035,N_32448,N_32843);
nand U34036 (N_34036,N_33877,N_33529);
or U34037 (N_34037,N_33782,N_32785);
or U34038 (N_34038,N_32271,N_33340);
or U34039 (N_34039,N_32937,N_32381);
xnor U34040 (N_34040,N_33074,N_32170);
or U34041 (N_34041,N_32254,N_32958);
or U34042 (N_34042,N_32425,N_32239);
and U34043 (N_34043,N_32255,N_33102);
nor U34044 (N_34044,N_32943,N_32322);
nand U34045 (N_34045,N_32027,N_32799);
nand U34046 (N_34046,N_32171,N_32514);
nand U34047 (N_34047,N_33702,N_32942);
nor U34048 (N_34048,N_32199,N_33054);
xnor U34049 (N_34049,N_33873,N_32278);
and U34050 (N_34050,N_32544,N_32293);
nor U34051 (N_34051,N_33058,N_32490);
and U34052 (N_34052,N_32212,N_33912);
xor U34053 (N_34053,N_33311,N_33047);
xor U34054 (N_34054,N_33716,N_33606);
xnor U34055 (N_34055,N_33598,N_33655);
nand U34056 (N_34056,N_32059,N_33991);
or U34057 (N_34057,N_32165,N_32782);
and U34058 (N_34058,N_32618,N_33964);
and U34059 (N_34059,N_33736,N_33949);
xor U34060 (N_34060,N_32262,N_33612);
or U34061 (N_34061,N_33176,N_33789);
xnor U34062 (N_34062,N_32226,N_33356);
nand U34063 (N_34063,N_33148,N_32619);
nor U34064 (N_34064,N_33933,N_32506);
nand U34065 (N_34065,N_32326,N_33684);
or U34066 (N_34066,N_32824,N_32249);
and U34067 (N_34067,N_33734,N_32728);
nor U34068 (N_34068,N_33399,N_32145);
and U34069 (N_34069,N_32368,N_33740);
and U34070 (N_34070,N_33320,N_33915);
nand U34071 (N_34071,N_33774,N_32695);
and U34072 (N_34072,N_33041,N_33888);
and U34073 (N_34073,N_32519,N_32614);
or U34074 (N_34074,N_33220,N_33330);
and U34075 (N_34075,N_32045,N_33378);
nand U34076 (N_34076,N_33885,N_33318);
xor U34077 (N_34077,N_32489,N_32159);
nand U34078 (N_34078,N_33430,N_33287);
xnor U34079 (N_34079,N_33584,N_32768);
nor U34080 (N_34080,N_33168,N_32918);
or U34081 (N_34081,N_32346,N_32702);
and U34082 (N_34082,N_33733,N_32749);
nand U34083 (N_34083,N_33741,N_32949);
or U34084 (N_34084,N_32984,N_32353);
and U34085 (N_34085,N_33502,N_32719);
or U34086 (N_34086,N_33276,N_32847);
or U34087 (N_34087,N_32788,N_33626);
xnor U34088 (N_34088,N_33152,N_33762);
and U34089 (N_34089,N_33910,N_32342);
nand U34090 (N_34090,N_33042,N_33331);
xor U34091 (N_34091,N_33832,N_32442);
nand U34092 (N_34092,N_33198,N_32172);
nor U34093 (N_34093,N_33478,N_32272);
nand U34094 (N_34094,N_32976,N_33243);
xor U34095 (N_34095,N_32892,N_32561);
nand U34096 (N_34096,N_33228,N_32667);
and U34097 (N_34097,N_32083,N_32318);
and U34098 (N_34098,N_33934,N_32870);
xnor U34099 (N_34099,N_32157,N_33669);
nand U34100 (N_34100,N_32674,N_32312);
nand U34101 (N_34101,N_32806,N_33167);
xnor U34102 (N_34102,N_32284,N_32040);
xnor U34103 (N_34103,N_32499,N_33937);
nor U34104 (N_34104,N_32812,N_32657);
and U34105 (N_34105,N_32273,N_32717);
nor U34106 (N_34106,N_33162,N_33987);
nand U34107 (N_34107,N_33186,N_32335);
nand U34108 (N_34108,N_32683,N_32969);
and U34109 (N_34109,N_33824,N_33301);
xnor U34110 (N_34110,N_32712,N_32380);
nand U34111 (N_34111,N_32537,N_32781);
nand U34112 (N_34112,N_33678,N_32966);
xnor U34113 (N_34113,N_33793,N_33822);
nor U34114 (N_34114,N_33978,N_32733);
nor U34115 (N_34115,N_32938,N_32513);
and U34116 (N_34116,N_32025,N_33798);
nor U34117 (N_34117,N_33253,N_33769);
or U34118 (N_34118,N_33113,N_33840);
xnor U34119 (N_34119,N_32316,N_32891);
nand U34120 (N_34120,N_32809,N_32395);
nand U34121 (N_34121,N_32961,N_32413);
xnor U34122 (N_34122,N_32432,N_33707);
nor U34123 (N_34123,N_33174,N_32336);
and U34124 (N_34124,N_32978,N_33270);
nor U34125 (N_34125,N_33022,N_33993);
xnor U34126 (N_34126,N_32191,N_33215);
nand U34127 (N_34127,N_32600,N_32037);
and U34128 (N_34128,N_32577,N_32839);
or U34129 (N_34129,N_33969,N_32258);
and U34130 (N_34130,N_32126,N_33384);
and U34131 (N_34131,N_33434,N_33357);
nand U34132 (N_34132,N_32210,N_32285);
nor U34133 (N_34133,N_33683,N_33803);
nand U34134 (N_34134,N_33752,N_32608);
and U34135 (N_34135,N_33570,N_32810);
xnor U34136 (N_34136,N_33713,N_32041);
nand U34137 (N_34137,N_32310,N_32595);
xor U34138 (N_34138,N_32769,N_32581);
nor U34139 (N_34139,N_32244,N_33857);
or U34140 (N_34140,N_33979,N_33652);
or U34141 (N_34141,N_32078,N_33021);
and U34142 (N_34142,N_33804,N_32545);
nor U34143 (N_34143,N_33305,N_33134);
or U34144 (N_34144,N_33348,N_32686);
xnor U34145 (N_34145,N_32012,N_33948);
nand U34146 (N_34146,N_32364,N_33362);
and U34147 (N_34147,N_32452,N_33552);
and U34148 (N_34148,N_33776,N_32510);
and U34149 (N_34149,N_33100,N_33585);
and U34150 (N_34150,N_33003,N_32721);
and U34151 (N_34151,N_33532,N_32206);
nor U34152 (N_34152,N_33862,N_33423);
or U34153 (N_34153,N_32731,N_33459);
nand U34154 (N_34154,N_33656,N_33238);
and U34155 (N_34155,N_33997,N_33269);
or U34156 (N_34156,N_32358,N_33105);
or U34157 (N_34157,N_32086,N_32885);
xnor U34158 (N_34158,N_32645,N_32687);
xor U34159 (N_34159,N_33420,N_33867);
xnor U34160 (N_34160,N_32689,N_32981);
or U34161 (N_34161,N_32582,N_32487);
xnor U34162 (N_34162,N_33551,N_33114);
and U34163 (N_34163,N_32662,N_33073);
nand U34164 (N_34164,N_33919,N_32174);
and U34165 (N_34165,N_33893,N_32959);
and U34166 (N_34166,N_32878,N_32016);
or U34167 (N_34167,N_32707,N_33932);
or U34168 (N_34168,N_32046,N_32241);
xnor U34169 (N_34169,N_32007,N_32439);
xor U34170 (N_34170,N_33445,N_32682);
nor U34171 (N_34171,N_33451,N_32043);
or U34172 (N_34172,N_32558,N_33363);
xnor U34173 (N_34173,N_32759,N_32047);
nand U34174 (N_34174,N_33170,N_32287);
xor U34175 (N_34175,N_33443,N_32089);
and U34176 (N_34176,N_33202,N_33281);
and U34177 (N_34177,N_32248,N_33515);
nand U34178 (N_34178,N_32071,N_32853);
or U34179 (N_34179,N_32833,N_33980);
and U34180 (N_34180,N_33659,N_32330);
nand U34181 (N_34181,N_32551,N_32975);
and U34182 (N_34182,N_32736,N_33842);
and U34183 (N_34183,N_32603,N_33057);
xnor U34184 (N_34184,N_33482,N_32356);
xor U34185 (N_34185,N_32252,N_32048);
and U34186 (N_34186,N_33179,N_32098);
xor U34187 (N_34187,N_33442,N_33242);
nand U34188 (N_34188,N_32327,N_33197);
nand U34189 (N_34189,N_32730,N_32178);
or U34190 (N_34190,N_32549,N_32488);
nand U34191 (N_34191,N_32668,N_33338);
and U34192 (N_34192,N_33872,N_33230);
nand U34193 (N_34193,N_33246,N_32020);
or U34194 (N_34194,N_33999,N_32548);
nor U34195 (N_34195,N_33078,N_33107);
nor U34196 (N_34196,N_33807,N_33615);
and U34197 (N_34197,N_32914,N_32181);
and U34198 (N_34198,N_32430,N_33719);
nand U34199 (N_34199,N_33636,N_32956);
or U34200 (N_34200,N_33641,N_32505);
and U34201 (N_34201,N_32398,N_32370);
nor U34202 (N_34202,N_32921,N_33925);
or U34203 (N_34203,N_33385,N_33159);
nand U34204 (N_34204,N_33914,N_32758);
and U34205 (N_34205,N_33063,N_33508);
nor U34206 (N_34206,N_33098,N_32375);
and U34207 (N_34207,N_32836,N_33942);
xnor U34208 (N_34208,N_32530,N_32651);
nand U34209 (N_34209,N_32522,N_33681);
nor U34210 (N_34210,N_32386,N_33846);
nor U34211 (N_34211,N_33810,N_32443);
nand U34212 (N_34212,N_32536,N_33699);
xnor U34213 (N_34213,N_33913,N_32323);
and U34214 (N_34214,N_32774,N_33927);
nor U34215 (N_34215,N_33376,N_33494);
xnor U34216 (N_34216,N_33265,N_32605);
xor U34217 (N_34217,N_32761,N_33571);
nand U34218 (N_34218,N_33972,N_32096);
and U34219 (N_34219,N_33540,N_32496);
nand U34220 (N_34220,N_32260,N_32186);
and U34221 (N_34221,N_32438,N_33049);
or U34222 (N_34222,N_32208,N_32141);
and U34223 (N_34223,N_32372,N_33044);
xnor U34224 (N_34224,N_32419,N_33369);
and U34225 (N_34225,N_33952,N_32905);
nand U34226 (N_34226,N_33347,N_32408);
nor U34227 (N_34227,N_32539,N_32069);
nand U34228 (N_34228,N_33638,N_33759);
and U34229 (N_34229,N_32404,N_33468);
xor U34230 (N_34230,N_33566,N_32989);
nand U34231 (N_34231,N_33510,N_32197);
xnor U34232 (N_34232,N_33319,N_32951);
xnor U34233 (N_34233,N_33815,N_33151);
and U34234 (N_34234,N_32571,N_33639);
xor U34235 (N_34235,N_33498,N_32660);
nand U34236 (N_34236,N_33216,N_33024);
or U34237 (N_34237,N_32161,N_32498);
or U34238 (N_34238,N_33030,N_32223);
nor U34239 (N_34239,N_33322,N_33409);
or U34240 (N_34240,N_33597,N_32869);
nor U34241 (N_34241,N_33858,N_32669);
or U34242 (N_34242,N_32795,N_33467);
nand U34243 (N_34243,N_32763,N_32678);
xor U34244 (N_34244,N_33522,N_32247);
nor U34245 (N_34245,N_33138,N_33110);
or U34246 (N_34246,N_33642,N_32679);
nand U34247 (N_34247,N_32715,N_32029);
and U34248 (N_34248,N_33260,N_32646);
and U34249 (N_34249,N_32392,N_33558);
or U34250 (N_34250,N_33088,N_32003);
nor U34251 (N_34251,N_33313,N_32004);
nand U34252 (N_34252,N_32094,N_32648);
and U34253 (N_34253,N_32279,N_32865);
xor U34254 (N_34254,N_33015,N_32923);
and U34255 (N_34255,N_32901,N_32328);
nor U34256 (N_34256,N_33561,N_32767);
xnor U34257 (N_34257,N_32431,N_32021);
nand U34258 (N_34258,N_32359,N_32305);
nor U34259 (N_34259,N_33249,N_33367);
nand U34260 (N_34260,N_33727,N_32531);
and U34261 (N_34261,N_33783,N_32753);
nand U34262 (N_34262,N_32150,N_32729);
or U34263 (N_34263,N_32129,N_33043);
nand U34264 (N_34264,N_33484,N_33791);
xor U34265 (N_34265,N_32057,N_33757);
and U34266 (N_34266,N_32240,N_33393);
xor U34267 (N_34267,N_32407,N_32124);
or U34268 (N_34268,N_32670,N_33630);
and U34269 (N_34269,N_33381,N_33332);
nor U34270 (N_34270,N_33140,N_32426);
nor U34271 (N_34271,N_32993,N_33519);
nand U34272 (N_34272,N_32820,N_33272);
or U34273 (N_34273,N_32030,N_32850);
or U34274 (N_34274,N_32180,N_32418);
and U34275 (N_34275,N_32598,N_33579);
nor U34276 (N_34276,N_33698,N_33818);
nor U34277 (N_34277,N_33448,N_32737);
xor U34278 (N_34278,N_33418,N_32387);
and U34279 (N_34279,N_32266,N_33663);
xor U34280 (N_34280,N_32664,N_32106);
nor U34281 (N_34281,N_32784,N_33245);
xor U34282 (N_34282,N_32579,N_33608);
nand U34283 (N_34283,N_33779,N_33436);
and U34284 (N_34284,N_33812,N_33239);
xnor U34285 (N_34285,N_32928,N_33543);
nand U34286 (N_34286,N_33499,N_32478);
xnor U34287 (N_34287,N_33291,N_33432);
xor U34288 (N_34288,N_32834,N_33462);
nand U34289 (N_34289,N_32705,N_33068);
xor U34290 (N_34290,N_33237,N_32475);
nor U34291 (N_34291,N_32904,N_33891);
or U34292 (N_34292,N_32347,N_33169);
or U34293 (N_34293,N_33673,N_33092);
nor U34294 (N_34294,N_32801,N_32576);
nand U34295 (N_34295,N_32967,N_32309);
or U34296 (N_34296,N_32000,N_32875);
and U34297 (N_34297,N_33071,N_32065);
nor U34298 (N_34298,N_32044,N_33814);
or U34299 (N_34299,N_33785,N_33266);
xor U34300 (N_34300,N_33723,N_32412);
nor U34301 (N_34301,N_32088,N_32385);
nor U34302 (N_34302,N_33528,N_32823);
and U34303 (N_34303,N_32066,N_33847);
nand U34304 (N_34304,N_33658,N_32099);
xnor U34305 (N_34305,N_32586,N_32776);
or U34306 (N_34306,N_32388,N_32563);
and U34307 (N_34307,N_33387,N_33075);
or U34308 (N_34308,N_33069,N_32570);
or U34309 (N_34309,N_32194,N_33006);
or U34310 (N_34310,N_33275,N_32585);
and U34311 (N_34311,N_33166,N_33813);
or U34312 (N_34312,N_33603,N_32319);
nand U34313 (N_34313,N_32243,N_33258);
or U34314 (N_34314,N_32081,N_32156);
nand U34315 (N_34315,N_33321,N_33557);
nor U34316 (N_34316,N_32143,N_32685);
or U34317 (N_34317,N_33072,N_32898);
or U34318 (N_34318,N_33465,N_32887);
nor U34319 (N_34319,N_32543,N_33225);
and U34320 (N_34320,N_33580,N_32032);
nor U34321 (N_34321,N_33886,N_33027);
nor U34322 (N_34322,N_33470,N_33559);
and U34323 (N_34323,N_32120,N_33521);
nand U34324 (N_34324,N_32821,N_33235);
nor U34325 (N_34325,N_33257,N_32103);
xor U34326 (N_34326,N_32814,N_32383);
or U34327 (N_34327,N_32659,N_33241);
nor U34328 (N_34328,N_33809,N_33029);
or U34329 (N_34329,N_32117,N_32031);
or U34330 (N_34330,N_32135,N_32234);
and U34331 (N_34331,N_33729,N_32207);
and U34332 (N_34332,N_33011,N_33836);
xnor U34333 (N_34333,N_33908,N_32770);
nor U34334 (N_34334,N_32826,N_33181);
nand U34335 (N_34335,N_33750,N_33161);
and U34336 (N_34336,N_33781,N_33084);
nand U34337 (N_34337,N_33086,N_32634);
or U34338 (N_34338,N_33300,N_33137);
xor U34339 (N_34339,N_32074,N_33226);
and U34340 (N_34340,N_32907,N_33602);
nor U34341 (N_34341,N_33419,N_32930);
nand U34342 (N_34342,N_32996,N_33977);
or U34343 (N_34343,N_32501,N_32518);
nand U34344 (N_34344,N_32973,N_33128);
nor U34345 (N_34345,N_32509,N_33704);
nand U34346 (N_34346,N_32593,N_32783);
nand U34347 (N_34347,N_32789,N_33590);
and U34348 (N_34348,N_32093,N_32049);
nor U34349 (N_34349,N_32100,N_32920);
or U34350 (N_34350,N_32533,N_33545);
xnor U34351 (N_34351,N_33328,N_33851);
xnor U34352 (N_34352,N_32136,N_33377);
and U34353 (N_34353,N_33175,N_33447);
nand U34354 (N_34354,N_32998,N_33268);
nand U34355 (N_34355,N_33696,N_33973);
nor U34356 (N_34356,N_32852,N_32752);
nand U34357 (N_34357,N_33045,N_32631);
nor U34358 (N_34358,N_33173,N_32201);
and U34359 (N_34359,N_32744,N_33854);
xnor U34360 (N_34360,N_33676,N_33007);
nor U34361 (N_34361,N_33085,N_33870);
xnor U34362 (N_34362,N_32787,N_33286);
nand U34363 (N_34363,N_33634,N_33737);
nor U34364 (N_34364,N_33806,N_33605);
or U34365 (N_34365,N_32345,N_32613);
nor U34366 (N_34366,N_33770,N_33936);
nor U34367 (N_34367,N_32653,N_33229);
and U34368 (N_34368,N_32882,N_32466);
or U34369 (N_34369,N_32297,N_33968);
or U34370 (N_34370,N_32493,N_33415);
xor U34371 (N_34371,N_32472,N_33201);
or U34372 (N_34372,N_33706,N_32308);
xnor U34373 (N_34373,N_32282,N_32945);
or U34374 (N_34374,N_33581,N_32591);
nor U34375 (N_34375,N_32231,N_33929);
nor U34376 (N_34376,N_32006,N_32512);
and U34377 (N_34377,N_33444,N_32290);
and U34378 (N_34378,N_32402,N_32390);
xnor U34379 (N_34379,N_32125,N_33456);
nor U34380 (N_34380,N_32780,N_33192);
nand U34381 (N_34381,N_33323,N_32013);
xor U34382 (N_34382,N_32857,N_32002);
or U34383 (N_34383,N_32056,N_32355);
nor U34384 (N_34384,N_33906,N_32841);
xnor U34385 (N_34385,N_33838,N_33171);
nor U34386 (N_34386,N_33953,N_32663);
or U34387 (N_34387,N_33217,N_32394);
nand U34388 (N_34388,N_32073,N_32957);
nor U34389 (N_34389,N_32894,N_33255);
nand U34390 (N_34390,N_33831,N_32175);
and U34391 (N_34391,N_33577,N_33576);
nor U34392 (N_34392,N_32818,N_33959);
xnor U34393 (N_34393,N_33868,N_32822);
or U34394 (N_34394,N_32863,N_33544);
or U34395 (N_34395,N_33637,N_32939);
and U34396 (N_34396,N_32130,N_32525);
nor U34397 (N_34397,N_32845,N_32023);
nand U34398 (N_34398,N_33089,N_33589);
xnor U34399 (N_34399,N_32229,N_32778);
nand U34400 (N_34400,N_32269,N_32219);
or U34401 (N_34401,N_32908,N_33271);
nor U34402 (N_34402,N_32872,N_33766);
nor U34403 (N_34403,N_32424,N_32846);
or U34404 (N_34404,N_33310,N_32362);
nand U34405 (N_34405,N_33172,N_33274);
or U34406 (N_34406,N_32888,N_33126);
nor U34407 (N_34407,N_32675,N_32160);
or U34408 (N_34408,N_33010,N_32464);
and U34409 (N_34409,N_32541,N_32743);
nor U34410 (N_34410,N_32521,N_33537);
and U34411 (N_34411,N_33595,N_33650);
nor U34412 (N_34412,N_33394,N_33714);
nand U34413 (N_34413,N_32699,N_33911);
xor U34414 (N_34414,N_33938,N_32444);
xnor U34415 (N_34415,N_33517,N_33435);
nor U34416 (N_34416,N_33550,N_33103);
or U34417 (N_34417,N_33541,N_33342);
nor U34418 (N_34418,N_32727,N_33017);
nand U34419 (N_34419,N_32734,N_32250);
nor U34420 (N_34420,N_32338,N_33306);
nor U34421 (N_34421,N_32352,N_33187);
nand U34422 (N_34422,N_32022,N_33304);
and U34423 (N_34423,N_32971,N_33879);
nand U34424 (N_34424,N_33374,N_33335);
xnor U34425 (N_34425,N_32445,N_32185);
nand U34426 (N_34426,N_33941,N_32236);
nor U34427 (N_34427,N_32709,N_33299);
or U34428 (N_34428,N_32680,N_33679);
nand U34429 (N_34429,N_33573,N_33250);
or U34430 (N_34430,N_32747,N_33380);
xor U34431 (N_34431,N_33124,N_33967);
nor U34432 (N_34432,N_33388,N_33853);
nor U34433 (N_34433,N_32283,N_32339);
and U34434 (N_34434,N_32511,N_33730);
xor U34435 (N_34435,N_32348,N_33777);
nor U34436 (N_34436,N_32379,N_33486);
or U34437 (N_34437,N_32855,N_32552);
xor U34438 (N_34438,N_33690,N_33118);
or U34439 (N_34439,N_32991,N_32647);
nor U34440 (N_34440,N_33816,N_33090);
nor U34441 (N_34441,N_33000,N_32367);
xor U34442 (N_34442,N_32245,N_32745);
xor U34443 (N_34443,N_32588,N_33096);
nand U34444 (N_34444,N_32147,N_32654);
or U34445 (N_34445,N_32410,N_33280);
or U34446 (N_34446,N_32369,N_33697);
xor U34447 (N_34447,N_33440,N_33871);
and U34448 (N_34448,N_33599,N_33620);
xor U34449 (N_34449,N_33661,N_33951);
nand U34450 (N_34450,N_33428,N_32427);
nor U34451 (N_34451,N_33117,N_33660);
nor U34452 (N_34452,N_32055,N_32008);
or U34453 (N_34453,N_33143,N_32909);
xor U34454 (N_34454,N_33691,N_33424);
or U34455 (N_34455,N_33469,N_32874);
or U34456 (N_34456,N_33962,N_33797);
nand U34457 (N_34457,N_33950,N_32118);
nand U34458 (N_34458,N_33700,N_32681);
nor U34459 (N_34459,N_32917,N_33316);
or U34460 (N_34460,N_33193,N_33829);
xnor U34461 (N_34461,N_33366,N_32566);
nand U34462 (N_34462,N_33329,N_33664);
nor U34463 (N_34463,N_32320,N_32698);
nand U34464 (N_34464,N_33361,N_32982);
or U34465 (N_34465,N_32481,N_33823);
xor U34466 (N_34466,N_33917,N_32458);
xor U34467 (N_34467,N_33233,N_32779);
nor U34468 (N_34468,N_33989,N_33901);
nor U34469 (N_34469,N_33182,N_33132);
nor U34470 (N_34470,N_33694,N_33326);
xnor U34471 (N_34471,N_33053,N_33523);
nand U34472 (N_34472,N_33725,N_32301);
nand U34473 (N_34473,N_33452,N_32457);
nand U34474 (N_34474,N_33668,N_33665);
nand U34475 (N_34475,N_33232,N_33839);
and U34476 (N_34476,N_32910,N_33212);
nor U34477 (N_34477,N_32963,N_33036);
and U34478 (N_34478,N_33218,N_33568);
nand U34479 (N_34479,N_33805,N_33227);
nor U34480 (N_34480,N_32819,N_32629);
or U34481 (N_34481,N_32798,N_33860);
nand U34482 (N_34482,N_33431,N_32915);
or U34483 (N_34483,N_33352,N_32622);
or U34484 (N_34484,N_33509,N_32714);
or U34485 (N_34485,N_33682,N_33627);
xor U34486 (N_34486,N_32880,N_33052);
xnor U34487 (N_34487,N_32830,N_33083);
or U34488 (N_34488,N_33726,N_32934);
or U34489 (N_34489,N_32351,N_32422);
nand U34490 (N_34490,N_32153,N_33285);
nor U34491 (N_34491,N_33881,N_33582);
or U34492 (N_34492,N_33046,N_32092);
or U34493 (N_34493,N_32343,N_32546);
xnor U34494 (N_34494,N_32451,N_33863);
nand U34495 (N_34495,N_32732,N_32039);
or U34496 (N_34496,N_33614,N_33038);
nand U34497 (N_34497,N_32064,N_33327);
and U34498 (N_34498,N_33120,N_33607);
nand U34499 (N_34499,N_32617,N_33715);
xor U34500 (N_34500,N_32691,N_32405);
xor U34501 (N_34501,N_33433,N_32371);
nand U34502 (N_34502,N_33028,N_33667);
nor U34503 (N_34503,N_33213,N_32726);
nor U34504 (N_34504,N_33943,N_33312);
or U34505 (N_34505,N_33370,N_32257);
xnor U34506 (N_34506,N_32879,N_32697);
or U34507 (N_34507,N_33758,N_32105);
xor U34508 (N_34508,N_33874,N_33427);
and U34509 (N_34509,N_32999,N_32026);
nor U34510 (N_34510,N_33251,N_33111);
or U34511 (N_34511,N_33693,N_32067);
and U34512 (N_34512,N_33984,N_33990);
xnor U34513 (N_34513,N_33214,N_32864);
or U34514 (N_34514,N_33530,N_32858);
xnor U34515 (N_34515,N_32416,N_33905);
and U34516 (N_34516,N_33578,N_33099);
nor U34517 (N_34517,N_33480,N_32532);
xnor U34518 (N_34518,N_33976,N_33014);
and U34519 (N_34519,N_33458,N_33895);
xnor U34520 (N_34520,N_33353,N_33533);
and U34521 (N_34521,N_32365,N_33056);
or U34522 (N_34522,N_32912,N_33156);
and U34523 (N_34523,N_33411,N_32376);
nand U34524 (N_34524,N_32122,N_32950);
and U34525 (N_34525,N_32246,N_32101);
nor U34526 (N_34526,N_32935,N_33267);
nor U34527 (N_34527,N_32173,N_33303);
xnor U34528 (N_34528,N_33031,N_33624);
and U34529 (N_34529,N_32137,N_32508);
xnor U34530 (N_34530,N_32594,N_33922);
or U34531 (N_34531,N_33918,N_32713);
or U34532 (N_34532,N_33189,N_33767);
nand U34533 (N_34533,N_32080,N_33209);
nand U34534 (N_34534,N_33645,N_32307);
and U34535 (N_34535,N_33464,N_33611);
and U34536 (N_34536,N_32277,N_32862);
nand U34537 (N_34537,N_33164,N_33104);
xor U34538 (N_34538,N_32952,N_32158);
xor U34539 (N_34539,N_32133,N_33142);
nor U34540 (N_34540,N_32677,N_33123);
and U34541 (N_34541,N_33749,N_32696);
nor U34542 (N_34542,N_33994,N_33294);
and U34543 (N_34543,N_33548,N_32467);
xnor U34544 (N_34544,N_32817,N_32138);
or U34545 (N_34545,N_33359,N_32502);
xor U34546 (N_34546,N_33188,N_32295);
nor U34547 (N_34547,N_32183,N_32760);
nor U34548 (N_34548,N_33333,N_33183);
nand U34549 (N_34549,N_32433,N_32868);
xor U34550 (N_34550,N_32010,N_32123);
and U34551 (N_34551,N_32220,N_32876);
xnor U34552 (N_34552,N_33325,N_32871);
and U34553 (N_34553,N_32861,N_33288);
nand U34554 (N_34554,N_33506,N_32940);
xnor U34555 (N_34555,N_33574,N_32673);
or U34556 (N_34556,N_33830,N_32251);
and U34557 (N_34557,N_32883,N_33125);
or U34558 (N_34558,N_33856,N_32192);
xor U34559 (N_34559,N_33012,N_33974);
and U34560 (N_34560,N_33389,N_32626);
nor U34561 (N_34561,N_32547,N_32473);
xnor U34562 (N_34562,N_33833,N_33406);
and U34563 (N_34563,N_33449,N_32149);
xnor U34564 (N_34564,N_32718,N_33339);
nor U34565 (N_34565,N_32557,N_32641);
nand U34566 (N_34566,N_32655,N_32350);
and U34567 (N_34567,N_32720,N_32773);
nor U34568 (N_34568,N_32741,N_33158);
xor U34569 (N_34569,N_32656,N_33562);
nand U34570 (N_34570,N_32476,N_33778);
and U34571 (N_34571,N_32060,N_33277);
nor U34572 (N_34572,N_32014,N_33640);
and U34573 (N_34573,N_32400,N_33077);
or U34574 (N_34574,N_33008,N_33722);
or U34575 (N_34575,N_32838,N_32196);
nor U34576 (N_34576,N_32128,N_32382);
nand U34577 (N_34577,N_33144,N_32163);
xor U34578 (N_34578,N_32377,N_32520);
and U34579 (N_34579,N_32528,N_32097);
or U34580 (N_34580,N_32253,N_33513);
or U34581 (N_34581,N_33703,N_33567);
xor U34582 (N_34582,N_32980,N_33738);
nand U34583 (N_34583,N_32911,N_33026);
and U34584 (N_34584,N_33903,N_33792);
or U34585 (N_34585,N_33391,N_33334);
nand U34586 (N_34586,N_32357,N_32373);
and U34587 (N_34587,N_33207,N_33855);
or U34588 (N_34588,N_32281,N_33492);
xor U34589 (N_34589,N_33109,N_32280);
nor U34590 (N_34590,N_33236,N_32294);
or U34591 (N_34591,N_32722,N_33983);
or U34592 (N_34592,N_32095,N_32748);
xor U34593 (N_34593,N_32401,N_33852);
nand U34594 (N_34594,N_33094,N_32643);
or U34595 (N_34595,N_32471,N_33059);
nand U34596 (N_34596,N_32110,N_32058);
nand U34597 (N_34597,N_33350,N_33150);
or U34598 (N_34598,N_33390,N_32633);
nand U34599 (N_34599,N_33375,N_33307);
nor U34600 (N_34600,N_33720,N_32762);
nand U34601 (N_34601,N_32754,N_32480);
xnor U34602 (N_34602,N_33995,N_33512);
and U34603 (N_34603,N_32529,N_32671);
xor U34604 (N_34604,N_32932,N_33939);
or U34605 (N_34605,N_33289,N_33283);
or U34606 (N_34606,N_32944,N_32454);
xor U34607 (N_34607,N_32494,N_33996);
nor U34608 (N_34608,N_32409,N_32463);
xor U34609 (N_34609,N_33820,N_33819);
or U34610 (N_34610,N_33554,N_32565);
xnor U34611 (N_34611,N_32797,N_33701);
and U34612 (N_34612,N_33817,N_32906);
and U34613 (N_34613,N_33849,N_33354);
xor U34614 (N_34614,N_32574,N_32119);
nor U34615 (N_34615,N_32990,N_32068);
and U34616 (N_34616,N_32925,N_33539);
or U34617 (N_34617,N_32146,N_32075);
nand U34618 (N_34618,N_32334,N_33446);
and U34619 (N_34619,N_32288,N_33500);
nand U34620 (N_34620,N_32337,N_32009);
and U34621 (N_34621,N_33177,N_33670);
and U34622 (N_34622,N_33475,N_33034);
nand U34623 (N_34623,N_33930,N_32640);
or U34624 (N_34624,N_33018,N_33402);
nor U34625 (N_34625,N_33859,N_33211);
nor U34626 (N_34626,N_33064,N_32151);
nor U34627 (N_34627,N_32017,N_33009);
nor U34628 (N_34628,N_32061,N_32179);
or U34629 (N_34629,N_32955,N_33617);
nor U34630 (N_34630,N_33958,N_33643);
nand U34631 (N_34631,N_33845,N_33050);
nand U34632 (N_34632,N_33349,N_32803);
nor U34633 (N_34633,N_33371,N_32154);
nor U34634 (N_34634,N_32903,N_33351);
nand U34635 (N_34635,N_33728,N_32423);
nor U34636 (N_34636,N_32168,N_32856);
nand U34637 (N_34637,N_33790,N_33493);
nor U34638 (N_34638,N_32983,N_32134);
nor U34639 (N_34639,N_32011,N_33956);
or U34640 (N_34640,N_32564,N_33601);
and U34641 (N_34641,N_33784,N_32112);
xor U34642 (N_34642,N_32933,N_33985);
and U34643 (N_34643,N_32470,N_33360);
xor U34644 (N_34644,N_32140,N_32115);
and U34645 (N_34645,N_32742,N_33080);
nor U34646 (N_34646,N_32620,N_32916);
nand U34647 (N_34647,N_32264,N_33631);
and U34648 (N_34648,N_32802,N_33051);
nand U34649 (N_34649,N_32517,N_32378);
and U34650 (N_34650,N_33685,N_33931);
and U34651 (N_34651,N_33709,N_32485);
or U34652 (N_34652,N_32015,N_33732);
or U34653 (N_34653,N_33254,N_32828);
xor U34654 (N_34654,N_33635,N_33717);
nand U34655 (N_34655,N_32082,N_33724);
and U34656 (N_34656,N_33115,N_33247);
nand U34657 (N_34657,N_33773,N_33745);
nor U34658 (N_34658,N_33954,N_32315);
nand U34659 (N_34659,N_32764,N_33221);
or U34660 (N_34660,N_33460,N_33534);
nor U34661 (N_34661,N_32019,N_32972);
nand U34662 (N_34662,N_32805,N_32276);
nor U34663 (N_34663,N_32946,N_33297);
or U34664 (N_34664,N_33344,N_33525);
xnor U34665 (N_34665,N_32321,N_32213);
and U34666 (N_34666,N_33383,N_33843);
or U34667 (N_34667,N_33542,N_32610);
nor U34668 (N_34668,N_33882,N_33203);
and U34669 (N_34669,N_32102,N_33801);
nor U34670 (N_34670,N_33248,N_33768);
xor U34671 (N_34671,N_33865,N_32195);
or U34672 (N_34672,N_33923,N_33588);
nand U34673 (N_34673,N_33160,N_32233);
and U34674 (N_34674,N_32970,N_33902);
or U34675 (N_34675,N_32018,N_32960);
xnor U34676 (N_34676,N_32070,N_33178);
nor U34677 (N_34677,N_32038,N_32639);
and U34678 (N_34678,N_33483,N_33924);
and U34679 (N_34679,N_32630,N_33416);
nand U34680 (N_34680,N_33892,N_33896);
nand U34681 (N_34681,N_33998,N_32666);
xor U34682 (N_34682,N_33644,N_32267);
or U34683 (N_34683,N_32182,N_33284);
and U34684 (N_34684,N_33675,N_32176);
or U34685 (N_34685,N_33206,N_32396);
and U34686 (N_34686,N_33586,N_32028);
nor U34687 (N_34687,N_32085,N_33407);
or U34688 (N_34688,N_32694,N_32205);
nand U34689 (N_34689,N_33324,N_32062);
nand U34690 (N_34690,N_33314,N_32311);
or U34691 (N_34691,N_33244,N_32936);
nor U34692 (N_34692,N_32455,N_32414);
nand U34693 (N_34693,N_32114,N_32575);
nand U34694 (N_34694,N_32926,N_32599);
or U34695 (N_34695,N_33223,N_33802);
nor U34696 (N_34696,N_32540,N_33628);
nor U34697 (N_34697,N_32775,N_32602);
nand U34698 (N_34698,N_33372,N_32261);
xor U34699 (N_34699,N_32435,N_33234);
nor U34700 (N_34700,N_33136,N_32860);
nand U34701 (N_34701,N_33712,N_32628);
and U34702 (N_34702,N_32036,N_32609);
or U34703 (N_34703,N_32224,N_32635);
nor U34704 (N_34704,N_32051,N_33453);
nor U34705 (N_34705,N_33563,N_33346);
or U34706 (N_34706,N_33466,N_33864);
xnor U34707 (N_34707,N_32483,N_32202);
xor U34708 (N_34708,N_32587,N_32623);
nand U34709 (N_34709,N_32800,N_32399);
or U34710 (N_34710,N_33002,N_33219);
nor U34711 (N_34711,N_32479,N_32867);
nand U34712 (N_34712,N_32187,N_32113);
nand U34713 (N_34713,N_33195,N_32446);
xor U34714 (N_34714,N_33772,N_32658);
or U34715 (N_34715,N_32450,N_32790);
and U34716 (N_34716,N_33004,N_32121);
xnor U34717 (N_34717,N_32127,N_32735);
and U34718 (N_34718,N_33205,N_33302);
nor U34719 (N_34719,N_33935,N_32535);
or U34720 (N_34720,N_32740,N_33549);
xnor U34721 (N_34721,N_32791,N_32034);
or U34722 (N_34722,N_33200,N_33695);
or U34723 (N_34723,N_33672,N_33067);
xor U34724 (N_34724,N_32341,N_32033);
xnor U34725 (N_34725,N_33616,N_32242);
and U34726 (N_34726,N_33259,N_33129);
nand U34727 (N_34727,N_33122,N_32986);
nand U34728 (N_34728,N_33992,N_33887);
nor U34729 (N_34729,N_32637,N_33721);
xor U34730 (N_34730,N_32461,N_32389);
and U34731 (N_34731,N_33112,N_33337);
and U34732 (N_34732,N_32896,N_33224);
xor U34733 (N_34733,N_33666,N_32214);
or U34734 (N_34734,N_33897,N_33422);
or U34735 (N_34735,N_33880,N_32724);
nor U34736 (N_34736,N_32270,N_33878);
or U34737 (N_34737,N_33505,N_32842);
and U34738 (N_34738,N_33916,N_33261);
and U34739 (N_34739,N_33410,N_32354);
or U34740 (N_34740,N_32237,N_33735);
nor U34741 (N_34741,N_32198,N_32221);
or U34742 (N_34742,N_33646,N_32142);
nor U34743 (N_34743,N_33742,N_32995);
nand U34744 (N_34744,N_33252,N_33292);
or U34745 (N_34745,N_33587,N_33504);
nor U34746 (N_34746,N_32676,N_32453);
and U34747 (N_34747,N_33290,N_33293);
nor U34748 (N_34748,N_32642,N_32592);
and U34749 (N_34749,N_32554,N_32804);
and U34750 (N_34750,N_33744,N_32001);
xnor U34751 (N_34751,N_32436,N_33538);
xor U34752 (N_34752,N_33503,N_32193);
or U34753 (N_34753,N_33988,N_33421);
nand U34754 (N_34754,N_32053,N_32304);
or U34755 (N_34755,N_32650,N_32661);
and U34756 (N_34756,N_32063,N_32589);
or U34757 (N_34757,N_33222,N_32924);
or U34758 (N_34758,N_33495,N_33379);
xor U34759 (N_34759,N_32393,N_32079);
and U34760 (N_34760,N_32216,N_33754);
or U34761 (N_34761,N_32289,N_32590);
xor U34762 (N_34762,N_33135,N_32268);
nor U34763 (N_34763,N_33476,N_33583);
and U34764 (N_34764,N_33687,N_32434);
nand U34765 (N_34765,N_32303,N_32162);
xor U34766 (N_34766,N_32503,N_33689);
nor U34767 (N_34767,N_32825,N_33477);
nand U34768 (N_34768,N_33796,N_32832);
nor U34769 (N_34769,N_32578,N_33618);
or U34770 (N_34770,N_33457,N_33091);
nor U34771 (N_34771,N_32190,N_33473);
nor U34772 (N_34772,N_32793,N_33488);
or U34773 (N_34773,N_32417,N_32325);
nand U34774 (N_34774,N_32792,N_32516);
and U34775 (N_34775,N_33108,N_32200);
and U34776 (N_34776,N_33705,N_33279);
and U34777 (N_34777,N_33960,N_33426);
xnor U34778 (N_34778,N_33355,N_33861);
nand U34779 (N_34779,N_33592,N_32567);
and U34780 (N_34780,N_33194,N_33560);
nand U34781 (N_34781,N_32090,N_32428);
nor U34782 (N_34782,N_32988,N_33130);
nor U34783 (N_34783,N_33441,N_32299);
xnor U34784 (N_34784,N_33827,N_32227);
xnor U34785 (N_34785,N_32701,N_33828);
xnor U34786 (N_34786,N_32152,N_33263);
and U34787 (N_34787,N_32167,N_32087);
nor U34788 (N_34788,N_32164,N_32238);
and U34789 (N_34789,N_32954,N_33947);
and U34790 (N_34790,N_33093,N_32462);
nor U34791 (N_34791,N_33671,N_33546);
nor U34792 (N_34792,N_33662,N_32189);
nand U34793 (N_34793,N_33397,N_33417);
nor U34794 (N_34794,N_32477,N_32979);
nand U34795 (N_34795,N_32829,N_32606);
nand U34796 (N_34796,N_32997,N_32716);
nor U34797 (N_34797,N_32313,N_32459);
nand U34798 (N_34798,N_33647,N_33536);
and U34799 (N_34799,N_33481,N_33926);
xnor U34800 (N_34800,N_33764,N_32968);
nand U34801 (N_34801,N_33163,N_32465);
or U34802 (N_34802,N_33760,N_32366);
nor U34803 (N_34803,N_33401,N_32527);
nor U34804 (N_34804,N_33343,N_32644);
and U34805 (N_34805,N_33591,N_33039);
and U34806 (N_34806,N_33516,N_32232);
and U34807 (N_34807,N_32550,N_32292);
or U34808 (N_34808,N_33622,N_33553);
nor U34809 (N_34809,N_32209,N_33395);
and U34810 (N_34810,N_32688,N_32116);
or U34811 (N_34811,N_33800,N_33844);
and U34812 (N_34812,N_33775,N_32542);
nor U34813 (N_34813,N_32786,N_33755);
nor U34814 (N_34814,N_32515,N_32931);
or U34815 (N_34815,N_33490,N_33514);
or U34816 (N_34816,N_32568,N_33743);
and U34817 (N_34817,N_32203,N_33055);
nor U34818 (N_34818,N_32859,N_32230);
and U34819 (N_34819,N_33688,N_33520);
xor U34820 (N_34820,N_32706,N_33060);
or U34821 (N_34821,N_33184,N_33295);
nor U34822 (N_34822,N_32035,N_33474);
nand U34823 (N_34823,N_33439,N_33032);
and U34824 (N_34824,N_32148,N_33524);
and U34825 (N_34825,N_33382,N_33535);
or U34826 (N_34826,N_33780,N_32374);
nand U34827 (N_34827,N_32886,N_33966);
xnor U34828 (N_34828,N_32665,N_33119);
and U34829 (N_34829,N_32739,N_33531);
and U34830 (N_34830,N_32211,N_33070);
and U34831 (N_34831,N_32155,N_32636);
and U34832 (N_34832,N_33336,N_33786);
nand U34833 (N_34833,N_32440,N_33153);
nor U34834 (N_34834,N_33569,N_33609);
xor U34835 (N_34835,N_33095,N_32851);
or U34836 (N_34836,N_33575,N_32108);
nand U34837 (N_34837,N_33133,N_33358);
nor U34838 (N_34838,N_33788,N_32166);
or U34839 (N_34839,N_33653,N_33900);
and U34840 (N_34840,N_33016,N_32902);
or U34841 (N_34841,N_32624,N_33157);
nand U34842 (N_34842,N_32873,N_33479);
nor U34843 (N_34843,N_32573,N_33106);
or U34844 (N_34844,N_33121,N_32274);
nand U34845 (N_34845,N_32612,N_32391);
xnor U34846 (N_34846,N_32225,N_33511);
nor U34847 (N_34847,N_32556,N_33154);
xor U34848 (N_34848,N_32555,N_33373);
nor U34849 (N_34849,N_33400,N_33345);
and U34850 (N_34850,N_32913,N_33037);
xor U34851 (N_34851,N_32534,N_33264);
or U34852 (N_34852,N_32621,N_33975);
nor U34853 (N_34853,N_32340,N_32569);
nor U34854 (N_34854,N_32965,N_33405);
xor U34855 (N_34855,N_32259,N_33035);
or U34856 (N_34856,N_32884,N_33471);
or U34857 (N_34857,N_33507,N_33398);
and U34858 (N_34858,N_32723,N_32900);
xnor U34859 (N_34859,N_33731,N_32672);
nor U34860 (N_34860,N_32893,N_32962);
and U34861 (N_34861,N_32746,N_32460);
nand U34862 (N_34862,N_33185,N_32977);
xor U34863 (N_34863,N_32306,N_33487);
xor U34864 (N_34864,N_33654,N_32403);
and U34865 (N_34865,N_32889,N_33594);
nand U34866 (N_34866,N_33403,N_33651);
nor U34867 (N_34867,N_33596,N_33572);
xnor U34868 (N_34868,N_33965,N_33081);
xnor U34869 (N_34869,N_32985,N_33296);
nand U34870 (N_34870,N_32559,N_33748);
nor U34871 (N_34871,N_33686,N_32607);
nor U34872 (N_34872,N_32693,N_32415);
nor U34873 (N_34873,N_33747,N_32052);
or U34874 (N_34874,N_33033,N_32468);
nand U34875 (N_34875,N_32831,N_33834);
and U34876 (N_34876,N_32738,N_33240);
or U34877 (N_34877,N_32625,N_32054);
xor U34878 (N_34878,N_33368,N_33771);
xor U34879 (N_34879,N_32497,N_32562);
xnor U34880 (N_34880,N_33518,N_32692);
nor U34881 (N_34881,N_33884,N_32384);
xnor U34882 (N_34882,N_32275,N_32333);
nand U34883 (N_34883,N_32500,N_32111);
nand U34884 (N_34884,N_32684,N_33621);
xnor U34885 (N_34885,N_33210,N_32139);
and U34886 (N_34886,N_33547,N_32361);
and U34887 (N_34887,N_32881,N_32484);
or U34888 (N_34888,N_33365,N_32597);
xnor U34889 (N_34889,N_32420,N_33710);
and U34890 (N_34890,N_33425,N_33692);
nand U34891 (N_34891,N_32580,N_33961);
nor U34892 (N_34892,N_32604,N_33013);
nand U34893 (N_34893,N_32076,N_32611);
nor U34894 (N_34894,N_32265,N_33485);
or U34895 (N_34895,N_32756,N_33155);
xnor U34896 (N_34896,N_32941,N_32710);
xnor U34897 (N_34897,N_32184,N_33564);
and U34898 (N_34898,N_32492,N_32596);
or U34899 (N_34899,N_32397,N_33082);
nand U34900 (N_34900,N_32107,N_33489);
nor U34901 (N_34901,N_33907,N_33048);
or U34902 (N_34902,N_32218,N_32495);
or U34903 (N_34903,N_32256,N_32835);
and U34904 (N_34904,N_33718,N_32994);
nor U34905 (N_34905,N_33491,N_33404);
xor U34906 (N_34906,N_32584,N_33165);
xnor U34907 (N_34907,N_33957,N_32638);
nand U34908 (N_34908,N_32601,N_32811);
nand U34909 (N_34909,N_32314,N_32144);
and U34910 (N_34910,N_33890,N_32132);
nand U34911 (N_34911,N_32771,N_32796);
or U34912 (N_34912,N_33526,N_33146);
and U34913 (N_34913,N_33386,N_32235);
xor U34914 (N_34914,N_32437,N_33711);
xnor U34915 (N_34915,N_32560,N_33145);
nand U34916 (N_34916,N_33848,N_32474);
nand U34917 (N_34917,N_33899,N_33455);
or U34918 (N_34918,N_32895,N_32005);
nand U34919 (N_34919,N_32077,N_33438);
and U34920 (N_34920,N_32228,N_32429);
nor U34921 (N_34921,N_33837,N_33308);
nand U34922 (N_34922,N_32992,N_33909);
xnor U34923 (N_34923,N_32897,N_33921);
and U34924 (N_34924,N_32411,N_32947);
xnor U34925 (N_34925,N_32572,N_32215);
and U34926 (N_34926,N_33204,N_33963);
nor U34927 (N_34927,N_32848,N_32317);
nor U34928 (N_34928,N_33298,N_32690);
and U34929 (N_34929,N_32649,N_33262);
and U34930 (N_34930,N_33981,N_33191);
nand U34931 (N_34931,N_32948,N_32899);
or U34932 (N_34932,N_33613,N_33256);
or U34933 (N_34933,N_32704,N_33001);
nand U34934 (N_34934,N_33945,N_33463);
nand U34935 (N_34935,N_33869,N_33883);
xnor U34936 (N_34936,N_33808,N_33680);
nor U34937 (N_34937,N_32849,N_33396);
or U34938 (N_34938,N_33131,N_32204);
or U34939 (N_34939,N_32987,N_33005);
or U34940 (N_34940,N_33023,N_32441);
nand U34941 (N_34941,N_32816,N_32104);
xnor U34942 (N_34942,N_33841,N_32131);
nand U34943 (N_34943,N_32024,N_32526);
xor U34944 (N_34944,N_32507,N_33898);
and U34945 (N_34945,N_32808,N_32491);
nand U34946 (N_34946,N_33649,N_33556);
and U34947 (N_34947,N_32072,N_33278);
or U34948 (N_34948,N_32750,N_32652);
nor U34949 (N_34949,N_33061,N_32324);
or U34950 (N_34950,N_33019,N_32091);
and U34951 (N_34951,N_32919,N_33632);
nand U34952 (N_34952,N_32953,N_33066);
nand U34953 (N_34953,N_33040,N_32447);
or U34954 (N_34954,N_32050,N_33593);
xnor U34955 (N_34955,N_32711,N_33761);
or U34956 (N_34956,N_33850,N_32344);
nand U34957 (N_34957,N_33763,N_33904);
or U34958 (N_34958,N_33940,N_33190);
xnor U34959 (N_34959,N_32725,N_33341);
and U34960 (N_34960,N_33025,N_33657);
and U34961 (N_34961,N_32349,N_32877);
nand U34962 (N_34962,N_33101,N_33946);
and U34963 (N_34963,N_32922,N_32291);
nand U34964 (N_34964,N_33765,N_33199);
and U34965 (N_34965,N_33097,N_33392);
nand U34966 (N_34966,N_32974,N_32456);
and U34967 (N_34967,N_32772,N_33610);
nor U34968 (N_34968,N_33141,N_33282);
or U34969 (N_34969,N_32524,N_33600);
nand U34970 (N_34970,N_32777,N_32300);
or U34971 (N_34971,N_32222,N_32302);
xor U34972 (N_34972,N_33147,N_32177);
nand U34973 (N_34973,N_32329,N_33986);
nor U34974 (N_34974,N_32807,N_33894);
or U34975 (N_34975,N_32583,N_33087);
xor U34976 (N_34976,N_33920,N_33633);
nor U34977 (N_34977,N_33648,N_32866);
xor U34978 (N_34978,N_32794,N_33496);
or U34979 (N_34979,N_33309,N_32486);
nand U34980 (N_34980,N_32469,N_32332);
xnor U34981 (N_34981,N_33149,N_32523);
nor U34982 (N_34982,N_33273,N_33461);
xor U34983 (N_34983,N_32538,N_32360);
nand U34984 (N_34984,N_33116,N_33889);
nor U34985 (N_34985,N_33971,N_33982);
or U34986 (N_34986,N_33414,N_33708);
or U34987 (N_34987,N_33527,N_32827);
nand U34988 (N_34988,N_33970,N_33501);
xnor U34989 (N_34989,N_32840,N_33876);
or U34990 (N_34990,N_32854,N_33751);
nand U34991 (N_34991,N_33619,N_32927);
nor U34992 (N_34992,N_32298,N_33795);
nand U34993 (N_34993,N_33062,N_33472);
nor U34994 (N_34994,N_32042,N_32708);
and U34995 (N_34995,N_32217,N_33825);
nand U34996 (N_34996,N_32084,N_32482);
and U34997 (N_34997,N_33674,N_33139);
xnor U34998 (N_34998,N_32632,N_32755);
nand U34999 (N_34999,N_32700,N_33497);
and U35000 (N_35000,N_32238,N_32211);
xor U35001 (N_35001,N_32343,N_32867);
xor U35002 (N_35002,N_33271,N_32452);
nor U35003 (N_35003,N_33070,N_32918);
xnor U35004 (N_35004,N_32952,N_33954);
nor U35005 (N_35005,N_32928,N_32652);
xnor U35006 (N_35006,N_33042,N_33692);
xor U35007 (N_35007,N_33839,N_33005);
nor U35008 (N_35008,N_33800,N_33200);
or U35009 (N_35009,N_32461,N_33119);
and U35010 (N_35010,N_32602,N_32427);
xnor U35011 (N_35011,N_32139,N_33730);
nand U35012 (N_35012,N_32765,N_32079);
xnor U35013 (N_35013,N_33626,N_32980);
xnor U35014 (N_35014,N_33050,N_32837);
nor U35015 (N_35015,N_33823,N_32652);
nor U35016 (N_35016,N_33997,N_33492);
nor U35017 (N_35017,N_33242,N_33257);
nand U35018 (N_35018,N_33850,N_32444);
and U35019 (N_35019,N_32940,N_32867);
and U35020 (N_35020,N_32332,N_33044);
nand U35021 (N_35021,N_32066,N_33222);
or U35022 (N_35022,N_32295,N_33264);
or U35023 (N_35023,N_33810,N_33902);
nor U35024 (N_35024,N_33056,N_33525);
and U35025 (N_35025,N_33279,N_32312);
xor U35026 (N_35026,N_33098,N_33202);
nand U35027 (N_35027,N_32299,N_33071);
xnor U35028 (N_35028,N_32708,N_33029);
or U35029 (N_35029,N_32066,N_33857);
xor U35030 (N_35030,N_32259,N_32837);
or U35031 (N_35031,N_32724,N_32027);
nand U35032 (N_35032,N_32881,N_32233);
nand U35033 (N_35033,N_33912,N_33172);
or U35034 (N_35034,N_32688,N_33930);
or U35035 (N_35035,N_33360,N_32644);
and U35036 (N_35036,N_33796,N_32002);
nand U35037 (N_35037,N_32981,N_32810);
or U35038 (N_35038,N_32774,N_33641);
nor U35039 (N_35039,N_33957,N_33524);
xnor U35040 (N_35040,N_33417,N_33335);
or U35041 (N_35041,N_32317,N_32272);
nor U35042 (N_35042,N_33775,N_33846);
xnor U35043 (N_35043,N_33943,N_32708);
and U35044 (N_35044,N_32276,N_32977);
nor U35045 (N_35045,N_33899,N_33785);
xnor U35046 (N_35046,N_32887,N_32843);
or U35047 (N_35047,N_32852,N_32173);
nor U35048 (N_35048,N_32657,N_33003);
or U35049 (N_35049,N_33792,N_32282);
or U35050 (N_35050,N_32435,N_32689);
or U35051 (N_35051,N_32455,N_32899);
and U35052 (N_35052,N_32138,N_33681);
and U35053 (N_35053,N_32304,N_33194);
nor U35054 (N_35054,N_33887,N_32543);
or U35055 (N_35055,N_33579,N_33687);
or U35056 (N_35056,N_32976,N_32249);
xor U35057 (N_35057,N_32005,N_33645);
nand U35058 (N_35058,N_33965,N_32452);
xnor U35059 (N_35059,N_32578,N_33010);
xor U35060 (N_35060,N_33559,N_32637);
and U35061 (N_35061,N_32385,N_33539);
or U35062 (N_35062,N_33639,N_32767);
and U35063 (N_35063,N_33030,N_32134);
xor U35064 (N_35064,N_33954,N_32885);
or U35065 (N_35065,N_33041,N_32743);
and U35066 (N_35066,N_33161,N_33344);
nand U35067 (N_35067,N_32463,N_33837);
nand U35068 (N_35068,N_32410,N_32727);
xor U35069 (N_35069,N_32389,N_32374);
xor U35070 (N_35070,N_32358,N_33164);
and U35071 (N_35071,N_33521,N_33542);
and U35072 (N_35072,N_32556,N_32692);
or U35073 (N_35073,N_33078,N_32987);
and U35074 (N_35074,N_32163,N_33387);
or U35075 (N_35075,N_33189,N_32611);
nand U35076 (N_35076,N_32569,N_32306);
or U35077 (N_35077,N_33926,N_32476);
nand U35078 (N_35078,N_33831,N_32867);
or U35079 (N_35079,N_33491,N_33605);
or U35080 (N_35080,N_33458,N_32756);
xnor U35081 (N_35081,N_32382,N_32753);
xor U35082 (N_35082,N_33927,N_32705);
or U35083 (N_35083,N_32693,N_32330);
or U35084 (N_35084,N_32119,N_33743);
and U35085 (N_35085,N_33663,N_32900);
nor U35086 (N_35086,N_33287,N_33069);
and U35087 (N_35087,N_32374,N_32131);
xnor U35088 (N_35088,N_32470,N_33088);
and U35089 (N_35089,N_32543,N_33651);
or U35090 (N_35090,N_32862,N_33061);
nor U35091 (N_35091,N_33456,N_32378);
xor U35092 (N_35092,N_33687,N_33532);
nand U35093 (N_35093,N_33373,N_33515);
nor U35094 (N_35094,N_32122,N_33254);
and U35095 (N_35095,N_32303,N_32824);
nand U35096 (N_35096,N_33757,N_33256);
and U35097 (N_35097,N_33872,N_33282);
xor U35098 (N_35098,N_33397,N_32462);
nor U35099 (N_35099,N_33327,N_33432);
nor U35100 (N_35100,N_33803,N_32508);
or U35101 (N_35101,N_32442,N_33041);
and U35102 (N_35102,N_32326,N_33978);
nand U35103 (N_35103,N_32790,N_33941);
nor U35104 (N_35104,N_32336,N_33567);
nand U35105 (N_35105,N_32011,N_33983);
and U35106 (N_35106,N_32336,N_32603);
nor U35107 (N_35107,N_33594,N_33710);
and U35108 (N_35108,N_32918,N_33947);
nor U35109 (N_35109,N_32560,N_33148);
xnor U35110 (N_35110,N_32319,N_33476);
nor U35111 (N_35111,N_32386,N_32421);
nor U35112 (N_35112,N_33609,N_33146);
nand U35113 (N_35113,N_32125,N_33884);
and U35114 (N_35114,N_33121,N_33812);
xor U35115 (N_35115,N_33822,N_33133);
xnor U35116 (N_35116,N_33212,N_33504);
nor U35117 (N_35117,N_32516,N_32863);
nor U35118 (N_35118,N_33853,N_33475);
and U35119 (N_35119,N_33600,N_32688);
xnor U35120 (N_35120,N_33785,N_32486);
xnor U35121 (N_35121,N_33655,N_33351);
or U35122 (N_35122,N_32782,N_32798);
nand U35123 (N_35123,N_32341,N_32158);
nand U35124 (N_35124,N_33484,N_33676);
and U35125 (N_35125,N_32623,N_33764);
nor U35126 (N_35126,N_32574,N_33118);
nand U35127 (N_35127,N_33959,N_33149);
nor U35128 (N_35128,N_32163,N_32528);
and U35129 (N_35129,N_32720,N_32019);
nand U35130 (N_35130,N_33469,N_32127);
nor U35131 (N_35131,N_32857,N_32166);
xnor U35132 (N_35132,N_32581,N_33204);
or U35133 (N_35133,N_32027,N_32591);
or U35134 (N_35134,N_33451,N_32269);
or U35135 (N_35135,N_33607,N_32515);
xnor U35136 (N_35136,N_33269,N_33864);
nor U35137 (N_35137,N_33332,N_32072);
or U35138 (N_35138,N_32343,N_32227);
or U35139 (N_35139,N_33285,N_32560);
nand U35140 (N_35140,N_33903,N_33407);
or U35141 (N_35141,N_32533,N_32411);
or U35142 (N_35142,N_33147,N_32470);
and U35143 (N_35143,N_32821,N_32052);
xor U35144 (N_35144,N_33811,N_33999);
or U35145 (N_35145,N_32427,N_32009);
nor U35146 (N_35146,N_32754,N_32019);
nor U35147 (N_35147,N_33041,N_33903);
and U35148 (N_35148,N_33892,N_32123);
and U35149 (N_35149,N_33773,N_33777);
nor U35150 (N_35150,N_33398,N_33322);
xnor U35151 (N_35151,N_32869,N_33874);
and U35152 (N_35152,N_33741,N_32123);
or U35153 (N_35153,N_33259,N_32849);
and U35154 (N_35154,N_32552,N_32687);
nand U35155 (N_35155,N_33704,N_32939);
and U35156 (N_35156,N_33511,N_33885);
xor U35157 (N_35157,N_32588,N_32126);
nor U35158 (N_35158,N_32453,N_32372);
or U35159 (N_35159,N_32712,N_33343);
xnor U35160 (N_35160,N_33863,N_32302);
xor U35161 (N_35161,N_32739,N_32752);
and U35162 (N_35162,N_33399,N_32869);
xnor U35163 (N_35163,N_32093,N_33001);
nor U35164 (N_35164,N_32509,N_33280);
xor U35165 (N_35165,N_33371,N_32006);
xnor U35166 (N_35166,N_33900,N_32826);
nor U35167 (N_35167,N_32767,N_32673);
nand U35168 (N_35168,N_32774,N_32770);
and U35169 (N_35169,N_33150,N_32750);
nand U35170 (N_35170,N_33942,N_32464);
xor U35171 (N_35171,N_32662,N_33750);
nand U35172 (N_35172,N_33597,N_33444);
xnor U35173 (N_35173,N_32935,N_32735);
nor U35174 (N_35174,N_33092,N_32796);
nand U35175 (N_35175,N_33481,N_33573);
xnor U35176 (N_35176,N_32738,N_32519);
nor U35177 (N_35177,N_33327,N_33495);
and U35178 (N_35178,N_33731,N_32801);
or U35179 (N_35179,N_32969,N_33347);
xor U35180 (N_35180,N_33103,N_33835);
xnor U35181 (N_35181,N_33743,N_33402);
and U35182 (N_35182,N_33179,N_33535);
xor U35183 (N_35183,N_33881,N_32374);
and U35184 (N_35184,N_32607,N_33383);
nand U35185 (N_35185,N_33036,N_33335);
nand U35186 (N_35186,N_33818,N_33387);
xnor U35187 (N_35187,N_32238,N_33801);
nor U35188 (N_35188,N_32385,N_33912);
nand U35189 (N_35189,N_32404,N_33533);
nand U35190 (N_35190,N_32402,N_32844);
and U35191 (N_35191,N_33548,N_32492);
nor U35192 (N_35192,N_32538,N_32072);
or U35193 (N_35193,N_33907,N_33791);
xor U35194 (N_35194,N_32362,N_33976);
xnor U35195 (N_35195,N_32704,N_33375);
nand U35196 (N_35196,N_33012,N_32412);
and U35197 (N_35197,N_32325,N_33395);
nor U35198 (N_35198,N_32510,N_33268);
nand U35199 (N_35199,N_32568,N_32224);
or U35200 (N_35200,N_33250,N_33449);
nor U35201 (N_35201,N_32092,N_32642);
and U35202 (N_35202,N_33145,N_33464);
or U35203 (N_35203,N_32512,N_32361);
nand U35204 (N_35204,N_33695,N_33039);
nand U35205 (N_35205,N_32089,N_32359);
nor U35206 (N_35206,N_32084,N_33894);
nor U35207 (N_35207,N_32129,N_32766);
nor U35208 (N_35208,N_33851,N_33924);
and U35209 (N_35209,N_32155,N_33913);
or U35210 (N_35210,N_33821,N_32672);
xnor U35211 (N_35211,N_32838,N_33085);
xor U35212 (N_35212,N_33861,N_33627);
xor U35213 (N_35213,N_32504,N_33524);
or U35214 (N_35214,N_32696,N_33712);
nor U35215 (N_35215,N_33585,N_32632);
xor U35216 (N_35216,N_32933,N_32938);
nor U35217 (N_35217,N_32654,N_32236);
or U35218 (N_35218,N_32093,N_33240);
nor U35219 (N_35219,N_32670,N_32022);
nor U35220 (N_35220,N_32179,N_32067);
and U35221 (N_35221,N_33774,N_32963);
xnor U35222 (N_35222,N_33803,N_32308);
or U35223 (N_35223,N_33467,N_33801);
nand U35224 (N_35224,N_33321,N_32341);
nand U35225 (N_35225,N_32667,N_33901);
xor U35226 (N_35226,N_33443,N_32146);
and U35227 (N_35227,N_32673,N_32847);
and U35228 (N_35228,N_33272,N_33682);
xnor U35229 (N_35229,N_32504,N_32591);
and U35230 (N_35230,N_33872,N_33798);
or U35231 (N_35231,N_33557,N_33084);
and U35232 (N_35232,N_32811,N_33325);
xor U35233 (N_35233,N_33824,N_32098);
and U35234 (N_35234,N_32445,N_32890);
nand U35235 (N_35235,N_33745,N_32806);
or U35236 (N_35236,N_32448,N_32545);
xor U35237 (N_35237,N_33709,N_32175);
or U35238 (N_35238,N_32834,N_33425);
or U35239 (N_35239,N_33808,N_32190);
xnor U35240 (N_35240,N_33239,N_32101);
or U35241 (N_35241,N_32035,N_33291);
and U35242 (N_35242,N_33064,N_32840);
and U35243 (N_35243,N_33844,N_32779);
or U35244 (N_35244,N_33138,N_32751);
nor U35245 (N_35245,N_33504,N_32212);
or U35246 (N_35246,N_33693,N_32348);
or U35247 (N_35247,N_33548,N_32542);
xnor U35248 (N_35248,N_32305,N_32883);
xor U35249 (N_35249,N_33215,N_33575);
and U35250 (N_35250,N_32367,N_32357);
nand U35251 (N_35251,N_32797,N_32625);
nand U35252 (N_35252,N_33597,N_32553);
or U35253 (N_35253,N_33916,N_32290);
or U35254 (N_35254,N_33535,N_33718);
or U35255 (N_35255,N_33441,N_33629);
and U35256 (N_35256,N_32248,N_33180);
xnor U35257 (N_35257,N_32563,N_33222);
or U35258 (N_35258,N_32189,N_32033);
or U35259 (N_35259,N_32613,N_33140);
xor U35260 (N_35260,N_32122,N_33553);
and U35261 (N_35261,N_32714,N_32646);
and U35262 (N_35262,N_32413,N_33319);
or U35263 (N_35263,N_33983,N_33939);
and U35264 (N_35264,N_33445,N_33497);
and U35265 (N_35265,N_32442,N_32911);
and U35266 (N_35266,N_32088,N_32039);
and U35267 (N_35267,N_32356,N_32539);
and U35268 (N_35268,N_32598,N_33439);
nand U35269 (N_35269,N_33662,N_32470);
nand U35270 (N_35270,N_32830,N_32341);
or U35271 (N_35271,N_32792,N_32842);
xnor U35272 (N_35272,N_32309,N_33290);
nand U35273 (N_35273,N_33997,N_33349);
nor U35274 (N_35274,N_32581,N_33901);
or U35275 (N_35275,N_33735,N_33383);
xor U35276 (N_35276,N_33247,N_33363);
nor U35277 (N_35277,N_32529,N_33976);
xor U35278 (N_35278,N_33860,N_32637);
or U35279 (N_35279,N_33471,N_32522);
nor U35280 (N_35280,N_33129,N_32392);
xnor U35281 (N_35281,N_33980,N_32205);
xnor U35282 (N_35282,N_32369,N_33262);
and U35283 (N_35283,N_32480,N_32970);
or U35284 (N_35284,N_33913,N_33035);
nand U35285 (N_35285,N_33590,N_33302);
or U35286 (N_35286,N_32705,N_33978);
nor U35287 (N_35287,N_32242,N_33441);
or U35288 (N_35288,N_33391,N_33006);
nand U35289 (N_35289,N_32538,N_33540);
nor U35290 (N_35290,N_33245,N_33530);
nor U35291 (N_35291,N_33904,N_32615);
or U35292 (N_35292,N_32023,N_33957);
or U35293 (N_35293,N_33673,N_33966);
or U35294 (N_35294,N_33308,N_33310);
xnor U35295 (N_35295,N_33644,N_32055);
nand U35296 (N_35296,N_32967,N_32264);
xnor U35297 (N_35297,N_32804,N_33954);
xor U35298 (N_35298,N_32200,N_33767);
and U35299 (N_35299,N_32450,N_32124);
and U35300 (N_35300,N_32911,N_32005);
nor U35301 (N_35301,N_32789,N_32267);
and U35302 (N_35302,N_32996,N_32957);
nand U35303 (N_35303,N_33739,N_32710);
nand U35304 (N_35304,N_33424,N_32676);
nand U35305 (N_35305,N_32668,N_33291);
or U35306 (N_35306,N_33583,N_32554);
or U35307 (N_35307,N_33709,N_32630);
xor U35308 (N_35308,N_33233,N_32720);
or U35309 (N_35309,N_32749,N_33414);
nor U35310 (N_35310,N_33043,N_33088);
xor U35311 (N_35311,N_33373,N_33697);
nand U35312 (N_35312,N_33325,N_32124);
nor U35313 (N_35313,N_33064,N_33819);
and U35314 (N_35314,N_32689,N_32549);
xnor U35315 (N_35315,N_32238,N_32848);
or U35316 (N_35316,N_32236,N_32509);
nand U35317 (N_35317,N_32007,N_33271);
xnor U35318 (N_35318,N_33632,N_32973);
or U35319 (N_35319,N_33424,N_33759);
xnor U35320 (N_35320,N_32149,N_33142);
nand U35321 (N_35321,N_33285,N_33008);
or U35322 (N_35322,N_32122,N_33870);
xnor U35323 (N_35323,N_32640,N_32728);
xor U35324 (N_35324,N_33307,N_32361);
xor U35325 (N_35325,N_33116,N_32821);
or U35326 (N_35326,N_33759,N_32459);
nand U35327 (N_35327,N_32159,N_32963);
or U35328 (N_35328,N_33061,N_32247);
nand U35329 (N_35329,N_33254,N_32074);
or U35330 (N_35330,N_32366,N_33548);
or U35331 (N_35331,N_32185,N_32848);
or U35332 (N_35332,N_32303,N_33924);
and U35333 (N_35333,N_32996,N_33157);
nand U35334 (N_35334,N_33963,N_33387);
and U35335 (N_35335,N_33673,N_33926);
xnor U35336 (N_35336,N_32949,N_32647);
nor U35337 (N_35337,N_33767,N_32578);
xnor U35338 (N_35338,N_32787,N_33177);
and U35339 (N_35339,N_33115,N_33984);
xor U35340 (N_35340,N_33058,N_33001);
or U35341 (N_35341,N_32496,N_33147);
xor U35342 (N_35342,N_32388,N_33361);
nand U35343 (N_35343,N_33419,N_32707);
nor U35344 (N_35344,N_32787,N_33200);
and U35345 (N_35345,N_32360,N_32248);
nor U35346 (N_35346,N_33239,N_33217);
and U35347 (N_35347,N_33255,N_32147);
or U35348 (N_35348,N_33022,N_33254);
or U35349 (N_35349,N_32727,N_33092);
or U35350 (N_35350,N_32506,N_33656);
or U35351 (N_35351,N_32639,N_32410);
and U35352 (N_35352,N_33486,N_33487);
or U35353 (N_35353,N_32547,N_33220);
nor U35354 (N_35354,N_32432,N_33366);
and U35355 (N_35355,N_32095,N_32552);
or U35356 (N_35356,N_32262,N_33436);
nor U35357 (N_35357,N_33016,N_32476);
nor U35358 (N_35358,N_33318,N_32571);
nand U35359 (N_35359,N_33676,N_32185);
nand U35360 (N_35360,N_33045,N_33836);
nand U35361 (N_35361,N_33165,N_32040);
nor U35362 (N_35362,N_32947,N_32513);
nand U35363 (N_35363,N_32272,N_33624);
nand U35364 (N_35364,N_32899,N_32125);
nand U35365 (N_35365,N_33466,N_33725);
and U35366 (N_35366,N_32877,N_32055);
or U35367 (N_35367,N_33084,N_32113);
and U35368 (N_35368,N_33534,N_32664);
nor U35369 (N_35369,N_32285,N_32522);
or U35370 (N_35370,N_32077,N_33536);
nor U35371 (N_35371,N_33795,N_33010);
or U35372 (N_35372,N_32672,N_32060);
xor U35373 (N_35373,N_33185,N_32786);
and U35374 (N_35374,N_33572,N_32718);
nor U35375 (N_35375,N_33063,N_32799);
nor U35376 (N_35376,N_32379,N_32320);
xor U35377 (N_35377,N_33528,N_33258);
and U35378 (N_35378,N_33919,N_32010);
nand U35379 (N_35379,N_33643,N_32352);
and U35380 (N_35380,N_33567,N_32133);
and U35381 (N_35381,N_32559,N_33418);
and U35382 (N_35382,N_33724,N_33787);
nand U35383 (N_35383,N_32658,N_32179);
nand U35384 (N_35384,N_33078,N_32958);
and U35385 (N_35385,N_33557,N_33746);
nor U35386 (N_35386,N_32241,N_33470);
or U35387 (N_35387,N_32765,N_33101);
and U35388 (N_35388,N_33280,N_33958);
or U35389 (N_35389,N_33835,N_33358);
xor U35390 (N_35390,N_33197,N_33176);
nand U35391 (N_35391,N_32089,N_32595);
or U35392 (N_35392,N_33186,N_33017);
nor U35393 (N_35393,N_32290,N_33278);
nor U35394 (N_35394,N_33726,N_33798);
or U35395 (N_35395,N_33843,N_33384);
nand U35396 (N_35396,N_32709,N_33453);
nand U35397 (N_35397,N_32663,N_32643);
or U35398 (N_35398,N_32012,N_33204);
xor U35399 (N_35399,N_33715,N_33435);
or U35400 (N_35400,N_32285,N_33667);
xor U35401 (N_35401,N_33859,N_32663);
xor U35402 (N_35402,N_33209,N_32813);
nand U35403 (N_35403,N_33658,N_32543);
and U35404 (N_35404,N_32357,N_33386);
nand U35405 (N_35405,N_32491,N_33251);
nor U35406 (N_35406,N_32905,N_33278);
and U35407 (N_35407,N_32887,N_32542);
nand U35408 (N_35408,N_32708,N_32525);
or U35409 (N_35409,N_32031,N_32318);
or U35410 (N_35410,N_32862,N_33210);
nand U35411 (N_35411,N_32263,N_33443);
and U35412 (N_35412,N_33970,N_33929);
or U35413 (N_35413,N_33254,N_32474);
nand U35414 (N_35414,N_32701,N_32871);
nand U35415 (N_35415,N_32389,N_33388);
or U35416 (N_35416,N_33927,N_32753);
nor U35417 (N_35417,N_33431,N_33479);
or U35418 (N_35418,N_33693,N_33560);
xor U35419 (N_35419,N_33190,N_32993);
nand U35420 (N_35420,N_33762,N_32556);
xor U35421 (N_35421,N_32413,N_33686);
or U35422 (N_35422,N_32961,N_33026);
or U35423 (N_35423,N_33039,N_32642);
xor U35424 (N_35424,N_33851,N_33743);
and U35425 (N_35425,N_33897,N_33790);
xnor U35426 (N_35426,N_33186,N_32015);
nand U35427 (N_35427,N_33229,N_32308);
xnor U35428 (N_35428,N_33032,N_33378);
or U35429 (N_35429,N_33081,N_33913);
xnor U35430 (N_35430,N_33829,N_33361);
or U35431 (N_35431,N_32170,N_32362);
nand U35432 (N_35432,N_32913,N_33824);
xor U35433 (N_35433,N_32347,N_33022);
nand U35434 (N_35434,N_32845,N_32759);
or U35435 (N_35435,N_32701,N_33610);
nor U35436 (N_35436,N_33297,N_33851);
xor U35437 (N_35437,N_33362,N_32362);
or U35438 (N_35438,N_32332,N_33591);
nand U35439 (N_35439,N_33305,N_33603);
and U35440 (N_35440,N_32381,N_33210);
nand U35441 (N_35441,N_33957,N_33100);
nand U35442 (N_35442,N_32272,N_32190);
nand U35443 (N_35443,N_32361,N_32380);
nand U35444 (N_35444,N_32288,N_32876);
xor U35445 (N_35445,N_33312,N_33219);
and U35446 (N_35446,N_32747,N_33878);
or U35447 (N_35447,N_33321,N_33072);
or U35448 (N_35448,N_32122,N_33827);
nor U35449 (N_35449,N_32879,N_33940);
xnor U35450 (N_35450,N_33698,N_33241);
nand U35451 (N_35451,N_33839,N_33272);
and U35452 (N_35452,N_33838,N_33108);
nand U35453 (N_35453,N_32647,N_32605);
nand U35454 (N_35454,N_33057,N_32759);
nand U35455 (N_35455,N_32359,N_33323);
nor U35456 (N_35456,N_32640,N_33599);
nor U35457 (N_35457,N_32566,N_32221);
and U35458 (N_35458,N_33855,N_33812);
or U35459 (N_35459,N_32427,N_32635);
nand U35460 (N_35460,N_32983,N_33422);
nand U35461 (N_35461,N_33271,N_32611);
nand U35462 (N_35462,N_32128,N_32549);
or U35463 (N_35463,N_32092,N_32188);
and U35464 (N_35464,N_32517,N_33771);
nor U35465 (N_35465,N_32848,N_32996);
xnor U35466 (N_35466,N_33686,N_32132);
nand U35467 (N_35467,N_32235,N_32732);
and U35468 (N_35468,N_32601,N_32251);
and U35469 (N_35469,N_32525,N_32706);
nand U35470 (N_35470,N_32925,N_33611);
nand U35471 (N_35471,N_32777,N_33190);
or U35472 (N_35472,N_32037,N_32061);
xor U35473 (N_35473,N_33772,N_33741);
and U35474 (N_35474,N_32824,N_33712);
or U35475 (N_35475,N_33358,N_33447);
xnor U35476 (N_35476,N_32212,N_33478);
xnor U35477 (N_35477,N_32921,N_33292);
nand U35478 (N_35478,N_33384,N_32367);
or U35479 (N_35479,N_33342,N_33952);
or U35480 (N_35480,N_33273,N_33855);
xor U35481 (N_35481,N_33196,N_32236);
nor U35482 (N_35482,N_32402,N_33743);
nand U35483 (N_35483,N_32763,N_33359);
xnor U35484 (N_35484,N_32804,N_33623);
nand U35485 (N_35485,N_33430,N_33624);
or U35486 (N_35486,N_32360,N_33907);
and U35487 (N_35487,N_33026,N_32380);
and U35488 (N_35488,N_33478,N_33233);
and U35489 (N_35489,N_33689,N_32066);
xor U35490 (N_35490,N_33764,N_33660);
xnor U35491 (N_35491,N_33130,N_32051);
or U35492 (N_35492,N_32844,N_33983);
nand U35493 (N_35493,N_33831,N_32808);
nor U35494 (N_35494,N_33792,N_33964);
and U35495 (N_35495,N_32892,N_33263);
or U35496 (N_35496,N_32813,N_33680);
and U35497 (N_35497,N_32019,N_32481);
xnor U35498 (N_35498,N_32748,N_32973);
xnor U35499 (N_35499,N_33845,N_32515);
nand U35500 (N_35500,N_33454,N_33993);
and U35501 (N_35501,N_32981,N_33991);
nor U35502 (N_35502,N_33531,N_33053);
and U35503 (N_35503,N_32457,N_32015);
and U35504 (N_35504,N_33414,N_33208);
xor U35505 (N_35505,N_33154,N_33373);
nand U35506 (N_35506,N_33456,N_33692);
nor U35507 (N_35507,N_33794,N_32773);
or U35508 (N_35508,N_33986,N_33379);
xnor U35509 (N_35509,N_32509,N_33991);
xnor U35510 (N_35510,N_33746,N_33206);
nor U35511 (N_35511,N_33724,N_33142);
or U35512 (N_35512,N_32661,N_33339);
nor U35513 (N_35513,N_33134,N_32996);
or U35514 (N_35514,N_32441,N_32695);
xnor U35515 (N_35515,N_32786,N_32571);
nor U35516 (N_35516,N_33643,N_33368);
xnor U35517 (N_35517,N_33860,N_32017);
nand U35518 (N_35518,N_32950,N_32031);
nor U35519 (N_35519,N_32951,N_32860);
or U35520 (N_35520,N_32280,N_32228);
xnor U35521 (N_35521,N_33663,N_32923);
nor U35522 (N_35522,N_32626,N_32968);
xnor U35523 (N_35523,N_33290,N_32444);
or U35524 (N_35524,N_32321,N_32973);
or U35525 (N_35525,N_33423,N_33522);
nand U35526 (N_35526,N_32310,N_33309);
or U35527 (N_35527,N_32499,N_32224);
nor U35528 (N_35528,N_33676,N_32250);
or U35529 (N_35529,N_32014,N_32778);
nor U35530 (N_35530,N_32736,N_33284);
xor U35531 (N_35531,N_33329,N_32773);
and U35532 (N_35532,N_33105,N_32445);
or U35533 (N_35533,N_32326,N_32501);
and U35534 (N_35534,N_32541,N_33401);
nor U35535 (N_35535,N_33630,N_33588);
or U35536 (N_35536,N_33312,N_32437);
and U35537 (N_35537,N_32006,N_32186);
or U35538 (N_35538,N_33041,N_33673);
nor U35539 (N_35539,N_33612,N_32423);
xnor U35540 (N_35540,N_33615,N_32490);
or U35541 (N_35541,N_33022,N_32190);
nor U35542 (N_35542,N_33975,N_32378);
and U35543 (N_35543,N_33491,N_33726);
or U35544 (N_35544,N_33017,N_33805);
nor U35545 (N_35545,N_33204,N_32238);
nor U35546 (N_35546,N_32553,N_33861);
nand U35547 (N_35547,N_33135,N_33427);
or U35548 (N_35548,N_33418,N_32388);
xnor U35549 (N_35549,N_32747,N_33441);
and U35550 (N_35550,N_32545,N_32644);
nor U35551 (N_35551,N_33185,N_33004);
and U35552 (N_35552,N_32605,N_32381);
nor U35553 (N_35553,N_32837,N_33458);
and U35554 (N_35554,N_33174,N_33096);
nor U35555 (N_35555,N_33656,N_33420);
or U35556 (N_35556,N_33823,N_33332);
or U35557 (N_35557,N_32860,N_32954);
nor U35558 (N_35558,N_33672,N_33859);
and U35559 (N_35559,N_33781,N_33419);
nor U35560 (N_35560,N_33154,N_32830);
or U35561 (N_35561,N_33269,N_32481);
or U35562 (N_35562,N_33016,N_33554);
xnor U35563 (N_35563,N_32520,N_32669);
xnor U35564 (N_35564,N_33814,N_33821);
nor U35565 (N_35565,N_32565,N_32836);
xor U35566 (N_35566,N_33425,N_32644);
nand U35567 (N_35567,N_33842,N_33861);
and U35568 (N_35568,N_33665,N_33522);
nor U35569 (N_35569,N_33894,N_33602);
nand U35570 (N_35570,N_32364,N_33935);
xor U35571 (N_35571,N_33882,N_33219);
xor U35572 (N_35572,N_32616,N_33900);
nand U35573 (N_35573,N_32202,N_33358);
xnor U35574 (N_35574,N_33250,N_33116);
nand U35575 (N_35575,N_33523,N_33774);
nor U35576 (N_35576,N_32568,N_33117);
nand U35577 (N_35577,N_33461,N_33748);
nor U35578 (N_35578,N_33288,N_33759);
or U35579 (N_35579,N_33518,N_32527);
nor U35580 (N_35580,N_32200,N_33071);
nand U35581 (N_35581,N_33145,N_33809);
xor U35582 (N_35582,N_32450,N_33829);
and U35583 (N_35583,N_33507,N_33892);
xor U35584 (N_35584,N_32343,N_33724);
nor U35585 (N_35585,N_32627,N_33519);
nand U35586 (N_35586,N_33877,N_32357);
nand U35587 (N_35587,N_33659,N_32786);
nor U35588 (N_35588,N_32921,N_33353);
nand U35589 (N_35589,N_32683,N_32657);
and U35590 (N_35590,N_33301,N_32543);
or U35591 (N_35591,N_33230,N_33045);
nor U35592 (N_35592,N_32177,N_32748);
nor U35593 (N_35593,N_32977,N_32948);
or U35594 (N_35594,N_32309,N_33632);
nor U35595 (N_35595,N_32712,N_32154);
xnor U35596 (N_35596,N_32298,N_32562);
nor U35597 (N_35597,N_33504,N_32806);
and U35598 (N_35598,N_33523,N_32272);
nor U35599 (N_35599,N_33458,N_33038);
nor U35600 (N_35600,N_32353,N_32667);
or U35601 (N_35601,N_32194,N_33757);
and U35602 (N_35602,N_32994,N_32035);
or U35603 (N_35603,N_33196,N_32037);
and U35604 (N_35604,N_32623,N_33882);
and U35605 (N_35605,N_32028,N_32527);
and U35606 (N_35606,N_33225,N_32121);
or U35607 (N_35607,N_32472,N_32250);
nor U35608 (N_35608,N_32242,N_32766);
or U35609 (N_35609,N_33046,N_33654);
and U35610 (N_35610,N_33075,N_33365);
or U35611 (N_35611,N_33732,N_32053);
nor U35612 (N_35612,N_32333,N_33605);
nand U35613 (N_35613,N_33920,N_33469);
and U35614 (N_35614,N_32056,N_32611);
xor U35615 (N_35615,N_33905,N_32877);
and U35616 (N_35616,N_32553,N_32699);
and U35617 (N_35617,N_32351,N_33483);
xnor U35618 (N_35618,N_33523,N_32904);
and U35619 (N_35619,N_33681,N_33767);
or U35620 (N_35620,N_32753,N_33853);
nand U35621 (N_35621,N_32210,N_33286);
or U35622 (N_35622,N_33135,N_33644);
or U35623 (N_35623,N_33984,N_33643);
nand U35624 (N_35624,N_32722,N_33497);
and U35625 (N_35625,N_32226,N_32720);
and U35626 (N_35626,N_32408,N_32843);
xnor U35627 (N_35627,N_33322,N_32559);
or U35628 (N_35628,N_32016,N_33589);
or U35629 (N_35629,N_33084,N_33639);
nor U35630 (N_35630,N_33881,N_32226);
or U35631 (N_35631,N_33522,N_32226);
or U35632 (N_35632,N_33443,N_32559);
xor U35633 (N_35633,N_32638,N_33718);
or U35634 (N_35634,N_32167,N_33164);
and U35635 (N_35635,N_32778,N_32256);
and U35636 (N_35636,N_33385,N_32388);
nand U35637 (N_35637,N_32786,N_33404);
xnor U35638 (N_35638,N_33676,N_32748);
nand U35639 (N_35639,N_33429,N_32730);
nand U35640 (N_35640,N_33336,N_32708);
xor U35641 (N_35641,N_32654,N_33396);
and U35642 (N_35642,N_33871,N_33739);
nand U35643 (N_35643,N_33428,N_32854);
xor U35644 (N_35644,N_32914,N_32794);
nor U35645 (N_35645,N_32966,N_32852);
nor U35646 (N_35646,N_33110,N_33361);
and U35647 (N_35647,N_32307,N_32052);
and U35648 (N_35648,N_33031,N_32271);
or U35649 (N_35649,N_32929,N_33532);
nor U35650 (N_35650,N_33941,N_33544);
nor U35651 (N_35651,N_33480,N_32530);
nand U35652 (N_35652,N_33276,N_32537);
or U35653 (N_35653,N_32308,N_33522);
nor U35654 (N_35654,N_33121,N_32105);
xor U35655 (N_35655,N_32262,N_33503);
nor U35656 (N_35656,N_32132,N_32050);
and U35657 (N_35657,N_32048,N_32202);
and U35658 (N_35658,N_32696,N_32694);
nor U35659 (N_35659,N_32401,N_32617);
xor U35660 (N_35660,N_32431,N_32986);
nor U35661 (N_35661,N_32815,N_32414);
nor U35662 (N_35662,N_32175,N_33394);
nor U35663 (N_35663,N_32910,N_32900);
or U35664 (N_35664,N_32969,N_32583);
xor U35665 (N_35665,N_32668,N_32384);
xor U35666 (N_35666,N_32707,N_33799);
or U35667 (N_35667,N_33124,N_33741);
nor U35668 (N_35668,N_32460,N_32291);
and U35669 (N_35669,N_33315,N_32235);
or U35670 (N_35670,N_33433,N_33789);
xor U35671 (N_35671,N_33410,N_32703);
xor U35672 (N_35672,N_33460,N_32842);
or U35673 (N_35673,N_32069,N_33979);
xor U35674 (N_35674,N_32971,N_32010);
or U35675 (N_35675,N_33804,N_32107);
nand U35676 (N_35676,N_33971,N_32604);
or U35677 (N_35677,N_32722,N_32319);
xor U35678 (N_35678,N_32375,N_33679);
or U35679 (N_35679,N_33700,N_33732);
nor U35680 (N_35680,N_33517,N_32838);
or U35681 (N_35681,N_32209,N_32366);
nor U35682 (N_35682,N_33898,N_32537);
nor U35683 (N_35683,N_33789,N_33578);
nor U35684 (N_35684,N_33089,N_33938);
nor U35685 (N_35685,N_33738,N_33008);
xor U35686 (N_35686,N_33733,N_33754);
and U35687 (N_35687,N_33912,N_33001);
and U35688 (N_35688,N_33838,N_32408);
xnor U35689 (N_35689,N_33671,N_32899);
nand U35690 (N_35690,N_33098,N_33948);
nor U35691 (N_35691,N_33196,N_33409);
and U35692 (N_35692,N_33734,N_32090);
or U35693 (N_35693,N_32828,N_32540);
and U35694 (N_35694,N_33347,N_32483);
and U35695 (N_35695,N_32087,N_33733);
nand U35696 (N_35696,N_33881,N_33174);
xor U35697 (N_35697,N_33356,N_32294);
and U35698 (N_35698,N_33157,N_32916);
or U35699 (N_35699,N_33626,N_32327);
nand U35700 (N_35700,N_32973,N_33242);
or U35701 (N_35701,N_33491,N_32461);
and U35702 (N_35702,N_33957,N_33979);
or U35703 (N_35703,N_32541,N_33310);
nand U35704 (N_35704,N_33405,N_32365);
nor U35705 (N_35705,N_33224,N_33663);
nor U35706 (N_35706,N_32437,N_33954);
or U35707 (N_35707,N_32216,N_33532);
or U35708 (N_35708,N_32313,N_32049);
or U35709 (N_35709,N_32488,N_33195);
or U35710 (N_35710,N_32563,N_32938);
xor U35711 (N_35711,N_33213,N_32199);
nor U35712 (N_35712,N_32495,N_33895);
xor U35713 (N_35713,N_33487,N_33836);
or U35714 (N_35714,N_32183,N_32274);
nand U35715 (N_35715,N_33377,N_33645);
nor U35716 (N_35716,N_32266,N_32146);
nand U35717 (N_35717,N_32748,N_33709);
or U35718 (N_35718,N_32879,N_33359);
nand U35719 (N_35719,N_32515,N_32571);
and U35720 (N_35720,N_32409,N_32998);
xnor U35721 (N_35721,N_33191,N_32605);
xnor U35722 (N_35722,N_32696,N_32257);
nor U35723 (N_35723,N_32081,N_32804);
xor U35724 (N_35724,N_32525,N_32260);
and U35725 (N_35725,N_33992,N_33296);
or U35726 (N_35726,N_32946,N_33527);
xor U35727 (N_35727,N_32540,N_32560);
nand U35728 (N_35728,N_33767,N_32168);
xnor U35729 (N_35729,N_33389,N_33301);
nor U35730 (N_35730,N_33270,N_33234);
nand U35731 (N_35731,N_33174,N_33196);
or U35732 (N_35732,N_33755,N_32155);
xnor U35733 (N_35733,N_33839,N_33371);
or U35734 (N_35734,N_32105,N_33451);
and U35735 (N_35735,N_32177,N_32481);
xor U35736 (N_35736,N_32165,N_32916);
nand U35737 (N_35737,N_32396,N_32420);
or U35738 (N_35738,N_32340,N_32210);
xor U35739 (N_35739,N_32702,N_32692);
nand U35740 (N_35740,N_32531,N_32530);
nand U35741 (N_35741,N_32631,N_32013);
xor U35742 (N_35742,N_33782,N_32530);
nand U35743 (N_35743,N_32844,N_33601);
or U35744 (N_35744,N_33399,N_32589);
xor U35745 (N_35745,N_33501,N_33825);
xnor U35746 (N_35746,N_33270,N_32127);
and U35747 (N_35747,N_33646,N_32626);
or U35748 (N_35748,N_32947,N_32204);
or U35749 (N_35749,N_33057,N_33116);
and U35750 (N_35750,N_33244,N_32853);
and U35751 (N_35751,N_33036,N_33350);
nor U35752 (N_35752,N_33637,N_33393);
xor U35753 (N_35753,N_33803,N_32931);
nand U35754 (N_35754,N_33800,N_32550);
xor U35755 (N_35755,N_33879,N_33122);
nor U35756 (N_35756,N_33849,N_33617);
nor U35757 (N_35757,N_33491,N_33463);
nand U35758 (N_35758,N_32171,N_32597);
and U35759 (N_35759,N_32664,N_32100);
nor U35760 (N_35760,N_33249,N_32315);
nor U35761 (N_35761,N_32904,N_33654);
or U35762 (N_35762,N_32998,N_32882);
and U35763 (N_35763,N_32352,N_32217);
xnor U35764 (N_35764,N_32710,N_33119);
or U35765 (N_35765,N_32381,N_33059);
nor U35766 (N_35766,N_33333,N_33012);
nor U35767 (N_35767,N_32689,N_32836);
xor U35768 (N_35768,N_33275,N_33788);
nand U35769 (N_35769,N_33124,N_33413);
xor U35770 (N_35770,N_33912,N_32159);
and U35771 (N_35771,N_33943,N_33564);
and U35772 (N_35772,N_33481,N_33821);
nor U35773 (N_35773,N_32082,N_32531);
and U35774 (N_35774,N_33989,N_33742);
nand U35775 (N_35775,N_33666,N_32124);
and U35776 (N_35776,N_32403,N_33813);
or U35777 (N_35777,N_32879,N_32947);
nor U35778 (N_35778,N_32744,N_32889);
nor U35779 (N_35779,N_33962,N_33446);
and U35780 (N_35780,N_32882,N_32029);
xor U35781 (N_35781,N_33273,N_32209);
xnor U35782 (N_35782,N_32545,N_32310);
nor U35783 (N_35783,N_32552,N_32784);
and U35784 (N_35784,N_33546,N_32291);
xor U35785 (N_35785,N_32822,N_32936);
nand U35786 (N_35786,N_33806,N_32505);
xor U35787 (N_35787,N_32010,N_33953);
or U35788 (N_35788,N_32337,N_32312);
nor U35789 (N_35789,N_33451,N_32095);
or U35790 (N_35790,N_33339,N_33224);
or U35791 (N_35791,N_33283,N_32146);
xnor U35792 (N_35792,N_32947,N_32647);
nor U35793 (N_35793,N_33929,N_32055);
nor U35794 (N_35794,N_33083,N_33201);
nand U35795 (N_35795,N_33798,N_32382);
xor U35796 (N_35796,N_33743,N_33329);
and U35797 (N_35797,N_33402,N_33290);
and U35798 (N_35798,N_32664,N_32103);
nand U35799 (N_35799,N_32092,N_32076);
and U35800 (N_35800,N_32234,N_32482);
or U35801 (N_35801,N_33310,N_33621);
or U35802 (N_35802,N_33869,N_32431);
nor U35803 (N_35803,N_33311,N_33962);
nor U35804 (N_35804,N_33001,N_33660);
or U35805 (N_35805,N_32350,N_32082);
nand U35806 (N_35806,N_33499,N_33456);
and U35807 (N_35807,N_33333,N_33309);
or U35808 (N_35808,N_33731,N_32257);
xnor U35809 (N_35809,N_32085,N_33257);
and U35810 (N_35810,N_33766,N_32382);
nor U35811 (N_35811,N_33554,N_33124);
nand U35812 (N_35812,N_32746,N_33563);
and U35813 (N_35813,N_32328,N_32568);
nor U35814 (N_35814,N_32159,N_33076);
or U35815 (N_35815,N_33342,N_33492);
xor U35816 (N_35816,N_32930,N_32489);
or U35817 (N_35817,N_32082,N_32442);
or U35818 (N_35818,N_33705,N_33810);
or U35819 (N_35819,N_32810,N_33891);
and U35820 (N_35820,N_33422,N_32372);
nand U35821 (N_35821,N_33426,N_32022);
and U35822 (N_35822,N_33938,N_33757);
nor U35823 (N_35823,N_33418,N_32714);
nand U35824 (N_35824,N_33059,N_33124);
or U35825 (N_35825,N_33943,N_32625);
xnor U35826 (N_35826,N_33679,N_33212);
nor U35827 (N_35827,N_33696,N_32218);
nand U35828 (N_35828,N_33655,N_32385);
and U35829 (N_35829,N_33290,N_32581);
or U35830 (N_35830,N_32115,N_32322);
nand U35831 (N_35831,N_32094,N_33871);
and U35832 (N_35832,N_32983,N_32695);
nor U35833 (N_35833,N_33410,N_33768);
xnor U35834 (N_35834,N_33786,N_32833);
xnor U35835 (N_35835,N_32744,N_33365);
or U35836 (N_35836,N_33848,N_33952);
or U35837 (N_35837,N_32869,N_33620);
or U35838 (N_35838,N_33282,N_32584);
xor U35839 (N_35839,N_33504,N_33353);
and U35840 (N_35840,N_33520,N_33578);
or U35841 (N_35841,N_33263,N_32210);
and U35842 (N_35842,N_33596,N_33802);
or U35843 (N_35843,N_32737,N_32187);
or U35844 (N_35844,N_33079,N_32847);
and U35845 (N_35845,N_33942,N_33981);
and U35846 (N_35846,N_33812,N_33849);
and U35847 (N_35847,N_33484,N_32186);
xor U35848 (N_35848,N_33756,N_32945);
xor U35849 (N_35849,N_32114,N_33841);
nand U35850 (N_35850,N_32113,N_32482);
or U35851 (N_35851,N_33419,N_32261);
nand U35852 (N_35852,N_33231,N_32018);
nor U35853 (N_35853,N_32657,N_33933);
and U35854 (N_35854,N_32573,N_33795);
nor U35855 (N_35855,N_32776,N_32487);
nor U35856 (N_35856,N_32941,N_33091);
xor U35857 (N_35857,N_33236,N_32805);
and U35858 (N_35858,N_33428,N_32036);
or U35859 (N_35859,N_33658,N_33125);
and U35860 (N_35860,N_33215,N_33922);
nor U35861 (N_35861,N_33851,N_32465);
nand U35862 (N_35862,N_33064,N_32734);
nand U35863 (N_35863,N_32476,N_33507);
nor U35864 (N_35864,N_33010,N_32444);
nand U35865 (N_35865,N_32747,N_33533);
nor U35866 (N_35866,N_33007,N_33405);
xor U35867 (N_35867,N_32732,N_32027);
nor U35868 (N_35868,N_33301,N_33963);
nand U35869 (N_35869,N_32725,N_33488);
and U35870 (N_35870,N_33219,N_33084);
nand U35871 (N_35871,N_32555,N_33052);
xnor U35872 (N_35872,N_33079,N_33105);
nand U35873 (N_35873,N_32132,N_32531);
and U35874 (N_35874,N_33639,N_33826);
nor U35875 (N_35875,N_33685,N_33367);
xnor U35876 (N_35876,N_33969,N_33860);
or U35877 (N_35877,N_33667,N_33560);
and U35878 (N_35878,N_33077,N_32213);
nor U35879 (N_35879,N_32101,N_33346);
and U35880 (N_35880,N_33368,N_33961);
nand U35881 (N_35881,N_33967,N_32491);
and U35882 (N_35882,N_33079,N_32059);
or U35883 (N_35883,N_33686,N_32049);
nand U35884 (N_35884,N_32253,N_32233);
or U35885 (N_35885,N_33828,N_33636);
nand U35886 (N_35886,N_32957,N_33538);
nand U35887 (N_35887,N_32286,N_32527);
xnor U35888 (N_35888,N_32932,N_32034);
nor U35889 (N_35889,N_33661,N_32845);
nand U35890 (N_35890,N_32369,N_32776);
nand U35891 (N_35891,N_33870,N_32867);
or U35892 (N_35892,N_33653,N_32907);
xnor U35893 (N_35893,N_32199,N_32031);
nand U35894 (N_35894,N_33077,N_32229);
nand U35895 (N_35895,N_33691,N_33060);
nor U35896 (N_35896,N_32066,N_33715);
and U35897 (N_35897,N_32139,N_33347);
nor U35898 (N_35898,N_32168,N_33528);
and U35899 (N_35899,N_32579,N_33167);
xor U35900 (N_35900,N_32640,N_33876);
nand U35901 (N_35901,N_33926,N_32394);
and U35902 (N_35902,N_33763,N_32118);
or U35903 (N_35903,N_32762,N_32203);
nand U35904 (N_35904,N_32524,N_32715);
and U35905 (N_35905,N_32790,N_33608);
nor U35906 (N_35906,N_33741,N_33852);
and U35907 (N_35907,N_33035,N_32890);
nand U35908 (N_35908,N_32570,N_32079);
or U35909 (N_35909,N_32522,N_32043);
or U35910 (N_35910,N_32904,N_33146);
xnor U35911 (N_35911,N_33213,N_32138);
and U35912 (N_35912,N_32603,N_32363);
nor U35913 (N_35913,N_33949,N_32928);
and U35914 (N_35914,N_32040,N_32650);
and U35915 (N_35915,N_32332,N_33622);
and U35916 (N_35916,N_33623,N_33053);
nor U35917 (N_35917,N_33310,N_33586);
nand U35918 (N_35918,N_32512,N_32723);
xnor U35919 (N_35919,N_32420,N_32778);
and U35920 (N_35920,N_32538,N_33953);
and U35921 (N_35921,N_33285,N_32889);
xnor U35922 (N_35922,N_33394,N_32090);
nor U35923 (N_35923,N_32759,N_33434);
xnor U35924 (N_35924,N_33871,N_32695);
and U35925 (N_35925,N_33344,N_33845);
xor U35926 (N_35926,N_33594,N_32244);
nand U35927 (N_35927,N_33253,N_32827);
and U35928 (N_35928,N_33635,N_33529);
or U35929 (N_35929,N_33206,N_33028);
xnor U35930 (N_35930,N_33852,N_33956);
xnor U35931 (N_35931,N_32283,N_33448);
xor U35932 (N_35932,N_33919,N_33360);
xnor U35933 (N_35933,N_33220,N_32964);
xor U35934 (N_35934,N_33284,N_32629);
or U35935 (N_35935,N_33758,N_32457);
or U35936 (N_35936,N_33912,N_32545);
xor U35937 (N_35937,N_32758,N_33709);
and U35938 (N_35938,N_33908,N_33757);
or U35939 (N_35939,N_32492,N_32486);
nand U35940 (N_35940,N_33848,N_33221);
nand U35941 (N_35941,N_32540,N_33787);
or U35942 (N_35942,N_33843,N_33728);
nand U35943 (N_35943,N_32184,N_32352);
nand U35944 (N_35944,N_33592,N_33096);
nand U35945 (N_35945,N_33131,N_32487);
nand U35946 (N_35946,N_32336,N_33259);
xor U35947 (N_35947,N_33317,N_33685);
nor U35948 (N_35948,N_32690,N_32014);
and U35949 (N_35949,N_32903,N_33146);
xor U35950 (N_35950,N_33450,N_32941);
xnor U35951 (N_35951,N_33225,N_32141);
and U35952 (N_35952,N_33162,N_32146);
xnor U35953 (N_35953,N_32406,N_32481);
xor U35954 (N_35954,N_33292,N_33654);
and U35955 (N_35955,N_32832,N_32804);
nor U35956 (N_35956,N_32757,N_32347);
nor U35957 (N_35957,N_33722,N_33667);
nor U35958 (N_35958,N_33523,N_32629);
nor U35959 (N_35959,N_33232,N_33389);
xor U35960 (N_35960,N_32503,N_32155);
xor U35961 (N_35961,N_32440,N_33984);
and U35962 (N_35962,N_33253,N_33586);
or U35963 (N_35963,N_32381,N_32138);
nor U35964 (N_35964,N_33585,N_33526);
xnor U35965 (N_35965,N_33556,N_33566);
xor U35966 (N_35966,N_32748,N_32371);
or U35967 (N_35967,N_33477,N_32417);
nor U35968 (N_35968,N_32350,N_33225);
xnor U35969 (N_35969,N_32579,N_32449);
nand U35970 (N_35970,N_32715,N_33879);
nand U35971 (N_35971,N_32274,N_32144);
nor U35972 (N_35972,N_32281,N_32055);
and U35973 (N_35973,N_33514,N_32393);
and U35974 (N_35974,N_32587,N_33423);
xnor U35975 (N_35975,N_32993,N_33494);
nand U35976 (N_35976,N_32246,N_33076);
or U35977 (N_35977,N_32761,N_33267);
nand U35978 (N_35978,N_32475,N_33456);
nor U35979 (N_35979,N_33387,N_32604);
and U35980 (N_35980,N_33745,N_33079);
xnor U35981 (N_35981,N_32095,N_33703);
nand U35982 (N_35982,N_32728,N_32920);
and U35983 (N_35983,N_32206,N_32983);
or U35984 (N_35984,N_33420,N_32131);
xnor U35985 (N_35985,N_32568,N_33699);
nor U35986 (N_35986,N_33432,N_33040);
xnor U35987 (N_35987,N_32348,N_32286);
xor U35988 (N_35988,N_33052,N_33371);
xnor U35989 (N_35989,N_32270,N_33504);
nor U35990 (N_35990,N_33157,N_33898);
xor U35991 (N_35991,N_32366,N_32386);
xor U35992 (N_35992,N_33797,N_33050);
and U35993 (N_35993,N_33527,N_32541);
nor U35994 (N_35994,N_33687,N_33206);
or U35995 (N_35995,N_32999,N_33369);
or U35996 (N_35996,N_33322,N_33752);
xor U35997 (N_35997,N_33662,N_33985);
xnor U35998 (N_35998,N_33517,N_32737);
xor U35999 (N_35999,N_33025,N_33049);
and U36000 (N_36000,N_35581,N_34319);
or U36001 (N_36001,N_34550,N_35768);
and U36002 (N_36002,N_34078,N_35019);
and U36003 (N_36003,N_35122,N_34137);
nor U36004 (N_36004,N_35337,N_35355);
or U36005 (N_36005,N_34810,N_34777);
or U36006 (N_36006,N_35309,N_34228);
nand U36007 (N_36007,N_35843,N_35054);
nand U36008 (N_36008,N_35953,N_35312);
and U36009 (N_36009,N_34034,N_35669);
nor U36010 (N_36010,N_35009,N_35363);
and U36011 (N_36011,N_34676,N_34757);
nand U36012 (N_36012,N_34576,N_34920);
xnor U36013 (N_36013,N_34555,N_35408);
nor U36014 (N_36014,N_35657,N_34043);
nor U36015 (N_36015,N_35992,N_35066);
and U36016 (N_36016,N_35892,N_35690);
and U36017 (N_36017,N_35274,N_34915);
nand U36018 (N_36018,N_34285,N_35960);
and U36019 (N_36019,N_35810,N_35488);
nor U36020 (N_36020,N_35152,N_35649);
or U36021 (N_36021,N_35084,N_34296);
and U36022 (N_36022,N_34792,N_35571);
xnor U36023 (N_36023,N_35787,N_35039);
or U36024 (N_36024,N_35117,N_35077);
or U36025 (N_36025,N_34141,N_35275);
nor U36026 (N_36026,N_34859,N_35942);
nor U36027 (N_36027,N_35530,N_35969);
or U36028 (N_36028,N_34683,N_35387);
xor U36029 (N_36029,N_34451,N_35986);
xnor U36030 (N_36030,N_34302,N_34601);
xor U36031 (N_36031,N_35006,N_34769);
nand U36032 (N_36032,N_35413,N_34875);
nor U36033 (N_36033,N_35265,N_35766);
and U36034 (N_36034,N_35906,N_34771);
or U36035 (N_36035,N_34347,N_34816);
or U36036 (N_36036,N_34329,N_35146);
and U36037 (N_36037,N_35799,N_35051);
and U36038 (N_36038,N_34307,N_34570);
nor U36039 (N_36039,N_35638,N_35923);
xor U36040 (N_36040,N_35391,N_35747);
and U36041 (N_36041,N_35439,N_34582);
and U36042 (N_36042,N_34866,N_35703);
xor U36043 (N_36043,N_34617,N_35852);
or U36044 (N_36044,N_34821,N_35813);
or U36045 (N_36045,N_34391,N_35620);
xnor U36046 (N_36046,N_35547,N_35036);
and U36047 (N_36047,N_35398,N_34912);
and U36048 (N_36048,N_35007,N_34359);
nor U36049 (N_36049,N_35695,N_35206);
or U36050 (N_36050,N_35842,N_34208);
nand U36051 (N_36051,N_35815,N_34877);
or U36052 (N_36052,N_35708,N_34348);
and U36053 (N_36053,N_34349,N_34313);
nor U36054 (N_36054,N_34626,N_34533);
nand U36055 (N_36055,N_35368,N_34179);
nor U36056 (N_36056,N_35110,N_35560);
xnor U36057 (N_36057,N_35893,N_35131);
and U36058 (N_36058,N_35797,N_34140);
or U36059 (N_36059,N_35691,N_35565);
xnor U36060 (N_36060,N_35882,N_35971);
xor U36061 (N_36061,N_34910,N_34764);
xnor U36062 (N_36062,N_35831,N_34428);
and U36063 (N_36063,N_34178,N_34463);
xnor U36064 (N_36064,N_35607,N_35151);
nor U36065 (N_36065,N_35144,N_34352);
nor U36066 (N_36066,N_35556,N_35168);
and U36067 (N_36067,N_34674,N_34196);
xor U36068 (N_36068,N_34580,N_34107);
nand U36069 (N_36069,N_34223,N_35042);
or U36070 (N_36070,N_34686,N_34464);
xnor U36071 (N_36071,N_35086,N_34725);
nor U36072 (N_36072,N_35466,N_34990);
and U36073 (N_36073,N_34204,N_35423);
nor U36074 (N_36074,N_34827,N_35235);
or U36075 (N_36075,N_35481,N_35771);
and U36076 (N_36076,N_34907,N_34603);
or U36077 (N_36077,N_35016,N_35229);
nor U36078 (N_36078,N_35934,N_35770);
or U36079 (N_36079,N_34691,N_34409);
and U36080 (N_36080,N_34526,N_34508);
nor U36081 (N_36081,N_35932,N_35908);
nand U36082 (N_36082,N_34500,N_35062);
or U36083 (N_36083,N_34088,N_35231);
nand U36084 (N_36084,N_34480,N_35411);
nand U36085 (N_36085,N_35385,N_35814);
and U36086 (N_36086,N_34211,N_34387);
xnor U36087 (N_36087,N_34786,N_34321);
nor U36088 (N_36088,N_35984,N_34744);
nand U36089 (N_36089,N_35271,N_35765);
or U36090 (N_36090,N_34331,N_34880);
or U36091 (N_36091,N_35078,N_35030);
or U36092 (N_36092,N_35660,N_34712);
and U36093 (N_36093,N_34728,N_35407);
xor U36094 (N_36094,N_35247,N_34344);
xnor U36095 (N_36095,N_35433,N_34644);
nor U36096 (N_36096,N_35314,N_34678);
nand U36097 (N_36097,N_34439,N_35748);
xnor U36098 (N_36098,N_34556,N_35327);
nor U36099 (N_36099,N_35313,N_34536);
or U36100 (N_36100,N_34099,N_35979);
xor U36101 (N_36101,N_34432,N_34899);
or U36102 (N_36102,N_35319,N_35197);
and U36103 (N_36103,N_34559,N_35844);
nor U36104 (N_36104,N_35501,N_34001);
nand U36105 (N_36105,N_34488,N_35092);
and U36106 (N_36106,N_35603,N_35273);
xor U36107 (N_36107,N_35344,N_35455);
nand U36108 (N_36108,N_34849,N_34087);
nor U36109 (N_36109,N_34896,N_35647);
nand U36110 (N_36110,N_34273,N_34578);
or U36111 (N_36111,N_35332,N_35448);
or U36112 (N_36112,N_34942,N_35622);
nand U36113 (N_36113,N_34950,N_35033);
nand U36114 (N_36114,N_35619,N_34798);
and U36115 (N_36115,N_34693,N_34783);
nand U36116 (N_36116,N_34024,N_35272);
nand U36117 (N_36117,N_34278,N_34962);
nand U36118 (N_36118,N_34665,N_35330);
nand U36119 (N_36119,N_35471,N_35203);
or U36120 (N_36120,N_34926,N_34322);
nand U36121 (N_36121,N_35359,N_34145);
or U36122 (N_36122,N_34188,N_35700);
and U36123 (N_36123,N_35219,N_35937);
xor U36124 (N_36124,N_34602,N_34294);
or U36125 (N_36125,N_34544,N_34660);
and U36126 (N_36126,N_35989,N_34510);
and U36127 (N_36127,N_35419,N_34354);
nand U36128 (N_36128,N_35749,N_35472);
and U36129 (N_36129,N_35060,N_34413);
xnor U36130 (N_36130,N_34543,N_35890);
xnor U36131 (N_36131,N_35237,N_35631);
nor U36132 (N_36132,N_35089,N_35477);
nor U36133 (N_36133,N_34879,N_35410);
or U36134 (N_36134,N_34969,N_34079);
or U36135 (N_36135,N_34721,N_34241);
or U36136 (N_36136,N_34637,N_34906);
nand U36137 (N_36137,N_35069,N_35339);
xor U36138 (N_36138,N_35948,N_34383);
xnor U36139 (N_36139,N_34641,N_35345);
xor U36140 (N_36140,N_34271,N_35106);
nand U36141 (N_36141,N_34070,N_34103);
and U36142 (N_36142,N_35280,N_35491);
xnor U36143 (N_36143,N_35524,N_35812);
and U36144 (N_36144,N_35927,N_35181);
or U36145 (N_36145,N_35268,N_34521);
nor U36146 (N_36146,N_34680,N_35982);
or U36147 (N_36147,N_35869,N_34606);
and U36148 (N_36148,N_35426,N_34856);
nor U36149 (N_36149,N_34668,N_35452);
and U36150 (N_36150,N_35511,N_35564);
or U36151 (N_36151,N_35162,N_34484);
nor U36152 (N_36152,N_34441,N_34889);
or U36153 (N_36153,N_34339,N_34921);
xor U36154 (N_36154,N_34945,N_35907);
nor U36155 (N_36155,N_35721,N_35136);
or U36156 (N_36156,N_34151,N_34068);
or U36157 (N_36157,N_35236,N_34939);
or U36158 (N_36158,N_34052,N_35075);
nor U36159 (N_36159,N_34826,N_35580);
nand U36160 (N_36160,N_34397,N_34876);
nand U36161 (N_36161,N_35329,N_34288);
nand U36162 (N_36162,N_34878,N_34191);
xor U36163 (N_36163,N_34624,N_35230);
and U36164 (N_36164,N_34527,N_35296);
xor U36165 (N_36165,N_35487,N_34963);
xnor U36166 (N_36166,N_34916,N_35712);
and U36167 (N_36167,N_35090,N_34564);
xor U36168 (N_36168,N_34454,N_35588);
and U36169 (N_36169,N_35990,N_35840);
nand U36170 (N_36170,N_35256,N_34724);
or U36171 (N_36171,N_35111,N_35824);
nand U36172 (N_36172,N_34973,N_35742);
xnor U36173 (N_36173,N_35114,N_34027);
xnor U36174 (N_36174,N_35284,N_35085);
nor U36175 (N_36175,N_34577,N_35196);
and U36176 (N_36176,N_34206,N_34420);
nand U36177 (N_36177,N_35262,N_35605);
nand U36178 (N_36178,N_34654,N_35393);
nor U36179 (N_36179,N_35474,N_34146);
xnor U36180 (N_36180,N_35017,N_35846);
nor U36181 (N_36181,N_34247,N_35267);
nor U36182 (N_36182,N_35753,N_34740);
nand U36183 (N_36183,N_34264,N_34529);
nor U36184 (N_36184,N_34845,N_35138);
or U36185 (N_36185,N_34108,N_34489);
xor U36186 (N_36186,N_35072,N_34227);
nor U36187 (N_36187,N_35772,N_34639);
nor U36188 (N_36188,N_35174,N_35563);
nand U36189 (N_36189,N_35397,N_35902);
xor U36190 (N_36190,N_35884,N_35277);
and U36191 (N_36191,N_34595,N_34540);
nand U36192 (N_36192,N_34888,N_34590);
nor U36193 (N_36193,N_34730,N_35709);
nor U36194 (N_36194,N_34496,N_34634);
nand U36195 (N_36195,N_34584,N_35755);
or U36196 (N_36196,N_35951,N_35848);
nor U36197 (N_36197,N_35653,N_34933);
nor U36198 (N_36198,N_34890,N_34064);
or U36199 (N_36199,N_34780,N_34987);
xor U36200 (N_36200,N_35671,N_35276);
or U36201 (N_36201,N_34325,N_34310);
or U36202 (N_36202,N_35324,N_35165);
xor U36203 (N_36203,N_34796,N_35128);
xnor U36204 (N_36204,N_35602,N_35743);
xor U36205 (N_36205,N_35762,N_34225);
or U36206 (N_36206,N_35298,N_35819);
nand U36207 (N_36207,N_35285,N_35282);
xnor U36208 (N_36208,N_34868,N_34411);
and U36209 (N_36209,N_34563,N_35055);
or U36210 (N_36210,N_35475,N_35454);
nand U36211 (N_36211,N_34162,N_34588);
nand U36212 (N_36212,N_34483,N_34265);
xor U36213 (N_36213,N_35751,N_34279);
nor U36214 (N_36214,N_34170,N_35167);
nand U36215 (N_36215,N_35912,N_34673);
xor U36216 (N_36216,N_34406,N_34793);
nor U36217 (N_36217,N_35034,N_35290);
and U36218 (N_36218,N_34884,N_35105);
or U36219 (N_36219,N_35680,N_34186);
nand U36220 (N_36220,N_34739,N_35803);
nand U36221 (N_36221,N_35909,N_34927);
xnor U36222 (N_36222,N_35716,N_34328);
nand U36223 (N_36223,N_35453,N_35401);
and U36224 (N_36224,N_35598,N_34938);
nor U36225 (N_36225,N_35470,N_34476);
or U36226 (N_36226,N_34605,N_34551);
or U36227 (N_36227,N_34971,N_34787);
and U36228 (N_36228,N_34373,N_34882);
nor U36229 (N_36229,N_35566,N_34158);
nor U36230 (N_36230,N_34532,N_35880);
or U36231 (N_36231,N_35378,N_35182);
nor U36232 (N_36232,N_35507,N_35479);
or U36233 (N_36233,N_34013,N_35014);
nor U36234 (N_36234,N_34004,N_34689);
nor U36235 (N_36235,N_35253,N_35379);
or U36236 (N_36236,N_35793,N_34525);
xor U36237 (N_36237,N_34459,N_34135);
or U36238 (N_36238,N_35301,N_35925);
nor U36239 (N_36239,N_34478,N_34604);
nand U36240 (N_36240,N_35694,N_34643);
xor U36241 (N_36241,N_35795,N_35013);
and U36242 (N_36242,N_34823,N_35866);
nor U36243 (N_36243,N_34440,N_34804);
nor U36244 (N_36244,N_35183,N_35210);
or U36245 (N_36245,N_34520,N_34364);
nor U36246 (N_36246,N_34185,N_35807);
xnor U36247 (N_36247,N_35510,N_34911);
and U36248 (N_36248,N_34066,N_35881);
xor U36249 (N_36249,N_35008,N_34200);
or U36250 (N_36250,N_35446,N_34295);
or U36251 (N_36251,N_34717,N_34812);
nand U36252 (N_36252,N_35946,N_34369);
xnor U36253 (N_36253,N_34873,N_34591);
xnor U36254 (N_36254,N_35922,N_35554);
or U36255 (N_36255,N_35279,N_34799);
xor U36256 (N_36256,N_35447,N_35593);
nor U36257 (N_36257,N_35873,N_35356);
nor U36258 (N_36258,N_35914,N_35321);
xor U36259 (N_36259,N_34988,N_34970);
xor U36260 (N_36260,N_35185,N_34198);
xor U36261 (N_36261,N_35246,N_34549);
xnor U36262 (N_36262,N_34118,N_35575);
xor U36263 (N_36263,N_34519,N_35630);
or U36264 (N_36264,N_34380,N_34977);
nor U36265 (N_36265,N_35916,N_34234);
or U36266 (N_36266,N_34233,N_34006);
and U36267 (N_36267,N_34281,N_35940);
or U36268 (N_36268,N_34240,N_34738);
xor U36269 (N_36269,N_34702,N_34197);
or U36270 (N_36270,N_35143,N_34610);
xor U36271 (N_36271,N_35546,N_35505);
xnor U36272 (N_36272,N_34424,N_34579);
or U36273 (N_36273,N_34030,N_35295);
and U36274 (N_36274,N_35140,N_34136);
or U36275 (N_36275,N_35692,N_34060);
nand U36276 (N_36276,N_35429,N_35839);
and U36277 (N_36277,N_34433,N_34524);
nor U36278 (N_36278,N_34415,N_35137);
xnor U36279 (N_36279,N_35050,N_34860);
or U36280 (N_36280,N_34401,N_34254);
nor U36281 (N_36281,N_34340,N_35370);
xor U36282 (N_36282,N_35970,N_34566);
nand U36283 (N_36283,N_34713,N_34572);
or U36284 (N_36284,N_34573,N_35957);
xor U36285 (N_36285,N_34893,N_35048);
or U36286 (N_36286,N_34897,N_34710);
and U36287 (N_36287,N_35888,N_34306);
nand U36288 (N_36288,N_34688,N_34018);
or U36289 (N_36289,N_34308,N_34954);
xor U36290 (N_36290,N_34023,N_35264);
or U36291 (N_36291,N_34327,N_34841);
or U36292 (N_36292,N_34160,N_34708);
nor U36293 (N_36293,N_34869,N_35905);
nand U36294 (N_36294,N_34377,N_35894);
and U36295 (N_36295,N_34669,N_35781);
and U36296 (N_36296,N_35561,N_34357);
or U36297 (N_36297,N_34941,N_35776);
nand U36298 (N_36298,N_35543,N_34913);
xnor U36299 (N_36299,N_35679,N_34129);
or U36300 (N_36300,N_35641,N_34423);
nand U36301 (N_36301,N_35896,N_35788);
nand U36302 (N_36302,N_34256,N_35107);
nor U36303 (N_36303,N_34502,N_35629);
nor U36304 (N_36304,N_35318,N_35664);
nor U36305 (N_36305,N_35040,N_34266);
nand U36306 (N_36306,N_34994,N_34919);
or U36307 (N_36307,N_35763,N_34671);
and U36308 (N_36308,N_34038,N_35412);
xor U36309 (N_36309,N_34119,N_34512);
and U36310 (N_36310,N_34305,N_35856);
nor U36311 (N_36311,N_35160,N_35886);
nand U36312 (N_36312,N_34967,N_35025);
and U36313 (N_36313,N_35129,N_34957);
and U36314 (N_36314,N_34600,N_35043);
or U36315 (N_36315,N_34366,N_34632);
nand U36316 (N_36316,N_35502,N_34737);
nor U36317 (N_36317,N_35931,N_34597);
and U36318 (N_36318,N_35158,N_35492);
or U36319 (N_36319,N_34917,N_34652);
xnor U36320 (N_36320,N_34486,N_35608);
nor U36321 (N_36321,N_34169,N_35464);
or U36322 (N_36322,N_34017,N_34163);
nor U36323 (N_36323,N_35021,N_35098);
or U36324 (N_36324,N_35764,N_35933);
nand U36325 (N_36325,N_34164,N_35746);
nor U36326 (N_36326,N_34210,N_35095);
and U36327 (N_36327,N_35949,N_35745);
nor U36328 (N_36328,N_34250,N_34336);
xnor U36329 (N_36329,N_35395,N_35585);
or U36330 (N_36330,N_35698,N_34057);
xor U36331 (N_36331,N_35835,N_34820);
nand U36332 (N_36332,N_35228,N_35540);
nand U36333 (N_36333,N_34040,N_35473);
nand U36334 (N_36334,N_35785,N_35968);
xnor U36335 (N_36335,N_34803,N_34097);
nand U36336 (N_36336,N_34147,N_35737);
nor U36337 (N_36337,N_34019,N_34855);
xor U36338 (N_36338,N_34286,N_34007);
and U36339 (N_36339,N_35650,N_35609);
xnor U36340 (N_36340,N_34337,N_34468);
nor U36341 (N_36341,N_34828,N_35670);
xor U36342 (N_36342,N_34785,N_34871);
nand U36343 (N_36343,N_34386,N_34358);
nand U36344 (N_36344,N_34898,N_35930);
and U36345 (N_36345,N_34334,N_34086);
or U36346 (N_36346,N_35861,N_35023);
and U36347 (N_36347,N_35241,N_35676);
nor U36348 (N_36348,N_35364,N_35738);
nor U36349 (N_36349,N_35809,N_35226);
nor U36350 (N_36350,N_34682,N_35517);
or U36351 (N_36351,N_35857,N_35833);
xor U36352 (N_36352,N_34113,N_35515);
nand U36353 (N_36353,N_34449,N_35616);
and U36354 (N_36354,N_34966,N_34640);
or U36355 (N_36355,N_35663,N_34650);
or U36356 (N_36356,N_34000,N_35555);
and U36357 (N_36357,N_34759,N_35335);
nor U36358 (N_36358,N_34231,N_35366);
or U36359 (N_36359,N_34784,N_34788);
and U36360 (N_36360,N_34132,N_34466);
or U36361 (N_36361,N_35333,N_35263);
and U36362 (N_36362,N_35444,N_34883);
nand U36363 (N_36363,N_34053,N_34155);
or U36364 (N_36364,N_34914,N_34090);
or U36365 (N_36365,N_34042,N_35214);
nand U36366 (N_36366,N_34649,N_35683);
and U36367 (N_36367,N_35245,N_35983);
xnor U36368 (N_36368,N_35950,N_34716);
and U36369 (N_36369,N_34100,N_34242);
xnor U36370 (N_36370,N_35482,N_34505);
nand U36371 (N_36371,N_34416,N_34367);
or U36372 (N_36372,N_35134,N_35340);
xor U36373 (N_36373,N_35065,N_35029);
xnor U36374 (N_36374,N_35283,N_34012);
xnor U36375 (N_36375,N_34159,N_34323);
and U36376 (N_36376,N_34473,N_35438);
xor U36377 (N_36377,N_34753,N_34861);
or U36378 (N_36378,N_35300,N_35323);
nor U36379 (N_36379,N_35775,N_35915);
and U36380 (N_36380,N_34209,N_34620);
or U36381 (N_36381,N_34677,N_35348);
and U36382 (N_36382,N_35760,N_34156);
nor U36383 (N_36383,N_34809,N_35727);
and U36384 (N_36384,N_35929,N_35792);
xor U36385 (N_36385,N_34045,N_34182);
nand U36386 (N_36386,N_34585,N_35678);
xnor U36387 (N_36387,N_35613,N_34244);
xnor U36388 (N_36388,N_35667,N_35921);
xnor U36389 (N_36389,N_35381,N_34684);
nor U36390 (N_36390,N_35503,N_34049);
and U36391 (N_36391,N_35082,N_35686);
and U36392 (N_36392,N_35287,N_35919);
or U36393 (N_36393,N_34157,N_34028);
nor U36394 (N_36394,N_34504,N_34944);
nand U36395 (N_36395,N_34404,N_35028);
nor U36396 (N_36396,N_34734,N_34438);
and U36397 (N_36397,N_35935,N_34080);
and U36398 (N_36398,N_34427,N_35123);
nand U36399 (N_36399,N_35701,N_34760);
and U36400 (N_36400,N_34341,N_34462);
and U36401 (N_36401,N_35222,N_34201);
nor U36402 (N_36402,N_34393,N_34983);
or U36403 (N_36403,N_35544,N_35903);
or U36404 (N_36404,N_35463,N_34048);
xor U36405 (N_36405,N_34122,N_34445);
nor U36406 (N_36406,N_35221,N_34862);
nand U36407 (N_36407,N_35514,N_34239);
nor U36408 (N_36408,N_34986,N_35533);
or U36409 (N_36409,N_35414,N_34335);
or U36410 (N_36410,N_35999,N_34951);
and U36411 (N_36411,N_34382,N_34324);
xnor U36412 (N_36412,N_34270,N_34457);
nand U36413 (N_36413,N_35046,N_35436);
or U36414 (N_36414,N_34928,N_34840);
nand U36415 (N_36415,N_35617,N_34695);
xnor U36416 (N_36416,N_34047,N_35673);
and U36417 (N_36417,N_35910,N_35526);
and U36418 (N_36418,N_35254,N_34022);
or U36419 (N_36419,N_34276,N_34732);
and U36420 (N_36420,N_34554,N_35154);
and U36421 (N_36421,N_34666,N_34607);
or U36422 (N_36422,N_35292,N_35855);
or U36423 (N_36423,N_35467,N_34645);
or U36424 (N_36424,N_34538,N_34565);
and U36425 (N_36425,N_35947,N_35244);
nor U36426 (N_36426,N_34735,N_35100);
xnor U36427 (N_36427,N_35595,N_35976);
and U36428 (N_36428,N_35791,N_35088);
nand U36429 (N_36429,N_34098,N_34356);
or U36430 (N_36430,N_34700,N_35723);
or U36431 (N_36431,N_34465,N_35227);
or U36432 (N_36432,N_34125,N_34332);
nand U36433 (N_36433,N_34779,N_35080);
or U36434 (N_36434,N_34586,N_34736);
nor U36435 (N_36435,N_35794,N_34104);
nand U36436 (N_36436,N_35572,N_34518);
xnor U36437 (N_36437,N_34093,N_35194);
nor U36438 (N_36438,N_34059,N_34199);
xnor U36439 (N_36439,N_34929,N_34283);
xor U36440 (N_36440,N_34035,N_35186);
nor U36441 (N_36441,N_35829,N_35594);
nand U36442 (N_36442,N_34282,N_35371);
and U36443 (N_36443,N_35315,N_35898);
or U36444 (N_36444,N_34979,N_35633);
and U36445 (N_36445,N_34854,N_34371);
or U36446 (N_36446,N_34515,N_34690);
nor U36447 (N_36447,N_35901,N_34263);
and U36448 (N_36448,N_34539,N_35952);
xnor U36449 (N_36449,N_35103,N_35782);
xnor U36450 (N_36450,N_34814,N_35003);
or U36451 (N_36451,N_34778,N_35035);
and U36452 (N_36452,N_34709,N_34835);
nand U36453 (N_36453,N_35218,N_35534);
or U36454 (N_36454,N_34943,N_35443);
or U36455 (N_36455,N_34338,N_35045);
and U36456 (N_36456,N_35827,N_35132);
nor U36457 (N_36457,N_35325,N_35331);
and U36458 (N_36458,N_34836,N_34569);
and U36459 (N_36459,N_34900,N_35420);
or U36460 (N_36460,N_34594,N_34032);
nor U36461 (N_36461,N_35451,N_35459);
nand U36462 (N_36462,N_35926,N_34036);
and U36463 (N_36463,N_34742,N_34268);
nand U36464 (N_36464,N_34701,N_35954);
or U36465 (N_36465,N_34016,N_35523);
or U36466 (N_36466,N_35442,N_35834);
or U36467 (N_36467,N_34870,N_34745);
nand U36468 (N_36468,N_34442,N_35118);
and U36469 (N_36469,N_34635,N_34455);
or U36470 (N_36470,N_35112,N_34202);
or U36471 (N_36471,N_35821,N_35317);
nor U36472 (N_36472,N_35557,N_34842);
or U36473 (N_36473,N_35462,N_34982);
xnor U36474 (N_36474,N_35156,N_35148);
nand U36475 (N_36475,N_34394,N_34999);
xor U36476 (N_36476,N_34167,N_35841);
xnor U36477 (N_36477,N_34523,N_34763);
and U36478 (N_36478,N_34694,N_34405);
nor U36479 (N_36479,N_35071,N_35600);
nand U36480 (N_36480,N_34940,N_34333);
nor U36481 (N_36481,N_34217,N_34894);
xor U36482 (N_36482,N_35399,N_35297);
nor U36483 (N_36483,N_35532,N_34984);
and U36484 (N_36484,N_34429,N_35512);
xor U36485 (N_36485,N_34011,N_35731);
xor U36486 (N_36486,N_35711,N_34936);
xor U36487 (N_36487,N_34997,N_35961);
or U36488 (N_36488,N_35542,N_34120);
nand U36489 (N_36489,N_34758,N_35405);
or U36490 (N_36490,N_35739,N_34485);
nand U36491 (N_36491,N_35991,N_34948);
nand U36492 (N_36492,N_35494,N_34838);
xnor U36493 (N_36493,N_35083,N_34472);
xor U36494 (N_36494,N_34959,N_35239);
xnor U36495 (N_36495,N_34507,N_34790);
nor U36496 (N_36496,N_35484,N_34008);
nor U36497 (N_36497,N_34667,N_34995);
nor U36498 (N_36498,N_35293,N_35707);
or U36499 (N_36499,N_34117,N_35212);
xnor U36500 (N_36500,N_34857,N_34316);
nor U36501 (N_36501,N_34575,N_34499);
nor U36502 (N_36502,N_35562,N_34831);
or U36503 (N_36503,N_34289,N_35538);
nand U36504 (N_36504,N_34166,N_34291);
or U36505 (N_36505,N_34370,N_35139);
nand U36506 (N_36506,N_35305,N_35553);
xor U36507 (N_36507,N_35718,N_34687);
nor U36508 (N_36508,N_34501,N_35918);
xor U36509 (N_36509,N_35975,N_34298);
nand U36510 (N_36510,N_34662,N_35885);
and U36511 (N_36511,N_34976,N_35769);
nand U36512 (N_36512,N_35115,N_34748);
nand U36513 (N_36513,N_34553,N_35980);
and U36514 (N_36514,N_35266,N_34075);
xnor U36515 (N_36515,N_35924,N_35779);
or U36516 (N_36516,N_35208,N_34255);
xnor U36517 (N_36517,N_34794,N_35962);
xnor U36518 (N_36518,N_34714,N_35658);
and U36519 (N_36519,N_35351,N_34243);
nor U36520 (N_36520,N_34450,N_35578);
xor U36521 (N_36521,N_35859,N_34353);
or U36522 (N_36522,N_35858,N_35281);
xnor U36523 (N_36523,N_35400,N_34245);
and U36524 (N_36524,N_35796,N_34458);
nand U36525 (N_36525,N_34627,N_34773);
and U36526 (N_36526,N_35874,N_35802);
nor U36527 (N_36527,N_34924,N_34622);
xnor U36528 (N_36528,N_34487,N_35644);
and U36529 (N_36529,N_35871,N_34062);
nor U36530 (N_36530,N_35224,N_35234);
or U36531 (N_36531,N_34084,N_35627);
nor U36532 (N_36532,N_34881,N_34096);
and U36533 (N_36533,N_34698,N_34619);
nand U36534 (N_36534,N_34629,N_34557);
nor U36535 (N_36535,N_35242,N_34046);
nor U36536 (N_36536,N_34902,N_35015);
xor U36537 (N_36537,N_34772,N_35959);
nor U36538 (N_36538,N_34214,N_34848);
nand U36539 (N_36539,N_35498,N_34762);
and U36540 (N_36540,N_35551,N_34259);
nand U36541 (N_36541,N_35830,N_34699);
nor U36542 (N_36542,N_35891,N_34418);
nand U36543 (N_36543,N_35406,N_35403);
nor U36544 (N_36544,N_35800,N_34885);
and U36545 (N_36545,N_35645,N_35939);
and U36546 (N_36546,N_35632,N_35685);
xnor U36547 (N_36547,N_34301,N_34608);
nor U36548 (N_36548,N_34275,N_35804);
or U36549 (N_36549,N_34776,N_35735);
and U36550 (N_36550,N_35611,N_34598);
and U36551 (N_36551,N_34002,N_35715);
nand U36552 (N_36552,N_34326,N_35087);
or U36553 (N_36553,N_35187,N_34203);
and U36554 (N_36554,N_34949,N_34355);
or U36555 (N_36555,N_34761,N_35125);
nand U36556 (N_36556,N_35497,N_34138);
nand U36557 (N_36557,N_34221,N_35116);
or U36558 (N_36558,N_34277,N_34946);
xnor U36559 (N_36559,N_35646,N_35291);
nand U36560 (N_36560,N_34832,N_35981);
xnor U36561 (N_36561,N_35099,N_35596);
or U36562 (N_36562,N_35207,N_35719);
nor U36563 (N_36563,N_35037,N_34083);
nor U36564 (N_36564,N_34363,N_35548);
xor U36565 (N_36565,N_34350,N_34131);
and U36566 (N_36566,N_34829,N_34453);
nor U36567 (N_36567,N_34697,N_34216);
nand U36568 (N_36568,N_35714,N_34041);
xor U36569 (N_36569,N_34446,N_35178);
or U36570 (N_36570,N_35101,N_35801);
or U36571 (N_36571,N_35702,N_34077);
and U36572 (N_36572,N_35361,N_34213);
and U36573 (N_36573,N_35574,N_35863);
and U36574 (N_36574,N_35064,N_34102);
nand U36575 (N_36575,N_35441,N_34830);
nand U36576 (N_36576,N_35161,N_35259);
xor U36577 (N_36577,N_35404,N_34651);
and U36578 (N_36578,N_35599,N_34765);
or U36579 (N_36579,N_34267,N_35648);
nor U36580 (N_36580,N_35465,N_35063);
nor U36581 (N_36581,N_35468,N_35637);
nor U36582 (N_36582,N_35820,N_35710);
nor U36583 (N_36583,N_35868,N_35175);
or U36584 (N_36584,N_34568,N_34139);
nand U36585 (N_36585,N_34300,N_35248);
nor U36586 (N_36586,N_35539,N_34503);
xor U36587 (N_36587,N_35618,N_35899);
or U36588 (N_36588,N_34351,N_35334);
nor U36589 (N_36589,N_35020,N_35357);
nor U36590 (N_36590,N_34297,N_35081);
or U36591 (N_36591,N_34567,N_35238);
or U36592 (N_36592,N_34031,N_35604);
and U36593 (N_36593,N_34646,N_34904);
or U36594 (N_36594,N_34426,N_35872);
xor U36595 (N_36595,N_35163,N_35496);
and U36596 (N_36596,N_34249,N_35978);
or U36597 (N_36597,N_34749,N_35102);
and U36598 (N_36598,N_34116,N_34101);
nand U36599 (N_36599,N_34768,N_34839);
nand U36600 (N_36600,N_34054,N_34766);
nand U36601 (N_36601,N_35730,N_34587);
or U36602 (N_36602,N_34747,N_34037);
and U36603 (N_36603,N_35286,N_35386);
and U36604 (N_36604,N_35260,N_34692);
nor U36605 (N_36605,N_34490,N_35320);
xnor U36606 (N_36606,N_34703,N_35659);
or U36607 (N_36607,N_35490,N_34781);
and U36608 (N_36608,N_34398,N_34562);
xor U36609 (N_36609,N_34109,N_35258);
and U36610 (N_36610,N_34891,N_35577);
xor U36611 (N_36611,N_34599,N_35149);
or U36612 (N_36612,N_34818,N_34630);
nor U36613 (N_36613,N_34726,N_35079);
or U36614 (N_36614,N_35853,N_35010);
nand U36615 (N_36615,N_35000,N_35392);
nand U36616 (N_36616,N_34092,N_35130);
nand U36617 (N_36617,N_34126,N_34867);
xor U36618 (N_36618,N_34051,N_35499);
nand U36619 (N_36619,N_35093,N_35427);
xnor U36620 (N_36620,N_34985,N_34299);
or U36621 (N_36621,N_35220,N_35688);
or U36622 (N_36622,N_34130,N_34447);
nor U36623 (N_36623,N_34851,N_35967);
and U36624 (N_36624,N_34516,N_34782);
and U36625 (N_36625,N_35166,N_34212);
nor U36626 (N_36626,N_34647,N_34317);
nand U36627 (N_36627,N_34152,N_35754);
and U36628 (N_36628,N_35252,N_35058);
and U36629 (N_36629,N_35699,N_34082);
xnor U36630 (N_36630,N_35153,N_35536);
xnor U36631 (N_36631,N_35875,N_35270);
or U36632 (N_36632,N_35624,N_34246);
and U36633 (N_36633,N_35904,N_34705);
nand U36634 (N_36634,N_35722,N_35249);
nor U36635 (N_36635,N_34376,N_35550);
and U36636 (N_36636,N_35535,N_34506);
and U36637 (N_36637,N_34509,N_34612);
and U36638 (N_36638,N_34180,N_35195);
xor U36639 (N_36639,N_35431,N_34530);
nor U36640 (N_36640,N_34303,N_34395);
or U36641 (N_36641,N_35876,N_34314);
or U36642 (N_36642,N_34304,N_34791);
or U36643 (N_36643,N_35583,N_35338);
and U36644 (N_36644,N_35150,N_34542);
nor U36645 (N_36645,N_34365,N_34010);
or U36646 (N_36646,N_35373,N_34552);
and U36647 (N_36647,N_35941,N_34653);
nand U36648 (N_36648,N_34173,N_34105);
or U36649 (N_36649,N_34410,N_35693);
nand U36650 (N_36650,N_35377,N_35074);
xor U36651 (N_36651,N_35059,N_35587);
xor U36652 (N_36652,N_34648,N_35311);
xnor U36653 (N_36653,N_34061,N_34795);
and U36654 (N_36654,N_35198,N_34805);
or U36655 (N_36655,N_35726,N_34574);
xor U36656 (N_36656,N_35750,N_35216);
and U36657 (N_36657,N_35592,N_35394);
or U36658 (N_36658,N_34611,N_35380);
nand U36659 (N_36659,N_35612,N_35654);
or U36660 (N_36660,N_34589,N_34494);
nand U36661 (N_36661,N_35350,N_35205);
or U36662 (N_36662,N_35987,N_34437);
nand U36663 (N_36663,N_34238,N_34696);
or U36664 (N_36664,N_34148,N_35303);
xor U36665 (N_36665,N_34961,N_34864);
nand U36666 (N_36666,N_35525,N_35666);
and U36667 (N_36667,N_34181,N_34252);
and U36668 (N_36668,N_34495,N_34127);
or U36669 (N_36669,N_35997,N_35360);
and U36670 (N_36670,N_35289,N_34149);
nor U36671 (N_36671,N_35837,N_35002);
nor U36672 (N_36672,N_35774,N_35193);
xnor U36673 (N_36673,N_34850,N_35516);
xor U36674 (N_36674,N_35545,N_35601);
nand U36675 (N_36675,N_34901,N_34378);
nor U36676 (N_36676,N_35870,N_35917);
nand U36677 (N_36677,N_35278,N_35460);
and U36678 (N_36678,N_34154,N_34375);
xor U36679 (N_36679,N_35142,N_35073);
nand U36680 (N_36680,N_35883,N_35428);
and U36681 (N_36681,N_35798,N_35269);
and U36682 (N_36682,N_35589,N_35591);
or U36683 (N_36683,N_35860,N_35145);
and U36684 (N_36684,N_34143,N_34858);
nand U36685 (N_36685,N_34903,N_34069);
nand U36686 (N_36686,N_34661,N_34545);
or U36687 (N_36687,N_35573,N_34421);
nor U36688 (N_36688,N_34153,N_34005);
nor U36689 (N_36689,N_35867,N_34479);
and U36690 (N_36690,N_35421,N_35159);
and U36691 (N_36691,N_34800,N_35651);
xor U36692 (N_36692,N_35031,N_35945);
or U36693 (N_36693,N_35251,N_35109);
or U36694 (N_36694,N_34293,N_35635);
xnor U36695 (N_36695,N_35308,N_34020);
or U36696 (N_36696,N_34558,N_35963);
xnor U36697 (N_36697,N_35586,N_35164);
nand U36698 (N_36698,N_34260,N_34414);
xnor U36699 (N_36699,N_35450,N_34592);
nand U36700 (N_36700,N_35567,N_35864);
xnor U36701 (N_36701,N_34968,N_35850);
nor U36702 (N_36702,N_35674,N_34150);
nor U36703 (N_36703,N_34396,N_35728);
and U36704 (N_36704,N_34908,N_35508);
or U36705 (N_36705,N_35897,N_34436);
nand U36706 (N_36706,N_35347,N_34360);
or U36707 (N_36707,N_35456,N_35636);
and U36708 (N_36708,N_35784,N_34616);
and U36709 (N_36709,N_34021,N_35172);
and U36710 (N_36710,N_34237,N_35041);
nor U36711 (N_36711,N_34727,N_34822);
and U36712 (N_36712,N_34315,N_35200);
or U36713 (N_36713,N_35180,N_34284);
nand U36714 (N_36714,N_34165,N_35661);
nor U36715 (N_36715,N_34392,N_34089);
or U36716 (N_36716,N_35372,N_34039);
xor U36717 (N_36717,N_35173,N_35920);
xnor U36718 (N_36718,N_34114,N_35818);
and U36719 (N_36719,N_34195,N_35761);
nand U36720 (N_36720,N_34422,N_34115);
xor U36721 (N_36721,N_35425,N_34847);
xor U36722 (N_36722,N_35549,N_35486);
and U36723 (N_36723,N_35675,N_35847);
xnor U36724 (N_36724,N_35384,N_35495);
nor U36725 (N_36725,N_35445,N_35326);
nor U36726 (N_36726,N_35988,N_34704);
and U36727 (N_36727,N_35354,N_35985);
and U36728 (N_36728,N_34220,N_34715);
or U36729 (N_36729,N_34583,N_35528);
and U36730 (N_36730,N_34679,N_35422);
and U36731 (N_36731,N_35121,N_34384);
nand U36732 (N_36732,N_34419,N_34953);
nor U36733 (N_36733,N_35211,N_35570);
and U36734 (N_36734,N_35038,N_35744);
or U36735 (N_36735,N_35005,N_35382);
xor U36736 (N_36736,N_34955,N_34824);
nor U36737 (N_36737,N_34681,N_35966);
or U36738 (N_36738,N_34205,N_34846);
xor U36739 (N_36739,N_34571,N_35358);
xnor U36740 (N_36740,N_34723,N_35302);
xnor U36741 (N_36741,N_35606,N_35108);
and U36742 (N_36742,N_35067,N_35133);
xnor U36743 (N_36743,N_34482,N_35944);
nor U36744 (N_36744,N_35733,N_35758);
xnor U36745 (N_36745,N_35169,N_34183);
or U36746 (N_36746,N_34817,N_34931);
or U36747 (N_36747,N_34535,N_34235);
or U36748 (N_36748,N_34513,N_35584);
nor U36749 (N_36749,N_34134,N_34311);
and U36750 (N_36750,N_35346,N_35026);
nand U36751 (N_36751,N_35457,N_35705);
xnor U36752 (N_36752,N_34222,N_35367);
xor U36753 (N_36753,N_35643,N_34189);
or U36754 (N_36754,N_35519,N_35878);
or U36755 (N_36755,N_34345,N_35192);
nor U36756 (N_36756,N_34399,N_35011);
nand U36757 (N_36757,N_35004,N_34361);
and U36758 (N_36758,N_34287,N_35135);
or U36759 (N_36759,N_35189,N_35889);
nor U36760 (N_36760,N_35724,N_34342);
xnor U36761 (N_36761,N_34412,N_35342);
nor U36762 (N_36762,N_34534,N_34972);
xnor U36763 (N_36763,N_35956,N_34947);
nand U36764 (N_36764,N_35811,N_35958);
nor U36765 (N_36765,N_34174,N_34318);
nor U36766 (N_36766,N_35094,N_35642);
nand U36767 (N_36767,N_34865,N_35199);
nor U36768 (N_36768,N_35826,N_35068);
nor U36769 (N_36769,N_34091,N_35662);
nor U36770 (N_36770,N_34176,N_34733);
nor U36771 (N_36771,N_35500,N_34443);
or U36772 (N_36772,N_35449,N_35849);
or U36773 (N_36773,N_34144,N_34932);
and U36774 (N_36774,N_34381,N_35955);
and U36775 (N_36775,N_35900,N_34343);
or U36776 (N_36776,N_34161,N_34657);
or U36777 (N_36777,N_34236,N_34905);
nand U36778 (N_36778,N_34067,N_34843);
nor U36779 (N_36779,N_35529,N_35854);
nor U36780 (N_36780,N_35232,N_35170);
and U36781 (N_36781,N_34111,N_35687);
or U36782 (N_36782,N_35365,N_35634);
xor U36783 (N_36783,N_35684,N_35097);
nand U36784 (N_36784,N_35823,N_35832);
and U36785 (N_36785,N_35489,N_34330);
nor U36786 (N_36786,N_35936,N_34470);
and U36787 (N_36787,N_34751,N_34292);
nand U36788 (N_36788,N_35943,N_35147);
nor U36789 (N_36789,N_35250,N_35729);
nand U36790 (N_36790,N_35049,N_35623);
xnor U36791 (N_36791,N_35240,N_35522);
nor U36792 (N_36792,N_35773,N_34224);
nand U36793 (N_36793,N_35822,N_35440);
xor U36794 (N_36794,N_35299,N_34815);
nor U36795 (N_36795,N_35582,N_34755);
nor U36796 (N_36796,N_34133,N_34388);
nand U36797 (N_36797,N_35640,N_34033);
nor U36798 (N_36798,N_35012,N_34980);
nor U36799 (N_36799,N_35928,N_35434);
or U36800 (N_36800,N_35126,N_35998);
nand U36801 (N_36801,N_34852,N_34514);
xnor U36802 (N_36802,N_34493,N_35417);
nor U36803 (N_36803,N_34718,N_34063);
nand U36804 (N_36804,N_34374,N_35838);
or U36805 (N_36805,N_34801,N_35288);
and U36806 (N_36806,N_34672,N_34797);
nor U36807 (N_36807,N_34491,N_35204);
or U36808 (N_36808,N_35862,N_35061);
or U36809 (N_36809,N_34175,N_35388);
or U36810 (N_36810,N_34312,N_35213);
nor U36811 (N_36811,N_35518,N_34253);
nand U36812 (N_36812,N_34232,N_35913);
or U36813 (N_36813,N_35478,N_34965);
nand U36814 (N_36814,N_35362,N_35091);
or U36815 (N_36815,N_35225,N_35022);
nand U36816 (N_36816,N_35736,N_34844);
nand U36817 (N_36817,N_34219,N_34731);
xor U36818 (N_36818,N_34750,N_35476);
or U36819 (N_36819,N_34806,N_35188);
xor U36820 (N_36820,N_35352,N_34121);
nor U36821 (N_36821,N_35047,N_35652);
or U36822 (N_36822,N_34009,N_34996);
nor U36823 (N_36823,N_35845,N_35375);
or U36824 (N_36824,N_34923,N_34628);
nor U36825 (N_36825,N_34581,N_35155);
nor U36826 (N_36826,N_34452,N_34517);
or U36827 (N_36827,N_34560,N_35977);
nor U36828 (N_36828,N_35911,N_34309);
and U36829 (N_36829,N_34071,N_35096);
and U36830 (N_36830,N_34475,N_35469);
nor U36831 (N_36831,N_34431,N_34477);
and U36832 (N_36832,N_34561,N_35177);
nor U36833 (N_36833,N_34964,N_34909);
xnor U36834 (N_36834,N_35217,N_34055);
or U36835 (N_36835,N_35336,N_35349);
nand U36836 (N_36836,N_35202,N_34746);
nor U36837 (N_36837,N_34863,N_34014);
xor U36838 (N_36838,N_35328,N_35052);
nand U36839 (N_36839,N_34930,N_35865);
nor U36840 (N_36840,N_34614,N_34741);
nor U36841 (N_36841,N_35409,N_34194);
nor U36842 (N_36842,N_35120,N_34664);
xor U36843 (N_36843,N_34073,N_34918);
xnor U36844 (N_36844,N_35141,N_35402);
nand U36845 (N_36845,N_34874,N_35461);
nand U36846 (N_36846,N_34050,N_35430);
nor U36847 (N_36847,N_35682,N_34807);
nand U36848 (N_36848,N_35621,N_35656);
xnor U36849 (N_36849,N_34095,N_34631);
xor U36850 (N_36850,N_34633,N_34471);
nor U36851 (N_36851,N_34767,N_35509);
or U36852 (N_36852,N_35480,N_34085);
or U36853 (N_36853,N_34026,N_34658);
or U36854 (N_36854,N_35614,N_34106);
xor U36855 (N_36855,N_34720,N_34003);
or U36856 (N_36856,N_34192,N_34190);
nand U36857 (N_36857,N_34989,N_35157);
xnor U36858 (N_36858,N_35806,N_34993);
xor U36859 (N_36859,N_34072,N_35390);
nor U36860 (N_36860,N_35418,N_34934);
or U36861 (N_36861,N_34663,N_34262);
nor U36862 (N_36862,N_34956,N_34460);
or U36863 (N_36863,N_35415,N_34444);
and U36864 (N_36864,N_35176,N_35119);
nand U36865 (N_36865,N_34659,N_35836);
and U36866 (N_36866,N_34636,N_35437);
nor U36867 (N_36867,N_34215,N_34789);
xnor U36868 (N_36868,N_35576,N_34368);
nor U36869 (N_36869,N_35383,N_34638);
nor U36870 (N_36870,N_34774,N_34992);
nand U36871 (N_36871,N_34142,N_35558);
and U36872 (N_36872,N_35223,N_35568);
nor U36873 (N_36873,N_35597,N_35615);
nand U36874 (N_36874,N_34656,N_35513);
nor U36875 (N_36875,N_34177,N_34528);
nor U36876 (N_36876,N_35341,N_35424);
nand U36877 (N_36877,N_34670,N_35713);
nand U36878 (N_36878,N_34895,N_35665);
xor U36879 (N_36879,N_35625,N_34722);
nand U36880 (N_36880,N_35938,N_35825);
and U36881 (N_36881,N_34998,N_34775);
or U36882 (N_36882,N_35389,N_34811);
and U36883 (N_36883,N_35018,N_34430);
and U36884 (N_36884,N_34808,N_34402);
nand U36885 (N_36885,N_34541,N_34015);
nor U36886 (N_36886,N_34400,N_34621);
nor U36887 (N_36887,N_35756,N_34613);
or U36888 (N_36888,N_34435,N_34872);
or U36889 (N_36889,N_35972,N_34802);
xnor U36890 (N_36890,N_35396,N_35759);
xnor U36891 (N_36891,N_35316,N_35783);
and U36892 (N_36892,N_34537,N_34290);
or U36893 (N_36893,N_35257,N_34925);
and U36894 (N_36894,N_34274,N_35527);
nor U36895 (N_36895,N_35628,N_34546);
nor U36896 (N_36896,N_35996,N_35374);
xor U36897 (N_36897,N_35672,N_34124);
xnor U36898 (N_36898,N_34258,N_35304);
nor U36899 (N_36899,N_35767,N_34408);
nor U36900 (N_36900,N_35696,N_34547);
nand U36901 (N_36901,N_34269,N_35704);
nand U36902 (N_36902,N_35559,N_34261);
nor U36903 (N_36903,N_35506,N_34481);
nand U36904 (N_36904,N_35310,N_35741);
nor U36905 (N_36905,N_35057,N_34974);
xnor U36906 (N_36906,N_35190,N_35626);
nand U36907 (N_36907,N_34609,N_35569);
nand U36908 (N_36908,N_35053,N_35689);
nand U36909 (N_36909,N_35752,N_34937);
xor U36910 (N_36910,N_34981,N_35215);
nand U36911 (N_36911,N_34819,N_35993);
xor U36912 (N_36912,N_34960,N_34675);
xnor U36913 (N_36913,N_35817,N_35777);
and U36914 (N_36914,N_34456,N_35579);
or U36915 (N_36915,N_35778,N_34044);
and U36916 (N_36916,N_34417,N_35056);
nand U36917 (N_36917,N_35541,N_35343);
or U36918 (N_36918,N_34935,N_34853);
and U36919 (N_36919,N_34251,N_35552);
nor U36920 (N_36920,N_35789,N_34025);
nor U36921 (N_36921,N_35717,N_34623);
nand U36922 (N_36922,N_34833,N_34596);
and U36923 (N_36923,N_34074,N_35964);
xnor U36924 (N_36924,N_34655,N_35780);
or U36925 (N_36925,N_34991,N_35369);
or U36926 (N_36926,N_34346,N_35306);
or U36927 (N_36927,N_35184,N_35113);
or U36928 (N_36928,N_34770,N_35032);
nor U36929 (N_36929,N_35376,N_34168);
nand U36930 (N_36930,N_35127,N_35734);
nand U36931 (N_36931,N_34548,N_35070);
nand U36932 (N_36932,N_35104,N_35973);
nand U36933 (N_36933,N_34975,N_35757);
and U36934 (N_36934,N_35322,N_34390);
nor U36935 (N_36935,N_34531,N_34257);
and U36936 (N_36936,N_34706,N_35076);
nand U36937 (N_36937,N_35697,N_34511);
nor U36938 (N_36938,N_35590,N_34171);
and U36939 (N_36939,N_34207,N_34522);
or U36940 (N_36940,N_35294,N_35994);
nor U36941 (N_36941,N_35681,N_34081);
nand U36942 (N_36942,N_35209,N_34892);
or U36943 (N_36943,N_34379,N_34407);
nor U36944 (N_36944,N_34187,N_35706);
nand U36945 (N_36945,N_35740,N_35485);
nand U36946 (N_36946,N_34729,N_34434);
or U36947 (N_36947,N_34743,N_35027);
nor U36948 (N_36948,N_35851,N_35124);
nand U36949 (N_36949,N_34461,N_34754);
nand U36950 (N_36950,N_35887,N_35677);
nand U36951 (N_36951,N_35537,N_35179);
or U36952 (N_36952,N_35435,N_35995);
xnor U36953 (N_36953,N_34837,N_34320);
or U36954 (N_36954,N_34230,N_34474);
nand U36955 (N_36955,N_34752,N_35493);
and U36956 (N_36956,N_35521,N_34707);
or U36957 (N_36957,N_34618,N_34065);
or U36958 (N_36958,N_34094,N_35610);
or U36959 (N_36959,N_34756,N_34922);
nand U36960 (N_36960,N_34625,N_35432);
nand U36961 (N_36961,N_35895,N_34719);
nor U36962 (N_36962,N_35520,N_35732);
nand U36963 (N_36963,N_34593,N_35655);
or U36964 (N_36964,N_34498,N_35353);
xnor U36965 (N_36965,N_34226,N_34978);
nand U36966 (N_36966,N_34029,N_35261);
or U36967 (N_36967,N_34403,N_34128);
nand U36968 (N_36968,N_35668,N_34076);
or U36969 (N_36969,N_35191,N_34642);
or U36970 (N_36970,N_35255,N_35458);
nor U36971 (N_36971,N_35720,N_35828);
and U36972 (N_36972,N_34389,N_34825);
or U36973 (N_36973,N_35307,N_35816);
nor U36974 (N_36974,N_34110,N_34229);
or U36975 (N_36975,N_34952,N_34123);
nor U36976 (N_36976,N_35024,N_35974);
and U36977 (N_36977,N_34615,N_35725);
nor U36978 (N_36978,N_34272,N_34497);
xor U36979 (N_36979,N_35243,N_34172);
xnor U36980 (N_36980,N_35877,N_34058);
xor U36981 (N_36981,N_35233,N_35201);
xnor U36982 (N_36982,N_35001,N_34112);
nor U36983 (N_36983,N_35416,N_35790);
or U36984 (N_36984,N_34193,N_34958);
or U36985 (N_36985,N_35639,N_34280);
nor U36986 (N_36986,N_34218,N_34385);
xnor U36987 (N_36987,N_34448,N_35531);
or U36988 (N_36988,N_34184,N_35805);
or U36989 (N_36989,N_35483,N_35044);
nand U36990 (N_36990,N_34425,N_35965);
nor U36991 (N_36991,N_35879,N_34372);
nand U36992 (N_36992,N_34887,N_35808);
nor U36993 (N_36993,N_35786,N_34248);
xor U36994 (N_36994,N_34467,N_34834);
and U36995 (N_36995,N_34492,N_34056);
and U36996 (N_36996,N_34711,N_34362);
nand U36997 (N_36997,N_35171,N_34886);
nand U36998 (N_36998,N_34685,N_34469);
or U36999 (N_36999,N_34813,N_35504);
nand U37000 (N_37000,N_35241,N_35002);
and U37001 (N_37001,N_35333,N_34908);
nor U37002 (N_37002,N_34952,N_35491);
and U37003 (N_37003,N_35745,N_34958);
or U37004 (N_37004,N_35620,N_35021);
or U37005 (N_37005,N_34210,N_35490);
and U37006 (N_37006,N_35834,N_35480);
nor U37007 (N_37007,N_35188,N_35577);
nor U37008 (N_37008,N_34911,N_35099);
nand U37009 (N_37009,N_34704,N_34497);
xor U37010 (N_37010,N_35295,N_35814);
and U37011 (N_37011,N_35250,N_34100);
nand U37012 (N_37012,N_35962,N_35271);
and U37013 (N_37013,N_34402,N_34187);
nand U37014 (N_37014,N_34539,N_35881);
nor U37015 (N_37015,N_35227,N_34526);
xor U37016 (N_37016,N_34104,N_34734);
nand U37017 (N_37017,N_34464,N_35127);
and U37018 (N_37018,N_34448,N_35808);
xor U37019 (N_37019,N_34092,N_34892);
and U37020 (N_37020,N_34083,N_34261);
xor U37021 (N_37021,N_34409,N_34664);
nor U37022 (N_37022,N_34601,N_35122);
and U37023 (N_37023,N_34394,N_34738);
xor U37024 (N_37024,N_35440,N_34920);
xnor U37025 (N_37025,N_34115,N_34564);
nand U37026 (N_37026,N_34094,N_35638);
nand U37027 (N_37027,N_34089,N_34546);
or U37028 (N_37028,N_35355,N_34357);
or U37029 (N_37029,N_34593,N_34947);
and U37030 (N_37030,N_35193,N_34274);
xnor U37031 (N_37031,N_35367,N_34327);
nor U37032 (N_37032,N_35138,N_34032);
xnor U37033 (N_37033,N_35452,N_35748);
nor U37034 (N_37034,N_34739,N_34258);
nand U37035 (N_37035,N_34059,N_34259);
nor U37036 (N_37036,N_35305,N_35496);
or U37037 (N_37037,N_34472,N_35114);
xor U37038 (N_37038,N_35168,N_34125);
nor U37039 (N_37039,N_35595,N_35381);
or U37040 (N_37040,N_35760,N_35848);
or U37041 (N_37041,N_35555,N_35290);
nand U37042 (N_37042,N_34315,N_35689);
and U37043 (N_37043,N_34279,N_35511);
and U37044 (N_37044,N_34404,N_35815);
and U37045 (N_37045,N_35155,N_35360);
xnor U37046 (N_37046,N_35832,N_35337);
and U37047 (N_37047,N_34040,N_35700);
and U37048 (N_37048,N_35143,N_35396);
or U37049 (N_37049,N_35698,N_34246);
and U37050 (N_37050,N_34564,N_34729);
and U37051 (N_37051,N_34766,N_35161);
nor U37052 (N_37052,N_34071,N_35015);
nor U37053 (N_37053,N_35020,N_35280);
xnor U37054 (N_37054,N_35353,N_34542);
or U37055 (N_37055,N_34699,N_34078);
nor U37056 (N_37056,N_35993,N_34577);
nand U37057 (N_37057,N_35196,N_34827);
nor U37058 (N_37058,N_35008,N_35661);
nor U37059 (N_37059,N_35035,N_34702);
and U37060 (N_37060,N_35839,N_34715);
or U37061 (N_37061,N_34233,N_35979);
or U37062 (N_37062,N_34001,N_34774);
xor U37063 (N_37063,N_34623,N_35812);
xor U37064 (N_37064,N_35197,N_35579);
xnor U37065 (N_37065,N_34466,N_35464);
xnor U37066 (N_37066,N_34200,N_34778);
nand U37067 (N_37067,N_35556,N_34359);
and U37068 (N_37068,N_35538,N_35536);
nand U37069 (N_37069,N_34217,N_35279);
and U37070 (N_37070,N_34511,N_35724);
or U37071 (N_37071,N_35962,N_35872);
xor U37072 (N_37072,N_35420,N_35773);
nor U37073 (N_37073,N_35702,N_34287);
xor U37074 (N_37074,N_34115,N_34837);
nand U37075 (N_37075,N_34397,N_34175);
nor U37076 (N_37076,N_34395,N_35915);
or U37077 (N_37077,N_34122,N_35333);
nand U37078 (N_37078,N_34860,N_35297);
or U37079 (N_37079,N_34221,N_35774);
and U37080 (N_37080,N_34717,N_34870);
nand U37081 (N_37081,N_34989,N_34012);
and U37082 (N_37082,N_35521,N_34733);
and U37083 (N_37083,N_35888,N_34216);
and U37084 (N_37084,N_34399,N_34905);
or U37085 (N_37085,N_35704,N_35516);
nand U37086 (N_37086,N_34849,N_34556);
nand U37087 (N_37087,N_35165,N_35784);
nor U37088 (N_37088,N_34095,N_35692);
or U37089 (N_37089,N_35864,N_34779);
xor U37090 (N_37090,N_35591,N_34324);
nand U37091 (N_37091,N_35713,N_35041);
nor U37092 (N_37092,N_34522,N_34945);
nand U37093 (N_37093,N_34914,N_35825);
nor U37094 (N_37094,N_35225,N_35911);
nand U37095 (N_37095,N_35197,N_34612);
xor U37096 (N_37096,N_35720,N_35785);
nor U37097 (N_37097,N_34089,N_35128);
xor U37098 (N_37098,N_35528,N_35422);
nor U37099 (N_37099,N_35880,N_35295);
nor U37100 (N_37100,N_34905,N_35976);
nor U37101 (N_37101,N_34794,N_34198);
nand U37102 (N_37102,N_35544,N_35674);
nand U37103 (N_37103,N_34488,N_34593);
xor U37104 (N_37104,N_34807,N_34193);
or U37105 (N_37105,N_34899,N_34125);
nor U37106 (N_37106,N_35318,N_34941);
xnor U37107 (N_37107,N_35817,N_34640);
or U37108 (N_37108,N_34100,N_35321);
xnor U37109 (N_37109,N_34424,N_34310);
nand U37110 (N_37110,N_34946,N_35343);
nor U37111 (N_37111,N_35885,N_35953);
nor U37112 (N_37112,N_34698,N_35303);
nor U37113 (N_37113,N_35164,N_35632);
nor U37114 (N_37114,N_35376,N_34267);
nor U37115 (N_37115,N_34313,N_34723);
or U37116 (N_37116,N_34165,N_34945);
xor U37117 (N_37117,N_35692,N_35781);
nand U37118 (N_37118,N_35923,N_35914);
or U37119 (N_37119,N_35605,N_35373);
and U37120 (N_37120,N_34894,N_35382);
and U37121 (N_37121,N_35076,N_35665);
nand U37122 (N_37122,N_34894,N_34376);
nor U37123 (N_37123,N_34910,N_35566);
or U37124 (N_37124,N_35385,N_34009);
xor U37125 (N_37125,N_34609,N_34128);
or U37126 (N_37126,N_35596,N_35077);
and U37127 (N_37127,N_34320,N_35625);
nand U37128 (N_37128,N_34495,N_35244);
xnor U37129 (N_37129,N_35816,N_35498);
or U37130 (N_37130,N_35938,N_34792);
and U37131 (N_37131,N_35437,N_35418);
or U37132 (N_37132,N_35918,N_34357);
xnor U37133 (N_37133,N_35768,N_34505);
and U37134 (N_37134,N_35504,N_35180);
xnor U37135 (N_37135,N_34769,N_34261);
nand U37136 (N_37136,N_34801,N_35592);
nor U37137 (N_37137,N_34523,N_35646);
nand U37138 (N_37138,N_35305,N_34095);
nor U37139 (N_37139,N_34694,N_35505);
and U37140 (N_37140,N_34683,N_35546);
nand U37141 (N_37141,N_34994,N_34849);
nand U37142 (N_37142,N_35812,N_34011);
or U37143 (N_37143,N_34069,N_34347);
xor U37144 (N_37144,N_35180,N_35967);
nor U37145 (N_37145,N_35822,N_34434);
or U37146 (N_37146,N_34143,N_34024);
and U37147 (N_37147,N_34156,N_35371);
and U37148 (N_37148,N_35868,N_35907);
nor U37149 (N_37149,N_34067,N_34382);
or U37150 (N_37150,N_35305,N_34004);
nor U37151 (N_37151,N_35469,N_35626);
and U37152 (N_37152,N_35055,N_35641);
and U37153 (N_37153,N_34921,N_34603);
nand U37154 (N_37154,N_34553,N_34373);
nand U37155 (N_37155,N_34057,N_34423);
nand U37156 (N_37156,N_35748,N_35658);
and U37157 (N_37157,N_34423,N_35873);
xnor U37158 (N_37158,N_34225,N_35609);
or U37159 (N_37159,N_35386,N_34891);
nor U37160 (N_37160,N_35680,N_34911);
or U37161 (N_37161,N_34717,N_34261);
or U37162 (N_37162,N_35397,N_34842);
and U37163 (N_37163,N_35758,N_34887);
nand U37164 (N_37164,N_34256,N_34643);
nand U37165 (N_37165,N_34533,N_34251);
or U37166 (N_37166,N_35534,N_35643);
nand U37167 (N_37167,N_35580,N_35138);
and U37168 (N_37168,N_35362,N_35278);
and U37169 (N_37169,N_34127,N_35258);
xor U37170 (N_37170,N_35322,N_35383);
and U37171 (N_37171,N_34401,N_34719);
nor U37172 (N_37172,N_35319,N_34838);
and U37173 (N_37173,N_35113,N_34463);
nand U37174 (N_37174,N_35699,N_35082);
nand U37175 (N_37175,N_34935,N_35627);
nor U37176 (N_37176,N_35629,N_34011);
and U37177 (N_37177,N_34487,N_35632);
nor U37178 (N_37178,N_35241,N_35009);
nor U37179 (N_37179,N_35396,N_35359);
nand U37180 (N_37180,N_34836,N_35880);
xor U37181 (N_37181,N_35450,N_35205);
or U37182 (N_37182,N_35871,N_34435);
nor U37183 (N_37183,N_35613,N_35735);
or U37184 (N_37184,N_34637,N_35229);
and U37185 (N_37185,N_35777,N_35932);
nand U37186 (N_37186,N_35769,N_34720);
or U37187 (N_37187,N_35760,N_34830);
nor U37188 (N_37188,N_35399,N_34488);
or U37189 (N_37189,N_35775,N_34649);
nor U37190 (N_37190,N_35427,N_35979);
or U37191 (N_37191,N_35442,N_34195);
and U37192 (N_37192,N_34264,N_35197);
and U37193 (N_37193,N_34311,N_35518);
or U37194 (N_37194,N_34430,N_35574);
xnor U37195 (N_37195,N_34480,N_34861);
nand U37196 (N_37196,N_34978,N_34802);
or U37197 (N_37197,N_34849,N_35056);
nand U37198 (N_37198,N_35367,N_35527);
xor U37199 (N_37199,N_35104,N_34448);
or U37200 (N_37200,N_35176,N_35089);
and U37201 (N_37201,N_35884,N_35816);
and U37202 (N_37202,N_35195,N_34367);
nor U37203 (N_37203,N_34130,N_34205);
xnor U37204 (N_37204,N_35200,N_34459);
nand U37205 (N_37205,N_35305,N_35058);
and U37206 (N_37206,N_35145,N_34631);
nor U37207 (N_37207,N_35686,N_34908);
xnor U37208 (N_37208,N_34695,N_35948);
and U37209 (N_37209,N_35115,N_35579);
or U37210 (N_37210,N_35934,N_34487);
nand U37211 (N_37211,N_34325,N_35678);
nor U37212 (N_37212,N_35902,N_34984);
xor U37213 (N_37213,N_34924,N_35200);
or U37214 (N_37214,N_35614,N_34581);
xor U37215 (N_37215,N_34338,N_34635);
nor U37216 (N_37216,N_35224,N_35867);
xnor U37217 (N_37217,N_35984,N_35321);
and U37218 (N_37218,N_34955,N_34235);
nand U37219 (N_37219,N_34044,N_35239);
nor U37220 (N_37220,N_34695,N_35499);
nand U37221 (N_37221,N_34168,N_35422);
nor U37222 (N_37222,N_35346,N_35771);
or U37223 (N_37223,N_34546,N_34651);
or U37224 (N_37224,N_34592,N_35284);
or U37225 (N_37225,N_34888,N_35282);
and U37226 (N_37226,N_34158,N_34885);
xnor U37227 (N_37227,N_34776,N_34380);
nand U37228 (N_37228,N_35965,N_34154);
xnor U37229 (N_37229,N_34793,N_34136);
or U37230 (N_37230,N_35930,N_35749);
xnor U37231 (N_37231,N_34890,N_35124);
or U37232 (N_37232,N_35590,N_34455);
xnor U37233 (N_37233,N_35339,N_35730);
nand U37234 (N_37234,N_34605,N_34714);
or U37235 (N_37235,N_34297,N_35236);
xnor U37236 (N_37236,N_35146,N_34032);
xnor U37237 (N_37237,N_34759,N_35942);
or U37238 (N_37238,N_34352,N_34849);
nor U37239 (N_37239,N_35538,N_34961);
nand U37240 (N_37240,N_34697,N_35478);
or U37241 (N_37241,N_35583,N_35420);
and U37242 (N_37242,N_35129,N_34689);
nor U37243 (N_37243,N_34804,N_35158);
and U37244 (N_37244,N_35902,N_34442);
nor U37245 (N_37245,N_34740,N_34799);
nor U37246 (N_37246,N_35844,N_35849);
xor U37247 (N_37247,N_35392,N_35612);
nor U37248 (N_37248,N_34866,N_35089);
xnor U37249 (N_37249,N_35768,N_35477);
or U37250 (N_37250,N_34037,N_34382);
or U37251 (N_37251,N_35036,N_35613);
or U37252 (N_37252,N_34317,N_35550);
nor U37253 (N_37253,N_34908,N_34733);
xor U37254 (N_37254,N_34131,N_35199);
nand U37255 (N_37255,N_34226,N_34332);
or U37256 (N_37256,N_35486,N_35115);
nand U37257 (N_37257,N_35909,N_34002);
or U37258 (N_37258,N_35558,N_34368);
or U37259 (N_37259,N_35727,N_34164);
or U37260 (N_37260,N_35283,N_34952);
and U37261 (N_37261,N_34950,N_35449);
xor U37262 (N_37262,N_35407,N_34207);
or U37263 (N_37263,N_34949,N_35356);
or U37264 (N_37264,N_35354,N_34973);
or U37265 (N_37265,N_34220,N_35113);
and U37266 (N_37266,N_35836,N_34277);
nand U37267 (N_37267,N_35716,N_34405);
nand U37268 (N_37268,N_34698,N_35314);
or U37269 (N_37269,N_34866,N_34195);
or U37270 (N_37270,N_35699,N_34772);
xor U37271 (N_37271,N_34109,N_35490);
nand U37272 (N_37272,N_34019,N_34425);
xnor U37273 (N_37273,N_35492,N_35085);
xnor U37274 (N_37274,N_34443,N_34253);
or U37275 (N_37275,N_34388,N_35889);
nor U37276 (N_37276,N_35348,N_34774);
nor U37277 (N_37277,N_35033,N_34565);
nand U37278 (N_37278,N_34895,N_34152);
nand U37279 (N_37279,N_34123,N_34106);
xnor U37280 (N_37280,N_35913,N_35232);
nor U37281 (N_37281,N_34406,N_34704);
and U37282 (N_37282,N_35967,N_35086);
and U37283 (N_37283,N_34774,N_34762);
and U37284 (N_37284,N_34071,N_34029);
xnor U37285 (N_37285,N_35280,N_34300);
and U37286 (N_37286,N_35862,N_34143);
or U37287 (N_37287,N_35510,N_34626);
and U37288 (N_37288,N_35911,N_34754);
nor U37289 (N_37289,N_34774,N_35774);
or U37290 (N_37290,N_34516,N_35533);
nand U37291 (N_37291,N_35544,N_35098);
and U37292 (N_37292,N_35252,N_34973);
and U37293 (N_37293,N_34126,N_34514);
nor U37294 (N_37294,N_35739,N_34410);
and U37295 (N_37295,N_34195,N_35614);
nand U37296 (N_37296,N_34026,N_34219);
nor U37297 (N_37297,N_34401,N_34510);
nand U37298 (N_37298,N_34095,N_34206);
or U37299 (N_37299,N_34504,N_34426);
nand U37300 (N_37300,N_34189,N_35284);
or U37301 (N_37301,N_34342,N_35007);
nor U37302 (N_37302,N_35217,N_35168);
and U37303 (N_37303,N_34736,N_34669);
and U37304 (N_37304,N_35319,N_35100);
nand U37305 (N_37305,N_34751,N_34674);
nand U37306 (N_37306,N_35031,N_34396);
or U37307 (N_37307,N_35989,N_34193);
nor U37308 (N_37308,N_34481,N_35994);
nand U37309 (N_37309,N_34091,N_34157);
and U37310 (N_37310,N_35629,N_35464);
nor U37311 (N_37311,N_34776,N_35167);
and U37312 (N_37312,N_35011,N_34135);
nor U37313 (N_37313,N_34694,N_35914);
or U37314 (N_37314,N_34281,N_35033);
or U37315 (N_37315,N_34859,N_35163);
and U37316 (N_37316,N_34262,N_34782);
nor U37317 (N_37317,N_34991,N_35014);
nor U37318 (N_37318,N_34469,N_34561);
or U37319 (N_37319,N_35167,N_35592);
nor U37320 (N_37320,N_35537,N_35167);
nor U37321 (N_37321,N_35865,N_34081);
nor U37322 (N_37322,N_34590,N_34446);
nor U37323 (N_37323,N_34393,N_34773);
nand U37324 (N_37324,N_34824,N_35609);
or U37325 (N_37325,N_35303,N_34653);
nor U37326 (N_37326,N_35509,N_35217);
nor U37327 (N_37327,N_35938,N_34192);
or U37328 (N_37328,N_35970,N_35317);
xnor U37329 (N_37329,N_35535,N_35457);
nor U37330 (N_37330,N_34300,N_34120);
or U37331 (N_37331,N_35317,N_35002);
nand U37332 (N_37332,N_35295,N_35305);
or U37333 (N_37333,N_34684,N_35903);
or U37334 (N_37334,N_35038,N_34512);
and U37335 (N_37335,N_34150,N_34338);
or U37336 (N_37336,N_35533,N_34339);
or U37337 (N_37337,N_35366,N_35382);
xor U37338 (N_37338,N_34266,N_34047);
and U37339 (N_37339,N_34922,N_35247);
or U37340 (N_37340,N_35938,N_35738);
and U37341 (N_37341,N_34644,N_34459);
xor U37342 (N_37342,N_34438,N_35723);
nand U37343 (N_37343,N_34008,N_34953);
or U37344 (N_37344,N_34267,N_34320);
nor U37345 (N_37345,N_34495,N_35979);
nand U37346 (N_37346,N_35941,N_34021);
xnor U37347 (N_37347,N_34993,N_34811);
or U37348 (N_37348,N_35415,N_35953);
or U37349 (N_37349,N_35997,N_34794);
or U37350 (N_37350,N_34338,N_34233);
nand U37351 (N_37351,N_35014,N_35987);
xnor U37352 (N_37352,N_34135,N_35047);
or U37353 (N_37353,N_34136,N_35825);
nor U37354 (N_37354,N_35920,N_35755);
or U37355 (N_37355,N_35126,N_34061);
nand U37356 (N_37356,N_34153,N_35194);
xnor U37357 (N_37357,N_35306,N_35617);
xor U37358 (N_37358,N_34524,N_35294);
xnor U37359 (N_37359,N_34705,N_35516);
nand U37360 (N_37360,N_35058,N_35876);
nor U37361 (N_37361,N_34124,N_34053);
or U37362 (N_37362,N_35172,N_35731);
or U37363 (N_37363,N_34454,N_35453);
nand U37364 (N_37364,N_34506,N_35855);
nor U37365 (N_37365,N_34495,N_34002);
nand U37366 (N_37366,N_35494,N_35163);
nand U37367 (N_37367,N_35072,N_34786);
and U37368 (N_37368,N_34710,N_34449);
nor U37369 (N_37369,N_34244,N_35767);
nor U37370 (N_37370,N_35555,N_34215);
nor U37371 (N_37371,N_34111,N_34893);
nand U37372 (N_37372,N_35163,N_35129);
nor U37373 (N_37373,N_35124,N_35167);
or U37374 (N_37374,N_34867,N_35446);
nand U37375 (N_37375,N_35282,N_34310);
nor U37376 (N_37376,N_34603,N_34301);
or U37377 (N_37377,N_35683,N_34129);
nand U37378 (N_37378,N_34847,N_35448);
nor U37379 (N_37379,N_35158,N_35508);
nand U37380 (N_37380,N_34183,N_35307);
nand U37381 (N_37381,N_34837,N_35612);
nor U37382 (N_37382,N_34168,N_34906);
and U37383 (N_37383,N_35384,N_34408);
xnor U37384 (N_37384,N_35154,N_35580);
and U37385 (N_37385,N_34659,N_35533);
xor U37386 (N_37386,N_35677,N_35917);
nor U37387 (N_37387,N_35327,N_35564);
and U37388 (N_37388,N_35393,N_34865);
or U37389 (N_37389,N_35821,N_35532);
nor U37390 (N_37390,N_35060,N_35303);
or U37391 (N_37391,N_34882,N_35004);
nor U37392 (N_37392,N_35562,N_35333);
or U37393 (N_37393,N_35481,N_35486);
or U37394 (N_37394,N_34831,N_34218);
or U37395 (N_37395,N_34274,N_35337);
nand U37396 (N_37396,N_35482,N_34753);
and U37397 (N_37397,N_35429,N_35510);
nand U37398 (N_37398,N_35782,N_35394);
nor U37399 (N_37399,N_35152,N_35254);
nand U37400 (N_37400,N_34752,N_35690);
nor U37401 (N_37401,N_35933,N_35395);
nand U37402 (N_37402,N_34815,N_35704);
nand U37403 (N_37403,N_35273,N_34969);
or U37404 (N_37404,N_35096,N_34024);
or U37405 (N_37405,N_34818,N_34038);
or U37406 (N_37406,N_35111,N_34203);
or U37407 (N_37407,N_34873,N_35713);
or U37408 (N_37408,N_35170,N_35648);
nand U37409 (N_37409,N_34100,N_34509);
nand U37410 (N_37410,N_35688,N_34032);
xnor U37411 (N_37411,N_35167,N_35438);
or U37412 (N_37412,N_34170,N_35129);
and U37413 (N_37413,N_34326,N_35587);
nor U37414 (N_37414,N_34288,N_35062);
or U37415 (N_37415,N_34055,N_35323);
xnor U37416 (N_37416,N_35065,N_35824);
nand U37417 (N_37417,N_35021,N_35759);
nand U37418 (N_37418,N_34087,N_35174);
and U37419 (N_37419,N_35885,N_34533);
or U37420 (N_37420,N_34507,N_35595);
xnor U37421 (N_37421,N_34659,N_34842);
nand U37422 (N_37422,N_35779,N_34955);
or U37423 (N_37423,N_34559,N_35383);
nand U37424 (N_37424,N_34995,N_35165);
nor U37425 (N_37425,N_34828,N_35622);
xor U37426 (N_37426,N_35656,N_35821);
nand U37427 (N_37427,N_35189,N_34437);
nor U37428 (N_37428,N_35916,N_34435);
and U37429 (N_37429,N_34119,N_35985);
xor U37430 (N_37430,N_35353,N_34977);
xor U37431 (N_37431,N_35864,N_35481);
nand U37432 (N_37432,N_34167,N_34719);
nor U37433 (N_37433,N_34467,N_35769);
and U37434 (N_37434,N_35660,N_34328);
xor U37435 (N_37435,N_35810,N_34563);
nor U37436 (N_37436,N_34880,N_35100);
nand U37437 (N_37437,N_35056,N_35289);
nor U37438 (N_37438,N_34427,N_35419);
nor U37439 (N_37439,N_34674,N_35933);
nor U37440 (N_37440,N_35274,N_35335);
nor U37441 (N_37441,N_34528,N_35333);
or U37442 (N_37442,N_35429,N_34347);
or U37443 (N_37443,N_35160,N_35147);
and U37444 (N_37444,N_34116,N_35469);
xnor U37445 (N_37445,N_35886,N_34298);
or U37446 (N_37446,N_34158,N_35564);
and U37447 (N_37447,N_35212,N_35131);
nand U37448 (N_37448,N_35850,N_35486);
and U37449 (N_37449,N_34219,N_34344);
and U37450 (N_37450,N_35232,N_34730);
nor U37451 (N_37451,N_34012,N_34026);
nor U37452 (N_37452,N_34305,N_35498);
and U37453 (N_37453,N_34994,N_35194);
xnor U37454 (N_37454,N_35234,N_35060);
nand U37455 (N_37455,N_35183,N_34068);
or U37456 (N_37456,N_35374,N_34279);
or U37457 (N_37457,N_35513,N_34933);
nand U37458 (N_37458,N_34796,N_34224);
or U37459 (N_37459,N_35437,N_34061);
nor U37460 (N_37460,N_35093,N_34510);
and U37461 (N_37461,N_34055,N_35874);
xnor U37462 (N_37462,N_34814,N_35311);
nand U37463 (N_37463,N_34081,N_35201);
nor U37464 (N_37464,N_35132,N_34055);
and U37465 (N_37465,N_35757,N_35289);
and U37466 (N_37466,N_35877,N_34875);
nand U37467 (N_37467,N_35963,N_34733);
nor U37468 (N_37468,N_35847,N_35432);
xnor U37469 (N_37469,N_34114,N_34078);
nand U37470 (N_37470,N_35803,N_34192);
or U37471 (N_37471,N_35566,N_34811);
xnor U37472 (N_37472,N_35100,N_35396);
nand U37473 (N_37473,N_35372,N_34172);
nor U37474 (N_37474,N_35473,N_35668);
or U37475 (N_37475,N_34589,N_35819);
nand U37476 (N_37476,N_34427,N_34753);
or U37477 (N_37477,N_34981,N_35434);
or U37478 (N_37478,N_34372,N_34719);
or U37479 (N_37479,N_34468,N_35273);
or U37480 (N_37480,N_34871,N_34226);
xor U37481 (N_37481,N_35959,N_34942);
or U37482 (N_37482,N_34386,N_34088);
or U37483 (N_37483,N_35944,N_34519);
nor U37484 (N_37484,N_34624,N_34587);
nor U37485 (N_37485,N_34066,N_35033);
or U37486 (N_37486,N_34402,N_34182);
and U37487 (N_37487,N_35015,N_34752);
nor U37488 (N_37488,N_34693,N_34695);
nor U37489 (N_37489,N_34934,N_34125);
xor U37490 (N_37490,N_35085,N_35099);
nand U37491 (N_37491,N_35254,N_34721);
xnor U37492 (N_37492,N_35879,N_35464);
and U37493 (N_37493,N_34096,N_35100);
and U37494 (N_37494,N_35710,N_35193);
and U37495 (N_37495,N_34067,N_34834);
xor U37496 (N_37496,N_35079,N_35518);
or U37497 (N_37497,N_34660,N_35184);
or U37498 (N_37498,N_35352,N_34594);
nand U37499 (N_37499,N_34192,N_35220);
and U37500 (N_37500,N_35151,N_35323);
nand U37501 (N_37501,N_34323,N_35032);
xor U37502 (N_37502,N_35527,N_34376);
or U37503 (N_37503,N_35992,N_35654);
nand U37504 (N_37504,N_35752,N_34214);
nor U37505 (N_37505,N_34129,N_34903);
xor U37506 (N_37506,N_35567,N_34627);
xnor U37507 (N_37507,N_34369,N_34358);
or U37508 (N_37508,N_35455,N_34355);
or U37509 (N_37509,N_34187,N_35955);
or U37510 (N_37510,N_34408,N_35688);
nor U37511 (N_37511,N_34794,N_35639);
xor U37512 (N_37512,N_34352,N_34205);
nand U37513 (N_37513,N_35292,N_34143);
xor U37514 (N_37514,N_34087,N_34768);
or U37515 (N_37515,N_34746,N_35572);
or U37516 (N_37516,N_35783,N_34562);
xor U37517 (N_37517,N_34201,N_34332);
nor U37518 (N_37518,N_34599,N_34049);
nor U37519 (N_37519,N_35452,N_35322);
nor U37520 (N_37520,N_35353,N_34577);
nand U37521 (N_37521,N_34493,N_34736);
or U37522 (N_37522,N_34542,N_34423);
and U37523 (N_37523,N_35832,N_35107);
and U37524 (N_37524,N_34140,N_35090);
nand U37525 (N_37525,N_35372,N_35108);
and U37526 (N_37526,N_34020,N_35311);
nand U37527 (N_37527,N_35478,N_34926);
nor U37528 (N_37528,N_35093,N_35088);
nor U37529 (N_37529,N_35548,N_35446);
and U37530 (N_37530,N_34181,N_35112);
or U37531 (N_37531,N_34256,N_34271);
nor U37532 (N_37532,N_34060,N_35454);
nand U37533 (N_37533,N_35160,N_35687);
xnor U37534 (N_37534,N_35607,N_34429);
nor U37535 (N_37535,N_34394,N_35614);
and U37536 (N_37536,N_35357,N_34651);
nand U37537 (N_37537,N_35032,N_35829);
and U37538 (N_37538,N_35518,N_34875);
nor U37539 (N_37539,N_35971,N_34170);
nor U37540 (N_37540,N_35181,N_35445);
or U37541 (N_37541,N_34752,N_35280);
nand U37542 (N_37542,N_34997,N_35692);
xor U37543 (N_37543,N_35268,N_35416);
and U37544 (N_37544,N_35428,N_34748);
and U37545 (N_37545,N_35522,N_35994);
xor U37546 (N_37546,N_34601,N_34309);
or U37547 (N_37547,N_35675,N_35917);
nor U37548 (N_37548,N_34251,N_34371);
nand U37549 (N_37549,N_34962,N_35594);
or U37550 (N_37550,N_35233,N_34096);
nor U37551 (N_37551,N_35074,N_35406);
nand U37552 (N_37552,N_34933,N_35609);
nand U37553 (N_37553,N_34065,N_34505);
xor U37554 (N_37554,N_34278,N_34379);
nand U37555 (N_37555,N_35215,N_34114);
xor U37556 (N_37556,N_34803,N_34875);
and U37557 (N_37557,N_35388,N_34955);
nand U37558 (N_37558,N_34092,N_35499);
nor U37559 (N_37559,N_35318,N_34721);
and U37560 (N_37560,N_34525,N_34119);
xor U37561 (N_37561,N_34095,N_34401);
nand U37562 (N_37562,N_34108,N_35855);
or U37563 (N_37563,N_35591,N_35750);
nor U37564 (N_37564,N_34414,N_34422);
xnor U37565 (N_37565,N_34433,N_34447);
nand U37566 (N_37566,N_35888,N_35729);
nor U37567 (N_37567,N_34195,N_34969);
or U37568 (N_37568,N_34841,N_35960);
nor U37569 (N_37569,N_35056,N_34040);
nor U37570 (N_37570,N_35552,N_34619);
nand U37571 (N_37571,N_35812,N_34424);
nand U37572 (N_37572,N_35369,N_34216);
or U37573 (N_37573,N_35433,N_35212);
nor U37574 (N_37574,N_34864,N_35541);
nand U37575 (N_37575,N_34286,N_34215);
nand U37576 (N_37576,N_35307,N_34883);
xor U37577 (N_37577,N_35289,N_34586);
or U37578 (N_37578,N_35468,N_35806);
nand U37579 (N_37579,N_35059,N_34046);
nor U37580 (N_37580,N_35776,N_34544);
and U37581 (N_37581,N_35329,N_35084);
and U37582 (N_37582,N_35760,N_34599);
or U37583 (N_37583,N_34950,N_34263);
and U37584 (N_37584,N_35452,N_35589);
and U37585 (N_37585,N_34295,N_34617);
xnor U37586 (N_37586,N_35818,N_35644);
nand U37587 (N_37587,N_35288,N_34051);
nor U37588 (N_37588,N_34781,N_35981);
nor U37589 (N_37589,N_35946,N_35165);
xor U37590 (N_37590,N_35725,N_34834);
nand U37591 (N_37591,N_35474,N_34024);
nand U37592 (N_37592,N_35003,N_34288);
and U37593 (N_37593,N_35823,N_35848);
nand U37594 (N_37594,N_34882,N_35301);
xor U37595 (N_37595,N_35674,N_34571);
xor U37596 (N_37596,N_34094,N_34007);
or U37597 (N_37597,N_34427,N_34990);
or U37598 (N_37598,N_34992,N_35526);
nand U37599 (N_37599,N_34856,N_34825);
nand U37600 (N_37600,N_34589,N_34536);
and U37601 (N_37601,N_34644,N_35562);
and U37602 (N_37602,N_34287,N_34482);
nor U37603 (N_37603,N_34927,N_34579);
xnor U37604 (N_37604,N_34626,N_34705);
or U37605 (N_37605,N_34909,N_34444);
and U37606 (N_37606,N_34235,N_34214);
and U37607 (N_37607,N_34130,N_35624);
xnor U37608 (N_37608,N_35903,N_35260);
or U37609 (N_37609,N_35623,N_35105);
xnor U37610 (N_37610,N_35490,N_34158);
or U37611 (N_37611,N_35714,N_34573);
nand U37612 (N_37612,N_34048,N_34412);
nor U37613 (N_37613,N_35454,N_34182);
xnor U37614 (N_37614,N_35915,N_35548);
xnor U37615 (N_37615,N_35848,N_34962);
nor U37616 (N_37616,N_35093,N_35044);
nor U37617 (N_37617,N_35126,N_35036);
nor U37618 (N_37618,N_35521,N_34187);
xor U37619 (N_37619,N_35648,N_34277);
or U37620 (N_37620,N_34142,N_35594);
nand U37621 (N_37621,N_35476,N_34537);
and U37622 (N_37622,N_35402,N_35031);
and U37623 (N_37623,N_35088,N_34576);
or U37624 (N_37624,N_35388,N_34537);
nor U37625 (N_37625,N_34253,N_34884);
nand U37626 (N_37626,N_34021,N_34308);
xor U37627 (N_37627,N_35195,N_34920);
nor U37628 (N_37628,N_34618,N_35913);
or U37629 (N_37629,N_34037,N_34413);
nand U37630 (N_37630,N_35566,N_35260);
nor U37631 (N_37631,N_35704,N_34972);
nor U37632 (N_37632,N_35140,N_35370);
or U37633 (N_37633,N_35878,N_35835);
nand U37634 (N_37634,N_34904,N_34736);
and U37635 (N_37635,N_34260,N_35865);
xnor U37636 (N_37636,N_34930,N_34959);
xnor U37637 (N_37637,N_35126,N_35474);
nand U37638 (N_37638,N_34132,N_34399);
or U37639 (N_37639,N_35027,N_35627);
nor U37640 (N_37640,N_35027,N_35638);
or U37641 (N_37641,N_35073,N_34491);
nor U37642 (N_37642,N_34702,N_35846);
or U37643 (N_37643,N_35343,N_35680);
and U37644 (N_37644,N_35142,N_34925);
nand U37645 (N_37645,N_34301,N_35861);
xor U37646 (N_37646,N_35593,N_35482);
nand U37647 (N_37647,N_34575,N_34358);
or U37648 (N_37648,N_35021,N_35326);
and U37649 (N_37649,N_34596,N_35461);
nor U37650 (N_37650,N_35018,N_34481);
xor U37651 (N_37651,N_35630,N_35328);
xor U37652 (N_37652,N_35443,N_35145);
and U37653 (N_37653,N_35299,N_34817);
nor U37654 (N_37654,N_35458,N_35581);
nand U37655 (N_37655,N_34114,N_34813);
nand U37656 (N_37656,N_35150,N_34627);
nor U37657 (N_37657,N_34286,N_34757);
and U37658 (N_37658,N_34630,N_35259);
and U37659 (N_37659,N_34989,N_34519);
and U37660 (N_37660,N_34853,N_35550);
xnor U37661 (N_37661,N_34779,N_34827);
xor U37662 (N_37662,N_34670,N_35394);
nor U37663 (N_37663,N_34159,N_35857);
xor U37664 (N_37664,N_34579,N_35109);
xnor U37665 (N_37665,N_34238,N_35032);
and U37666 (N_37666,N_35518,N_34959);
xor U37667 (N_37667,N_35096,N_34446);
xor U37668 (N_37668,N_34265,N_34429);
or U37669 (N_37669,N_35655,N_35091);
or U37670 (N_37670,N_35697,N_34793);
or U37671 (N_37671,N_35451,N_35648);
xnor U37672 (N_37672,N_34256,N_35963);
nand U37673 (N_37673,N_35138,N_35783);
xnor U37674 (N_37674,N_34040,N_35072);
nand U37675 (N_37675,N_34920,N_35050);
nand U37676 (N_37676,N_35218,N_34728);
and U37677 (N_37677,N_34222,N_34293);
nor U37678 (N_37678,N_35350,N_34794);
nand U37679 (N_37679,N_35767,N_35017);
and U37680 (N_37680,N_35159,N_35987);
xnor U37681 (N_37681,N_35335,N_35088);
and U37682 (N_37682,N_35522,N_34350);
nor U37683 (N_37683,N_35473,N_34107);
or U37684 (N_37684,N_35458,N_34066);
or U37685 (N_37685,N_35066,N_35510);
and U37686 (N_37686,N_34178,N_35594);
xnor U37687 (N_37687,N_35719,N_35433);
nand U37688 (N_37688,N_34818,N_34797);
and U37689 (N_37689,N_34927,N_34522);
nor U37690 (N_37690,N_35086,N_35325);
nor U37691 (N_37691,N_35255,N_35147);
or U37692 (N_37692,N_34153,N_35596);
or U37693 (N_37693,N_34517,N_35306);
nor U37694 (N_37694,N_34732,N_35218);
and U37695 (N_37695,N_35245,N_34095);
nand U37696 (N_37696,N_34641,N_34254);
or U37697 (N_37697,N_34108,N_34674);
and U37698 (N_37698,N_34587,N_35489);
xor U37699 (N_37699,N_35484,N_35548);
nand U37700 (N_37700,N_35366,N_34960);
and U37701 (N_37701,N_34427,N_35933);
nand U37702 (N_37702,N_35214,N_35561);
or U37703 (N_37703,N_34493,N_35507);
xnor U37704 (N_37704,N_34521,N_34948);
xnor U37705 (N_37705,N_34404,N_35112);
nand U37706 (N_37706,N_34699,N_34532);
nor U37707 (N_37707,N_35662,N_35886);
or U37708 (N_37708,N_34247,N_35645);
or U37709 (N_37709,N_35867,N_35194);
or U37710 (N_37710,N_34434,N_34303);
or U37711 (N_37711,N_35080,N_34967);
and U37712 (N_37712,N_34273,N_34758);
nor U37713 (N_37713,N_35393,N_35760);
and U37714 (N_37714,N_34143,N_34426);
or U37715 (N_37715,N_35927,N_34878);
or U37716 (N_37716,N_35050,N_34291);
and U37717 (N_37717,N_35890,N_34989);
and U37718 (N_37718,N_35178,N_34688);
or U37719 (N_37719,N_35695,N_35330);
nand U37720 (N_37720,N_34842,N_34347);
xnor U37721 (N_37721,N_34413,N_34618);
nand U37722 (N_37722,N_34842,N_34162);
nor U37723 (N_37723,N_35104,N_35561);
nor U37724 (N_37724,N_34790,N_34134);
or U37725 (N_37725,N_34864,N_34865);
and U37726 (N_37726,N_35226,N_35787);
or U37727 (N_37727,N_35799,N_35738);
and U37728 (N_37728,N_35977,N_34442);
and U37729 (N_37729,N_34322,N_35244);
and U37730 (N_37730,N_34028,N_35509);
nor U37731 (N_37731,N_35064,N_34113);
or U37732 (N_37732,N_35128,N_35254);
or U37733 (N_37733,N_35711,N_34823);
xnor U37734 (N_37734,N_34697,N_35977);
or U37735 (N_37735,N_35624,N_34841);
nor U37736 (N_37736,N_34026,N_34387);
nand U37737 (N_37737,N_35622,N_35733);
and U37738 (N_37738,N_34492,N_35365);
nor U37739 (N_37739,N_34025,N_35213);
xor U37740 (N_37740,N_35690,N_35979);
nor U37741 (N_37741,N_34422,N_34686);
nor U37742 (N_37742,N_35943,N_35684);
and U37743 (N_37743,N_34296,N_34676);
and U37744 (N_37744,N_35760,N_35318);
or U37745 (N_37745,N_34871,N_35394);
nor U37746 (N_37746,N_34539,N_35254);
and U37747 (N_37747,N_35985,N_35291);
or U37748 (N_37748,N_34663,N_34952);
nand U37749 (N_37749,N_35341,N_35782);
and U37750 (N_37750,N_34911,N_35657);
and U37751 (N_37751,N_34475,N_34560);
nand U37752 (N_37752,N_35945,N_34210);
nand U37753 (N_37753,N_34253,N_35260);
nand U37754 (N_37754,N_34679,N_35927);
and U37755 (N_37755,N_34775,N_34069);
xnor U37756 (N_37756,N_35011,N_35746);
or U37757 (N_37757,N_34288,N_34598);
xor U37758 (N_37758,N_34819,N_34870);
or U37759 (N_37759,N_35920,N_34411);
and U37760 (N_37760,N_34054,N_35787);
or U37761 (N_37761,N_35694,N_35970);
xnor U37762 (N_37762,N_34218,N_35837);
nand U37763 (N_37763,N_35597,N_34452);
xor U37764 (N_37764,N_35238,N_34399);
nor U37765 (N_37765,N_34527,N_35174);
or U37766 (N_37766,N_34049,N_34505);
xnor U37767 (N_37767,N_34790,N_34619);
or U37768 (N_37768,N_35248,N_34507);
xnor U37769 (N_37769,N_35860,N_34030);
xnor U37770 (N_37770,N_35569,N_34414);
and U37771 (N_37771,N_34154,N_35186);
and U37772 (N_37772,N_34648,N_34497);
nor U37773 (N_37773,N_35306,N_34501);
xnor U37774 (N_37774,N_35158,N_35162);
and U37775 (N_37775,N_34989,N_35806);
nor U37776 (N_37776,N_34363,N_35828);
nand U37777 (N_37777,N_34500,N_35966);
and U37778 (N_37778,N_35743,N_35439);
or U37779 (N_37779,N_34588,N_34520);
nand U37780 (N_37780,N_35223,N_34787);
and U37781 (N_37781,N_35578,N_34031);
xor U37782 (N_37782,N_35669,N_35815);
nor U37783 (N_37783,N_34358,N_34604);
nor U37784 (N_37784,N_35713,N_34924);
or U37785 (N_37785,N_34229,N_35286);
nand U37786 (N_37786,N_35812,N_35720);
or U37787 (N_37787,N_35600,N_35500);
or U37788 (N_37788,N_35856,N_35244);
xnor U37789 (N_37789,N_35511,N_34845);
or U37790 (N_37790,N_35819,N_35066);
nor U37791 (N_37791,N_35573,N_35706);
nor U37792 (N_37792,N_35724,N_34754);
xor U37793 (N_37793,N_34731,N_34343);
xor U37794 (N_37794,N_35353,N_35356);
xor U37795 (N_37795,N_34687,N_34236);
xnor U37796 (N_37796,N_35422,N_35295);
or U37797 (N_37797,N_35173,N_35320);
xnor U37798 (N_37798,N_35441,N_34567);
xnor U37799 (N_37799,N_34418,N_34677);
xor U37800 (N_37800,N_34812,N_35801);
or U37801 (N_37801,N_35805,N_34387);
nand U37802 (N_37802,N_35188,N_34600);
or U37803 (N_37803,N_35562,N_34824);
and U37804 (N_37804,N_35162,N_35289);
nand U37805 (N_37805,N_34854,N_35162);
nor U37806 (N_37806,N_34094,N_34534);
xor U37807 (N_37807,N_35269,N_35400);
and U37808 (N_37808,N_35961,N_34994);
and U37809 (N_37809,N_34583,N_35629);
nor U37810 (N_37810,N_34865,N_35681);
nor U37811 (N_37811,N_34632,N_35995);
nor U37812 (N_37812,N_35331,N_35645);
xor U37813 (N_37813,N_35567,N_35092);
xnor U37814 (N_37814,N_35618,N_35507);
nand U37815 (N_37815,N_35603,N_35727);
nor U37816 (N_37816,N_35210,N_34821);
and U37817 (N_37817,N_34147,N_35854);
xor U37818 (N_37818,N_34127,N_34087);
nor U37819 (N_37819,N_34690,N_35344);
or U37820 (N_37820,N_35989,N_35410);
or U37821 (N_37821,N_34527,N_35491);
xnor U37822 (N_37822,N_35013,N_34284);
nor U37823 (N_37823,N_35039,N_34912);
xnor U37824 (N_37824,N_35825,N_34769);
or U37825 (N_37825,N_34760,N_34700);
and U37826 (N_37826,N_34340,N_35274);
nand U37827 (N_37827,N_34806,N_34566);
xnor U37828 (N_37828,N_34616,N_34387);
xor U37829 (N_37829,N_34011,N_35964);
or U37830 (N_37830,N_35384,N_35915);
or U37831 (N_37831,N_35702,N_35144);
xnor U37832 (N_37832,N_34917,N_34628);
or U37833 (N_37833,N_35931,N_35650);
nand U37834 (N_37834,N_34884,N_35954);
nand U37835 (N_37835,N_35410,N_34669);
nor U37836 (N_37836,N_35166,N_34967);
xnor U37837 (N_37837,N_34917,N_34751);
or U37838 (N_37838,N_34052,N_34239);
xnor U37839 (N_37839,N_34987,N_34673);
nand U37840 (N_37840,N_35174,N_35739);
xnor U37841 (N_37841,N_34663,N_35486);
xnor U37842 (N_37842,N_35345,N_34008);
and U37843 (N_37843,N_35325,N_35102);
or U37844 (N_37844,N_35975,N_35225);
nor U37845 (N_37845,N_34004,N_34138);
nand U37846 (N_37846,N_34925,N_34932);
xor U37847 (N_37847,N_35348,N_35605);
and U37848 (N_37848,N_35214,N_35031);
xor U37849 (N_37849,N_34834,N_34717);
or U37850 (N_37850,N_35922,N_35919);
xnor U37851 (N_37851,N_34325,N_35121);
or U37852 (N_37852,N_34940,N_35175);
xor U37853 (N_37853,N_34056,N_35446);
nor U37854 (N_37854,N_35176,N_35388);
nand U37855 (N_37855,N_35028,N_35496);
and U37856 (N_37856,N_35246,N_34072);
or U37857 (N_37857,N_34283,N_34047);
nor U37858 (N_37858,N_34585,N_34309);
nand U37859 (N_37859,N_34045,N_34243);
nand U37860 (N_37860,N_35541,N_34134);
or U37861 (N_37861,N_34221,N_34539);
nor U37862 (N_37862,N_34655,N_35146);
nand U37863 (N_37863,N_35643,N_35777);
nand U37864 (N_37864,N_35244,N_34732);
nand U37865 (N_37865,N_35111,N_35611);
nor U37866 (N_37866,N_35055,N_35220);
nand U37867 (N_37867,N_34966,N_35266);
nand U37868 (N_37868,N_34817,N_34124);
nor U37869 (N_37869,N_34469,N_34644);
or U37870 (N_37870,N_35324,N_34278);
nor U37871 (N_37871,N_35056,N_35089);
nor U37872 (N_37872,N_35702,N_35587);
nor U37873 (N_37873,N_35047,N_35806);
or U37874 (N_37874,N_35552,N_35806);
nand U37875 (N_37875,N_34997,N_35812);
xor U37876 (N_37876,N_35240,N_35963);
nor U37877 (N_37877,N_34979,N_34479);
xor U37878 (N_37878,N_35847,N_34239);
nor U37879 (N_37879,N_34835,N_35899);
or U37880 (N_37880,N_34368,N_35532);
and U37881 (N_37881,N_34435,N_34722);
nand U37882 (N_37882,N_34720,N_35279);
nand U37883 (N_37883,N_35209,N_35537);
nand U37884 (N_37884,N_34543,N_35854);
nand U37885 (N_37885,N_35241,N_35547);
and U37886 (N_37886,N_35577,N_35128);
nand U37887 (N_37887,N_35690,N_34461);
and U37888 (N_37888,N_34615,N_35873);
and U37889 (N_37889,N_34705,N_34578);
nor U37890 (N_37890,N_35944,N_34025);
and U37891 (N_37891,N_34721,N_35705);
and U37892 (N_37892,N_34029,N_35935);
nor U37893 (N_37893,N_34650,N_35695);
and U37894 (N_37894,N_34976,N_35839);
nand U37895 (N_37895,N_34552,N_34675);
and U37896 (N_37896,N_35847,N_34944);
or U37897 (N_37897,N_34847,N_35334);
and U37898 (N_37898,N_34176,N_34376);
or U37899 (N_37899,N_35492,N_34490);
and U37900 (N_37900,N_35704,N_35269);
xor U37901 (N_37901,N_34876,N_34879);
xor U37902 (N_37902,N_35154,N_34234);
xnor U37903 (N_37903,N_34682,N_35425);
and U37904 (N_37904,N_34219,N_34293);
and U37905 (N_37905,N_34499,N_35022);
and U37906 (N_37906,N_35888,N_35332);
nand U37907 (N_37907,N_34176,N_34192);
and U37908 (N_37908,N_34085,N_35537);
or U37909 (N_37909,N_35880,N_35781);
nand U37910 (N_37910,N_34303,N_34419);
xnor U37911 (N_37911,N_34464,N_34618);
nor U37912 (N_37912,N_35677,N_34581);
nor U37913 (N_37913,N_35470,N_35974);
nor U37914 (N_37914,N_34366,N_34298);
nand U37915 (N_37915,N_34802,N_35488);
xnor U37916 (N_37916,N_34941,N_35127);
nor U37917 (N_37917,N_35503,N_34072);
nor U37918 (N_37918,N_35459,N_34565);
xor U37919 (N_37919,N_35922,N_35068);
nand U37920 (N_37920,N_35877,N_34800);
nor U37921 (N_37921,N_35200,N_34759);
nor U37922 (N_37922,N_34354,N_34158);
or U37923 (N_37923,N_34481,N_34967);
nand U37924 (N_37924,N_34759,N_35427);
xor U37925 (N_37925,N_35886,N_34386);
xnor U37926 (N_37926,N_35407,N_34404);
or U37927 (N_37927,N_34463,N_35469);
nand U37928 (N_37928,N_34200,N_34269);
nor U37929 (N_37929,N_34119,N_34674);
xnor U37930 (N_37930,N_35818,N_34721);
or U37931 (N_37931,N_34735,N_35232);
xor U37932 (N_37932,N_35551,N_34551);
xor U37933 (N_37933,N_35788,N_35431);
or U37934 (N_37934,N_35626,N_35069);
and U37935 (N_37935,N_35921,N_34120);
or U37936 (N_37936,N_35172,N_34539);
nand U37937 (N_37937,N_34005,N_35374);
nand U37938 (N_37938,N_35135,N_35879);
or U37939 (N_37939,N_34793,N_34961);
and U37940 (N_37940,N_34376,N_34833);
nand U37941 (N_37941,N_34169,N_35584);
and U37942 (N_37942,N_34237,N_35223);
and U37943 (N_37943,N_35200,N_34347);
and U37944 (N_37944,N_35994,N_35329);
nor U37945 (N_37945,N_35476,N_35522);
or U37946 (N_37946,N_35189,N_35835);
and U37947 (N_37947,N_35617,N_34741);
xor U37948 (N_37948,N_35091,N_35082);
and U37949 (N_37949,N_34673,N_35326);
nand U37950 (N_37950,N_34351,N_35074);
nor U37951 (N_37951,N_35974,N_34482);
nand U37952 (N_37952,N_35453,N_35966);
xnor U37953 (N_37953,N_35204,N_34986);
nor U37954 (N_37954,N_35044,N_34614);
nand U37955 (N_37955,N_35645,N_34527);
nand U37956 (N_37956,N_34636,N_35802);
nand U37957 (N_37957,N_35503,N_34522);
nand U37958 (N_37958,N_35976,N_35284);
nor U37959 (N_37959,N_35826,N_34485);
and U37960 (N_37960,N_35397,N_34889);
nor U37961 (N_37961,N_34674,N_35747);
xnor U37962 (N_37962,N_34544,N_34682);
xnor U37963 (N_37963,N_34918,N_34061);
nand U37964 (N_37964,N_35032,N_34780);
xnor U37965 (N_37965,N_34283,N_34575);
or U37966 (N_37966,N_34330,N_34361);
and U37967 (N_37967,N_34221,N_34727);
or U37968 (N_37968,N_34238,N_35756);
nor U37969 (N_37969,N_34464,N_35438);
xnor U37970 (N_37970,N_35211,N_34122);
nor U37971 (N_37971,N_34865,N_35280);
or U37972 (N_37972,N_34163,N_35788);
xnor U37973 (N_37973,N_35761,N_34143);
nor U37974 (N_37974,N_35702,N_34036);
or U37975 (N_37975,N_35825,N_34232);
and U37976 (N_37976,N_34912,N_35227);
or U37977 (N_37977,N_35821,N_35356);
nand U37978 (N_37978,N_35672,N_35287);
and U37979 (N_37979,N_34564,N_35988);
xor U37980 (N_37980,N_34208,N_34194);
nand U37981 (N_37981,N_34442,N_34893);
nor U37982 (N_37982,N_35742,N_35926);
nand U37983 (N_37983,N_35178,N_34929);
or U37984 (N_37984,N_34035,N_35156);
and U37985 (N_37985,N_35303,N_35704);
xor U37986 (N_37986,N_35399,N_35832);
or U37987 (N_37987,N_35372,N_34725);
nor U37988 (N_37988,N_34126,N_35950);
and U37989 (N_37989,N_34687,N_35375);
nand U37990 (N_37990,N_35080,N_34626);
or U37991 (N_37991,N_34065,N_34737);
xor U37992 (N_37992,N_35735,N_34757);
xnor U37993 (N_37993,N_35769,N_35143);
nor U37994 (N_37994,N_34618,N_34479);
or U37995 (N_37995,N_34258,N_35772);
or U37996 (N_37996,N_35765,N_35705);
nor U37997 (N_37997,N_35929,N_35053);
xor U37998 (N_37998,N_34314,N_34304);
nor U37999 (N_37999,N_34262,N_34698);
nor U38000 (N_38000,N_37302,N_36023);
xnor U38001 (N_38001,N_37863,N_37184);
nor U38002 (N_38002,N_36237,N_37736);
xor U38003 (N_38003,N_36810,N_36929);
or U38004 (N_38004,N_37940,N_37014);
or U38005 (N_38005,N_37102,N_37269);
nor U38006 (N_38006,N_36848,N_37732);
and U38007 (N_38007,N_36471,N_36343);
nand U38008 (N_38008,N_37376,N_37679);
nand U38009 (N_38009,N_36521,N_37566);
or U38010 (N_38010,N_36233,N_37455);
or U38011 (N_38011,N_36268,N_37946);
nand U38012 (N_38012,N_36325,N_36622);
xor U38013 (N_38013,N_36407,N_36254);
or U38014 (N_38014,N_36024,N_36862);
nand U38015 (N_38015,N_37359,N_37999);
nand U38016 (N_38016,N_36116,N_36297);
nor U38017 (N_38017,N_36164,N_36844);
nor U38018 (N_38018,N_36758,N_36732);
or U38019 (N_38019,N_37320,N_37172);
or U38020 (N_38020,N_37664,N_36835);
xor U38021 (N_38021,N_37332,N_36993);
nor U38022 (N_38022,N_37991,N_37143);
nand U38023 (N_38023,N_36368,N_37174);
or U38024 (N_38024,N_37258,N_37669);
nor U38025 (N_38025,N_37207,N_36861);
xor U38026 (N_38026,N_36406,N_36387);
xnor U38027 (N_38027,N_36624,N_36229);
and U38028 (N_38028,N_37949,N_36634);
nor U38029 (N_38029,N_37276,N_36887);
nand U38030 (N_38030,N_37009,N_37074);
nor U38031 (N_38031,N_37414,N_36126);
nor U38032 (N_38032,N_36917,N_37809);
or U38033 (N_38033,N_37213,N_36720);
or U38034 (N_38034,N_37812,N_36985);
nand U38035 (N_38035,N_36014,N_37824);
or U38036 (N_38036,N_37981,N_36974);
nor U38037 (N_38037,N_37587,N_36678);
nand U38038 (N_38038,N_36599,N_36376);
nand U38039 (N_38039,N_36592,N_36777);
nor U38040 (N_38040,N_37186,N_36136);
nand U38041 (N_38041,N_37839,N_37987);
nand U38042 (N_38042,N_37154,N_37973);
and U38043 (N_38043,N_37619,N_37611);
and U38044 (N_38044,N_37557,N_37864);
or U38045 (N_38045,N_36837,N_37179);
nand U38046 (N_38046,N_37032,N_36053);
and U38047 (N_38047,N_36517,N_36561);
nor U38048 (N_38048,N_36933,N_36138);
or U38049 (N_38049,N_37261,N_37432);
xor U38050 (N_38050,N_36943,N_36415);
nand U38051 (N_38051,N_37115,N_37251);
or U38052 (N_38052,N_36260,N_37831);
xnor U38053 (N_38053,N_36977,N_37869);
and U38054 (N_38054,N_36869,N_37028);
and U38055 (N_38055,N_36265,N_37485);
nand U38056 (N_38056,N_36157,N_37390);
xnor U38057 (N_38057,N_37694,N_37397);
nand U38058 (N_38058,N_37726,N_36896);
or U38059 (N_38059,N_36401,N_37707);
and U38060 (N_38060,N_36082,N_36477);
or U38061 (N_38061,N_36209,N_36289);
xor U38062 (N_38062,N_37626,N_36762);
xnor U38063 (N_38063,N_36286,N_36476);
xor U38064 (N_38064,N_36315,N_36152);
nand U38065 (N_38065,N_36399,N_37110);
or U38066 (N_38066,N_37042,N_36095);
nand U38067 (N_38067,N_37017,N_37459);
or U38068 (N_38068,N_36058,N_37328);
nor U38069 (N_38069,N_36834,N_36290);
xor U38070 (N_38070,N_36306,N_37590);
and U38071 (N_38071,N_37501,N_37807);
or U38072 (N_38072,N_37189,N_36267);
nand U38073 (N_38073,N_36059,N_37099);
nand U38074 (N_38074,N_37684,N_36191);
xnor U38075 (N_38075,N_36203,N_37625);
nor U38076 (N_38076,N_37272,N_37943);
or U38077 (N_38077,N_37550,N_36804);
xnor U38078 (N_38078,N_36990,N_37280);
and U38079 (N_38079,N_37303,N_36466);
xor U38080 (N_38080,N_37479,N_36020);
nor U38081 (N_38081,N_36405,N_37537);
xor U38082 (N_38082,N_36270,N_36201);
and U38083 (N_38083,N_37313,N_36960);
nor U38084 (N_38084,N_37446,N_36035);
nand U38085 (N_38085,N_36587,N_36514);
xnor U38086 (N_38086,N_36404,N_37615);
nand U38087 (N_38087,N_36937,N_37621);
nand U38088 (N_38088,N_36668,N_36833);
nand U38089 (N_38089,N_36319,N_37784);
or U38090 (N_38090,N_36602,N_36432);
xnor U38091 (N_38091,N_36066,N_36108);
and U38092 (N_38092,N_37416,N_36934);
nand U38093 (N_38093,N_36253,N_37434);
nand U38094 (N_38094,N_37702,N_37494);
and U38095 (N_38095,N_36391,N_37541);
or U38096 (N_38096,N_37342,N_37122);
nand U38097 (N_38097,N_36045,N_37796);
and U38098 (N_38098,N_36904,N_37523);
nand U38099 (N_38099,N_37935,N_37388);
xnor U38100 (N_38100,N_37551,N_37651);
xnor U38101 (N_38101,N_36748,N_37472);
or U38102 (N_38102,N_37356,N_37780);
xnor U38103 (N_38103,N_37751,N_36515);
nor U38104 (N_38104,N_37959,N_36076);
and U38105 (N_38105,N_36706,N_37828);
nor U38106 (N_38106,N_36802,N_37294);
and U38107 (N_38107,N_36940,N_36222);
or U38108 (N_38108,N_36344,N_37062);
nor U38109 (N_38109,N_36760,N_36147);
nand U38110 (N_38110,N_36021,N_37173);
nor U38111 (N_38111,N_37358,N_36868);
xnor U38112 (N_38112,N_36109,N_36601);
or U38113 (N_38113,N_36845,N_37465);
and U38114 (N_38114,N_36296,N_37212);
xnor U38115 (N_38115,N_36796,N_36825);
nand U38116 (N_38116,N_36957,N_37483);
and U38117 (N_38117,N_37617,N_36687);
and U38118 (N_38118,N_36712,N_36107);
and U38119 (N_38119,N_36828,N_37354);
nand U38120 (N_38120,N_36033,N_37244);
nand U38121 (N_38121,N_37422,N_37881);
xor U38122 (N_38122,N_36840,N_36250);
nand U38123 (N_38123,N_36853,N_37387);
or U38124 (N_38124,N_37867,N_36044);
xor U38125 (N_38125,N_37560,N_37289);
and U38126 (N_38126,N_36008,N_37841);
xor U38127 (N_38127,N_37101,N_37937);
and U38128 (N_38128,N_37366,N_36999);
xnor U38129 (N_38129,N_36909,N_36353);
and U38130 (N_38130,N_37347,N_37141);
nand U38131 (N_38131,N_37435,N_37854);
xnor U38132 (N_38132,N_37445,N_37539);
nand U38133 (N_38133,N_36631,N_37048);
and U38134 (N_38134,N_36574,N_36529);
and U38135 (N_38135,N_36996,N_36124);
xor U38136 (N_38136,N_36936,N_36794);
or U38137 (N_38137,N_36646,N_37673);
or U38138 (N_38138,N_36499,N_36006);
and U38139 (N_38139,N_37984,N_36811);
or U38140 (N_38140,N_36071,N_36459);
and U38141 (N_38141,N_36503,N_37768);
or U38142 (N_38142,N_36623,N_37199);
xor U38143 (N_38143,N_36185,N_37668);
and U38144 (N_38144,N_36806,N_36410);
nor U38145 (N_38145,N_37486,N_37908);
xnor U38146 (N_38146,N_36751,N_37793);
and U38147 (N_38147,N_37293,N_37589);
or U38148 (N_38148,N_37939,N_36475);
xor U38149 (N_38149,N_37852,N_36483);
nand U38150 (N_38150,N_37708,N_36617);
nand U38151 (N_38151,N_36571,N_37473);
xor U38152 (N_38152,N_36952,N_36017);
xor U38153 (N_38153,N_37083,N_36255);
nand U38154 (N_38154,N_36986,N_37309);
xnor U38155 (N_38155,N_36154,N_36779);
nand U38156 (N_38156,N_37629,N_36543);
and U38157 (N_38157,N_36172,N_36615);
xor U38158 (N_38158,N_36140,N_36573);
nand U38159 (N_38159,N_37267,N_37871);
and U38160 (N_38160,N_37635,N_37021);
xnor U38161 (N_38161,N_37470,N_36893);
nor U38162 (N_38162,N_36606,N_36433);
or U38163 (N_38163,N_36106,N_37866);
or U38164 (N_38164,N_36040,N_37755);
xor U38165 (N_38165,N_37531,N_37774);
nand U38166 (N_38166,N_37068,N_36118);
nand U38167 (N_38167,N_36616,N_37515);
xnor U38168 (N_38168,N_36776,N_36962);
nor U38169 (N_38169,N_37795,N_37067);
and U38170 (N_38170,N_36507,N_37420);
and U38171 (N_38171,N_36660,N_36239);
nor U38172 (N_38172,N_37507,N_37652);
xor U38173 (N_38173,N_37331,N_37106);
or U38174 (N_38174,N_37004,N_36866);
and U38175 (N_38175,N_36068,N_37686);
nand U38176 (N_38176,N_37311,N_37941);
xnor U38177 (N_38177,N_36864,N_37606);
or U38178 (N_38178,N_36036,N_36644);
and U38179 (N_38179,N_37257,N_36009);
nand U38180 (N_38180,N_37133,N_36658);
xnor U38181 (N_38181,N_37874,N_37412);
or U38182 (N_38182,N_36520,N_36754);
nand U38183 (N_38183,N_37138,N_37884);
and U38184 (N_38184,N_37654,N_36394);
and U38185 (N_38185,N_37733,N_36998);
nor U38186 (N_38186,N_36490,N_37777);
xor U38187 (N_38187,N_36161,N_36183);
xnor U38188 (N_38188,N_37306,N_36771);
xor U38189 (N_38189,N_37970,N_37558);
or U38190 (N_38190,N_36534,N_36019);
nor U38191 (N_38191,N_37705,N_36655);
nand U38192 (N_38192,N_37570,N_36348);
nand U38193 (N_38193,N_37450,N_36558);
nand U38194 (N_38194,N_36346,N_36080);
xor U38195 (N_38195,N_37909,N_37646);
xor U38196 (N_38196,N_37933,N_36431);
nor U38197 (N_38197,N_36682,N_36288);
or U38198 (N_38198,N_37967,N_36084);
nor U38199 (N_38199,N_37020,N_36285);
nor U38200 (N_38200,N_37075,N_37128);
nand U38201 (N_38201,N_37156,N_37781);
nor U38202 (N_38202,N_37591,N_36261);
xnor U38203 (N_38203,N_36843,N_36247);
or U38204 (N_38204,N_37339,N_37369);
nor U38205 (N_38205,N_36241,N_36951);
nor U38206 (N_38206,N_37197,N_37948);
nor U38207 (N_38207,N_37081,N_36892);
and U38208 (N_38208,N_37428,N_37256);
xor U38209 (N_38209,N_36565,N_37988);
nor U38210 (N_38210,N_36753,N_36377);
and U38211 (N_38211,N_36357,N_36980);
or U38212 (N_38212,N_36264,N_36438);
xor U38213 (N_38213,N_37748,N_37527);
and U38214 (N_38214,N_36412,N_36860);
and U38215 (N_38215,N_37975,N_37892);
and U38216 (N_38216,N_36470,N_37015);
nor U38217 (N_38217,N_37936,N_37518);
or U38218 (N_38218,N_36204,N_37301);
nand U38219 (N_38219,N_36046,N_36362);
and U38220 (N_38220,N_36497,N_37082);
nor U38221 (N_38221,N_37957,N_36910);
xor U38222 (N_38222,N_36293,N_37016);
or U38223 (N_38223,N_36689,N_37030);
and U38224 (N_38224,N_36820,N_36114);
xnor U38225 (N_38225,N_37103,N_37182);
xnor U38226 (N_38226,N_37219,N_36303);
xnor U38227 (N_38227,N_37964,N_36756);
nand U38228 (N_38228,N_37150,N_36211);
and U38229 (N_38229,N_37752,N_36926);
nor U38230 (N_38230,N_36322,N_37756);
nand U38231 (N_38231,N_36620,N_36890);
nand U38232 (N_38232,N_36179,N_36025);
xor U38233 (N_38233,N_36461,N_36484);
nor U38234 (N_38234,N_36567,N_36151);
and U38235 (N_38235,N_36047,N_37057);
nand U38236 (N_38236,N_36105,N_36944);
nor U38237 (N_38237,N_37319,N_36971);
xnor U38238 (N_38238,N_37125,N_36938);
or U38239 (N_38239,N_36345,N_36425);
nor U38240 (N_38240,N_37166,N_36428);
and U38241 (N_38241,N_37209,N_37399);
xor U38242 (N_38242,N_37146,N_37353);
xor U38243 (N_38243,N_37721,N_36783);
xor U38244 (N_38244,N_36468,N_37047);
nand U38245 (N_38245,N_37253,N_37105);
or U38246 (N_38246,N_37323,N_37955);
xor U38247 (N_38247,N_36628,N_36175);
and U38248 (N_38248,N_36048,N_37167);
and U38249 (N_38249,N_36457,N_36367);
or U38250 (N_38250,N_36454,N_36294);
nor U38251 (N_38251,N_36436,N_37547);
or U38252 (N_38252,N_37231,N_36453);
or U38253 (N_38253,N_37490,N_36347);
xor U38254 (N_38254,N_37906,N_36532);
xor U38255 (N_38255,N_37198,N_36123);
and U38256 (N_38256,N_37805,N_36111);
xor U38257 (N_38257,N_37297,N_37642);
nor U38258 (N_38258,N_37623,N_36973);
nand U38259 (N_38259,N_37120,N_37903);
or U38260 (N_38260,N_36088,N_36667);
xor U38261 (N_38261,N_37535,N_36186);
nand U38262 (N_38262,N_36767,N_36472);
xor U38263 (N_38263,N_36130,N_37282);
nor U38264 (N_38264,N_36257,N_36330);
xnor U38265 (N_38265,N_37893,N_36182);
nand U38266 (N_38266,N_36536,N_37475);
nand U38267 (N_38267,N_36016,N_37093);
or U38268 (N_38268,N_36988,N_36994);
and U38269 (N_38269,N_37976,N_36739);
and U38270 (N_38270,N_36078,N_37861);
nand U38271 (N_38271,N_37430,N_36932);
and U38272 (N_38272,N_37980,N_36277);
xor U38273 (N_38273,N_37529,N_36366);
xnor U38274 (N_38274,N_37767,N_36452);
xor U38275 (N_38275,N_37891,N_37840);
nand U38276 (N_38276,N_36649,N_36530);
and U38277 (N_38277,N_36137,N_36546);
xor U38278 (N_38278,N_36654,N_37215);
or U38279 (N_38279,N_37211,N_37208);
xor U38280 (N_38280,N_36456,N_36057);
or U38281 (N_38281,N_37917,N_36077);
nor U38282 (N_38282,N_37990,N_36800);
nand U38283 (N_38283,N_37951,N_36830);
xnor U38284 (N_38284,N_36384,N_37779);
or U38285 (N_38285,N_37210,N_36488);
or U38286 (N_38286,N_36721,N_37640);
nor U38287 (N_38287,N_37985,N_36018);
or U38288 (N_38288,N_36437,N_37098);
nand U38289 (N_38289,N_36727,N_37913);
or U38290 (N_38290,N_36763,N_36772);
and U38291 (N_38291,N_36846,N_36128);
xor U38292 (N_38292,N_37500,N_36626);
and U38293 (N_38293,N_37860,N_36564);
xnor U38294 (N_38294,N_36312,N_37790);
nor U38295 (N_38295,N_37438,N_37696);
xor U38296 (N_38296,N_37401,N_37914);
or U38297 (N_38297,N_37380,N_36923);
or U38298 (N_38298,N_37938,N_37722);
nor U38299 (N_38299,N_37757,N_37018);
nor U38300 (N_38300,N_37723,N_37743);
or U38301 (N_38301,N_37436,N_36273);
nor U38302 (N_38302,N_36693,N_37806);
and U38303 (N_38303,N_37711,N_36092);
or U38304 (N_38304,N_36907,N_37540);
xnor U38305 (N_38305,N_36842,N_37569);
xnor U38306 (N_38306,N_37419,N_37672);
nor U38307 (N_38307,N_37274,N_37317);
nand U38308 (N_38308,N_36978,N_37247);
nand U38309 (N_38309,N_36585,N_36508);
xor U38310 (N_38310,N_37682,N_36956);
or U38311 (N_38311,N_36263,N_37895);
nor U38312 (N_38312,N_36174,N_36226);
xnor U38313 (N_38313,N_37063,N_36618);
nor U38314 (N_38314,N_37859,N_37411);
or U38315 (N_38315,N_36555,N_36176);
xor U38316 (N_38316,N_37066,N_36880);
and U38317 (N_38317,N_37204,N_36695);
or U38318 (N_38318,N_37942,N_37266);
nand U38319 (N_38319,N_37088,N_36121);
or U38320 (N_38320,N_36112,N_36955);
or U38321 (N_38321,N_36908,N_37229);
and U38322 (N_38322,N_36948,N_36575);
and U38323 (N_38323,N_37375,N_36370);
nor U38324 (N_38324,N_36075,N_36413);
and U38325 (N_38325,N_37384,N_36418);
nor U38326 (N_38326,N_37457,N_36663);
and U38327 (N_38327,N_37264,N_37202);
nand U38328 (N_38328,N_36232,N_37548);
nand U38329 (N_38329,N_37160,N_37162);
nor U38330 (N_38330,N_37993,N_36403);
and U38331 (N_38331,N_36984,N_36153);
or U38332 (N_38332,N_36709,N_36146);
nand U38333 (N_38333,N_36921,N_36785);
xnor U38334 (N_38334,N_36166,N_36967);
nand U38335 (N_38335,N_37534,N_36746);
nand U38336 (N_38336,N_36559,N_36870);
nand U38337 (N_38337,N_37118,N_37553);
xnor U38338 (N_38338,N_37627,N_36474);
or U38339 (N_38339,N_36479,N_36552);
nand U38340 (N_38340,N_36248,N_36676);
and U38341 (N_38341,N_37753,N_36005);
xnor U38342 (N_38342,N_37151,N_37729);
and U38343 (N_38343,N_37050,N_36291);
and U38344 (N_38344,N_37952,N_37766);
and U38345 (N_38345,N_37578,N_37348);
or U38346 (N_38346,N_36188,N_36691);
xnor U38347 (N_38347,N_36583,N_37546);
xnor U38348 (N_38348,N_37761,N_36298);
and U38349 (N_38349,N_36013,N_36621);
xor U38350 (N_38350,N_37602,N_37883);
xnor U38351 (N_38351,N_37950,N_37246);
and U38352 (N_38352,N_37504,N_36549);
xor U38353 (N_38353,N_37055,N_36886);
xor U38354 (N_38354,N_37789,N_37396);
and U38355 (N_38355,N_37327,N_36451);
nor U38356 (N_38356,N_37349,N_37144);
nor U38357 (N_38357,N_37600,N_36749);
nor U38358 (N_38358,N_36321,N_37023);
nor U38359 (N_38359,N_37441,N_36374);
or U38360 (N_38360,N_36714,N_36307);
and U38361 (N_38361,N_37239,N_37314);
or U38362 (N_38362,N_37706,N_37573);
and U38363 (N_38363,N_36604,N_36510);
nor U38364 (N_38364,N_36177,N_37300);
nand U38365 (N_38365,N_36317,N_37690);
xor U38366 (N_38366,N_37810,N_37899);
nor U38367 (N_38367,N_37870,N_37265);
or U38368 (N_38368,N_37851,N_36323);
xor U38369 (N_38369,N_36947,N_37155);
or U38370 (N_38370,N_37811,N_36449);
xor U38371 (N_38371,N_36939,N_37372);
xor U38372 (N_38372,N_36141,N_36832);
xor U38373 (N_38373,N_36029,N_37808);
and U38374 (N_38374,N_37214,N_36899);
or U38375 (N_38375,N_37206,N_37510);
xor U38376 (N_38376,N_37394,N_37008);
or U38377 (N_38377,N_37292,N_36494);
nand U38378 (N_38378,N_36897,N_37176);
or U38379 (N_38379,N_36213,N_37759);
or U38380 (N_38380,N_36478,N_37355);
nor U38381 (N_38381,N_37901,N_37056);
xnor U38382 (N_38382,N_37846,N_36110);
nor U38383 (N_38383,N_36089,N_36160);
nor U38384 (N_38384,N_36102,N_37410);
xnor U38385 (N_38385,N_36653,N_37561);
xor U38386 (N_38386,N_37177,N_37368);
nand U38387 (N_38387,N_36769,N_36411);
xnor U38388 (N_38388,N_37613,N_37928);
nor U38389 (N_38389,N_37581,N_36504);
nor U38390 (N_38390,N_36424,N_36310);
or U38391 (N_38391,N_36557,N_37966);
or U38392 (N_38392,N_36526,N_36389);
xnor U38393 (N_38393,N_36770,N_36826);
and U38394 (N_38394,N_36196,N_36512);
or U38395 (N_38395,N_36647,N_37147);
nand U38396 (N_38396,N_37749,N_36755);
nor U38397 (N_38397,N_36664,N_36607);
nor U38398 (N_38398,N_37498,N_37429);
nor U38399 (N_38399,N_36100,N_37270);
nand U38400 (N_38400,N_37709,N_37491);
xor U38401 (N_38401,N_36184,N_36795);
or U38402 (N_38402,N_37769,N_36895);
or U38403 (N_38403,N_37844,N_36619);
or U38404 (N_38404,N_36450,N_36591);
nand U38405 (N_38405,N_36115,N_37787);
or U38406 (N_38406,N_36383,N_36903);
nand U38407 (N_38407,N_36919,N_37754);
nor U38408 (N_38408,N_36819,N_36673);
xor U38409 (N_38409,N_37877,N_36032);
nand U38410 (N_38410,N_37737,N_36822);
xnor U38411 (N_38411,N_36349,N_37005);
and U38412 (N_38412,N_37001,N_37575);
and U38413 (N_38413,N_37816,N_36614);
or U38414 (N_38414,N_37637,N_37163);
or U38415 (N_38415,N_37739,N_36827);
xor U38416 (N_38416,N_36600,N_37232);
xor U38417 (N_38417,N_36473,N_36747);
or U38418 (N_38418,N_37997,N_36657);
xor U38419 (N_38419,N_37078,N_37853);
xnor U38420 (N_38420,N_37471,N_36788);
xnor U38421 (N_38421,N_36198,N_37094);
nor U38422 (N_38422,N_37727,N_37567);
and U38423 (N_38423,N_36836,N_37452);
nand U38424 (N_38424,N_37760,N_36231);
or U38425 (N_38425,N_36632,N_36959);
or U38426 (N_38426,N_37788,N_37284);
nand U38427 (N_38427,N_36354,N_37373);
xor U38428 (N_38428,N_36545,N_36731);
nor U38429 (N_38429,N_37580,N_36636);
and U38430 (N_38430,N_37765,N_36275);
or U38431 (N_38431,N_36675,N_36421);
and U38432 (N_38432,N_36928,N_36234);
nand U38433 (N_38433,N_37670,N_37910);
xor U38434 (N_38434,N_36331,N_36305);
xnor U38435 (N_38435,N_37944,N_37059);
and U38436 (N_38436,N_36379,N_37227);
and U38437 (N_38437,N_37108,N_37250);
or U38438 (N_38438,N_36839,N_36611);
and U38439 (N_38439,N_37724,N_37821);
and U38440 (N_38440,N_37362,N_37169);
nor U38441 (N_38441,N_36790,N_36324);
nand U38442 (N_38442,N_37834,N_37890);
and U38443 (N_38443,N_36417,N_36011);
xnor U38444 (N_38444,N_36638,N_37130);
or U38445 (N_38445,N_37312,N_37818);
or U38446 (N_38446,N_37351,N_36181);
and U38447 (N_38447,N_36003,N_36945);
nand U38448 (N_38448,N_37403,N_36086);
or U38449 (N_38449,N_36259,N_36134);
nor U38450 (N_38450,N_36171,N_36236);
and U38451 (N_38451,N_37091,N_37113);
xnor U38452 (N_38452,N_36042,N_36094);
or U38453 (N_38453,N_36408,N_37140);
or U38454 (N_38454,N_37220,N_37862);
or U38455 (N_38455,N_37268,N_36878);
nor U38456 (N_38456,N_37181,N_36801);
nor U38457 (N_38457,N_36395,N_36272);
and U38458 (N_38458,N_36652,N_37947);
xnor U38459 (N_38459,N_36439,N_36659);
xnor U38460 (N_38460,N_37666,N_36576);
xnor U38461 (N_38461,N_37555,N_36043);
nor U38462 (N_38462,N_36780,N_36007);
xnor U38463 (N_38463,N_37413,N_37880);
xor U38464 (N_38464,N_37868,N_37655);
and U38465 (N_38465,N_37927,N_37636);
nor U38466 (N_38466,N_37524,N_37357);
or U38467 (N_38467,N_36584,N_36158);
and U38468 (N_38468,N_36527,N_37803);
or U38469 (N_38469,N_37377,N_36073);
and U38470 (N_38470,N_36429,N_36975);
xnor U38471 (N_38471,N_36462,N_37404);
nand U38472 (N_38472,N_36339,N_36015);
nor U38473 (N_38473,N_37885,N_37334);
or U38474 (N_38474,N_37601,N_36665);
xnor U38475 (N_38475,N_37389,N_37006);
xor U38476 (N_38476,N_36744,N_36946);
or U38477 (N_38477,N_37386,N_37681);
or U38478 (N_38478,N_37418,N_37907);
xnor U38479 (N_38479,N_36651,N_37982);
or U38480 (N_38480,N_36969,N_37833);
and U38481 (N_38481,N_37563,N_36210);
nor U38482 (N_38482,N_36093,N_36309);
nand U38483 (N_38483,N_37750,N_37659);
nor U38484 (N_38484,N_36375,N_36361);
xnor U38485 (N_38485,N_37433,N_36096);
and U38486 (N_38486,N_37241,N_36240);
nand U38487 (N_38487,N_37638,N_36097);
nand U38488 (N_38488,N_36884,N_37425);
nand U38489 (N_38489,N_36335,N_37379);
or U38490 (N_38490,N_37308,N_37603);
and U38491 (N_38491,N_37665,N_37352);
nand U38492 (N_38492,N_36012,N_36279);
nand U38493 (N_38493,N_36441,N_37090);
nand U38494 (N_38494,N_36580,N_37089);
and U38495 (N_38495,N_37010,N_36519);
nand U38496 (N_38496,N_37287,N_36807);
and U38497 (N_38497,N_37667,N_37661);
and U38498 (N_38498,N_37195,N_36246);
and U38499 (N_38499,N_37911,N_36717);
or U38500 (N_38500,N_36352,N_37164);
and U38501 (N_38501,N_37924,N_37631);
and U38502 (N_38502,N_37782,N_36726);
xnor U38503 (N_38503,N_37785,N_36742);
nor U38504 (N_38504,N_36393,N_36067);
nand U38505 (N_38505,N_36050,N_37026);
or U38506 (N_38506,N_37764,N_37142);
nor U38507 (N_38507,N_36511,N_37053);
nor U38508 (N_38508,N_37556,N_36301);
nand U38509 (N_38509,N_37378,N_37337);
nand U38510 (N_38510,N_36207,N_36730);
nor U38511 (N_38511,N_37238,N_36091);
and U38512 (N_38512,N_37597,N_37513);
nand U38513 (N_38513,N_37674,N_36435);
nor U38514 (N_38514,N_36900,N_36873);
and U38515 (N_38515,N_37582,N_36480);
or U38516 (N_38516,N_37585,N_37039);
nand U38517 (N_38517,N_36027,N_37117);
nor U38518 (N_38518,N_37983,N_37634);
nor U38519 (N_38519,N_36821,N_36139);
or U38520 (N_38520,N_37499,N_37643);
nor U38521 (N_38521,N_36596,N_37461);
nor U38522 (N_38522,N_36690,N_36931);
or U38523 (N_38523,N_36541,N_36481);
nand U38524 (N_38524,N_37649,N_37084);
or U38525 (N_38525,N_36090,N_36442);
xnor U38526 (N_38526,N_36752,N_36064);
nor U38527 (N_38527,N_37526,N_37095);
nor U38528 (N_38528,N_37598,N_36206);
nor U38529 (N_38529,N_37364,N_37458);
nand U38530 (N_38530,N_36789,N_37183);
nand U38531 (N_38531,N_37190,N_36823);
nor U38532 (N_38532,N_37149,N_36735);
and U38533 (N_38533,N_37002,N_37979);
or U38534 (N_38534,N_37382,N_37596);
xor U38535 (N_38535,N_36165,N_36518);
and U38536 (N_38536,N_36148,N_36104);
nand U38537 (N_38537,N_36156,N_37747);
nor U38538 (N_38538,N_36063,N_37791);
nand U38539 (N_38539,N_37007,N_37505);
nor U38540 (N_38540,N_36911,N_36797);
or U38541 (N_38541,N_36872,N_37153);
and U38542 (N_38542,N_37444,N_37409);
xnor U38543 (N_38543,N_36491,N_37716);
and U38544 (N_38544,N_36195,N_37165);
nand U38545 (N_38545,N_36740,N_36320);
nand U38546 (N_38546,N_36528,N_37639);
nor U38547 (N_38547,N_37579,N_37571);
and U38548 (N_38548,N_37076,N_36083);
nor U38549 (N_38549,N_37407,N_37431);
nor U38550 (N_38550,N_37468,N_37516);
nor U38551 (N_38551,N_36793,N_36637);
nand U38552 (N_38552,N_37963,N_36002);
nor U38553 (N_38553,N_36129,N_37157);
xnor U38554 (N_38554,N_37819,N_37205);
xnor U38555 (N_38555,N_37235,N_37281);
xnor U38556 (N_38556,N_36901,N_37406);
and U38557 (N_38557,N_37283,N_37677);
nor U38558 (N_38558,N_36455,N_37912);
xor U38559 (N_38559,N_37676,N_37887);
and U38560 (N_38560,N_36132,N_37124);
nand U38561 (N_38561,N_36738,N_36278);
xnor U38562 (N_38562,N_36876,N_36467);
xnor U38563 (N_38563,N_36113,N_36863);
nor U38564 (N_38564,N_37064,N_37464);
or U38565 (N_38565,N_37324,N_36276);
nor U38566 (N_38566,N_36891,N_37203);
nor U38567 (N_38567,N_37079,N_37478);
nand U38568 (N_38568,N_36028,N_37929);
or U38569 (N_38569,N_37495,N_37720);
and U38570 (N_38570,N_37630,N_36034);
or U38571 (N_38571,N_36099,N_36685);
nand U38572 (N_38572,N_36538,N_37236);
nand U38573 (N_38573,N_37632,N_37715);
nor U38574 (N_38574,N_36803,N_37998);
nand U38575 (N_38575,N_37735,N_36143);
and U38576 (N_38576,N_37827,N_37427);
xor U38577 (N_38577,N_36879,N_36694);
and U38578 (N_38578,N_37678,N_37593);
xor U38579 (N_38579,N_36258,N_37506);
and U38580 (N_38580,N_36818,N_36463);
or U38581 (N_38581,N_37439,N_36674);
or U38582 (N_38582,N_37657,N_37290);
xnor U38583 (N_38583,N_36784,N_37037);
and U38584 (N_38584,N_37921,N_37307);
or U38585 (N_38585,N_36841,N_37318);
or U38586 (N_38586,N_36242,N_36681);
and U38587 (N_38587,N_37288,N_36283);
nand U38588 (N_38588,N_37221,N_36650);
xor U38589 (N_38589,N_37145,N_36913);
and U38590 (N_38590,N_36953,N_36851);
nand U38591 (N_38591,N_37583,N_37240);
xnor U38592 (N_38592,N_37092,N_37346);
or U38593 (N_38593,N_36669,N_36648);
or U38594 (N_38594,N_37545,N_36218);
nand U38595 (N_38595,N_36142,N_36392);
nor U38596 (N_38596,N_36949,N_37586);
nand U38597 (N_38597,N_36072,N_36163);
nand U38598 (N_38598,N_36051,N_36958);
and U38599 (N_38599,N_36965,N_37763);
and U38600 (N_38600,N_37622,N_37111);
xnor U38601 (N_38601,N_37758,N_37194);
nand U38602 (N_38602,N_36101,N_36365);
nor U38603 (N_38603,N_36062,N_36460);
xnor U38604 (N_38604,N_37857,N_37228);
nand U38605 (N_38605,N_36799,N_37918);
and U38606 (N_38606,N_37391,N_36125);
or U38607 (N_38607,N_37878,N_37826);
nand U38608 (N_38608,N_37363,N_36194);
or U38609 (N_38609,N_37476,N_37837);
and U38610 (N_38610,N_37799,N_36224);
nand U38611 (N_38611,N_37178,N_36641);
xor U38612 (N_38612,N_36214,N_36482);
and U38613 (N_38613,N_37977,N_36629);
nand U38614 (N_38614,N_37894,N_36420);
nand U38615 (N_38615,N_36235,N_37695);
xor U38616 (N_38616,N_37503,N_37725);
xnor U38617 (N_38617,N_37474,N_36625);
and U38618 (N_38618,N_36373,N_37159);
nor U38619 (N_38619,N_37691,N_36877);
nand U38620 (N_38620,N_36854,N_36544);
xnor U38621 (N_38621,N_37873,N_37045);
xnor U38622 (N_38622,N_37060,N_37426);
and U38623 (N_38623,N_36539,N_37820);
xnor U38624 (N_38624,N_36326,N_37070);
nor U38625 (N_38625,N_36696,N_36871);
xor U38626 (N_38626,N_37038,N_37259);
nand U38627 (N_38627,N_37033,N_36905);
nor U38628 (N_38628,N_36723,N_37517);
xnor U38629 (N_38629,N_37776,N_37856);
or U38630 (N_38630,N_37134,N_37511);
nor U38631 (N_38631,N_37322,N_36505);
nand U38632 (N_38632,N_36220,N_36577);
and U38633 (N_38633,N_36223,N_37011);
nor U38634 (N_38634,N_36227,N_37338);
and U38635 (N_38635,N_36757,N_36612);
xor U38636 (N_38636,N_36447,N_36423);
xnor U38637 (N_38637,N_36513,N_37592);
nand U38638 (N_38638,N_36060,N_37734);
or U38639 (N_38639,N_36922,N_37609);
nor U38640 (N_38640,N_37934,N_37978);
nand U38641 (N_38641,N_37919,N_37393);
and U38642 (N_38642,N_37956,N_36551);
nand U38643 (N_38643,N_36244,N_36888);
nor U38644 (N_38644,N_37663,N_37180);
xnor U38645 (N_38645,N_37193,N_37989);
nor U38646 (N_38646,N_37797,N_36976);
xor U38647 (N_38647,N_36409,N_36671);
or U38648 (N_38648,N_36200,N_37624);
nand U38649 (N_38649,N_36486,N_36282);
or U38650 (N_38650,N_37242,N_36643);
or U38651 (N_38651,N_37000,N_37469);
xnor U38652 (N_38652,N_36364,N_37442);
or U38653 (N_38653,N_37365,N_37405);
nand U38654 (N_38654,N_36595,N_36914);
xor U38655 (N_38655,N_36808,N_36065);
and U38656 (N_38656,N_36787,N_36197);
or U38657 (N_38657,N_36656,N_37136);
xor U38658 (N_38658,N_36496,N_37168);
nor U38659 (N_38659,N_37572,N_37344);
xnor U38660 (N_38660,N_36509,N_37520);
or U38661 (N_38661,N_36316,N_36444);
and U38662 (N_38662,N_37607,N_37620);
and U38663 (N_38663,N_36707,N_36838);
xor U38664 (N_38664,N_37986,N_37565);
and U38665 (N_38665,N_36701,N_36135);
nand U38666 (N_38666,N_37321,N_36026);
nor U38667 (N_38667,N_36328,N_37965);
nand U38668 (N_38668,N_36711,N_37522);
and U38669 (N_38669,N_36569,N_36855);
and U38670 (N_38670,N_37644,N_37509);
xnor U38671 (N_38671,N_36180,N_36190);
nand U38672 (N_38672,N_37271,N_37704);
and U38673 (N_38673,N_36085,N_37285);
or U38674 (N_38674,N_36563,N_37838);
xor U38675 (N_38675,N_37326,N_36719);
xnor U38676 (N_38676,N_36422,N_37171);
nor U38677 (N_38677,N_37482,N_36173);
xnor U38678 (N_38678,N_37158,N_36145);
and U38679 (N_38679,N_36292,N_37316);
and U38680 (N_38680,N_36608,N_36249);
nor U38681 (N_38681,N_36849,N_37916);
or U38682 (N_38682,N_36284,N_37683);
nor U38683 (N_38683,N_36768,N_37329);
or U38684 (N_38684,N_37296,N_36252);
or U38685 (N_38685,N_37595,N_37350);
nor U38686 (N_38686,N_37648,N_36350);
xor U38687 (N_38687,N_37467,N_36041);
nand U38688 (N_38688,N_36774,N_37783);
or U38689 (N_38689,N_37310,N_36489);
xnor U38690 (N_38690,N_37594,N_37061);
xnor U38691 (N_38691,N_37879,N_36351);
nor U38692 (N_38692,N_36889,N_36765);
and U38693 (N_38693,N_36692,N_36684);
nor U38694 (N_38694,N_37466,N_36764);
xor U38695 (N_38695,N_36736,N_36728);
nand U38696 (N_38696,N_36337,N_37371);
nor U38697 (N_38697,N_36131,N_36699);
nand U38698 (N_38698,N_37069,N_36725);
and U38699 (N_38699,N_36371,N_36927);
nand U38700 (N_38700,N_37487,N_36448);
nand U38701 (N_38701,N_37528,N_37845);
or U38702 (N_38702,N_37542,N_36363);
and U38703 (N_38703,N_37448,N_36859);
nor U38704 (N_38704,N_36314,N_37974);
nand U38705 (N_38705,N_36982,N_37519);
xnor U38706 (N_38706,N_37086,N_36493);
nor U38707 (N_38707,N_37135,N_37121);
or U38708 (N_38708,N_36498,N_36598);
or U38709 (N_38709,N_36581,N_37360);
nand U38710 (N_38710,N_37254,N_37223);
or U38711 (N_38711,N_36713,N_36502);
and U38712 (N_38712,N_37188,N_36440);
and U38713 (N_38713,N_36991,N_37675);
nor U38714 (N_38714,N_36791,N_37044);
xor U38715 (N_38715,N_36679,N_37544);
xnor U38716 (N_38716,N_37496,N_36722);
nor U38717 (N_38717,N_37532,N_37829);
xor U38718 (N_38718,N_36781,N_37814);
xnor U38719 (N_38719,N_37395,N_37051);
nor U38720 (N_38720,N_37492,N_36342);
xnor U38721 (N_38721,N_36069,N_37080);
or U38722 (N_38722,N_37299,N_37961);
nor U38723 (N_38723,N_37291,N_37484);
or U38724 (N_38724,N_37129,N_36169);
nor U38725 (N_38725,N_37453,N_37514);
nor U38726 (N_38726,N_36189,N_36954);
or U38727 (N_38727,N_36666,N_36464);
and U38728 (N_38728,N_36212,N_37543);
or U38729 (N_38729,N_36961,N_37460);
nor U38730 (N_38730,N_37226,N_36586);
nor U38731 (N_38731,N_36597,N_36492);
or U38732 (N_38732,N_37538,N_37552);
or U38733 (N_38733,N_36883,N_36381);
xor U38734 (N_38734,N_37052,N_37417);
nand U38735 (N_38735,N_37699,N_37900);
nand U38736 (N_38736,N_36603,N_37850);
nand U38737 (N_38737,N_37836,N_37564);
nor U38738 (N_38738,N_36798,N_36495);
xor U38739 (N_38739,N_36686,N_36906);
and U38740 (N_38740,N_36817,N_37340);
xor U38741 (N_38741,N_37187,N_37237);
nor U38742 (N_38742,N_37367,N_37139);
nor U38743 (N_38743,N_36167,N_36912);
or U38744 (N_38744,N_37073,N_36199);
or U38745 (N_38745,N_36332,N_37969);
nand U38746 (N_38746,N_36434,N_36159);
nor U38747 (N_38747,N_36170,N_37343);
nor U38748 (N_38748,N_37508,N_36589);
or U38749 (N_38749,N_36778,N_36500);
and U38750 (N_38750,N_36038,N_37031);
nand U38751 (N_38751,N_36397,N_37333);
nand U38752 (N_38752,N_36302,N_37463);
nor U38753 (N_38753,N_37192,N_36885);
xnor U38754 (N_38754,N_36710,N_37116);
nor U38755 (N_38755,N_37647,N_37481);
nand U38756 (N_38756,N_36295,N_36318);
nand U38757 (N_38757,N_37714,N_36039);
nand U38758 (N_38758,N_37489,N_36524);
xnor U38759 (N_38759,N_36055,N_37043);
xnor U38760 (N_38760,N_37131,N_36380);
nor U38761 (N_38761,N_36426,N_36698);
xor U38762 (N_38762,N_37058,N_36733);
nor U38763 (N_38763,N_36149,N_37713);
nor U38764 (N_38764,N_36941,N_36560);
and U38765 (N_38765,N_36630,N_36119);
xor U38766 (N_38766,N_37279,N_37786);
or U38767 (N_38767,N_36338,N_37325);
nand U38768 (N_38768,N_37249,N_37813);
nand U38769 (N_38769,N_36358,N_37132);
or U38770 (N_38770,N_37886,N_36824);
and U38771 (N_38771,N_36225,N_36155);
xnor U38772 (N_38772,N_37741,N_36992);
nor U38773 (N_38773,N_37025,N_37577);
and U38774 (N_38774,N_37710,N_36715);
or U38775 (N_38775,N_37902,N_37454);
nor U38776 (N_38776,N_37930,N_36256);
nand U38777 (N_38777,N_36205,N_36056);
xnor U38778 (N_38778,N_37252,N_37096);
nand U38779 (N_38779,N_37104,N_36550);
nor U38780 (N_38780,N_36281,N_37731);
and U38781 (N_38781,N_37650,N_36465);
or U38782 (N_38782,N_37662,N_37745);
or U38783 (N_38783,N_36271,N_36816);
xnor U38784 (N_38784,N_37041,N_37576);
xnor U38785 (N_38785,N_37170,N_37896);
or U38786 (N_38786,N_36979,N_36542);
xor U38787 (N_38787,N_37335,N_36582);
nand U38788 (N_38788,N_37584,N_37065);
nor U38789 (N_38789,N_37437,N_36972);
nand U38790 (N_38790,N_37286,N_37653);
and U38791 (N_38791,N_37109,N_37415);
nor U38792 (N_38792,N_37019,N_37855);
and U38793 (N_38793,N_36079,N_36458);
and U38794 (N_38794,N_36070,N_36202);
and U38795 (N_38795,N_36127,N_36966);
nand U38796 (N_38796,N_37689,N_36313);
xnor U38797 (N_38797,N_36813,N_36266);
nor U38798 (N_38798,N_37022,N_36388);
nand U38799 (N_38799,N_37148,N_36516);
and U38800 (N_38800,N_36081,N_37127);
nand U38801 (N_38801,N_37385,N_37962);
and U38802 (N_38802,N_36300,N_36568);
xor U38803 (N_38803,N_37295,N_36274);
nor U38804 (N_38804,N_37029,N_36385);
and U38805 (N_38805,N_36964,N_36579);
nand U38806 (N_38806,N_36287,N_37794);
nor U38807 (N_38807,N_36761,N_37599);
xor U38808 (N_38808,N_37616,N_37843);
or U38809 (N_38809,N_36120,N_37003);
nor U38810 (N_38810,N_36087,N_37605);
nand U38811 (N_38811,N_37865,N_37027);
xnor U38812 (N_38812,N_36995,N_37968);
or U38813 (N_38813,N_37054,N_37718);
and U38814 (N_38814,N_36187,N_36847);
nand U38815 (N_38815,N_36759,N_36308);
nor U38816 (N_38816,N_37738,N_37554);
and U38817 (N_38817,N_36010,N_37685);
and U38818 (N_38818,N_37196,N_37013);
nand U38819 (N_38819,N_37559,N_37931);
nand U38820 (N_38820,N_37245,N_36037);
nand U38821 (N_38821,N_37608,N_37770);
nand U38822 (N_38822,N_37077,N_37298);
nor U38823 (N_38823,N_36865,N_36680);
nand U38824 (N_38824,N_37304,N_36419);
xor U38825 (N_38825,N_37100,N_37374);
or U38826 (N_38826,N_36697,N_37954);
and U38827 (N_38827,N_37530,N_36572);
xnor U38828 (N_38828,N_36882,N_36304);
and U38829 (N_38829,N_36269,N_36230);
and U38830 (N_38830,N_37097,N_37512);
xnor U38831 (N_38831,N_36782,N_36670);
nand U38832 (N_38832,N_37218,N_36262);
xor U38833 (N_38833,N_37533,N_36708);
and U38834 (N_38834,N_36705,N_36553);
or U38835 (N_38835,N_36745,N_37849);
and U38836 (N_38836,N_36997,N_36786);
nor U38837 (N_38837,N_37848,N_36642);
or U38838 (N_38838,N_37574,N_37275);
and U38839 (N_38839,N_37612,N_37995);
and U38840 (N_38840,N_36430,N_36369);
or U38841 (N_38841,N_36766,N_36924);
or U38842 (N_38842,N_37225,N_36372);
nand U38843 (N_38843,N_36874,N_37400);
xnor U38844 (N_38844,N_36831,N_37771);
or U38845 (N_38845,N_36168,N_37536);
and U38846 (N_38846,N_37443,N_37341);
or U38847 (N_38847,N_37521,N_36333);
xor U38848 (N_38848,N_36875,N_37697);
xor U38849 (N_38849,N_37085,N_37255);
or U38850 (N_38850,N_36775,N_36216);
xnor U38851 (N_38851,N_37958,N_36192);
or U38852 (N_38852,N_36378,N_37703);
or U38853 (N_38853,N_37217,N_37847);
or U38854 (N_38854,N_37815,N_37687);
nand U38855 (N_38855,N_37361,N_37876);
xor U38856 (N_38856,N_37447,N_37832);
and U38857 (N_38857,N_37222,N_36867);
nand U38858 (N_38858,N_37036,N_36537);
nand U38859 (N_38859,N_37243,N_37107);
or U38860 (N_38860,N_36355,N_37746);
or U38861 (N_38861,N_37277,N_36925);
xnor U38862 (N_38862,N_37549,N_36336);
nor U38863 (N_38863,N_37712,N_37421);
and U38864 (N_38864,N_37119,N_37688);
nor U38865 (N_38865,N_36238,N_36402);
xnor U38866 (N_38866,N_36609,N_36724);
and U38867 (N_38867,N_37875,N_36805);
or U38868 (N_38868,N_37456,N_37772);
or U38869 (N_38869,N_36639,N_36178);
and U38870 (N_38870,N_37920,N_37717);
xnor U38871 (N_38871,N_37263,N_37730);
xnor U38872 (N_38872,N_36857,N_36506);
or U38873 (N_38873,N_37462,N_36340);
or U38874 (N_38874,N_37922,N_37762);
nand U38875 (N_38875,N_37440,N_37305);
nor U38876 (N_38876,N_37992,N_36562);
nand U38877 (N_38877,N_36396,N_36280);
nor U38878 (N_38878,N_36640,N_37693);
and U38879 (N_38879,N_36593,N_37830);
and U38880 (N_38880,N_36613,N_36703);
or U38881 (N_38881,N_37191,N_37680);
nor U38882 (N_38882,N_36902,N_37497);
nand U38883 (N_38883,N_37201,N_36117);
nand U38884 (N_38884,N_37040,N_37872);
nand U38885 (N_38885,N_36554,N_37802);
and U38886 (N_38886,N_37112,N_37804);
xnor U38887 (N_38887,N_37915,N_36970);
or U38888 (N_38888,N_37345,N_36704);
or U38889 (N_38889,N_36989,N_37370);
nor U38890 (N_38890,N_36968,N_36382);
nand U38891 (N_38891,N_37701,N_36311);
xor U38892 (N_38892,N_36548,N_36852);
nand U38893 (N_38893,N_37588,N_37888);
and U38894 (N_38894,N_36221,N_37656);
and U38895 (N_38895,N_36356,N_37925);
nand U38896 (N_38896,N_36750,N_36566);
nand U38897 (N_38897,N_36916,N_37200);
or U38898 (N_38898,N_37402,N_36400);
xor U38899 (N_38899,N_36702,N_37898);
xnor U38900 (N_38900,N_37451,N_37798);
or U38901 (N_38901,N_36547,N_36228);
nand U38902 (N_38902,N_36898,N_36215);
nand U38903 (N_38903,N_37618,N_36193);
nand U38904 (N_38904,N_36540,N_37398);
xor U38905 (N_38905,N_36588,N_37262);
nor U38906 (N_38906,N_37126,N_36590);
or U38907 (N_38907,N_37273,N_36208);
xor U38908 (N_38908,N_37175,N_37645);
nor U38909 (N_38909,N_36627,N_36525);
or U38910 (N_38910,N_36523,N_37825);
nor U38911 (N_38911,N_36856,N_37161);
nor U38912 (N_38912,N_36661,N_36645);
nand U38913 (N_38913,N_36737,N_37224);
nand U38914 (N_38914,N_37087,N_37248);
and U38915 (N_38915,N_37904,N_37719);
and U38916 (N_38916,N_37012,N_36061);
nand U38917 (N_38917,N_37614,N_36683);
and U38918 (N_38918,N_37932,N_36445);
xnor U38919 (N_38919,N_36443,N_36398);
xnor U38920 (N_38920,N_36812,N_37568);
nor U38921 (N_38921,N_37137,N_36729);
nor U38922 (N_38922,N_36734,N_37778);
nor U38923 (N_38923,N_37858,N_37960);
and U38924 (N_38924,N_37801,N_36251);
or U38925 (N_38925,N_36950,N_37842);
xor U38926 (N_38926,N_36773,N_36743);
xnor U38927 (N_38927,N_37049,N_37493);
and U38928 (N_38928,N_37330,N_36531);
or U38929 (N_38929,N_36533,N_36792);
and U38930 (N_38930,N_36416,N_36716);
or U38931 (N_38931,N_36103,N_36427);
or U38932 (N_38932,N_37477,N_36386);
xnor U38933 (N_38933,N_37034,N_37972);
nand U38934 (N_38934,N_37800,N_36881);
xnor U38935 (N_38935,N_36815,N_37449);
and U38936 (N_38936,N_36850,N_36935);
and U38937 (N_38937,N_37480,N_36360);
nor U38938 (N_38938,N_37315,N_36469);
and U38939 (N_38939,N_36219,N_37905);
xnor U38940 (N_38940,N_36217,N_36334);
or U38941 (N_38941,N_37889,N_37424);
and U38942 (N_38942,N_36049,N_36359);
nor U38943 (N_38943,N_37562,N_37024);
and U38944 (N_38944,N_36052,N_36983);
or U38945 (N_38945,N_37381,N_37234);
nor U38946 (N_38946,N_36485,N_36920);
nand U38947 (N_38947,N_36662,N_37692);
xor U38948 (N_38948,N_37046,N_37926);
and U38949 (N_38949,N_36578,N_37072);
nand U38950 (N_38950,N_37923,N_37502);
and U38951 (N_38951,N_36963,N_37700);
or U38952 (N_38952,N_36942,N_36610);
nand U38953 (N_38953,N_36718,N_36329);
and U38954 (N_38954,N_37945,N_36501);
xnor U38955 (N_38955,N_36570,N_37035);
or U38956 (N_38956,N_37383,N_37996);
or U38957 (N_38957,N_36829,N_36688);
or U38958 (N_38958,N_37658,N_36243);
xnor U38959 (N_38959,N_37628,N_36001);
xnor U38960 (N_38960,N_36031,N_37488);
or U38961 (N_38961,N_36741,N_36133);
and U38962 (N_38962,N_36522,N_37823);
or U38963 (N_38963,N_37882,N_36341);
xor U38964 (N_38964,N_37953,N_37775);
and U38965 (N_38965,N_36535,N_36144);
and U38966 (N_38966,N_36594,N_36414);
or U38967 (N_38967,N_37773,N_36809);
xor U38968 (N_38968,N_37835,N_37071);
xor U38969 (N_38969,N_36390,N_37278);
and U38970 (N_38970,N_37740,N_36915);
and U38971 (N_38971,N_36700,N_37230);
xor U38972 (N_38972,N_36054,N_36030);
nor U38973 (N_38973,N_36918,N_36930);
and U38974 (N_38974,N_37408,N_37152);
or U38975 (N_38975,N_36672,N_37971);
and U38976 (N_38976,N_37185,N_37641);
xor U38977 (N_38977,N_37336,N_36981);
and U38978 (N_38978,N_37260,N_37233);
or U38979 (N_38979,N_36004,N_36245);
xnor U38980 (N_38980,N_37114,N_37423);
nand U38981 (N_38981,N_37897,N_36633);
or U38982 (N_38982,N_36858,N_36022);
or U38983 (N_38983,N_36987,N_37216);
or U38984 (N_38984,N_36299,N_37744);
or U38985 (N_38985,N_36894,N_36814);
and U38986 (N_38986,N_36000,N_37728);
or U38987 (N_38987,N_36074,N_37660);
nand U38988 (N_38988,N_37817,N_37633);
nor U38989 (N_38989,N_36446,N_36122);
or U38990 (N_38990,N_36556,N_37671);
nand U38991 (N_38991,N_36677,N_36150);
and U38992 (N_38992,N_36635,N_36487);
nand U38993 (N_38993,N_37525,N_36605);
nor U38994 (N_38994,N_37994,N_37742);
xnor U38995 (N_38995,N_37123,N_37610);
or U38996 (N_38996,N_37792,N_36098);
nand U38997 (N_38997,N_36327,N_37822);
nand U38998 (N_38998,N_36162,N_37698);
xnor U38999 (N_38999,N_37604,N_37392);
nand U39000 (N_39000,N_36135,N_37290);
and U39001 (N_39001,N_37686,N_37675);
nand U39002 (N_39002,N_37600,N_37812);
nor U39003 (N_39003,N_37707,N_37376);
xnor U39004 (N_39004,N_36479,N_36032);
xnor U39005 (N_39005,N_37615,N_37753);
and U39006 (N_39006,N_37964,N_37590);
nand U39007 (N_39007,N_36071,N_36717);
nand U39008 (N_39008,N_37255,N_37448);
nor U39009 (N_39009,N_36126,N_36808);
xor U39010 (N_39010,N_36314,N_37595);
xnor U39011 (N_39011,N_37546,N_36633);
or U39012 (N_39012,N_36053,N_36397);
or U39013 (N_39013,N_37655,N_37728);
nand U39014 (N_39014,N_36087,N_37898);
nor U39015 (N_39015,N_37428,N_36998);
and U39016 (N_39016,N_37173,N_37333);
xnor U39017 (N_39017,N_36119,N_36015);
or U39018 (N_39018,N_37726,N_37340);
nor U39019 (N_39019,N_36479,N_37225);
or U39020 (N_39020,N_36394,N_37307);
xnor U39021 (N_39021,N_36342,N_36965);
or U39022 (N_39022,N_37774,N_37956);
xnor U39023 (N_39023,N_36011,N_36877);
or U39024 (N_39024,N_37285,N_36261);
xor U39025 (N_39025,N_37323,N_36049);
or U39026 (N_39026,N_37638,N_37910);
and U39027 (N_39027,N_36956,N_36692);
and U39028 (N_39028,N_37299,N_36408);
nor U39029 (N_39029,N_37350,N_37426);
and U39030 (N_39030,N_36349,N_36718);
nor U39031 (N_39031,N_37232,N_36911);
or U39032 (N_39032,N_37776,N_37523);
xor U39033 (N_39033,N_36603,N_37256);
and U39034 (N_39034,N_36644,N_36899);
nand U39035 (N_39035,N_36398,N_37413);
nor U39036 (N_39036,N_36167,N_37956);
nor U39037 (N_39037,N_36309,N_37255);
nor U39038 (N_39038,N_37770,N_37350);
nor U39039 (N_39039,N_37217,N_36531);
xor U39040 (N_39040,N_37955,N_36617);
nand U39041 (N_39041,N_37946,N_36543);
or U39042 (N_39042,N_36137,N_36746);
nor U39043 (N_39043,N_36230,N_36834);
and U39044 (N_39044,N_36171,N_36911);
xnor U39045 (N_39045,N_36683,N_37956);
nor U39046 (N_39046,N_37705,N_37568);
and U39047 (N_39047,N_37698,N_37106);
nor U39048 (N_39048,N_36722,N_36749);
xor U39049 (N_39049,N_37664,N_36214);
xor U39050 (N_39050,N_37625,N_36535);
or U39051 (N_39051,N_36099,N_37434);
or U39052 (N_39052,N_36402,N_36098);
nand U39053 (N_39053,N_36343,N_36467);
nor U39054 (N_39054,N_36354,N_36187);
or U39055 (N_39055,N_37340,N_37730);
or U39056 (N_39056,N_36702,N_36343);
xor U39057 (N_39057,N_37362,N_37674);
and U39058 (N_39058,N_36229,N_37972);
nor U39059 (N_39059,N_37424,N_37248);
and U39060 (N_39060,N_37402,N_37982);
nor U39061 (N_39061,N_36823,N_37602);
or U39062 (N_39062,N_36343,N_37704);
xnor U39063 (N_39063,N_37782,N_37097);
xor U39064 (N_39064,N_37681,N_36571);
or U39065 (N_39065,N_36078,N_36074);
xnor U39066 (N_39066,N_37322,N_37420);
nor U39067 (N_39067,N_36077,N_36440);
nor U39068 (N_39068,N_37408,N_37529);
or U39069 (N_39069,N_36837,N_37913);
xnor U39070 (N_39070,N_37134,N_37013);
nor U39071 (N_39071,N_36854,N_37610);
nor U39072 (N_39072,N_36725,N_36445);
or U39073 (N_39073,N_37389,N_37092);
and U39074 (N_39074,N_36014,N_36066);
and U39075 (N_39075,N_36346,N_36950);
or U39076 (N_39076,N_36510,N_36613);
and U39077 (N_39077,N_37567,N_37401);
nor U39078 (N_39078,N_37507,N_36454);
or U39079 (N_39079,N_36829,N_36015);
nand U39080 (N_39080,N_37405,N_37423);
and U39081 (N_39081,N_37255,N_37482);
xor U39082 (N_39082,N_37196,N_36620);
and U39083 (N_39083,N_36426,N_37571);
or U39084 (N_39084,N_37537,N_36763);
nor U39085 (N_39085,N_36238,N_36650);
xnor U39086 (N_39086,N_37643,N_36672);
or U39087 (N_39087,N_37856,N_36312);
or U39088 (N_39088,N_36390,N_37820);
or U39089 (N_39089,N_37402,N_37812);
nor U39090 (N_39090,N_37953,N_36436);
nor U39091 (N_39091,N_36159,N_36148);
nor U39092 (N_39092,N_36011,N_37853);
xnor U39093 (N_39093,N_37881,N_36495);
or U39094 (N_39094,N_37361,N_36976);
xnor U39095 (N_39095,N_36720,N_37985);
xnor U39096 (N_39096,N_37402,N_36568);
nor U39097 (N_39097,N_36161,N_36180);
or U39098 (N_39098,N_36565,N_37803);
nand U39099 (N_39099,N_36420,N_36327);
or U39100 (N_39100,N_36108,N_36608);
nor U39101 (N_39101,N_37866,N_36417);
nand U39102 (N_39102,N_36173,N_37110);
and U39103 (N_39103,N_37331,N_37663);
xor U39104 (N_39104,N_37721,N_36641);
nand U39105 (N_39105,N_37047,N_36345);
xnor U39106 (N_39106,N_36952,N_36572);
or U39107 (N_39107,N_37862,N_37303);
and U39108 (N_39108,N_36315,N_36269);
xor U39109 (N_39109,N_36544,N_37305);
and U39110 (N_39110,N_37036,N_36812);
xnor U39111 (N_39111,N_37481,N_37056);
and U39112 (N_39112,N_37242,N_37788);
or U39113 (N_39113,N_37524,N_37325);
and U39114 (N_39114,N_36328,N_36579);
or U39115 (N_39115,N_36439,N_37891);
or U39116 (N_39116,N_37324,N_36952);
and U39117 (N_39117,N_37331,N_37327);
or U39118 (N_39118,N_36271,N_36286);
or U39119 (N_39119,N_36016,N_36997);
and U39120 (N_39120,N_37338,N_37551);
xor U39121 (N_39121,N_36049,N_37547);
nand U39122 (N_39122,N_37383,N_36584);
nand U39123 (N_39123,N_37505,N_37221);
nor U39124 (N_39124,N_36568,N_36317);
xor U39125 (N_39125,N_36837,N_36036);
or U39126 (N_39126,N_36493,N_37737);
nand U39127 (N_39127,N_36732,N_36256);
and U39128 (N_39128,N_37517,N_36607);
xnor U39129 (N_39129,N_36141,N_37483);
and U39130 (N_39130,N_37311,N_37202);
nor U39131 (N_39131,N_37668,N_36427);
or U39132 (N_39132,N_36471,N_37371);
xor U39133 (N_39133,N_36153,N_36525);
or U39134 (N_39134,N_37756,N_37383);
and U39135 (N_39135,N_37278,N_36833);
nand U39136 (N_39136,N_37452,N_36214);
and U39137 (N_39137,N_37970,N_37554);
nand U39138 (N_39138,N_37149,N_37073);
and U39139 (N_39139,N_37617,N_36361);
nor U39140 (N_39140,N_37451,N_37981);
nand U39141 (N_39141,N_36086,N_37502);
nand U39142 (N_39142,N_37744,N_37867);
nand U39143 (N_39143,N_36733,N_36411);
nand U39144 (N_39144,N_37588,N_37643);
or U39145 (N_39145,N_36851,N_37097);
nor U39146 (N_39146,N_36493,N_36300);
or U39147 (N_39147,N_36086,N_37315);
nor U39148 (N_39148,N_36455,N_36223);
nand U39149 (N_39149,N_37518,N_37349);
nor U39150 (N_39150,N_36322,N_37669);
xnor U39151 (N_39151,N_36548,N_36721);
nor U39152 (N_39152,N_37824,N_37619);
or U39153 (N_39153,N_36783,N_37964);
nand U39154 (N_39154,N_36901,N_37681);
nor U39155 (N_39155,N_37697,N_36981);
nor U39156 (N_39156,N_36574,N_37789);
nand U39157 (N_39157,N_36826,N_36870);
and U39158 (N_39158,N_36650,N_36085);
nor U39159 (N_39159,N_37136,N_36493);
nor U39160 (N_39160,N_36543,N_37150);
xnor U39161 (N_39161,N_36229,N_37008);
nand U39162 (N_39162,N_36125,N_36932);
nand U39163 (N_39163,N_37324,N_36464);
or U39164 (N_39164,N_36552,N_37642);
xor U39165 (N_39165,N_37725,N_37333);
and U39166 (N_39166,N_37814,N_36369);
xor U39167 (N_39167,N_36982,N_36343);
nor U39168 (N_39168,N_37520,N_36890);
and U39169 (N_39169,N_36469,N_37852);
and U39170 (N_39170,N_36807,N_36934);
and U39171 (N_39171,N_36999,N_37518);
xor U39172 (N_39172,N_36204,N_36143);
nand U39173 (N_39173,N_37501,N_36556);
nand U39174 (N_39174,N_36549,N_37061);
nand U39175 (N_39175,N_36417,N_37285);
xor U39176 (N_39176,N_36533,N_36523);
nand U39177 (N_39177,N_36948,N_37650);
nor U39178 (N_39178,N_37320,N_36418);
xnor U39179 (N_39179,N_36918,N_37892);
xnor U39180 (N_39180,N_36542,N_37187);
nand U39181 (N_39181,N_37991,N_37696);
nor U39182 (N_39182,N_36694,N_37094);
nand U39183 (N_39183,N_36035,N_36517);
xor U39184 (N_39184,N_37004,N_36346);
and U39185 (N_39185,N_36882,N_37742);
nor U39186 (N_39186,N_37368,N_36623);
xnor U39187 (N_39187,N_36513,N_37749);
and U39188 (N_39188,N_37445,N_36735);
and U39189 (N_39189,N_37197,N_36944);
or U39190 (N_39190,N_37826,N_36107);
or U39191 (N_39191,N_37075,N_36047);
and U39192 (N_39192,N_36045,N_36333);
or U39193 (N_39193,N_36025,N_36621);
and U39194 (N_39194,N_36912,N_37137);
xor U39195 (N_39195,N_37958,N_37138);
nand U39196 (N_39196,N_37320,N_36171);
nand U39197 (N_39197,N_37935,N_37954);
or U39198 (N_39198,N_37190,N_36620);
nor U39199 (N_39199,N_36602,N_37065);
and U39200 (N_39200,N_37315,N_36869);
and U39201 (N_39201,N_36123,N_36024);
nand U39202 (N_39202,N_36354,N_37362);
nor U39203 (N_39203,N_37539,N_37826);
nand U39204 (N_39204,N_37335,N_37512);
xnor U39205 (N_39205,N_36490,N_36684);
or U39206 (N_39206,N_36612,N_37978);
nor U39207 (N_39207,N_36508,N_37118);
and U39208 (N_39208,N_37363,N_36669);
or U39209 (N_39209,N_36863,N_36480);
nand U39210 (N_39210,N_37785,N_37275);
nand U39211 (N_39211,N_37603,N_36220);
nand U39212 (N_39212,N_36969,N_36716);
or U39213 (N_39213,N_37407,N_36016);
or U39214 (N_39214,N_36720,N_36694);
and U39215 (N_39215,N_37263,N_36672);
xor U39216 (N_39216,N_37173,N_36428);
or U39217 (N_39217,N_36559,N_37766);
or U39218 (N_39218,N_36514,N_36170);
or U39219 (N_39219,N_37441,N_36676);
or U39220 (N_39220,N_36881,N_36709);
or U39221 (N_39221,N_36828,N_37063);
and U39222 (N_39222,N_37777,N_36030);
and U39223 (N_39223,N_37101,N_36270);
nor U39224 (N_39224,N_37714,N_37651);
nand U39225 (N_39225,N_37755,N_37939);
and U39226 (N_39226,N_36208,N_37802);
xor U39227 (N_39227,N_37124,N_36456);
and U39228 (N_39228,N_37768,N_37335);
or U39229 (N_39229,N_36549,N_36332);
and U39230 (N_39230,N_36608,N_37887);
nand U39231 (N_39231,N_36660,N_36453);
nand U39232 (N_39232,N_36682,N_36913);
or U39233 (N_39233,N_36569,N_36650);
or U39234 (N_39234,N_37854,N_36347);
or U39235 (N_39235,N_37238,N_37995);
nand U39236 (N_39236,N_36700,N_37168);
nor U39237 (N_39237,N_36605,N_36724);
xor U39238 (N_39238,N_37892,N_37102);
xor U39239 (N_39239,N_37586,N_36769);
or U39240 (N_39240,N_37666,N_37263);
nor U39241 (N_39241,N_37218,N_37729);
or U39242 (N_39242,N_37087,N_37053);
and U39243 (N_39243,N_37196,N_37925);
nand U39244 (N_39244,N_37232,N_36684);
or U39245 (N_39245,N_36137,N_36975);
xnor U39246 (N_39246,N_36369,N_37067);
xor U39247 (N_39247,N_36478,N_36011);
nand U39248 (N_39248,N_36611,N_36025);
nor U39249 (N_39249,N_37265,N_36561);
nand U39250 (N_39250,N_36118,N_37778);
and U39251 (N_39251,N_36898,N_36876);
nor U39252 (N_39252,N_37668,N_37920);
nor U39253 (N_39253,N_36595,N_37902);
nor U39254 (N_39254,N_36065,N_36719);
nor U39255 (N_39255,N_37913,N_36853);
or U39256 (N_39256,N_37742,N_36137);
and U39257 (N_39257,N_36490,N_37811);
nor U39258 (N_39258,N_37991,N_36140);
or U39259 (N_39259,N_36336,N_36537);
nand U39260 (N_39260,N_37962,N_37485);
and U39261 (N_39261,N_37760,N_36314);
nor U39262 (N_39262,N_37053,N_36864);
nor U39263 (N_39263,N_37035,N_37779);
nand U39264 (N_39264,N_37647,N_36248);
xnor U39265 (N_39265,N_37643,N_36929);
and U39266 (N_39266,N_36309,N_36561);
or U39267 (N_39267,N_36838,N_36915);
xor U39268 (N_39268,N_36592,N_37285);
and U39269 (N_39269,N_36801,N_37974);
xnor U39270 (N_39270,N_37927,N_37036);
nand U39271 (N_39271,N_37925,N_36046);
and U39272 (N_39272,N_36243,N_37216);
and U39273 (N_39273,N_36122,N_37985);
nand U39274 (N_39274,N_36723,N_37037);
nand U39275 (N_39275,N_37154,N_37128);
xnor U39276 (N_39276,N_36681,N_36503);
or U39277 (N_39277,N_37659,N_36922);
xor U39278 (N_39278,N_36949,N_36446);
nor U39279 (N_39279,N_36588,N_36460);
or U39280 (N_39280,N_37700,N_37216);
nand U39281 (N_39281,N_36790,N_37692);
nand U39282 (N_39282,N_37527,N_36996);
and U39283 (N_39283,N_37051,N_37638);
xnor U39284 (N_39284,N_37797,N_37848);
nor U39285 (N_39285,N_37507,N_37349);
nand U39286 (N_39286,N_36708,N_37534);
and U39287 (N_39287,N_36973,N_37924);
nor U39288 (N_39288,N_36943,N_36813);
nand U39289 (N_39289,N_36626,N_36285);
and U39290 (N_39290,N_37280,N_36505);
or U39291 (N_39291,N_36623,N_36140);
xnor U39292 (N_39292,N_37683,N_37740);
xnor U39293 (N_39293,N_36645,N_36743);
nand U39294 (N_39294,N_37938,N_36164);
nor U39295 (N_39295,N_36727,N_37921);
nand U39296 (N_39296,N_36033,N_37386);
xnor U39297 (N_39297,N_37649,N_37991);
nor U39298 (N_39298,N_36182,N_37565);
nor U39299 (N_39299,N_37116,N_36390);
nand U39300 (N_39300,N_37458,N_37864);
nand U39301 (N_39301,N_36355,N_36196);
or U39302 (N_39302,N_36759,N_37696);
xnor U39303 (N_39303,N_36232,N_37959);
xnor U39304 (N_39304,N_37580,N_37104);
or U39305 (N_39305,N_36586,N_37169);
nor U39306 (N_39306,N_37347,N_37149);
nand U39307 (N_39307,N_36807,N_37085);
or U39308 (N_39308,N_37135,N_36315);
nand U39309 (N_39309,N_37086,N_36697);
nor U39310 (N_39310,N_36038,N_36892);
nand U39311 (N_39311,N_36148,N_37157);
nor U39312 (N_39312,N_37133,N_36150);
nand U39313 (N_39313,N_36769,N_37142);
nand U39314 (N_39314,N_36624,N_37078);
or U39315 (N_39315,N_37278,N_37016);
and U39316 (N_39316,N_37477,N_37333);
xor U39317 (N_39317,N_36941,N_36381);
nor U39318 (N_39318,N_37460,N_37252);
and U39319 (N_39319,N_36666,N_37707);
xor U39320 (N_39320,N_36205,N_37587);
xnor U39321 (N_39321,N_37959,N_37706);
nand U39322 (N_39322,N_36862,N_37586);
xor U39323 (N_39323,N_37570,N_37130);
nand U39324 (N_39324,N_37150,N_36468);
xnor U39325 (N_39325,N_37173,N_37331);
nand U39326 (N_39326,N_37382,N_37124);
nor U39327 (N_39327,N_37929,N_36826);
nand U39328 (N_39328,N_37406,N_36005);
or U39329 (N_39329,N_37586,N_36753);
or U39330 (N_39330,N_37467,N_36258);
xor U39331 (N_39331,N_36937,N_37063);
or U39332 (N_39332,N_36960,N_37133);
nand U39333 (N_39333,N_37215,N_36493);
nand U39334 (N_39334,N_36574,N_36025);
or U39335 (N_39335,N_37328,N_36780);
nor U39336 (N_39336,N_36608,N_37269);
or U39337 (N_39337,N_36496,N_36563);
nand U39338 (N_39338,N_36849,N_36855);
nand U39339 (N_39339,N_37317,N_37332);
and U39340 (N_39340,N_36102,N_37349);
nor U39341 (N_39341,N_37016,N_36374);
xnor U39342 (N_39342,N_36466,N_36173);
nor U39343 (N_39343,N_37440,N_36717);
nor U39344 (N_39344,N_36863,N_37747);
or U39345 (N_39345,N_37101,N_36145);
or U39346 (N_39346,N_36395,N_36190);
xor U39347 (N_39347,N_36681,N_37776);
or U39348 (N_39348,N_36278,N_37958);
and U39349 (N_39349,N_37440,N_37964);
xnor U39350 (N_39350,N_37320,N_36702);
nand U39351 (N_39351,N_37835,N_36837);
nand U39352 (N_39352,N_37609,N_36109);
xor U39353 (N_39353,N_37625,N_36071);
xnor U39354 (N_39354,N_37746,N_36968);
nor U39355 (N_39355,N_37948,N_36017);
nand U39356 (N_39356,N_37042,N_37060);
and U39357 (N_39357,N_36649,N_37526);
nand U39358 (N_39358,N_36441,N_37069);
nor U39359 (N_39359,N_36498,N_37319);
or U39360 (N_39360,N_36185,N_36343);
nand U39361 (N_39361,N_37130,N_36234);
and U39362 (N_39362,N_37395,N_36209);
nor U39363 (N_39363,N_36789,N_37114);
nor U39364 (N_39364,N_37293,N_36782);
xnor U39365 (N_39365,N_36794,N_36183);
and U39366 (N_39366,N_37642,N_36922);
xor U39367 (N_39367,N_36796,N_37675);
or U39368 (N_39368,N_37540,N_36729);
or U39369 (N_39369,N_37267,N_36164);
nor U39370 (N_39370,N_36310,N_36493);
nor U39371 (N_39371,N_37107,N_36365);
nor U39372 (N_39372,N_36462,N_37126);
and U39373 (N_39373,N_36190,N_37995);
or U39374 (N_39374,N_36007,N_36657);
nand U39375 (N_39375,N_37806,N_36289);
nor U39376 (N_39376,N_36297,N_36249);
nor U39377 (N_39377,N_36820,N_36987);
or U39378 (N_39378,N_36503,N_36841);
and U39379 (N_39379,N_36970,N_37927);
nor U39380 (N_39380,N_37001,N_36215);
and U39381 (N_39381,N_37859,N_37434);
nand U39382 (N_39382,N_37005,N_36937);
and U39383 (N_39383,N_36759,N_36914);
and U39384 (N_39384,N_36426,N_36673);
xor U39385 (N_39385,N_36649,N_37392);
nor U39386 (N_39386,N_37261,N_36213);
and U39387 (N_39387,N_37629,N_36927);
nand U39388 (N_39388,N_36412,N_37948);
and U39389 (N_39389,N_36345,N_37511);
xor U39390 (N_39390,N_37613,N_37557);
nand U39391 (N_39391,N_37153,N_36373);
or U39392 (N_39392,N_37766,N_36913);
nand U39393 (N_39393,N_37493,N_36642);
xnor U39394 (N_39394,N_36080,N_37406);
xor U39395 (N_39395,N_36895,N_37660);
nand U39396 (N_39396,N_36868,N_36949);
nor U39397 (N_39397,N_37017,N_37223);
and U39398 (N_39398,N_36903,N_36307);
nor U39399 (N_39399,N_36482,N_36495);
and U39400 (N_39400,N_36555,N_36630);
and U39401 (N_39401,N_37030,N_37520);
or U39402 (N_39402,N_37158,N_37508);
or U39403 (N_39403,N_37170,N_37962);
nor U39404 (N_39404,N_37278,N_36373);
nor U39405 (N_39405,N_37539,N_37521);
nand U39406 (N_39406,N_37518,N_37857);
or U39407 (N_39407,N_37446,N_36525);
nor U39408 (N_39408,N_36237,N_36590);
or U39409 (N_39409,N_36986,N_36950);
nand U39410 (N_39410,N_36846,N_36922);
nand U39411 (N_39411,N_37295,N_36046);
xor U39412 (N_39412,N_36409,N_36922);
nor U39413 (N_39413,N_37978,N_37666);
nand U39414 (N_39414,N_37120,N_37476);
and U39415 (N_39415,N_37062,N_37572);
xor U39416 (N_39416,N_37360,N_37476);
xor U39417 (N_39417,N_37886,N_37046);
or U39418 (N_39418,N_36551,N_36575);
and U39419 (N_39419,N_37075,N_37045);
nor U39420 (N_39420,N_36363,N_36173);
nand U39421 (N_39421,N_37644,N_36934);
nand U39422 (N_39422,N_37319,N_36440);
xor U39423 (N_39423,N_37450,N_36140);
nand U39424 (N_39424,N_36553,N_36728);
or U39425 (N_39425,N_37362,N_36127);
and U39426 (N_39426,N_36837,N_37917);
nand U39427 (N_39427,N_37532,N_36373);
or U39428 (N_39428,N_37306,N_36798);
xor U39429 (N_39429,N_36157,N_36220);
xor U39430 (N_39430,N_37994,N_37703);
or U39431 (N_39431,N_37440,N_37676);
and U39432 (N_39432,N_37924,N_36287);
and U39433 (N_39433,N_37866,N_37541);
xnor U39434 (N_39434,N_37719,N_37238);
nor U39435 (N_39435,N_36678,N_36656);
nor U39436 (N_39436,N_37191,N_36227);
and U39437 (N_39437,N_36609,N_37238);
xnor U39438 (N_39438,N_37416,N_37997);
nor U39439 (N_39439,N_37833,N_37086);
or U39440 (N_39440,N_37383,N_36241);
or U39441 (N_39441,N_36047,N_36207);
or U39442 (N_39442,N_36532,N_36323);
nor U39443 (N_39443,N_37850,N_37792);
or U39444 (N_39444,N_37894,N_36435);
or U39445 (N_39445,N_37423,N_37145);
or U39446 (N_39446,N_37661,N_37579);
nand U39447 (N_39447,N_37549,N_36717);
nor U39448 (N_39448,N_37650,N_36916);
and U39449 (N_39449,N_37437,N_37564);
nand U39450 (N_39450,N_36174,N_36515);
or U39451 (N_39451,N_36331,N_36995);
and U39452 (N_39452,N_37866,N_37534);
and U39453 (N_39453,N_36207,N_37246);
and U39454 (N_39454,N_36540,N_37312);
and U39455 (N_39455,N_37133,N_37927);
nor U39456 (N_39456,N_37512,N_36904);
xnor U39457 (N_39457,N_36316,N_36985);
and U39458 (N_39458,N_37684,N_36277);
xnor U39459 (N_39459,N_37987,N_37188);
xor U39460 (N_39460,N_37216,N_36006);
and U39461 (N_39461,N_37022,N_36344);
nand U39462 (N_39462,N_37970,N_36015);
or U39463 (N_39463,N_36884,N_37193);
or U39464 (N_39464,N_37879,N_37417);
or U39465 (N_39465,N_37004,N_37372);
and U39466 (N_39466,N_36273,N_37067);
nand U39467 (N_39467,N_36663,N_36892);
nor U39468 (N_39468,N_37416,N_36292);
nor U39469 (N_39469,N_36681,N_36350);
nor U39470 (N_39470,N_36129,N_37023);
or U39471 (N_39471,N_37065,N_36185);
nand U39472 (N_39472,N_36480,N_36777);
or U39473 (N_39473,N_37068,N_36543);
or U39474 (N_39474,N_37352,N_37279);
or U39475 (N_39475,N_36330,N_36966);
or U39476 (N_39476,N_37842,N_36600);
xnor U39477 (N_39477,N_36286,N_37047);
nand U39478 (N_39478,N_36740,N_36310);
nor U39479 (N_39479,N_37758,N_37221);
and U39480 (N_39480,N_37470,N_36952);
xor U39481 (N_39481,N_36207,N_36559);
nand U39482 (N_39482,N_36948,N_36559);
nand U39483 (N_39483,N_37787,N_36069);
xnor U39484 (N_39484,N_37538,N_36199);
and U39485 (N_39485,N_36458,N_36119);
and U39486 (N_39486,N_37290,N_36241);
nor U39487 (N_39487,N_37009,N_37555);
and U39488 (N_39488,N_36205,N_36698);
and U39489 (N_39489,N_36507,N_36016);
xor U39490 (N_39490,N_37625,N_36263);
xnor U39491 (N_39491,N_37840,N_36689);
and U39492 (N_39492,N_37977,N_37799);
and U39493 (N_39493,N_36672,N_37478);
nor U39494 (N_39494,N_36454,N_36221);
or U39495 (N_39495,N_37858,N_37547);
nor U39496 (N_39496,N_37789,N_36761);
nor U39497 (N_39497,N_36958,N_37393);
nand U39498 (N_39498,N_36936,N_37315);
xor U39499 (N_39499,N_37103,N_37713);
xor U39500 (N_39500,N_36221,N_37740);
and U39501 (N_39501,N_37970,N_36387);
nor U39502 (N_39502,N_36335,N_37035);
and U39503 (N_39503,N_37392,N_37080);
xor U39504 (N_39504,N_37672,N_37804);
nand U39505 (N_39505,N_37495,N_36752);
nor U39506 (N_39506,N_37791,N_37150);
nor U39507 (N_39507,N_36188,N_37311);
nor U39508 (N_39508,N_36456,N_36390);
or U39509 (N_39509,N_36758,N_36880);
nand U39510 (N_39510,N_37532,N_36866);
nor U39511 (N_39511,N_37159,N_36886);
nor U39512 (N_39512,N_37576,N_36485);
nor U39513 (N_39513,N_36429,N_37316);
nor U39514 (N_39514,N_36551,N_37399);
and U39515 (N_39515,N_36055,N_37902);
nor U39516 (N_39516,N_36012,N_36370);
nand U39517 (N_39517,N_37188,N_37802);
nand U39518 (N_39518,N_36547,N_37868);
or U39519 (N_39519,N_37466,N_37188);
or U39520 (N_39520,N_37690,N_36994);
and U39521 (N_39521,N_37603,N_37933);
nand U39522 (N_39522,N_37033,N_36752);
nor U39523 (N_39523,N_36601,N_37586);
nand U39524 (N_39524,N_37325,N_37671);
or U39525 (N_39525,N_37800,N_36958);
or U39526 (N_39526,N_37321,N_36842);
nand U39527 (N_39527,N_37652,N_36186);
xnor U39528 (N_39528,N_36010,N_37751);
and U39529 (N_39529,N_37205,N_36987);
xor U39530 (N_39530,N_36004,N_36184);
nor U39531 (N_39531,N_37580,N_37182);
or U39532 (N_39532,N_37827,N_37029);
nor U39533 (N_39533,N_36702,N_36297);
nor U39534 (N_39534,N_36091,N_36070);
or U39535 (N_39535,N_37430,N_37638);
xor U39536 (N_39536,N_36038,N_37414);
or U39537 (N_39537,N_37652,N_36867);
xor U39538 (N_39538,N_37995,N_36877);
or U39539 (N_39539,N_37194,N_36767);
xnor U39540 (N_39540,N_36102,N_36447);
or U39541 (N_39541,N_37350,N_36486);
xor U39542 (N_39542,N_36181,N_36392);
or U39543 (N_39543,N_36319,N_36475);
xnor U39544 (N_39544,N_37235,N_37823);
or U39545 (N_39545,N_36229,N_37721);
xor U39546 (N_39546,N_37111,N_37559);
or U39547 (N_39547,N_36118,N_37978);
or U39548 (N_39548,N_36121,N_37451);
nor U39549 (N_39549,N_37848,N_36825);
xnor U39550 (N_39550,N_37767,N_37035);
nand U39551 (N_39551,N_36814,N_37314);
nand U39552 (N_39552,N_36956,N_37528);
and U39553 (N_39553,N_37433,N_37616);
nand U39554 (N_39554,N_37884,N_36000);
or U39555 (N_39555,N_36777,N_36941);
or U39556 (N_39556,N_36884,N_36804);
and U39557 (N_39557,N_37285,N_37503);
nor U39558 (N_39558,N_37962,N_36399);
nand U39559 (N_39559,N_36146,N_36830);
xnor U39560 (N_39560,N_37526,N_36772);
xnor U39561 (N_39561,N_37386,N_37844);
and U39562 (N_39562,N_36338,N_37006);
and U39563 (N_39563,N_37781,N_37735);
xor U39564 (N_39564,N_36633,N_37660);
nor U39565 (N_39565,N_36117,N_36736);
or U39566 (N_39566,N_37716,N_37757);
and U39567 (N_39567,N_37136,N_36334);
and U39568 (N_39568,N_36366,N_37639);
or U39569 (N_39569,N_37668,N_36331);
xnor U39570 (N_39570,N_36476,N_37439);
and U39571 (N_39571,N_37854,N_37600);
nand U39572 (N_39572,N_37671,N_37032);
or U39573 (N_39573,N_37641,N_37765);
nor U39574 (N_39574,N_36782,N_36380);
and U39575 (N_39575,N_36618,N_36636);
and U39576 (N_39576,N_36351,N_37949);
and U39577 (N_39577,N_36499,N_36136);
and U39578 (N_39578,N_36076,N_37646);
and U39579 (N_39579,N_37365,N_37133);
xnor U39580 (N_39580,N_36194,N_37847);
and U39581 (N_39581,N_37348,N_37977);
nand U39582 (N_39582,N_36672,N_36420);
nand U39583 (N_39583,N_36358,N_36109);
nor U39584 (N_39584,N_36765,N_37818);
xnor U39585 (N_39585,N_37633,N_37882);
xor U39586 (N_39586,N_36400,N_37174);
xnor U39587 (N_39587,N_36906,N_37246);
and U39588 (N_39588,N_37038,N_36983);
and U39589 (N_39589,N_37230,N_36187);
nor U39590 (N_39590,N_36028,N_37423);
nor U39591 (N_39591,N_36727,N_36827);
nor U39592 (N_39592,N_37668,N_36406);
or U39593 (N_39593,N_37806,N_37598);
xnor U39594 (N_39594,N_37560,N_37466);
nor U39595 (N_39595,N_36391,N_37783);
xor U39596 (N_39596,N_36129,N_37215);
nand U39597 (N_39597,N_36172,N_37839);
nand U39598 (N_39598,N_37541,N_37468);
or U39599 (N_39599,N_36567,N_36576);
nor U39600 (N_39600,N_36900,N_36020);
and U39601 (N_39601,N_36890,N_37379);
nor U39602 (N_39602,N_37371,N_36149);
xnor U39603 (N_39603,N_36621,N_36192);
and U39604 (N_39604,N_36145,N_37975);
nor U39605 (N_39605,N_36071,N_36960);
xnor U39606 (N_39606,N_36197,N_37686);
xor U39607 (N_39607,N_36503,N_36760);
nor U39608 (N_39608,N_37438,N_36929);
and U39609 (N_39609,N_36791,N_37175);
nand U39610 (N_39610,N_36122,N_37471);
nand U39611 (N_39611,N_37062,N_36363);
nand U39612 (N_39612,N_36988,N_36647);
nand U39613 (N_39613,N_36718,N_37282);
nand U39614 (N_39614,N_36476,N_36982);
nor U39615 (N_39615,N_37903,N_36792);
nand U39616 (N_39616,N_37164,N_36057);
and U39617 (N_39617,N_36183,N_37412);
nand U39618 (N_39618,N_37237,N_37525);
nor U39619 (N_39619,N_37751,N_37581);
nor U39620 (N_39620,N_37614,N_37564);
nor U39621 (N_39621,N_36732,N_36253);
and U39622 (N_39622,N_36642,N_37490);
and U39623 (N_39623,N_37959,N_37855);
and U39624 (N_39624,N_37214,N_36847);
xnor U39625 (N_39625,N_36164,N_37133);
nor U39626 (N_39626,N_36820,N_36734);
xor U39627 (N_39627,N_36785,N_37237);
and U39628 (N_39628,N_36187,N_36292);
and U39629 (N_39629,N_37651,N_37355);
or U39630 (N_39630,N_37021,N_37970);
xor U39631 (N_39631,N_36180,N_37702);
and U39632 (N_39632,N_36072,N_36600);
and U39633 (N_39633,N_37823,N_36058);
or U39634 (N_39634,N_36396,N_36238);
nand U39635 (N_39635,N_36963,N_37357);
xnor U39636 (N_39636,N_36092,N_37025);
and U39637 (N_39637,N_36793,N_37736);
xor U39638 (N_39638,N_36766,N_37959);
nor U39639 (N_39639,N_36488,N_37509);
or U39640 (N_39640,N_37819,N_36989);
and U39641 (N_39641,N_36606,N_37658);
nand U39642 (N_39642,N_37479,N_37629);
xor U39643 (N_39643,N_36940,N_37753);
or U39644 (N_39644,N_37625,N_37255);
and U39645 (N_39645,N_36133,N_36462);
xor U39646 (N_39646,N_37085,N_36373);
or U39647 (N_39647,N_36925,N_36224);
nand U39648 (N_39648,N_36698,N_37154);
xnor U39649 (N_39649,N_36829,N_37199);
nor U39650 (N_39650,N_37392,N_37558);
nor U39651 (N_39651,N_37175,N_37081);
or U39652 (N_39652,N_37695,N_37217);
or U39653 (N_39653,N_36604,N_36014);
and U39654 (N_39654,N_36041,N_36002);
or U39655 (N_39655,N_36933,N_37005);
nor U39656 (N_39656,N_37055,N_37358);
nor U39657 (N_39657,N_36789,N_36173);
nand U39658 (N_39658,N_37844,N_36758);
or U39659 (N_39659,N_36944,N_37716);
xor U39660 (N_39660,N_36730,N_37989);
and U39661 (N_39661,N_37945,N_37614);
or U39662 (N_39662,N_37327,N_36979);
nand U39663 (N_39663,N_36254,N_36735);
nor U39664 (N_39664,N_37026,N_37041);
nand U39665 (N_39665,N_36543,N_36414);
nor U39666 (N_39666,N_36034,N_36746);
and U39667 (N_39667,N_36842,N_36772);
nor U39668 (N_39668,N_36010,N_37330);
nand U39669 (N_39669,N_36891,N_36728);
nand U39670 (N_39670,N_37710,N_36794);
nand U39671 (N_39671,N_36316,N_37133);
nor U39672 (N_39672,N_37000,N_37495);
and U39673 (N_39673,N_37890,N_36570);
xnor U39674 (N_39674,N_36165,N_36725);
and U39675 (N_39675,N_37064,N_36341);
nand U39676 (N_39676,N_36719,N_37408);
nand U39677 (N_39677,N_36183,N_36120);
and U39678 (N_39678,N_37990,N_36914);
xor U39679 (N_39679,N_37017,N_37934);
nor U39680 (N_39680,N_36078,N_36949);
xor U39681 (N_39681,N_37784,N_36384);
and U39682 (N_39682,N_37214,N_36233);
nor U39683 (N_39683,N_36087,N_36656);
or U39684 (N_39684,N_36016,N_36059);
and U39685 (N_39685,N_37015,N_37086);
or U39686 (N_39686,N_37233,N_37741);
and U39687 (N_39687,N_37453,N_36745);
xnor U39688 (N_39688,N_37245,N_36146);
nand U39689 (N_39689,N_37632,N_36158);
and U39690 (N_39690,N_36733,N_36792);
nor U39691 (N_39691,N_36252,N_36159);
or U39692 (N_39692,N_36656,N_36651);
or U39693 (N_39693,N_36292,N_36516);
nand U39694 (N_39694,N_36715,N_37129);
nand U39695 (N_39695,N_36887,N_37296);
nor U39696 (N_39696,N_36368,N_37439);
nor U39697 (N_39697,N_37766,N_36092);
nand U39698 (N_39698,N_37140,N_37190);
xor U39699 (N_39699,N_36464,N_37225);
nor U39700 (N_39700,N_37084,N_36009);
nor U39701 (N_39701,N_36162,N_37880);
nand U39702 (N_39702,N_36075,N_37953);
xnor U39703 (N_39703,N_36158,N_37790);
and U39704 (N_39704,N_36561,N_36925);
nand U39705 (N_39705,N_37226,N_36642);
and U39706 (N_39706,N_36669,N_37399);
or U39707 (N_39707,N_37680,N_36926);
xor U39708 (N_39708,N_37783,N_36958);
xor U39709 (N_39709,N_36320,N_37894);
and U39710 (N_39710,N_37749,N_37021);
xnor U39711 (N_39711,N_37223,N_36746);
nor U39712 (N_39712,N_36371,N_36226);
or U39713 (N_39713,N_36045,N_37614);
or U39714 (N_39714,N_36770,N_37162);
xnor U39715 (N_39715,N_37473,N_36716);
nor U39716 (N_39716,N_36742,N_37283);
nand U39717 (N_39717,N_37379,N_37340);
nor U39718 (N_39718,N_37397,N_36004);
nand U39719 (N_39719,N_36287,N_37603);
nor U39720 (N_39720,N_36159,N_36237);
nor U39721 (N_39721,N_37731,N_37671);
or U39722 (N_39722,N_36032,N_36381);
nor U39723 (N_39723,N_36035,N_37378);
xor U39724 (N_39724,N_36502,N_36936);
nand U39725 (N_39725,N_36709,N_37286);
nand U39726 (N_39726,N_36495,N_37159);
nand U39727 (N_39727,N_36240,N_37288);
nand U39728 (N_39728,N_37895,N_36159);
nand U39729 (N_39729,N_36893,N_36857);
nand U39730 (N_39730,N_37940,N_37079);
nand U39731 (N_39731,N_37773,N_37580);
or U39732 (N_39732,N_37218,N_37830);
and U39733 (N_39733,N_36884,N_37058);
nand U39734 (N_39734,N_37508,N_37934);
or U39735 (N_39735,N_36515,N_37371);
nand U39736 (N_39736,N_37877,N_36215);
nand U39737 (N_39737,N_36228,N_37695);
or U39738 (N_39738,N_36996,N_37578);
nor U39739 (N_39739,N_37221,N_36752);
nand U39740 (N_39740,N_36434,N_36637);
nand U39741 (N_39741,N_36445,N_37378);
nor U39742 (N_39742,N_37551,N_36123);
nor U39743 (N_39743,N_36406,N_37576);
or U39744 (N_39744,N_36737,N_36247);
and U39745 (N_39745,N_37045,N_37813);
xnor U39746 (N_39746,N_36825,N_37918);
nor U39747 (N_39747,N_37801,N_37732);
xor U39748 (N_39748,N_36979,N_37299);
or U39749 (N_39749,N_36099,N_37084);
xor U39750 (N_39750,N_37163,N_37299);
nand U39751 (N_39751,N_36009,N_36056);
nor U39752 (N_39752,N_36078,N_37062);
and U39753 (N_39753,N_37008,N_37931);
nor U39754 (N_39754,N_36818,N_36777);
nor U39755 (N_39755,N_36571,N_37691);
nor U39756 (N_39756,N_36128,N_37726);
or U39757 (N_39757,N_36613,N_37464);
xor U39758 (N_39758,N_37399,N_36862);
nand U39759 (N_39759,N_37613,N_36697);
nand U39760 (N_39760,N_36189,N_36207);
or U39761 (N_39761,N_37207,N_37451);
nor U39762 (N_39762,N_36350,N_37942);
xnor U39763 (N_39763,N_37725,N_37933);
or U39764 (N_39764,N_36640,N_37386);
and U39765 (N_39765,N_37147,N_37573);
or U39766 (N_39766,N_37975,N_37565);
xnor U39767 (N_39767,N_37555,N_36071);
xnor U39768 (N_39768,N_37648,N_36086);
nand U39769 (N_39769,N_36045,N_36538);
or U39770 (N_39770,N_37047,N_36626);
nor U39771 (N_39771,N_36038,N_36755);
or U39772 (N_39772,N_36683,N_36204);
and U39773 (N_39773,N_36455,N_36089);
or U39774 (N_39774,N_37846,N_37931);
nand U39775 (N_39775,N_36202,N_36473);
xnor U39776 (N_39776,N_37616,N_36614);
nand U39777 (N_39777,N_37147,N_36889);
or U39778 (N_39778,N_37648,N_36791);
xor U39779 (N_39779,N_37213,N_36906);
xnor U39780 (N_39780,N_37428,N_36929);
nand U39781 (N_39781,N_36300,N_36401);
and U39782 (N_39782,N_36574,N_36382);
xnor U39783 (N_39783,N_36013,N_36624);
nor U39784 (N_39784,N_37101,N_37023);
nand U39785 (N_39785,N_36512,N_37730);
and U39786 (N_39786,N_36916,N_37380);
or U39787 (N_39787,N_36352,N_37573);
nor U39788 (N_39788,N_36374,N_36668);
or U39789 (N_39789,N_36459,N_37035);
xnor U39790 (N_39790,N_36260,N_37546);
and U39791 (N_39791,N_36046,N_36048);
and U39792 (N_39792,N_36644,N_37658);
xnor U39793 (N_39793,N_37901,N_37557);
and U39794 (N_39794,N_36934,N_36302);
or U39795 (N_39795,N_37453,N_36494);
nor U39796 (N_39796,N_36056,N_36260);
or U39797 (N_39797,N_37829,N_37698);
xnor U39798 (N_39798,N_36242,N_37236);
nand U39799 (N_39799,N_37591,N_37420);
and U39800 (N_39800,N_37968,N_36733);
or U39801 (N_39801,N_36152,N_37416);
nand U39802 (N_39802,N_37061,N_37067);
nor U39803 (N_39803,N_37265,N_37940);
nor U39804 (N_39804,N_36033,N_36172);
xnor U39805 (N_39805,N_37559,N_36040);
or U39806 (N_39806,N_36235,N_37544);
xnor U39807 (N_39807,N_37912,N_37439);
or U39808 (N_39808,N_36711,N_36004);
nand U39809 (N_39809,N_37946,N_37524);
nand U39810 (N_39810,N_37719,N_36119);
and U39811 (N_39811,N_36351,N_37822);
nor U39812 (N_39812,N_36344,N_36908);
nor U39813 (N_39813,N_37419,N_36433);
and U39814 (N_39814,N_36810,N_36060);
nor U39815 (N_39815,N_37506,N_37977);
or U39816 (N_39816,N_37826,N_36837);
and U39817 (N_39817,N_36935,N_36920);
nor U39818 (N_39818,N_36831,N_36346);
and U39819 (N_39819,N_37738,N_37776);
nor U39820 (N_39820,N_36182,N_37158);
nand U39821 (N_39821,N_36653,N_37670);
nand U39822 (N_39822,N_36441,N_36492);
and U39823 (N_39823,N_36787,N_37777);
or U39824 (N_39824,N_36843,N_36570);
nor U39825 (N_39825,N_36031,N_36190);
xnor U39826 (N_39826,N_36215,N_36496);
and U39827 (N_39827,N_37526,N_37024);
nand U39828 (N_39828,N_36527,N_37077);
nand U39829 (N_39829,N_37693,N_36167);
nand U39830 (N_39830,N_36404,N_36336);
nor U39831 (N_39831,N_37059,N_36250);
and U39832 (N_39832,N_36530,N_36450);
or U39833 (N_39833,N_36286,N_37999);
nand U39834 (N_39834,N_36073,N_37125);
nand U39835 (N_39835,N_37085,N_36617);
nand U39836 (N_39836,N_37156,N_37879);
or U39837 (N_39837,N_37669,N_36770);
xor U39838 (N_39838,N_37129,N_37951);
or U39839 (N_39839,N_36137,N_36455);
nor U39840 (N_39840,N_36745,N_36192);
xor U39841 (N_39841,N_37077,N_37973);
or U39842 (N_39842,N_37851,N_37829);
xor U39843 (N_39843,N_37833,N_37834);
and U39844 (N_39844,N_36328,N_36639);
nand U39845 (N_39845,N_36998,N_37203);
nor U39846 (N_39846,N_37493,N_37879);
or U39847 (N_39847,N_36263,N_36056);
or U39848 (N_39848,N_37136,N_37017);
xnor U39849 (N_39849,N_37660,N_36841);
xor U39850 (N_39850,N_37819,N_37042);
xnor U39851 (N_39851,N_37899,N_37767);
nand U39852 (N_39852,N_37805,N_37071);
or U39853 (N_39853,N_36572,N_37644);
and U39854 (N_39854,N_37600,N_37872);
nand U39855 (N_39855,N_37147,N_37719);
nand U39856 (N_39856,N_37784,N_36851);
nor U39857 (N_39857,N_37471,N_36704);
or U39858 (N_39858,N_37831,N_36964);
xor U39859 (N_39859,N_37824,N_36119);
nor U39860 (N_39860,N_37415,N_37982);
and U39861 (N_39861,N_37022,N_37150);
xnor U39862 (N_39862,N_36279,N_36319);
nand U39863 (N_39863,N_36359,N_37669);
nand U39864 (N_39864,N_37772,N_37134);
nand U39865 (N_39865,N_37587,N_37823);
and U39866 (N_39866,N_37210,N_36762);
nand U39867 (N_39867,N_36499,N_37247);
or U39868 (N_39868,N_37202,N_36161);
nand U39869 (N_39869,N_37189,N_36903);
nand U39870 (N_39870,N_36636,N_36841);
nor U39871 (N_39871,N_36612,N_37024);
or U39872 (N_39872,N_36919,N_37314);
nor U39873 (N_39873,N_36369,N_36788);
and U39874 (N_39874,N_37301,N_36217);
xnor U39875 (N_39875,N_36824,N_37696);
or U39876 (N_39876,N_37439,N_37148);
or U39877 (N_39877,N_36293,N_36718);
nand U39878 (N_39878,N_36184,N_37529);
nand U39879 (N_39879,N_36156,N_36206);
nor U39880 (N_39880,N_37043,N_37138);
or U39881 (N_39881,N_37398,N_36235);
nand U39882 (N_39882,N_37426,N_36518);
xnor U39883 (N_39883,N_36293,N_36507);
xor U39884 (N_39884,N_37501,N_37259);
nand U39885 (N_39885,N_37921,N_37663);
and U39886 (N_39886,N_37163,N_36490);
and U39887 (N_39887,N_36805,N_36303);
or U39888 (N_39888,N_36766,N_37566);
nor U39889 (N_39889,N_37464,N_37520);
xor U39890 (N_39890,N_37616,N_37989);
or U39891 (N_39891,N_37788,N_36503);
and U39892 (N_39892,N_36954,N_37404);
and U39893 (N_39893,N_37917,N_36927);
and U39894 (N_39894,N_37865,N_36423);
xor U39895 (N_39895,N_37143,N_37653);
or U39896 (N_39896,N_36837,N_37807);
and U39897 (N_39897,N_36800,N_36516);
and U39898 (N_39898,N_37144,N_37302);
or U39899 (N_39899,N_37416,N_37532);
nand U39900 (N_39900,N_36217,N_36540);
nand U39901 (N_39901,N_37801,N_37193);
nor U39902 (N_39902,N_37934,N_37041);
nand U39903 (N_39903,N_37975,N_37545);
or U39904 (N_39904,N_37822,N_37268);
xnor U39905 (N_39905,N_37685,N_37478);
or U39906 (N_39906,N_37548,N_37539);
and U39907 (N_39907,N_36897,N_37023);
nand U39908 (N_39908,N_36776,N_37347);
and U39909 (N_39909,N_37224,N_37401);
nand U39910 (N_39910,N_36114,N_36407);
nand U39911 (N_39911,N_36410,N_37138);
nor U39912 (N_39912,N_36439,N_37830);
and U39913 (N_39913,N_37311,N_37449);
and U39914 (N_39914,N_36114,N_37119);
or U39915 (N_39915,N_37440,N_36721);
or U39916 (N_39916,N_36566,N_36155);
xor U39917 (N_39917,N_36508,N_37601);
or U39918 (N_39918,N_36835,N_37274);
and U39919 (N_39919,N_37813,N_37352);
nor U39920 (N_39920,N_36076,N_36823);
and U39921 (N_39921,N_37274,N_37977);
xor U39922 (N_39922,N_36070,N_37365);
and U39923 (N_39923,N_36684,N_37850);
nor U39924 (N_39924,N_37650,N_37389);
nand U39925 (N_39925,N_36153,N_36830);
or U39926 (N_39926,N_37304,N_36543);
nor U39927 (N_39927,N_36682,N_37382);
xor U39928 (N_39928,N_37342,N_37038);
nor U39929 (N_39929,N_36998,N_36815);
xor U39930 (N_39930,N_36216,N_37996);
nor U39931 (N_39931,N_37811,N_36042);
xnor U39932 (N_39932,N_36636,N_37833);
and U39933 (N_39933,N_36017,N_37513);
and U39934 (N_39934,N_37974,N_36876);
or U39935 (N_39935,N_37699,N_37748);
xnor U39936 (N_39936,N_36591,N_36986);
xnor U39937 (N_39937,N_37903,N_37614);
xor U39938 (N_39938,N_37570,N_37509);
xor U39939 (N_39939,N_37473,N_36116);
xor U39940 (N_39940,N_37644,N_36446);
xor U39941 (N_39941,N_37916,N_36618);
and U39942 (N_39942,N_36784,N_37942);
nor U39943 (N_39943,N_36545,N_36674);
xor U39944 (N_39944,N_36018,N_37781);
nor U39945 (N_39945,N_37579,N_36149);
or U39946 (N_39946,N_36771,N_36497);
and U39947 (N_39947,N_36885,N_36696);
or U39948 (N_39948,N_37767,N_37282);
xnor U39949 (N_39949,N_36508,N_37654);
nor U39950 (N_39950,N_37789,N_37959);
nor U39951 (N_39951,N_36713,N_36629);
xnor U39952 (N_39952,N_36082,N_37282);
and U39953 (N_39953,N_36851,N_36003);
xor U39954 (N_39954,N_36635,N_37676);
xnor U39955 (N_39955,N_37735,N_36859);
or U39956 (N_39956,N_37522,N_37110);
nor U39957 (N_39957,N_37490,N_37941);
or U39958 (N_39958,N_36329,N_36358);
nand U39959 (N_39959,N_37133,N_37777);
nand U39960 (N_39960,N_36992,N_36092);
nand U39961 (N_39961,N_37808,N_37257);
and U39962 (N_39962,N_37421,N_37300);
nand U39963 (N_39963,N_37417,N_36942);
or U39964 (N_39964,N_36429,N_37347);
nand U39965 (N_39965,N_36147,N_37217);
or U39966 (N_39966,N_36798,N_36763);
xnor U39967 (N_39967,N_37811,N_37212);
or U39968 (N_39968,N_36312,N_36897);
xnor U39969 (N_39969,N_36104,N_36439);
and U39970 (N_39970,N_36059,N_37990);
and U39971 (N_39971,N_36930,N_36133);
nand U39972 (N_39972,N_37193,N_36277);
or U39973 (N_39973,N_37796,N_37246);
or U39974 (N_39974,N_37505,N_36613);
nor U39975 (N_39975,N_36758,N_37255);
xor U39976 (N_39976,N_36978,N_36035);
nor U39977 (N_39977,N_36952,N_37220);
nand U39978 (N_39978,N_37973,N_37203);
and U39979 (N_39979,N_37834,N_37921);
nor U39980 (N_39980,N_37405,N_37278);
nor U39981 (N_39981,N_37270,N_37508);
xor U39982 (N_39982,N_36039,N_36413);
nor U39983 (N_39983,N_37446,N_36779);
nor U39984 (N_39984,N_37123,N_37443);
and U39985 (N_39985,N_37140,N_36867);
xnor U39986 (N_39986,N_36458,N_36289);
xnor U39987 (N_39987,N_36072,N_36867);
nand U39988 (N_39988,N_37082,N_37023);
nand U39989 (N_39989,N_37473,N_37897);
or U39990 (N_39990,N_37973,N_37490);
nor U39991 (N_39991,N_36982,N_37242);
or U39992 (N_39992,N_37667,N_37333);
nand U39993 (N_39993,N_36624,N_36280);
or U39994 (N_39994,N_37139,N_37351);
nor U39995 (N_39995,N_36782,N_36303);
xnor U39996 (N_39996,N_36109,N_36053);
xor U39997 (N_39997,N_36608,N_37066);
nand U39998 (N_39998,N_37381,N_36399);
or U39999 (N_39999,N_36314,N_37031);
and U40000 (N_40000,N_39806,N_39490);
nor U40001 (N_40001,N_39299,N_38142);
or U40002 (N_40002,N_39439,N_39457);
nor U40003 (N_40003,N_38800,N_39406);
nor U40004 (N_40004,N_39470,N_38160);
nor U40005 (N_40005,N_38239,N_38143);
nand U40006 (N_40006,N_38762,N_38335);
xor U40007 (N_40007,N_39221,N_38657);
nand U40008 (N_40008,N_38483,N_38985);
xor U40009 (N_40009,N_38784,N_39564);
nand U40010 (N_40010,N_39360,N_38659);
nand U40011 (N_40011,N_39953,N_38253);
nor U40012 (N_40012,N_38796,N_39990);
or U40013 (N_40013,N_39204,N_39570);
xor U40014 (N_40014,N_38058,N_38471);
xor U40015 (N_40015,N_38599,N_38674);
nand U40016 (N_40016,N_38653,N_38922);
nand U40017 (N_40017,N_38581,N_39844);
or U40018 (N_40018,N_38202,N_38215);
nor U40019 (N_40019,N_39502,N_38013);
nor U40020 (N_40020,N_39504,N_39617);
or U40021 (N_40021,N_39975,N_39563);
or U40022 (N_40022,N_39209,N_39545);
nand U40023 (N_40023,N_39555,N_39270);
xnor U40024 (N_40024,N_38692,N_38145);
nand U40025 (N_40025,N_39069,N_39973);
or U40026 (N_40026,N_39155,N_38363);
nand U40027 (N_40027,N_39551,N_39843);
or U40028 (N_40028,N_39829,N_39860);
and U40029 (N_40029,N_39359,N_38908);
xnor U40030 (N_40030,N_38693,N_39768);
and U40031 (N_40031,N_39669,N_39903);
nor U40032 (N_40032,N_38466,N_38056);
or U40033 (N_40033,N_39626,N_39809);
xnor U40034 (N_40034,N_38604,N_38696);
and U40035 (N_40035,N_39871,N_38989);
xnor U40036 (N_40036,N_38356,N_39110);
or U40037 (N_40037,N_38726,N_38181);
nand U40038 (N_40038,N_39425,N_38544);
nand U40039 (N_40039,N_38209,N_39097);
and U40040 (N_40040,N_39275,N_38462);
or U40041 (N_40041,N_39734,N_38447);
and U40042 (N_40042,N_39991,N_39639);
or U40043 (N_40043,N_39552,N_38357);
or U40044 (N_40044,N_39194,N_39647);
nand U40045 (N_40045,N_38470,N_38963);
xor U40046 (N_40046,N_38074,N_38857);
xnor U40047 (N_40047,N_38804,N_39652);
nor U40048 (N_40048,N_39598,N_38860);
xor U40049 (N_40049,N_39489,N_38981);
nor U40050 (N_40050,N_39696,N_39873);
nor U40051 (N_40051,N_39213,N_38545);
or U40052 (N_40052,N_39288,N_39586);
nor U40053 (N_40053,N_38083,N_39324);
nand U40054 (N_40054,N_38438,N_38130);
or U40055 (N_40055,N_38161,N_39841);
nor U40056 (N_40056,N_38348,N_38894);
nand U40057 (N_40057,N_38073,N_39503);
or U40058 (N_40058,N_39158,N_38861);
and U40059 (N_40059,N_38248,N_39648);
nand U40060 (N_40060,N_39154,N_38064);
or U40061 (N_40061,N_38311,N_39087);
and U40062 (N_40062,N_39801,N_38071);
nor U40063 (N_40063,N_38264,N_39114);
xnor U40064 (N_40064,N_38088,N_38267);
xor U40065 (N_40065,N_39714,N_38178);
nand U40066 (N_40066,N_38733,N_38694);
xnor U40067 (N_40067,N_39113,N_38139);
xnor U40068 (N_40068,N_39842,N_38243);
nand U40069 (N_40069,N_38467,N_38876);
nor U40070 (N_40070,N_39635,N_38306);
nor U40071 (N_40071,N_38537,N_39199);
and U40072 (N_40072,N_38761,N_39085);
or U40073 (N_40073,N_39468,N_39845);
nor U40074 (N_40074,N_38159,N_39337);
xor U40075 (N_40075,N_38944,N_38059);
or U40076 (N_40076,N_39314,N_38309);
nor U40077 (N_40077,N_38385,N_39574);
xor U40078 (N_40078,N_38360,N_38988);
xor U40079 (N_40079,N_39320,N_38703);
or U40080 (N_40080,N_39680,N_39001);
xnor U40081 (N_40081,N_39893,N_39536);
xnor U40082 (N_40082,N_39569,N_39079);
nand U40083 (N_40083,N_39746,N_39910);
nand U40084 (N_40084,N_38872,N_38710);
xor U40085 (N_40085,N_38927,N_39804);
nor U40086 (N_40086,N_38384,N_38967);
nand U40087 (N_40087,N_39813,N_39447);
xnor U40088 (N_40088,N_38389,N_39814);
nor U40089 (N_40089,N_39957,N_39775);
nor U40090 (N_40090,N_39041,N_38259);
xnor U40091 (N_40091,N_38719,N_38245);
or U40092 (N_40092,N_39721,N_39119);
or U40093 (N_40093,N_38204,N_38421);
nand U40094 (N_40094,N_39779,N_39044);
and U40095 (N_40095,N_39345,N_38051);
and U40096 (N_40096,N_39753,N_39277);
or U40097 (N_40097,N_38287,N_38042);
or U40098 (N_40098,N_38153,N_38140);
or U40099 (N_40099,N_38839,N_38551);
nor U40100 (N_40100,N_39784,N_39152);
and U40101 (N_40101,N_38247,N_39442);
nand U40102 (N_40102,N_38075,N_39864);
or U40103 (N_40103,N_38716,N_39733);
xnor U40104 (N_40104,N_39189,N_39538);
or U40105 (N_40105,N_39177,N_38543);
and U40106 (N_40106,N_39679,N_39583);
or U40107 (N_40107,N_39467,N_39747);
nor U40108 (N_40108,N_38125,N_38878);
nor U40109 (N_40109,N_39237,N_38100);
or U40110 (N_40110,N_39043,N_39322);
or U40111 (N_40111,N_39748,N_38144);
xor U40112 (N_40112,N_38034,N_38899);
xor U40113 (N_40113,N_39151,N_38958);
nand U40114 (N_40114,N_39413,N_39946);
nand U40115 (N_40115,N_38523,N_38501);
nand U40116 (N_40116,N_38330,N_39026);
nor U40117 (N_40117,N_38082,N_39281);
and U40118 (N_40118,N_38399,N_38270);
nand U40119 (N_40119,N_38835,N_39274);
and U40120 (N_40120,N_38709,N_39913);
nor U40121 (N_40121,N_39115,N_39854);
nand U40122 (N_40122,N_38195,N_38177);
nand U40123 (N_40123,N_38162,N_38532);
nor U40124 (N_40124,N_38921,N_39445);
or U40125 (N_40125,N_38187,N_39614);
nor U40126 (N_40126,N_38624,N_39762);
or U40127 (N_40127,N_38858,N_38031);
nand U40128 (N_40128,N_38240,N_39018);
nand U40129 (N_40129,N_39620,N_38738);
xnor U40130 (N_40130,N_39928,N_39098);
nor U40131 (N_40131,N_38821,N_38920);
xnor U40132 (N_40132,N_38369,N_38035);
nor U40133 (N_40133,N_39348,N_39571);
or U40134 (N_40134,N_39109,N_38156);
or U40135 (N_40135,N_38969,N_39601);
or U40136 (N_40136,N_39223,N_38990);
or U40137 (N_40137,N_39798,N_39567);
nand U40138 (N_40138,N_38234,N_39219);
nor U40139 (N_40139,N_38103,N_38011);
xor U40140 (N_40140,N_38806,N_39046);
nand U40141 (N_40141,N_38705,N_39476);
or U40142 (N_40142,N_38318,N_39452);
and U40143 (N_40143,N_38069,N_39145);
nor U40144 (N_40144,N_38896,N_38208);
nand U40145 (N_40145,N_39157,N_38026);
nand U40146 (N_40146,N_38179,N_38236);
nand U40147 (N_40147,N_39770,N_38475);
nand U40148 (N_40148,N_38729,N_38603);
nand U40149 (N_40149,N_38233,N_38200);
nand U40150 (N_40150,N_39883,N_38732);
xor U40151 (N_40151,N_38898,N_39279);
nor U40152 (N_40152,N_39278,N_39783);
nand U40153 (N_40153,N_39141,N_38948);
nand U40154 (N_40154,N_39610,N_39391);
and U40155 (N_40155,N_38822,N_39589);
xnor U40156 (N_40156,N_38353,N_39282);
nand U40157 (N_40157,N_39054,N_38002);
xnor U40158 (N_40158,N_39584,N_38323);
xnor U40159 (N_40159,N_39901,N_38676);
nand U40160 (N_40160,N_38910,N_39495);
and U40161 (N_40161,N_39068,N_38246);
or U40162 (N_40162,N_39911,N_39165);
and U40163 (N_40163,N_38201,N_38009);
and U40164 (N_40164,N_38128,N_38783);
and U40165 (N_40165,N_38020,N_39848);
or U40166 (N_40166,N_39700,N_38104);
nor U40167 (N_40167,N_38146,N_38403);
nor U40168 (N_40168,N_39838,N_38527);
or U40169 (N_40169,N_39764,N_39805);
and U40170 (N_40170,N_38352,N_38167);
nand U40171 (N_40171,N_38884,N_38266);
nor U40172 (N_40172,N_39186,N_39437);
nand U40173 (N_40173,N_39292,N_38480);
or U40174 (N_40174,N_39658,N_38423);
xnor U40175 (N_40175,N_39821,N_39232);
nand U40176 (N_40176,N_39318,N_38408);
nor U40177 (N_40177,N_38788,N_38049);
and U40178 (N_40178,N_38137,N_38307);
or U40179 (N_40179,N_38117,N_39884);
nor U40180 (N_40180,N_38736,N_39301);
nor U40181 (N_40181,N_38956,N_39710);
nor U40182 (N_40182,N_39865,N_38756);
xor U40183 (N_40183,N_38645,N_38824);
nand U40184 (N_40184,N_38123,N_38238);
xor U40185 (N_40185,N_38608,N_39531);
or U40186 (N_40186,N_39673,N_39047);
xnor U40187 (N_40187,N_38606,N_39429);
and U40188 (N_40188,N_39855,N_38838);
nor U40189 (N_40189,N_39577,N_38873);
nor U40190 (N_40190,N_39866,N_38598);
nor U40191 (N_40191,N_39167,N_39212);
nor U40192 (N_40192,N_39859,N_39815);
nor U40193 (N_40193,N_39267,N_38818);
nor U40194 (N_40194,N_38627,N_39817);
nor U40195 (N_40195,N_39233,N_38803);
nand U40196 (N_40196,N_38514,N_39183);
or U40197 (N_40197,N_38378,N_39641);
nor U40198 (N_40198,N_39729,N_38715);
nand U40199 (N_40199,N_39365,N_39256);
nor U40200 (N_40200,N_38664,N_39440);
nor U40201 (N_40201,N_39972,N_39987);
or U40202 (N_40202,N_39311,N_39168);
nor U40203 (N_40203,N_39794,N_39058);
or U40204 (N_40204,N_38095,N_39364);
nand U40205 (N_40205,N_39180,N_39600);
or U40206 (N_40206,N_38684,N_38512);
and U40207 (N_40207,N_39251,N_38834);
and U40208 (N_40208,N_39590,N_39244);
nor U40209 (N_40209,N_39675,N_38890);
or U40210 (N_40210,N_38326,N_39431);
and U40211 (N_40211,N_38015,N_38063);
xor U40212 (N_40212,N_38583,N_38749);
nand U40213 (N_40213,N_38122,N_39833);
nor U40214 (N_40214,N_39788,N_39171);
nor U40215 (N_40215,N_38984,N_39191);
nor U40216 (N_40216,N_39510,N_39162);
and U40217 (N_40217,N_38638,N_39464);
or U40218 (N_40218,N_38443,N_38040);
xnor U40219 (N_40219,N_39613,N_38735);
xor U40220 (N_40220,N_38019,N_38205);
nand U40221 (N_40221,N_38991,N_39943);
nor U40222 (N_40222,N_38650,N_38740);
or U40223 (N_40223,N_38765,N_39965);
xnor U40224 (N_40224,N_39433,N_39507);
nor U40225 (N_40225,N_38157,N_39917);
nor U40226 (N_40226,N_39882,N_39184);
nor U40227 (N_40227,N_38265,N_39377);
xnor U40228 (N_40228,N_39238,N_38983);
xor U40229 (N_40229,N_38014,N_38312);
and U40230 (N_40230,N_38376,N_38327);
nor U40231 (N_40231,N_38704,N_38502);
nand U40232 (N_40232,N_38281,N_39636);
nand U40233 (N_40233,N_39397,N_39560);
nand U40234 (N_40234,N_39646,N_38531);
nor U40235 (N_40235,N_38972,N_38560);
nor U40236 (N_40236,N_39343,N_39637);
or U40237 (N_40237,N_38743,N_38428);
nand U40238 (N_40238,N_38007,N_39607);
xor U40239 (N_40239,N_39053,N_39438);
nand U40240 (N_40240,N_39019,N_38024);
and U40241 (N_40241,N_39422,N_38955);
xor U40242 (N_40242,N_38728,N_39615);
xnor U40243 (N_40243,N_38488,N_38744);
xnor U40244 (N_40244,N_39492,N_39816);
and U40245 (N_40245,N_38493,N_38552);
or U40246 (N_40246,N_39938,N_39619);
xor U40247 (N_40247,N_39543,N_38637);
nor U40248 (N_40248,N_39969,N_39056);
nand U40249 (N_40249,N_39872,N_39588);
xnor U40250 (N_40250,N_39924,N_39090);
nor U40251 (N_40251,N_38135,N_39683);
nand U40252 (N_40252,N_38329,N_39720);
xor U40253 (N_40253,N_38010,N_38597);
or U40254 (N_40254,N_39082,N_38962);
nand U40255 (N_40255,N_39653,N_39395);
nand U40256 (N_40256,N_39549,N_38118);
nor U40257 (N_40257,N_39136,N_38998);
xor U40258 (N_40258,N_39978,N_38620);
or U40259 (N_40259,N_39891,N_38395);
and U40260 (N_40260,N_38717,N_39491);
xnor U40261 (N_40261,N_38321,N_39206);
and U40262 (N_40262,N_39914,N_38305);
nand U40263 (N_40263,N_38947,N_38206);
nor U40264 (N_40264,N_38254,N_39667);
nor U40265 (N_40265,N_39055,N_38302);
nor U40266 (N_40266,N_38616,N_38382);
and U40267 (N_40267,N_39367,N_39532);
xor U40268 (N_40268,N_39419,N_39120);
nor U40269 (N_40269,N_38448,N_38439);
and U40270 (N_40270,N_38757,N_38271);
xnor U40271 (N_40271,N_39511,N_38524);
nor U40272 (N_40272,N_38646,N_38119);
nor U40273 (N_40273,N_38096,N_38180);
nand U40274 (N_40274,N_38987,N_38381);
nand U40275 (N_40275,N_38897,N_38970);
nor U40276 (N_40276,N_38252,N_39064);
and U40277 (N_40277,N_39936,N_38614);
or U40278 (N_40278,N_39899,N_39678);
nor U40279 (N_40279,N_39245,N_38050);
nand U40280 (N_40280,N_39606,N_39017);
nand U40281 (N_40281,N_38222,N_39803);
or U40282 (N_40282,N_38000,N_39919);
and U40283 (N_40283,N_39926,N_39888);
nand U40284 (N_40284,N_38299,N_39628);
nand U40285 (N_40285,N_39366,N_39172);
nor U40286 (N_40286,N_38005,N_38176);
xnor U40287 (N_40287,N_39622,N_38794);
and U40288 (N_40288,N_38742,N_38244);
nor U40289 (N_40289,N_39908,N_39602);
or U40290 (N_40290,N_39448,N_38182);
nand U40291 (N_40291,N_39923,N_39287);
xnor U40292 (N_40292,N_38847,N_39934);
or U40293 (N_40293,N_39554,N_38351);
or U40294 (N_40294,N_38332,N_38632);
and U40295 (N_40295,N_38843,N_38212);
and U40296 (N_40296,N_38775,N_38361);
and U40297 (N_40297,N_39897,N_39568);
or U40298 (N_40298,N_39161,N_39688);
and U40299 (N_40299,N_38345,N_39105);
nor U40300 (N_40300,N_39780,N_38585);
xnor U40301 (N_40301,N_39722,N_38044);
nor U40302 (N_40302,N_38168,N_39674);
and U40303 (N_40303,N_39654,N_38458);
xnor U40304 (N_40304,N_38164,N_38030);
or U40305 (N_40305,N_39716,N_39566);
nor U40306 (N_40306,N_38094,N_38489);
and U40307 (N_40307,N_39333,N_38549);
xnor U40308 (N_40308,N_39271,N_38567);
or U40309 (N_40309,N_38224,N_38372);
xnor U40310 (N_40310,N_38805,N_39501);
nor U40311 (N_40311,N_39493,N_39336);
nor U40312 (N_40312,N_39417,N_38786);
xnor U40313 (N_40313,N_38365,N_39181);
nor U40314 (N_40314,N_38116,N_38782);
nand U40315 (N_40315,N_39796,N_38194);
or U40316 (N_40316,N_38937,N_38640);
or U40317 (N_40317,N_38768,N_39272);
nor U40318 (N_40318,N_39912,N_39192);
and U40319 (N_40319,N_38262,N_39403);
nand U40320 (N_40320,N_39084,N_38880);
nand U40321 (N_40321,N_39744,N_38230);
nand U40322 (N_40322,N_38893,N_38126);
xor U40323 (N_40323,N_39410,N_39527);
or U40324 (N_40324,N_38464,N_38417);
nor U40325 (N_40325,N_39955,N_39078);
and U40326 (N_40326,N_38420,N_39095);
xnor U40327 (N_40327,N_38280,N_38586);
and U40328 (N_40328,N_38338,N_39239);
or U40329 (N_40329,N_38691,N_39684);
or U40330 (N_40330,N_39100,N_38066);
nand U40331 (N_40331,N_38919,N_39045);
nor U40332 (N_40332,N_38902,N_39966);
nand U40333 (N_40333,N_39285,N_39605);
nor U40334 (N_40334,N_38690,N_39217);
nand U40335 (N_40335,N_38151,N_38155);
nand U40336 (N_40336,N_38097,N_38136);
nor U40337 (N_40337,N_39922,N_39418);
and U40338 (N_40338,N_39240,N_38868);
and U40339 (N_40339,N_39689,N_39944);
and U40340 (N_40340,N_39302,N_38076);
or U40341 (N_40341,N_39642,N_39659);
nand U40342 (N_40342,N_38279,N_38473);
and U40343 (N_40343,N_38386,N_38546);
or U40344 (N_40344,N_39396,N_38257);
xor U40345 (N_40345,N_38669,N_39300);
and U40346 (N_40346,N_39825,N_38808);
nand U40347 (N_40347,N_39315,N_38982);
and U40348 (N_40348,N_38763,N_39792);
nor U40349 (N_40349,N_38186,N_38322);
or U40350 (N_40350,N_39608,N_39284);
xnor U40351 (N_40351,N_38398,N_39486);
nor U40352 (N_40352,N_38656,N_39231);
nand U40353 (N_40353,N_39159,N_39303);
or U40354 (N_40354,N_39852,N_38402);
or U40355 (N_40355,N_38701,N_38641);
nor U40356 (N_40356,N_39144,N_38476);
xnor U40357 (N_40357,N_39030,N_38840);
and U40358 (N_40358,N_39828,N_39008);
nor U40359 (N_40359,N_39827,N_38029);
or U40360 (N_40360,N_38296,N_38085);
or U40361 (N_40361,N_38943,N_38485);
xnor U40362 (N_40362,N_39885,N_39867);
or U40363 (N_40363,N_39541,N_38541);
nand U40364 (N_40364,N_38255,N_38667);
and U40365 (N_40365,N_38272,N_39952);
nor U40366 (N_40366,N_39443,N_39236);
xnor U40367 (N_40367,N_39508,N_39035);
or U40368 (N_40368,N_39374,N_38359);
and U40369 (N_40369,N_38405,N_39208);
nand U40370 (N_40370,N_39879,N_39909);
nand U40371 (N_40371,N_39986,N_39640);
and U40372 (N_40372,N_39297,N_38131);
and U40373 (N_40373,N_39581,N_39392);
nand U40374 (N_40374,N_38150,N_39173);
or U40375 (N_40375,N_39453,N_39945);
and U40376 (N_40376,N_38555,N_39627);
xor U40377 (N_40377,N_39461,N_38877);
nand U40378 (N_40378,N_39743,N_39497);
or U40379 (N_40379,N_38333,N_38343);
xor U40380 (N_40380,N_38855,N_38630);
or U40381 (N_40381,N_38456,N_39023);
xor U40382 (N_40382,N_38241,N_38120);
nor U40383 (N_40383,N_39709,N_38568);
or U40384 (N_40384,N_39771,N_39465);
and U40385 (N_40385,N_38436,N_39967);
nor U40386 (N_40386,N_38750,N_39383);
and U40387 (N_40387,N_39609,N_39338);
or U40388 (N_40388,N_38487,N_39370);
xnor U40389 (N_40389,N_39594,N_39170);
and U40390 (N_40390,N_39964,N_38218);
nand U40391 (N_40391,N_39993,N_38079);
nor U40392 (N_40392,N_38953,N_38820);
nand U40393 (N_40393,N_39649,N_38086);
xnor U40394 (N_40394,N_38440,N_38346);
or U40395 (N_40395,N_39052,N_39892);
xor U40396 (N_40396,N_39824,N_39656);
xor U40397 (N_40397,N_38089,N_39147);
and U40398 (N_40398,N_38507,N_39262);
or U40399 (N_40399,N_38284,N_38777);
and U40400 (N_40400,N_38127,N_39755);
or U40401 (N_40401,N_38611,N_39307);
nor U40402 (N_40402,N_38844,N_38992);
or U40403 (N_40403,N_38766,N_39858);
or U40404 (N_40404,N_39960,N_39006);
and U40405 (N_40405,N_39820,N_39948);
and U40406 (N_40406,N_38625,N_39176);
or U40407 (N_40407,N_39049,N_38711);
xnor U40408 (N_40408,N_38169,N_38509);
xor U40409 (N_40409,N_39756,N_38354);
xnor U40410 (N_40410,N_39863,N_38134);
nor U40411 (N_40411,N_39742,N_38666);
and U40412 (N_40412,N_39346,N_38959);
or U40413 (N_40413,N_39612,N_38769);
nor U40414 (N_40414,N_38368,N_39668);
or U40415 (N_40415,N_39188,N_39561);
nor U40416 (N_40416,N_38787,N_38629);
nor U40417 (N_40417,N_38547,N_38022);
xor U40418 (N_40418,N_39411,N_39799);
nor U40419 (N_40419,N_38228,N_38748);
and U40420 (N_40420,N_38203,N_39718);
and U40421 (N_40421,N_39676,N_39483);
nor U40422 (N_40422,N_38250,N_39394);
and U40423 (N_40423,N_39791,N_38883);
nand U40424 (N_40424,N_38773,N_38141);
or U40425 (N_40425,N_38377,N_39487);
nor U40426 (N_40426,N_39076,N_39539);
nor U40427 (N_40427,N_39787,N_38687);
and U40428 (N_40428,N_39013,N_38310);
nor U40429 (N_40429,N_38269,N_39514);
and U40430 (N_40430,N_39988,N_38498);
or U40431 (N_40431,N_38154,N_39134);
xor U40432 (N_40432,N_39379,N_38098);
nor U40433 (N_40433,N_39557,N_38871);
or U40434 (N_40434,N_39632,N_38041);
nand U40435 (N_40435,N_39915,N_38655);
and U40436 (N_40436,N_39057,N_39469);
nand U40437 (N_40437,N_39273,N_39071);
nand U40438 (N_40438,N_38971,N_39512);
nor U40439 (N_40439,N_38198,N_39496);
nand U40440 (N_40440,N_38949,N_39701);
or U40441 (N_40441,N_38791,N_39585);
and U40442 (N_40442,N_38665,N_39774);
nor U40443 (N_40443,N_38996,N_38274);
nor U40444 (N_40444,N_39547,N_38952);
or U40445 (N_40445,N_38565,N_38227);
or U40446 (N_40446,N_39840,N_38431);
nor U40447 (N_40447,N_38484,N_39623);
or U40448 (N_40448,N_39137,N_38404);
and U40449 (N_40449,N_39313,N_38685);
nand U40450 (N_40450,N_39003,N_38454);
nand U40451 (N_40451,N_38383,N_39093);
nor U40452 (N_40452,N_39225,N_39761);
and U40453 (N_40453,N_38047,N_38336);
nand U40454 (N_40454,N_39752,N_38950);
nand U40455 (N_40455,N_38392,N_38472);
xnor U40456 (N_40456,N_38138,N_38522);
xnor U40457 (N_40457,N_39878,N_39725);
nand U40458 (N_40458,N_39998,N_38276);
xnor U40459 (N_40459,N_38216,N_38295);
or U40460 (N_40460,N_38845,N_38435);
or U40461 (N_40461,N_39012,N_38023);
nand U40462 (N_40462,N_38842,N_38973);
xnor U40463 (N_40463,N_39671,N_39254);
nand U40464 (N_40464,N_38450,N_39382);
or U40465 (N_40465,N_39712,N_38165);
nand U40466 (N_40466,N_38342,N_39331);
and U40467 (N_40467,N_38574,N_39319);
nand U40468 (N_40468,N_39772,N_39822);
or U40469 (N_40469,N_39014,N_38289);
xnor U40470 (N_40470,N_38718,N_39022);
nor U40471 (N_40471,N_39408,N_39525);
or U40472 (N_40472,N_38379,N_39399);
xnor U40473 (N_40473,N_38500,N_39449);
and U40474 (N_40474,N_38980,N_39516);
and U40475 (N_40475,N_39918,N_38976);
nand U40476 (N_40476,N_39427,N_38770);
or U40477 (N_40477,N_39478,N_39995);
or U40478 (N_40478,N_39222,N_39687);
and U40479 (N_40479,N_38366,N_38698);
and U40480 (N_40480,N_39187,N_38207);
and U40481 (N_40481,N_39959,N_38424);
xor U40482 (N_40482,N_39127,N_39389);
nand U40483 (N_40483,N_39846,N_39528);
or U40484 (N_40484,N_38815,N_38801);
or U40485 (N_40485,N_39706,N_39498);
nor U40486 (N_40486,N_38457,N_38776);
xnor U40487 (N_40487,N_38874,N_38590);
nand U40488 (N_40488,N_38412,N_39895);
nor U40489 (N_40489,N_38866,N_38340);
or U40490 (N_40490,N_38525,N_38810);
and U40491 (N_40491,N_39618,N_38539);
nand U40492 (N_40492,N_38746,N_38562);
xor U40493 (N_40493,N_39662,N_38401);
and U40494 (N_40494,N_39670,N_39645);
xor U40495 (N_40495,N_38290,N_38045);
xnor U40496 (N_40496,N_39378,N_39558);
and U40497 (N_40497,N_39708,N_38018);
nand U40498 (N_40498,N_39738,N_38622);
xnor U40499 (N_40499,N_38652,N_38764);
or U40500 (N_40500,N_38699,N_39129);
and U40501 (N_40501,N_39759,N_39664);
and U40502 (N_40502,N_38587,N_39434);
xor U40503 (N_40503,N_38394,N_39139);
nor U40504 (N_40504,N_39368,N_38660);
or U40505 (N_40505,N_39979,N_39573);
or U40506 (N_40506,N_38760,N_38939);
nand U40507 (N_40507,N_38152,N_38563);
xor U40508 (N_40508,N_39112,N_38631);
xnor U40509 (N_40509,N_39506,N_39800);
nand U40510 (N_40510,N_39310,N_39138);
nor U40511 (N_40511,N_39665,N_38111);
xnor U40512 (N_40512,N_38720,N_39685);
xnor U40513 (N_40513,N_39037,N_38495);
xnor U40514 (N_40514,N_38191,N_39309);
xor U40515 (N_40515,N_39412,N_39146);
nor U40516 (N_40516,N_39421,N_39451);
nand U40517 (N_40517,N_39715,N_38957);
nor U40518 (N_40518,N_39724,N_39556);
nor U40519 (N_40519,N_39094,N_38906);
and U40520 (N_40520,N_38429,N_38077);
and U40521 (N_40521,N_39067,N_39500);
nor U40522 (N_40522,N_39705,N_39243);
nor U40523 (N_40523,N_38173,N_38451);
or U40524 (N_40524,N_38712,N_38602);
xor U40525 (N_40525,N_38807,N_38968);
xnor U40526 (N_40526,N_39351,N_39686);
nor U40527 (N_40527,N_39007,N_39207);
and U40528 (N_40528,N_38008,N_38430);
nor U40529 (N_40529,N_39340,N_39518);
and U40530 (N_40530,N_38977,N_38158);
and U40531 (N_40531,N_39059,N_39677);
and U40532 (N_40532,N_38538,N_38651);
nor U40533 (N_40533,N_38928,N_39795);
or U40534 (N_40534,N_38298,N_38021);
or U40535 (N_40535,N_39790,N_38938);
and U40536 (N_40536,N_39435,N_39849);
nor U40537 (N_40537,N_38946,N_39666);
xnor U40538 (N_40538,N_39591,N_39296);
nor U40539 (N_40539,N_39133,N_39235);
nand U40540 (N_40540,N_38400,N_38390);
and U40541 (N_40541,N_38612,N_39060);
or U40542 (N_40542,N_39713,N_39450);
and U40543 (N_40543,N_38864,N_38817);
nand U40544 (N_40544,N_39736,N_39477);
and U40545 (N_40545,N_39234,N_39371);
or U40546 (N_40546,N_39737,N_38528);
nor U40547 (N_40547,N_38190,N_38293);
and U40548 (N_40548,N_39335,N_39341);
and U40549 (N_40549,N_38995,N_38175);
xor U40550 (N_40550,N_38496,N_39125);
nor U40551 (N_40551,N_39111,N_39326);
nor U40552 (N_40552,N_39940,N_38174);
nand U40553 (N_40553,N_39968,N_39381);
nor U40554 (N_40554,N_38979,N_39931);
xor U40555 (N_40555,N_39248,N_39850);
or U40556 (N_40556,N_39777,N_39031);
and U40557 (N_40557,N_39929,N_38584);
and U40558 (N_40558,N_39428,N_38273);
nor U40559 (N_40559,N_38115,N_39016);
nand U40560 (N_40560,N_39376,N_38017);
xnor U40561 (N_40561,N_38752,N_38869);
or U40562 (N_40562,N_39459,N_39096);
and U40563 (N_40563,N_39631,N_39416);
or U40564 (N_40564,N_38486,N_38109);
nand U40565 (N_40565,N_38261,N_39107);
xnor U40566 (N_40566,N_39582,N_38197);
and U40567 (N_40567,N_39894,N_39075);
nor U40568 (N_40568,N_38609,N_39540);
xnor U40569 (N_40569,N_39179,N_38231);
and U40570 (N_40570,N_38533,N_39005);
and U40571 (N_40571,N_38529,N_39242);
nor U40572 (N_40572,N_38268,N_38785);
and U40573 (N_40573,N_38588,N_39681);
nand U40574 (N_40574,N_38648,N_38682);
and U40575 (N_40575,N_38445,N_38798);
and U40576 (N_40576,N_39066,N_38062);
nor U40577 (N_40577,N_38758,N_38607);
or U40578 (N_40578,N_39424,N_38433);
xor U40579 (N_40579,N_39835,N_39826);
nand U40580 (N_40580,N_38774,N_38680);
xor U40581 (N_40581,N_39887,N_38413);
xor U40582 (N_40582,N_38441,N_39387);
or U40583 (N_40583,N_38039,N_39400);
nor U40584 (N_40584,N_39999,N_39344);
xor U40585 (N_40585,N_39741,N_39463);
and U40586 (N_40586,N_39404,N_39950);
and U40587 (N_40587,N_39749,N_39870);
nor U40588 (N_40588,N_39259,N_39655);
xnor U40589 (N_40589,N_38556,N_38739);
or U40590 (N_40590,N_39135,N_38121);
and U40591 (N_40591,N_38677,N_38028);
or U40592 (N_40592,N_39198,N_39731);
or U40593 (N_40593,N_39981,N_38778);
nor U40594 (N_40594,N_39205,N_38724);
nand U40595 (N_40595,N_38826,N_39559);
and U40596 (N_40596,N_38781,N_39789);
nor U40597 (N_40597,N_38065,N_38105);
or U40598 (N_40598,N_39033,N_38344);
and U40599 (N_40599,N_39578,N_38924);
nor U40600 (N_40600,N_39011,N_39526);
and U40601 (N_40601,N_38589,N_38576);
and U40602 (N_40602,N_39861,N_38886);
or U40603 (N_40603,N_39323,N_38578);
nand U40604 (N_40604,N_38478,N_38499);
or U40605 (N_40605,N_38580,N_39032);
or U40606 (N_40606,N_39260,N_39321);
or U40607 (N_40607,N_38730,N_39148);
nor U40608 (N_40608,N_38819,N_39763);
xnor U40609 (N_40609,N_39550,N_39727);
xor U40610 (N_40610,N_38492,N_39160);
and U40611 (N_40611,N_39956,N_38813);
or U40612 (N_40612,N_38966,N_38449);
xor U40613 (N_40613,N_38370,N_39357);
xor U40614 (N_40614,N_38829,N_39036);
and U40615 (N_40615,N_38315,N_38755);
nor U40616 (N_40616,N_39200,N_38931);
xor U40617 (N_40617,N_38341,N_39839);
or U40618 (N_40618,N_38217,N_38935);
xnor U40619 (N_40619,N_39488,N_38461);
nand U40620 (N_40620,N_38909,N_39592);
and U40621 (N_40621,N_38636,N_39758);
and U40622 (N_40622,N_38288,N_39316);
or U40623 (N_40623,N_38933,N_39572);
or U40624 (N_40624,N_38923,N_38006);
and U40625 (N_40625,N_38316,N_38993);
or U40626 (N_40626,N_38654,N_38542);
nor U40627 (N_40627,N_38016,N_39086);
nand U40628 (N_40628,N_38661,N_38380);
nor U40629 (N_40629,N_39896,N_39402);
and U40630 (N_40630,N_39024,N_38572);
nand U40631 (N_40631,N_38792,N_39750);
or U40632 (N_40632,N_39980,N_38833);
or U40633 (N_40633,N_39130,N_38148);
xnor U40634 (N_40634,N_39650,N_39797);
nand U40635 (N_40635,N_39328,N_39089);
or U40636 (N_40636,N_39740,N_39717);
and U40637 (N_40637,N_39983,N_38623);
nor U40638 (N_40638,N_39904,N_39985);
nor U40639 (N_40639,N_39294,N_38112);
nor U40640 (N_40640,N_38772,N_39099);
or U40641 (N_40641,N_38827,N_38304);
nor U40642 (N_40642,N_38504,N_39295);
nand U40643 (N_40643,N_38841,N_39386);
or U40644 (N_40644,N_39697,N_39745);
and U40645 (N_40645,N_39754,N_39063);
nor U40646 (N_40646,N_39441,N_39916);
and U40647 (N_40647,N_38670,N_38301);
and U40648 (N_40648,N_38723,N_39651);
nand U40649 (N_40649,N_38617,N_38591);
and U40650 (N_40650,N_38561,N_39009);
nand U40651 (N_40651,N_38721,N_38836);
nor U40652 (N_40652,N_38668,N_38517);
nor U40653 (N_40653,N_38540,N_38673);
nor U40654 (N_40654,N_39118,N_39958);
and U40655 (N_40655,N_39485,N_38263);
nand U40656 (N_40656,N_38221,N_39472);
nand U40657 (N_40657,N_38940,N_38601);
nand U40658 (N_40658,N_38291,N_38184);
xor U40659 (N_40659,N_39455,N_39781);
nor U40660 (N_40660,N_39692,N_39021);
nand U40661 (N_40661,N_39811,N_39390);
and U40662 (N_40662,N_39264,N_39881);
nor U40663 (N_40663,N_38513,N_38491);
and U40664 (N_40664,N_39230,N_39070);
nand U40665 (N_40665,N_38452,N_38932);
or U40666 (N_40666,N_39039,N_38520);
xor U40667 (N_40667,N_39874,N_38107);
nand U40668 (N_40668,N_39218,N_39920);
and U40669 (N_40669,N_38510,N_38057);
or U40670 (N_40670,N_38848,N_38865);
and U40671 (N_40671,N_39862,N_38225);
nor U40672 (N_40672,N_39890,N_39121);
nor U40673 (N_40673,N_38814,N_39175);
xor U40674 (N_40674,N_38978,N_39481);
and U40675 (N_40675,N_38942,N_39116);
and U40676 (N_40676,N_39249,N_39268);
nand U40677 (N_40677,N_38463,N_39339);
nor U40678 (N_40678,N_39877,N_38901);
nand U40679 (N_40679,N_38012,N_39203);
nor U40680 (N_40680,N_39553,N_38697);
and U40681 (N_40681,N_39580,N_38550);
or U40682 (N_40682,N_39304,N_38516);
xor U40683 (N_40683,N_38954,N_38916);
nand U40684 (N_40684,N_38892,N_38455);
nand U40685 (N_40685,N_38830,N_39250);
nor U40686 (N_40686,N_38172,N_39994);
nand U40687 (N_40687,N_39728,N_38052);
and U40688 (N_40688,N_39726,N_39760);
nand U40689 (N_40689,N_38211,N_38411);
xor U40690 (N_40690,N_39393,N_39542);
or U40691 (N_40691,N_38852,N_39185);
xor U40692 (N_40692,N_39776,N_38149);
and U40693 (N_40693,N_39823,N_38713);
nor U40694 (N_40694,N_38442,N_39830);
nor U40695 (N_40695,N_38559,N_38745);
or U40696 (N_40696,N_38647,N_39996);
or U40697 (N_40697,N_38494,N_38799);
nand U40698 (N_40698,N_39027,N_39757);
nand U40699 (N_40699,N_38941,N_38679);
and U40700 (N_40700,N_38465,N_38754);
or U40701 (N_40701,N_39375,N_38859);
nand U40702 (N_40702,N_38090,N_38900);
nand U40703 (N_40703,N_39793,N_39050);
or U40704 (N_40704,N_39927,N_38319);
and U40705 (N_40705,N_39597,N_39474);
and U40706 (N_40706,N_39088,N_38615);
xor U40707 (N_40707,N_38393,N_38882);
nand U40708 (N_40708,N_39475,N_39565);
nor U40709 (N_40709,N_39369,N_39334);
xnor U40710 (N_40710,N_39951,N_38727);
nand U40711 (N_40711,N_38566,N_39812);
nand U40712 (N_40712,N_39509,N_38460);
and U40713 (N_40713,N_38469,N_39342);
and U40714 (N_40714,N_39935,N_39291);
xnor U40715 (N_40715,N_39868,N_39436);
xnor U40716 (N_40716,N_38557,N_39704);
nor U40717 (N_40717,N_38303,N_39266);
nor U40718 (N_40718,N_39521,N_38053);
or U40719 (N_40719,N_39471,N_39458);
xor U40720 (N_40720,N_38628,N_39432);
or U40721 (N_40721,N_39699,N_38965);
xnor U40722 (N_40722,N_39004,N_38771);
nor U40723 (N_40723,N_39595,N_38132);
nor U40724 (N_40724,N_39286,N_38907);
nor U40725 (N_40725,N_38853,N_39661);
nor U40726 (N_40726,N_38634,N_39992);
nor U40727 (N_40727,N_39305,N_39290);
or U40728 (N_40728,N_38425,N_38851);
xnor U40729 (N_40729,N_38282,N_39080);
nor U40730 (N_40730,N_38831,N_38570);
and U40731 (N_40731,N_39767,N_38407);
or U40732 (N_40732,N_39971,N_39548);
nor U40733 (N_40733,N_38593,N_38278);
or U40734 (N_40734,N_39216,N_38964);
or U40735 (N_40735,N_39241,N_39104);
and U40736 (N_40736,N_38235,N_39482);
nor U40737 (N_40737,N_38915,N_39197);
xor U40738 (N_40738,N_39178,N_38875);
and U40739 (N_40739,N_38553,N_38579);
or U40740 (N_40740,N_39289,N_39730);
xor U40741 (N_40741,N_38453,N_38795);
and U40742 (N_40742,N_39265,N_38106);
nor U40743 (N_40743,N_39751,N_39042);
nand U40744 (N_40744,N_38663,N_38355);
xor U40745 (N_40745,N_38870,N_39802);
xor U40746 (N_40746,N_39466,N_39544);
nor U40747 (N_40747,N_38903,N_38867);
or U40748 (N_40748,N_38226,N_39140);
or U40749 (N_40749,N_39153,N_38862);
nand U40750 (N_40750,N_39051,N_38025);
or U40751 (N_40751,N_38639,N_38432);
xnor U40752 (N_40752,N_38102,N_39163);
nor U40753 (N_40753,N_39131,N_38508);
nand U40754 (N_40754,N_39970,N_38414);
and U40755 (N_40755,N_39117,N_39214);
and U40756 (N_40756,N_39048,N_38334);
or U40757 (N_40757,N_38337,N_38129);
or U40758 (N_40758,N_39535,N_38171);
nor U40759 (N_40759,N_39077,N_38644);
nor U40760 (N_40760,N_38926,N_38070);
xor U40761 (N_40761,N_39616,N_38038);
nand U40762 (N_40762,N_39444,N_38714);
and U40763 (N_40763,N_38325,N_39638);
or U40764 (N_40764,N_38055,N_38997);
xor U40765 (N_40765,N_38422,N_39081);
and U40766 (N_40766,N_38828,N_38232);
xnor U40767 (N_40767,N_38427,N_38387);
nand U40768 (N_40768,N_38426,N_38081);
or U40769 (N_40769,N_39832,N_39246);
nand U40770 (N_40770,N_39298,N_38518);
and U40771 (N_40771,N_39347,N_39906);
and U40772 (N_40772,N_39202,N_38734);
and U40773 (N_40773,N_38199,N_39902);
nor U40774 (N_40774,N_39480,N_38686);
or U40775 (N_40775,N_38060,N_38374);
or U40776 (N_40776,N_38072,N_39479);
nand U40777 (N_40777,N_38446,N_39576);
nor U40778 (N_40778,N_39108,N_39308);
or U40779 (N_40779,N_38350,N_39603);
nand U40780 (N_40780,N_39898,N_38912);
xor U40781 (N_40781,N_39034,N_39575);
and U40782 (N_40782,N_39523,N_38242);
xor U40783 (N_40783,N_38708,N_38554);
nand U40784 (N_40784,N_38737,N_39961);
and U40785 (N_40785,N_38596,N_39258);
or U40786 (N_40786,N_38093,N_39530);
or U40787 (N_40787,N_38592,N_39786);
and U40788 (N_40788,N_38497,N_39210);
xor U40789 (N_40789,N_38832,N_39002);
xnor U40790 (N_40790,N_38854,N_38147);
and U40791 (N_40791,N_38418,N_39040);
nor U40792 (N_40792,N_39834,N_38099);
nand U40793 (N_40793,N_39905,N_39372);
nand U40794 (N_40794,N_39124,N_39765);
nor U40795 (N_40795,N_38092,N_39907);
xor U40796 (N_40796,N_39810,N_39634);
or U40797 (N_40797,N_38468,N_39886);
xnor U40798 (N_40798,N_38535,N_39587);
or U40799 (N_40799,N_39269,N_38396);
nor U40800 (N_40800,N_39837,N_39182);
xnor U40801 (N_40801,N_38283,N_38371);
nand U40802 (N_40802,N_39819,N_39356);
nand U40803 (N_40803,N_38879,N_38416);
or U40804 (N_40804,N_39630,N_39312);
nor U40805 (N_40805,N_38613,N_38213);
or U40806 (N_40806,N_38409,N_39515);
xor U40807 (N_40807,N_39407,N_38837);
and U40808 (N_40808,N_39122,N_39423);
and U40809 (N_40809,N_38358,N_39963);
xnor U40810 (N_40810,N_39954,N_39362);
and U40811 (N_40811,N_38521,N_39327);
xnor U40812 (N_40812,N_38027,N_39430);
nor U40813 (N_40813,N_39962,N_39593);
or U40814 (N_40814,N_39384,N_38917);
xnor U40815 (N_40815,N_38582,N_39723);
nand U40816 (N_40816,N_38397,N_39579);
nor U40817 (N_40817,N_38317,N_38188);
nor U40818 (N_40818,N_39933,N_39529);
or U40819 (N_40819,N_39317,N_38605);
and U40820 (N_40820,N_39693,N_38986);
xor U40821 (N_40821,N_38087,N_38887);
or U40822 (N_40822,N_39350,N_38675);
nor U40823 (N_40823,N_39190,N_38600);
or U40824 (N_40824,N_39921,N_39010);
or U40825 (N_40825,N_38558,N_39150);
or U40826 (N_40826,N_39038,N_38286);
xnor U40827 (N_40827,N_38863,N_38678);
nor U40828 (N_40828,N_39132,N_38519);
nand U40829 (N_40829,N_39363,N_39164);
or U40830 (N_40830,N_38388,N_39769);
and U40831 (N_40831,N_38084,N_38681);
and U40832 (N_40832,N_39519,N_39773);
or U40833 (N_40833,N_38474,N_39702);
or U40834 (N_40834,N_38702,N_38505);
nand U40835 (N_40835,N_38571,N_39373);
or U40836 (N_40836,N_38477,N_39534);
nand U40837 (N_40837,N_39169,N_38220);
nor U40838 (N_40838,N_39329,N_38649);
nand U40839 (N_40839,N_39255,N_39414);
xnor U40840 (N_40840,N_39690,N_38929);
nand U40841 (N_40841,N_39126,N_38548);
or U40842 (N_40842,N_38731,N_38481);
or U40843 (N_40843,N_39143,N_39091);
xor U40844 (N_40844,N_39101,N_38033);
and U40845 (N_40845,N_38037,N_39517);
and U40846 (N_40846,N_38809,N_39405);
nor U40847 (N_40847,N_38700,N_39252);
nand U40848 (N_40848,N_39401,N_39380);
nand U40849 (N_40849,N_38891,N_38003);
and U40850 (N_40850,N_39707,N_38536);
and U40851 (N_40851,N_38889,N_38314);
and U40852 (N_40852,N_38214,N_39349);
nand U40853 (N_40853,N_38895,N_38577);
xnor U40854 (N_40854,N_39083,N_39257);
xnor U40855 (N_40855,N_38913,N_39869);
xor U40856 (N_40856,N_39657,N_39694);
nand U40857 (N_40857,N_38275,N_39072);
nor U40858 (N_40858,N_39621,N_39853);
and U40859 (N_40859,N_39857,N_38419);
nand U40860 (N_40860,N_38534,N_38229);
nand U40861 (N_40861,N_39103,N_39398);
and U40862 (N_40862,N_38575,N_39174);
nand U40863 (N_40863,N_39735,N_39524);
or U40864 (N_40864,N_38994,N_38856);
nor U40865 (N_40865,N_39984,N_39446);
xnor U40866 (N_40866,N_39976,N_39889);
nor U40867 (N_40867,N_38113,N_39261);
or U40868 (N_40868,N_38945,N_39719);
nand U40869 (N_40869,N_38658,N_38444);
xor U40870 (N_40870,N_38067,N_39682);
or U40871 (N_40871,N_39385,N_39925);
xor U40872 (N_40872,N_38124,N_39025);
and U40873 (N_40873,N_38789,N_38635);
xnor U40874 (N_40874,N_38223,N_39332);
nor U40875 (N_40875,N_39462,N_39494);
and U40876 (N_40876,N_39513,N_39695);
or U40877 (N_40877,N_38642,N_38320);
and U40878 (N_40878,N_38331,N_38308);
xnor U40879 (N_40879,N_38911,N_39142);
nor U40880 (N_40880,N_38741,N_38249);
nor U40881 (N_40881,N_38626,N_39807);
xnor U40882 (N_40882,N_38375,N_38482);
nor U40883 (N_40883,N_38277,N_38619);
nor U40884 (N_40884,N_38068,N_39624);
or U40885 (N_40885,N_38960,N_39942);
nand U40886 (N_40886,N_39106,N_39388);
xnor U40887 (N_40887,N_38662,N_38101);
nor U40888 (N_40888,N_39201,N_39836);
nor U40889 (N_40889,N_39196,N_38391);
or U40890 (N_40890,N_39456,N_38048);
xor U40891 (N_40891,N_38364,N_39020);
nor U40892 (N_40892,N_38193,N_38170);
xnor U40893 (N_40893,N_38043,N_38210);
xnor U40894 (N_40894,N_38285,N_39361);
and U40895 (N_40895,N_38166,N_39633);
xnor U40896 (N_40896,N_39711,N_38300);
and U40897 (N_40897,N_38925,N_39739);
and U40898 (N_40898,N_39672,N_39880);
or U40899 (N_40899,N_39460,N_39876);
nor U40900 (N_40900,N_38258,N_38812);
xnor U40901 (N_40901,N_38610,N_38511);
or U40902 (N_40902,N_39625,N_39330);
nor U40903 (N_40903,N_39505,N_39354);
xnor U40904 (N_40904,N_39596,N_38196);
or U40905 (N_40905,N_39939,N_39520);
or U40906 (N_40906,N_38707,N_39941);
nand U40907 (N_40907,N_38618,N_39283);
xor U40908 (N_40908,N_38918,N_39785);
and U40909 (N_40909,N_39522,N_38885);
or U40910 (N_40910,N_38373,N_39947);
or U40911 (N_40911,N_38324,N_38192);
xnor U40912 (N_40912,N_38347,N_38503);
xor U40913 (N_40913,N_39703,N_38930);
nor U40914 (N_40914,N_39974,N_38564);
xor U40915 (N_40915,N_38725,N_39074);
and U40916 (N_40916,N_38961,N_38237);
and U40917 (N_40917,N_38046,N_39599);
and U40918 (N_40918,N_38779,N_38706);
nor U40919 (N_40919,N_38406,N_38780);
or U40920 (N_40920,N_38415,N_38689);
or U40921 (N_40921,N_39306,N_38189);
or U40922 (N_40922,N_38251,N_38850);
nand U40923 (N_40923,N_38849,N_39875);
or U40924 (N_40924,N_39484,N_38569);
nor U40925 (N_40925,N_39280,N_39211);
nand U40926 (N_40926,N_38114,N_38936);
xor U40927 (N_40927,N_39604,N_38767);
or U40928 (N_40928,N_39325,N_38753);
nor U40929 (N_40929,N_39065,N_38479);
or U40930 (N_40930,N_38001,N_38515);
and U40931 (N_40931,N_38260,N_39166);
xnor U40932 (N_40932,N_38683,N_38793);
or U40933 (N_40933,N_39426,N_38643);
and U40934 (N_40934,N_39691,N_38108);
and U40935 (N_40935,N_39546,N_39355);
or U40936 (N_40936,N_39409,N_38823);
nor U40937 (N_40937,N_39937,N_38297);
xnor U40938 (N_40938,N_39818,N_39352);
xor U40939 (N_40939,N_39533,N_39782);
xnor U40940 (N_40940,N_38362,N_38339);
and U40941 (N_40941,N_39644,N_39276);
or U40942 (N_40942,N_39454,N_39851);
and U40943 (N_40943,N_38975,N_38594);
xor U40944 (N_40944,N_39611,N_39092);
xor U40945 (N_40945,N_39149,N_39015);
xor U40946 (N_40946,N_38004,N_39061);
nor U40947 (N_40947,N_39473,N_38695);
xor U40948 (N_40948,N_39228,N_38816);
and U40949 (N_40949,N_39128,N_38526);
xor U40950 (N_40950,N_39847,N_39195);
nand U40951 (N_40951,N_38811,N_38328);
xor U40952 (N_40952,N_38185,N_38671);
nor U40953 (N_40953,N_38999,N_38091);
nand U40954 (N_40954,N_38061,N_38573);
nand U40955 (N_40955,N_38349,N_38294);
or U40956 (N_40956,N_39215,N_39029);
nand U40957 (N_40957,N_39073,N_38437);
nor U40958 (N_40958,N_38802,N_39629);
and U40959 (N_40959,N_38054,N_38797);
nand U40960 (N_40960,N_38888,N_38313);
and U40961 (N_40961,N_38790,N_39263);
and U40962 (N_40962,N_39499,N_39663);
nor U40963 (N_40963,N_39932,N_38459);
nand U40964 (N_40964,N_39643,N_38110);
or U40965 (N_40965,N_38905,N_39989);
nand U40966 (N_40966,N_39415,N_38751);
nor U40967 (N_40967,N_39000,N_39900);
xnor U40968 (N_40968,N_39358,N_38036);
nor U40969 (N_40969,N_39808,N_38722);
nand U40970 (N_40970,N_39102,N_38934);
nor U40971 (N_40971,N_39353,N_39224);
nand U40972 (N_40972,N_38219,N_39766);
nand U40973 (N_40973,N_39156,N_39930);
and U40974 (N_40974,N_38434,N_38621);
xor U40975 (N_40975,N_39247,N_38183);
and U40976 (N_40976,N_38530,N_39977);
xor U40977 (N_40977,N_38974,N_39220);
nand U40978 (N_40978,N_38633,N_39253);
and U40979 (N_40979,N_38914,N_39229);
or U40980 (N_40980,N_38759,N_38951);
or U40981 (N_40981,N_38595,N_39562);
nor U40982 (N_40982,N_39997,N_39537);
and U40983 (N_40983,N_38747,N_39856);
or U40984 (N_40984,N_39226,N_39227);
nor U40985 (N_40985,N_38506,N_39982);
or U40986 (N_40986,N_39732,N_38163);
nor U40987 (N_40987,N_38825,N_39193);
nor U40988 (N_40988,N_39028,N_39698);
xor U40989 (N_40989,N_38256,N_38032);
and U40990 (N_40990,N_39831,N_38292);
nand U40991 (N_40991,N_38688,N_38080);
nand U40992 (N_40992,N_38133,N_39420);
xor U40993 (N_40993,N_38881,N_38410);
nor U40994 (N_40994,N_39949,N_38904);
nor U40995 (N_40995,N_38672,N_38490);
nor U40996 (N_40996,N_38846,N_39778);
and U40997 (N_40997,N_39293,N_38367);
and U40998 (N_40998,N_39123,N_39062);
and U40999 (N_40999,N_38078,N_39660);
or U41000 (N_41000,N_38231,N_38653);
nand U41001 (N_41001,N_38725,N_39419);
xnor U41002 (N_41002,N_39150,N_38952);
nand U41003 (N_41003,N_39813,N_39978);
xor U41004 (N_41004,N_39227,N_39499);
nor U41005 (N_41005,N_38535,N_39553);
and U41006 (N_41006,N_39854,N_39941);
xor U41007 (N_41007,N_38324,N_39735);
nor U41008 (N_41008,N_39428,N_38412);
xor U41009 (N_41009,N_39190,N_39806);
nor U41010 (N_41010,N_39046,N_39494);
nand U41011 (N_41011,N_39542,N_39766);
nand U41012 (N_41012,N_39559,N_39027);
nand U41013 (N_41013,N_39930,N_38721);
and U41014 (N_41014,N_39584,N_39183);
nor U41015 (N_41015,N_39656,N_39313);
nand U41016 (N_41016,N_38803,N_39243);
or U41017 (N_41017,N_39235,N_39114);
nor U41018 (N_41018,N_38732,N_39095);
nand U41019 (N_41019,N_38842,N_38570);
nand U41020 (N_41020,N_39695,N_39068);
or U41021 (N_41021,N_38390,N_38486);
and U41022 (N_41022,N_39312,N_39537);
nor U41023 (N_41023,N_38622,N_39504);
nor U41024 (N_41024,N_38308,N_39200);
xnor U41025 (N_41025,N_38121,N_39383);
xor U41026 (N_41026,N_38360,N_39958);
nor U41027 (N_41027,N_39033,N_39123);
and U41028 (N_41028,N_38389,N_39983);
nor U41029 (N_41029,N_38756,N_39531);
and U41030 (N_41030,N_39983,N_38557);
nor U41031 (N_41031,N_39942,N_38050);
nand U41032 (N_41032,N_38402,N_39542);
and U41033 (N_41033,N_38209,N_39341);
and U41034 (N_41034,N_38125,N_39794);
xor U41035 (N_41035,N_39462,N_39954);
or U41036 (N_41036,N_39800,N_39251);
and U41037 (N_41037,N_38016,N_38396);
nand U41038 (N_41038,N_38966,N_39773);
xnor U41039 (N_41039,N_38293,N_38189);
and U41040 (N_41040,N_39247,N_38077);
nor U41041 (N_41041,N_38343,N_39384);
nand U41042 (N_41042,N_38586,N_38871);
xnor U41043 (N_41043,N_39479,N_38094);
nor U41044 (N_41044,N_38602,N_39236);
xor U41045 (N_41045,N_39839,N_39899);
nor U41046 (N_41046,N_39711,N_38018);
nand U41047 (N_41047,N_38487,N_38852);
xnor U41048 (N_41048,N_38026,N_38783);
and U41049 (N_41049,N_39693,N_38748);
nor U41050 (N_41050,N_38756,N_38023);
nand U41051 (N_41051,N_39294,N_38079);
nor U41052 (N_41052,N_38384,N_39033);
xor U41053 (N_41053,N_38949,N_38627);
or U41054 (N_41054,N_39631,N_39084);
and U41055 (N_41055,N_38464,N_39743);
nand U41056 (N_41056,N_39892,N_39869);
nor U41057 (N_41057,N_38162,N_39735);
or U41058 (N_41058,N_38304,N_39790);
and U41059 (N_41059,N_39848,N_39605);
or U41060 (N_41060,N_38747,N_38640);
or U41061 (N_41061,N_39522,N_38543);
or U41062 (N_41062,N_39032,N_38861);
nand U41063 (N_41063,N_38310,N_39206);
and U41064 (N_41064,N_39571,N_39382);
and U41065 (N_41065,N_39781,N_38404);
or U41066 (N_41066,N_39752,N_39898);
and U41067 (N_41067,N_39725,N_39883);
nand U41068 (N_41068,N_39857,N_39338);
and U41069 (N_41069,N_38207,N_39759);
xor U41070 (N_41070,N_38865,N_38447);
nand U41071 (N_41071,N_38800,N_39624);
or U41072 (N_41072,N_38495,N_39959);
xnor U41073 (N_41073,N_39793,N_38515);
or U41074 (N_41074,N_39356,N_39237);
nand U41075 (N_41075,N_38385,N_39272);
or U41076 (N_41076,N_39042,N_38509);
or U41077 (N_41077,N_39069,N_38540);
nand U41078 (N_41078,N_39177,N_39503);
and U41079 (N_41079,N_38465,N_39682);
nor U41080 (N_41080,N_38116,N_39019);
nand U41081 (N_41081,N_39303,N_38963);
or U41082 (N_41082,N_38482,N_38931);
and U41083 (N_41083,N_38976,N_39042);
nor U41084 (N_41084,N_38169,N_39672);
nor U41085 (N_41085,N_39422,N_38222);
nor U41086 (N_41086,N_38270,N_39032);
and U41087 (N_41087,N_38449,N_39189);
or U41088 (N_41088,N_38590,N_39896);
xor U41089 (N_41089,N_38791,N_38276);
nor U41090 (N_41090,N_39765,N_39146);
nor U41091 (N_41091,N_39029,N_38245);
or U41092 (N_41092,N_39325,N_38641);
and U41093 (N_41093,N_38832,N_38375);
nor U41094 (N_41094,N_38182,N_38880);
nand U41095 (N_41095,N_38648,N_39055);
nor U41096 (N_41096,N_38156,N_39782);
xnor U41097 (N_41097,N_38692,N_38488);
nor U41098 (N_41098,N_39132,N_39419);
nor U41099 (N_41099,N_38324,N_38920);
and U41100 (N_41100,N_38122,N_39776);
nor U41101 (N_41101,N_39546,N_38400);
xor U41102 (N_41102,N_38226,N_38856);
xnor U41103 (N_41103,N_39632,N_39553);
nand U41104 (N_41104,N_39886,N_39664);
nand U41105 (N_41105,N_38743,N_38890);
nand U41106 (N_41106,N_38290,N_38952);
or U41107 (N_41107,N_39476,N_39439);
or U41108 (N_41108,N_38536,N_39056);
nor U41109 (N_41109,N_38092,N_39913);
or U41110 (N_41110,N_38767,N_39767);
nor U41111 (N_41111,N_38834,N_39032);
or U41112 (N_41112,N_38137,N_38434);
xnor U41113 (N_41113,N_38604,N_38529);
nor U41114 (N_41114,N_38988,N_38436);
xnor U41115 (N_41115,N_39497,N_38933);
xnor U41116 (N_41116,N_38411,N_39571);
xor U41117 (N_41117,N_39291,N_38971);
or U41118 (N_41118,N_39615,N_39021);
nor U41119 (N_41119,N_38254,N_39170);
and U41120 (N_41120,N_39488,N_39528);
or U41121 (N_41121,N_38915,N_39456);
and U41122 (N_41122,N_39593,N_38559);
or U41123 (N_41123,N_38129,N_39187);
or U41124 (N_41124,N_39455,N_39093);
nor U41125 (N_41125,N_39296,N_38823);
nand U41126 (N_41126,N_39417,N_38099);
or U41127 (N_41127,N_39874,N_38886);
nand U41128 (N_41128,N_39614,N_39021);
nand U41129 (N_41129,N_39207,N_38178);
and U41130 (N_41130,N_39604,N_39244);
and U41131 (N_41131,N_38519,N_38180);
or U41132 (N_41132,N_39619,N_38044);
or U41133 (N_41133,N_39957,N_38992);
or U41134 (N_41134,N_39685,N_38536);
nand U41135 (N_41135,N_38709,N_39658);
nor U41136 (N_41136,N_38878,N_38910);
nor U41137 (N_41137,N_38462,N_38337);
nand U41138 (N_41138,N_39143,N_38313);
nand U41139 (N_41139,N_38445,N_38762);
nor U41140 (N_41140,N_38347,N_38420);
or U41141 (N_41141,N_39682,N_39367);
xnor U41142 (N_41142,N_39863,N_39206);
or U41143 (N_41143,N_38146,N_38416);
xor U41144 (N_41144,N_39818,N_38428);
and U41145 (N_41145,N_39193,N_38159);
or U41146 (N_41146,N_38351,N_39940);
nand U41147 (N_41147,N_39434,N_38170);
nor U41148 (N_41148,N_38782,N_38345);
xnor U41149 (N_41149,N_38473,N_39617);
nand U41150 (N_41150,N_39838,N_38976);
and U41151 (N_41151,N_39334,N_38858);
nor U41152 (N_41152,N_39165,N_39651);
and U41153 (N_41153,N_39333,N_39099);
nor U41154 (N_41154,N_38811,N_39557);
nor U41155 (N_41155,N_38545,N_38099);
nor U41156 (N_41156,N_38764,N_38486);
and U41157 (N_41157,N_39893,N_39961);
and U41158 (N_41158,N_38066,N_39532);
xor U41159 (N_41159,N_39549,N_38555);
nor U41160 (N_41160,N_39217,N_39728);
xor U41161 (N_41161,N_39095,N_38407);
nand U41162 (N_41162,N_38815,N_38252);
nor U41163 (N_41163,N_39255,N_39287);
or U41164 (N_41164,N_38956,N_39587);
xnor U41165 (N_41165,N_39456,N_38134);
xor U41166 (N_41166,N_38025,N_38984);
xnor U41167 (N_41167,N_38430,N_38901);
nor U41168 (N_41168,N_38520,N_38079);
xor U41169 (N_41169,N_38846,N_38738);
nand U41170 (N_41170,N_38974,N_38216);
nor U41171 (N_41171,N_38672,N_38891);
or U41172 (N_41172,N_39710,N_39067);
nor U41173 (N_41173,N_38880,N_38029);
nor U41174 (N_41174,N_39751,N_39940);
or U41175 (N_41175,N_39921,N_39610);
xor U41176 (N_41176,N_38106,N_39323);
or U41177 (N_41177,N_39608,N_38556);
or U41178 (N_41178,N_38033,N_38635);
nor U41179 (N_41179,N_38203,N_39418);
nor U41180 (N_41180,N_39468,N_38083);
xor U41181 (N_41181,N_38352,N_39612);
nand U41182 (N_41182,N_38374,N_38774);
nor U41183 (N_41183,N_39247,N_39613);
or U41184 (N_41184,N_39107,N_39562);
nand U41185 (N_41185,N_39355,N_38635);
nand U41186 (N_41186,N_38080,N_38911);
xor U41187 (N_41187,N_38215,N_39521);
nor U41188 (N_41188,N_38187,N_39416);
nor U41189 (N_41189,N_39130,N_38420);
nor U41190 (N_41190,N_39151,N_38472);
and U41191 (N_41191,N_39843,N_38997);
or U41192 (N_41192,N_39415,N_38342);
nand U41193 (N_41193,N_38557,N_39382);
and U41194 (N_41194,N_38198,N_39199);
and U41195 (N_41195,N_38520,N_38513);
or U41196 (N_41196,N_39076,N_39446);
nand U41197 (N_41197,N_38562,N_39820);
and U41198 (N_41198,N_38604,N_38585);
nand U41199 (N_41199,N_38129,N_39259);
or U41200 (N_41200,N_39416,N_38010);
nor U41201 (N_41201,N_39460,N_39034);
or U41202 (N_41202,N_38191,N_39795);
and U41203 (N_41203,N_39417,N_38200);
nand U41204 (N_41204,N_39519,N_39171);
xnor U41205 (N_41205,N_39057,N_38356);
or U41206 (N_41206,N_39848,N_39754);
xnor U41207 (N_41207,N_38392,N_38727);
nor U41208 (N_41208,N_38537,N_38815);
nor U41209 (N_41209,N_38754,N_38628);
or U41210 (N_41210,N_38680,N_39155);
nor U41211 (N_41211,N_38031,N_38629);
xnor U41212 (N_41212,N_38048,N_39176);
nand U41213 (N_41213,N_38903,N_38938);
xnor U41214 (N_41214,N_39751,N_38840);
or U41215 (N_41215,N_39622,N_38691);
or U41216 (N_41216,N_38144,N_38001);
xnor U41217 (N_41217,N_39213,N_39732);
nor U41218 (N_41218,N_39475,N_39733);
nor U41219 (N_41219,N_38865,N_38085);
xnor U41220 (N_41220,N_39951,N_39736);
nand U41221 (N_41221,N_39903,N_38513);
nand U41222 (N_41222,N_38304,N_39060);
nor U41223 (N_41223,N_39898,N_39114);
or U41224 (N_41224,N_39874,N_38543);
xor U41225 (N_41225,N_38759,N_38743);
nand U41226 (N_41226,N_39749,N_38748);
or U41227 (N_41227,N_38172,N_38417);
xnor U41228 (N_41228,N_39464,N_38492);
nor U41229 (N_41229,N_38283,N_39308);
xor U41230 (N_41230,N_38357,N_38673);
and U41231 (N_41231,N_38735,N_38751);
and U41232 (N_41232,N_38549,N_39783);
xor U41233 (N_41233,N_38892,N_38423);
xor U41234 (N_41234,N_39275,N_39527);
nand U41235 (N_41235,N_38781,N_39910);
nor U41236 (N_41236,N_39708,N_38887);
and U41237 (N_41237,N_38856,N_38502);
nand U41238 (N_41238,N_38222,N_38878);
nand U41239 (N_41239,N_39967,N_38525);
nor U41240 (N_41240,N_38957,N_38563);
nor U41241 (N_41241,N_39062,N_38574);
xnor U41242 (N_41242,N_38743,N_39991);
nor U41243 (N_41243,N_38098,N_39538);
or U41244 (N_41244,N_38695,N_38294);
nor U41245 (N_41245,N_39301,N_38944);
and U41246 (N_41246,N_38350,N_39129);
nand U41247 (N_41247,N_39240,N_38837);
nor U41248 (N_41248,N_38562,N_38276);
nand U41249 (N_41249,N_39949,N_38490);
nand U41250 (N_41250,N_38329,N_39492);
nor U41251 (N_41251,N_39453,N_38231);
xnor U41252 (N_41252,N_38482,N_39254);
and U41253 (N_41253,N_39125,N_39622);
and U41254 (N_41254,N_39377,N_38065);
xor U41255 (N_41255,N_39305,N_39489);
xnor U41256 (N_41256,N_38924,N_38161);
nand U41257 (N_41257,N_38285,N_39349);
nand U41258 (N_41258,N_39931,N_39398);
or U41259 (N_41259,N_38148,N_38432);
and U41260 (N_41260,N_38623,N_39668);
or U41261 (N_41261,N_38189,N_38051);
xor U41262 (N_41262,N_39561,N_39123);
xor U41263 (N_41263,N_39647,N_39726);
xnor U41264 (N_41264,N_39492,N_38443);
and U41265 (N_41265,N_39357,N_39210);
nor U41266 (N_41266,N_38611,N_38433);
or U41267 (N_41267,N_38903,N_38629);
xnor U41268 (N_41268,N_38801,N_39867);
nand U41269 (N_41269,N_39678,N_38163);
nor U41270 (N_41270,N_39986,N_39627);
and U41271 (N_41271,N_38988,N_38150);
nand U41272 (N_41272,N_38500,N_38696);
nand U41273 (N_41273,N_39722,N_39032);
xnor U41274 (N_41274,N_38289,N_39294);
or U41275 (N_41275,N_38950,N_39482);
and U41276 (N_41276,N_38597,N_38724);
nor U41277 (N_41277,N_39073,N_39598);
nand U41278 (N_41278,N_39772,N_38353);
or U41279 (N_41279,N_38087,N_39094);
or U41280 (N_41280,N_39497,N_38633);
nand U41281 (N_41281,N_39386,N_38727);
and U41282 (N_41282,N_38198,N_38011);
xor U41283 (N_41283,N_38274,N_39390);
nand U41284 (N_41284,N_39558,N_38717);
nand U41285 (N_41285,N_39318,N_38253);
nor U41286 (N_41286,N_39241,N_39011);
or U41287 (N_41287,N_39688,N_38528);
or U41288 (N_41288,N_39832,N_38341);
or U41289 (N_41289,N_38474,N_38997);
xnor U41290 (N_41290,N_38938,N_38030);
or U41291 (N_41291,N_38949,N_39415);
or U41292 (N_41292,N_38498,N_38381);
xnor U41293 (N_41293,N_38056,N_38938);
and U41294 (N_41294,N_39206,N_38012);
nand U41295 (N_41295,N_38414,N_39204);
or U41296 (N_41296,N_39361,N_39328);
nor U41297 (N_41297,N_39503,N_39915);
xor U41298 (N_41298,N_38695,N_38709);
nand U41299 (N_41299,N_38318,N_38832);
and U41300 (N_41300,N_39818,N_39129);
nor U41301 (N_41301,N_38231,N_39444);
nor U41302 (N_41302,N_38306,N_39169);
nand U41303 (N_41303,N_39282,N_39133);
and U41304 (N_41304,N_38861,N_38811);
and U41305 (N_41305,N_39293,N_39129);
nand U41306 (N_41306,N_39592,N_38105);
xor U41307 (N_41307,N_38349,N_39738);
or U41308 (N_41308,N_38940,N_38502);
or U41309 (N_41309,N_38499,N_38557);
xor U41310 (N_41310,N_38232,N_39678);
or U41311 (N_41311,N_39618,N_38027);
or U41312 (N_41312,N_39306,N_39960);
xor U41313 (N_41313,N_38308,N_39048);
and U41314 (N_41314,N_39766,N_39257);
and U41315 (N_41315,N_38470,N_39423);
nor U41316 (N_41316,N_39795,N_38384);
nand U41317 (N_41317,N_38326,N_39637);
or U41318 (N_41318,N_39891,N_38541);
and U41319 (N_41319,N_38664,N_39485);
or U41320 (N_41320,N_39498,N_38335);
nor U41321 (N_41321,N_39448,N_38075);
xnor U41322 (N_41322,N_38488,N_39130);
nor U41323 (N_41323,N_39825,N_38133);
and U41324 (N_41324,N_38375,N_39791);
nor U41325 (N_41325,N_38426,N_39730);
nand U41326 (N_41326,N_39327,N_38032);
or U41327 (N_41327,N_38392,N_38559);
nand U41328 (N_41328,N_39458,N_39758);
xor U41329 (N_41329,N_38652,N_39011);
xnor U41330 (N_41330,N_39889,N_38429);
xor U41331 (N_41331,N_39781,N_39989);
or U41332 (N_41332,N_39700,N_39178);
and U41333 (N_41333,N_38826,N_38741);
xnor U41334 (N_41334,N_39059,N_39457);
nor U41335 (N_41335,N_38049,N_38692);
and U41336 (N_41336,N_38635,N_39958);
nor U41337 (N_41337,N_38364,N_38766);
nand U41338 (N_41338,N_38156,N_39395);
nand U41339 (N_41339,N_38647,N_39350);
or U41340 (N_41340,N_38758,N_38941);
nand U41341 (N_41341,N_38397,N_39346);
nor U41342 (N_41342,N_38785,N_39130);
nor U41343 (N_41343,N_38983,N_38632);
and U41344 (N_41344,N_39840,N_38422);
or U41345 (N_41345,N_38286,N_38675);
or U41346 (N_41346,N_39178,N_38993);
or U41347 (N_41347,N_38427,N_38946);
and U41348 (N_41348,N_39947,N_38765);
nand U41349 (N_41349,N_39613,N_39220);
and U41350 (N_41350,N_39876,N_39216);
nor U41351 (N_41351,N_39512,N_39285);
xnor U41352 (N_41352,N_39982,N_39758);
nor U41353 (N_41353,N_39005,N_38165);
or U41354 (N_41354,N_39953,N_39702);
or U41355 (N_41355,N_38723,N_38077);
and U41356 (N_41356,N_39576,N_38573);
nor U41357 (N_41357,N_39379,N_38626);
or U41358 (N_41358,N_38488,N_38224);
nor U41359 (N_41359,N_39563,N_39068);
nand U41360 (N_41360,N_39962,N_39724);
nand U41361 (N_41361,N_38153,N_38790);
nor U41362 (N_41362,N_38652,N_38976);
nand U41363 (N_41363,N_39344,N_39256);
and U41364 (N_41364,N_38832,N_38369);
and U41365 (N_41365,N_39590,N_39498);
and U41366 (N_41366,N_39614,N_38005);
and U41367 (N_41367,N_38095,N_38975);
nand U41368 (N_41368,N_38377,N_39194);
nand U41369 (N_41369,N_39965,N_38876);
nand U41370 (N_41370,N_38850,N_39465);
or U41371 (N_41371,N_39939,N_39749);
and U41372 (N_41372,N_39925,N_38018);
nor U41373 (N_41373,N_38869,N_38483);
and U41374 (N_41374,N_38911,N_39547);
xor U41375 (N_41375,N_38698,N_38302);
and U41376 (N_41376,N_38652,N_39116);
nand U41377 (N_41377,N_39865,N_39816);
nor U41378 (N_41378,N_39142,N_38318);
or U41379 (N_41379,N_38838,N_39279);
xnor U41380 (N_41380,N_39757,N_39849);
xor U41381 (N_41381,N_39170,N_39265);
nor U41382 (N_41382,N_39467,N_38712);
xor U41383 (N_41383,N_38827,N_38540);
and U41384 (N_41384,N_38618,N_39655);
xnor U41385 (N_41385,N_38151,N_39190);
or U41386 (N_41386,N_39423,N_39205);
xor U41387 (N_41387,N_39438,N_39269);
nand U41388 (N_41388,N_38928,N_39077);
or U41389 (N_41389,N_39333,N_39066);
xnor U41390 (N_41390,N_39595,N_39714);
nor U41391 (N_41391,N_38456,N_38850);
and U41392 (N_41392,N_38325,N_39714);
xnor U41393 (N_41393,N_38685,N_39050);
nor U41394 (N_41394,N_39712,N_39492);
or U41395 (N_41395,N_38670,N_38893);
nor U41396 (N_41396,N_39701,N_38133);
nor U41397 (N_41397,N_38097,N_39717);
or U41398 (N_41398,N_38741,N_38446);
or U41399 (N_41399,N_39179,N_38864);
or U41400 (N_41400,N_38063,N_39233);
or U41401 (N_41401,N_39645,N_38148);
nand U41402 (N_41402,N_38631,N_38589);
nand U41403 (N_41403,N_38789,N_39124);
or U41404 (N_41404,N_39636,N_38923);
nor U41405 (N_41405,N_38192,N_38537);
xnor U41406 (N_41406,N_38442,N_39194);
and U41407 (N_41407,N_39816,N_38590);
xnor U41408 (N_41408,N_38828,N_38455);
and U41409 (N_41409,N_38971,N_39863);
or U41410 (N_41410,N_38855,N_38076);
or U41411 (N_41411,N_39482,N_38433);
and U41412 (N_41412,N_38716,N_38204);
or U41413 (N_41413,N_38493,N_38476);
nand U41414 (N_41414,N_39450,N_38646);
or U41415 (N_41415,N_39450,N_39380);
nand U41416 (N_41416,N_38125,N_39027);
nand U41417 (N_41417,N_38388,N_38302);
nand U41418 (N_41418,N_39716,N_38485);
or U41419 (N_41419,N_38925,N_38936);
nor U41420 (N_41420,N_39528,N_39860);
xor U41421 (N_41421,N_38298,N_39498);
nor U41422 (N_41422,N_39551,N_39469);
xor U41423 (N_41423,N_39179,N_38590);
and U41424 (N_41424,N_38690,N_39483);
nand U41425 (N_41425,N_39432,N_38309);
nand U41426 (N_41426,N_39993,N_39040);
xnor U41427 (N_41427,N_38763,N_38331);
xnor U41428 (N_41428,N_39435,N_38936);
nor U41429 (N_41429,N_39293,N_38513);
and U41430 (N_41430,N_39969,N_39698);
and U41431 (N_41431,N_38606,N_39872);
nor U41432 (N_41432,N_39669,N_38463);
nand U41433 (N_41433,N_38723,N_38953);
or U41434 (N_41434,N_39603,N_38217);
or U41435 (N_41435,N_39759,N_39112);
nand U41436 (N_41436,N_38536,N_39402);
nor U41437 (N_41437,N_38936,N_38883);
nor U41438 (N_41438,N_39453,N_39880);
nor U41439 (N_41439,N_38408,N_38232);
nor U41440 (N_41440,N_39125,N_39733);
nand U41441 (N_41441,N_38178,N_39901);
xnor U41442 (N_41442,N_38742,N_39375);
and U41443 (N_41443,N_39660,N_39206);
nand U41444 (N_41444,N_39847,N_39909);
or U41445 (N_41445,N_38575,N_38920);
or U41446 (N_41446,N_39149,N_38865);
or U41447 (N_41447,N_38647,N_39009);
nand U41448 (N_41448,N_38834,N_38480);
nor U41449 (N_41449,N_38915,N_38965);
xor U41450 (N_41450,N_38436,N_38335);
nor U41451 (N_41451,N_39235,N_38082);
nor U41452 (N_41452,N_39348,N_38887);
xor U41453 (N_41453,N_39016,N_38604);
and U41454 (N_41454,N_39588,N_38101);
or U41455 (N_41455,N_38169,N_39783);
xnor U41456 (N_41456,N_38411,N_38978);
and U41457 (N_41457,N_39696,N_39495);
nor U41458 (N_41458,N_38947,N_38813);
xor U41459 (N_41459,N_39117,N_38966);
nand U41460 (N_41460,N_39375,N_38207);
xnor U41461 (N_41461,N_39275,N_39535);
nand U41462 (N_41462,N_39071,N_38839);
nor U41463 (N_41463,N_39416,N_38792);
xor U41464 (N_41464,N_38915,N_39758);
and U41465 (N_41465,N_38140,N_39894);
nor U41466 (N_41466,N_39342,N_38118);
or U41467 (N_41467,N_38442,N_38433);
nand U41468 (N_41468,N_38492,N_39189);
xor U41469 (N_41469,N_38118,N_38312);
nand U41470 (N_41470,N_39349,N_39734);
nor U41471 (N_41471,N_38892,N_38290);
or U41472 (N_41472,N_38793,N_38061);
and U41473 (N_41473,N_38388,N_38186);
nor U41474 (N_41474,N_38252,N_39724);
nand U41475 (N_41475,N_39925,N_38358);
nor U41476 (N_41476,N_38745,N_38321);
xnor U41477 (N_41477,N_39241,N_39608);
nand U41478 (N_41478,N_39586,N_39540);
nor U41479 (N_41479,N_39133,N_38174);
and U41480 (N_41480,N_38351,N_38329);
nor U41481 (N_41481,N_38414,N_38781);
nand U41482 (N_41482,N_39327,N_38755);
nand U41483 (N_41483,N_38122,N_39046);
or U41484 (N_41484,N_39836,N_39318);
xnor U41485 (N_41485,N_38149,N_38817);
nor U41486 (N_41486,N_38461,N_38590);
or U41487 (N_41487,N_39084,N_38852);
and U41488 (N_41488,N_38252,N_39782);
nor U41489 (N_41489,N_39302,N_39386);
xnor U41490 (N_41490,N_39275,N_39801);
xnor U41491 (N_41491,N_38402,N_39334);
xnor U41492 (N_41492,N_38003,N_39931);
xor U41493 (N_41493,N_38180,N_39282);
nor U41494 (N_41494,N_38811,N_39046);
nand U41495 (N_41495,N_38149,N_38477);
and U41496 (N_41496,N_39787,N_38053);
nor U41497 (N_41497,N_39693,N_39114);
nor U41498 (N_41498,N_39331,N_39790);
xnor U41499 (N_41499,N_38155,N_38758);
and U41500 (N_41500,N_39479,N_38671);
and U41501 (N_41501,N_38008,N_38841);
xor U41502 (N_41502,N_39318,N_39326);
xor U41503 (N_41503,N_38576,N_39494);
nand U41504 (N_41504,N_38837,N_39737);
nor U41505 (N_41505,N_38377,N_38446);
and U41506 (N_41506,N_39430,N_39455);
xor U41507 (N_41507,N_39946,N_38179);
xor U41508 (N_41508,N_38953,N_39219);
nand U41509 (N_41509,N_39178,N_38089);
nor U41510 (N_41510,N_39499,N_39683);
xnor U41511 (N_41511,N_39093,N_39074);
nor U41512 (N_41512,N_38357,N_39212);
nand U41513 (N_41513,N_38562,N_38870);
or U41514 (N_41514,N_39639,N_38416);
or U41515 (N_41515,N_38185,N_38765);
and U41516 (N_41516,N_38461,N_39151);
nor U41517 (N_41517,N_38832,N_38167);
nand U41518 (N_41518,N_38282,N_38686);
xnor U41519 (N_41519,N_38814,N_38002);
xnor U41520 (N_41520,N_39914,N_38619);
nor U41521 (N_41521,N_39758,N_38712);
nor U41522 (N_41522,N_38186,N_39067);
or U41523 (N_41523,N_38031,N_38916);
xnor U41524 (N_41524,N_39400,N_39132);
xor U41525 (N_41525,N_38986,N_38838);
nand U41526 (N_41526,N_38988,N_39595);
nand U41527 (N_41527,N_38903,N_39963);
nor U41528 (N_41528,N_39383,N_39998);
xor U41529 (N_41529,N_38803,N_39481);
or U41530 (N_41530,N_39421,N_39550);
or U41531 (N_41531,N_39207,N_39491);
or U41532 (N_41532,N_38897,N_38606);
nand U41533 (N_41533,N_39907,N_39111);
nand U41534 (N_41534,N_38738,N_39894);
nor U41535 (N_41535,N_38755,N_39104);
nor U41536 (N_41536,N_38451,N_39388);
and U41537 (N_41537,N_39224,N_39144);
or U41538 (N_41538,N_39347,N_39633);
and U41539 (N_41539,N_38544,N_39966);
xnor U41540 (N_41540,N_38137,N_39259);
nor U41541 (N_41541,N_38806,N_38704);
nand U41542 (N_41542,N_38106,N_38107);
nand U41543 (N_41543,N_39452,N_38381);
nor U41544 (N_41544,N_39020,N_38587);
or U41545 (N_41545,N_39243,N_39792);
nand U41546 (N_41546,N_39934,N_38431);
or U41547 (N_41547,N_39763,N_38860);
nand U41548 (N_41548,N_39040,N_38840);
or U41549 (N_41549,N_38267,N_38369);
xor U41550 (N_41550,N_39639,N_39737);
nor U41551 (N_41551,N_38106,N_38667);
or U41552 (N_41552,N_38530,N_39233);
xor U41553 (N_41553,N_38831,N_38590);
xor U41554 (N_41554,N_38927,N_38892);
or U41555 (N_41555,N_39483,N_38226);
nand U41556 (N_41556,N_38858,N_39389);
xnor U41557 (N_41557,N_38369,N_38363);
or U41558 (N_41558,N_39622,N_39652);
and U41559 (N_41559,N_39576,N_38562);
xnor U41560 (N_41560,N_39624,N_39287);
nand U41561 (N_41561,N_39611,N_39970);
nand U41562 (N_41562,N_38453,N_38097);
and U41563 (N_41563,N_38808,N_39908);
nor U41564 (N_41564,N_38381,N_39696);
and U41565 (N_41565,N_39659,N_39178);
xnor U41566 (N_41566,N_39696,N_38683);
and U41567 (N_41567,N_38776,N_38400);
or U41568 (N_41568,N_38169,N_38892);
nand U41569 (N_41569,N_38248,N_38361);
nor U41570 (N_41570,N_39329,N_38762);
or U41571 (N_41571,N_38958,N_39984);
nand U41572 (N_41572,N_39025,N_39510);
and U41573 (N_41573,N_38291,N_39920);
nand U41574 (N_41574,N_38293,N_39481);
or U41575 (N_41575,N_38713,N_39213);
nor U41576 (N_41576,N_39201,N_38620);
nand U41577 (N_41577,N_39153,N_38979);
nor U41578 (N_41578,N_38393,N_39643);
or U41579 (N_41579,N_38389,N_39916);
nand U41580 (N_41580,N_38554,N_39390);
nand U41581 (N_41581,N_39400,N_39342);
and U41582 (N_41582,N_39618,N_39039);
nand U41583 (N_41583,N_39360,N_38165);
xnor U41584 (N_41584,N_38142,N_38446);
and U41585 (N_41585,N_39497,N_38023);
or U41586 (N_41586,N_39548,N_39206);
nor U41587 (N_41587,N_39348,N_39250);
or U41588 (N_41588,N_39616,N_38739);
nor U41589 (N_41589,N_39799,N_39604);
nand U41590 (N_41590,N_39585,N_39768);
or U41591 (N_41591,N_38679,N_38426);
xnor U41592 (N_41592,N_39853,N_38870);
xor U41593 (N_41593,N_38330,N_38759);
nand U41594 (N_41594,N_38491,N_38247);
xnor U41595 (N_41595,N_39825,N_38895);
nand U41596 (N_41596,N_39670,N_38765);
nor U41597 (N_41597,N_39277,N_39013);
and U41598 (N_41598,N_39439,N_38231);
and U41599 (N_41599,N_38443,N_38618);
and U41600 (N_41600,N_38560,N_39809);
or U41601 (N_41601,N_39526,N_39673);
or U41602 (N_41602,N_38024,N_39465);
nand U41603 (N_41603,N_39993,N_38791);
nor U41604 (N_41604,N_38421,N_38736);
xor U41605 (N_41605,N_38402,N_38993);
nor U41606 (N_41606,N_39965,N_38007);
nor U41607 (N_41607,N_39539,N_39734);
nand U41608 (N_41608,N_39067,N_39608);
nand U41609 (N_41609,N_38779,N_39837);
nand U41610 (N_41610,N_39726,N_39942);
nor U41611 (N_41611,N_39909,N_38032);
nor U41612 (N_41612,N_39978,N_38454);
or U41613 (N_41613,N_38829,N_38431);
nor U41614 (N_41614,N_39237,N_38421);
and U41615 (N_41615,N_39586,N_39866);
xor U41616 (N_41616,N_39687,N_38532);
or U41617 (N_41617,N_38988,N_39765);
or U41618 (N_41618,N_38626,N_38131);
nor U41619 (N_41619,N_38808,N_38662);
and U41620 (N_41620,N_39782,N_39919);
xor U41621 (N_41621,N_38049,N_38253);
or U41622 (N_41622,N_39443,N_39648);
nand U41623 (N_41623,N_39518,N_39085);
or U41624 (N_41624,N_38975,N_38568);
and U41625 (N_41625,N_38318,N_39712);
nor U41626 (N_41626,N_38961,N_39874);
and U41627 (N_41627,N_38779,N_38769);
and U41628 (N_41628,N_39707,N_38097);
or U41629 (N_41629,N_38212,N_39665);
and U41630 (N_41630,N_38120,N_39221);
nor U41631 (N_41631,N_38975,N_39517);
nor U41632 (N_41632,N_39829,N_38176);
or U41633 (N_41633,N_38325,N_38473);
or U41634 (N_41634,N_38522,N_38551);
nand U41635 (N_41635,N_39516,N_38143);
nor U41636 (N_41636,N_39433,N_38269);
and U41637 (N_41637,N_38807,N_38068);
nor U41638 (N_41638,N_38828,N_38986);
nor U41639 (N_41639,N_38297,N_39688);
xnor U41640 (N_41640,N_38184,N_38384);
nor U41641 (N_41641,N_38680,N_38099);
nand U41642 (N_41642,N_38664,N_39005);
or U41643 (N_41643,N_39957,N_39056);
nand U41644 (N_41644,N_38858,N_38748);
and U41645 (N_41645,N_38607,N_39653);
nand U41646 (N_41646,N_38656,N_38818);
or U41647 (N_41647,N_39551,N_38582);
nor U41648 (N_41648,N_38899,N_39258);
nor U41649 (N_41649,N_39873,N_38507);
nand U41650 (N_41650,N_39688,N_38915);
and U41651 (N_41651,N_39884,N_38152);
nand U41652 (N_41652,N_39115,N_39665);
xor U41653 (N_41653,N_39550,N_38380);
or U41654 (N_41654,N_38848,N_38819);
and U41655 (N_41655,N_38638,N_38403);
and U41656 (N_41656,N_39770,N_38558);
nor U41657 (N_41657,N_39365,N_39246);
or U41658 (N_41658,N_39913,N_39213);
or U41659 (N_41659,N_39690,N_39300);
or U41660 (N_41660,N_39498,N_39633);
nor U41661 (N_41661,N_39781,N_38912);
nor U41662 (N_41662,N_38790,N_38044);
xnor U41663 (N_41663,N_38851,N_39351);
and U41664 (N_41664,N_39275,N_38770);
and U41665 (N_41665,N_39760,N_38655);
nor U41666 (N_41666,N_38059,N_38217);
or U41667 (N_41667,N_39184,N_39632);
and U41668 (N_41668,N_39107,N_38519);
or U41669 (N_41669,N_39740,N_39822);
or U41670 (N_41670,N_39818,N_38414);
nor U41671 (N_41671,N_39976,N_38406);
nand U41672 (N_41672,N_38644,N_39637);
xor U41673 (N_41673,N_39622,N_39718);
xor U41674 (N_41674,N_38966,N_39778);
nor U41675 (N_41675,N_39322,N_38694);
nand U41676 (N_41676,N_38681,N_38665);
nand U41677 (N_41677,N_38657,N_38565);
or U41678 (N_41678,N_39449,N_38415);
nor U41679 (N_41679,N_39350,N_38534);
nand U41680 (N_41680,N_38536,N_38241);
nand U41681 (N_41681,N_38620,N_39519);
or U41682 (N_41682,N_38730,N_39750);
xor U41683 (N_41683,N_39245,N_39258);
or U41684 (N_41684,N_38964,N_38180);
nor U41685 (N_41685,N_39508,N_38854);
nor U41686 (N_41686,N_39196,N_38662);
nor U41687 (N_41687,N_39322,N_38442);
and U41688 (N_41688,N_38785,N_39715);
nor U41689 (N_41689,N_38961,N_39276);
and U41690 (N_41690,N_39212,N_38187);
nand U41691 (N_41691,N_38063,N_39778);
xor U41692 (N_41692,N_39178,N_38680);
xor U41693 (N_41693,N_38310,N_38515);
nor U41694 (N_41694,N_39905,N_38985);
or U41695 (N_41695,N_39470,N_38166);
xnor U41696 (N_41696,N_39118,N_39896);
nand U41697 (N_41697,N_39769,N_38368);
and U41698 (N_41698,N_38794,N_38087);
xnor U41699 (N_41699,N_38628,N_38933);
nor U41700 (N_41700,N_38309,N_38185);
or U41701 (N_41701,N_39420,N_38708);
or U41702 (N_41702,N_38866,N_39084);
nand U41703 (N_41703,N_39891,N_38698);
nand U41704 (N_41704,N_38559,N_38742);
and U41705 (N_41705,N_39898,N_39194);
or U41706 (N_41706,N_39148,N_39035);
xor U41707 (N_41707,N_38822,N_39161);
nand U41708 (N_41708,N_39686,N_38229);
xor U41709 (N_41709,N_39074,N_39748);
or U41710 (N_41710,N_38125,N_39641);
or U41711 (N_41711,N_38983,N_39127);
or U41712 (N_41712,N_39673,N_39741);
or U41713 (N_41713,N_39730,N_39856);
nand U41714 (N_41714,N_39409,N_39468);
nor U41715 (N_41715,N_38162,N_39693);
nor U41716 (N_41716,N_39526,N_38688);
or U41717 (N_41717,N_38876,N_39181);
nand U41718 (N_41718,N_39240,N_38883);
nor U41719 (N_41719,N_39372,N_38064);
or U41720 (N_41720,N_38109,N_38560);
and U41721 (N_41721,N_38158,N_38115);
and U41722 (N_41722,N_38158,N_38617);
and U41723 (N_41723,N_38536,N_38103);
nor U41724 (N_41724,N_38093,N_38662);
nand U41725 (N_41725,N_38253,N_39766);
and U41726 (N_41726,N_39906,N_39099);
nor U41727 (N_41727,N_39211,N_39132);
nand U41728 (N_41728,N_39621,N_38497);
nand U41729 (N_41729,N_38010,N_39888);
or U41730 (N_41730,N_38030,N_39782);
or U41731 (N_41731,N_38873,N_38760);
and U41732 (N_41732,N_39208,N_39727);
nor U41733 (N_41733,N_38715,N_38693);
or U41734 (N_41734,N_38493,N_39572);
or U41735 (N_41735,N_38628,N_38661);
nand U41736 (N_41736,N_39150,N_38578);
or U41737 (N_41737,N_38241,N_38430);
or U41738 (N_41738,N_38356,N_38315);
xor U41739 (N_41739,N_39488,N_39602);
xnor U41740 (N_41740,N_38863,N_38220);
or U41741 (N_41741,N_39522,N_38370);
nor U41742 (N_41742,N_38914,N_39137);
nor U41743 (N_41743,N_39000,N_39845);
or U41744 (N_41744,N_39680,N_38776);
nor U41745 (N_41745,N_39682,N_39418);
xnor U41746 (N_41746,N_39525,N_38501);
nand U41747 (N_41747,N_39865,N_39500);
nand U41748 (N_41748,N_38648,N_39470);
and U41749 (N_41749,N_39685,N_38143);
and U41750 (N_41750,N_39417,N_39950);
and U41751 (N_41751,N_39020,N_38120);
xor U41752 (N_41752,N_38100,N_39456);
and U41753 (N_41753,N_39489,N_39875);
or U41754 (N_41754,N_39929,N_39042);
and U41755 (N_41755,N_38835,N_38321);
or U41756 (N_41756,N_39213,N_38520);
or U41757 (N_41757,N_38075,N_38993);
xor U41758 (N_41758,N_39402,N_38468);
xnor U41759 (N_41759,N_38932,N_39321);
or U41760 (N_41760,N_38176,N_38624);
nor U41761 (N_41761,N_39162,N_39867);
nor U41762 (N_41762,N_39866,N_38008);
xor U41763 (N_41763,N_39172,N_39531);
and U41764 (N_41764,N_38830,N_38070);
nor U41765 (N_41765,N_38033,N_38658);
nand U41766 (N_41766,N_38076,N_38356);
nor U41767 (N_41767,N_39572,N_39919);
and U41768 (N_41768,N_38498,N_38969);
and U41769 (N_41769,N_39809,N_38123);
and U41770 (N_41770,N_38807,N_39586);
or U41771 (N_41771,N_38502,N_38340);
or U41772 (N_41772,N_38844,N_38075);
or U41773 (N_41773,N_39867,N_38057);
nand U41774 (N_41774,N_38583,N_38766);
nor U41775 (N_41775,N_38252,N_39627);
nor U41776 (N_41776,N_39520,N_38875);
xnor U41777 (N_41777,N_39383,N_38859);
nor U41778 (N_41778,N_38247,N_38386);
xor U41779 (N_41779,N_38659,N_39653);
and U41780 (N_41780,N_39601,N_38994);
nand U41781 (N_41781,N_38247,N_38156);
nand U41782 (N_41782,N_38370,N_38083);
nand U41783 (N_41783,N_38287,N_38525);
nand U41784 (N_41784,N_39792,N_39245);
nand U41785 (N_41785,N_38265,N_39801);
nor U41786 (N_41786,N_39941,N_39202);
xnor U41787 (N_41787,N_39574,N_39031);
and U41788 (N_41788,N_38650,N_39665);
or U41789 (N_41789,N_39466,N_38055);
or U41790 (N_41790,N_39950,N_39598);
or U41791 (N_41791,N_38797,N_38439);
or U41792 (N_41792,N_39244,N_38451);
nor U41793 (N_41793,N_38484,N_39274);
or U41794 (N_41794,N_38242,N_39886);
xnor U41795 (N_41795,N_39511,N_38779);
nand U41796 (N_41796,N_38676,N_39114);
nand U41797 (N_41797,N_38255,N_39615);
nor U41798 (N_41798,N_39865,N_39697);
and U41799 (N_41799,N_38350,N_38299);
nor U41800 (N_41800,N_39043,N_39668);
xor U41801 (N_41801,N_39522,N_39194);
nand U41802 (N_41802,N_38609,N_38373);
nor U41803 (N_41803,N_38602,N_38568);
and U41804 (N_41804,N_38817,N_39028);
or U41805 (N_41805,N_38639,N_39714);
and U41806 (N_41806,N_38259,N_39873);
or U41807 (N_41807,N_39534,N_39361);
and U41808 (N_41808,N_38524,N_38787);
or U41809 (N_41809,N_39381,N_38204);
nand U41810 (N_41810,N_39607,N_39928);
xor U41811 (N_41811,N_39468,N_38164);
xnor U41812 (N_41812,N_39516,N_38053);
xnor U41813 (N_41813,N_39586,N_38677);
or U41814 (N_41814,N_38172,N_39880);
nand U41815 (N_41815,N_38953,N_38176);
xor U41816 (N_41816,N_38410,N_39004);
nor U41817 (N_41817,N_39602,N_39766);
xor U41818 (N_41818,N_38592,N_39512);
nand U41819 (N_41819,N_38891,N_39582);
and U41820 (N_41820,N_38780,N_39074);
nand U41821 (N_41821,N_38150,N_39179);
and U41822 (N_41822,N_39825,N_39480);
or U41823 (N_41823,N_39193,N_39385);
and U41824 (N_41824,N_39387,N_39227);
and U41825 (N_41825,N_39476,N_39226);
and U41826 (N_41826,N_38786,N_39322);
nor U41827 (N_41827,N_38263,N_38892);
and U41828 (N_41828,N_38097,N_39744);
xor U41829 (N_41829,N_38329,N_38804);
xnor U41830 (N_41830,N_38766,N_38005);
nand U41831 (N_41831,N_38011,N_38669);
and U41832 (N_41832,N_38289,N_39049);
nor U41833 (N_41833,N_39847,N_39964);
xor U41834 (N_41834,N_39245,N_38790);
nand U41835 (N_41835,N_38602,N_39947);
nand U41836 (N_41836,N_38380,N_39188);
and U41837 (N_41837,N_39371,N_39904);
nor U41838 (N_41838,N_38484,N_39813);
and U41839 (N_41839,N_39471,N_38319);
xor U41840 (N_41840,N_38595,N_38478);
and U41841 (N_41841,N_39108,N_39299);
nor U41842 (N_41842,N_39525,N_38978);
nand U41843 (N_41843,N_39456,N_38807);
and U41844 (N_41844,N_39242,N_38390);
nor U41845 (N_41845,N_38519,N_38682);
nor U41846 (N_41846,N_38803,N_38162);
xor U41847 (N_41847,N_39236,N_39749);
and U41848 (N_41848,N_39252,N_39499);
nor U41849 (N_41849,N_38547,N_38849);
and U41850 (N_41850,N_38037,N_39165);
nand U41851 (N_41851,N_38930,N_39314);
and U41852 (N_41852,N_39555,N_38456);
and U41853 (N_41853,N_39305,N_38244);
or U41854 (N_41854,N_39484,N_39105);
and U41855 (N_41855,N_39212,N_38035);
or U41856 (N_41856,N_39539,N_39613);
xnor U41857 (N_41857,N_39476,N_38713);
or U41858 (N_41858,N_38504,N_39021);
nor U41859 (N_41859,N_39873,N_38566);
and U41860 (N_41860,N_39598,N_39792);
nor U41861 (N_41861,N_39320,N_38049);
or U41862 (N_41862,N_38978,N_39238);
and U41863 (N_41863,N_38393,N_38958);
and U41864 (N_41864,N_38810,N_38386);
nor U41865 (N_41865,N_38414,N_39983);
or U41866 (N_41866,N_38193,N_38135);
xor U41867 (N_41867,N_39180,N_38348);
or U41868 (N_41868,N_39435,N_39047);
and U41869 (N_41869,N_39747,N_38378);
or U41870 (N_41870,N_39314,N_38740);
xnor U41871 (N_41871,N_38697,N_38605);
xor U41872 (N_41872,N_38064,N_38571);
or U41873 (N_41873,N_39482,N_39190);
nand U41874 (N_41874,N_38879,N_39856);
and U41875 (N_41875,N_38867,N_39916);
or U41876 (N_41876,N_38412,N_38433);
nor U41877 (N_41877,N_38787,N_39184);
nand U41878 (N_41878,N_39634,N_39262);
nor U41879 (N_41879,N_39109,N_39150);
or U41880 (N_41880,N_39303,N_38758);
or U41881 (N_41881,N_38557,N_39225);
or U41882 (N_41882,N_38656,N_38621);
xnor U41883 (N_41883,N_38132,N_39503);
nand U41884 (N_41884,N_38030,N_39511);
nand U41885 (N_41885,N_39133,N_38293);
and U41886 (N_41886,N_38852,N_39168);
or U41887 (N_41887,N_39318,N_39331);
nand U41888 (N_41888,N_39613,N_39040);
or U41889 (N_41889,N_38181,N_39958);
nand U41890 (N_41890,N_39549,N_39717);
nand U41891 (N_41891,N_39597,N_38390);
or U41892 (N_41892,N_39070,N_39002);
xnor U41893 (N_41893,N_38989,N_38605);
nor U41894 (N_41894,N_38678,N_39859);
and U41895 (N_41895,N_38487,N_39934);
xor U41896 (N_41896,N_39987,N_39745);
and U41897 (N_41897,N_39337,N_39284);
or U41898 (N_41898,N_39741,N_39627);
nand U41899 (N_41899,N_39880,N_38217);
xor U41900 (N_41900,N_39405,N_39415);
and U41901 (N_41901,N_38908,N_38100);
and U41902 (N_41902,N_38670,N_39315);
nand U41903 (N_41903,N_38981,N_39252);
or U41904 (N_41904,N_39334,N_38541);
xnor U41905 (N_41905,N_38879,N_38698);
nand U41906 (N_41906,N_38536,N_38683);
or U41907 (N_41907,N_39981,N_39269);
and U41908 (N_41908,N_38106,N_38218);
xnor U41909 (N_41909,N_38396,N_38504);
xor U41910 (N_41910,N_39053,N_38625);
and U41911 (N_41911,N_39911,N_38117);
and U41912 (N_41912,N_38262,N_38490);
nor U41913 (N_41913,N_38726,N_39439);
xor U41914 (N_41914,N_38025,N_38192);
nand U41915 (N_41915,N_39832,N_38929);
and U41916 (N_41916,N_39924,N_38905);
nand U41917 (N_41917,N_38029,N_39703);
nand U41918 (N_41918,N_39077,N_38486);
and U41919 (N_41919,N_39513,N_39227);
nor U41920 (N_41920,N_39333,N_39447);
nand U41921 (N_41921,N_38861,N_38924);
xor U41922 (N_41922,N_39271,N_38588);
xor U41923 (N_41923,N_38069,N_38448);
xnor U41924 (N_41924,N_39598,N_38604);
nor U41925 (N_41925,N_39873,N_39505);
nor U41926 (N_41926,N_39554,N_38369);
or U41927 (N_41927,N_38354,N_39853);
and U41928 (N_41928,N_39330,N_38937);
nor U41929 (N_41929,N_38359,N_39058);
and U41930 (N_41930,N_38973,N_38157);
xnor U41931 (N_41931,N_38951,N_38426);
nand U41932 (N_41932,N_38867,N_39056);
xnor U41933 (N_41933,N_39390,N_39414);
or U41934 (N_41934,N_39000,N_39762);
and U41935 (N_41935,N_38336,N_39865);
and U41936 (N_41936,N_38126,N_38794);
or U41937 (N_41937,N_39714,N_39958);
nand U41938 (N_41938,N_38104,N_38950);
xnor U41939 (N_41939,N_39145,N_38258);
nor U41940 (N_41940,N_39389,N_39894);
and U41941 (N_41941,N_39218,N_38746);
xnor U41942 (N_41942,N_38825,N_38497);
and U41943 (N_41943,N_39974,N_38116);
nor U41944 (N_41944,N_38097,N_39044);
xor U41945 (N_41945,N_39622,N_38313);
and U41946 (N_41946,N_38365,N_39844);
and U41947 (N_41947,N_39915,N_39490);
or U41948 (N_41948,N_39633,N_38987);
and U41949 (N_41949,N_38660,N_38400);
nor U41950 (N_41950,N_39450,N_38033);
nand U41951 (N_41951,N_38262,N_39441);
nor U41952 (N_41952,N_39501,N_38314);
xor U41953 (N_41953,N_38768,N_39132);
or U41954 (N_41954,N_39530,N_39810);
or U41955 (N_41955,N_39844,N_39083);
nand U41956 (N_41956,N_38974,N_38079);
xnor U41957 (N_41957,N_39587,N_38049);
nor U41958 (N_41958,N_39749,N_39183);
and U41959 (N_41959,N_38745,N_38498);
or U41960 (N_41960,N_39520,N_39574);
nand U41961 (N_41961,N_38919,N_39556);
nand U41962 (N_41962,N_39524,N_38944);
nor U41963 (N_41963,N_39469,N_38443);
and U41964 (N_41964,N_38667,N_38494);
and U41965 (N_41965,N_39290,N_38023);
nand U41966 (N_41966,N_39921,N_39194);
xor U41967 (N_41967,N_39696,N_39860);
nand U41968 (N_41968,N_39311,N_39228);
and U41969 (N_41969,N_39684,N_38099);
xnor U41970 (N_41970,N_38185,N_38313);
nand U41971 (N_41971,N_38192,N_38198);
xor U41972 (N_41972,N_38834,N_38639);
xor U41973 (N_41973,N_39189,N_39587);
nand U41974 (N_41974,N_39262,N_38502);
or U41975 (N_41975,N_39168,N_38607);
xor U41976 (N_41976,N_39856,N_38025);
xor U41977 (N_41977,N_38881,N_38096);
nand U41978 (N_41978,N_39108,N_38360);
and U41979 (N_41979,N_39858,N_39683);
nand U41980 (N_41980,N_38365,N_39137);
nor U41981 (N_41981,N_38932,N_39984);
nand U41982 (N_41982,N_39647,N_39278);
nand U41983 (N_41983,N_38260,N_39366);
xor U41984 (N_41984,N_38787,N_38954);
and U41985 (N_41985,N_39566,N_39601);
nand U41986 (N_41986,N_39810,N_38638);
nor U41987 (N_41987,N_38047,N_39372);
and U41988 (N_41988,N_38730,N_39876);
nor U41989 (N_41989,N_39308,N_38595);
xnor U41990 (N_41990,N_39277,N_39423);
xnor U41991 (N_41991,N_39858,N_39497);
and U41992 (N_41992,N_39416,N_39835);
xnor U41993 (N_41993,N_39329,N_38658);
xor U41994 (N_41994,N_39947,N_38125);
nand U41995 (N_41995,N_39283,N_38453);
nor U41996 (N_41996,N_38120,N_39134);
nor U41997 (N_41997,N_39775,N_38002);
nand U41998 (N_41998,N_39153,N_39121);
or U41999 (N_41999,N_39230,N_38100);
nand U42000 (N_42000,N_40999,N_41967);
xnor U42001 (N_42001,N_41301,N_41884);
and U42002 (N_42002,N_40537,N_41325);
and U42003 (N_42003,N_40680,N_40446);
nand U42004 (N_42004,N_41579,N_40890);
and U42005 (N_42005,N_40551,N_40158);
nand U42006 (N_42006,N_41187,N_41762);
nor U42007 (N_42007,N_40529,N_41974);
xnor U42008 (N_42008,N_40755,N_40809);
nor U42009 (N_42009,N_41130,N_41870);
or U42010 (N_42010,N_41033,N_41944);
nor U42011 (N_42011,N_40093,N_40946);
and U42012 (N_42012,N_40577,N_40459);
nand U42013 (N_42013,N_40117,N_41175);
and U42014 (N_42014,N_41633,N_41165);
nand U42015 (N_42015,N_41132,N_41802);
nor U42016 (N_42016,N_40321,N_40985);
nor U42017 (N_42017,N_40535,N_41695);
nor U42018 (N_42018,N_41184,N_41515);
xor U42019 (N_42019,N_41010,N_40236);
or U42020 (N_42020,N_40269,N_40258);
or U42021 (N_42021,N_41101,N_40700);
nand U42022 (N_42022,N_40880,N_41277);
nor U42023 (N_42023,N_40043,N_41985);
or U42024 (N_42024,N_41908,N_40637);
nand U42025 (N_42025,N_40540,N_40346);
xnor U42026 (N_42026,N_40007,N_41648);
xor U42027 (N_42027,N_40076,N_40353);
and U42028 (N_42028,N_40653,N_40203);
nor U42029 (N_42029,N_41414,N_41264);
nand U42030 (N_42030,N_40275,N_41440);
nand U42031 (N_42031,N_40285,N_41980);
or U42032 (N_42032,N_40591,N_40307);
nand U42033 (N_42033,N_41972,N_41361);
nor U42034 (N_42034,N_40197,N_40479);
or U42035 (N_42035,N_41774,N_41464);
nand U42036 (N_42036,N_41926,N_40761);
nand U42037 (N_42037,N_40658,N_40305);
nor U42038 (N_42038,N_40705,N_41917);
and U42039 (N_42039,N_40463,N_41534);
nand U42040 (N_42040,N_40092,N_40026);
nor U42041 (N_42041,N_41211,N_40378);
nand U42042 (N_42042,N_41072,N_40478);
and U42043 (N_42043,N_40775,N_41900);
nand U42044 (N_42044,N_40186,N_41653);
or U42045 (N_42045,N_40221,N_41268);
nor U42046 (N_42046,N_41871,N_41588);
and U42047 (N_42047,N_40679,N_41895);
nor U42048 (N_42048,N_41749,N_40831);
nor U42049 (N_42049,N_40640,N_41109);
xor U42050 (N_42050,N_41161,N_40748);
and U42051 (N_42051,N_40993,N_41842);
nand U42052 (N_42052,N_41990,N_41496);
nand U42053 (N_42053,N_40575,N_40785);
xnor U42054 (N_42054,N_41129,N_41643);
nand U42055 (N_42055,N_41903,N_41634);
nand U42056 (N_42056,N_41032,N_40832);
and U42057 (N_42057,N_41910,N_41083);
xor U42058 (N_42058,N_41878,N_41997);
xnor U42059 (N_42059,N_40528,N_41351);
xor U42060 (N_42060,N_41355,N_40808);
and U42061 (N_42061,N_40308,N_40019);
nor U42062 (N_42062,N_40558,N_40143);
nor U42063 (N_42063,N_41396,N_41710);
xnor U42064 (N_42064,N_40797,N_41216);
or U42065 (N_42065,N_40228,N_40233);
nand U42066 (N_42066,N_41332,N_40161);
xnor U42067 (N_42067,N_41035,N_40933);
xnor U42068 (N_42068,N_40202,N_40854);
or U42069 (N_42069,N_41862,N_40014);
xor U42070 (N_42070,N_41584,N_41891);
or U42071 (N_42071,N_41416,N_41454);
nor U42072 (N_42072,N_41673,N_40681);
nor U42073 (N_42073,N_40187,N_40821);
nand U42074 (N_42074,N_41546,N_40904);
and U42075 (N_42075,N_40834,N_41307);
nand U42076 (N_42076,N_40249,N_40441);
or U42077 (N_42077,N_41100,N_41973);
xor U42078 (N_42078,N_41274,N_41754);
and U42079 (N_42079,N_40507,N_40215);
nor U42080 (N_42080,N_41732,N_40099);
nand U42081 (N_42081,N_41838,N_40235);
nor U42082 (N_42082,N_40656,N_40648);
nor U42083 (N_42083,N_41806,N_41205);
and U42084 (N_42084,N_41867,N_40815);
and U42085 (N_42085,N_41408,N_41093);
nor U42086 (N_42086,N_41920,N_40980);
or U42087 (N_42087,N_40853,N_41568);
or U42088 (N_42088,N_41436,N_41906);
xnor U42089 (N_42089,N_41660,N_41026);
nor U42090 (N_42090,N_41577,N_41209);
nand U42091 (N_42091,N_40623,N_41131);
and U42092 (N_42092,N_41106,N_41280);
xnor U42093 (N_42093,N_40747,N_41882);
and U42094 (N_42094,N_40484,N_41137);
xnor U42095 (N_42095,N_41552,N_40082);
nor U42096 (N_42096,N_40098,N_41113);
nand U42097 (N_42097,N_40363,N_41993);
nor U42098 (N_42098,N_40872,N_41497);
nand U42099 (N_42099,N_40435,N_40807);
or U42100 (N_42100,N_41984,N_40886);
or U42101 (N_42101,N_41225,N_41108);
xnor U42102 (N_42102,N_40572,N_41748);
or U42103 (N_42103,N_40131,N_41699);
xor U42104 (N_42104,N_41037,N_40817);
nand U42105 (N_42105,N_41146,N_40505);
and U42106 (N_42106,N_41659,N_40369);
nand U42107 (N_42107,N_41369,N_41321);
xnor U42108 (N_42108,N_41279,N_41423);
or U42109 (N_42109,N_41265,N_40184);
xor U42110 (N_42110,N_41843,N_41350);
nor U42111 (N_42111,N_40749,N_41684);
or U42112 (N_42112,N_41599,N_40111);
or U42113 (N_42113,N_41581,N_41485);
nand U42114 (N_42114,N_40960,N_41319);
xor U42115 (N_42115,N_40472,N_41860);
or U42116 (N_42116,N_41704,N_41480);
nand U42117 (N_42117,N_40325,N_40366);
and U42118 (N_42118,N_40642,N_41153);
and U42119 (N_42119,N_40934,N_40181);
or U42120 (N_42120,N_40217,N_40343);
nor U42121 (N_42121,N_40109,N_41305);
nand U42122 (N_42122,N_41442,N_41460);
and U42123 (N_42123,N_40199,N_40911);
nor U42124 (N_42124,N_41134,N_40085);
nor U42125 (N_42125,N_40518,N_40995);
and U42126 (N_42126,N_40284,N_41831);
nand U42127 (N_42127,N_40750,N_41893);
nand U42128 (N_42128,N_41455,N_40768);
nor U42129 (N_42129,N_41326,N_40298);
nor U42130 (N_42130,N_41253,N_41041);
nor U42131 (N_42131,N_40283,N_41387);
nor U42132 (N_42132,N_41038,N_40892);
nor U42133 (N_42133,N_41829,N_40268);
or U42134 (N_42134,N_41742,N_40108);
or U42135 (N_42135,N_41335,N_41705);
nand U42136 (N_42136,N_41328,N_41202);
or U42137 (N_42137,N_41294,N_41885);
xnor U42138 (N_42138,N_41846,N_40708);
nand U42139 (N_42139,N_40138,N_41536);
and U42140 (N_42140,N_40274,N_40135);
nand U42141 (N_42141,N_40465,N_41304);
and U42142 (N_42142,N_40864,N_41786);
xor U42143 (N_42143,N_41345,N_40481);
and U42144 (N_42144,N_40517,N_41323);
nand U42145 (N_42145,N_40922,N_40220);
nand U42146 (N_42146,N_41662,N_41218);
nor U42147 (N_42147,N_41507,N_40859);
or U42148 (N_42148,N_40595,N_40030);
and U42149 (N_42149,N_41942,N_40665);
nor U42150 (N_42150,N_40898,N_40483);
and U42151 (N_42151,N_40494,N_40907);
xnor U42152 (N_42152,N_41687,N_40846);
nand U42153 (N_42153,N_41303,N_41815);
xnor U42154 (N_42154,N_40924,N_41619);
nand U42155 (N_42155,N_40431,N_40418);
or U42156 (N_42156,N_41399,N_40801);
nand U42157 (N_42157,N_40800,N_41804);
nand U42158 (N_42158,N_41276,N_41024);
nand U42159 (N_42159,N_41805,N_40090);
and U42160 (N_42160,N_40185,N_40051);
and U42161 (N_42161,N_41376,N_40234);
or U42162 (N_42162,N_40248,N_40611);
nand U42163 (N_42163,N_41880,N_40614);
nand U42164 (N_42164,N_41835,N_40002);
and U42165 (N_42165,N_41567,N_41943);
nor U42166 (N_42166,N_40627,N_41776);
nand U42167 (N_42167,N_41682,N_41939);
and U42168 (N_42168,N_40089,N_41254);
or U42169 (N_42169,N_40332,N_40594);
nand U42170 (N_42170,N_40501,N_40256);
nor U42171 (N_42171,N_41911,N_40348);
xor U42172 (N_42172,N_41426,N_41593);
nand U42173 (N_42173,N_40789,N_41002);
and U42174 (N_42174,N_40096,N_40949);
or U42175 (N_42175,N_40230,N_40688);
nand U42176 (N_42176,N_40027,N_40687);
nand U42177 (N_42177,N_41606,N_40986);
nor U42178 (N_42178,N_40061,N_41813);
nand U42179 (N_42179,N_41011,N_40136);
xor U42180 (N_42180,N_40715,N_41925);
xnor U42181 (N_42181,N_40176,N_41630);
or U42182 (N_42182,N_41412,N_40499);
and U42183 (N_42183,N_40387,N_41050);
and U42184 (N_42184,N_41528,N_41170);
nand U42185 (N_42185,N_40432,N_40842);
xnor U42186 (N_42186,N_41084,N_41192);
nor U42187 (N_42187,N_41152,N_41622);
or U42188 (N_42188,N_41573,N_40436);
and U42189 (N_42189,N_41763,N_40262);
and U42190 (N_42190,N_40416,N_40402);
xor U42191 (N_42191,N_41022,N_41063);
xnor U42192 (N_42192,N_41245,N_41081);
nand U42193 (N_42193,N_40331,N_41722);
or U42194 (N_42194,N_40790,N_40941);
nand U42195 (N_42195,N_41291,N_40413);
and U42196 (N_42196,N_41201,N_41766);
xor U42197 (N_42197,N_40426,N_40520);
xnor U42198 (N_42198,N_40991,N_41339);
or U42199 (N_42199,N_40368,N_40504);
xnor U42200 (N_42200,N_40023,N_41178);
nor U42201 (N_42201,N_41310,N_41384);
and U42202 (N_42202,N_40403,N_40327);
nor U42203 (N_42203,N_41255,N_40984);
nor U42204 (N_42204,N_41126,N_41243);
or U42205 (N_42205,N_41260,N_41466);
xnor U42206 (N_42206,N_40471,N_40502);
nand U42207 (N_42207,N_40758,N_41611);
and U42208 (N_42208,N_41847,N_41923);
and U42209 (N_42209,N_41927,N_40401);
or U42210 (N_42210,N_40253,N_40695);
and U42211 (N_42211,N_40174,N_40812);
nand U42212 (N_42212,N_41270,N_41822);
or U42213 (N_42213,N_41015,N_40393);
nand U42214 (N_42214,N_40850,N_40448);
and U42215 (N_42215,N_41750,N_40699);
xnor U42216 (N_42216,N_41760,N_40464);
and U42217 (N_42217,N_41263,N_40914);
and U42218 (N_42218,N_41337,N_40500);
nand U42219 (N_42219,N_40003,N_41744);
xnor U42220 (N_42220,N_41734,N_40370);
nor U42221 (N_42221,N_41889,N_40616);
and U42222 (N_42222,N_40190,N_41685);
nor U42223 (N_42223,N_40796,N_40457);
or U42224 (N_42224,N_40686,N_40983);
and U42225 (N_42225,N_40303,N_40996);
xor U42226 (N_42226,N_40057,N_41628);
or U42227 (N_42227,N_41338,N_41945);
nor U42228 (N_42228,N_40811,N_41217);
xor U42229 (N_42229,N_41551,N_40382);
nand U42230 (N_42230,N_41086,N_41433);
or U42231 (N_42231,N_40598,N_40314);
nor U42232 (N_42232,N_41220,N_40804);
nor U42233 (N_42233,N_41148,N_41259);
nor U42234 (N_42234,N_41755,N_41444);
or U42235 (N_42235,N_40279,N_41400);
xor U42236 (N_42236,N_40490,N_40814);
xnor U42237 (N_42237,N_41071,N_41068);
xor U42238 (N_42238,N_41697,N_40706);
nor U42239 (N_42239,N_40791,N_41533);
xor U42240 (N_42240,N_40810,N_40588);
or U42241 (N_42241,N_41652,N_40852);
nor U42242 (N_42242,N_41213,N_41262);
xnor U42243 (N_42243,N_40018,N_41793);
nor U42244 (N_42244,N_41865,N_41392);
or U42245 (N_42245,N_40944,N_40482);
or U42246 (N_42246,N_40458,N_41575);
nand U42247 (N_42247,N_40820,N_40153);
and U42248 (N_42248,N_41090,N_40795);
nor U42249 (N_42249,N_40127,N_41459);
and U42250 (N_42250,N_40940,N_41495);
nand U42251 (N_42251,N_40103,N_40523);
nand U42252 (N_42252,N_40963,N_40264);
and U42253 (N_42253,N_40330,N_40506);
xnor U42254 (N_42254,N_41798,N_41239);
xnor U42255 (N_42255,N_41664,N_41164);
nand U42256 (N_42256,N_41646,N_41448);
xnor U42257 (N_42257,N_41393,N_41680);
nand U42258 (N_42258,N_40145,N_41471);
and U42259 (N_42259,N_41128,N_41641);
nand U42260 (N_42260,N_41686,N_40473);
xor U42261 (N_42261,N_41663,N_41529);
nand U42262 (N_42262,N_41757,N_40081);
xnor U42263 (N_42263,N_40979,N_40447);
nor U42264 (N_42264,N_41238,N_40175);
and U42265 (N_42265,N_41645,N_40666);
or U42266 (N_42266,N_41513,N_40516);
nand U42267 (N_42267,N_40169,N_41316);
or U42268 (N_42268,N_41941,N_40969);
or U42269 (N_42269,N_41905,N_41897);
nor U42270 (N_42270,N_41812,N_40349);
nand U42271 (N_42271,N_41506,N_41147);
nand U42272 (N_42272,N_40602,N_40736);
and U42273 (N_42273,N_40966,N_40851);
or U42274 (N_42274,N_40573,N_40819);
nor U42275 (N_42275,N_41912,N_41095);
nor U42276 (N_42276,N_41127,N_40876);
nor U42277 (N_42277,N_40882,N_40086);
or U42278 (N_42278,N_40603,N_40272);
nor U42279 (N_42279,N_41117,N_41367);
and U42280 (N_42280,N_41182,N_41009);
nor U42281 (N_42281,N_40075,N_41918);
and U42282 (N_42282,N_41676,N_40137);
xor U42283 (N_42283,N_40772,N_41703);
nor U42284 (N_42284,N_41091,N_41518);
nand U42285 (N_42285,N_40313,N_41018);
and U42286 (N_42286,N_41708,N_41157);
and U42287 (N_42287,N_41062,N_40396);
nor U42288 (N_42288,N_41904,N_41549);
xnor U42289 (N_42289,N_40713,N_41288);
nor U42290 (N_42290,N_41767,N_41234);
nand U42291 (N_42291,N_40917,N_41696);
and U42292 (N_42292,N_40204,N_40212);
or U42293 (N_42293,N_40668,N_40031);
or U42294 (N_42294,N_40771,N_41978);
nor U42295 (N_42295,N_41782,N_41428);
or U42296 (N_42296,N_40429,N_40545);
nor U42297 (N_42297,N_41560,N_40840);
xnor U42298 (N_42298,N_41194,N_41368);
xnor U42299 (N_42299,N_41737,N_40802);
nor U42300 (N_42300,N_40530,N_41907);
nor U42301 (N_42301,N_40693,N_41728);
or U42302 (N_42302,N_41258,N_41559);
and U42303 (N_42303,N_40878,N_40879);
or U42304 (N_42304,N_41096,N_41693);
nand U42305 (N_42305,N_41932,N_41269);
or U42306 (N_42306,N_41407,N_40865);
or U42307 (N_42307,N_41456,N_41226);
nor U42308 (N_42308,N_41076,N_40194);
nand U42309 (N_42309,N_41045,N_40400);
nand U42310 (N_42310,N_41052,N_41059);
or U42311 (N_42311,N_41200,N_40408);
nand U42312 (N_42312,N_40113,N_40420);
nor U42313 (N_42313,N_40277,N_41429);
and U42314 (N_42314,N_41372,N_41342);
xor U42315 (N_42315,N_40677,N_41597);
or U42316 (N_42316,N_40838,N_40580);
or U42317 (N_42317,N_41668,N_41293);
nor U42318 (N_42318,N_40129,N_40013);
xnor U42319 (N_42319,N_41284,N_40025);
nand U42320 (N_42320,N_40242,N_41629);
nor U42321 (N_42321,N_40259,N_40751);
nor U42322 (N_42322,N_41300,N_41143);
nor U42323 (N_42323,N_40856,N_40060);
and U42324 (N_42324,N_41298,N_41406);
or U42325 (N_42325,N_41807,N_41717);
xor U42326 (N_42326,N_40581,N_41810);
nand U42327 (N_42327,N_41215,N_40824);
xnor U42328 (N_42328,N_41803,N_41458);
or U42329 (N_42329,N_41447,N_40844);
xnor U42330 (N_42330,N_40813,N_40229);
nand U42331 (N_42331,N_41166,N_41241);
xor U42332 (N_42332,N_40883,N_40377);
xnor U42333 (N_42333,N_40462,N_40849);
or U42334 (N_42334,N_40689,N_41701);
nand U42335 (N_42335,N_41856,N_41866);
nor U42336 (N_42336,N_40391,N_40992);
nor U42337 (N_42337,N_40753,N_40938);
xnor U42338 (N_42338,N_41681,N_40439);
xnor U42339 (N_42339,N_41505,N_40740);
and U42340 (N_42340,N_41118,N_40663);
and U42341 (N_42341,N_40958,N_41720);
or U42342 (N_42342,N_40972,N_40365);
xnor U42343 (N_42343,N_41364,N_41275);
xnor U42344 (N_42344,N_40388,N_41638);
nand U42345 (N_42345,N_40769,N_41948);
nor U42346 (N_42346,N_41759,N_40643);
or U42347 (N_42347,N_40041,N_41098);
nor U42348 (N_42348,N_40427,N_40599);
nor U42349 (N_42349,N_40238,N_41609);
and U42350 (N_42350,N_41079,N_40798);
nand U42351 (N_42351,N_40536,N_41543);
or U42352 (N_42352,N_41819,N_41540);
or U42353 (N_42353,N_41857,N_40592);
xnor U42354 (N_42354,N_40543,N_40988);
nor U42355 (N_42355,N_40503,N_41104);
xor U42356 (N_42356,N_40288,N_40652);
nor U42357 (N_42357,N_40243,N_41056);
nor U42358 (N_42358,N_41612,N_40373);
xor U42359 (N_42359,N_41107,N_41979);
or U42360 (N_42360,N_41613,N_41424);
and U42361 (N_42361,N_40214,N_40716);
and U42362 (N_42362,N_40962,N_40049);
nor U42363 (N_42363,N_40509,N_40563);
and U42364 (N_42364,N_40557,N_41249);
nand U42365 (N_42365,N_40344,N_40151);
xnor U42366 (N_42366,N_41289,N_40128);
xor U42367 (N_42367,N_40615,N_40936);
nor U42368 (N_42368,N_41395,N_41620);
xor U42369 (N_42369,N_40302,N_40104);
and U42370 (N_42370,N_41844,N_41743);
or U42371 (N_42371,N_40183,N_40742);
and U42372 (N_42372,N_40894,N_40714);
or U42373 (N_42373,N_40725,N_41898);
nor U42374 (N_42374,N_40281,N_40244);
xor U42375 (N_42375,N_41252,N_41761);
nand U42376 (N_42376,N_41061,N_41587);
and U42377 (N_42377,N_41473,N_40449);
and U42378 (N_42378,N_40045,N_40641);
or U42379 (N_42379,N_41527,N_40380);
or U42380 (N_42380,N_40570,N_41541);
nor U42381 (N_42381,N_41975,N_41883);
and U42382 (N_42382,N_41768,N_40394);
or U42383 (N_42383,N_41353,N_40015);
nand U42384 (N_42384,N_40955,N_40745);
nor U42385 (N_42385,N_41003,N_41186);
xnor U42386 (N_42386,N_40696,N_41503);
and U42387 (N_42387,N_41794,N_40254);
and U42388 (N_42388,N_41378,N_40897);
nor U42389 (N_42389,N_40632,N_41834);
nor U42390 (N_42390,N_40126,N_41933);
or U42391 (N_42391,N_40260,N_40793);
xor U42392 (N_42392,N_41021,N_40177);
or U42393 (N_42393,N_40885,N_40247);
and U42394 (N_42394,N_41115,N_40858);
xnor U42395 (N_42395,N_40562,N_41434);
nor U42396 (N_42396,N_41935,N_41196);
xnor U42397 (N_42397,N_40336,N_40857);
xnor U42398 (N_42398,N_41491,N_40896);
or U42399 (N_42399,N_40222,N_40806);
nand U42400 (N_42400,N_41913,N_40160);
nor U42401 (N_42401,N_40120,N_41566);
and U42402 (N_42402,N_41116,N_41419);
nor U42403 (N_42403,N_40364,N_41343);
and U42404 (N_42404,N_41179,N_40782);
nor U42405 (N_42405,N_40361,N_40765);
nor U42406 (N_42406,N_40692,N_40803);
and U42407 (N_42407,N_40062,N_40029);
nor U42408 (N_42408,N_40701,N_40087);
nand U42409 (N_42409,N_41493,N_40450);
xnor U42410 (N_42410,N_41881,N_40333);
or U42411 (N_42411,N_41644,N_40867);
and U42412 (N_42412,N_40510,N_41349);
xor U42413 (N_42413,N_40836,N_41075);
nand U42414 (N_42414,N_40477,N_40100);
nand U42415 (N_42415,N_40163,N_41616);
or U42416 (N_42416,N_41859,N_40855);
or U42417 (N_42417,N_41029,N_40399);
nor U42418 (N_42418,N_41538,N_40913);
or U42419 (N_42419,N_40756,N_40959);
xnor U42420 (N_42420,N_40767,N_41219);
xor U42421 (N_42421,N_41949,N_41047);
nor U42422 (N_42422,N_40487,N_41632);
nor U42423 (N_42423,N_41365,N_41017);
xor U42424 (N_42424,N_40871,N_40146);
nor U42425 (N_42425,N_41631,N_40094);
nand U42426 (N_42426,N_41988,N_40485);
xor U42427 (N_42427,N_41607,N_40355);
nor U42428 (N_42428,N_41640,N_40240);
and U42429 (N_42429,N_40266,N_41565);
xnor U42430 (N_42430,N_40651,N_41402);
nor U42431 (N_42431,N_41715,N_40132);
nand U42432 (N_42432,N_41572,N_41639);
nor U42433 (N_42433,N_41752,N_41498);
nor U42434 (N_42434,N_40779,N_41863);
nand U42435 (N_42435,N_41785,N_41313);
nor U42436 (N_42436,N_40662,N_41778);
or U42437 (N_42437,N_40350,N_41080);
nor U42438 (N_42438,N_40633,N_40626);
nor U42439 (N_42439,N_41675,N_40712);
nand U42440 (N_42440,N_40763,N_41043);
xnor U42441 (N_42441,N_40182,N_40923);
and U42442 (N_42442,N_41901,N_40273);
and U42443 (N_42443,N_41141,N_41446);
or U42444 (N_42444,N_41452,N_41899);
nand U42445 (N_42445,N_41162,N_40975);
or U42446 (N_42446,N_41770,N_41726);
nand U42447 (N_42447,N_40607,N_40527);
or U42448 (N_42448,N_41741,N_40531);
xnor U42449 (N_42449,N_40406,N_41235);
nand U42450 (N_42450,N_41067,N_41030);
and U42451 (N_42451,N_40173,N_40180);
or U42452 (N_42452,N_41591,N_41698);
or U42453 (N_42453,N_40935,N_41013);
or U42454 (N_42454,N_40189,N_41937);
or U42455 (N_42455,N_41360,N_40971);
nor U42456 (N_42456,N_41404,N_41702);
nand U42457 (N_42457,N_40550,N_41799);
nor U42458 (N_42458,N_41624,N_40048);
and U42459 (N_42459,N_40583,N_41122);
nor U42460 (N_42460,N_41180,N_40737);
nor U42461 (N_42461,N_41007,N_40522);
or U42462 (N_42462,N_40707,N_40335);
xnor U42463 (N_42463,N_41828,N_41183);
nand U42464 (N_42464,N_41228,N_41700);
nor U42465 (N_42465,N_40956,N_40080);
nand U42466 (N_42466,N_40625,N_41145);
and U42467 (N_42467,N_40028,N_41501);
nor U42468 (N_42468,N_40629,N_41914);
and U42469 (N_42469,N_41853,N_40990);
xnor U42470 (N_42470,N_40334,N_41986);
nand U42471 (N_42471,N_41657,N_41909);
or U42472 (N_42472,N_40847,N_41329);
or U42473 (N_42473,N_41415,N_40600);
or U42474 (N_42474,N_40612,N_41962);
nand U42475 (N_42475,N_40157,N_40287);
or U42476 (N_42476,N_41677,N_41092);
and U42477 (N_42477,N_40064,N_40881);
and U42478 (N_42478,N_40360,N_41099);
xnor U42479 (N_42479,N_40034,N_41042);
nor U42480 (N_42480,N_40390,N_40912);
nor U42481 (N_42481,N_40567,N_40694);
xnor U42482 (N_42482,N_40731,N_41136);
xor U42483 (N_42483,N_40282,N_40300);
nor U42484 (N_42484,N_40826,N_40827);
nand U42485 (N_42485,N_40553,N_40188);
nand U42486 (N_42486,N_40141,N_41309);
or U42487 (N_42487,N_40965,N_41461);
nor U42488 (N_42488,N_40142,N_41492);
and U42489 (N_42489,N_40056,N_40409);
nor U42490 (N_42490,N_40460,N_40050);
nand U42491 (N_42491,N_41626,N_41547);
nand U42492 (N_42492,N_40650,N_41796);
xnor U42493 (N_42493,N_41951,N_40799);
xor U42494 (N_42494,N_40862,N_40674);
nor U42495 (N_42495,N_41417,N_41221);
and U42496 (N_42496,N_40209,N_40513);
nor U42497 (N_42497,N_40434,N_40555);
and U42498 (N_42498,N_40711,N_40424);
and U42499 (N_42499,N_41087,N_41210);
or U42500 (N_42500,N_41678,N_41504);
nand U42501 (N_42501,N_40263,N_41478);
nand U42502 (N_42502,N_40371,N_41089);
xor U42503 (N_42503,N_41690,N_41636);
or U42504 (N_42504,N_41998,N_40646);
and U42505 (N_42505,N_41248,N_41637);
xor U42506 (N_42506,N_41191,N_40746);
xor U42507 (N_42507,N_40474,N_40915);
nand U42508 (N_42508,N_40576,N_40942);
nand U42509 (N_42509,N_40042,N_41851);
and U42510 (N_42510,N_41273,N_40784);
xnor U42511 (N_42511,N_41324,N_41520);
or U42512 (N_42512,N_41500,N_40559);
nor U42513 (N_42513,N_41525,N_40571);
and U42514 (N_42514,N_41040,N_40304);
or U42515 (N_42515,N_40179,N_41207);
xnor U42516 (N_42516,N_40978,N_41066);
nand U42517 (N_42517,N_40430,N_40375);
and U42518 (N_42518,N_40372,N_41839);
nand U42519 (N_42519,N_40928,N_41133);
or U42520 (N_42520,N_41023,N_41614);
xnor U42521 (N_42521,N_40299,N_41919);
and U42522 (N_42522,N_40816,N_41212);
or U42523 (N_42523,N_40232,N_41787);
nor U42524 (N_42524,N_41380,N_40359);
and U42525 (N_42525,N_41103,N_41105);
or U42526 (N_42526,N_40152,N_41227);
and U42527 (N_42527,N_40743,N_40069);
and U42528 (N_42528,N_41282,N_40193);
nand U42529 (N_42529,N_41124,N_40548);
and U42530 (N_42530,N_40738,N_40584);
xor U42531 (N_42531,N_40001,N_40412);
nand U42532 (N_42532,N_41151,N_41832);
xnor U42533 (N_42533,N_41203,N_40066);
or U42534 (N_42534,N_41875,N_41902);
nor U42535 (N_42535,N_40004,N_41172);
nor U42536 (N_42536,N_40021,N_41751);
nor U42537 (N_42537,N_41771,N_40397);
nand U42538 (N_42538,N_41073,N_41094);
and U42539 (N_42539,N_40601,N_40297);
xor U42540 (N_42540,N_40385,N_41333);
and U42541 (N_42541,N_41430,N_41450);
nor U42542 (N_42542,N_41576,N_40443);
nand U42543 (N_42543,N_41991,N_41672);
nand U42544 (N_42544,N_41818,N_41457);
xnor U42545 (N_42545,N_40618,N_41156);
xnor U42546 (N_42546,N_40676,N_40829);
nor U42547 (N_42547,N_40054,N_41358);
nor U42548 (N_42548,N_40683,N_40491);
and U42549 (N_42549,N_40660,N_41474);
xnor U42550 (N_42550,N_40889,N_40469);
nor U42551 (N_42551,N_40937,N_41589);
nor U42552 (N_42552,N_40352,N_41601);
nand U42553 (N_42553,N_41223,N_40067);
and U42554 (N_42554,N_41692,N_41841);
nor U42555 (N_42555,N_40140,N_40669);
xor U42556 (N_42556,N_40376,N_40525);
and U42557 (N_42557,N_41283,N_41311);
and U42558 (N_42558,N_40398,N_41476);
and U42559 (N_42559,N_41027,N_40118);
nand U42560 (N_42560,N_41173,N_40381);
and U42561 (N_42561,N_40875,N_41229);
nand U42562 (N_42562,N_40930,N_41558);
xor U42563 (N_42563,N_40110,N_41821);
nor U42564 (N_42564,N_41727,N_40148);
nand U42565 (N_42565,N_41453,N_41382);
nor U42566 (N_42566,N_40639,N_41623);
and U42567 (N_42567,N_41049,N_41051);
nand U42568 (N_42568,N_40167,N_40392);
and U42569 (N_42569,N_41598,N_40454);
xor U42570 (N_42570,N_41438,N_40245);
or U42571 (N_42571,N_41874,N_41377);
nor U42572 (N_42572,N_41656,N_40835);
nor U42573 (N_42573,N_40568,N_41649);
xor U42574 (N_42574,N_41195,N_40542);
and U42575 (N_42575,N_41879,N_41855);
or U42576 (N_42576,N_40951,N_41074);
xor U42577 (N_42577,N_41669,N_41366);
and U42578 (N_42578,N_40967,N_40901);
nand U42579 (N_42579,N_41512,N_41197);
and U42580 (N_42580,N_41363,N_40556);
nand U42581 (N_42581,N_40010,N_41479);
nor U42582 (N_42582,N_40931,N_41435);
and U42583 (N_42583,N_40943,N_40741);
and U42584 (N_42584,N_40453,N_41729);
and U42585 (N_42585,N_40033,N_41781);
or U42586 (N_42586,N_41386,N_41112);
nor U42587 (N_42587,N_40475,N_40684);
nand U42588 (N_42588,N_40617,N_40047);
xnor U42589 (N_42589,N_40579,N_41463);
xor U42590 (N_42590,N_41371,N_40224);
or U42591 (N_42591,N_41797,N_41666);
or U42592 (N_42592,N_41198,N_41475);
and U42593 (N_42593,N_41296,N_41848);
xnor U42594 (N_42594,N_40925,N_41952);
nand U42595 (N_42595,N_41469,N_40178);
or U42596 (N_42596,N_40645,N_41484);
nor U42597 (N_42597,N_41970,N_40171);
nand U42598 (N_42598,N_40317,N_40671);
and U42599 (N_42599,N_40476,N_41405);
nor U42600 (N_42600,N_40130,N_40968);
nand U42601 (N_42601,N_40417,N_40586);
nor U42602 (N_42602,N_40899,N_40078);
and U42603 (N_42603,N_40734,N_40918);
xor U42604 (N_42604,N_41222,N_41600);
nand U42605 (N_42605,N_41635,N_40016);
nand U42606 (N_42606,N_41765,N_40073);
or U42607 (N_42607,N_40239,N_40906);
and U42608 (N_42608,N_41740,N_41472);
and U42609 (N_42609,N_40326,N_40608);
nor U42610 (N_42610,N_40425,N_41557);
or U42611 (N_42611,N_40621,N_40306);
and U42612 (N_42612,N_40201,N_41348);
or U42613 (N_42613,N_41031,N_40323);
nor U42614 (N_42614,N_40910,N_40316);
xnor U42615 (N_42615,N_40328,N_41779);
nand U42616 (N_42616,N_41140,N_41214);
and U42617 (N_42617,N_40083,N_40549);
and U42618 (N_42618,N_41896,N_41057);
nand U42619 (N_42619,N_41964,N_40873);
nor U42620 (N_42620,N_40636,N_40884);
nor U42621 (N_42621,N_40539,N_41667);
or U42622 (N_42622,N_41957,N_40389);
xor U42623 (N_42623,N_40112,N_40532);
or U42624 (N_42624,N_40337,N_41982);
and U42625 (N_42625,N_41155,N_41486);
nand U42626 (N_42626,N_40071,N_40869);
nor U42627 (N_42627,N_40726,N_41783);
nand U42628 (N_42628,N_41563,N_40164);
xnor U42629 (N_42629,N_41230,N_41554);
nor U42630 (N_42630,N_40964,N_41745);
and U42631 (N_42631,N_40597,N_40916);
or U42632 (N_42632,N_41374,N_41938);
xor U42633 (N_42633,N_41679,N_40997);
nand U42634 (N_42634,N_41562,N_41604);
and U42635 (N_42635,N_41169,N_40752);
nor U42636 (N_42636,N_41608,N_41825);
xnor U42637 (N_42637,N_40511,N_40495);
or U42638 (N_42638,N_41502,N_40690);
xnor U42639 (N_42639,N_41647,N_40005);
or U42640 (N_42640,N_41242,N_40544);
nand U42641 (N_42641,N_41961,N_40150);
and U42642 (N_42642,N_41921,N_41250);
and U42643 (N_42643,N_40628,N_40404);
and U42644 (N_42644,N_41594,N_41537);
nand U42645 (N_42645,N_41683,N_40419);
xnor U42646 (N_42646,N_40115,N_41490);
and U42647 (N_42647,N_40624,N_41174);
and U42648 (N_42648,N_40207,N_41302);
xor U42649 (N_42649,N_40945,N_40783);
nand U42650 (N_42650,N_41826,N_41381);
nand U42651 (N_42651,N_40318,N_40927);
nor U42652 (N_42652,N_40139,N_41955);
nor U42653 (N_42653,N_41758,N_40981);
xnor U42654 (N_42654,N_40270,N_40052);
xnor U42655 (N_42655,N_41344,N_41272);
and U42656 (N_42656,N_40957,N_40496);
nand U42657 (N_42657,N_41849,N_40428);
or U42658 (N_42658,N_41036,N_41441);
and U42659 (N_42659,N_40102,N_40065);
nand U42660 (N_42660,N_41689,N_40379);
nand U42661 (N_42661,N_40486,N_41582);
xnor U42662 (N_42662,N_40895,N_40982);
and U42663 (N_42663,N_41418,N_40311);
xnor U42664 (N_42664,N_41924,N_41160);
nand U42665 (N_42665,N_40585,N_40265);
or U42666 (N_42666,N_41069,N_40823);
nor U42667 (N_42667,N_41034,N_40074);
nand U42668 (N_42668,N_41809,N_41391);
or U42669 (N_42669,N_41295,N_40560);
xnor U42670 (N_42670,N_41733,N_40691);
xor U42671 (N_42671,N_40438,N_41487);
and U42672 (N_42672,N_40866,N_40710);
and U42673 (N_42673,N_41204,N_41953);
nor U42674 (N_42674,N_40661,N_41443);
xnor U42675 (N_42675,N_40703,N_40084);
nand U42676 (N_42676,N_40079,N_40198);
nand U42677 (N_42677,N_40040,N_41596);
nor U42678 (N_42678,N_41655,N_41330);
nand U42679 (N_42679,N_41780,N_41795);
nor U42680 (N_42680,N_41769,N_41738);
xor U42681 (N_42681,N_41347,N_41931);
and U42682 (N_42682,N_41286,N_40124);
xnor U42683 (N_42683,N_40672,N_41651);
nor U42684 (N_42684,N_40077,N_40456);
nor U42685 (N_42685,N_41314,N_41954);
nor U42686 (N_42686,N_40206,N_40547);
xnor U42687 (N_42687,N_41409,N_41425);
nand U42688 (N_42688,N_41306,N_40774);
nand U42689 (N_42689,N_41370,N_40480);
or U42690 (N_42690,N_40841,N_41688);
nor U42691 (N_42691,N_41176,N_40024);
nor U42692 (N_42692,N_41583,N_41465);
nand U42693 (N_42693,N_40405,N_40744);
xor U42694 (N_42694,N_41578,N_41149);
nand U42695 (N_42695,N_40467,N_40442);
or U42696 (N_42696,N_41929,N_40644);
nor U42697 (N_42697,N_40566,N_41085);
or U42698 (N_42698,N_41336,N_41539);
or U42699 (N_42699,N_40329,N_40932);
or U42700 (N_42700,N_41421,N_41411);
nand U42701 (N_42701,N_40290,N_41006);
nor U42702 (N_42702,N_41872,N_40704);
xnor U42703 (N_42703,N_41482,N_41489);
nand U42704 (N_42704,N_40825,N_41661);
xnor U42705 (N_42705,N_40670,N_40338);
xnor U42706 (N_42706,N_41773,N_40231);
and U42707 (N_42707,N_40762,N_41060);
and U42708 (N_42708,N_40097,N_41168);
nor U42709 (N_42709,N_40754,N_40719);
xor U42710 (N_42710,N_40470,N_41877);
xor U42711 (N_42711,N_40514,N_40818);
and U42712 (N_42712,N_40168,N_40606);
or U42713 (N_42713,N_40970,N_40919);
nand U42714 (N_42714,N_40721,N_41994);
nand U42715 (N_42715,N_41969,N_41691);
or U42716 (N_42716,N_41756,N_41511);
nor U42717 (N_42717,N_41420,N_41530);
nand U42718 (N_42718,N_41928,N_40589);
and U42719 (N_42719,N_40837,N_41327);
and U42720 (N_42720,N_40466,N_41777);
nand U42721 (N_42721,N_40008,N_40324);
nor U42722 (N_42722,N_41285,N_41398);
nor U42723 (N_42723,N_41542,N_40200);
or U42724 (N_42724,N_40526,N_41139);
nor U42725 (N_42725,N_41005,N_40533);
and U42726 (N_42726,N_41873,N_41256);
xnor U42727 (N_42727,N_40309,N_41064);
nand U42728 (N_42728,N_40046,N_41642);
or U42729 (N_42729,N_41334,N_40718);
xnor U42730 (N_42730,N_40893,N_41154);
and U42731 (N_42731,N_40165,N_41965);
nor U42732 (N_42732,N_41008,N_40134);
nor U42733 (N_42733,N_41526,N_41671);
xnor U42734 (N_42734,N_41055,N_41340);
and U42735 (N_42735,N_40170,N_41102);
nand U42736 (N_42736,N_40116,N_41864);
xnor U42737 (N_42737,N_40622,N_40166);
xnor U42738 (N_42738,N_41956,N_41389);
or U42739 (N_42739,N_41449,N_41508);
xnor U42740 (N_42740,N_41595,N_41237);
or U42741 (N_42741,N_40578,N_40044);
nand U42742 (N_42742,N_40805,N_40356);
or U42743 (N_42743,N_40730,N_40787);
or U42744 (N_42744,N_40345,N_41394);
xnor U42745 (N_42745,N_41468,N_40386);
nand U42746 (N_42746,N_40091,N_40410);
nor U42747 (N_42747,N_41292,N_41379);
xnor U42748 (N_42748,N_40552,N_40739);
or U42749 (N_42749,N_40994,N_41058);
nor U42750 (N_42750,N_40121,N_41922);
and U42751 (N_42751,N_40433,N_40210);
nor U42752 (N_42752,N_40257,N_40411);
xnor U42753 (N_42753,N_41375,N_40294);
xor U42754 (N_42754,N_40208,N_40415);
xnor U42755 (N_42755,N_40192,N_41996);
and U42756 (N_42756,N_41586,N_41724);
and U42757 (N_42757,N_41947,N_40541);
or U42758 (N_42758,N_41357,N_41494);
nor U42759 (N_42759,N_40223,N_41000);
nor U42760 (N_42760,N_41971,N_40216);
xor U42761 (N_42761,N_41261,N_40630);
or U42762 (N_42762,N_40973,N_40123);
nand U42763 (N_42763,N_40340,N_40205);
xnor U42764 (N_42764,N_41892,N_41966);
xor U42765 (N_42765,N_40929,N_40271);
nand U42766 (N_42766,N_40159,N_41561);
or U42767 (N_42767,N_41983,N_40357);
or U42768 (N_42768,N_40423,N_41341);
and U42769 (N_42769,N_41354,N_40702);
nand U42770 (N_42770,N_41208,N_40211);
xor U42771 (N_42771,N_41625,N_41711);
or U42772 (N_42772,N_41735,N_40947);
nand U42773 (N_42773,N_41120,N_41915);
or U42774 (N_42774,N_41850,N_40843);
nor U42775 (N_42775,N_40301,N_41125);
or U42776 (N_42776,N_41001,N_40276);
nor U42777 (N_42777,N_40144,N_41764);
xor U42778 (N_42778,N_40667,N_41097);
or U42779 (N_42779,N_41004,N_40455);
or U42780 (N_42780,N_40149,N_40735);
and U42781 (N_42781,N_41308,N_40521);
nor U42782 (N_42782,N_40421,N_40237);
nand U42783 (N_42783,N_41618,N_41224);
nand U42784 (N_42784,N_41020,N_41111);
nand U42785 (N_42785,N_41236,N_41852);
and U42786 (N_42786,N_40909,N_41934);
and U42787 (N_42787,N_41723,N_40998);
or U42788 (N_42788,N_41401,N_40685);
nor U42789 (N_42789,N_41352,N_40320);
or U42790 (N_42790,N_40546,N_40887);
nor U42791 (N_42791,N_40122,N_41775);
xor U42792 (N_42792,N_40000,N_40250);
nor U42793 (N_42793,N_40038,N_41792);
or U42794 (N_42794,N_40921,N_41362);
and U42795 (N_42795,N_41747,N_40974);
and U42796 (N_42796,N_41278,N_40383);
and U42797 (N_42797,N_40635,N_41359);
xor U42798 (N_42798,N_40678,N_40764);
and U42799 (N_42799,N_40868,N_40822);
and U42800 (N_42800,N_41739,N_41854);
and U42801 (N_42801,N_40068,N_40792);
or U42802 (N_42802,N_40489,N_41658);
xnor U42803 (N_42803,N_41833,N_40213);
and U42804 (N_42804,N_40950,N_40032);
or U42805 (N_42805,N_41356,N_40770);
or U42806 (N_42806,N_41886,N_40395);
or U42807 (N_42807,N_41571,N_40848);
and U42808 (N_42808,N_41706,N_41163);
and U42809 (N_42809,N_40341,N_40727);
xor U42810 (N_42810,N_40172,N_40006);
or U42811 (N_42811,N_41271,N_40058);
nor U42812 (N_42812,N_40786,N_41930);
nand U42813 (N_42813,N_41876,N_41916);
xnor U42814 (N_42814,N_40227,N_41290);
nor U42815 (N_42815,N_40733,N_41028);
nor U42816 (N_42816,N_41413,N_41976);
xnor U42817 (N_42817,N_40561,N_40292);
xnor U42818 (N_42818,N_41823,N_41548);
nor U42819 (N_42819,N_40384,N_40191);
or U42820 (N_42820,N_41654,N_41016);
or U42821 (N_42821,N_41046,N_40620);
nand U42822 (N_42822,N_40125,N_40697);
nand U42823 (N_42823,N_40720,N_40020);
or U42824 (N_42824,N_40362,N_40114);
and U42825 (N_42825,N_41053,N_41694);
and U42826 (N_42826,N_41590,N_40709);
xor U42827 (N_42827,N_41709,N_41784);
nand U42828 (N_42828,N_40565,N_40251);
nand U42829 (N_42829,N_40226,N_41840);
xor U42830 (N_42830,N_41868,N_41992);
and U42831 (N_42831,N_40839,N_40512);
or U42832 (N_42832,N_41940,N_41403);
nand U42833 (N_42833,N_40773,N_41390);
nor U42834 (N_42834,N_40310,N_41730);
nand U42835 (N_42835,N_41445,N_40036);
nor U42836 (N_42836,N_41824,N_41522);
nand U42837 (N_42837,N_41012,N_41297);
xnor U42838 (N_42838,N_41890,N_40154);
nand U42839 (N_42839,N_41958,N_40053);
nor U42840 (N_42840,N_41462,N_41317);
nor U42841 (N_42841,N_40631,N_40728);
or U42842 (N_42842,N_40655,N_40295);
or U42843 (N_42843,N_41574,N_40780);
nor U42844 (N_42844,N_41244,N_41524);
nand U42845 (N_42845,N_41510,N_41427);
or U42846 (N_42846,N_40989,N_40017);
nor U42847 (N_42847,N_40903,N_41065);
nor U42848 (N_42848,N_40613,N_41177);
and U42849 (N_42849,N_41158,N_41963);
xor U42850 (N_42850,N_41206,N_41240);
and U42851 (N_42851,N_40891,N_40833);
and U42852 (N_42852,N_41665,N_40638);
or U42853 (N_42853,N_40444,N_41816);
nand U42854 (N_42854,N_40619,N_41432);
nand U42855 (N_42855,N_41817,N_40088);
and U42856 (N_42856,N_41451,N_41716);
and U42857 (N_42857,N_41231,N_40059);
and U42858 (N_42858,N_40647,N_40218);
nand U42859 (N_42859,N_41553,N_40155);
xnor U42860 (N_42860,N_40267,N_41320);
xor U42861 (N_42861,N_40682,N_41514);
xnor U42862 (N_42862,N_40534,N_40977);
or U42863 (N_42863,N_40564,N_40445);
nor U42864 (N_42864,N_40604,N_40593);
nand U42865 (N_42865,N_40845,N_40952);
nor U42866 (N_42866,N_41257,N_40587);
nor U42867 (N_42867,N_40673,N_40698);
and U42868 (N_42868,N_40659,N_41199);
nor U42869 (N_42869,N_40241,N_41820);
or U42870 (N_42870,N_41287,N_41788);
nor U42871 (N_42871,N_40322,N_40723);
or U42872 (N_42872,N_40939,N_41621);
and U42873 (N_42873,N_41861,N_40414);
nor U42874 (N_42874,N_40374,N_41523);
nand U42875 (N_42875,N_40452,N_41346);
nor U42876 (N_42876,N_41981,N_40101);
nand U42877 (N_42877,N_40554,N_40657);
nor U42878 (N_42878,N_40654,N_41570);
or U42879 (N_42879,N_40351,N_40860);
or U42880 (N_42880,N_40195,N_40574);
or U42881 (N_42881,N_41718,N_41617);
xor U42882 (N_42882,N_41121,N_41088);
xnor U42883 (N_42883,N_41535,N_41070);
nor U42884 (N_42884,N_41712,N_40877);
and U42885 (N_42885,N_40072,N_40492);
or U42886 (N_42886,N_40828,N_40729);
xor U42887 (N_42887,N_40162,N_40296);
or U42888 (N_42888,N_40493,N_41119);
nor U42889 (N_42889,N_40451,N_40976);
and U42890 (N_42890,N_41077,N_41731);
and U42891 (N_42891,N_40367,N_41532);
or U42892 (N_42892,N_41481,N_40497);
nor U42893 (N_42893,N_40009,N_41650);
and U42894 (N_42894,N_40609,N_41246);
xor U42895 (N_42895,N_41789,N_40905);
nor U42896 (N_42896,N_40095,N_40012);
nor U42897 (N_42897,N_41185,N_40610);
or U42898 (N_42898,N_41193,N_40196);
nand U42899 (N_42899,N_41385,N_41233);
nand U42900 (N_42900,N_41373,N_41266);
or U42901 (N_42901,N_40035,N_40590);
nor U42902 (N_42902,N_41048,N_41517);
nor U42903 (N_42903,N_40255,N_40760);
nor U42904 (N_42904,N_41968,N_40757);
and U42905 (N_42905,N_41888,N_41550);
nor U42906 (N_42906,N_41159,N_41602);
nand U42907 (N_42907,N_41150,N_40948);
nand U42908 (N_42908,N_40246,N_41019);
nor U42909 (N_42909,N_41946,N_40781);
xor U42910 (N_42910,N_41887,N_40759);
and U42911 (N_42911,N_41736,N_40777);
nor U42912 (N_42912,N_40874,N_40649);
xnor U42913 (N_42913,N_41138,N_41585);
xor U42914 (N_42914,N_40519,N_41322);
nor U42915 (N_42915,N_40252,N_40954);
xnor U42916 (N_42916,N_40953,N_41837);
and U42917 (N_42917,N_40900,N_41811);
nor U42918 (N_42918,N_40063,N_41959);
or U42919 (N_42919,N_41331,N_41707);
xnor U42920 (N_42920,N_41627,N_41232);
nand U42921 (N_42921,N_41190,N_41388);
nor U42922 (N_42922,N_40315,N_41555);
nand U42923 (N_42923,N_40732,N_40039);
nand U42924 (N_42924,N_40498,N_41437);
nand U42925 (N_42925,N_41188,N_40422);
nor U42926 (N_42926,N_40440,N_40861);
and U42927 (N_42927,N_40717,N_41987);
nand U42928 (N_42928,N_40830,N_40766);
xor U42929 (N_42929,N_41439,N_40070);
nand U42930 (N_42930,N_41569,N_41753);
xor U42931 (N_42931,N_41516,N_41830);
nor U42932 (N_42932,N_41251,N_40022);
and U42933 (N_42933,N_40342,N_40055);
and U42934 (N_42934,N_40219,N_40278);
and U42935 (N_42935,N_41791,N_40133);
xor U42936 (N_42936,N_41189,N_40569);
nand U42937 (N_42937,N_41719,N_40156);
or U42938 (N_42938,N_41488,N_41827);
or U42939 (N_42939,N_40794,N_41592);
or U42940 (N_42940,N_40407,N_40788);
xor U42941 (N_42941,N_40722,N_41790);
xor U42942 (N_42942,N_40987,N_40280);
or U42943 (N_42943,N_41531,N_41281);
or U42944 (N_42944,N_41603,N_41431);
nand U42945 (N_42945,N_41312,N_41142);
and U42946 (N_42946,N_41564,N_41318);
xnor U42947 (N_42947,N_40147,N_41894);
or U42948 (N_42948,N_41858,N_40107);
nand U42949 (N_42949,N_41078,N_41615);
or U42950 (N_42950,N_41772,N_41545);
nand U42951 (N_42951,N_41422,N_41467);
or U42952 (N_42952,N_41110,N_40437);
nand U42953 (N_42953,N_40358,N_40778);
or U42954 (N_42954,N_41721,N_41544);
or U42955 (N_42955,N_41044,N_40289);
nand U42956 (N_42956,N_41054,N_40582);
xnor U42957 (N_42957,N_41247,N_41114);
and U42958 (N_42958,N_41499,N_40596);
xnor U42959 (N_42959,N_40776,N_40888);
xnor U42960 (N_42960,N_41801,N_40926);
xor U42961 (N_42961,N_41509,N_41267);
nand U42962 (N_42962,N_41960,N_41995);
xor U42963 (N_42963,N_40347,N_40354);
or U42964 (N_42964,N_40261,N_41725);
and U42965 (N_42965,N_40037,N_40119);
nand U42966 (N_42966,N_40724,N_40339);
and U42967 (N_42967,N_41836,N_40605);
or U42968 (N_42968,N_41800,N_41605);
xor U42969 (N_42969,N_40902,N_40293);
nor U42970 (N_42970,N_40920,N_40961);
nor U42971 (N_42971,N_40291,N_40664);
and U42972 (N_42972,N_40634,N_41977);
nor U42973 (N_42973,N_41470,N_41674);
nand U42974 (N_42974,N_41171,N_41610);
xor U42975 (N_42975,N_41014,N_41713);
nand U42976 (N_42976,N_40488,N_41181);
xor U42977 (N_42977,N_40538,N_41869);
or U42978 (N_42978,N_41580,N_40312);
xnor U42979 (N_42979,N_41383,N_41397);
nand U42980 (N_42980,N_41410,N_40468);
or U42981 (N_42981,N_40908,N_41144);
or U42982 (N_42982,N_40675,N_41746);
xnor U42983 (N_42983,N_41483,N_41814);
or U42984 (N_42984,N_40508,N_40011);
nand U42985 (N_42985,N_41299,N_40524);
nor U42986 (N_42986,N_41989,N_41039);
and U42987 (N_42987,N_41808,N_40319);
nor U42988 (N_42988,N_41477,N_41670);
xor U42989 (N_42989,N_41135,N_41999);
nand U42990 (N_42990,N_40863,N_41950);
xor U42991 (N_42991,N_41123,N_40225);
nand U42992 (N_42992,N_40461,N_40105);
and U42993 (N_42993,N_40106,N_40515);
and U42994 (N_42994,N_41936,N_41025);
nand U42995 (N_42995,N_41315,N_41845);
or U42996 (N_42996,N_41519,N_41082);
or U42997 (N_42997,N_40286,N_41714);
xor U42998 (N_42998,N_41556,N_41521);
xor U42999 (N_42999,N_41167,N_40870);
and U43000 (N_43000,N_41413,N_40600);
nor U43001 (N_43001,N_41854,N_40034);
and U43002 (N_43002,N_40477,N_41997);
or U43003 (N_43003,N_40863,N_40853);
and U43004 (N_43004,N_41271,N_41430);
nand U43005 (N_43005,N_41824,N_41042);
xor U43006 (N_43006,N_41177,N_40556);
nand U43007 (N_43007,N_40571,N_41508);
xor U43008 (N_43008,N_40161,N_40246);
and U43009 (N_43009,N_41301,N_40974);
or U43010 (N_43010,N_40036,N_40071);
or U43011 (N_43011,N_40376,N_40139);
xnor U43012 (N_43012,N_41810,N_41305);
nor U43013 (N_43013,N_41915,N_41242);
nand U43014 (N_43014,N_41890,N_41337);
and U43015 (N_43015,N_40049,N_40310);
nand U43016 (N_43016,N_40854,N_40747);
nand U43017 (N_43017,N_41398,N_41530);
nand U43018 (N_43018,N_40063,N_41865);
xor U43019 (N_43019,N_40179,N_40173);
nand U43020 (N_43020,N_41285,N_40138);
or U43021 (N_43021,N_41773,N_41479);
xnor U43022 (N_43022,N_41955,N_41732);
xor U43023 (N_43023,N_40303,N_40226);
or U43024 (N_43024,N_41712,N_40976);
xor U43025 (N_43025,N_40547,N_40132);
nand U43026 (N_43026,N_41988,N_40748);
nand U43027 (N_43027,N_41519,N_41859);
and U43028 (N_43028,N_40853,N_40069);
and U43029 (N_43029,N_41115,N_40630);
xnor U43030 (N_43030,N_40510,N_40279);
and U43031 (N_43031,N_40014,N_41649);
xnor U43032 (N_43032,N_40656,N_40836);
nand U43033 (N_43033,N_40613,N_41998);
and U43034 (N_43034,N_40345,N_41891);
xor U43035 (N_43035,N_40736,N_41310);
xor U43036 (N_43036,N_40534,N_40378);
and U43037 (N_43037,N_41162,N_41941);
and U43038 (N_43038,N_40834,N_40271);
nand U43039 (N_43039,N_40591,N_40296);
nor U43040 (N_43040,N_40061,N_40745);
or U43041 (N_43041,N_40936,N_40530);
xnor U43042 (N_43042,N_40670,N_41466);
xor U43043 (N_43043,N_41714,N_40362);
and U43044 (N_43044,N_40131,N_41473);
nand U43045 (N_43045,N_40608,N_41431);
nand U43046 (N_43046,N_40440,N_40988);
nand U43047 (N_43047,N_40074,N_40322);
or U43048 (N_43048,N_40915,N_40042);
and U43049 (N_43049,N_41167,N_40812);
xnor U43050 (N_43050,N_41413,N_41854);
and U43051 (N_43051,N_41584,N_40740);
and U43052 (N_43052,N_41633,N_41701);
nor U43053 (N_43053,N_41673,N_40987);
nand U43054 (N_43054,N_41291,N_41102);
nand U43055 (N_43055,N_41648,N_41526);
nand U43056 (N_43056,N_41511,N_40535);
or U43057 (N_43057,N_40468,N_41985);
nor U43058 (N_43058,N_41830,N_41987);
and U43059 (N_43059,N_40854,N_41724);
xor U43060 (N_43060,N_40033,N_41319);
xnor U43061 (N_43061,N_40144,N_40197);
and U43062 (N_43062,N_41934,N_41861);
nand U43063 (N_43063,N_40656,N_41462);
nor U43064 (N_43064,N_40631,N_40456);
or U43065 (N_43065,N_41085,N_41972);
or U43066 (N_43066,N_41917,N_40282);
xor U43067 (N_43067,N_40790,N_40678);
nand U43068 (N_43068,N_41389,N_41009);
nor U43069 (N_43069,N_40817,N_41642);
nand U43070 (N_43070,N_41129,N_41336);
or U43071 (N_43071,N_41401,N_40983);
nor U43072 (N_43072,N_40497,N_40779);
xor U43073 (N_43073,N_40994,N_41853);
nand U43074 (N_43074,N_41522,N_40336);
xor U43075 (N_43075,N_41835,N_40583);
nand U43076 (N_43076,N_41118,N_40707);
and U43077 (N_43077,N_40811,N_41575);
xnor U43078 (N_43078,N_40856,N_41679);
nand U43079 (N_43079,N_41254,N_40426);
nand U43080 (N_43080,N_41856,N_41416);
or U43081 (N_43081,N_40450,N_41642);
xnor U43082 (N_43082,N_41062,N_40158);
and U43083 (N_43083,N_41919,N_41630);
or U43084 (N_43084,N_41633,N_41496);
and U43085 (N_43085,N_40638,N_41025);
nor U43086 (N_43086,N_40399,N_40889);
xor U43087 (N_43087,N_41393,N_41644);
and U43088 (N_43088,N_41468,N_40362);
or U43089 (N_43089,N_41014,N_40633);
nand U43090 (N_43090,N_40392,N_41425);
and U43091 (N_43091,N_40093,N_40763);
xnor U43092 (N_43092,N_41791,N_40367);
nor U43093 (N_43093,N_41969,N_41430);
xnor U43094 (N_43094,N_40682,N_41106);
xor U43095 (N_43095,N_40303,N_41733);
nand U43096 (N_43096,N_40818,N_41244);
and U43097 (N_43097,N_41603,N_41993);
nand U43098 (N_43098,N_41231,N_40245);
nand U43099 (N_43099,N_41552,N_40356);
nor U43100 (N_43100,N_40625,N_40410);
nand U43101 (N_43101,N_40076,N_41281);
nand U43102 (N_43102,N_40973,N_41556);
nand U43103 (N_43103,N_41576,N_40633);
nand U43104 (N_43104,N_41041,N_40691);
nand U43105 (N_43105,N_40869,N_41751);
xnor U43106 (N_43106,N_41118,N_40601);
xor U43107 (N_43107,N_40948,N_40033);
xor U43108 (N_43108,N_40048,N_41581);
and U43109 (N_43109,N_41027,N_41957);
or U43110 (N_43110,N_41850,N_40738);
nor U43111 (N_43111,N_40497,N_40658);
xor U43112 (N_43112,N_41395,N_41025);
xor U43113 (N_43113,N_41495,N_41367);
nor U43114 (N_43114,N_40661,N_40607);
xnor U43115 (N_43115,N_40357,N_41730);
or U43116 (N_43116,N_40876,N_41840);
or U43117 (N_43117,N_40387,N_40340);
nor U43118 (N_43118,N_40336,N_40043);
nand U43119 (N_43119,N_40933,N_40816);
and U43120 (N_43120,N_41625,N_41334);
and U43121 (N_43121,N_41195,N_40900);
and U43122 (N_43122,N_40752,N_41310);
nand U43123 (N_43123,N_40363,N_40900);
or U43124 (N_43124,N_41193,N_40863);
or U43125 (N_43125,N_40172,N_40578);
or U43126 (N_43126,N_41142,N_40477);
xor U43127 (N_43127,N_40477,N_40918);
or U43128 (N_43128,N_41132,N_40798);
nor U43129 (N_43129,N_40431,N_40374);
xnor U43130 (N_43130,N_40705,N_40232);
and U43131 (N_43131,N_41477,N_41639);
xor U43132 (N_43132,N_40996,N_41094);
or U43133 (N_43133,N_41537,N_41333);
nand U43134 (N_43134,N_40906,N_41014);
nand U43135 (N_43135,N_40696,N_40497);
and U43136 (N_43136,N_41746,N_40933);
xnor U43137 (N_43137,N_41823,N_40247);
nor U43138 (N_43138,N_40099,N_41154);
or U43139 (N_43139,N_40198,N_41049);
nor U43140 (N_43140,N_41255,N_41208);
or U43141 (N_43141,N_41978,N_41437);
nand U43142 (N_43142,N_41576,N_40295);
or U43143 (N_43143,N_40794,N_40370);
nor U43144 (N_43144,N_41373,N_41544);
or U43145 (N_43145,N_40102,N_40279);
xor U43146 (N_43146,N_40690,N_40782);
xnor U43147 (N_43147,N_40021,N_40160);
or U43148 (N_43148,N_41951,N_41344);
nand U43149 (N_43149,N_41305,N_41286);
nand U43150 (N_43150,N_41373,N_41109);
nor U43151 (N_43151,N_40835,N_41457);
nand U43152 (N_43152,N_40432,N_41647);
and U43153 (N_43153,N_41981,N_41785);
and U43154 (N_43154,N_41317,N_41325);
xnor U43155 (N_43155,N_41540,N_40496);
or U43156 (N_43156,N_40563,N_40364);
xor U43157 (N_43157,N_40994,N_41014);
xor U43158 (N_43158,N_41543,N_41009);
nor U43159 (N_43159,N_40543,N_41097);
nor U43160 (N_43160,N_41746,N_41818);
and U43161 (N_43161,N_40761,N_40068);
and U43162 (N_43162,N_40371,N_41574);
or U43163 (N_43163,N_40602,N_40386);
nand U43164 (N_43164,N_40470,N_40542);
or U43165 (N_43165,N_40740,N_41348);
and U43166 (N_43166,N_40216,N_40517);
xor U43167 (N_43167,N_41931,N_41538);
nand U43168 (N_43168,N_41495,N_40804);
and U43169 (N_43169,N_40634,N_40154);
nand U43170 (N_43170,N_40323,N_40750);
nand U43171 (N_43171,N_41270,N_40603);
xnor U43172 (N_43172,N_40833,N_40245);
or U43173 (N_43173,N_40236,N_40525);
nand U43174 (N_43174,N_40780,N_41314);
and U43175 (N_43175,N_41906,N_40344);
nor U43176 (N_43176,N_41677,N_40768);
nand U43177 (N_43177,N_40586,N_41321);
nand U43178 (N_43178,N_40795,N_41466);
xnor U43179 (N_43179,N_40248,N_40445);
nor U43180 (N_43180,N_41420,N_41911);
and U43181 (N_43181,N_40380,N_41730);
nor U43182 (N_43182,N_40728,N_40711);
and U43183 (N_43183,N_40886,N_40481);
xor U43184 (N_43184,N_41556,N_41374);
nand U43185 (N_43185,N_41167,N_41941);
nand U43186 (N_43186,N_41202,N_40720);
xnor U43187 (N_43187,N_40946,N_40529);
nand U43188 (N_43188,N_41466,N_40522);
xor U43189 (N_43189,N_41535,N_40709);
or U43190 (N_43190,N_41437,N_41820);
nand U43191 (N_43191,N_40755,N_41748);
nand U43192 (N_43192,N_40823,N_41717);
nor U43193 (N_43193,N_40393,N_41734);
nand U43194 (N_43194,N_40960,N_40683);
xnor U43195 (N_43195,N_40116,N_41035);
and U43196 (N_43196,N_41234,N_41135);
xnor U43197 (N_43197,N_41819,N_41767);
nor U43198 (N_43198,N_40367,N_40058);
nand U43199 (N_43199,N_41207,N_40485);
xor U43200 (N_43200,N_40514,N_41367);
nand U43201 (N_43201,N_40530,N_40286);
xor U43202 (N_43202,N_40116,N_41439);
xor U43203 (N_43203,N_40057,N_40492);
or U43204 (N_43204,N_41058,N_40753);
xor U43205 (N_43205,N_41892,N_41676);
nor U43206 (N_43206,N_40932,N_40033);
and U43207 (N_43207,N_41395,N_40173);
or U43208 (N_43208,N_41956,N_40811);
nand U43209 (N_43209,N_41039,N_41350);
nor U43210 (N_43210,N_40542,N_41928);
or U43211 (N_43211,N_40414,N_40303);
or U43212 (N_43212,N_40048,N_40644);
or U43213 (N_43213,N_41465,N_40919);
nor U43214 (N_43214,N_40597,N_40337);
or U43215 (N_43215,N_41946,N_41555);
or U43216 (N_43216,N_41883,N_41681);
nand U43217 (N_43217,N_41375,N_40259);
xnor U43218 (N_43218,N_40519,N_41523);
nand U43219 (N_43219,N_41271,N_40179);
xnor U43220 (N_43220,N_40145,N_41321);
and U43221 (N_43221,N_41319,N_41222);
and U43222 (N_43222,N_41805,N_40140);
and U43223 (N_43223,N_40456,N_40788);
or U43224 (N_43224,N_41725,N_41945);
or U43225 (N_43225,N_40213,N_41955);
or U43226 (N_43226,N_40532,N_41677);
nand U43227 (N_43227,N_40788,N_40891);
xor U43228 (N_43228,N_41419,N_40401);
or U43229 (N_43229,N_40203,N_40204);
and U43230 (N_43230,N_41581,N_40107);
nor U43231 (N_43231,N_40034,N_40688);
nor U43232 (N_43232,N_40427,N_41730);
and U43233 (N_43233,N_41370,N_41145);
or U43234 (N_43234,N_40664,N_40237);
nand U43235 (N_43235,N_40902,N_41548);
nand U43236 (N_43236,N_41693,N_41310);
xnor U43237 (N_43237,N_40665,N_41123);
nor U43238 (N_43238,N_41530,N_41311);
or U43239 (N_43239,N_40293,N_41508);
nand U43240 (N_43240,N_41872,N_41070);
nand U43241 (N_43241,N_40620,N_40169);
nand U43242 (N_43242,N_41667,N_41270);
or U43243 (N_43243,N_41035,N_40098);
nand U43244 (N_43244,N_41744,N_41669);
and U43245 (N_43245,N_41340,N_41393);
or U43246 (N_43246,N_40458,N_41266);
or U43247 (N_43247,N_40444,N_40747);
xor U43248 (N_43248,N_40841,N_41698);
nand U43249 (N_43249,N_40680,N_40066);
nor U43250 (N_43250,N_40610,N_41711);
or U43251 (N_43251,N_41552,N_41109);
or U43252 (N_43252,N_41620,N_40114);
or U43253 (N_43253,N_40662,N_41707);
nor U43254 (N_43254,N_41709,N_40614);
and U43255 (N_43255,N_41063,N_40603);
and U43256 (N_43256,N_40545,N_40248);
and U43257 (N_43257,N_40266,N_40403);
xor U43258 (N_43258,N_41468,N_41520);
and U43259 (N_43259,N_40314,N_41217);
and U43260 (N_43260,N_41868,N_40080);
nor U43261 (N_43261,N_41132,N_41324);
nor U43262 (N_43262,N_40833,N_40682);
nand U43263 (N_43263,N_41451,N_41514);
xnor U43264 (N_43264,N_41811,N_40181);
or U43265 (N_43265,N_40999,N_40799);
and U43266 (N_43266,N_41608,N_40544);
or U43267 (N_43267,N_41580,N_41844);
nor U43268 (N_43268,N_40410,N_41166);
xnor U43269 (N_43269,N_41627,N_40571);
xnor U43270 (N_43270,N_40085,N_40487);
nor U43271 (N_43271,N_41713,N_40441);
or U43272 (N_43272,N_40013,N_40699);
nand U43273 (N_43273,N_40300,N_40800);
xnor U43274 (N_43274,N_40179,N_40644);
nor U43275 (N_43275,N_41905,N_40258);
nor U43276 (N_43276,N_41072,N_41809);
xor U43277 (N_43277,N_40421,N_40448);
or U43278 (N_43278,N_40439,N_41053);
or U43279 (N_43279,N_41067,N_41114);
nor U43280 (N_43280,N_41798,N_40935);
nand U43281 (N_43281,N_41980,N_40195);
or U43282 (N_43282,N_41178,N_40356);
nand U43283 (N_43283,N_41823,N_40262);
xnor U43284 (N_43284,N_41508,N_40015);
or U43285 (N_43285,N_41019,N_40525);
and U43286 (N_43286,N_40631,N_41499);
xnor U43287 (N_43287,N_40148,N_41540);
nand U43288 (N_43288,N_40196,N_41195);
nand U43289 (N_43289,N_41262,N_41508);
xnor U43290 (N_43290,N_40920,N_40335);
nor U43291 (N_43291,N_41181,N_40458);
or U43292 (N_43292,N_41185,N_41348);
nor U43293 (N_43293,N_40836,N_41035);
or U43294 (N_43294,N_41039,N_40716);
and U43295 (N_43295,N_41134,N_40070);
nand U43296 (N_43296,N_40775,N_41545);
and U43297 (N_43297,N_41229,N_40100);
nor U43298 (N_43298,N_41463,N_40071);
and U43299 (N_43299,N_40902,N_40358);
nor U43300 (N_43300,N_40516,N_41489);
nor U43301 (N_43301,N_40114,N_41880);
and U43302 (N_43302,N_40011,N_41801);
and U43303 (N_43303,N_41966,N_41000);
and U43304 (N_43304,N_41354,N_41811);
and U43305 (N_43305,N_40618,N_40621);
and U43306 (N_43306,N_40384,N_40642);
xnor U43307 (N_43307,N_40202,N_40208);
nand U43308 (N_43308,N_40199,N_40477);
nor U43309 (N_43309,N_41490,N_41311);
xnor U43310 (N_43310,N_41451,N_40435);
or U43311 (N_43311,N_41630,N_41024);
xnor U43312 (N_43312,N_40980,N_40397);
or U43313 (N_43313,N_41206,N_40311);
nand U43314 (N_43314,N_40844,N_40386);
or U43315 (N_43315,N_41978,N_40434);
xor U43316 (N_43316,N_40923,N_40261);
or U43317 (N_43317,N_40659,N_41635);
xor U43318 (N_43318,N_40863,N_41196);
nor U43319 (N_43319,N_41016,N_41316);
or U43320 (N_43320,N_41765,N_40602);
nand U43321 (N_43321,N_41650,N_41970);
nand U43322 (N_43322,N_40128,N_41412);
or U43323 (N_43323,N_41750,N_41499);
or U43324 (N_43324,N_40804,N_40244);
nor U43325 (N_43325,N_41362,N_40843);
or U43326 (N_43326,N_41678,N_40783);
xor U43327 (N_43327,N_41891,N_41768);
or U43328 (N_43328,N_41529,N_41349);
or U43329 (N_43329,N_40376,N_41284);
nand U43330 (N_43330,N_40101,N_41925);
nand U43331 (N_43331,N_41039,N_41826);
xor U43332 (N_43332,N_40496,N_40921);
nand U43333 (N_43333,N_40500,N_41750);
or U43334 (N_43334,N_40419,N_41717);
and U43335 (N_43335,N_41899,N_41314);
xnor U43336 (N_43336,N_41195,N_41101);
or U43337 (N_43337,N_41640,N_41470);
nor U43338 (N_43338,N_40317,N_41767);
nor U43339 (N_43339,N_41623,N_41017);
xor U43340 (N_43340,N_41730,N_41393);
or U43341 (N_43341,N_41133,N_41926);
nor U43342 (N_43342,N_40257,N_40702);
or U43343 (N_43343,N_41281,N_40090);
and U43344 (N_43344,N_41431,N_41478);
or U43345 (N_43345,N_40062,N_41532);
nor U43346 (N_43346,N_41706,N_41041);
and U43347 (N_43347,N_41380,N_41283);
and U43348 (N_43348,N_40331,N_40396);
xnor U43349 (N_43349,N_41789,N_40851);
xor U43350 (N_43350,N_41411,N_40127);
and U43351 (N_43351,N_40742,N_40014);
xor U43352 (N_43352,N_40607,N_40852);
nand U43353 (N_43353,N_41481,N_41733);
or U43354 (N_43354,N_40927,N_41711);
nand U43355 (N_43355,N_41641,N_41807);
nor U43356 (N_43356,N_41519,N_41202);
nand U43357 (N_43357,N_41995,N_40570);
nor U43358 (N_43358,N_41984,N_41735);
and U43359 (N_43359,N_41090,N_40356);
nor U43360 (N_43360,N_40816,N_40547);
nor U43361 (N_43361,N_40893,N_40112);
or U43362 (N_43362,N_41814,N_41748);
or U43363 (N_43363,N_40229,N_41950);
nor U43364 (N_43364,N_41007,N_41691);
nor U43365 (N_43365,N_41179,N_40977);
xor U43366 (N_43366,N_40161,N_41594);
or U43367 (N_43367,N_41230,N_41843);
xnor U43368 (N_43368,N_41856,N_40905);
xor U43369 (N_43369,N_41065,N_41846);
and U43370 (N_43370,N_40612,N_41361);
nand U43371 (N_43371,N_41161,N_41120);
nor U43372 (N_43372,N_40403,N_41037);
xnor U43373 (N_43373,N_40153,N_40309);
and U43374 (N_43374,N_40083,N_41198);
nand U43375 (N_43375,N_40695,N_41030);
nor U43376 (N_43376,N_41360,N_41226);
nor U43377 (N_43377,N_40885,N_40105);
and U43378 (N_43378,N_40230,N_41017);
and U43379 (N_43379,N_40123,N_41796);
nor U43380 (N_43380,N_40338,N_40382);
nand U43381 (N_43381,N_40971,N_40120);
xnor U43382 (N_43382,N_41821,N_41358);
nor U43383 (N_43383,N_41137,N_40432);
and U43384 (N_43384,N_41496,N_40868);
nand U43385 (N_43385,N_40464,N_40895);
xnor U43386 (N_43386,N_40788,N_40835);
nand U43387 (N_43387,N_41837,N_40386);
nor U43388 (N_43388,N_41210,N_40971);
and U43389 (N_43389,N_41442,N_41934);
xnor U43390 (N_43390,N_40267,N_41132);
and U43391 (N_43391,N_40858,N_41225);
nor U43392 (N_43392,N_40888,N_40588);
or U43393 (N_43393,N_41315,N_40288);
or U43394 (N_43394,N_40286,N_41130);
xor U43395 (N_43395,N_41017,N_40203);
and U43396 (N_43396,N_40127,N_41080);
xor U43397 (N_43397,N_40552,N_41121);
nand U43398 (N_43398,N_40229,N_41022);
nand U43399 (N_43399,N_41888,N_41330);
nand U43400 (N_43400,N_40746,N_41257);
nand U43401 (N_43401,N_40417,N_40387);
xnor U43402 (N_43402,N_41385,N_40673);
and U43403 (N_43403,N_41468,N_40535);
nand U43404 (N_43404,N_41254,N_41421);
nor U43405 (N_43405,N_40560,N_41769);
nand U43406 (N_43406,N_41825,N_40362);
or U43407 (N_43407,N_41638,N_41144);
and U43408 (N_43408,N_40962,N_41509);
or U43409 (N_43409,N_40240,N_40435);
nand U43410 (N_43410,N_41215,N_41089);
or U43411 (N_43411,N_41733,N_41594);
xor U43412 (N_43412,N_40092,N_40787);
xor U43413 (N_43413,N_40455,N_40500);
xnor U43414 (N_43414,N_40992,N_40244);
and U43415 (N_43415,N_40371,N_40842);
or U43416 (N_43416,N_41979,N_40891);
and U43417 (N_43417,N_40148,N_40344);
nand U43418 (N_43418,N_41439,N_40432);
nor U43419 (N_43419,N_41644,N_40129);
nor U43420 (N_43420,N_41947,N_40670);
nor U43421 (N_43421,N_41497,N_40951);
or U43422 (N_43422,N_41496,N_40638);
or U43423 (N_43423,N_40017,N_40783);
xor U43424 (N_43424,N_41196,N_41814);
nor U43425 (N_43425,N_41344,N_41716);
nand U43426 (N_43426,N_40533,N_40218);
nand U43427 (N_43427,N_40813,N_40828);
xnor U43428 (N_43428,N_40096,N_41382);
nor U43429 (N_43429,N_40963,N_41118);
or U43430 (N_43430,N_41094,N_41896);
xor U43431 (N_43431,N_41227,N_41151);
xor U43432 (N_43432,N_40505,N_41470);
nor U43433 (N_43433,N_41669,N_41183);
nor U43434 (N_43434,N_41815,N_40680);
nor U43435 (N_43435,N_40834,N_40120);
and U43436 (N_43436,N_40859,N_40132);
nand U43437 (N_43437,N_40769,N_41641);
or U43438 (N_43438,N_41577,N_41609);
xnor U43439 (N_43439,N_40711,N_41679);
or U43440 (N_43440,N_40595,N_40404);
and U43441 (N_43441,N_40999,N_40098);
or U43442 (N_43442,N_40529,N_41695);
nor U43443 (N_43443,N_41122,N_40469);
nor U43444 (N_43444,N_40753,N_41792);
nor U43445 (N_43445,N_41038,N_40715);
nor U43446 (N_43446,N_41440,N_41983);
nand U43447 (N_43447,N_41094,N_40533);
nand U43448 (N_43448,N_41152,N_41434);
or U43449 (N_43449,N_40493,N_41609);
xnor U43450 (N_43450,N_41634,N_40500);
and U43451 (N_43451,N_41331,N_41267);
xor U43452 (N_43452,N_40304,N_40724);
xnor U43453 (N_43453,N_41255,N_41322);
xor U43454 (N_43454,N_41392,N_40159);
nor U43455 (N_43455,N_40568,N_41586);
xnor U43456 (N_43456,N_40982,N_41262);
xor U43457 (N_43457,N_40487,N_40143);
and U43458 (N_43458,N_41590,N_40352);
xnor U43459 (N_43459,N_41772,N_40921);
nor U43460 (N_43460,N_40386,N_41780);
or U43461 (N_43461,N_40155,N_41476);
and U43462 (N_43462,N_40558,N_41251);
nand U43463 (N_43463,N_40373,N_40015);
nand U43464 (N_43464,N_40805,N_40404);
nor U43465 (N_43465,N_41783,N_40813);
nand U43466 (N_43466,N_41956,N_40501);
xnor U43467 (N_43467,N_40734,N_40117);
or U43468 (N_43468,N_41844,N_40989);
xor U43469 (N_43469,N_40285,N_41784);
nand U43470 (N_43470,N_40990,N_41687);
xnor U43471 (N_43471,N_40289,N_41292);
nand U43472 (N_43472,N_40329,N_41773);
or U43473 (N_43473,N_40209,N_41918);
and U43474 (N_43474,N_41072,N_41730);
xor U43475 (N_43475,N_41447,N_41914);
nor U43476 (N_43476,N_40445,N_41166);
xnor U43477 (N_43477,N_41946,N_40322);
and U43478 (N_43478,N_40632,N_41982);
xnor U43479 (N_43479,N_40230,N_41996);
and U43480 (N_43480,N_41495,N_41744);
nor U43481 (N_43481,N_41821,N_41732);
nor U43482 (N_43482,N_41821,N_40175);
xor U43483 (N_43483,N_40908,N_41563);
or U43484 (N_43484,N_41391,N_41683);
nor U43485 (N_43485,N_40763,N_40258);
or U43486 (N_43486,N_41332,N_40360);
or U43487 (N_43487,N_41155,N_40004);
or U43488 (N_43488,N_40979,N_40863);
nor U43489 (N_43489,N_40945,N_40053);
nor U43490 (N_43490,N_40713,N_40417);
and U43491 (N_43491,N_40611,N_41861);
nand U43492 (N_43492,N_41768,N_40430);
xor U43493 (N_43493,N_40652,N_40619);
and U43494 (N_43494,N_40011,N_41744);
and U43495 (N_43495,N_40078,N_41282);
nand U43496 (N_43496,N_40075,N_41171);
nand U43497 (N_43497,N_40891,N_40652);
or U43498 (N_43498,N_40269,N_40802);
and U43499 (N_43499,N_41250,N_40590);
nor U43500 (N_43500,N_41428,N_40244);
xor U43501 (N_43501,N_41664,N_40838);
nand U43502 (N_43502,N_40787,N_41751);
or U43503 (N_43503,N_41985,N_40027);
xnor U43504 (N_43504,N_41948,N_41809);
or U43505 (N_43505,N_40387,N_41094);
or U43506 (N_43506,N_41293,N_40198);
nor U43507 (N_43507,N_40592,N_41352);
nor U43508 (N_43508,N_41783,N_40687);
or U43509 (N_43509,N_40578,N_40766);
or U43510 (N_43510,N_41600,N_40712);
nor U43511 (N_43511,N_40332,N_41260);
and U43512 (N_43512,N_40074,N_41461);
and U43513 (N_43513,N_41288,N_40470);
and U43514 (N_43514,N_40570,N_40195);
nor U43515 (N_43515,N_40078,N_40267);
xnor U43516 (N_43516,N_40338,N_40546);
nand U43517 (N_43517,N_41336,N_40186);
xnor U43518 (N_43518,N_40781,N_41277);
nand U43519 (N_43519,N_40392,N_41848);
or U43520 (N_43520,N_40849,N_40570);
xor U43521 (N_43521,N_40513,N_41810);
nor U43522 (N_43522,N_40882,N_41850);
nor U43523 (N_43523,N_41933,N_41226);
or U43524 (N_43524,N_40773,N_40983);
or U43525 (N_43525,N_41440,N_41539);
and U43526 (N_43526,N_41188,N_40635);
or U43527 (N_43527,N_40052,N_40677);
nand U43528 (N_43528,N_40417,N_40401);
xor U43529 (N_43529,N_40619,N_40337);
nor U43530 (N_43530,N_41893,N_41480);
nor U43531 (N_43531,N_41669,N_40344);
or U43532 (N_43532,N_41212,N_40167);
nand U43533 (N_43533,N_41077,N_40678);
and U43534 (N_43534,N_41025,N_40305);
xor U43535 (N_43535,N_40588,N_41261);
nand U43536 (N_43536,N_41706,N_40377);
xnor U43537 (N_43537,N_40524,N_40127);
xor U43538 (N_43538,N_41553,N_41082);
nand U43539 (N_43539,N_41935,N_40492);
nand U43540 (N_43540,N_41003,N_41970);
and U43541 (N_43541,N_41863,N_41315);
nand U43542 (N_43542,N_40488,N_40549);
or U43543 (N_43543,N_41405,N_41818);
and U43544 (N_43544,N_41961,N_41342);
xor U43545 (N_43545,N_40537,N_40281);
and U43546 (N_43546,N_40258,N_41882);
nand U43547 (N_43547,N_41007,N_41484);
nand U43548 (N_43548,N_40679,N_40073);
and U43549 (N_43549,N_41307,N_40771);
and U43550 (N_43550,N_40577,N_41848);
and U43551 (N_43551,N_41320,N_41239);
nor U43552 (N_43552,N_41447,N_40003);
or U43553 (N_43553,N_40915,N_40798);
xnor U43554 (N_43554,N_40817,N_41381);
nand U43555 (N_43555,N_40724,N_41754);
and U43556 (N_43556,N_40332,N_41650);
nand U43557 (N_43557,N_41109,N_40062);
xor U43558 (N_43558,N_41915,N_41276);
nand U43559 (N_43559,N_40288,N_41133);
xnor U43560 (N_43560,N_41987,N_41816);
xnor U43561 (N_43561,N_40583,N_41652);
nor U43562 (N_43562,N_41707,N_40283);
nor U43563 (N_43563,N_40412,N_41199);
or U43564 (N_43564,N_40388,N_41632);
nand U43565 (N_43565,N_41238,N_41222);
nand U43566 (N_43566,N_41652,N_40434);
and U43567 (N_43567,N_41580,N_41266);
or U43568 (N_43568,N_41838,N_40574);
nand U43569 (N_43569,N_41051,N_41790);
or U43570 (N_43570,N_41300,N_40108);
or U43571 (N_43571,N_40611,N_40239);
nand U43572 (N_43572,N_40185,N_40522);
xnor U43573 (N_43573,N_40315,N_41194);
or U43574 (N_43574,N_41786,N_41401);
nor U43575 (N_43575,N_40860,N_41979);
nor U43576 (N_43576,N_41179,N_41467);
and U43577 (N_43577,N_41582,N_40233);
xor U43578 (N_43578,N_40008,N_40489);
nor U43579 (N_43579,N_40622,N_40280);
nor U43580 (N_43580,N_41582,N_40948);
and U43581 (N_43581,N_40574,N_41842);
nand U43582 (N_43582,N_41713,N_40455);
or U43583 (N_43583,N_41376,N_40414);
nor U43584 (N_43584,N_41238,N_40363);
or U43585 (N_43585,N_41504,N_41934);
and U43586 (N_43586,N_40538,N_41778);
and U43587 (N_43587,N_40527,N_40032);
nor U43588 (N_43588,N_40836,N_41373);
xnor U43589 (N_43589,N_41839,N_40504);
nor U43590 (N_43590,N_41323,N_41869);
and U43591 (N_43591,N_40299,N_41215);
nand U43592 (N_43592,N_40727,N_41036);
or U43593 (N_43593,N_40616,N_41842);
and U43594 (N_43594,N_40829,N_40974);
or U43595 (N_43595,N_40204,N_41470);
xor U43596 (N_43596,N_40082,N_41341);
nor U43597 (N_43597,N_41411,N_41821);
nand U43598 (N_43598,N_40917,N_40082);
nand U43599 (N_43599,N_41422,N_40321);
xnor U43600 (N_43600,N_40845,N_40549);
or U43601 (N_43601,N_40832,N_40836);
and U43602 (N_43602,N_41202,N_40911);
xor U43603 (N_43603,N_40749,N_41419);
and U43604 (N_43604,N_40629,N_40524);
and U43605 (N_43605,N_41591,N_40036);
nand U43606 (N_43606,N_41959,N_41459);
and U43607 (N_43607,N_40552,N_41211);
nor U43608 (N_43608,N_41171,N_41220);
and U43609 (N_43609,N_41537,N_41248);
nor U43610 (N_43610,N_40424,N_40026);
nor U43611 (N_43611,N_41423,N_40772);
nor U43612 (N_43612,N_40894,N_41003);
xor U43613 (N_43613,N_40450,N_40628);
or U43614 (N_43614,N_40653,N_40132);
nor U43615 (N_43615,N_40931,N_40146);
or U43616 (N_43616,N_40711,N_40099);
nor U43617 (N_43617,N_41470,N_41261);
nand U43618 (N_43618,N_41001,N_40739);
or U43619 (N_43619,N_41678,N_41021);
nand U43620 (N_43620,N_41491,N_40445);
nand U43621 (N_43621,N_41395,N_41229);
nand U43622 (N_43622,N_41745,N_41148);
and U43623 (N_43623,N_40489,N_40765);
nor U43624 (N_43624,N_41173,N_40650);
nor U43625 (N_43625,N_41866,N_40680);
or U43626 (N_43626,N_41293,N_40372);
or U43627 (N_43627,N_40681,N_40237);
nand U43628 (N_43628,N_40237,N_41717);
or U43629 (N_43629,N_41993,N_41798);
nand U43630 (N_43630,N_40031,N_40943);
and U43631 (N_43631,N_41689,N_41913);
and U43632 (N_43632,N_41842,N_41348);
nor U43633 (N_43633,N_41298,N_41748);
nor U43634 (N_43634,N_40643,N_40544);
xor U43635 (N_43635,N_41354,N_40163);
nand U43636 (N_43636,N_41416,N_40751);
nor U43637 (N_43637,N_40130,N_40906);
and U43638 (N_43638,N_41010,N_40883);
nand U43639 (N_43639,N_40590,N_41466);
nand U43640 (N_43640,N_40561,N_40190);
xor U43641 (N_43641,N_41274,N_40291);
xor U43642 (N_43642,N_41043,N_41704);
nand U43643 (N_43643,N_41731,N_41175);
nand U43644 (N_43644,N_41805,N_40778);
nor U43645 (N_43645,N_40938,N_41395);
and U43646 (N_43646,N_41841,N_40031);
nand U43647 (N_43647,N_41545,N_40474);
xnor U43648 (N_43648,N_41229,N_40024);
nand U43649 (N_43649,N_41502,N_41169);
or U43650 (N_43650,N_41007,N_41950);
or U43651 (N_43651,N_41163,N_40802);
nand U43652 (N_43652,N_40335,N_41637);
xnor U43653 (N_43653,N_40971,N_40374);
and U43654 (N_43654,N_41452,N_40902);
nor U43655 (N_43655,N_41637,N_41118);
nand U43656 (N_43656,N_41625,N_40595);
and U43657 (N_43657,N_40148,N_41287);
nand U43658 (N_43658,N_40089,N_41594);
xnor U43659 (N_43659,N_41040,N_41722);
and U43660 (N_43660,N_40979,N_40500);
xor U43661 (N_43661,N_41561,N_40881);
and U43662 (N_43662,N_40282,N_41705);
nor U43663 (N_43663,N_41471,N_40352);
nor U43664 (N_43664,N_40429,N_40409);
and U43665 (N_43665,N_40576,N_41962);
nor U43666 (N_43666,N_41669,N_41055);
xnor U43667 (N_43667,N_40511,N_41202);
and U43668 (N_43668,N_41111,N_41290);
nand U43669 (N_43669,N_41323,N_41129);
or U43670 (N_43670,N_40255,N_40071);
or U43671 (N_43671,N_40715,N_41270);
nor U43672 (N_43672,N_41831,N_40524);
nor U43673 (N_43673,N_40856,N_40508);
and U43674 (N_43674,N_41489,N_41348);
nor U43675 (N_43675,N_41788,N_41952);
xnor U43676 (N_43676,N_41636,N_41104);
nand U43677 (N_43677,N_41759,N_40701);
or U43678 (N_43678,N_41709,N_41926);
and U43679 (N_43679,N_41805,N_41233);
nor U43680 (N_43680,N_40953,N_41769);
xor U43681 (N_43681,N_41426,N_41989);
xnor U43682 (N_43682,N_41966,N_41124);
xnor U43683 (N_43683,N_41798,N_41766);
xor U43684 (N_43684,N_41495,N_41555);
xor U43685 (N_43685,N_41477,N_40639);
nand U43686 (N_43686,N_40556,N_41611);
nor U43687 (N_43687,N_41736,N_41176);
xor U43688 (N_43688,N_41254,N_40704);
or U43689 (N_43689,N_41993,N_40291);
nand U43690 (N_43690,N_41271,N_40330);
nor U43691 (N_43691,N_40739,N_41784);
or U43692 (N_43692,N_40797,N_40481);
or U43693 (N_43693,N_41103,N_40437);
xnor U43694 (N_43694,N_41419,N_41554);
nand U43695 (N_43695,N_41448,N_41230);
xnor U43696 (N_43696,N_41805,N_40656);
nand U43697 (N_43697,N_40017,N_41051);
xor U43698 (N_43698,N_41339,N_41528);
nor U43699 (N_43699,N_41655,N_41425);
xor U43700 (N_43700,N_41444,N_41075);
nand U43701 (N_43701,N_41622,N_41841);
nand U43702 (N_43702,N_41067,N_41671);
xor U43703 (N_43703,N_40457,N_41560);
xor U43704 (N_43704,N_40797,N_40142);
or U43705 (N_43705,N_41193,N_40991);
and U43706 (N_43706,N_40873,N_40953);
or U43707 (N_43707,N_41835,N_41328);
or U43708 (N_43708,N_40707,N_40360);
nor U43709 (N_43709,N_41794,N_41682);
nor U43710 (N_43710,N_41171,N_41257);
and U43711 (N_43711,N_40689,N_40532);
nor U43712 (N_43712,N_41895,N_40204);
or U43713 (N_43713,N_40920,N_41104);
nor U43714 (N_43714,N_40417,N_41922);
xnor U43715 (N_43715,N_41239,N_40541);
and U43716 (N_43716,N_40051,N_40013);
nor U43717 (N_43717,N_41781,N_40649);
or U43718 (N_43718,N_41732,N_40638);
xnor U43719 (N_43719,N_40074,N_41770);
nand U43720 (N_43720,N_40658,N_41194);
xor U43721 (N_43721,N_40656,N_41029);
or U43722 (N_43722,N_41810,N_40408);
nand U43723 (N_43723,N_40947,N_41120);
or U43724 (N_43724,N_40936,N_41234);
and U43725 (N_43725,N_41014,N_41117);
xnor U43726 (N_43726,N_40642,N_41857);
or U43727 (N_43727,N_40865,N_41106);
nor U43728 (N_43728,N_40320,N_40122);
xnor U43729 (N_43729,N_41126,N_41857);
nor U43730 (N_43730,N_40855,N_41406);
nand U43731 (N_43731,N_41509,N_41093);
nor U43732 (N_43732,N_41672,N_41055);
and U43733 (N_43733,N_40510,N_40800);
xnor U43734 (N_43734,N_41091,N_41460);
nand U43735 (N_43735,N_40981,N_40920);
and U43736 (N_43736,N_40494,N_40093);
or U43737 (N_43737,N_41442,N_40654);
xnor U43738 (N_43738,N_40099,N_41308);
or U43739 (N_43739,N_41741,N_41402);
nand U43740 (N_43740,N_41107,N_41971);
and U43741 (N_43741,N_41224,N_40777);
nor U43742 (N_43742,N_41436,N_41600);
nand U43743 (N_43743,N_41188,N_41876);
and U43744 (N_43744,N_40000,N_41490);
nand U43745 (N_43745,N_40134,N_40885);
nor U43746 (N_43746,N_41176,N_41979);
nor U43747 (N_43747,N_41295,N_41317);
or U43748 (N_43748,N_41998,N_41810);
xnor U43749 (N_43749,N_40934,N_41347);
and U43750 (N_43750,N_41021,N_40275);
or U43751 (N_43751,N_40397,N_41852);
and U43752 (N_43752,N_40044,N_41410);
xnor U43753 (N_43753,N_41153,N_41956);
nand U43754 (N_43754,N_41213,N_41543);
and U43755 (N_43755,N_40979,N_41862);
or U43756 (N_43756,N_41923,N_40446);
nand U43757 (N_43757,N_41056,N_41325);
nor U43758 (N_43758,N_40292,N_41697);
xor U43759 (N_43759,N_41419,N_41724);
xnor U43760 (N_43760,N_40248,N_40192);
and U43761 (N_43761,N_40722,N_40017);
xnor U43762 (N_43762,N_40180,N_40649);
xnor U43763 (N_43763,N_40041,N_41534);
nor U43764 (N_43764,N_40118,N_40097);
nand U43765 (N_43765,N_40330,N_40190);
xor U43766 (N_43766,N_41780,N_41788);
xor U43767 (N_43767,N_41465,N_40500);
and U43768 (N_43768,N_41148,N_41452);
or U43769 (N_43769,N_41278,N_41496);
and U43770 (N_43770,N_41530,N_40537);
and U43771 (N_43771,N_40527,N_40479);
xor U43772 (N_43772,N_41781,N_40089);
xnor U43773 (N_43773,N_40956,N_40857);
and U43774 (N_43774,N_40695,N_40605);
nand U43775 (N_43775,N_40025,N_40073);
nor U43776 (N_43776,N_40631,N_41876);
nand U43777 (N_43777,N_41844,N_40056);
and U43778 (N_43778,N_40533,N_40002);
xnor U43779 (N_43779,N_40944,N_40141);
nand U43780 (N_43780,N_40702,N_40258);
and U43781 (N_43781,N_41104,N_41423);
nand U43782 (N_43782,N_41594,N_40138);
nand U43783 (N_43783,N_41245,N_41147);
and U43784 (N_43784,N_41110,N_40410);
xnor U43785 (N_43785,N_41171,N_41450);
or U43786 (N_43786,N_40203,N_40642);
or U43787 (N_43787,N_40441,N_41533);
or U43788 (N_43788,N_41469,N_40137);
nand U43789 (N_43789,N_40752,N_41203);
xor U43790 (N_43790,N_41714,N_41280);
and U43791 (N_43791,N_40321,N_40742);
nor U43792 (N_43792,N_40072,N_40320);
nor U43793 (N_43793,N_41824,N_40079);
and U43794 (N_43794,N_40593,N_41405);
nand U43795 (N_43795,N_41292,N_40456);
nand U43796 (N_43796,N_40961,N_41672);
and U43797 (N_43797,N_40933,N_41446);
xor U43798 (N_43798,N_40407,N_41008);
xnor U43799 (N_43799,N_40023,N_41900);
nor U43800 (N_43800,N_40089,N_41337);
or U43801 (N_43801,N_41435,N_40362);
nor U43802 (N_43802,N_40815,N_41765);
nor U43803 (N_43803,N_41876,N_40094);
or U43804 (N_43804,N_40235,N_41589);
nor U43805 (N_43805,N_40879,N_40697);
nor U43806 (N_43806,N_40297,N_41607);
xnor U43807 (N_43807,N_40857,N_40426);
and U43808 (N_43808,N_40273,N_40931);
nand U43809 (N_43809,N_41246,N_41970);
xor U43810 (N_43810,N_41528,N_41929);
or U43811 (N_43811,N_41981,N_41545);
xnor U43812 (N_43812,N_41331,N_40615);
nand U43813 (N_43813,N_40437,N_41322);
and U43814 (N_43814,N_41222,N_41507);
nand U43815 (N_43815,N_41552,N_40455);
nor U43816 (N_43816,N_40815,N_40693);
or U43817 (N_43817,N_40910,N_40736);
nor U43818 (N_43818,N_41164,N_40567);
nand U43819 (N_43819,N_40960,N_40355);
and U43820 (N_43820,N_40598,N_41967);
and U43821 (N_43821,N_41785,N_41532);
and U43822 (N_43822,N_40770,N_41556);
xor U43823 (N_43823,N_40357,N_41479);
nand U43824 (N_43824,N_41905,N_41073);
nor U43825 (N_43825,N_41198,N_40416);
or U43826 (N_43826,N_40689,N_41361);
and U43827 (N_43827,N_41866,N_40225);
nand U43828 (N_43828,N_41729,N_40518);
nand U43829 (N_43829,N_40938,N_41287);
and U43830 (N_43830,N_40716,N_41341);
xnor U43831 (N_43831,N_41133,N_41972);
or U43832 (N_43832,N_41603,N_40411);
xnor U43833 (N_43833,N_41075,N_40510);
or U43834 (N_43834,N_41466,N_40281);
and U43835 (N_43835,N_40047,N_41170);
nor U43836 (N_43836,N_41790,N_41218);
or U43837 (N_43837,N_40584,N_40751);
nand U43838 (N_43838,N_40700,N_41928);
or U43839 (N_43839,N_41072,N_41922);
nand U43840 (N_43840,N_40204,N_40634);
nand U43841 (N_43841,N_40328,N_41329);
xor U43842 (N_43842,N_40584,N_40314);
nand U43843 (N_43843,N_40986,N_41416);
nand U43844 (N_43844,N_40390,N_40425);
nor U43845 (N_43845,N_41293,N_40052);
xor U43846 (N_43846,N_40131,N_40717);
nor U43847 (N_43847,N_40352,N_40489);
nand U43848 (N_43848,N_41191,N_40183);
xor U43849 (N_43849,N_40628,N_41119);
or U43850 (N_43850,N_41260,N_41728);
nand U43851 (N_43851,N_40512,N_41995);
and U43852 (N_43852,N_41525,N_40835);
nand U43853 (N_43853,N_41347,N_41813);
nor U43854 (N_43854,N_40555,N_41524);
nand U43855 (N_43855,N_41604,N_40996);
nor U43856 (N_43856,N_40740,N_40458);
nor U43857 (N_43857,N_40545,N_40554);
and U43858 (N_43858,N_40286,N_40576);
or U43859 (N_43859,N_40925,N_40673);
and U43860 (N_43860,N_40332,N_41343);
nor U43861 (N_43861,N_40380,N_41324);
nand U43862 (N_43862,N_40083,N_40692);
nand U43863 (N_43863,N_41396,N_41064);
xnor U43864 (N_43864,N_40753,N_41555);
nor U43865 (N_43865,N_41298,N_41391);
xnor U43866 (N_43866,N_41760,N_41051);
nor U43867 (N_43867,N_40494,N_40346);
or U43868 (N_43868,N_41036,N_41692);
nand U43869 (N_43869,N_40647,N_40577);
xnor U43870 (N_43870,N_41128,N_40322);
nand U43871 (N_43871,N_40203,N_40680);
and U43872 (N_43872,N_40926,N_41167);
and U43873 (N_43873,N_41281,N_41830);
xor U43874 (N_43874,N_41976,N_40518);
and U43875 (N_43875,N_40673,N_41506);
or U43876 (N_43876,N_40217,N_40119);
nor U43877 (N_43877,N_41973,N_41693);
nor U43878 (N_43878,N_40183,N_40488);
or U43879 (N_43879,N_41740,N_40810);
xnor U43880 (N_43880,N_40263,N_41610);
nor U43881 (N_43881,N_40713,N_41962);
and U43882 (N_43882,N_41177,N_41268);
and U43883 (N_43883,N_40420,N_40030);
or U43884 (N_43884,N_41813,N_40187);
or U43885 (N_43885,N_40301,N_41918);
nand U43886 (N_43886,N_41160,N_40053);
xnor U43887 (N_43887,N_41668,N_41287);
xnor U43888 (N_43888,N_41497,N_41684);
and U43889 (N_43889,N_40648,N_41679);
or U43890 (N_43890,N_41167,N_40334);
nor U43891 (N_43891,N_40001,N_41654);
nor U43892 (N_43892,N_41013,N_41121);
nor U43893 (N_43893,N_40829,N_41355);
xor U43894 (N_43894,N_40861,N_41794);
and U43895 (N_43895,N_41754,N_40476);
or U43896 (N_43896,N_41552,N_40565);
and U43897 (N_43897,N_41166,N_41849);
nor U43898 (N_43898,N_40853,N_41542);
nand U43899 (N_43899,N_41855,N_40026);
or U43900 (N_43900,N_41959,N_41501);
nand U43901 (N_43901,N_40368,N_40083);
nor U43902 (N_43902,N_41702,N_41055);
and U43903 (N_43903,N_41427,N_40739);
xor U43904 (N_43904,N_41605,N_41472);
or U43905 (N_43905,N_41922,N_40230);
nand U43906 (N_43906,N_41608,N_40329);
xnor U43907 (N_43907,N_40507,N_40183);
xor U43908 (N_43908,N_40128,N_40673);
nand U43909 (N_43909,N_40778,N_40272);
or U43910 (N_43910,N_41269,N_40043);
xnor U43911 (N_43911,N_40712,N_40261);
nor U43912 (N_43912,N_40817,N_40497);
nand U43913 (N_43913,N_40095,N_40144);
nand U43914 (N_43914,N_40201,N_40512);
or U43915 (N_43915,N_41208,N_40839);
or U43916 (N_43916,N_40683,N_41722);
nor U43917 (N_43917,N_41694,N_40816);
or U43918 (N_43918,N_41269,N_40019);
and U43919 (N_43919,N_40546,N_40912);
xnor U43920 (N_43920,N_40744,N_41866);
nand U43921 (N_43921,N_41238,N_40481);
nand U43922 (N_43922,N_40960,N_41674);
or U43923 (N_43923,N_41281,N_41420);
or U43924 (N_43924,N_41158,N_40954);
and U43925 (N_43925,N_41111,N_41380);
or U43926 (N_43926,N_40777,N_41029);
and U43927 (N_43927,N_40336,N_40756);
and U43928 (N_43928,N_41857,N_41540);
xor U43929 (N_43929,N_40100,N_41727);
nor U43930 (N_43930,N_40557,N_41509);
nand U43931 (N_43931,N_40297,N_40240);
nor U43932 (N_43932,N_41858,N_40932);
nand U43933 (N_43933,N_41479,N_40078);
and U43934 (N_43934,N_40441,N_41100);
nor U43935 (N_43935,N_40506,N_40025);
or U43936 (N_43936,N_40542,N_40638);
xor U43937 (N_43937,N_41689,N_41777);
nand U43938 (N_43938,N_41523,N_40999);
or U43939 (N_43939,N_41676,N_40289);
xnor U43940 (N_43940,N_41056,N_41924);
nand U43941 (N_43941,N_41311,N_40588);
nand U43942 (N_43942,N_40217,N_41104);
or U43943 (N_43943,N_41194,N_40075);
or U43944 (N_43944,N_41237,N_41880);
xnor U43945 (N_43945,N_41286,N_40892);
xor U43946 (N_43946,N_41617,N_40570);
nor U43947 (N_43947,N_40193,N_41067);
xor U43948 (N_43948,N_40054,N_41472);
nand U43949 (N_43949,N_40509,N_41616);
or U43950 (N_43950,N_41194,N_41736);
nor U43951 (N_43951,N_40057,N_41946);
and U43952 (N_43952,N_41752,N_41093);
nand U43953 (N_43953,N_40728,N_40765);
or U43954 (N_43954,N_40088,N_40073);
and U43955 (N_43955,N_40624,N_40137);
xnor U43956 (N_43956,N_40911,N_41673);
or U43957 (N_43957,N_40440,N_40523);
or U43958 (N_43958,N_40879,N_41400);
and U43959 (N_43959,N_41992,N_41067);
and U43960 (N_43960,N_40595,N_40183);
nor U43961 (N_43961,N_40905,N_41666);
nor U43962 (N_43962,N_41385,N_40099);
xor U43963 (N_43963,N_41998,N_40197);
xnor U43964 (N_43964,N_41160,N_40780);
nand U43965 (N_43965,N_41315,N_40734);
nor U43966 (N_43966,N_40471,N_40518);
xor U43967 (N_43967,N_41996,N_41101);
nor U43968 (N_43968,N_41751,N_41161);
xnor U43969 (N_43969,N_41076,N_41768);
nand U43970 (N_43970,N_40386,N_40879);
xnor U43971 (N_43971,N_40064,N_40762);
xor U43972 (N_43972,N_40842,N_41357);
or U43973 (N_43973,N_41837,N_40564);
or U43974 (N_43974,N_40518,N_40550);
nand U43975 (N_43975,N_41862,N_40848);
nor U43976 (N_43976,N_40957,N_40545);
xor U43977 (N_43977,N_40885,N_40958);
and U43978 (N_43978,N_41259,N_41863);
and U43979 (N_43979,N_41090,N_41099);
nor U43980 (N_43980,N_40058,N_40633);
nor U43981 (N_43981,N_41408,N_41095);
or U43982 (N_43982,N_41000,N_40482);
or U43983 (N_43983,N_40847,N_41868);
xor U43984 (N_43984,N_41810,N_40941);
nor U43985 (N_43985,N_40876,N_40501);
or U43986 (N_43986,N_40359,N_41733);
xnor U43987 (N_43987,N_41513,N_41039);
nor U43988 (N_43988,N_40369,N_40675);
or U43989 (N_43989,N_40697,N_41829);
and U43990 (N_43990,N_41906,N_41151);
xnor U43991 (N_43991,N_40927,N_41116);
and U43992 (N_43992,N_41846,N_41683);
and U43993 (N_43993,N_41628,N_40874);
and U43994 (N_43994,N_40493,N_41089);
and U43995 (N_43995,N_40233,N_41778);
nand U43996 (N_43996,N_41266,N_40633);
and U43997 (N_43997,N_40421,N_41002);
nand U43998 (N_43998,N_40614,N_40108);
xnor U43999 (N_43999,N_40048,N_40595);
and U44000 (N_44000,N_43794,N_43109);
xor U44001 (N_44001,N_42650,N_43746);
nor U44002 (N_44002,N_42010,N_43936);
or U44003 (N_44003,N_43185,N_43826);
nor U44004 (N_44004,N_43581,N_42320);
and U44005 (N_44005,N_43086,N_43543);
and U44006 (N_44006,N_43881,N_43623);
or U44007 (N_44007,N_43559,N_43619);
xnor U44008 (N_44008,N_42441,N_42791);
and U44009 (N_44009,N_42052,N_42272);
or U44010 (N_44010,N_42995,N_43478);
xnor U44011 (N_44011,N_42790,N_43470);
or U44012 (N_44012,N_42962,N_43073);
and U44013 (N_44013,N_42903,N_42321);
nor U44014 (N_44014,N_43747,N_42128);
nand U44015 (N_44015,N_42420,N_43588);
xnor U44016 (N_44016,N_42901,N_43615);
and U44017 (N_44017,N_42848,N_42846);
xnor U44018 (N_44018,N_42851,N_42681);
nor U44019 (N_44019,N_43359,N_42544);
or U44020 (N_44020,N_42311,N_43914);
or U44021 (N_44021,N_42286,N_42063);
xor U44022 (N_44022,N_43129,N_42364);
and U44023 (N_44023,N_42159,N_43560);
nand U44024 (N_44024,N_43864,N_42331);
and U44025 (N_44025,N_42349,N_42122);
xor U44026 (N_44026,N_43898,N_42685);
and U44027 (N_44027,N_43490,N_42862);
and U44028 (N_44028,N_42729,N_42066);
nand U44029 (N_44029,N_42202,N_42383);
xor U44030 (N_44030,N_42587,N_43203);
nand U44031 (N_44031,N_43516,N_43396);
nor U44032 (N_44032,N_42016,N_43280);
nand U44033 (N_44033,N_43110,N_43819);
and U44034 (N_44034,N_42037,N_42354);
nand U44035 (N_44035,N_42671,N_43117);
xor U44036 (N_44036,N_42188,N_43800);
xor U44037 (N_44037,N_42779,N_43392);
xnor U44038 (N_44038,N_43617,N_43944);
or U44039 (N_44039,N_43813,N_42280);
or U44040 (N_44040,N_43575,N_43756);
and U44041 (N_44041,N_43252,N_42234);
nor U44042 (N_44042,N_42812,N_43569);
nor U44043 (N_44043,N_42330,N_43026);
xnor U44044 (N_44044,N_43867,N_42160);
nand U44045 (N_44045,N_42764,N_42020);
xnor U44046 (N_44046,N_42568,N_42881);
nor U44047 (N_44047,N_42821,N_42961);
or U44048 (N_44048,N_42357,N_42071);
nand U44049 (N_44049,N_42422,N_43532);
and U44050 (N_44050,N_42703,N_42186);
nand U44051 (N_44051,N_43048,N_43178);
xor U44052 (N_44052,N_42001,N_43750);
xor U44053 (N_44053,N_43765,N_43610);
nand U44054 (N_44054,N_42336,N_42949);
nand U44055 (N_44055,N_43933,N_43691);
nor U44056 (N_44056,N_43554,N_43498);
and U44057 (N_44057,N_43266,N_42893);
and U44058 (N_44058,N_42913,N_42784);
nor U44059 (N_44059,N_42100,N_43851);
nor U44060 (N_44060,N_43449,N_42545);
or U44061 (N_44061,N_43485,N_42968);
and U44062 (N_44062,N_42528,N_42561);
and U44063 (N_44063,N_43915,N_42424);
nor U44064 (N_44064,N_42612,N_42377);
nor U44065 (N_44065,N_43150,N_42825);
nor U44066 (N_44066,N_43010,N_43297);
or U44067 (N_44067,N_42167,N_43494);
xor U44068 (N_44068,N_43477,N_42939);
nand U44069 (N_44069,N_43093,N_42363);
nand U44070 (N_44070,N_42482,N_43163);
and U44071 (N_44071,N_42566,N_42917);
nor U44072 (N_44072,N_42132,N_43320);
nor U44073 (N_44073,N_42556,N_42055);
xnor U44074 (N_44074,N_42410,N_42290);
or U44075 (N_44075,N_43698,N_43334);
xnor U44076 (N_44076,N_43500,N_42533);
xnor U44077 (N_44077,N_43351,N_42299);
nor U44078 (N_44078,N_42237,N_42476);
nor U44079 (N_44079,N_43005,N_43829);
xnor U44080 (N_44080,N_43835,N_42109);
xnor U44081 (N_44081,N_42498,N_43620);
and U44082 (N_44082,N_43285,N_42595);
xnor U44083 (N_44083,N_42250,N_43440);
xnor U44084 (N_44084,N_42008,N_43932);
nand U44085 (N_44085,N_43384,N_42976);
nor U44086 (N_44086,N_42885,N_43597);
and U44087 (N_44087,N_42666,N_42753);
nand U44088 (N_44088,N_43029,N_42627);
nor U44089 (N_44089,N_42975,N_42038);
xor U44090 (N_44090,N_42600,N_42499);
nand U44091 (N_44091,N_43357,N_42850);
or U44092 (N_44092,N_43790,N_42376);
and U44093 (N_44093,N_43966,N_42573);
nand U44094 (N_44094,N_42054,N_43792);
nor U44095 (N_44095,N_42073,N_42553);
and U44096 (N_44096,N_43605,N_42496);
xnor U44097 (N_44097,N_43101,N_42249);
nand U44098 (N_44098,N_43999,N_43885);
nand U44099 (N_44099,N_42183,N_42447);
and U44100 (N_44100,N_43626,N_43870);
and U44101 (N_44101,N_42623,N_42657);
or U44102 (N_44102,N_43327,N_43902);
nor U44103 (N_44103,N_42242,N_43804);
or U44104 (N_44104,N_43095,N_43282);
xor U44105 (N_44105,N_43856,N_43555);
nor U44106 (N_44106,N_43279,N_43678);
or U44107 (N_44107,N_42700,N_43045);
xnor U44108 (N_44108,N_43293,N_43237);
and U44109 (N_44109,N_43793,N_42548);
or U44110 (N_44110,N_42590,N_43727);
and U44111 (N_44111,N_42271,N_42270);
and U44112 (N_44112,N_42429,N_42333);
nor U44113 (N_44113,N_42516,N_42085);
and U44114 (N_44114,N_42105,N_42187);
or U44115 (N_44115,N_42797,N_43164);
xor U44116 (N_44116,N_43680,N_42162);
and U44117 (N_44117,N_43425,N_43947);
nor U44118 (N_44118,N_43133,N_42788);
or U44119 (N_44119,N_43186,N_42839);
nand U44120 (N_44120,N_42506,N_43833);
or U44121 (N_44121,N_43616,N_42597);
xor U44122 (N_44122,N_43503,N_43290);
xnor U44123 (N_44123,N_42796,N_43319);
nand U44124 (N_44124,N_43462,N_43955);
and U44125 (N_44125,N_43367,N_43996);
nand U44126 (N_44126,N_42425,N_42200);
and U44127 (N_44127,N_43775,N_43378);
and U44128 (N_44128,N_43228,N_42987);
nor U44129 (N_44129,N_43510,N_43791);
xor U44130 (N_44130,N_42990,N_42385);
or U44131 (N_44131,N_43968,N_42281);
and U44132 (N_44132,N_43493,N_42395);
xnor U44133 (N_44133,N_42136,N_42580);
xnor U44134 (N_44134,N_43466,N_42389);
nand U44135 (N_44135,N_43066,N_42309);
nor U44136 (N_44136,N_43568,N_42660);
xor U44137 (N_44137,N_43768,N_42719);
or U44138 (N_44138,N_42701,N_43948);
nor U44139 (N_44139,N_42798,N_42992);
or U44140 (N_44140,N_43895,N_42969);
nand U44141 (N_44141,N_43135,N_43081);
nor U44142 (N_44142,N_42427,N_43637);
and U44143 (N_44143,N_42841,N_42318);
nand U44144 (N_44144,N_43130,N_43607);
and U44145 (N_44145,N_42758,N_43337);
xor U44146 (N_44146,N_42978,N_42459);
or U44147 (N_44147,N_42130,N_43217);
nor U44148 (N_44148,N_42248,N_42562);
or U44149 (N_44149,N_42900,N_42106);
xor U44150 (N_44150,N_42475,N_43356);
xnor U44151 (N_44151,N_43580,N_43660);
xnor U44152 (N_44152,N_42835,N_43148);
nor U44153 (N_44153,N_43094,N_43139);
and U44154 (N_44154,N_42801,N_43309);
nor U44155 (N_44155,N_43564,N_42140);
and U44156 (N_44156,N_43257,N_43938);
or U44157 (N_44157,N_43521,N_43984);
nor U44158 (N_44158,N_43064,N_42637);
nand U44159 (N_44159,N_43585,N_42807);
or U44160 (N_44160,N_42435,N_43731);
nand U44161 (N_44161,N_43738,N_42342);
nor U44162 (N_44162,N_42945,N_43424);
xor U44163 (N_44163,N_43937,N_43145);
nor U44164 (N_44164,N_42994,N_43215);
or U44165 (N_44165,N_43177,N_43253);
or U44166 (N_44166,N_42190,N_42076);
nand U44167 (N_44167,N_43664,N_43945);
or U44168 (N_44168,N_42951,N_43998);
nor U44169 (N_44169,N_42093,N_43815);
nand U44170 (N_44170,N_42743,N_42633);
or U44171 (N_44171,N_43739,N_43157);
xnor U44172 (N_44172,N_43767,N_42166);
xnor U44173 (N_44173,N_43656,N_42569);
and U44174 (N_44174,N_42501,N_42911);
xnor U44175 (N_44175,N_43014,N_43371);
xnor U44176 (N_44176,N_43138,N_43111);
xnor U44177 (N_44177,N_43539,N_43410);
and U44178 (N_44178,N_43483,N_42138);
nand U44179 (N_44179,N_43050,N_42683);
or U44180 (N_44180,N_42479,N_43069);
nand U44181 (N_44181,N_42003,N_42325);
nor U44182 (N_44182,N_43526,N_42956);
or U44183 (N_44183,N_42492,N_43283);
xor U44184 (N_44184,N_42736,N_43085);
and U44185 (N_44185,N_42679,N_42469);
or U44186 (N_44186,N_43394,N_42936);
or U44187 (N_44187,N_42039,N_42793);
or U44188 (N_44188,N_43547,N_43603);
or U44189 (N_44189,N_42704,N_43803);
or U44190 (N_44190,N_43070,N_43962);
and U44191 (N_44191,N_43456,N_42329);
or U44192 (N_44192,N_42111,N_42495);
or U44193 (N_44193,N_43659,N_43508);
or U44194 (N_44194,N_42036,N_42474);
nor U44195 (N_44195,N_43134,N_42006);
nor U44196 (N_44196,N_42135,N_42705);
nand U44197 (N_44197,N_42858,N_43687);
or U44198 (N_44198,N_42842,N_42440);
and U44199 (N_44199,N_42150,N_42769);
nand U44200 (N_44200,N_42210,N_43906);
nand U44201 (N_44201,N_43207,N_43305);
nand U44202 (N_44202,N_43464,N_42824);
and U44203 (N_44203,N_42301,N_43180);
nand U44204 (N_44204,N_43191,N_42374);
nor U44205 (N_44205,N_42129,N_42776);
nand U44206 (N_44206,N_43919,N_42442);
nor U44207 (N_44207,N_42531,N_42125);
or U44208 (N_44208,N_42172,N_43595);
xnor U44209 (N_44209,N_42965,N_43920);
nor U44210 (N_44210,N_43719,N_43296);
xnor U44211 (N_44211,N_43504,N_42816);
nand U44212 (N_44212,N_43635,N_43324);
xor U44213 (N_44213,N_43254,N_42861);
xnor U44214 (N_44214,N_42235,N_43685);
xnor U44215 (N_44215,N_43972,N_43929);
xor U44216 (N_44216,N_42689,N_42878);
and U44217 (N_44217,N_43225,N_42870);
or U44218 (N_44218,N_43949,N_43567);
or U44219 (N_44219,N_43156,N_42292);
or U44220 (N_44220,N_43748,N_43183);
xnor U44221 (N_44221,N_42225,N_42998);
xnor U44222 (N_44222,N_43866,N_42883);
or U44223 (N_44223,N_43231,N_43954);
or U44224 (N_44224,N_42397,N_43771);
or U44225 (N_44225,N_43175,N_42198);
nand U44226 (N_44226,N_43074,N_42431);
and U44227 (N_44227,N_42403,N_43862);
xnor U44228 (N_44228,N_43571,N_43628);
or U44229 (N_44229,N_42691,N_43737);
nand U44230 (N_44230,N_43412,N_42749);
xor U44231 (N_44231,N_43300,N_42742);
nor U44232 (N_44232,N_42601,N_43428);
nor U44233 (N_44233,N_42507,N_42768);
nor U44234 (N_44234,N_43801,N_43281);
nand U44235 (N_44235,N_42727,N_42350);
xnor U44236 (N_44236,N_42702,N_43028);
nand U44237 (N_44237,N_43128,N_43315);
or U44238 (N_44238,N_42196,N_42613);
xor U44239 (N_44239,N_42687,N_42262);
or U44240 (N_44240,N_42386,N_42536);
and U44241 (N_44241,N_42438,N_43787);
xor U44242 (N_44242,N_43781,N_42145);
nand U44243 (N_44243,N_43452,N_42811);
or U44244 (N_44244,N_42251,N_43570);
and U44245 (N_44245,N_43956,N_42457);
xor U44246 (N_44246,N_43480,N_43876);
xor U44247 (N_44247,N_42762,N_42061);
nand U44248 (N_44248,N_43322,N_43162);
and U44249 (N_44249,N_42169,N_42607);
nand U44250 (N_44250,N_42411,N_43629);
nand U44251 (N_44251,N_43318,N_42274);
or U44252 (N_44252,N_43181,N_43335);
or U44253 (N_44253,N_43648,N_43592);
and U44254 (N_44254,N_42107,N_43649);
and U44255 (N_44255,N_42387,N_43423);
nand U44256 (N_44256,N_42699,N_42959);
and U44257 (N_44257,N_43868,N_43900);
xnor U44258 (N_44258,N_43836,N_42971);
or U44259 (N_44259,N_43248,N_43522);
nand U44260 (N_44260,N_43276,N_42737);
and U44261 (N_44261,N_42582,N_43224);
and U44262 (N_44262,N_43350,N_43475);
or U44263 (N_44263,N_42339,N_43502);
nor U44264 (N_44264,N_43251,N_42682);
and U44265 (N_44265,N_42478,N_42899);
xnor U44266 (N_44266,N_43090,N_42437);
nor U44267 (N_44267,N_42337,N_43942);
nand U44268 (N_44268,N_42511,N_42831);
nand U44269 (N_44269,N_42306,N_43770);
nor U44270 (N_44270,N_42345,N_42289);
nand U44271 (N_44271,N_42487,N_42078);
nand U44272 (N_44272,N_43882,N_42777);
or U44273 (N_44273,N_43921,N_43506);
nor U44274 (N_44274,N_43857,N_42904);
nor U44275 (N_44275,N_43472,N_42979);
xnor U44276 (N_44276,N_43651,N_43816);
nor U44277 (N_44277,N_42112,N_43030);
nand U44278 (N_44278,N_43210,N_43223);
and U44279 (N_44279,N_42676,N_42113);
xnor U44280 (N_44280,N_42034,N_42754);
nand U44281 (N_44281,N_43684,N_42184);
nor U44282 (N_44282,N_43294,N_42708);
or U44283 (N_44283,N_42258,N_42445);
or U44284 (N_44284,N_43059,N_43814);
and U44285 (N_44285,N_43764,N_42964);
or U44286 (N_44286,N_43463,N_42018);
nor U44287 (N_44287,N_42880,N_43697);
xnor U44288 (N_44288,N_43980,N_43288);
and U44289 (N_44289,N_42030,N_43089);
nand U44290 (N_44290,N_42739,N_43476);
xor U44291 (N_44291,N_42191,N_42912);
nand U44292 (N_44292,N_42888,N_43076);
or U44293 (N_44293,N_42277,N_42486);
nor U44294 (N_44294,N_42514,N_42715);
and U44295 (N_44295,N_43336,N_42099);
nor U44296 (N_44296,N_42649,N_42223);
or U44297 (N_44297,N_43034,N_43380);
nand U44298 (N_44298,N_43729,N_42011);
xnor U44299 (N_44299,N_42177,N_43549);
or U44300 (N_44300,N_43012,N_42022);
or U44301 (N_44301,N_43267,N_42077);
xor U44302 (N_44302,N_43811,N_43721);
and U44303 (N_44303,N_42810,N_43891);
or U44304 (N_44304,N_43013,N_42396);
or U44305 (N_44305,N_43716,N_43896);
and U44306 (N_44306,N_42415,N_42952);
or U44307 (N_44307,N_43658,N_42763);
xor U44308 (N_44308,N_42829,N_43890);
xor U44309 (N_44309,N_43916,N_42470);
and U44310 (N_44310,N_42228,N_43981);
and U44311 (N_44311,N_43880,N_43007);
and U44312 (N_44312,N_43489,N_43507);
nor U44313 (N_44313,N_42584,N_43971);
xor U44314 (N_44314,N_42837,N_43271);
xnor U44315 (N_44315,N_42468,N_43259);
nor U44316 (N_44316,N_42639,N_43136);
and U44317 (N_44317,N_43757,N_43390);
or U44318 (N_44318,N_43796,N_43116);
nand U44319 (N_44319,N_42503,N_42830);
xor U44320 (N_44320,N_43517,N_43190);
nand U44321 (N_44321,N_42259,N_43328);
and U44322 (N_44322,N_43146,N_43732);
nand U44323 (N_44323,N_42282,N_43105);
xor U44324 (N_44324,N_43065,N_43467);
nand U44325 (N_44325,N_43670,N_42362);
and U44326 (N_44326,N_42631,N_42895);
and U44327 (N_44327,N_42133,N_43840);
and U44328 (N_44328,N_43272,N_43079);
nand U44329 (N_44329,N_42239,N_42803);
and U44330 (N_44330,N_43859,N_42693);
and U44331 (N_44331,N_43379,N_42246);
xor U44332 (N_44332,N_42694,N_42103);
and U44333 (N_44333,N_42869,N_43373);
nand U44334 (N_44334,N_42142,N_42080);
nand U44335 (N_44335,N_42902,N_42581);
nor U44336 (N_44336,N_43389,N_43983);
xnor U44337 (N_44337,N_43017,N_42680);
nor U44338 (N_44338,N_42655,N_43703);
and U44339 (N_44339,N_42269,N_43255);
xor U44340 (N_44340,N_42575,N_43743);
nand U44341 (N_44341,N_42799,N_42592);
nand U44342 (N_44342,N_42589,N_42929);
xor U44343 (N_44343,N_43877,N_42019);
xnor U44344 (N_44344,N_42448,N_43016);
or U44345 (N_44345,N_42672,N_43348);
nor U44346 (N_44346,N_42009,N_42608);
nand U44347 (N_44347,N_43123,N_42338);
or U44348 (N_44348,N_43075,N_42341);
xnor U44349 (N_44349,N_42024,N_42173);
or U44350 (N_44350,N_43661,N_43313);
nand U44351 (N_44351,N_43641,N_43221);
and U44352 (N_44352,N_43544,N_43542);
nor U44353 (N_44353,N_43758,N_42370);
xor U44354 (N_44354,N_42300,N_42148);
nand U44355 (N_44355,N_42565,N_43406);
xor U44356 (N_44356,N_43941,N_42875);
nor U44357 (N_44357,N_42443,N_42314);
nand U44358 (N_44358,N_42104,N_43256);
xor U44359 (N_44359,N_42868,N_42460);
and U44360 (N_44360,N_43830,N_42351);
and U44361 (N_44361,N_43031,N_43928);
and U44362 (N_44362,N_43715,N_42897);
and U44363 (N_44363,N_42604,N_42490);
nor U44364 (N_44364,N_43198,N_42454);
and U44365 (N_44365,N_42116,N_43201);
nor U44366 (N_44366,N_43170,N_43446);
xnor U44367 (N_44367,N_43250,N_43846);
and U44368 (N_44368,N_42759,N_43039);
nand U44369 (N_44369,N_43754,N_43609);
and U44370 (N_44370,N_43922,N_42989);
nand U44371 (N_44371,N_43683,N_42273);
and U44372 (N_44372,N_42193,N_43473);
and U44373 (N_44373,N_43416,N_42973);
nor U44374 (N_44374,N_42373,N_42464);
nor U44375 (N_44375,N_42838,N_43888);
xnor U44376 (N_44376,N_42252,N_42890);
xor U44377 (N_44377,N_43167,N_43258);
nand U44378 (N_44378,N_43565,N_42730);
or U44379 (N_44379,N_42508,N_43142);
nand U44380 (N_44380,N_43329,N_42937);
nor U44381 (N_44381,N_43749,N_42712);
or U44382 (N_44382,N_42728,N_42047);
nor U44383 (N_44383,N_42371,N_43077);
xnor U44384 (N_44384,N_42761,N_42738);
nor U44385 (N_44385,N_43484,N_43205);
nand U44386 (N_44386,N_43558,N_43151);
or U44387 (N_44387,N_43291,N_43622);
nand U44388 (N_44388,N_43707,N_42845);
nand U44389 (N_44389,N_43875,N_43227);
xor U44390 (N_44390,N_42662,N_42233);
nand U44391 (N_44391,N_42527,N_42361);
nor U44392 (N_44392,N_43244,N_42170);
nand U44393 (N_44393,N_42360,N_42781);
xor U44394 (N_44394,N_43098,N_42620);
nand U44395 (N_44395,N_42583,N_43194);
and U44396 (N_44396,N_42118,N_42045);
nand U44397 (N_44397,N_43479,N_43342);
or U44398 (N_44398,N_43573,N_42205);
or U44399 (N_44399,N_43091,N_43638);
nand U44400 (N_44400,N_42795,N_42178);
or U44401 (N_44401,N_43718,N_42640);
xor U44402 (N_44402,N_42356,N_42540);
xor U44403 (N_44403,N_42471,N_43451);
xor U44404 (N_44404,N_42408,N_43935);
or U44405 (N_44405,N_42452,N_43192);
and U44406 (N_44406,N_42591,N_42050);
and U44407 (N_44407,N_43889,N_42918);
nand U44408 (N_44408,N_43509,N_43530);
and U44409 (N_44409,N_43711,N_43583);
nand U44410 (N_44410,N_43120,N_42643);
or U44411 (N_44411,N_43572,N_43911);
nand U44412 (N_44412,N_43439,N_42384);
nor U44413 (N_44413,N_43369,N_43673);
and U44414 (N_44414,N_42211,N_42161);
and U44415 (N_44415,N_43165,N_42375);
xor U44416 (N_44416,N_42168,N_43520);
or U44417 (N_44417,N_43021,N_43112);
xor U44418 (N_44418,N_42787,N_43923);
and U44419 (N_44419,N_42433,N_42741);
xor U44420 (N_44420,N_42174,N_43270);
nor U44421 (N_44421,N_43200,N_43505);
xnor U44422 (N_44422,N_43666,N_42155);
nand U44423 (N_44423,N_43084,N_42353);
or U44424 (N_44424,N_42653,N_43100);
nand U44425 (N_44425,N_43127,N_42084);
nor U44426 (N_44426,N_43442,N_42451);
or U44427 (N_44427,N_42843,N_42532);
and U44428 (N_44428,N_42865,N_42021);
or U44429 (N_44429,N_42227,N_43360);
or U44430 (N_44430,N_43799,N_42734);
nand U44431 (N_44431,N_42243,N_43041);
xnor U44432 (N_44432,N_43323,N_43704);
xor U44433 (N_44433,N_43437,N_42098);
nand U44434 (N_44434,N_42863,N_42755);
nand U44435 (N_44435,N_42131,N_43429);
nand U44436 (N_44436,N_42040,N_42997);
nor U44437 (N_44437,N_43858,N_42955);
and U44438 (N_44438,N_42630,N_42075);
or U44439 (N_44439,N_42770,N_42418);
or U44440 (N_44440,N_43784,N_42877);
nand U44441 (N_44441,N_43679,N_43820);
and U44442 (N_44442,N_42149,N_43058);
xor U44443 (N_44443,N_42571,N_42352);
or U44444 (N_44444,N_42785,N_43046);
nand U44445 (N_44445,N_43632,N_42558);
and U44446 (N_44446,N_42453,N_42417);
nand U44447 (N_44447,N_43752,N_43497);
or U44448 (N_44448,N_43753,N_42023);
nor U44449 (N_44449,N_42578,N_43436);
and U44450 (N_44450,N_42626,N_43910);
nor U44451 (N_44451,N_43925,N_42709);
or U44452 (N_44452,N_42988,N_42725);
nand U44453 (N_44453,N_42152,N_43982);
or U44454 (N_44454,N_42594,N_42731);
and U44455 (N_44455,N_42856,N_43161);
nand U44456 (N_44456,N_43419,N_43003);
and U44457 (N_44457,N_42780,N_42542);
nor U44458 (N_44458,N_43556,N_42378);
xnor U44459 (N_44459,N_42636,N_42399);
xor U44460 (N_44460,N_43667,N_43339);
nor U44461 (N_44461,N_42879,N_43032);
xnor U44462 (N_44462,N_43843,N_42004);
nor U44463 (N_44463,N_42413,N_42804);
xor U44464 (N_44464,N_42894,N_43907);
and U44465 (N_44465,N_43519,N_42313);
xnor U44466 (N_44466,N_42089,N_43408);
or U44467 (N_44467,N_43438,N_42467);
or U44468 (N_44468,N_42910,N_43712);
nor U44469 (N_44469,N_42214,N_43345);
nand U44470 (N_44470,N_43887,N_42144);
and U44471 (N_44471,N_42081,N_43459);
nor U44472 (N_44472,N_43080,N_42002);
and U44473 (N_44473,N_42534,N_43690);
or U44474 (N_44474,N_42238,N_42293);
and U44475 (N_44475,N_43960,N_42772);
xor U44476 (N_44476,N_43674,N_42247);
nand U44477 (N_44477,N_43579,N_43140);
or U44478 (N_44478,N_42154,N_42156);
xnor U44479 (N_44479,N_43642,N_43103);
or U44480 (N_44480,N_42745,N_42195);
xor U44481 (N_44481,N_43788,N_43533);
or U44482 (N_44482,N_42049,N_43158);
or U44483 (N_44483,N_42664,N_43855);
nor U44484 (N_44484,N_43088,N_43681);
and U44485 (N_44485,N_42493,N_42999);
xor U44486 (N_44486,N_43640,N_43263);
or U44487 (N_44487,N_42669,N_43153);
or U44488 (N_44488,N_43481,N_42284);
or U44489 (N_44489,N_42412,N_42266);
nand U44490 (N_44490,N_42450,N_43049);
and U44491 (N_44491,N_43939,N_43193);
and U44492 (N_44492,N_43783,N_42175);
xnor U44493 (N_44493,N_43126,N_42058);
nand U44494 (N_44494,N_43332,N_42596);
and U44495 (N_44495,N_43722,N_43047);
and U44496 (N_44496,N_43606,N_42072);
nand U44497 (N_44497,N_43529,N_43114);
xnor U44498 (N_44498,N_43734,N_43119);
nand U44499 (N_44499,N_43330,N_42127);
and U44500 (N_44500,N_42358,N_42151);
or U44501 (N_44501,N_42485,N_43381);
nor U44502 (N_44502,N_43358,N_43950);
xnor U44503 (N_44503,N_42053,N_43967);
xor U44504 (N_44504,N_42813,N_42483);
nor U44505 (N_44505,N_43368,N_42307);
or U44506 (N_44506,N_42382,N_43848);
xor U44507 (N_44507,N_43426,N_42206);
xnor U44508 (N_44508,N_42744,N_42042);
or U44509 (N_44509,N_42853,N_43824);
and U44510 (N_44510,N_42808,N_42938);
and U44511 (N_44511,N_42097,N_43022);
nand U44512 (N_44512,N_42934,N_42044);
and U44513 (N_44513,N_42792,N_43613);
or U44514 (N_44514,N_42933,N_42647);
nand U44515 (N_44515,N_42983,N_43973);
xnor U44516 (N_44516,N_43688,N_43728);
and U44517 (N_44517,N_42232,N_42593);
or U44518 (N_44518,N_42823,N_43229);
nor U44519 (N_44519,N_42675,N_42889);
and U44520 (N_44520,N_42254,N_43934);
or U44521 (N_44521,N_43701,N_43534);
xnor U44522 (N_44522,N_42421,N_43853);
nand U44523 (N_44523,N_43386,N_42222);
nor U44524 (N_44524,N_43152,N_43435);
xor U44525 (N_44525,N_43693,N_43405);
xnor U44526 (N_44526,N_42276,N_42041);
xnor U44527 (N_44527,N_42552,N_43474);
and U44528 (N_44528,N_43773,N_43994);
and U44529 (N_44529,N_42529,N_42818);
nor U44530 (N_44530,N_42654,N_43492);
nand U44531 (N_44531,N_43874,N_43247);
nor U44532 (N_44532,N_42398,N_42984);
nand U44533 (N_44533,N_43314,N_42614);
nor U44534 (N_44534,N_42182,N_42543);
xor U44535 (N_44535,N_43959,N_42291);
nand U44536 (N_44536,N_43166,N_43125);
or U44537 (N_44537,N_43759,N_42794);
and U44538 (N_44538,N_43705,N_43845);
xor U44539 (N_44539,N_42697,N_42944);
xnor U44540 (N_44540,N_43551,N_43370);
xnor U44541 (N_44541,N_43924,N_42165);
xor U44542 (N_44542,N_43009,N_42366);
xor U44543 (N_44543,N_43837,N_43841);
nand U44544 (N_44544,N_42515,N_43197);
xor U44545 (N_44545,N_43160,N_43700);
nand U44546 (N_44546,N_42550,N_42481);
or U44547 (N_44547,N_43216,N_42555);
or U44548 (N_44548,N_42379,N_43665);
or U44549 (N_44549,N_42381,N_42456);
nand U44550 (N_44550,N_43187,N_43677);
or U44551 (N_44551,N_43869,N_43432);
nor U44552 (N_44552,N_43755,N_43527);
xnor U44553 (N_44553,N_43672,N_42632);
or U44554 (N_44554,N_43696,N_42651);
or U44555 (N_44555,N_43430,N_43052);
and U44556 (N_44556,N_42392,N_42414);
xor U44557 (N_44557,N_42782,N_43714);
nor U44558 (N_44558,N_43795,N_43951);
nor U44559 (N_44559,N_42692,N_43427);
and U44560 (N_44560,N_43445,N_43892);
xnor U44561 (N_44561,N_42826,N_42295);
or U44562 (N_44562,N_43639,N_42240);
xor U44563 (N_44563,N_43008,N_42365);
xor U44564 (N_44564,N_42605,N_43035);
or U44565 (N_44565,N_42602,N_43172);
nand U44566 (N_44566,N_43141,N_42551);
and U44567 (N_44567,N_43733,N_42844);
nand U44568 (N_44568,N_43067,N_43054);
or U44569 (N_44569,N_42430,N_43709);
nand U44570 (N_44570,N_42340,N_43550);
and U44571 (N_44571,N_42579,N_42139);
or U44572 (N_44572,N_42176,N_43132);
and U44573 (N_44573,N_42783,N_43978);
xor U44574 (N_44574,N_43897,N_42027);
nand U44575 (N_44575,N_42560,N_42947);
nor U44576 (N_44576,N_42088,N_42245);
nor U44577 (N_44577,N_42642,N_43202);
nand U44578 (N_44578,N_42598,N_42263);
and U44579 (N_44579,N_42404,N_42372);
and U44580 (N_44580,N_43115,N_43208);
or U44581 (N_44581,N_43849,N_43647);
nand U44582 (N_44582,N_42898,N_42684);
nor U44583 (N_44583,N_43289,N_42517);
and U44584 (N_44584,N_42327,N_42960);
xor U44585 (N_44585,N_43222,N_43211);
nand U44586 (N_44586,N_43310,N_42094);
nor U44587 (N_44587,N_42110,N_43810);
and U44588 (N_44588,N_42446,N_42663);
and U44589 (N_44589,N_43692,N_42199);
nor U44590 (N_44590,N_42733,N_43860);
or U44591 (N_44591,N_42261,N_43985);
nand U44592 (N_44592,N_43387,N_43831);
xnor U44593 (N_44593,N_42192,N_43461);
nor U44594 (N_44594,N_43196,N_42028);
nand U44595 (N_44595,N_43286,N_43671);
xnor U44596 (N_44596,N_43798,N_42153);
nor U44597 (N_44597,N_42919,N_43561);
nand U44598 (N_44598,N_42718,N_43852);
nor U44599 (N_44599,N_43663,N_42615);
nor U44600 (N_44600,N_42108,N_42477);
nor U44601 (N_44601,N_43577,N_42686);
nor U44602 (N_44602,N_42032,N_42060);
nor U44603 (N_44603,N_43511,N_42673);
xnor U44604 (N_44604,N_43209,N_43636);
or U44605 (N_44605,N_42201,N_42120);
xor U44606 (N_44606,N_42713,N_43176);
and U44607 (N_44607,N_42541,N_43689);
xor U44608 (N_44608,N_43122,N_43706);
or U44609 (N_44609,N_42380,N_42489);
xnor U44610 (N_44610,N_43099,N_43491);
xnor U44611 (N_44611,N_43953,N_42069);
and U44612 (N_44612,N_42817,N_42090);
xor U44613 (N_44613,N_42574,N_43295);
nor U44614 (N_44614,N_43361,N_43469);
nor U44615 (N_44615,N_43524,N_43601);
and U44616 (N_44616,N_42279,N_43587);
xor U44617 (N_44617,N_43062,N_43545);
nand U44618 (N_44618,N_42674,N_42907);
xor U44619 (N_44619,N_43886,N_43374);
and U44620 (N_44620,N_43087,N_43243);
and U44621 (N_44621,N_43741,N_42624);
nor U44622 (N_44622,N_42391,N_43147);
and U44623 (N_44623,N_42622,N_43388);
xnor U44624 (N_44624,N_42606,N_43908);
xor U44625 (N_44625,N_42416,N_43501);
and U44626 (N_44626,N_42621,N_42547);
nor U44627 (N_44627,N_43979,N_42896);
or U44628 (N_44628,N_43593,N_42892);
and U44629 (N_44629,N_42970,N_43044);
nor U44630 (N_44630,N_42735,N_43917);
nor U44631 (N_44631,N_43965,N_43131);
nor U44632 (N_44632,N_42564,N_42208);
xnor U44633 (N_44633,N_43990,N_43218);
or U44634 (N_44634,N_42625,N_42980);
xor U44635 (N_44635,N_43992,N_43092);
xnor U44636 (N_44636,N_43071,N_43537);
nand U44637 (N_44637,N_43195,N_42359);
nor U44638 (N_44638,N_43655,N_42974);
xnor U44639 (N_44639,N_43249,N_42977);
nand U44640 (N_44640,N_43171,N_43015);
xor U44641 (N_44641,N_43991,N_42134);
xor U44642 (N_44642,N_43051,N_42789);
nand U44643 (N_44643,N_42059,N_43108);
nand U44644 (N_44644,N_42932,N_43591);
or U44645 (N_44645,N_42778,N_42257);
nor U44646 (N_44646,N_43850,N_42434);
nand U44647 (N_44647,N_42219,N_42832);
xnor U44648 (N_44648,N_43913,N_42645);
xor U44649 (N_44649,N_43179,N_42950);
or U44650 (N_44650,N_43024,N_43961);
xor U44651 (N_44651,N_42312,N_42696);
xor U44652 (N_44652,N_42126,N_42163);
or U44653 (N_44653,N_43602,N_42079);
or U44654 (N_44654,N_43219,N_42226);
and U44655 (N_44655,N_43847,N_42957);
and U44656 (N_44656,N_42695,N_42335);
or U44657 (N_44657,N_43624,N_43989);
and U44658 (N_44658,N_42665,N_42854);
xnor U44659 (N_44659,N_42143,N_43362);
nor U44660 (N_44660,N_43861,N_43001);
or U44661 (N_44661,N_42220,N_43488);
and U44662 (N_44662,N_42723,N_42926);
and U44663 (N_44663,N_42963,N_43525);
nor U44664 (N_44664,N_42616,N_42287);
xor U44665 (N_44665,N_42628,N_43988);
nor U44666 (N_44666,N_43365,N_42935);
or U44667 (N_44667,N_42819,N_42260);
and U44668 (N_44668,N_42588,N_42599);
and U44669 (N_44669,N_42305,N_43952);
or U44670 (N_44670,N_43457,N_42610);
xnor U44671 (N_44671,N_43298,N_42067);
xor U44672 (N_44672,N_43654,N_42814);
or U44673 (N_44673,N_42472,N_43018);
and U44674 (N_44674,N_43072,N_43789);
nand U44675 (N_44675,N_42634,N_43546);
and U44676 (N_44676,N_43594,N_43307);
and U44677 (N_44677,N_42224,N_42343);
or U44678 (N_44678,N_43987,N_43879);
nand U44679 (N_44679,N_43531,N_42026);
xor U44680 (N_44680,N_43144,N_42298);
nand U44681 (N_44681,N_43668,N_42057);
or U44682 (N_44682,N_42367,N_43724);
xnor U44683 (N_44683,N_43233,N_43274);
xor U44684 (N_44684,N_43818,N_42317);
nor U44685 (N_44685,N_43458,N_43772);
and U44686 (N_44686,N_42255,N_43809);
xor U44687 (N_44687,N_43899,N_42923);
xnor U44688 (N_44688,N_43155,N_43515);
nor U44689 (N_44689,N_42721,N_43317);
or U44690 (N_44690,N_43301,N_42388);
nand U44691 (N_44691,N_42958,N_42720);
xnor U44692 (N_44692,N_43612,N_43400);
nand U44693 (N_44693,N_42426,N_42916);
nor U44694 (N_44694,N_42436,N_42310);
xnor U44695 (N_44695,N_43725,N_43278);
and U44696 (N_44696,N_42491,N_42524);
nor U44697 (N_44697,N_43037,N_42171);
and U44698 (N_44698,N_42576,N_42092);
xnor U44699 (N_44699,N_43113,N_43401);
xor U44700 (N_44700,N_43865,N_43576);
and U44701 (N_44701,N_43808,N_43631);
nand U44702 (N_44702,N_42732,N_43496);
nor U44703 (N_44703,N_43970,N_42015);
nand U44704 (N_44704,N_42488,N_43827);
or U44705 (N_44705,N_43805,N_43265);
and U44706 (N_44706,N_42941,N_42834);
and U44707 (N_44707,N_43599,N_42369);
xor U44708 (N_44708,N_42644,N_42805);
or U44709 (N_44709,N_42005,N_43854);
xnor U44710 (N_44710,N_43653,N_43471);
nor U44711 (N_44711,N_43844,N_42827);
xnor U44712 (N_44712,N_43260,N_43863);
nor U44713 (N_44713,N_43302,N_42750);
nand U44714 (N_44714,N_42668,N_43033);
or U44715 (N_44715,N_43338,N_43352);
nand U44716 (N_44716,N_42638,N_42748);
and U44717 (N_44717,N_43417,N_42539);
and U44718 (N_44718,N_42521,N_43444);
nand U44719 (N_44719,N_43232,N_42847);
nor U44720 (N_44720,N_43590,N_42146);
xor U44721 (N_44721,N_42500,N_42181);
xnor U44722 (N_44722,N_43536,N_43235);
xnor U44723 (N_44723,N_43118,N_43766);
and U44724 (N_44724,N_43385,N_42572);
and U44725 (N_44725,N_43055,N_43553);
nor U44726 (N_44726,N_42000,N_43723);
nor U44727 (N_44727,N_42082,N_43448);
xor U44728 (N_44728,N_43744,N_42771);
xor U44729 (N_44729,N_43695,N_42502);
nand U44730 (N_44730,N_43261,N_42635);
xor U44731 (N_44731,N_42095,N_42064);
nand U44732 (N_44732,N_42617,N_43434);
nand U44733 (N_44733,N_42953,N_42267);
nand U44734 (N_44734,N_42401,N_42216);
nand U44735 (N_44735,N_43273,N_43630);
xnor U44736 (N_44736,N_43242,N_42229);
nor U44737 (N_44737,N_42711,N_42928);
nand U44738 (N_44738,N_42197,N_42074);
nor U44739 (N_44739,N_43431,N_43023);
nor U44740 (N_44740,N_42688,N_43769);
nor U44741 (N_44741,N_42390,N_42577);
or U44742 (N_44742,N_43969,N_42866);
nand U44743 (N_44743,N_43331,N_43931);
xnor U44744 (N_44744,N_43822,N_43000);
or U44745 (N_44745,N_42480,N_43004);
xor U44746 (N_44746,N_43596,N_42315);
xnor U44747 (N_44747,N_43621,N_43713);
xnor U44748 (N_44748,N_43823,N_43997);
or U44749 (N_44749,N_42137,N_43940);
or U44750 (N_44750,N_42554,N_43686);
nand U44751 (N_44751,N_43785,N_43828);
xor U44752 (N_44752,N_43407,N_43383);
nor U44753 (N_44753,N_42035,N_43234);
or U44754 (N_44754,N_42991,N_42463);
or U44755 (N_44755,N_42559,N_43717);
nand U44756 (N_44756,N_42849,N_42316);
or U44757 (N_44757,N_43441,N_42872);
and U44758 (N_44758,N_42449,N_42920);
and U44759 (N_44759,N_43574,N_42207);
nand U44760 (N_44760,N_42164,N_43107);
and U44761 (N_44761,N_42658,N_43774);
nand U44762 (N_44762,N_43239,N_42972);
or U44763 (N_44763,N_42465,N_42619);
nor U44764 (N_44764,N_43468,N_42722);
or U44765 (N_44765,N_43708,N_43343);
and U44766 (N_44766,N_43975,N_43730);
nor U44767 (N_44767,N_42931,N_42766);
nor U44768 (N_44768,N_42603,N_42029);
and U44769 (N_44769,N_42840,N_42236);
and U44770 (N_44770,N_42707,N_42925);
xor U44771 (N_44771,N_42586,N_42406);
nor U44772 (N_44772,N_43742,N_43562);
nand U44773 (N_44773,N_43382,N_42303);
nor U44774 (N_44774,N_43676,N_43042);
and U44775 (N_44775,N_43548,N_43002);
nand U44776 (N_44776,N_42661,N_43779);
and U44777 (N_44777,N_43646,N_43325);
or U44778 (N_44778,N_42194,N_43414);
nor U44779 (N_44779,N_42563,N_43838);
and U44780 (N_44780,N_43974,N_42800);
and U44781 (N_44781,N_43482,N_43096);
nand U44782 (N_44782,N_43986,N_42505);
nand U44783 (N_44783,N_42549,N_43589);
or U44784 (N_44784,N_43236,N_43871);
nand U44785 (N_44785,N_43159,N_43777);
xor U44786 (N_44786,N_43220,N_42546);
xor U44787 (N_44787,N_42123,N_42747);
and U44788 (N_44788,N_43751,N_43460);
and U44789 (N_44789,N_42522,N_43745);
and U44790 (N_44790,N_43149,N_42033);
nor U44791 (N_44791,N_43326,N_43761);
or U44792 (N_44792,N_42428,N_42439);
or U44793 (N_44793,N_42221,N_42648);
xor U44794 (N_44794,N_42884,N_43104);
or U44795 (N_44795,N_42117,N_42458);
and U44796 (N_44796,N_42646,N_43415);
or U44797 (N_44797,N_42473,N_43883);
nor U44798 (N_44798,N_42906,N_42942);
xor U44799 (N_44799,N_43669,N_43633);
xor U44800 (N_44800,N_43063,N_42760);
and U44801 (N_44801,N_43878,N_43465);
xor U44802 (N_44802,N_43946,N_42567);
and U44803 (N_44803,N_42946,N_43292);
xnor U44804 (N_44804,N_43901,N_43341);
xnor U44805 (N_44805,N_43344,N_43614);
nor U44806 (N_44806,N_42203,N_43413);
or U44807 (N_44807,N_42520,N_42773);
xnor U44808 (N_44808,N_43395,N_43366);
xnor U44809 (N_44809,N_43662,N_42185);
and U44810 (N_44810,N_42025,N_42215);
xor U44811 (N_44811,N_42954,N_42419);
nor U44812 (N_44812,N_43409,N_42886);
or U44813 (N_44813,N_43842,N_42656);
or U44814 (N_44814,N_42537,N_42217);
nor U44815 (N_44815,N_43873,N_43340);
nand U44816 (N_44816,N_42774,N_42659);
xnor U44817 (N_44817,N_43682,N_42836);
nand U44818 (N_44818,N_42557,N_43964);
and U44819 (N_44819,N_42751,N_43523);
xnor U44820 (N_44820,N_42717,N_42124);
xor U44821 (N_44821,N_43311,N_42828);
or U44822 (N_44822,N_42996,N_43038);
nand U44823 (N_44823,N_42678,N_43834);
nand U44824 (N_44824,N_43391,N_43977);
and U44825 (N_44825,N_43894,N_42091);
and U44826 (N_44826,N_43552,N_43487);
xnor U44827 (N_44827,N_42740,N_43287);
nor U44828 (N_44828,N_43905,N_43903);
nor U44829 (N_44829,N_43760,N_42065);
nand U44830 (N_44830,N_43238,N_42855);
and U44831 (N_44831,N_42915,N_42882);
xor U44832 (N_44832,N_43040,N_43726);
xnor U44833 (N_44833,N_42526,N_42405);
and U44834 (N_44834,N_42806,N_42504);
nand U44835 (N_44835,N_43512,N_43586);
and U44836 (N_44836,N_42409,N_43443);
and U44837 (N_44837,N_42943,N_43600);
and U44838 (N_44838,N_42966,N_43275);
xnor U44839 (N_44839,N_43097,N_43563);
nor U44840 (N_44840,N_43312,N_42497);
and U44841 (N_44841,N_42056,N_42786);
nor U44842 (N_44842,N_42423,N_43912);
nand U44843 (N_44843,N_42876,N_43541);
nor U44844 (N_44844,N_42484,N_42319);
xnor U44845 (N_44845,N_42513,N_42914);
and U44846 (N_44846,N_42031,N_42324);
xor U44847 (N_44847,N_42859,N_43182);
nand U44848 (N_44848,N_42538,N_42180);
xor U44849 (N_44849,N_42466,N_43068);
nor U44850 (N_44850,N_43364,N_42244);
xor U44851 (N_44851,N_43174,N_43644);
and U44852 (N_44852,N_43710,N_42752);
nand U44853 (N_44853,N_43782,N_43433);
xor U44854 (N_44854,N_42864,N_43825);
and U44855 (N_44855,N_42241,N_43304);
xor U44856 (N_44856,N_42981,N_42323);
nand U44857 (N_44857,N_42158,N_42706);
nand U44858 (N_44858,N_42302,N_43321);
and U44859 (N_44859,N_43188,N_43214);
and U44860 (N_44860,N_43839,N_42014);
xnor U44861 (N_44861,N_42874,N_43786);
nor U44862 (N_44862,N_42212,N_42462);
or U44863 (N_44863,N_42141,N_43154);
or U44864 (N_44864,N_43106,N_42101);
nand U44865 (N_44865,N_42746,N_42288);
xor U44866 (N_44866,N_42652,N_43377);
nor U44867 (N_44867,N_43762,N_42402);
and U44868 (N_44868,N_42218,N_42283);
or U44869 (N_44869,N_43316,N_42618);
nand U44870 (N_44870,N_42046,N_43020);
and U44871 (N_44871,N_42523,N_42927);
or U44872 (N_44872,N_43993,N_43308);
xnor U44873 (N_44873,N_42297,N_43268);
or U44874 (N_44874,N_43376,N_42204);
nand U44875 (N_44875,N_42512,N_42346);
nor U44876 (N_44876,N_43740,N_42641);
or U44877 (N_44877,N_43643,N_43893);
xor U44878 (N_44878,N_42062,N_42667);
xnor U44879 (N_44879,N_42518,N_42924);
and U44880 (N_44880,N_43375,N_43060);
nand U44881 (N_44881,N_42407,N_42986);
nor U44882 (N_44882,N_42724,N_43102);
nand U44883 (N_44883,N_43036,N_42822);
nand U44884 (N_44884,N_43832,N_42867);
nand U44885 (N_44885,N_43213,N_43264);
nor U44886 (N_44886,N_42767,N_42887);
or U44887 (N_44887,N_42852,N_43354);
and U44888 (N_44888,N_42278,N_43025);
nor U44889 (N_44889,N_43735,N_43398);
nand U44890 (N_44890,N_43927,N_42400);
and U44891 (N_44891,N_43061,N_42609);
nand U44892 (N_44892,N_43057,N_43299);
or U44893 (N_44893,N_43121,N_42726);
and U44894 (N_44894,N_43082,N_43806);
and U44895 (N_44895,N_43652,N_42119);
xnor U44896 (N_44896,N_42909,N_42012);
or U44897 (N_44897,N_43604,N_43797);
xnor U44898 (N_44898,N_43650,N_43495);
nand U44899 (N_44899,N_43269,N_42394);
and U44900 (N_44900,N_43780,N_42670);
xnor U44901 (N_44901,N_43184,N_43675);
nor U44902 (N_44902,N_42275,N_43535);
nor U44903 (N_44903,N_43189,N_42921);
xnor U44904 (N_44904,N_42698,N_42775);
nor U44905 (N_44905,N_43226,N_42347);
xor U44906 (N_44906,N_42922,N_42147);
nor U44907 (N_44907,N_42322,N_42765);
or U44908 (N_44908,N_43078,N_43930);
nor U44909 (N_44909,N_43124,N_43420);
and U44910 (N_44910,N_43720,N_42535);
and U44911 (N_44911,N_43926,N_43943);
or U44912 (N_44912,N_43402,N_43347);
nor U44913 (N_44913,N_43817,N_42048);
nor U44914 (N_44914,N_43627,N_42525);
nor U44915 (N_44915,N_43262,N_42940);
xor U44916 (N_44916,N_42268,N_42179);
or U44917 (N_44917,N_42115,N_43245);
xnor U44918 (N_44918,N_42873,N_42871);
xnor U44919 (N_44919,N_43995,N_42231);
nor U44920 (N_44920,N_43333,N_43598);
nor U44921 (N_44921,N_43212,N_43027);
xor U44922 (N_44922,N_43776,N_43918);
or U44923 (N_44923,N_42757,N_42264);
nand U44924 (N_44924,N_42102,N_43566);
xnor U44925 (N_44925,N_43240,N_42294);
xor U44926 (N_44926,N_42509,N_43812);
nor U44927 (N_44927,N_43206,N_42157);
xor U44928 (N_44928,N_43447,N_42332);
and U44929 (N_44929,N_42833,N_42209);
nand U44930 (N_44930,N_42444,N_43204);
nor U44931 (N_44931,N_43763,N_42017);
and U44932 (N_44932,N_42510,N_43241);
xor U44933 (N_44933,N_43346,N_43540);
or U44934 (N_44934,N_43404,N_42368);
and U44935 (N_44935,N_43303,N_42334);
or U44936 (N_44936,N_42121,N_42982);
nand U44937 (N_44937,N_42519,N_43645);
and U44938 (N_44938,N_43582,N_43043);
nand U44939 (N_44939,N_42013,N_43625);
nor U44940 (N_44940,N_42285,N_42815);
or U44941 (N_44941,N_43957,N_42677);
and U44942 (N_44942,N_43056,N_42455);
and U44943 (N_44943,N_42070,N_43608);
nor U44944 (N_44944,N_43976,N_42908);
xor U44945 (N_44945,N_42189,N_42348);
xor U44946 (N_44946,N_42857,N_42304);
nor U44947 (N_44947,N_42355,N_43143);
xor U44948 (N_44948,N_43019,N_42043);
nand U44949 (N_44949,N_43513,N_42087);
nor U44950 (N_44950,N_42611,N_42051);
nand U44951 (N_44951,N_42328,N_42326);
and U44952 (N_44952,N_43909,N_43557);
nor U44953 (N_44953,N_43006,N_43807);
nor U44954 (N_44954,N_43528,N_42432);
nor U44955 (N_44955,N_43694,N_43657);
or U44956 (N_44956,N_43518,N_42967);
or U44957 (N_44957,N_43411,N_43372);
nand U44958 (N_44958,N_42710,N_42756);
or U44959 (N_44959,N_42570,N_43349);
xnor U44960 (N_44960,N_43778,N_42985);
nand U44961 (N_44961,N_43173,N_43399);
nand U44962 (N_44962,N_43355,N_43499);
and U44963 (N_44963,N_43199,N_43284);
or U44964 (N_44964,N_42714,N_42265);
nor U44965 (N_44965,N_43584,N_42993);
nand U44966 (N_44966,N_42802,N_42083);
or U44967 (N_44967,N_42296,N_43246);
and U44968 (N_44968,N_43053,N_43421);
nand U44969 (N_44969,N_43455,N_42891);
nor U44970 (N_44970,N_42716,N_43083);
nor U44971 (N_44971,N_42930,N_43958);
or U44972 (N_44972,N_43454,N_43230);
nor U44973 (N_44973,N_43702,N_43137);
xor U44974 (N_44974,N_43514,N_42860);
nand U44975 (N_44975,N_43618,N_43538);
nand U44976 (N_44976,N_42948,N_42230);
nor U44977 (N_44977,N_43011,N_43363);
xnor U44978 (N_44978,N_43422,N_42629);
nand U44979 (N_44979,N_43486,N_42820);
xnor U44980 (N_44980,N_42213,N_43821);
and U44981 (N_44981,N_43168,N_43353);
and U44982 (N_44982,N_42253,N_42393);
xor U44983 (N_44983,N_43578,N_43699);
nor U44984 (N_44984,N_43393,N_43277);
xor U44985 (N_44985,N_42256,N_43872);
and U44986 (N_44986,N_43418,N_43802);
or U44987 (N_44987,N_43403,N_43904);
nand U44988 (N_44988,N_42344,N_43397);
nand U44989 (N_44989,N_42068,N_43450);
or U44990 (N_44990,N_42494,N_43634);
nand U44991 (N_44991,N_42461,N_43306);
xnor U44992 (N_44992,N_43611,N_43736);
nand U44993 (N_44993,N_42530,N_42086);
or U44994 (N_44994,N_42308,N_43453);
and U44995 (N_44995,N_42690,N_42007);
nor U44996 (N_44996,N_42585,N_43884);
nor U44997 (N_44997,N_43169,N_43963);
nor U44998 (N_44998,N_42114,N_42809);
and U44999 (N_44999,N_42905,N_42096);
nand U45000 (N_45000,N_43342,N_43730);
and U45001 (N_45001,N_43598,N_42025);
or U45002 (N_45002,N_43722,N_42726);
xor U45003 (N_45003,N_42498,N_42005);
and U45004 (N_45004,N_42870,N_43266);
or U45005 (N_45005,N_43285,N_43354);
nor U45006 (N_45006,N_42996,N_42024);
nand U45007 (N_45007,N_43032,N_42966);
nand U45008 (N_45008,N_42486,N_43544);
and U45009 (N_45009,N_42709,N_43022);
and U45010 (N_45010,N_43586,N_42447);
and U45011 (N_45011,N_42332,N_42263);
and U45012 (N_45012,N_42020,N_42639);
or U45013 (N_45013,N_42326,N_43834);
or U45014 (N_45014,N_43391,N_42709);
nand U45015 (N_45015,N_42781,N_43849);
nor U45016 (N_45016,N_42315,N_43286);
nand U45017 (N_45017,N_43889,N_42366);
and U45018 (N_45018,N_42347,N_42115);
or U45019 (N_45019,N_42053,N_42280);
nand U45020 (N_45020,N_42950,N_43351);
nand U45021 (N_45021,N_43171,N_43718);
xnor U45022 (N_45022,N_42602,N_42532);
nand U45023 (N_45023,N_43734,N_43231);
xor U45024 (N_45024,N_42949,N_43447);
nor U45025 (N_45025,N_43260,N_43557);
xnor U45026 (N_45026,N_43411,N_42369);
nor U45027 (N_45027,N_43100,N_42103);
xor U45028 (N_45028,N_43083,N_43626);
nor U45029 (N_45029,N_42109,N_42595);
or U45030 (N_45030,N_42487,N_43001);
or U45031 (N_45031,N_42269,N_42921);
xnor U45032 (N_45032,N_42570,N_42131);
xnor U45033 (N_45033,N_42676,N_43216);
or U45034 (N_45034,N_42995,N_43284);
nand U45035 (N_45035,N_43565,N_43805);
nor U45036 (N_45036,N_43914,N_42725);
and U45037 (N_45037,N_43298,N_43356);
nor U45038 (N_45038,N_42120,N_43066);
or U45039 (N_45039,N_42915,N_43937);
xnor U45040 (N_45040,N_43295,N_42057);
or U45041 (N_45041,N_43640,N_42560);
or U45042 (N_45042,N_42587,N_43825);
or U45043 (N_45043,N_43521,N_43355);
xnor U45044 (N_45044,N_42865,N_42987);
and U45045 (N_45045,N_42601,N_42595);
nor U45046 (N_45046,N_42072,N_42085);
or U45047 (N_45047,N_42439,N_42016);
or U45048 (N_45048,N_43249,N_43247);
and U45049 (N_45049,N_43429,N_42054);
nand U45050 (N_45050,N_43682,N_43679);
nand U45051 (N_45051,N_42518,N_43502);
xnor U45052 (N_45052,N_42532,N_43644);
nor U45053 (N_45053,N_42360,N_42389);
nand U45054 (N_45054,N_42708,N_43037);
xnor U45055 (N_45055,N_42214,N_42978);
and U45056 (N_45056,N_43453,N_43098);
and U45057 (N_45057,N_42312,N_43984);
nor U45058 (N_45058,N_42879,N_43033);
or U45059 (N_45059,N_42922,N_43120);
xor U45060 (N_45060,N_42117,N_43883);
nor U45061 (N_45061,N_43720,N_43630);
nor U45062 (N_45062,N_43829,N_43315);
and U45063 (N_45063,N_42628,N_42276);
and U45064 (N_45064,N_43229,N_43389);
xor U45065 (N_45065,N_43176,N_42911);
or U45066 (N_45066,N_43990,N_43729);
or U45067 (N_45067,N_42647,N_42903);
and U45068 (N_45068,N_42756,N_42036);
nand U45069 (N_45069,N_42060,N_43618);
and U45070 (N_45070,N_43433,N_42389);
xor U45071 (N_45071,N_43774,N_43257);
and U45072 (N_45072,N_43379,N_42924);
and U45073 (N_45073,N_42887,N_42043);
and U45074 (N_45074,N_43425,N_43152);
and U45075 (N_45075,N_42557,N_43182);
and U45076 (N_45076,N_42905,N_42392);
xnor U45077 (N_45077,N_43097,N_43386);
nand U45078 (N_45078,N_43193,N_42289);
or U45079 (N_45079,N_42557,N_42419);
nor U45080 (N_45080,N_42169,N_42841);
xnor U45081 (N_45081,N_42113,N_42353);
xnor U45082 (N_45082,N_43911,N_42239);
or U45083 (N_45083,N_43933,N_42927);
nor U45084 (N_45084,N_43252,N_43479);
xor U45085 (N_45085,N_42712,N_43272);
or U45086 (N_45086,N_43306,N_42761);
xor U45087 (N_45087,N_43532,N_42455);
xnor U45088 (N_45088,N_42120,N_42169);
xnor U45089 (N_45089,N_42736,N_42334);
nand U45090 (N_45090,N_42438,N_43211);
and U45091 (N_45091,N_43681,N_43443);
nor U45092 (N_45092,N_43503,N_43766);
xnor U45093 (N_45093,N_43966,N_43936);
nand U45094 (N_45094,N_42643,N_42584);
xnor U45095 (N_45095,N_43547,N_42325);
nor U45096 (N_45096,N_43433,N_43856);
and U45097 (N_45097,N_43330,N_42194);
xor U45098 (N_45098,N_42334,N_43870);
or U45099 (N_45099,N_43567,N_43130);
xnor U45100 (N_45100,N_42174,N_42446);
and U45101 (N_45101,N_42845,N_42389);
or U45102 (N_45102,N_43155,N_43254);
xnor U45103 (N_45103,N_42933,N_42668);
nand U45104 (N_45104,N_42690,N_42624);
and U45105 (N_45105,N_43803,N_42115);
nor U45106 (N_45106,N_43254,N_43667);
and U45107 (N_45107,N_42524,N_43093);
nand U45108 (N_45108,N_43623,N_42390);
xor U45109 (N_45109,N_43480,N_43537);
nand U45110 (N_45110,N_43115,N_43491);
or U45111 (N_45111,N_42539,N_43896);
nor U45112 (N_45112,N_42448,N_42003);
and U45113 (N_45113,N_43320,N_43066);
xor U45114 (N_45114,N_42353,N_43891);
or U45115 (N_45115,N_43880,N_43475);
or U45116 (N_45116,N_43396,N_43803);
and U45117 (N_45117,N_42058,N_43563);
and U45118 (N_45118,N_43346,N_43577);
xor U45119 (N_45119,N_42475,N_43911);
nor U45120 (N_45120,N_43804,N_42580);
nor U45121 (N_45121,N_42055,N_43019);
nand U45122 (N_45122,N_43827,N_42279);
nor U45123 (N_45123,N_43590,N_43948);
nor U45124 (N_45124,N_43215,N_42745);
xnor U45125 (N_45125,N_43973,N_42002);
and U45126 (N_45126,N_42197,N_43998);
nor U45127 (N_45127,N_42659,N_42641);
nand U45128 (N_45128,N_43535,N_42167);
nand U45129 (N_45129,N_42931,N_42164);
xor U45130 (N_45130,N_43821,N_42092);
nor U45131 (N_45131,N_42051,N_42976);
xnor U45132 (N_45132,N_43992,N_42448);
nand U45133 (N_45133,N_43093,N_43920);
and U45134 (N_45134,N_42707,N_43089);
xor U45135 (N_45135,N_43401,N_43116);
nor U45136 (N_45136,N_43391,N_43658);
nand U45137 (N_45137,N_42212,N_43092);
nand U45138 (N_45138,N_43000,N_43595);
xor U45139 (N_45139,N_43075,N_42365);
or U45140 (N_45140,N_43273,N_42728);
nor U45141 (N_45141,N_43770,N_43782);
nor U45142 (N_45142,N_42604,N_43323);
nand U45143 (N_45143,N_42730,N_43503);
nor U45144 (N_45144,N_43294,N_42085);
xnor U45145 (N_45145,N_42395,N_42306);
or U45146 (N_45146,N_43561,N_42869);
and U45147 (N_45147,N_42708,N_43986);
xor U45148 (N_45148,N_42448,N_43793);
xnor U45149 (N_45149,N_42843,N_43828);
nand U45150 (N_45150,N_42490,N_43388);
or U45151 (N_45151,N_42275,N_43298);
or U45152 (N_45152,N_42709,N_43299);
xnor U45153 (N_45153,N_42877,N_42692);
nand U45154 (N_45154,N_42596,N_43248);
xnor U45155 (N_45155,N_43081,N_42395);
and U45156 (N_45156,N_43953,N_43779);
nor U45157 (N_45157,N_42333,N_42121);
and U45158 (N_45158,N_42670,N_43138);
nand U45159 (N_45159,N_42671,N_42941);
nor U45160 (N_45160,N_43750,N_42286);
nor U45161 (N_45161,N_43114,N_43290);
nor U45162 (N_45162,N_42237,N_42650);
xor U45163 (N_45163,N_42732,N_42020);
and U45164 (N_45164,N_43193,N_42092);
nor U45165 (N_45165,N_42473,N_43466);
nor U45166 (N_45166,N_43813,N_43466);
nand U45167 (N_45167,N_43813,N_43997);
nand U45168 (N_45168,N_43443,N_43239);
and U45169 (N_45169,N_42687,N_43534);
nor U45170 (N_45170,N_42902,N_42625);
and U45171 (N_45171,N_43866,N_42041);
and U45172 (N_45172,N_43779,N_43939);
or U45173 (N_45173,N_43917,N_42104);
or U45174 (N_45174,N_42295,N_42520);
nand U45175 (N_45175,N_42619,N_43991);
nor U45176 (N_45176,N_42203,N_43033);
or U45177 (N_45177,N_43641,N_43880);
xor U45178 (N_45178,N_42135,N_43530);
and U45179 (N_45179,N_42018,N_43576);
and U45180 (N_45180,N_42988,N_42358);
xnor U45181 (N_45181,N_43690,N_42812);
and U45182 (N_45182,N_43730,N_42426);
or U45183 (N_45183,N_43412,N_42188);
nand U45184 (N_45184,N_42940,N_42527);
nand U45185 (N_45185,N_42451,N_42298);
nor U45186 (N_45186,N_43483,N_42365);
nor U45187 (N_45187,N_43455,N_43134);
and U45188 (N_45188,N_43549,N_42304);
or U45189 (N_45189,N_43417,N_43793);
and U45190 (N_45190,N_42569,N_42124);
xnor U45191 (N_45191,N_43400,N_42232);
nand U45192 (N_45192,N_43624,N_43663);
nor U45193 (N_45193,N_42017,N_43550);
nand U45194 (N_45194,N_42502,N_43793);
and U45195 (N_45195,N_42946,N_42491);
nor U45196 (N_45196,N_43577,N_43780);
nor U45197 (N_45197,N_42729,N_42443);
nand U45198 (N_45198,N_42633,N_43120);
or U45199 (N_45199,N_43960,N_42973);
nor U45200 (N_45200,N_43135,N_43998);
xor U45201 (N_45201,N_43398,N_42829);
or U45202 (N_45202,N_43307,N_43187);
nor U45203 (N_45203,N_43152,N_42527);
xor U45204 (N_45204,N_42304,N_42323);
and U45205 (N_45205,N_42224,N_42380);
and U45206 (N_45206,N_43528,N_42337);
xnor U45207 (N_45207,N_43028,N_43119);
nand U45208 (N_45208,N_42807,N_42914);
nand U45209 (N_45209,N_42135,N_42046);
or U45210 (N_45210,N_42857,N_42095);
or U45211 (N_45211,N_42369,N_42990);
nand U45212 (N_45212,N_42971,N_43994);
xor U45213 (N_45213,N_42531,N_43103);
or U45214 (N_45214,N_43909,N_42765);
nor U45215 (N_45215,N_43585,N_43706);
nand U45216 (N_45216,N_43742,N_42109);
or U45217 (N_45217,N_42878,N_42266);
xor U45218 (N_45218,N_43542,N_43353);
xnor U45219 (N_45219,N_42664,N_43877);
or U45220 (N_45220,N_42860,N_43984);
and U45221 (N_45221,N_42631,N_42164);
nor U45222 (N_45222,N_42757,N_43364);
nor U45223 (N_45223,N_43192,N_42637);
xor U45224 (N_45224,N_42173,N_43200);
or U45225 (N_45225,N_42928,N_42095);
and U45226 (N_45226,N_43009,N_43277);
and U45227 (N_45227,N_42986,N_42138);
xnor U45228 (N_45228,N_43656,N_43124);
xnor U45229 (N_45229,N_42008,N_42356);
nand U45230 (N_45230,N_43458,N_42199);
and U45231 (N_45231,N_43389,N_43165);
or U45232 (N_45232,N_43824,N_42935);
or U45233 (N_45233,N_42157,N_42617);
xnor U45234 (N_45234,N_42925,N_43790);
or U45235 (N_45235,N_43517,N_43048);
xnor U45236 (N_45236,N_43060,N_42708);
nor U45237 (N_45237,N_43652,N_43587);
nand U45238 (N_45238,N_43499,N_43597);
nand U45239 (N_45239,N_42042,N_42397);
and U45240 (N_45240,N_43598,N_42266);
nor U45241 (N_45241,N_43573,N_42440);
xnor U45242 (N_45242,N_43276,N_43119);
and U45243 (N_45243,N_42372,N_43232);
and U45244 (N_45244,N_43215,N_43846);
or U45245 (N_45245,N_42076,N_42978);
nor U45246 (N_45246,N_42167,N_42717);
xor U45247 (N_45247,N_43632,N_43595);
xor U45248 (N_45248,N_43893,N_43148);
nand U45249 (N_45249,N_43122,N_42514);
xor U45250 (N_45250,N_42145,N_43802);
and U45251 (N_45251,N_43552,N_42613);
or U45252 (N_45252,N_43571,N_42712);
and U45253 (N_45253,N_43015,N_42374);
or U45254 (N_45254,N_42634,N_42149);
and U45255 (N_45255,N_43121,N_42474);
or U45256 (N_45256,N_42716,N_42348);
or U45257 (N_45257,N_43219,N_42180);
and U45258 (N_45258,N_42233,N_43991);
xor U45259 (N_45259,N_42801,N_43772);
xnor U45260 (N_45260,N_42798,N_42401);
and U45261 (N_45261,N_43845,N_42524);
or U45262 (N_45262,N_43353,N_43935);
or U45263 (N_45263,N_42597,N_43639);
and U45264 (N_45264,N_42720,N_43258);
xor U45265 (N_45265,N_42034,N_43216);
nand U45266 (N_45266,N_42208,N_43242);
nand U45267 (N_45267,N_43747,N_42808);
xor U45268 (N_45268,N_42033,N_42086);
xor U45269 (N_45269,N_42306,N_43488);
and U45270 (N_45270,N_42523,N_42664);
nand U45271 (N_45271,N_43399,N_42254);
xor U45272 (N_45272,N_42152,N_42492);
and U45273 (N_45273,N_42226,N_42423);
or U45274 (N_45274,N_42427,N_42038);
nor U45275 (N_45275,N_43084,N_43017);
or U45276 (N_45276,N_42474,N_43873);
and U45277 (N_45277,N_43049,N_43002);
xnor U45278 (N_45278,N_42599,N_42559);
and U45279 (N_45279,N_43475,N_43087);
nand U45280 (N_45280,N_42274,N_43722);
xor U45281 (N_45281,N_42550,N_43131);
and U45282 (N_45282,N_43426,N_43692);
or U45283 (N_45283,N_42579,N_43471);
xnor U45284 (N_45284,N_43260,N_43677);
or U45285 (N_45285,N_43816,N_43533);
nor U45286 (N_45286,N_43603,N_43845);
or U45287 (N_45287,N_42633,N_42769);
or U45288 (N_45288,N_42341,N_43788);
nor U45289 (N_45289,N_42279,N_42946);
and U45290 (N_45290,N_42507,N_42060);
nor U45291 (N_45291,N_42663,N_42046);
and U45292 (N_45292,N_42185,N_42079);
or U45293 (N_45293,N_42954,N_43964);
nor U45294 (N_45294,N_43468,N_42571);
or U45295 (N_45295,N_42593,N_43138);
nand U45296 (N_45296,N_43248,N_42876);
or U45297 (N_45297,N_43319,N_42717);
or U45298 (N_45298,N_42837,N_43064);
nor U45299 (N_45299,N_43200,N_42685);
nor U45300 (N_45300,N_42106,N_43805);
or U45301 (N_45301,N_42730,N_42450);
nor U45302 (N_45302,N_43716,N_43500);
xor U45303 (N_45303,N_42148,N_43113);
xor U45304 (N_45304,N_43283,N_42267);
nor U45305 (N_45305,N_43531,N_43105);
and U45306 (N_45306,N_43831,N_43879);
xnor U45307 (N_45307,N_42355,N_43224);
or U45308 (N_45308,N_43952,N_42523);
xnor U45309 (N_45309,N_43215,N_42123);
and U45310 (N_45310,N_43467,N_43003);
nor U45311 (N_45311,N_42229,N_43345);
nor U45312 (N_45312,N_42640,N_42459);
xnor U45313 (N_45313,N_43686,N_42531);
xnor U45314 (N_45314,N_43199,N_43853);
xor U45315 (N_45315,N_43515,N_43791);
and U45316 (N_45316,N_42693,N_43480);
nor U45317 (N_45317,N_42954,N_43841);
nor U45318 (N_45318,N_42736,N_42794);
nand U45319 (N_45319,N_42465,N_42456);
and U45320 (N_45320,N_43808,N_42317);
xor U45321 (N_45321,N_42099,N_42868);
nand U45322 (N_45322,N_42478,N_42265);
nand U45323 (N_45323,N_43707,N_42882);
nand U45324 (N_45324,N_43671,N_43973);
xnor U45325 (N_45325,N_42521,N_42168);
and U45326 (N_45326,N_42546,N_43965);
nand U45327 (N_45327,N_43622,N_42993);
and U45328 (N_45328,N_43669,N_43322);
nor U45329 (N_45329,N_42280,N_42036);
or U45330 (N_45330,N_43089,N_43484);
and U45331 (N_45331,N_43705,N_42481);
and U45332 (N_45332,N_43767,N_43551);
or U45333 (N_45333,N_42027,N_43453);
xor U45334 (N_45334,N_43292,N_43861);
and U45335 (N_45335,N_42064,N_42724);
xor U45336 (N_45336,N_42219,N_43409);
or U45337 (N_45337,N_43517,N_42233);
and U45338 (N_45338,N_43558,N_42224);
and U45339 (N_45339,N_42364,N_43150);
nand U45340 (N_45340,N_42866,N_43448);
nor U45341 (N_45341,N_43172,N_42268);
nand U45342 (N_45342,N_42956,N_43813);
nand U45343 (N_45343,N_42747,N_42830);
nor U45344 (N_45344,N_43394,N_42821);
nor U45345 (N_45345,N_42326,N_43838);
nand U45346 (N_45346,N_43660,N_42886);
nor U45347 (N_45347,N_43554,N_42846);
nor U45348 (N_45348,N_43811,N_43037);
nand U45349 (N_45349,N_43530,N_43130);
or U45350 (N_45350,N_43946,N_43091);
nor U45351 (N_45351,N_43628,N_43688);
nor U45352 (N_45352,N_42077,N_43123);
xor U45353 (N_45353,N_43028,N_43959);
xor U45354 (N_45354,N_42877,N_42147);
xnor U45355 (N_45355,N_42429,N_43871);
nor U45356 (N_45356,N_43749,N_42589);
and U45357 (N_45357,N_42606,N_43922);
nor U45358 (N_45358,N_42891,N_43784);
nor U45359 (N_45359,N_42733,N_43862);
nor U45360 (N_45360,N_42156,N_42380);
or U45361 (N_45361,N_42404,N_43662);
xor U45362 (N_45362,N_42769,N_43706);
nand U45363 (N_45363,N_42663,N_43546);
xnor U45364 (N_45364,N_42716,N_42330);
xnor U45365 (N_45365,N_43433,N_43496);
xor U45366 (N_45366,N_42395,N_43626);
xor U45367 (N_45367,N_42423,N_43194);
xor U45368 (N_45368,N_42441,N_42260);
and U45369 (N_45369,N_42108,N_43624);
and U45370 (N_45370,N_43373,N_43267);
and U45371 (N_45371,N_42463,N_43051);
xor U45372 (N_45372,N_42385,N_43390);
or U45373 (N_45373,N_42935,N_42014);
xnor U45374 (N_45374,N_42219,N_43525);
xor U45375 (N_45375,N_42499,N_43675);
nand U45376 (N_45376,N_43110,N_42880);
nor U45377 (N_45377,N_43049,N_42597);
or U45378 (N_45378,N_42886,N_43726);
and U45379 (N_45379,N_43442,N_43248);
nand U45380 (N_45380,N_43422,N_42447);
nor U45381 (N_45381,N_42176,N_43755);
or U45382 (N_45382,N_43422,N_42199);
nor U45383 (N_45383,N_42357,N_43306);
or U45384 (N_45384,N_43283,N_42741);
or U45385 (N_45385,N_42714,N_43274);
nand U45386 (N_45386,N_42074,N_42324);
and U45387 (N_45387,N_42550,N_42011);
nand U45388 (N_45388,N_43719,N_42093);
or U45389 (N_45389,N_43221,N_43287);
nand U45390 (N_45390,N_42950,N_43239);
xor U45391 (N_45391,N_43954,N_43985);
xnor U45392 (N_45392,N_43672,N_42587);
nand U45393 (N_45393,N_43228,N_43488);
xor U45394 (N_45394,N_43885,N_42230);
nand U45395 (N_45395,N_42937,N_43247);
xor U45396 (N_45396,N_42334,N_43196);
and U45397 (N_45397,N_42569,N_42242);
nand U45398 (N_45398,N_43936,N_42681);
nor U45399 (N_45399,N_42033,N_43555);
nand U45400 (N_45400,N_42198,N_42629);
nand U45401 (N_45401,N_42490,N_42200);
or U45402 (N_45402,N_42254,N_43805);
xor U45403 (N_45403,N_42421,N_43622);
and U45404 (N_45404,N_43415,N_42265);
nand U45405 (N_45405,N_42069,N_42685);
xnor U45406 (N_45406,N_42709,N_42534);
nand U45407 (N_45407,N_42251,N_42234);
nor U45408 (N_45408,N_42186,N_43842);
nor U45409 (N_45409,N_43223,N_42500);
nand U45410 (N_45410,N_42852,N_42769);
and U45411 (N_45411,N_42282,N_42345);
nor U45412 (N_45412,N_42927,N_43096);
and U45413 (N_45413,N_43925,N_42834);
and U45414 (N_45414,N_42295,N_43631);
nor U45415 (N_45415,N_42247,N_43210);
xor U45416 (N_45416,N_43282,N_43681);
nor U45417 (N_45417,N_43345,N_43698);
xor U45418 (N_45418,N_43398,N_42490);
or U45419 (N_45419,N_42176,N_43505);
or U45420 (N_45420,N_43682,N_43012);
nor U45421 (N_45421,N_43931,N_43950);
or U45422 (N_45422,N_43719,N_43755);
xor U45423 (N_45423,N_43248,N_43951);
nand U45424 (N_45424,N_43206,N_43234);
nand U45425 (N_45425,N_42421,N_42140);
or U45426 (N_45426,N_42307,N_42253);
and U45427 (N_45427,N_43739,N_43864);
nor U45428 (N_45428,N_43063,N_42381);
nand U45429 (N_45429,N_42791,N_42164);
xnor U45430 (N_45430,N_43180,N_42056);
or U45431 (N_45431,N_42723,N_42656);
nand U45432 (N_45432,N_42668,N_42334);
or U45433 (N_45433,N_42832,N_43516);
and U45434 (N_45434,N_43695,N_43748);
nor U45435 (N_45435,N_43823,N_42553);
xor U45436 (N_45436,N_42570,N_43986);
nor U45437 (N_45437,N_42449,N_43331);
or U45438 (N_45438,N_43019,N_42832);
nand U45439 (N_45439,N_42848,N_42079);
nand U45440 (N_45440,N_43900,N_43305);
xnor U45441 (N_45441,N_43725,N_42435);
nor U45442 (N_45442,N_43862,N_43221);
and U45443 (N_45443,N_42365,N_43737);
nor U45444 (N_45444,N_43677,N_43284);
and U45445 (N_45445,N_43254,N_43393);
nand U45446 (N_45446,N_42315,N_42196);
nor U45447 (N_45447,N_43299,N_43990);
or U45448 (N_45448,N_43118,N_43820);
nor U45449 (N_45449,N_43217,N_42174);
and U45450 (N_45450,N_43444,N_43669);
nor U45451 (N_45451,N_42301,N_43267);
or U45452 (N_45452,N_42716,N_43519);
and U45453 (N_45453,N_42383,N_43929);
nand U45454 (N_45454,N_42824,N_42846);
and U45455 (N_45455,N_42480,N_43064);
nor U45456 (N_45456,N_43222,N_42974);
or U45457 (N_45457,N_43421,N_43765);
and U45458 (N_45458,N_42343,N_42775);
nor U45459 (N_45459,N_42964,N_43034);
or U45460 (N_45460,N_43571,N_42296);
nor U45461 (N_45461,N_43116,N_43441);
nor U45462 (N_45462,N_43267,N_42800);
and U45463 (N_45463,N_43049,N_43540);
xnor U45464 (N_45464,N_42656,N_42705);
or U45465 (N_45465,N_42863,N_42073);
nor U45466 (N_45466,N_42168,N_43074);
and U45467 (N_45467,N_42200,N_43144);
nand U45468 (N_45468,N_42573,N_42433);
and U45469 (N_45469,N_43303,N_42685);
nor U45470 (N_45470,N_42438,N_43297);
or U45471 (N_45471,N_43985,N_43232);
nand U45472 (N_45472,N_43376,N_43976);
or U45473 (N_45473,N_42385,N_42400);
nand U45474 (N_45474,N_43216,N_42973);
nor U45475 (N_45475,N_42412,N_42208);
nor U45476 (N_45476,N_42866,N_42766);
or U45477 (N_45477,N_42053,N_43649);
xnor U45478 (N_45478,N_42971,N_42545);
nor U45479 (N_45479,N_43501,N_42324);
nand U45480 (N_45480,N_42979,N_42926);
and U45481 (N_45481,N_43742,N_43136);
xor U45482 (N_45482,N_42356,N_43860);
xnor U45483 (N_45483,N_43312,N_43239);
and U45484 (N_45484,N_43761,N_43193);
nor U45485 (N_45485,N_42209,N_43437);
xnor U45486 (N_45486,N_43805,N_42684);
nand U45487 (N_45487,N_42710,N_42141);
or U45488 (N_45488,N_42999,N_43903);
nor U45489 (N_45489,N_43563,N_42138);
nor U45490 (N_45490,N_42114,N_43272);
or U45491 (N_45491,N_42160,N_43893);
nor U45492 (N_45492,N_42192,N_43416);
or U45493 (N_45493,N_42121,N_42937);
or U45494 (N_45494,N_43374,N_42909);
and U45495 (N_45495,N_42957,N_42687);
xnor U45496 (N_45496,N_43164,N_42693);
nand U45497 (N_45497,N_43865,N_42652);
nand U45498 (N_45498,N_43219,N_42848);
nor U45499 (N_45499,N_42622,N_42100);
xnor U45500 (N_45500,N_43892,N_42965);
nand U45501 (N_45501,N_43926,N_42069);
or U45502 (N_45502,N_42332,N_42392);
nand U45503 (N_45503,N_43735,N_42188);
or U45504 (N_45504,N_43418,N_43878);
nor U45505 (N_45505,N_43417,N_43192);
xor U45506 (N_45506,N_43351,N_43920);
nor U45507 (N_45507,N_43826,N_42227);
nand U45508 (N_45508,N_42425,N_43216);
nand U45509 (N_45509,N_43874,N_43002);
and U45510 (N_45510,N_43065,N_43835);
xnor U45511 (N_45511,N_42853,N_43223);
and U45512 (N_45512,N_43744,N_42494);
or U45513 (N_45513,N_42555,N_43195);
xnor U45514 (N_45514,N_43910,N_43434);
xor U45515 (N_45515,N_43283,N_42102);
or U45516 (N_45516,N_43945,N_42884);
and U45517 (N_45517,N_43445,N_43008);
and U45518 (N_45518,N_42876,N_42044);
and U45519 (N_45519,N_42987,N_42738);
xor U45520 (N_45520,N_42127,N_43636);
or U45521 (N_45521,N_43723,N_42626);
nor U45522 (N_45522,N_42380,N_42438);
nor U45523 (N_45523,N_42650,N_42689);
xor U45524 (N_45524,N_42878,N_42320);
and U45525 (N_45525,N_42448,N_42738);
xor U45526 (N_45526,N_42029,N_43408);
or U45527 (N_45527,N_43402,N_43835);
xnor U45528 (N_45528,N_43224,N_43270);
xnor U45529 (N_45529,N_42219,N_43216);
and U45530 (N_45530,N_43039,N_43367);
or U45531 (N_45531,N_43977,N_42892);
and U45532 (N_45532,N_42108,N_42158);
nand U45533 (N_45533,N_43945,N_42369);
and U45534 (N_45534,N_43127,N_43033);
or U45535 (N_45535,N_43534,N_42088);
and U45536 (N_45536,N_42856,N_43328);
nand U45537 (N_45537,N_43047,N_42275);
xnor U45538 (N_45538,N_43780,N_42510);
xnor U45539 (N_45539,N_42000,N_43827);
nand U45540 (N_45540,N_43316,N_42973);
nand U45541 (N_45541,N_42261,N_43249);
xor U45542 (N_45542,N_43729,N_42465);
xor U45543 (N_45543,N_42562,N_43523);
xnor U45544 (N_45544,N_43711,N_42592);
or U45545 (N_45545,N_43585,N_42908);
and U45546 (N_45546,N_43741,N_43716);
xnor U45547 (N_45547,N_42219,N_43504);
and U45548 (N_45548,N_42953,N_43779);
nand U45549 (N_45549,N_42962,N_42222);
or U45550 (N_45550,N_43427,N_43734);
and U45551 (N_45551,N_43687,N_43812);
xor U45552 (N_45552,N_43410,N_42402);
nand U45553 (N_45553,N_43365,N_43507);
xor U45554 (N_45554,N_43230,N_43810);
nand U45555 (N_45555,N_43171,N_43089);
nor U45556 (N_45556,N_42328,N_42538);
nor U45557 (N_45557,N_42976,N_43187);
xor U45558 (N_45558,N_43799,N_43532);
xnor U45559 (N_45559,N_42454,N_42924);
nor U45560 (N_45560,N_43793,N_43798);
nand U45561 (N_45561,N_42945,N_42984);
nand U45562 (N_45562,N_42176,N_43800);
nand U45563 (N_45563,N_42291,N_43542);
xor U45564 (N_45564,N_43258,N_42125);
and U45565 (N_45565,N_42051,N_42090);
and U45566 (N_45566,N_42327,N_43815);
and U45567 (N_45567,N_42695,N_42677);
xor U45568 (N_45568,N_43658,N_42711);
nor U45569 (N_45569,N_43893,N_42044);
and U45570 (N_45570,N_42323,N_43769);
or U45571 (N_45571,N_42255,N_42115);
and U45572 (N_45572,N_43651,N_42206);
xnor U45573 (N_45573,N_43528,N_42110);
or U45574 (N_45574,N_42736,N_43942);
or U45575 (N_45575,N_42068,N_43537);
nand U45576 (N_45576,N_42244,N_42908);
nor U45577 (N_45577,N_42713,N_43443);
nand U45578 (N_45578,N_42936,N_42038);
and U45579 (N_45579,N_43938,N_42245);
or U45580 (N_45580,N_43979,N_43068);
or U45581 (N_45581,N_42366,N_42028);
nor U45582 (N_45582,N_42497,N_43482);
nor U45583 (N_45583,N_43942,N_43821);
xor U45584 (N_45584,N_43178,N_43380);
nand U45585 (N_45585,N_43120,N_42765);
and U45586 (N_45586,N_42847,N_43867);
xnor U45587 (N_45587,N_42154,N_43333);
nand U45588 (N_45588,N_43189,N_42088);
xnor U45589 (N_45589,N_43340,N_43507);
and U45590 (N_45590,N_43794,N_42417);
nand U45591 (N_45591,N_42692,N_43793);
xnor U45592 (N_45592,N_43578,N_43714);
xor U45593 (N_45593,N_43195,N_42821);
and U45594 (N_45594,N_42443,N_43227);
and U45595 (N_45595,N_42365,N_42061);
nand U45596 (N_45596,N_42381,N_42179);
xnor U45597 (N_45597,N_43910,N_43783);
nor U45598 (N_45598,N_42932,N_42839);
xor U45599 (N_45599,N_42790,N_43187);
xnor U45600 (N_45600,N_43760,N_42170);
xnor U45601 (N_45601,N_42318,N_42224);
xnor U45602 (N_45602,N_42503,N_42241);
nor U45603 (N_45603,N_43489,N_43886);
nand U45604 (N_45604,N_42152,N_42672);
nand U45605 (N_45605,N_42256,N_43963);
or U45606 (N_45606,N_43117,N_43310);
xor U45607 (N_45607,N_43978,N_43304);
and U45608 (N_45608,N_43673,N_42867);
nor U45609 (N_45609,N_43760,N_42737);
nand U45610 (N_45610,N_42790,N_43723);
nor U45611 (N_45611,N_42542,N_43541);
nor U45612 (N_45612,N_42199,N_42313);
nand U45613 (N_45613,N_43275,N_43693);
nor U45614 (N_45614,N_42452,N_43358);
xnor U45615 (N_45615,N_42169,N_43153);
nor U45616 (N_45616,N_42566,N_42798);
nor U45617 (N_45617,N_42766,N_43182);
xnor U45618 (N_45618,N_42167,N_42031);
or U45619 (N_45619,N_43923,N_42923);
nor U45620 (N_45620,N_43737,N_43945);
xor U45621 (N_45621,N_42491,N_42996);
and U45622 (N_45622,N_43172,N_43621);
xor U45623 (N_45623,N_43244,N_43839);
nor U45624 (N_45624,N_42026,N_42849);
nand U45625 (N_45625,N_42728,N_42060);
nand U45626 (N_45626,N_42247,N_42312);
and U45627 (N_45627,N_42621,N_42622);
or U45628 (N_45628,N_42725,N_42745);
nor U45629 (N_45629,N_42677,N_42889);
and U45630 (N_45630,N_42831,N_43759);
nor U45631 (N_45631,N_42996,N_43634);
and U45632 (N_45632,N_42356,N_43463);
nand U45633 (N_45633,N_43250,N_42162);
or U45634 (N_45634,N_43211,N_42274);
and U45635 (N_45635,N_43520,N_43490);
nand U45636 (N_45636,N_42778,N_42613);
xnor U45637 (N_45637,N_43094,N_43741);
nand U45638 (N_45638,N_43684,N_43734);
xor U45639 (N_45639,N_43285,N_43475);
nor U45640 (N_45640,N_43951,N_42644);
or U45641 (N_45641,N_42804,N_42430);
nand U45642 (N_45642,N_43193,N_42087);
xor U45643 (N_45643,N_42889,N_43315);
nor U45644 (N_45644,N_42716,N_43931);
nor U45645 (N_45645,N_42890,N_43485);
nand U45646 (N_45646,N_42823,N_42117);
nor U45647 (N_45647,N_43403,N_43388);
xnor U45648 (N_45648,N_42399,N_43288);
and U45649 (N_45649,N_43989,N_42926);
nand U45650 (N_45650,N_42050,N_43562);
nand U45651 (N_45651,N_42184,N_43745);
xor U45652 (N_45652,N_43515,N_43655);
nand U45653 (N_45653,N_43788,N_42103);
or U45654 (N_45654,N_43081,N_42677);
nor U45655 (N_45655,N_43122,N_43699);
or U45656 (N_45656,N_43759,N_42693);
and U45657 (N_45657,N_43287,N_42575);
xnor U45658 (N_45658,N_43568,N_42000);
nor U45659 (N_45659,N_43996,N_42838);
xnor U45660 (N_45660,N_42233,N_43798);
xnor U45661 (N_45661,N_42553,N_42533);
xnor U45662 (N_45662,N_42340,N_43420);
nor U45663 (N_45663,N_43731,N_42418);
nand U45664 (N_45664,N_42304,N_42161);
and U45665 (N_45665,N_43408,N_43270);
and U45666 (N_45666,N_43992,N_42408);
or U45667 (N_45667,N_42685,N_42122);
nor U45668 (N_45668,N_42615,N_42706);
nand U45669 (N_45669,N_42524,N_43456);
nand U45670 (N_45670,N_42350,N_42614);
or U45671 (N_45671,N_42577,N_42692);
nor U45672 (N_45672,N_43642,N_43716);
or U45673 (N_45673,N_42826,N_43023);
nand U45674 (N_45674,N_42851,N_42161);
and U45675 (N_45675,N_42160,N_43707);
xor U45676 (N_45676,N_42452,N_42426);
nand U45677 (N_45677,N_43770,N_42746);
nor U45678 (N_45678,N_43514,N_42312);
xnor U45679 (N_45679,N_42981,N_43763);
nor U45680 (N_45680,N_42283,N_42950);
or U45681 (N_45681,N_42355,N_43856);
nor U45682 (N_45682,N_43899,N_42695);
and U45683 (N_45683,N_42547,N_42483);
nand U45684 (N_45684,N_42747,N_43824);
nand U45685 (N_45685,N_42951,N_42549);
and U45686 (N_45686,N_42544,N_42706);
xnor U45687 (N_45687,N_42280,N_42049);
and U45688 (N_45688,N_43766,N_43574);
and U45689 (N_45689,N_42135,N_43621);
xnor U45690 (N_45690,N_43304,N_42396);
and U45691 (N_45691,N_42253,N_43335);
and U45692 (N_45692,N_43412,N_42139);
nand U45693 (N_45693,N_43428,N_43275);
nand U45694 (N_45694,N_43908,N_43883);
xnor U45695 (N_45695,N_43787,N_42909);
or U45696 (N_45696,N_42083,N_42397);
xnor U45697 (N_45697,N_42443,N_42552);
xnor U45698 (N_45698,N_42048,N_43438);
xor U45699 (N_45699,N_43658,N_42094);
or U45700 (N_45700,N_42802,N_43475);
or U45701 (N_45701,N_43986,N_42303);
xor U45702 (N_45702,N_43689,N_42387);
nor U45703 (N_45703,N_42049,N_43378);
nand U45704 (N_45704,N_43930,N_42882);
or U45705 (N_45705,N_43606,N_42812);
xnor U45706 (N_45706,N_42274,N_43904);
nand U45707 (N_45707,N_43396,N_43818);
and U45708 (N_45708,N_43485,N_42073);
nor U45709 (N_45709,N_43898,N_42773);
or U45710 (N_45710,N_43753,N_43267);
xor U45711 (N_45711,N_43593,N_43456);
xor U45712 (N_45712,N_42803,N_43226);
nor U45713 (N_45713,N_42016,N_42749);
xnor U45714 (N_45714,N_43157,N_43999);
nand U45715 (N_45715,N_43198,N_43362);
nand U45716 (N_45716,N_42910,N_42005);
nor U45717 (N_45717,N_43437,N_42772);
xor U45718 (N_45718,N_43691,N_42471);
xnor U45719 (N_45719,N_42702,N_42431);
or U45720 (N_45720,N_42268,N_42976);
nand U45721 (N_45721,N_43652,N_42648);
or U45722 (N_45722,N_42396,N_43400);
and U45723 (N_45723,N_43624,N_43656);
and U45724 (N_45724,N_42806,N_43418);
nor U45725 (N_45725,N_43321,N_43723);
or U45726 (N_45726,N_42188,N_42370);
nand U45727 (N_45727,N_42778,N_42229);
nand U45728 (N_45728,N_43200,N_42497);
or U45729 (N_45729,N_42708,N_42373);
nand U45730 (N_45730,N_43042,N_43843);
nor U45731 (N_45731,N_42601,N_42461);
nand U45732 (N_45732,N_42834,N_42912);
nor U45733 (N_45733,N_43511,N_43753);
xor U45734 (N_45734,N_42975,N_42361);
nand U45735 (N_45735,N_42294,N_43424);
or U45736 (N_45736,N_42778,N_42722);
nand U45737 (N_45737,N_42064,N_43700);
nand U45738 (N_45738,N_43577,N_42744);
or U45739 (N_45739,N_43627,N_42493);
or U45740 (N_45740,N_42550,N_42333);
and U45741 (N_45741,N_43307,N_43055);
or U45742 (N_45742,N_42475,N_42255);
and U45743 (N_45743,N_42056,N_43470);
nand U45744 (N_45744,N_43013,N_42011);
and U45745 (N_45745,N_42331,N_43520);
and U45746 (N_45746,N_43083,N_42879);
or U45747 (N_45747,N_42929,N_43974);
nand U45748 (N_45748,N_43018,N_43659);
and U45749 (N_45749,N_43721,N_42166);
and U45750 (N_45750,N_42284,N_42137);
and U45751 (N_45751,N_43388,N_42145);
xor U45752 (N_45752,N_42796,N_42736);
nor U45753 (N_45753,N_43340,N_43210);
xnor U45754 (N_45754,N_43301,N_42152);
nor U45755 (N_45755,N_42331,N_43701);
nor U45756 (N_45756,N_43760,N_42645);
xnor U45757 (N_45757,N_42855,N_43398);
or U45758 (N_45758,N_42215,N_43480);
xor U45759 (N_45759,N_42989,N_43056);
nor U45760 (N_45760,N_43653,N_43942);
xor U45761 (N_45761,N_42259,N_43501);
nand U45762 (N_45762,N_43103,N_43928);
nor U45763 (N_45763,N_42907,N_43886);
nand U45764 (N_45764,N_43161,N_43468);
nand U45765 (N_45765,N_43406,N_43034);
nand U45766 (N_45766,N_43863,N_43979);
nor U45767 (N_45767,N_42488,N_42666);
nor U45768 (N_45768,N_42582,N_42288);
nor U45769 (N_45769,N_43172,N_43148);
nand U45770 (N_45770,N_42333,N_43312);
nor U45771 (N_45771,N_42123,N_43942);
nor U45772 (N_45772,N_43836,N_43966);
or U45773 (N_45773,N_43057,N_42323);
nor U45774 (N_45774,N_42165,N_42251);
xor U45775 (N_45775,N_42863,N_43156);
nor U45776 (N_45776,N_42395,N_42534);
nor U45777 (N_45777,N_42449,N_42395);
nor U45778 (N_45778,N_43984,N_42335);
nor U45779 (N_45779,N_42192,N_42942);
or U45780 (N_45780,N_43855,N_43026);
and U45781 (N_45781,N_43714,N_42138);
nor U45782 (N_45782,N_43128,N_43903);
nand U45783 (N_45783,N_42563,N_42266);
nand U45784 (N_45784,N_42974,N_43019);
and U45785 (N_45785,N_42602,N_42642);
or U45786 (N_45786,N_42499,N_42530);
nand U45787 (N_45787,N_42918,N_43745);
xor U45788 (N_45788,N_42549,N_43515);
xor U45789 (N_45789,N_42357,N_42847);
nor U45790 (N_45790,N_42572,N_43010);
and U45791 (N_45791,N_43566,N_42265);
xnor U45792 (N_45792,N_42084,N_43005);
or U45793 (N_45793,N_43684,N_43070);
and U45794 (N_45794,N_43377,N_43879);
and U45795 (N_45795,N_42554,N_42154);
and U45796 (N_45796,N_42721,N_43096);
nor U45797 (N_45797,N_43200,N_43764);
xnor U45798 (N_45798,N_42089,N_42984);
or U45799 (N_45799,N_43078,N_42562);
xor U45800 (N_45800,N_43621,N_42772);
nand U45801 (N_45801,N_42098,N_42103);
or U45802 (N_45802,N_42302,N_43440);
xnor U45803 (N_45803,N_42622,N_42609);
or U45804 (N_45804,N_42036,N_42260);
and U45805 (N_45805,N_43458,N_42941);
nand U45806 (N_45806,N_42451,N_43963);
and U45807 (N_45807,N_42345,N_42922);
and U45808 (N_45808,N_42558,N_42418);
nor U45809 (N_45809,N_42041,N_43074);
xnor U45810 (N_45810,N_43622,N_43821);
nand U45811 (N_45811,N_43139,N_43644);
or U45812 (N_45812,N_42782,N_43369);
or U45813 (N_45813,N_42781,N_43382);
nand U45814 (N_45814,N_43256,N_43194);
and U45815 (N_45815,N_42142,N_42289);
nand U45816 (N_45816,N_42669,N_42736);
xor U45817 (N_45817,N_42454,N_42944);
nand U45818 (N_45818,N_43486,N_42392);
xor U45819 (N_45819,N_42026,N_42503);
and U45820 (N_45820,N_42425,N_42766);
and U45821 (N_45821,N_42606,N_43580);
and U45822 (N_45822,N_43936,N_42817);
nor U45823 (N_45823,N_42829,N_43049);
nand U45824 (N_45824,N_43173,N_42967);
nand U45825 (N_45825,N_42261,N_42428);
or U45826 (N_45826,N_43132,N_42297);
xor U45827 (N_45827,N_42168,N_42780);
xnor U45828 (N_45828,N_42024,N_42921);
and U45829 (N_45829,N_43921,N_43313);
and U45830 (N_45830,N_42587,N_43613);
nor U45831 (N_45831,N_43813,N_42885);
or U45832 (N_45832,N_42125,N_43789);
nand U45833 (N_45833,N_42444,N_43963);
xnor U45834 (N_45834,N_42838,N_42282);
nand U45835 (N_45835,N_42552,N_42676);
nand U45836 (N_45836,N_43679,N_42404);
xor U45837 (N_45837,N_43465,N_42905);
nor U45838 (N_45838,N_43423,N_42300);
and U45839 (N_45839,N_42435,N_42706);
or U45840 (N_45840,N_43861,N_43705);
or U45841 (N_45841,N_43888,N_43304);
xor U45842 (N_45842,N_42440,N_43528);
or U45843 (N_45843,N_43813,N_43745);
and U45844 (N_45844,N_43366,N_43333);
and U45845 (N_45845,N_43054,N_43999);
and U45846 (N_45846,N_42033,N_42316);
and U45847 (N_45847,N_43999,N_42080);
and U45848 (N_45848,N_42632,N_42605);
and U45849 (N_45849,N_42443,N_43335);
xnor U45850 (N_45850,N_42472,N_42967);
nor U45851 (N_45851,N_43318,N_43884);
nand U45852 (N_45852,N_43738,N_42544);
nor U45853 (N_45853,N_43576,N_43602);
or U45854 (N_45854,N_42743,N_42322);
xor U45855 (N_45855,N_43171,N_43062);
and U45856 (N_45856,N_42273,N_43262);
nor U45857 (N_45857,N_43813,N_42955);
nand U45858 (N_45858,N_42171,N_43932);
and U45859 (N_45859,N_42939,N_43404);
or U45860 (N_45860,N_42442,N_42459);
nor U45861 (N_45861,N_43354,N_43685);
nor U45862 (N_45862,N_43586,N_43615);
nor U45863 (N_45863,N_43083,N_42922);
nand U45864 (N_45864,N_43178,N_42667);
nor U45865 (N_45865,N_42325,N_42937);
or U45866 (N_45866,N_42591,N_42828);
nor U45867 (N_45867,N_42342,N_42360);
and U45868 (N_45868,N_43138,N_43671);
and U45869 (N_45869,N_43282,N_42892);
nand U45870 (N_45870,N_43538,N_43388);
xnor U45871 (N_45871,N_43206,N_42674);
and U45872 (N_45872,N_42670,N_42364);
xor U45873 (N_45873,N_43584,N_42210);
and U45874 (N_45874,N_43590,N_43555);
and U45875 (N_45875,N_43330,N_43507);
xnor U45876 (N_45876,N_43569,N_43122);
and U45877 (N_45877,N_42262,N_43672);
nand U45878 (N_45878,N_43791,N_42334);
nand U45879 (N_45879,N_43894,N_43089);
nor U45880 (N_45880,N_43297,N_43264);
xor U45881 (N_45881,N_43767,N_43688);
nor U45882 (N_45882,N_43601,N_43598);
nor U45883 (N_45883,N_43923,N_43880);
xnor U45884 (N_45884,N_43389,N_42772);
nand U45885 (N_45885,N_43623,N_43486);
or U45886 (N_45886,N_43339,N_43984);
nor U45887 (N_45887,N_42799,N_43671);
and U45888 (N_45888,N_43714,N_43246);
nand U45889 (N_45889,N_42582,N_42338);
and U45890 (N_45890,N_43550,N_42321);
nor U45891 (N_45891,N_43434,N_43870);
nor U45892 (N_45892,N_43619,N_43237);
and U45893 (N_45893,N_42533,N_43447);
or U45894 (N_45894,N_43961,N_42345);
nand U45895 (N_45895,N_43519,N_42839);
nand U45896 (N_45896,N_42836,N_42658);
or U45897 (N_45897,N_43693,N_43009);
and U45898 (N_45898,N_42749,N_43706);
and U45899 (N_45899,N_42508,N_42333);
and U45900 (N_45900,N_42033,N_43977);
or U45901 (N_45901,N_43459,N_42528);
xnor U45902 (N_45902,N_43429,N_43893);
xnor U45903 (N_45903,N_43452,N_43151);
nor U45904 (N_45904,N_42793,N_42459);
xor U45905 (N_45905,N_43712,N_43998);
xor U45906 (N_45906,N_42973,N_43573);
xor U45907 (N_45907,N_43974,N_42897);
and U45908 (N_45908,N_42603,N_42807);
nand U45909 (N_45909,N_43205,N_42795);
or U45910 (N_45910,N_42252,N_43835);
xor U45911 (N_45911,N_42893,N_43189);
nand U45912 (N_45912,N_43536,N_42496);
nor U45913 (N_45913,N_42162,N_42523);
and U45914 (N_45914,N_42942,N_42589);
nor U45915 (N_45915,N_42118,N_42229);
and U45916 (N_45916,N_42755,N_42256);
nor U45917 (N_45917,N_43446,N_43540);
and U45918 (N_45918,N_42169,N_43531);
or U45919 (N_45919,N_43528,N_43056);
xnor U45920 (N_45920,N_42424,N_42698);
xnor U45921 (N_45921,N_43459,N_43896);
and U45922 (N_45922,N_42529,N_42614);
nand U45923 (N_45923,N_42561,N_42796);
xor U45924 (N_45924,N_43035,N_43906);
xor U45925 (N_45925,N_42948,N_42325);
nor U45926 (N_45926,N_42373,N_42238);
nand U45927 (N_45927,N_42107,N_42086);
or U45928 (N_45928,N_43418,N_42455);
or U45929 (N_45929,N_42043,N_43995);
nor U45930 (N_45930,N_43068,N_43376);
xnor U45931 (N_45931,N_42504,N_43743);
nand U45932 (N_45932,N_42505,N_43176);
xnor U45933 (N_45933,N_43977,N_42133);
nor U45934 (N_45934,N_43983,N_43632);
nor U45935 (N_45935,N_43752,N_42064);
and U45936 (N_45936,N_42264,N_43914);
and U45937 (N_45937,N_42043,N_43864);
or U45938 (N_45938,N_43769,N_42386);
xor U45939 (N_45939,N_43891,N_42133);
nor U45940 (N_45940,N_42022,N_43358);
nor U45941 (N_45941,N_42268,N_43443);
nor U45942 (N_45942,N_42646,N_43072);
nand U45943 (N_45943,N_42740,N_43985);
nand U45944 (N_45944,N_42051,N_43036);
xnor U45945 (N_45945,N_43261,N_42292);
and U45946 (N_45946,N_42155,N_43887);
nor U45947 (N_45947,N_43336,N_42340);
xor U45948 (N_45948,N_42716,N_42353);
nand U45949 (N_45949,N_43404,N_43949);
and U45950 (N_45950,N_43408,N_43903);
or U45951 (N_45951,N_43284,N_43094);
and U45952 (N_45952,N_43058,N_42496);
nor U45953 (N_45953,N_42674,N_42406);
nand U45954 (N_45954,N_43198,N_43174);
nor U45955 (N_45955,N_43100,N_42913);
and U45956 (N_45956,N_42187,N_43873);
nor U45957 (N_45957,N_42404,N_42975);
nand U45958 (N_45958,N_43332,N_43596);
nand U45959 (N_45959,N_42283,N_42357);
and U45960 (N_45960,N_42835,N_43172);
and U45961 (N_45961,N_42590,N_43910);
xnor U45962 (N_45962,N_43714,N_42273);
and U45963 (N_45963,N_43013,N_42440);
nor U45964 (N_45964,N_42865,N_42509);
nand U45965 (N_45965,N_42462,N_42524);
xnor U45966 (N_45966,N_42032,N_42006);
and U45967 (N_45967,N_43242,N_42433);
and U45968 (N_45968,N_42561,N_42210);
and U45969 (N_45969,N_43664,N_42395);
or U45970 (N_45970,N_42855,N_43754);
and U45971 (N_45971,N_43769,N_43100);
xnor U45972 (N_45972,N_43576,N_42978);
nor U45973 (N_45973,N_43851,N_42857);
nand U45974 (N_45974,N_43904,N_43670);
and U45975 (N_45975,N_42542,N_42642);
or U45976 (N_45976,N_42219,N_42298);
and U45977 (N_45977,N_43737,N_43887);
and U45978 (N_45978,N_43052,N_42000);
nand U45979 (N_45979,N_43231,N_43704);
or U45980 (N_45980,N_43640,N_43108);
nand U45981 (N_45981,N_42022,N_43638);
xnor U45982 (N_45982,N_43443,N_42870);
and U45983 (N_45983,N_43749,N_43958);
nand U45984 (N_45984,N_43328,N_42778);
and U45985 (N_45985,N_43202,N_42993);
or U45986 (N_45986,N_43084,N_43929);
nand U45987 (N_45987,N_43194,N_43411);
and U45988 (N_45988,N_43685,N_42329);
and U45989 (N_45989,N_42540,N_43385);
and U45990 (N_45990,N_42873,N_42691);
and U45991 (N_45991,N_42519,N_42886);
nor U45992 (N_45992,N_42555,N_42988);
nand U45993 (N_45993,N_43935,N_42051);
and U45994 (N_45994,N_42525,N_42037);
and U45995 (N_45995,N_43619,N_43711);
xnor U45996 (N_45996,N_43333,N_43209);
nor U45997 (N_45997,N_42489,N_42243);
nand U45998 (N_45998,N_42649,N_42495);
and U45999 (N_45999,N_42926,N_43286);
xnor U46000 (N_46000,N_45713,N_44671);
nand U46001 (N_46001,N_45469,N_44791);
or U46002 (N_46002,N_45594,N_44117);
and U46003 (N_46003,N_44169,N_44527);
and U46004 (N_46004,N_45473,N_45726);
or U46005 (N_46005,N_44057,N_44596);
xnor U46006 (N_46006,N_45347,N_45183);
or U46007 (N_46007,N_45845,N_45328);
or U46008 (N_46008,N_44160,N_44093);
nand U46009 (N_46009,N_44719,N_44357);
xnor U46010 (N_46010,N_45716,N_44101);
and U46011 (N_46011,N_44733,N_45455);
or U46012 (N_46012,N_44276,N_44022);
nand U46013 (N_46013,N_44996,N_45582);
nor U46014 (N_46014,N_44396,N_44935);
xnor U46015 (N_46015,N_44892,N_44282);
and U46016 (N_46016,N_44312,N_44107);
nor U46017 (N_46017,N_45191,N_45229);
nor U46018 (N_46018,N_45207,N_44395);
nand U46019 (N_46019,N_44466,N_44777);
nand U46020 (N_46020,N_45854,N_45882);
and U46021 (N_46021,N_44685,N_44030);
nand U46022 (N_46022,N_44492,N_44321);
or U46023 (N_46023,N_44518,N_45098);
xnor U46024 (N_46024,N_44289,N_44953);
xnor U46025 (N_46025,N_44054,N_45568);
or U46026 (N_46026,N_44698,N_44069);
xor U46027 (N_46027,N_44666,N_44509);
and U46028 (N_46028,N_44503,N_45069);
nand U46029 (N_46029,N_45619,N_44484);
nor U46030 (N_46030,N_45932,N_44701);
nand U46031 (N_46031,N_44523,N_45419);
nor U46032 (N_46032,N_44916,N_44991);
and U46033 (N_46033,N_45024,N_44674);
or U46034 (N_46034,N_44738,N_44894);
nand U46035 (N_46035,N_45113,N_45530);
and U46036 (N_46036,N_45873,N_44797);
nand U46037 (N_46037,N_45685,N_44658);
nand U46038 (N_46038,N_45858,N_44864);
or U46039 (N_46039,N_44244,N_44035);
nand U46040 (N_46040,N_45536,N_44432);
and U46041 (N_46041,N_44802,N_45775);
nand U46042 (N_46042,N_44016,N_44852);
or U46043 (N_46043,N_45879,N_44636);
and U46044 (N_46044,N_45427,N_44304);
or U46045 (N_46045,N_44973,N_45357);
xor U46046 (N_46046,N_44988,N_44415);
nand U46047 (N_46047,N_44898,N_45373);
nand U46048 (N_46048,N_45399,N_44552);
or U46049 (N_46049,N_44440,N_44232);
and U46050 (N_46050,N_45111,N_45012);
and U46051 (N_46051,N_45596,N_44125);
and U46052 (N_46052,N_44389,N_44655);
or U46053 (N_46053,N_45956,N_44296);
xor U46054 (N_46054,N_45548,N_44362);
or U46055 (N_46055,N_44015,N_44669);
nand U46056 (N_46056,N_45146,N_45015);
or U46057 (N_46057,N_44618,N_44019);
or U46058 (N_46058,N_45417,N_45239);
xnor U46059 (N_46059,N_44416,N_44253);
or U46060 (N_46060,N_45063,N_44786);
xnor U46061 (N_46061,N_44082,N_45360);
or U46062 (N_46062,N_45276,N_44600);
xor U46063 (N_46063,N_45231,N_45168);
nor U46064 (N_46064,N_44757,N_45245);
and U46065 (N_46065,N_44681,N_44340);
nand U46066 (N_46066,N_45566,N_45562);
and U46067 (N_46067,N_44540,N_44794);
and U46068 (N_46068,N_44303,N_45539);
nor U46069 (N_46069,N_44859,N_45254);
or U46070 (N_46070,N_44453,N_44041);
xnor U46071 (N_46071,N_45210,N_44103);
nand U46072 (N_46072,N_44122,N_44162);
or U46073 (N_46073,N_44240,N_45284);
nand U46074 (N_46074,N_45592,N_44447);
and U46075 (N_46075,N_44997,N_45478);
or U46076 (N_46076,N_44670,N_45159);
xnor U46077 (N_46077,N_45553,N_44872);
nand U46078 (N_46078,N_45382,N_45540);
nor U46079 (N_46079,N_44286,N_44207);
nand U46080 (N_46080,N_45929,N_44422);
xnor U46081 (N_46081,N_45390,N_44487);
nor U46082 (N_46082,N_45126,N_45940);
nand U46083 (N_46083,N_45808,N_45060);
nor U46084 (N_46084,N_45326,N_45564);
xor U46085 (N_46085,N_45470,N_44577);
and U46086 (N_46086,N_44405,N_44641);
or U46087 (N_46087,N_44011,N_44407);
or U46088 (N_46088,N_44203,N_45735);
nand U46089 (N_46089,N_45188,N_44426);
xor U46090 (N_46090,N_44564,N_45740);
nand U46091 (N_46091,N_45767,N_44629);
or U46092 (N_46092,N_45179,N_44573);
or U46093 (N_46093,N_45701,N_44936);
xor U46094 (N_46094,N_45192,N_45908);
and U46095 (N_46095,N_44993,N_45538);
and U46096 (N_46096,N_45796,N_44624);
and U46097 (N_46097,N_44141,N_45466);
xnor U46098 (N_46098,N_45717,N_45097);
or U46099 (N_46099,N_45675,N_44753);
xor U46100 (N_46100,N_45105,N_45080);
nor U46101 (N_46101,N_45591,N_44186);
and U46102 (N_46102,N_45616,N_44344);
nor U46103 (N_46103,N_45385,N_44404);
and U46104 (N_46104,N_44586,N_45017);
and U46105 (N_46105,N_44110,N_44451);
nand U46106 (N_46106,N_45081,N_45635);
nor U46107 (N_46107,N_45110,N_44234);
nor U46108 (N_46108,N_44455,N_45046);
and U46109 (N_46109,N_44144,N_44164);
or U46110 (N_46110,N_45176,N_45861);
and U46111 (N_46111,N_44848,N_45516);
and U46112 (N_46112,N_44963,N_45715);
nor U46113 (N_46113,N_44410,N_45802);
xor U46114 (N_46114,N_45617,N_44114);
nor U46115 (N_46115,N_44010,N_45480);
nor U46116 (N_46116,N_45039,N_45282);
and U46117 (N_46117,N_44243,N_44832);
nand U46118 (N_46118,N_44364,N_45345);
nor U46119 (N_46119,N_44984,N_44877);
or U46120 (N_46120,N_45242,N_44033);
or U46121 (N_46121,N_45070,N_45145);
xnor U46122 (N_46122,N_45124,N_45006);
xnor U46123 (N_46123,N_44367,N_44982);
nor U46124 (N_46124,N_45651,N_45263);
and U46125 (N_46125,N_45226,N_45919);
nand U46126 (N_46126,N_44772,N_45278);
xor U46127 (N_46127,N_45147,N_45428);
and U46128 (N_46128,N_45321,N_45313);
xnor U46129 (N_46129,N_44842,N_45163);
and U46130 (N_46130,N_45283,N_44065);
xnor U46131 (N_46131,N_45687,N_45184);
and U46132 (N_46132,N_45318,N_45728);
or U46133 (N_46133,N_44014,N_45247);
nand U46134 (N_46134,N_45950,N_44421);
nor U46135 (N_46135,N_44866,N_44025);
xor U46136 (N_46136,N_45037,N_44970);
or U46137 (N_46137,N_44081,N_44210);
and U46138 (N_46138,N_44941,N_45340);
xnor U46139 (N_46139,N_44768,N_44076);
and U46140 (N_46140,N_45156,N_44088);
xnor U46141 (N_46141,N_45319,N_45777);
nand U46142 (N_46142,N_44420,N_44098);
nand U46143 (N_46143,N_45464,N_45452);
or U46144 (N_46144,N_44132,N_45927);
nand U46145 (N_46145,N_44204,N_45487);
or U46146 (N_46146,N_45605,N_45630);
xnor U46147 (N_46147,N_45165,N_45508);
xor U46148 (N_46148,N_45814,N_45523);
and U46149 (N_46149,N_44750,N_44783);
nor U46150 (N_46150,N_44385,N_44836);
nor U46151 (N_46151,N_45511,N_45601);
xnor U46152 (N_46152,N_44817,N_45604);
nand U46153 (N_46153,N_44940,N_44878);
xnor U46154 (N_46154,N_45439,N_44155);
or U46155 (N_46155,N_45211,N_44247);
xor U46156 (N_46156,N_45640,N_44476);
xnor U46157 (N_46157,N_44902,N_44221);
xor U46158 (N_46158,N_44879,N_45067);
nor U46159 (N_46159,N_44761,N_45141);
nand U46160 (N_46160,N_45085,N_45691);
nor U46161 (N_46161,N_45106,N_45270);
nor U46162 (N_46162,N_44029,N_45661);
or U46163 (N_46163,N_45968,N_45585);
xnor U46164 (N_46164,N_44501,N_44006);
and U46165 (N_46165,N_45410,N_44793);
or U46166 (N_46166,N_45108,N_45557);
or U46167 (N_46167,N_45036,N_45569);
nand U46168 (N_46168,N_44901,N_44598);
nor U46169 (N_46169,N_45057,N_45303);
and U46170 (N_46170,N_44273,N_44885);
or U46171 (N_46171,N_45750,N_44510);
nor U46172 (N_46172,N_45338,N_45797);
nor U46173 (N_46173,N_45670,N_45894);
nor U46174 (N_46174,N_44821,N_44258);
and U46175 (N_46175,N_45380,N_45680);
nand U46176 (N_46176,N_44754,N_45718);
and U46177 (N_46177,N_45415,N_45895);
nand U46178 (N_46178,N_44855,N_45368);
xor U46179 (N_46179,N_44089,N_44507);
nor U46180 (N_46180,N_44539,N_44739);
nor U46181 (N_46181,N_44264,N_44736);
or U46182 (N_46182,N_45101,N_44012);
or U46183 (N_46183,N_45626,N_44708);
xor U46184 (N_46184,N_44283,N_45751);
nor U46185 (N_46185,N_44024,N_44966);
nor U46186 (N_46186,N_45369,N_45838);
or U46187 (N_46187,N_44020,N_45921);
and U46188 (N_46188,N_45412,N_44061);
and U46189 (N_46189,N_44597,N_44956);
and U46190 (N_46190,N_44692,N_45019);
nor U46191 (N_46191,N_44735,N_44327);
and U46192 (N_46192,N_45479,N_45926);
xnor U46193 (N_46193,N_45975,N_45093);
nand U46194 (N_46194,N_44462,N_45910);
nor U46195 (N_46195,N_45265,N_44086);
nand U46196 (N_46196,N_45228,N_45458);
xor U46197 (N_46197,N_45120,N_44555);
nor U46198 (N_46198,N_45565,N_44444);
or U46199 (N_46199,N_45999,N_44652);
and U46200 (N_46200,N_44109,N_44119);
or U46201 (N_46201,N_45864,N_44134);
or U46202 (N_46202,N_44166,N_44860);
or U46203 (N_46203,N_45534,N_45256);
nor U46204 (N_46204,N_44818,N_44686);
and U46205 (N_46205,N_45001,N_45227);
nor U46206 (N_46206,N_45641,N_45799);
nand U46207 (N_46207,N_44128,N_44514);
or U46208 (N_46208,N_44371,N_45957);
nor U46209 (N_46209,N_44197,N_44644);
and U46210 (N_46210,N_44625,N_44500);
xnor U46211 (N_46211,N_45118,N_44260);
nor U46212 (N_46212,N_44580,N_45709);
and U46213 (N_46213,N_44633,N_44252);
or U46214 (N_46214,N_45138,N_45669);
and U46215 (N_46215,N_44788,N_44657);
or U46216 (N_46216,N_45638,N_45496);
xor U46217 (N_46217,N_44691,N_45613);
xnor U46218 (N_46218,N_45599,N_44498);
and U46219 (N_46219,N_45376,N_45885);
xnor U46220 (N_46220,N_44298,N_45995);
xor U46221 (N_46221,N_44206,N_45727);
nand U46222 (N_46222,N_45878,N_44152);
nor U46223 (N_46223,N_44399,N_45408);
and U46224 (N_46224,N_44148,N_44464);
nand U46225 (N_46225,N_44095,N_45367);
nand U46226 (N_46226,N_44102,N_45035);
nand U46227 (N_46227,N_45693,N_44388);
nor U46228 (N_46228,N_45383,N_44201);
xor U46229 (N_46229,N_45436,N_45988);
or U46230 (N_46230,N_44463,N_44962);
and U46231 (N_46231,N_45520,N_45847);
or U46232 (N_46232,N_44502,N_45870);
nor U46233 (N_46233,N_45075,N_44828);
nor U46234 (N_46234,N_45286,N_45459);
nor U46235 (N_46235,N_44397,N_44957);
and U46236 (N_46236,N_45959,N_44331);
nand U46237 (N_46237,N_44827,N_44205);
or U46238 (N_46238,N_45765,N_45759);
nor U46239 (N_46239,N_44229,N_45296);
and U46240 (N_46240,N_44146,N_44071);
and U46241 (N_46241,N_45082,N_45426);
or U46242 (N_46242,N_45089,N_45418);
or U46243 (N_46243,N_45705,N_44716);
nand U46244 (N_46244,N_44048,N_45474);
nor U46245 (N_46245,N_44759,N_44789);
or U46246 (N_46246,N_44700,N_45945);
nand U46247 (N_46247,N_44680,N_44883);
or U46248 (N_46248,N_44194,N_45495);
and U46249 (N_46249,N_45658,N_44895);
nor U46250 (N_46250,N_44917,N_44468);
xor U46251 (N_46251,N_45062,N_45502);
and U46252 (N_46252,N_45632,N_44383);
xnor U46253 (N_46253,N_44001,N_45757);
nor U46254 (N_46254,N_44635,N_45552);
xor U46255 (N_46255,N_44324,N_45501);
and U46256 (N_46256,N_44335,N_45339);
nand U46257 (N_46257,N_44411,N_45515);
nand U46258 (N_46258,N_45800,N_44108);
nor U46259 (N_46259,N_44223,N_45951);
or U46260 (N_46260,N_44561,N_44734);
or U46261 (N_46261,N_44461,N_44649);
xor U46262 (N_46262,N_44773,N_44530);
xor U46263 (N_46263,N_45308,N_44366);
and U46264 (N_46264,N_45529,N_45241);
nand U46265 (N_46265,N_44077,N_44712);
xnor U46266 (N_46266,N_45807,N_45322);
and U46267 (N_46267,N_44419,N_45964);
or U46268 (N_46268,N_44925,N_44373);
nand U46269 (N_46269,N_44978,N_45642);
or U46270 (N_46270,N_44816,N_44241);
nor U46271 (N_46271,N_45337,N_44696);
or U46272 (N_46272,N_44452,N_44630);
and U46273 (N_46273,N_44516,N_44413);
or U46274 (N_46274,N_45262,N_45300);
or U46275 (N_46275,N_45813,N_45551);
or U46276 (N_46276,N_44265,N_44480);
nor U46277 (N_46277,N_44653,N_45009);
nor U46278 (N_46278,N_45510,N_45084);
and U46279 (N_46279,N_44728,N_44104);
nor U46280 (N_46280,N_45679,N_45220);
xnor U46281 (N_46281,N_44427,N_45724);
and U46282 (N_46282,N_45776,N_44121);
xnor U46283 (N_46283,N_44938,N_44812);
nand U46284 (N_46284,N_44271,N_44460);
nor U46285 (N_46285,N_45237,N_45817);
nor U46286 (N_46286,N_45104,N_44292);
xor U46287 (N_46287,N_44270,N_44356);
xor U46288 (N_46288,N_44058,N_45987);
nor U46289 (N_46289,N_45151,N_44178);
xor U46290 (N_46290,N_45633,N_45305);
or U46291 (N_46291,N_44880,N_45665);
nor U46292 (N_46292,N_44952,N_44640);
and U46293 (N_46293,N_44031,N_44918);
or U46294 (N_46294,N_45584,N_45273);
nand U46295 (N_46295,N_44801,N_45819);
nor U46296 (N_46296,N_44912,N_44435);
and U46297 (N_46297,N_44406,N_44100);
nor U46298 (N_46298,N_44319,N_44483);
xnor U46299 (N_46299,N_45781,N_44697);
xnor U46300 (N_46300,N_45792,N_44050);
nor U46301 (N_46301,N_45846,N_45857);
and U46302 (N_46302,N_44308,N_45589);
or U46303 (N_46303,N_45622,N_44780);
nor U46304 (N_46304,N_44343,N_45682);
nand U46305 (N_46305,N_45832,N_45181);
and U46306 (N_46306,N_45881,N_44560);
xnor U46307 (N_46307,N_44809,N_44932);
or U46308 (N_46308,N_45411,N_44847);
nor U46309 (N_46309,N_45875,N_44747);
and U46310 (N_46310,N_44151,N_44578);
and U46311 (N_46311,N_44158,N_44939);
and U46312 (N_46312,N_44980,N_45645);
nand U46313 (N_46313,N_44379,N_45899);
nor U46314 (N_46314,N_44659,N_44147);
or U46315 (N_46315,N_44961,N_45774);
and U46316 (N_46316,N_44209,N_44375);
nand U46317 (N_46317,N_44893,N_45876);
or U46318 (N_46318,N_44450,N_44922);
xnor U46319 (N_46319,N_45747,N_45966);
nand U46320 (N_46320,N_45998,N_44135);
xor U46321 (N_46321,N_44665,N_44694);
nand U46322 (N_46322,N_45737,N_45433);
and U46323 (N_46323,N_45913,N_44843);
or U46324 (N_46324,N_45830,N_44714);
xnor U46325 (N_46325,N_45791,N_45153);
nor U46326 (N_46326,N_45489,N_44611);
and U46327 (N_46327,N_44631,N_44349);
or U46328 (N_46328,N_45550,N_44546);
nor U46329 (N_46329,N_45016,N_44913);
nand U46330 (N_46330,N_45051,N_45066);
and U46331 (N_46331,N_45196,N_45484);
or U46332 (N_46332,N_45289,N_44589);
or U46333 (N_46333,N_45342,N_44575);
or U46334 (N_46334,N_45704,N_44796);
nand U46335 (N_46335,N_44565,N_45805);
xor U46336 (N_46336,N_44705,N_44439);
xor U46337 (N_46337,N_44478,N_44376);
and U46338 (N_46338,N_44212,N_44288);
xor U46339 (N_46339,N_45107,N_45782);
or U46340 (N_46340,N_45855,N_44336);
xnor U46341 (N_46341,N_45423,N_45821);
xor U46342 (N_46342,N_45405,N_44491);
nand U46343 (N_46343,N_44968,N_44261);
or U46344 (N_46344,N_44784,N_44185);
nor U46345 (N_46345,N_45352,N_45744);
nand U46346 (N_46346,N_44599,N_44521);
or U46347 (N_46347,N_44612,N_45071);
nand U46348 (N_46348,N_45361,N_45435);
and U46349 (N_46349,N_45370,N_45272);
nor U46350 (N_46350,N_45355,N_45403);
and U46351 (N_46351,N_44238,N_44703);
and U46352 (N_46352,N_44688,N_45203);
nor U46353 (N_46353,N_45918,N_44920);
xor U46354 (N_46354,N_44187,N_45497);
or U46355 (N_46355,N_45162,N_44008);
and U46356 (N_46356,N_44442,N_44948);
or U46357 (N_46357,N_45912,N_45023);
or U46358 (N_46358,N_44944,N_45264);
nor U46359 (N_46359,N_45201,N_45099);
xor U46360 (N_46360,N_44059,N_45462);
nand U46361 (N_46361,N_45083,N_45903);
xnor U46362 (N_46362,N_44237,N_45150);
or U46363 (N_46363,N_45917,N_44829);
or U46364 (N_46364,N_44930,N_45218);
and U46365 (N_46365,N_45059,N_44255);
and U46366 (N_46366,N_44156,N_45664);
xor U46367 (N_46367,N_45233,N_44554);
or U46368 (N_46368,N_45374,N_45969);
or U46369 (N_46369,N_44026,N_45637);
nor U46370 (N_46370,N_45698,N_44277);
nor U46371 (N_46371,N_45209,N_44525);
nor U46372 (N_46372,N_45652,N_45213);
xnor U46373 (N_46373,N_45135,N_45004);
and U46374 (N_46374,N_45989,N_45749);
nor U46375 (N_46375,N_45974,N_45301);
and U46376 (N_46376,N_45820,N_45180);
or U46377 (N_46377,N_44695,N_45058);
and U46378 (N_46378,N_44831,N_44519);
nor U46379 (N_46379,N_44806,N_44825);
xnor U46380 (N_46380,N_44841,N_45437);
nand U46381 (N_46381,N_45279,N_45030);
or U46382 (N_46382,N_45133,N_44737);
and U46383 (N_46383,N_45772,N_45790);
nand U46384 (N_46384,N_44648,N_44372);
and U46385 (N_46385,N_45505,N_44196);
xor U46386 (N_46386,N_44486,N_45260);
xnor U46387 (N_46387,N_45297,N_45152);
nor U46388 (N_46388,N_45798,N_45033);
nor U46389 (N_46389,N_45973,N_45315);
xnor U46390 (N_46390,N_45666,N_45692);
nor U46391 (N_46391,N_44105,N_44013);
and U46392 (N_46392,N_44544,N_45102);
or U46393 (N_46393,N_45031,N_44333);
nor U46394 (N_46394,N_45499,N_44218);
xor U46395 (N_46395,N_44541,N_45028);
xor U46396 (N_46396,N_45068,N_44769);
xnor U46397 (N_46397,N_44840,N_45331);
xnor U46398 (N_46398,N_45131,N_44605);
nor U46399 (N_46399,N_44091,N_44745);
or U46400 (N_46400,N_45714,N_44181);
xor U46401 (N_46401,N_44834,N_45886);
and U46402 (N_46402,N_45554,N_45555);
nand U46403 (N_46403,N_45689,N_44365);
nor U46404 (N_46404,N_45366,N_45429);
xor U46405 (N_46405,N_45577,N_44726);
and U46406 (N_46406,N_44219,N_45826);
or U46407 (N_46407,N_45663,N_45200);
nand U46408 (N_46408,N_44979,N_44380);
nand U46409 (N_46409,N_45509,N_45323);
or U46410 (N_46410,N_44911,N_45456);
and U46411 (N_46411,N_45268,N_44428);
nand U46412 (N_46412,N_45007,N_45833);
xor U46413 (N_46413,N_44094,N_45696);
or U46414 (N_46414,N_44274,N_45444);
xor U46415 (N_46415,N_44792,N_44358);
and U46416 (N_46416,N_44933,N_45103);
nor U46417 (N_46417,N_44326,N_44672);
and U46418 (N_46418,N_45137,N_45281);
nor U46419 (N_46419,N_45513,N_44165);
xnor U46420 (N_46420,N_44200,N_44746);
nor U46421 (N_46421,N_44943,N_45401);
nor U46422 (N_46422,N_45578,N_44313);
and U46423 (N_46423,N_45848,N_44437);
and U46424 (N_46424,N_45825,N_44459);
nand U46425 (N_46425,N_44711,N_45954);
and U46426 (N_46426,N_45116,N_44715);
xor U46427 (N_46427,N_45924,N_45381);
nor U46428 (N_46428,N_45982,N_45134);
or U46429 (N_46429,N_45525,N_45871);
or U46430 (N_46430,N_44039,N_45365);
or U46431 (N_46431,N_45384,N_45904);
nor U46432 (N_46432,N_44551,N_45087);
nand U46433 (N_46433,N_44369,N_44338);
nand U46434 (N_46434,N_44067,N_44352);
nor U46435 (N_46435,N_45603,N_45117);
nor U46436 (N_46436,N_45330,N_44246);
or U46437 (N_46437,N_45615,N_44713);
nor U46438 (N_46438,N_45450,N_45754);
nand U46439 (N_46439,N_44080,N_45933);
nand U46440 (N_46440,N_44638,N_44301);
nand U46441 (N_46441,N_45026,N_45483);
and U46442 (N_46442,N_45556,N_45748);
or U46443 (N_46443,N_45732,N_44469);
xnor U46444 (N_46444,N_44056,N_45896);
and U46445 (N_46445,N_45606,N_45404);
nor U46446 (N_46446,N_44386,N_45646);
xnor U46447 (N_46447,N_45096,N_44656);
and U46448 (N_46448,N_44136,N_45961);
or U46449 (N_46449,N_44053,N_45041);
and U46450 (N_46450,N_45533,N_45029);
and U46451 (N_46451,N_45863,N_44608);
or U46452 (N_46452,N_45543,N_45362);
nor U46453 (N_46453,N_45518,N_45938);
and U46454 (N_46454,N_44224,N_44348);
nor U46455 (N_46455,N_44927,N_45977);
xnor U46456 (N_46456,N_44975,N_45320);
nand U46457 (N_46457,N_45842,N_45874);
or U46458 (N_46458,N_44009,N_44785);
nor U46459 (N_46459,N_44646,N_45022);
nor U46460 (N_46460,N_44250,N_44875);
xnor U46461 (N_46461,N_44471,N_44300);
and U46462 (N_46462,N_45816,N_44323);
xor U46463 (N_46463,N_45400,N_44284);
nor U46464 (N_46464,N_44438,N_45432);
or U46465 (N_46465,N_45546,N_45743);
and U46466 (N_46466,N_44424,N_45193);
or U46467 (N_46467,N_45052,N_44871);
xor U46468 (N_46468,N_45048,N_44867);
and U46469 (N_46469,N_45407,N_45173);
or U46470 (N_46470,N_45343,N_45441);
or U46471 (N_46471,N_45222,N_45699);
and U46472 (N_46472,N_44003,N_44990);
or U46473 (N_46473,N_44470,N_45843);
and U46474 (N_46474,N_45088,N_45773);
nand U46475 (N_46475,N_45425,N_45761);
nor U46476 (N_46476,N_45558,N_44934);
or U46477 (N_46477,N_45572,N_44562);
or U46478 (N_46478,N_44899,N_45676);
or U46479 (N_46479,N_44766,N_44675);
and U46480 (N_46480,N_45130,N_45413);
xnor U46481 (N_46481,N_45719,N_44779);
and U46482 (N_46482,N_44342,N_44064);
xnor U46483 (N_46483,N_44189,N_45609);
nor U46484 (N_46484,N_44914,N_44002);
nand U46485 (N_46485,N_44449,N_44310);
nor U46486 (N_46486,N_45259,N_45225);
or U46487 (N_46487,N_44645,N_45334);
xnor U46488 (N_46488,N_45522,N_45657);
or U46489 (N_46489,N_45742,N_44846);
and U46490 (N_46490,N_45711,N_44066);
nand U46491 (N_46491,N_44294,N_44131);
nor U46492 (N_46492,N_45818,N_44495);
or U46493 (N_46493,N_44778,N_45027);
and U46494 (N_46494,N_45752,N_44628);
nand U46495 (N_46495,N_45795,N_45449);
or U46496 (N_46496,N_45311,N_44316);
and U46497 (N_46497,N_45293,N_45471);
nand U46498 (N_46498,N_45779,N_45898);
nand U46499 (N_46499,N_45236,N_45936);
nand U46500 (N_46500,N_44374,N_44921);
and U46501 (N_46501,N_45980,N_45299);
nor U46502 (N_46502,N_45739,N_44999);
xnor U46503 (N_46503,N_44838,N_44070);
and U46504 (N_46504,N_45127,N_44722);
nand U46505 (N_46505,N_45831,N_44865);
and U46506 (N_46506,N_45290,N_44613);
nor U46507 (N_46507,N_44524,N_45010);
nand U46508 (N_46508,N_45040,N_44176);
or U46509 (N_46509,N_44572,N_45608);
and U46510 (N_46510,N_44904,N_44063);
xor U46511 (N_46511,N_45055,N_44393);
xor U46512 (N_46512,N_45884,N_44721);
nor U46513 (N_46513,N_44445,N_45667);
nand U46514 (N_46514,N_44254,N_45461);
or U46515 (N_46515,N_45182,N_45703);
nor U46516 (N_46516,N_45335,N_45690);
or U46517 (N_46517,N_45223,N_45128);
nor U46518 (N_46518,N_45000,N_45288);
nand U46519 (N_46519,N_44443,N_44355);
xor U46520 (N_46520,N_45688,N_44161);
xor U46521 (N_46521,N_44729,N_45371);
xor U46522 (N_46522,N_45045,N_45860);
xor U46523 (N_46523,N_45198,N_45937);
nor U46524 (N_46524,N_44903,N_45139);
or U46525 (N_46525,N_45827,N_45043);
nand U46526 (N_46526,N_45490,N_45597);
nor U46527 (N_46527,N_44740,N_45442);
or U46528 (N_46528,N_44537,N_44826);
xor U46529 (N_46529,N_44637,N_45764);
nand U46530 (N_46530,N_45379,N_44891);
nor U46531 (N_46531,N_45285,N_45916);
xor U46532 (N_46532,N_44805,N_45414);
nor U46533 (N_46533,N_44322,N_44868);
and U46534 (N_46534,N_45158,N_45560);
or U46535 (N_46535,N_45324,N_45888);
xnor U46536 (N_46536,N_45901,N_44425);
nand U46537 (N_46537,N_45756,N_44418);
nand U46538 (N_46538,N_45346,N_44731);
nor U46539 (N_46539,N_44488,N_44085);
xor U46540 (N_46540,N_45674,N_45660);
nand U46541 (N_46541,N_45378,N_45386);
xor U46542 (N_46542,N_44857,N_45803);
xnor U46543 (N_46543,N_44370,N_44643);
nor U46544 (N_46544,N_45157,N_44559);
nand U46545 (N_46545,N_44873,N_45018);
or U46546 (N_46546,N_44835,N_45736);
nor U46547 (N_46547,N_44116,N_45160);
nor U46548 (N_46548,N_45454,N_45880);
or U46549 (N_46549,N_45434,N_44267);
and U46550 (N_46550,N_45762,N_45295);
and U46551 (N_46551,N_44143,N_45465);
xor U46552 (N_46552,N_44869,N_45890);
xor U46553 (N_46553,N_44320,N_44617);
and U46554 (N_46554,N_45784,N_45234);
nand U46555 (N_46555,N_44803,N_45477);
xor U46556 (N_46556,N_45806,N_44634);
nor U46557 (N_46557,N_44391,N_45574);
and U46558 (N_46558,N_44142,N_45907);
and U46559 (N_46559,N_45364,N_45388);
and U46560 (N_46560,N_44710,N_44339);
nand U46561 (N_46561,N_45673,N_45769);
nor U46562 (N_46562,N_44018,N_44130);
or U46563 (N_46563,N_45563,N_44190);
nand U46564 (N_46564,N_44632,N_44765);
nor U46565 (N_46565,N_44998,N_44361);
nor U46566 (N_46566,N_44467,N_45889);
nand U46567 (N_46567,N_45984,N_45712);
or U46568 (N_46568,N_45486,N_45148);
and U46569 (N_46569,N_45573,N_45498);
nor U46570 (N_46570,N_45650,N_45061);
and U46571 (N_46571,N_44538,N_44621);
xor U46572 (N_46572,N_44799,N_44907);
or U46573 (N_46573,N_44398,N_45387);
nor U46574 (N_46574,N_44668,N_44236);
nand U46575 (N_46575,N_44822,N_45186);
nand U46576 (N_46576,N_45446,N_45504);
nand U46577 (N_46577,N_44664,N_44179);
nor U46578 (N_46578,N_45042,N_44639);
nand U46579 (N_46579,N_44227,N_44231);
and U46580 (N_46580,N_44511,N_44256);
or U46581 (N_46581,N_45287,N_44167);
nor U46582 (N_46582,N_44170,N_44756);
nand U46583 (N_46583,N_44262,N_44281);
and U46584 (N_46584,N_44707,N_44900);
nor U46585 (N_46585,N_44763,N_44400);
nand U46586 (N_46586,N_44987,N_44302);
xnor U46587 (N_46587,N_44760,N_44568);
or U46588 (N_46588,N_45252,N_44730);
nor U46589 (N_46589,N_45476,N_45869);
xor U46590 (N_46590,N_44034,N_45115);
or U46591 (N_46591,N_45868,N_45482);
and U46592 (N_46592,N_45839,N_44242);
or U46593 (N_46593,N_45431,N_44804);
nor U46594 (N_46594,N_44454,N_45389);
nand U46595 (N_46595,N_45997,N_45034);
or U46596 (N_46596,N_44693,N_44810);
xor U46597 (N_46597,N_44923,N_45235);
nand U46598 (N_46598,N_45094,N_44354);
and U46599 (N_46599,N_44268,N_44127);
nor U46600 (N_46600,N_45187,N_45671);
or U46601 (N_46601,N_45783,N_44607);
nor U46602 (N_46602,N_45922,N_44775);
nor U46603 (N_46603,N_45994,N_45208);
xnor U46604 (N_46604,N_45327,N_45507);
or U46605 (N_46605,N_45702,N_45493);
nand U46606 (N_46606,N_44235,N_44290);
nor U46607 (N_46607,N_44299,N_45468);
xor U46608 (N_46608,N_45955,N_45212);
xnor U46609 (N_46609,N_45358,N_44441);
nor U46610 (N_46610,N_45586,N_44888);
nor U46611 (N_46611,N_44278,N_44285);
or U46612 (N_46612,N_44023,N_45077);
nor U46613 (N_46613,N_44660,N_45341);
xor U46614 (N_46614,N_45393,N_44942);
xor U46615 (N_46615,N_45587,N_44043);
nor U46616 (N_46616,N_44021,N_44099);
nor U46617 (N_46617,N_45588,N_44897);
xor U46618 (N_46618,N_44309,N_45451);
and U46619 (N_46619,N_44175,N_45271);
or U46620 (N_46620,N_45494,N_45100);
or U46621 (N_46621,N_44073,N_45377);
xnor U46622 (N_46622,N_45733,N_45746);
xnor U46623 (N_46623,N_44615,N_45570);
and U46624 (N_46624,N_44330,N_44795);
and U46625 (N_46625,N_44515,N_44584);
or U46626 (N_46626,N_45620,N_44965);
and U46627 (N_46627,N_44755,N_45611);
and U46628 (N_46628,N_44072,N_44862);
nand U46629 (N_46629,N_44594,N_44532);
and U46630 (N_46630,N_45232,N_44725);
and U46631 (N_46631,N_44489,N_45953);
nand U46632 (N_46632,N_45392,N_45050);
nor U46633 (N_46633,N_44188,N_45258);
and U46634 (N_46634,N_45644,N_45144);
or U46635 (N_46635,N_45038,N_45793);
nor U46636 (N_46636,N_44220,N_44702);
or U46637 (N_46637,N_44040,N_44819);
or U46638 (N_46638,N_45810,N_44602);
and U46639 (N_46639,N_44601,N_44228);
and U46640 (N_46640,N_45535,N_45614);
nor U46641 (N_46641,N_45985,N_44662);
xnor U46642 (N_46642,N_45815,N_44679);
and U46643 (N_46643,N_45243,N_44115);
xor U46644 (N_46644,N_44213,N_44198);
or U46645 (N_46645,N_45629,N_44138);
nand U46646 (N_46646,N_45887,N_44172);
and U46647 (N_46647,N_45707,N_45255);
xnor U46648 (N_46648,N_45304,N_45763);
nor U46649 (N_46649,N_44332,N_45925);
nand U46650 (N_46650,N_45911,N_45005);
and U46651 (N_46651,N_45143,N_45544);
xnor U46652 (N_46652,N_45829,N_45409);
or U46653 (N_46653,N_44183,N_45920);
or U46654 (N_46654,N_44727,N_45298);
xnor U46655 (N_46655,N_45627,N_45154);
xor U46656 (N_46656,N_44038,N_44482);
and U46657 (N_46657,N_44090,N_44603);
xor U46658 (N_46658,N_45930,N_45576);
xnor U46659 (N_46659,N_45541,N_44216);
xnor U46660 (N_46660,N_44334,N_45571);
or U46661 (N_46661,N_44954,N_44060);
nor U46662 (N_46662,N_44150,N_44774);
or U46663 (N_46663,N_44049,N_45170);
nand U46664 (N_46664,N_45593,N_44305);
or U46665 (N_46665,N_44971,N_44173);
and U46666 (N_46666,N_44742,N_44297);
or U46667 (N_46667,N_44678,N_45453);
nand U46668 (N_46668,N_45789,N_45109);
or U46669 (N_46669,N_44126,N_45521);
or U46670 (N_46670,N_44360,N_44306);
xor U46671 (N_46671,N_44910,N_44837);
or U46672 (N_46672,N_45149,N_44433);
and U46673 (N_46673,N_44853,N_45194);
xnor U46674 (N_46674,N_45697,N_44931);
and U46675 (N_46675,N_45730,N_45694);
and U46676 (N_46676,N_44699,N_45219);
or U46677 (N_46677,N_44481,N_45760);
and U46678 (N_46678,N_44208,N_44642);
nor U46679 (N_46679,N_45310,N_44472);
or U46680 (N_46680,N_45112,N_44157);
nand U46681 (N_46681,N_44163,N_44046);
xnor U46682 (N_46682,N_44677,N_45850);
and U46683 (N_46683,N_45325,N_44359);
or U46684 (N_46684,N_44967,N_45090);
nor U46685 (N_46685,N_44647,N_45741);
nor U46686 (N_46686,N_44193,N_44531);
and U46687 (N_46687,N_45836,N_44896);
nand U46688 (N_46688,N_44989,N_45923);
xor U46689 (N_46689,N_44663,N_45185);
or U46690 (N_46690,N_44620,N_44522);
and U46691 (N_46691,N_44390,N_45700);
or U46692 (N_46692,N_44287,N_44651);
or U46693 (N_46693,N_45332,N_45729);
and U46694 (N_46694,N_44906,N_45448);
nor U46695 (N_46695,N_44353,N_44499);
nand U46696 (N_46696,N_45915,N_44876);
xnor U46697 (N_46697,N_45877,N_45844);
or U46698 (N_46698,N_45824,N_45656);
nand U46699 (N_46699,N_44550,N_45356);
xor U46700 (N_46700,N_44570,N_44528);
xnor U46701 (N_46701,N_44329,N_44226);
nor U46702 (N_46702,N_44870,N_45607);
nand U46703 (N_46703,N_45786,N_45171);
and U46704 (N_46704,N_45678,N_45722);
or U46705 (N_46705,N_45893,N_44566);
and U46706 (N_46706,N_45948,N_44113);
and U46707 (N_46707,N_44177,N_44517);
nor U46708 (N_46708,N_44798,N_45240);
nor U46709 (N_46709,N_44654,N_45943);
or U46710 (N_46710,N_44800,N_44808);
nor U46711 (N_46711,N_44490,N_45396);
or U46712 (N_46712,N_44964,N_44820);
or U46713 (N_46713,N_45065,N_44485);
xnor U46714 (N_46714,N_45725,N_44547);
nor U46715 (N_46715,N_45856,N_44446);
nor U46716 (N_46716,N_44960,N_45600);
xnor U46717 (N_46717,N_45532,N_45095);
xor U46718 (N_46718,N_45828,N_45914);
nor U46719 (N_46719,N_45900,N_44858);
and U46720 (N_46720,N_44771,N_45967);
and U46721 (N_46721,N_44667,N_45492);
or U46722 (N_46722,N_45475,N_45841);
nor U46723 (N_46723,N_44833,N_44926);
or U46724 (N_46724,N_45197,N_45460);
and U46725 (N_46725,N_45189,N_44762);
nand U46726 (N_46726,N_45064,N_45025);
xnor U46727 (N_46727,N_45561,N_45512);
nand U46728 (N_46728,N_44830,N_44861);
xnor U46729 (N_46729,N_45309,N_44622);
xor U46730 (N_46730,N_44251,N_44744);
and U46731 (N_46731,N_44814,N_45837);
nand U46732 (N_46732,N_45939,N_45244);
or U46733 (N_46733,N_44120,N_45883);
nand U46734 (N_46734,N_45517,N_45996);
nor U46735 (N_46735,N_45269,N_45391);
xnor U46736 (N_46736,N_45053,N_44770);
or U46737 (N_46737,N_45136,N_44087);
xor U46738 (N_46738,N_44473,N_44137);
nor U46739 (N_46739,N_45481,N_44767);
or U46740 (N_46740,N_44610,N_45463);
or U46741 (N_46741,N_45834,N_44387);
or U46742 (N_46742,N_44529,N_45866);
and U46743 (N_46743,N_44363,N_44909);
nand U46744 (N_46744,N_45990,N_45787);
or U46745 (N_46745,N_45092,N_45121);
xor U46746 (N_46746,N_44815,N_44430);
or U46747 (N_46747,N_44096,N_44394);
nor U46748 (N_46748,N_45314,N_45447);
xor U46749 (N_46749,N_45002,N_44248);
nor U46750 (N_46750,N_44849,N_45906);
or U46751 (N_46751,N_44650,N_45734);
nor U46752 (N_46752,N_45545,N_44295);
or U46753 (N_46753,N_44106,N_44751);
and U46754 (N_46754,N_45668,N_44781);
nand U46755 (N_46755,N_45809,N_44946);
nand U46756 (N_46756,N_44269,N_44341);
or U46757 (N_46757,N_44140,N_45549);
and U46758 (N_46758,N_44881,N_44042);
nand U46759 (N_46759,N_45942,N_44811);
xnor U46760 (N_46760,N_45250,N_44856);
nand U46761 (N_46761,N_45811,N_44513);
xnor U46762 (N_46762,N_44854,N_44474);
and U46763 (N_46763,N_45215,N_44000);
or U46764 (N_46764,N_44257,N_44199);
nand U46765 (N_46765,N_45647,N_44409);
or U46766 (N_46766,N_45859,N_44279);
nor U46767 (N_46767,N_44084,N_45172);
nand U46768 (N_46768,N_45851,N_44506);
xnor U46769 (N_46769,N_45983,N_44192);
or U46770 (N_46770,N_44346,N_44548);
or U46771 (N_46771,N_45812,N_44112);
nand U46772 (N_46772,N_45422,N_44585);
or U46773 (N_46773,N_45217,N_44717);
nand U46774 (N_46774,N_44986,N_44919);
nor U46775 (N_46775,N_44623,N_45952);
xor U46776 (N_46776,N_45169,N_45020);
nand U46777 (N_46777,N_45934,N_44661);
or U46778 (N_46778,N_45420,N_44718);
nand U46779 (N_46779,N_45261,N_45780);
nand U46780 (N_46780,N_45178,N_44764);
or U46781 (N_46781,N_45079,N_44275);
or U46782 (N_46782,N_45949,N_45306);
xnor U46783 (N_46783,N_44676,N_45440);
xor U46784 (N_46784,N_44683,N_44475);
or U46785 (N_46785,N_44436,N_44887);
nor U46786 (N_46786,N_44412,N_44494);
nor U46787 (N_46787,N_45350,N_44690);
nor U46788 (N_46788,N_44051,N_45114);
or U46789 (N_46789,N_44741,N_44378);
xor U46790 (N_46790,N_45125,N_44032);
or U46791 (N_46791,N_44230,N_45947);
and U46792 (N_46792,N_44616,N_44083);
nand U46793 (N_46793,N_44673,N_44263);
xnor U46794 (N_46794,N_44037,N_44174);
xnor U46795 (N_46795,N_44890,N_45348);
nand U46796 (N_46796,N_44245,N_45662);
xor U46797 (N_46797,N_44092,N_44315);
nor U46798 (N_46798,N_44458,N_45979);
nand U46799 (N_46799,N_45047,N_45013);
nor U46800 (N_46800,N_44882,N_45547);
nand U46801 (N_46801,N_44317,N_44139);
and U46802 (N_46802,N_44604,N_45397);
and U46803 (N_46803,N_44272,N_45202);
or U46804 (N_46804,N_44824,N_44958);
nand U46805 (N_46805,N_45849,N_45438);
or U46806 (N_46806,N_44807,N_44969);
nand U46807 (N_46807,N_44567,N_45049);
xor U46808 (N_46808,N_45014,N_45528);
nor U46809 (N_46809,N_44595,N_45537);
nor U46810 (N_46810,N_45897,N_44047);
and U46811 (N_46811,N_45054,N_44401);
xnor U46812 (N_46812,N_45872,N_45359);
xnor U46813 (N_46813,N_45643,N_45402);
or U46814 (N_46814,N_44028,N_45623);
nand U46815 (N_46815,N_45579,N_44776);
nand U46816 (N_46816,N_45794,N_44068);
or U46817 (N_46817,N_44184,N_44614);
nor U46818 (N_46818,N_45008,N_45257);
or U46819 (N_46819,N_45902,N_45349);
xor U46820 (N_46820,N_44571,N_45238);
or U46821 (N_46821,N_45853,N_45353);
xnor U46822 (N_46822,N_45970,N_44583);
and U46823 (N_46823,N_44929,N_45155);
nor U46824 (N_46824,N_44558,N_45672);
nor U46825 (N_46825,N_45648,N_44154);
xnor U46826 (N_46826,N_45344,N_44974);
nor U46827 (N_46827,N_45580,N_44111);
xnor U46828 (N_46828,N_44579,N_45214);
xor U46829 (N_46829,N_44291,N_45190);
nor U46830 (N_46830,N_44129,N_44027);
nor U46831 (N_46831,N_45354,N_44017);
xor U46832 (N_46832,N_44574,N_44587);
and U46833 (N_46833,N_44591,N_45801);
nand U46834 (N_46834,N_45074,N_44239);
nand U46835 (N_46835,N_44311,N_45527);
nand U46836 (N_46836,N_44222,N_44512);
and U46837 (N_46837,N_45804,N_45710);
nor U46838 (N_46838,N_45972,N_45329);
nor U46839 (N_46839,N_44844,N_45958);
nand U46840 (N_46840,N_44619,N_44994);
nand U46841 (N_46841,N_45129,N_45336);
xor U46842 (N_46842,N_44945,N_45275);
and U46843 (N_46843,N_45443,N_45177);
nor U46844 (N_46844,N_45519,N_44985);
and U46845 (N_46845,N_44706,N_44977);
xor U46846 (N_46846,N_44749,N_45631);
nand U46847 (N_46847,N_45738,N_44497);
xor U46848 (N_46848,N_44217,N_44609);
or U46849 (N_46849,N_45634,N_45768);
or U46850 (N_46850,N_45683,N_45753);
or U46851 (N_46851,N_44863,N_45221);
nand U46852 (N_46852,N_45655,N_45583);
xor U46853 (N_46853,N_45581,N_45333);
xnor U46854 (N_46854,N_44182,N_44787);
nand U46855 (N_46855,N_45758,N_44949);
nor U46856 (N_46856,N_44496,N_44724);
and U46857 (N_46857,N_45072,N_45978);
nor U46858 (N_46858,N_44005,N_44429);
nand U46859 (N_46859,N_45266,N_45430);
nor U46860 (N_46860,N_44790,N_44408);
and U46861 (N_46861,N_44908,N_45044);
nor U46862 (N_46862,N_45684,N_45398);
nand U46863 (N_46863,N_44392,N_45770);
xnor U46864 (N_46864,N_45624,N_45991);
nor U46865 (N_46865,N_44191,N_44709);
xor U46866 (N_46866,N_44947,N_45840);
and U46867 (N_46867,N_45140,N_45993);
and U46868 (N_46868,N_45174,N_45246);
nand U46869 (N_46869,N_45312,N_45277);
and U46870 (N_46870,N_45292,N_45394);
and U46871 (N_46871,N_45230,N_44758);
and U46872 (N_46872,N_44145,N_45852);
nor U46873 (N_46873,N_45406,N_45823);
and U46874 (N_46874,N_45745,N_44180);
xnor U46875 (N_46875,N_45294,N_44905);
nand U46876 (N_46876,N_44118,N_44504);
nor U46877 (N_46877,N_44590,N_44149);
or U46878 (N_46878,N_44123,N_45625);
nand U46879 (N_46879,N_45056,N_45526);
nand U46880 (N_46880,N_45935,N_45612);
nor U46881 (N_46881,N_45003,N_45788);
or U46882 (N_46882,N_44581,N_44687);
xnor U46883 (N_46883,N_45122,N_44318);
xnor U46884 (N_46884,N_44748,N_44593);
xnor U46885 (N_46885,N_45251,N_44133);
nor U46886 (N_46886,N_44074,N_45161);
nor U46887 (N_46887,N_44720,N_44915);
xnor U46888 (N_46888,N_45659,N_45021);
xnor U46889 (N_46889,N_44924,N_44351);
and U46890 (N_46890,N_45567,N_45941);
and U46891 (N_46891,N_44874,N_45835);
nand U46892 (N_46892,N_44976,N_45416);
and U46893 (N_46893,N_45199,N_45598);
and U46894 (N_46894,N_44384,N_45590);
nor U46895 (N_46895,N_45862,N_45307);
nor U46896 (N_46896,N_45708,N_45175);
nand U46897 (N_46897,N_44328,N_44992);
nor U46898 (N_46898,N_44377,N_44036);
nor U46899 (N_46899,N_44403,N_44233);
xor U46900 (N_46900,N_45867,N_44007);
nor U46901 (N_46901,N_44345,N_44682);
or U46902 (N_46902,N_44983,N_45636);
and U46903 (N_46903,N_45086,N_45032);
or U46904 (N_46904,N_44549,N_44536);
nand U46905 (N_46905,N_44171,N_44563);
xor U46906 (N_46906,N_45695,N_45865);
xor U46907 (N_46907,N_44381,N_45500);
or U46908 (N_46908,N_44159,N_45649);
xnor U46909 (N_46909,N_44782,N_45976);
or U46910 (N_46910,N_44280,N_44479);
nand U46911 (N_46911,N_45639,N_45575);
or U46912 (N_46912,N_45677,N_44314);
and U46913 (N_46913,N_44543,N_45302);
or U46914 (N_46914,N_44704,N_45909);
nor U46915 (N_46915,N_44557,N_45216);
xor U46916 (N_46916,N_45472,N_44457);
nand U46917 (N_46917,N_44723,N_45280);
nand U46918 (N_46918,N_44582,N_44689);
nand U46919 (N_46919,N_44535,N_44423);
and U46920 (N_46920,N_44465,N_45249);
or U46921 (N_46921,N_45167,N_44097);
nand U46922 (N_46922,N_45822,N_44368);
and U46923 (N_46923,N_45731,N_44606);
nand U46924 (N_46924,N_44045,N_45206);
nor U46925 (N_46925,N_45467,N_45960);
nor U46926 (N_46926,N_44337,N_44884);
nor U46927 (N_46927,N_44545,N_45981);
xor U46928 (N_46928,N_45073,N_44075);
or U46929 (N_46929,N_44569,N_45931);
nor U46930 (N_46930,N_44325,N_45992);
nand U46931 (N_46931,N_44556,N_44417);
nand U46932 (N_46932,N_44382,N_45653);
nand U46933 (N_46933,N_44456,N_44950);
xor U46934 (N_46934,N_45457,N_45785);
nand U46935 (N_46935,N_45485,N_45253);
and U46936 (N_46936,N_44955,N_44078);
nor U46937 (N_46937,N_44972,N_45681);
xor U46938 (N_46938,N_45531,N_44684);
or U46939 (N_46939,N_44526,N_45986);
or U46940 (N_46940,N_45621,N_44434);
or U46941 (N_46941,N_44214,N_44508);
or U46942 (N_46942,N_44981,N_44249);
or U46943 (N_46943,N_45618,N_44431);
nor U46944 (N_46944,N_45164,N_45628);
nand U46945 (N_46945,N_44414,N_44813);
nor U46946 (N_46946,N_45351,N_44850);
xnor U46947 (N_46947,N_45946,N_45123);
and U46948 (N_46948,N_44266,N_45766);
nor U46949 (N_46949,N_44004,N_45317);
and U46950 (N_46950,N_45971,N_45132);
nor U46951 (N_46951,N_44493,N_44937);
and U46952 (N_46952,N_45195,N_44477);
nor U46953 (N_46953,N_45491,N_44202);
nand U46954 (N_46954,N_45488,N_45078);
nor U46955 (N_46955,N_45142,N_45424);
xor U46956 (N_46956,N_45119,N_44588);
or U46957 (N_46957,N_45248,N_44576);
or U46958 (N_46958,N_44889,N_45274);
and U46959 (N_46959,N_45204,N_45905);
nor U46960 (N_46960,N_44062,N_45363);
nand U46961 (N_46961,N_44347,N_44627);
xnor U46962 (N_46962,N_45720,N_44350);
nand U46963 (N_46963,N_45375,N_45559);
or U46964 (N_46964,N_44951,N_44886);
or U46965 (N_46965,N_44195,N_44215);
xor U46966 (N_46966,N_45011,N_44520);
nor U46967 (N_46967,N_44448,N_44995);
and U46968 (N_46968,N_44307,N_45723);
xor U46969 (N_46969,N_44553,N_45372);
nand U46970 (N_46970,N_44124,N_44928);
or U46971 (N_46971,N_44542,N_45928);
xor U46972 (N_46972,N_45944,N_44402);
nand U46973 (N_46973,N_44959,N_44845);
or U46974 (N_46974,N_45686,N_45965);
xnor U46975 (N_46975,N_44752,N_45595);
and U46976 (N_46976,N_45891,N_44533);
xnor U46977 (N_46977,N_45721,N_45395);
nor U46978 (N_46978,N_44052,N_45091);
or U46979 (N_46979,N_44259,N_45654);
xor U46980 (N_46980,N_45962,N_45166);
and U46981 (N_46981,N_44293,N_44079);
nand U46982 (N_46982,N_45602,N_45205);
and U46983 (N_46983,N_44055,N_45291);
nand U46984 (N_46984,N_45963,N_44592);
or U46985 (N_46985,N_45755,N_44743);
or U46986 (N_46986,N_45316,N_45445);
nand U46987 (N_46987,N_45503,N_45224);
and U46988 (N_46988,N_44211,N_45778);
xnor U46989 (N_46989,N_45076,N_44168);
xor U46990 (N_46990,N_44505,N_44823);
and U46991 (N_46991,N_44839,N_45267);
xnor U46992 (N_46992,N_45610,N_44626);
nand U46993 (N_46993,N_44732,N_44225);
nand U46994 (N_46994,N_45506,N_45706);
and U46995 (N_46995,N_44534,N_44153);
nor U46996 (N_46996,N_45892,N_45542);
xnor U46997 (N_46997,N_45514,N_44044);
xor U46998 (N_46998,N_45524,N_45421);
nor U46999 (N_46999,N_44851,N_45771);
or U47000 (N_47000,N_45865,N_45190);
nor U47001 (N_47001,N_44933,N_45042);
and U47002 (N_47002,N_45491,N_45574);
or U47003 (N_47003,N_45701,N_44989);
nor U47004 (N_47004,N_45293,N_45967);
xnor U47005 (N_47005,N_44057,N_44108);
nand U47006 (N_47006,N_45008,N_45786);
nand U47007 (N_47007,N_45555,N_44520);
and U47008 (N_47008,N_45185,N_44717);
and U47009 (N_47009,N_45700,N_45666);
or U47010 (N_47010,N_44528,N_45379);
or U47011 (N_47011,N_44190,N_44259);
xor U47012 (N_47012,N_45215,N_45692);
nor U47013 (N_47013,N_45266,N_45230);
xnor U47014 (N_47014,N_44588,N_44663);
or U47015 (N_47015,N_44919,N_44521);
or U47016 (N_47016,N_44678,N_45130);
or U47017 (N_47017,N_45629,N_45330);
or U47018 (N_47018,N_45836,N_44557);
nand U47019 (N_47019,N_44076,N_44349);
and U47020 (N_47020,N_45890,N_45072);
nor U47021 (N_47021,N_44450,N_45989);
nand U47022 (N_47022,N_44826,N_45331);
xor U47023 (N_47023,N_44823,N_44970);
nor U47024 (N_47024,N_44229,N_44492);
xnor U47025 (N_47025,N_44260,N_45459);
nor U47026 (N_47026,N_45289,N_44199);
and U47027 (N_47027,N_44060,N_45758);
and U47028 (N_47028,N_44960,N_45245);
and U47029 (N_47029,N_44345,N_44928);
nand U47030 (N_47030,N_45358,N_45175);
nand U47031 (N_47031,N_44036,N_45947);
xor U47032 (N_47032,N_44411,N_45498);
and U47033 (N_47033,N_45443,N_45812);
or U47034 (N_47034,N_44554,N_44873);
nor U47035 (N_47035,N_45481,N_44824);
xnor U47036 (N_47036,N_45689,N_44651);
and U47037 (N_47037,N_44076,N_44930);
nor U47038 (N_47038,N_44538,N_45013);
nor U47039 (N_47039,N_45869,N_45129);
xnor U47040 (N_47040,N_44638,N_44571);
nor U47041 (N_47041,N_45767,N_44639);
nand U47042 (N_47042,N_44218,N_45721);
nand U47043 (N_47043,N_44769,N_45928);
nor U47044 (N_47044,N_45762,N_44983);
nand U47045 (N_47045,N_44102,N_45675);
nand U47046 (N_47046,N_44971,N_44965);
nand U47047 (N_47047,N_44267,N_45950);
nor U47048 (N_47048,N_44056,N_44615);
nand U47049 (N_47049,N_44999,N_44436);
xnor U47050 (N_47050,N_44874,N_44901);
nand U47051 (N_47051,N_45810,N_45045);
or U47052 (N_47052,N_44050,N_45342);
or U47053 (N_47053,N_44567,N_45656);
nor U47054 (N_47054,N_45609,N_44731);
and U47055 (N_47055,N_45190,N_44252);
xor U47056 (N_47056,N_44685,N_45425);
nand U47057 (N_47057,N_44051,N_44693);
nor U47058 (N_47058,N_45706,N_45875);
and U47059 (N_47059,N_45575,N_45733);
and U47060 (N_47060,N_45174,N_45450);
nand U47061 (N_47061,N_44977,N_44529);
nor U47062 (N_47062,N_44195,N_45381);
or U47063 (N_47063,N_44701,N_44933);
nor U47064 (N_47064,N_44775,N_44274);
nand U47065 (N_47065,N_45256,N_45561);
nor U47066 (N_47066,N_45969,N_45757);
xnor U47067 (N_47067,N_44019,N_45039);
nor U47068 (N_47068,N_44221,N_45136);
or U47069 (N_47069,N_44353,N_44235);
and U47070 (N_47070,N_45157,N_45523);
nor U47071 (N_47071,N_45689,N_45355);
and U47072 (N_47072,N_45177,N_45980);
or U47073 (N_47073,N_44556,N_45228);
nor U47074 (N_47074,N_45699,N_44966);
nand U47075 (N_47075,N_44399,N_44229);
nand U47076 (N_47076,N_45416,N_45610);
nor U47077 (N_47077,N_45111,N_45810);
and U47078 (N_47078,N_44035,N_45006);
xor U47079 (N_47079,N_45701,N_45320);
nand U47080 (N_47080,N_45061,N_44738);
xnor U47081 (N_47081,N_44840,N_45855);
xor U47082 (N_47082,N_44520,N_45742);
and U47083 (N_47083,N_45421,N_45389);
xor U47084 (N_47084,N_45882,N_45562);
nor U47085 (N_47085,N_45330,N_45852);
xnor U47086 (N_47086,N_44801,N_44392);
and U47087 (N_47087,N_44322,N_44416);
nand U47088 (N_47088,N_44478,N_44577);
xor U47089 (N_47089,N_45403,N_45505);
and U47090 (N_47090,N_45053,N_44041);
xor U47091 (N_47091,N_45093,N_44709);
nand U47092 (N_47092,N_44048,N_44481);
xnor U47093 (N_47093,N_44110,N_45100);
and U47094 (N_47094,N_45228,N_44162);
or U47095 (N_47095,N_44298,N_44783);
xnor U47096 (N_47096,N_45358,N_44734);
xnor U47097 (N_47097,N_45120,N_45327);
and U47098 (N_47098,N_44328,N_44868);
nand U47099 (N_47099,N_44795,N_45063);
nor U47100 (N_47100,N_45251,N_44997);
or U47101 (N_47101,N_45118,N_45530);
nand U47102 (N_47102,N_45428,N_45934);
and U47103 (N_47103,N_44067,N_44173);
nor U47104 (N_47104,N_44849,N_45482);
and U47105 (N_47105,N_45349,N_45861);
xor U47106 (N_47106,N_45890,N_45795);
nor U47107 (N_47107,N_44988,N_45483);
nand U47108 (N_47108,N_45655,N_45012);
or U47109 (N_47109,N_44979,N_45479);
and U47110 (N_47110,N_44646,N_44298);
nand U47111 (N_47111,N_44961,N_45380);
or U47112 (N_47112,N_44763,N_45581);
and U47113 (N_47113,N_45199,N_44530);
or U47114 (N_47114,N_44857,N_45023);
and U47115 (N_47115,N_44812,N_44035);
nor U47116 (N_47116,N_44409,N_45427);
nand U47117 (N_47117,N_44236,N_44186);
or U47118 (N_47118,N_44697,N_45299);
xor U47119 (N_47119,N_45821,N_44233);
nor U47120 (N_47120,N_45192,N_45131);
xor U47121 (N_47121,N_44488,N_45587);
xor U47122 (N_47122,N_45940,N_44464);
and U47123 (N_47123,N_44967,N_45280);
nor U47124 (N_47124,N_44600,N_45273);
and U47125 (N_47125,N_44243,N_44241);
nor U47126 (N_47126,N_44713,N_44817);
nor U47127 (N_47127,N_45859,N_45232);
and U47128 (N_47128,N_45628,N_44080);
and U47129 (N_47129,N_45099,N_44050);
or U47130 (N_47130,N_44636,N_44398);
or U47131 (N_47131,N_45880,N_45639);
xnor U47132 (N_47132,N_44128,N_44628);
and U47133 (N_47133,N_45581,N_45313);
or U47134 (N_47134,N_45355,N_44436);
and U47135 (N_47135,N_44195,N_45053);
nor U47136 (N_47136,N_45168,N_44114);
and U47137 (N_47137,N_44816,N_45496);
xor U47138 (N_47138,N_44067,N_45207);
nor U47139 (N_47139,N_44326,N_44730);
or U47140 (N_47140,N_44104,N_45093);
or U47141 (N_47141,N_44014,N_45988);
xor U47142 (N_47142,N_45134,N_44642);
or U47143 (N_47143,N_44266,N_44400);
and U47144 (N_47144,N_45873,N_44763);
and U47145 (N_47145,N_45576,N_44774);
and U47146 (N_47146,N_44236,N_45060);
and U47147 (N_47147,N_45299,N_44422);
nand U47148 (N_47148,N_45383,N_45218);
or U47149 (N_47149,N_44499,N_44306);
xnor U47150 (N_47150,N_44335,N_44475);
nand U47151 (N_47151,N_44248,N_44277);
nor U47152 (N_47152,N_45286,N_44642);
xor U47153 (N_47153,N_44894,N_45486);
nand U47154 (N_47154,N_45097,N_45346);
and U47155 (N_47155,N_45623,N_44130);
or U47156 (N_47156,N_45926,N_44252);
xor U47157 (N_47157,N_44221,N_45203);
nor U47158 (N_47158,N_44130,N_45488);
xor U47159 (N_47159,N_45474,N_45672);
nor U47160 (N_47160,N_45004,N_44143);
and U47161 (N_47161,N_44438,N_44072);
xnor U47162 (N_47162,N_44945,N_44417);
and U47163 (N_47163,N_44635,N_45209);
nor U47164 (N_47164,N_45989,N_45656);
and U47165 (N_47165,N_44723,N_45524);
nand U47166 (N_47166,N_45577,N_44656);
nor U47167 (N_47167,N_44428,N_45189);
or U47168 (N_47168,N_44906,N_45253);
and U47169 (N_47169,N_44505,N_45681);
and U47170 (N_47170,N_45670,N_44927);
nand U47171 (N_47171,N_45186,N_44353);
nor U47172 (N_47172,N_45575,N_45396);
nor U47173 (N_47173,N_45546,N_45432);
and U47174 (N_47174,N_44100,N_44978);
nor U47175 (N_47175,N_45817,N_44020);
xor U47176 (N_47176,N_44982,N_45148);
nor U47177 (N_47177,N_44953,N_45015);
nor U47178 (N_47178,N_45936,N_44700);
and U47179 (N_47179,N_44629,N_44138);
or U47180 (N_47180,N_44978,N_44202);
nor U47181 (N_47181,N_45218,N_45251);
xor U47182 (N_47182,N_45439,N_45375);
and U47183 (N_47183,N_44238,N_45373);
and U47184 (N_47184,N_45680,N_45156);
nand U47185 (N_47185,N_44243,N_44297);
nor U47186 (N_47186,N_44943,N_44068);
xor U47187 (N_47187,N_45669,N_45816);
or U47188 (N_47188,N_45486,N_45878);
or U47189 (N_47189,N_45708,N_44326);
nor U47190 (N_47190,N_45517,N_44942);
nand U47191 (N_47191,N_45929,N_45555);
nand U47192 (N_47192,N_45740,N_44821);
nand U47193 (N_47193,N_44669,N_45380);
nand U47194 (N_47194,N_45305,N_44384);
or U47195 (N_47195,N_44808,N_45675);
or U47196 (N_47196,N_44541,N_45122);
nor U47197 (N_47197,N_45173,N_45350);
or U47198 (N_47198,N_45974,N_44347);
nor U47199 (N_47199,N_45495,N_45235);
nand U47200 (N_47200,N_44643,N_45955);
nand U47201 (N_47201,N_45000,N_44695);
or U47202 (N_47202,N_45264,N_44004);
or U47203 (N_47203,N_44633,N_45594);
nand U47204 (N_47204,N_44539,N_44514);
or U47205 (N_47205,N_44069,N_45882);
and U47206 (N_47206,N_44752,N_45188);
or U47207 (N_47207,N_45461,N_45383);
nor U47208 (N_47208,N_45165,N_44059);
and U47209 (N_47209,N_45035,N_45976);
nor U47210 (N_47210,N_45721,N_44658);
nor U47211 (N_47211,N_44176,N_44652);
nor U47212 (N_47212,N_45013,N_44856);
nand U47213 (N_47213,N_44265,N_45997);
or U47214 (N_47214,N_44188,N_44391);
and U47215 (N_47215,N_44812,N_45606);
and U47216 (N_47216,N_45280,N_45208);
or U47217 (N_47217,N_44962,N_45090);
nand U47218 (N_47218,N_44527,N_44533);
and U47219 (N_47219,N_45389,N_45095);
nand U47220 (N_47220,N_44471,N_44886);
xnor U47221 (N_47221,N_44046,N_45434);
nor U47222 (N_47222,N_44173,N_44793);
and U47223 (N_47223,N_45076,N_45689);
nand U47224 (N_47224,N_45265,N_44265);
and U47225 (N_47225,N_44862,N_45464);
nand U47226 (N_47226,N_45403,N_45003);
or U47227 (N_47227,N_45217,N_44721);
and U47228 (N_47228,N_44957,N_44407);
xor U47229 (N_47229,N_44665,N_44991);
xnor U47230 (N_47230,N_44939,N_45323);
nand U47231 (N_47231,N_44307,N_44603);
xor U47232 (N_47232,N_45914,N_44796);
nand U47233 (N_47233,N_44895,N_45623);
and U47234 (N_47234,N_44421,N_45665);
xnor U47235 (N_47235,N_44671,N_44751);
nand U47236 (N_47236,N_44126,N_44976);
or U47237 (N_47237,N_45751,N_45117);
and U47238 (N_47238,N_45396,N_45837);
nor U47239 (N_47239,N_44092,N_44962);
xor U47240 (N_47240,N_45820,N_45752);
xor U47241 (N_47241,N_45342,N_44993);
nand U47242 (N_47242,N_45300,N_45180);
and U47243 (N_47243,N_45123,N_44823);
and U47244 (N_47244,N_45242,N_44704);
or U47245 (N_47245,N_45726,N_45495);
and U47246 (N_47246,N_44723,N_44212);
xnor U47247 (N_47247,N_45232,N_44037);
and U47248 (N_47248,N_44650,N_45517);
or U47249 (N_47249,N_45564,N_44045);
nand U47250 (N_47250,N_45771,N_45512);
and U47251 (N_47251,N_44755,N_45332);
or U47252 (N_47252,N_44345,N_44470);
xnor U47253 (N_47253,N_44092,N_45437);
or U47254 (N_47254,N_44452,N_45733);
nand U47255 (N_47255,N_45617,N_44815);
and U47256 (N_47256,N_44254,N_44865);
or U47257 (N_47257,N_45068,N_45569);
and U47258 (N_47258,N_44711,N_45572);
or U47259 (N_47259,N_45473,N_44365);
or U47260 (N_47260,N_44670,N_44986);
xnor U47261 (N_47261,N_44051,N_44738);
and U47262 (N_47262,N_44460,N_45165);
nor U47263 (N_47263,N_45786,N_44695);
and U47264 (N_47264,N_45806,N_45348);
nor U47265 (N_47265,N_45280,N_45345);
xor U47266 (N_47266,N_45503,N_44357);
nand U47267 (N_47267,N_44700,N_45089);
nand U47268 (N_47268,N_44354,N_45315);
and U47269 (N_47269,N_45354,N_44130);
or U47270 (N_47270,N_45191,N_44678);
and U47271 (N_47271,N_45240,N_45690);
xor U47272 (N_47272,N_45043,N_44395);
and U47273 (N_47273,N_44334,N_45645);
nor U47274 (N_47274,N_44288,N_44297);
or U47275 (N_47275,N_45395,N_44114);
and U47276 (N_47276,N_44183,N_44854);
nand U47277 (N_47277,N_44714,N_44663);
nor U47278 (N_47278,N_45890,N_45660);
xor U47279 (N_47279,N_44319,N_44019);
nor U47280 (N_47280,N_44447,N_45921);
or U47281 (N_47281,N_45321,N_45096);
xnor U47282 (N_47282,N_45518,N_44255);
nand U47283 (N_47283,N_44323,N_44071);
and U47284 (N_47284,N_44485,N_44319);
and U47285 (N_47285,N_45428,N_45637);
or U47286 (N_47286,N_45106,N_44689);
nor U47287 (N_47287,N_44785,N_45937);
or U47288 (N_47288,N_44055,N_44736);
nor U47289 (N_47289,N_45331,N_45256);
or U47290 (N_47290,N_45592,N_45535);
nor U47291 (N_47291,N_45603,N_45252);
nor U47292 (N_47292,N_44802,N_45789);
or U47293 (N_47293,N_45944,N_44696);
nand U47294 (N_47294,N_44888,N_45455);
nand U47295 (N_47295,N_45258,N_45937);
nor U47296 (N_47296,N_44875,N_44801);
nand U47297 (N_47297,N_44207,N_45824);
nor U47298 (N_47298,N_45715,N_45291);
xnor U47299 (N_47299,N_45814,N_44928);
nor U47300 (N_47300,N_44108,N_45615);
nor U47301 (N_47301,N_45040,N_44526);
and U47302 (N_47302,N_45076,N_44390);
nand U47303 (N_47303,N_44075,N_45589);
and U47304 (N_47304,N_44188,N_44056);
and U47305 (N_47305,N_44601,N_45619);
or U47306 (N_47306,N_45615,N_45203);
nor U47307 (N_47307,N_44654,N_45289);
or U47308 (N_47308,N_44786,N_44705);
nand U47309 (N_47309,N_44860,N_45310);
xor U47310 (N_47310,N_45578,N_45039);
nor U47311 (N_47311,N_45909,N_45097);
nand U47312 (N_47312,N_44230,N_44480);
xor U47313 (N_47313,N_44772,N_44182);
nor U47314 (N_47314,N_45223,N_44751);
and U47315 (N_47315,N_44295,N_45266);
xnor U47316 (N_47316,N_44315,N_45568);
nor U47317 (N_47317,N_45954,N_45077);
or U47318 (N_47318,N_44828,N_45402);
nand U47319 (N_47319,N_44021,N_45765);
or U47320 (N_47320,N_45121,N_44833);
and U47321 (N_47321,N_45224,N_44982);
or U47322 (N_47322,N_45891,N_44430);
nor U47323 (N_47323,N_45066,N_45068);
nor U47324 (N_47324,N_44218,N_44171);
and U47325 (N_47325,N_45544,N_45808);
or U47326 (N_47326,N_44229,N_45681);
or U47327 (N_47327,N_44105,N_45305);
xnor U47328 (N_47328,N_44776,N_45119);
and U47329 (N_47329,N_45881,N_45598);
or U47330 (N_47330,N_44427,N_44370);
xnor U47331 (N_47331,N_44841,N_45454);
and U47332 (N_47332,N_45091,N_45621);
xnor U47333 (N_47333,N_45516,N_45022);
xor U47334 (N_47334,N_45113,N_44947);
nor U47335 (N_47335,N_45571,N_45391);
xor U47336 (N_47336,N_45971,N_44177);
nand U47337 (N_47337,N_44360,N_44117);
nor U47338 (N_47338,N_45796,N_45577);
xnor U47339 (N_47339,N_45056,N_45683);
xnor U47340 (N_47340,N_44164,N_45214);
nor U47341 (N_47341,N_45175,N_44897);
and U47342 (N_47342,N_45415,N_44558);
and U47343 (N_47343,N_44669,N_44886);
xnor U47344 (N_47344,N_45146,N_44543);
nor U47345 (N_47345,N_45037,N_44259);
nand U47346 (N_47346,N_45504,N_44698);
or U47347 (N_47347,N_44838,N_45632);
and U47348 (N_47348,N_45354,N_44110);
and U47349 (N_47349,N_44182,N_44352);
or U47350 (N_47350,N_44277,N_45308);
nand U47351 (N_47351,N_44666,N_45926);
and U47352 (N_47352,N_44304,N_45191);
or U47353 (N_47353,N_45966,N_45828);
nand U47354 (N_47354,N_45924,N_45497);
nand U47355 (N_47355,N_44158,N_45344);
xnor U47356 (N_47356,N_45203,N_44300);
and U47357 (N_47357,N_45296,N_44886);
xnor U47358 (N_47358,N_44792,N_44913);
or U47359 (N_47359,N_45688,N_45469);
or U47360 (N_47360,N_44253,N_44533);
xnor U47361 (N_47361,N_45174,N_45577);
nand U47362 (N_47362,N_44746,N_45978);
xnor U47363 (N_47363,N_45079,N_45462);
nand U47364 (N_47364,N_45072,N_44033);
nor U47365 (N_47365,N_44435,N_44617);
xor U47366 (N_47366,N_44171,N_44898);
or U47367 (N_47367,N_45384,N_44474);
nor U47368 (N_47368,N_44661,N_44397);
nor U47369 (N_47369,N_44902,N_44836);
nor U47370 (N_47370,N_44776,N_44516);
xor U47371 (N_47371,N_45518,N_44130);
and U47372 (N_47372,N_44346,N_45214);
nor U47373 (N_47373,N_45259,N_44284);
and U47374 (N_47374,N_44879,N_45250);
xor U47375 (N_47375,N_45358,N_44364);
nand U47376 (N_47376,N_45389,N_45073);
or U47377 (N_47377,N_44232,N_44332);
or U47378 (N_47378,N_45132,N_44251);
nand U47379 (N_47379,N_44046,N_44275);
nand U47380 (N_47380,N_45392,N_45352);
and U47381 (N_47381,N_45535,N_45776);
nand U47382 (N_47382,N_45514,N_45158);
and U47383 (N_47383,N_44019,N_45453);
or U47384 (N_47384,N_45733,N_44241);
xor U47385 (N_47385,N_45970,N_44161);
or U47386 (N_47386,N_44237,N_45892);
nor U47387 (N_47387,N_45920,N_44488);
or U47388 (N_47388,N_45836,N_45825);
nand U47389 (N_47389,N_44411,N_45315);
xnor U47390 (N_47390,N_44375,N_45915);
or U47391 (N_47391,N_45739,N_44920);
or U47392 (N_47392,N_45203,N_44587);
xnor U47393 (N_47393,N_45857,N_44427);
xor U47394 (N_47394,N_44059,N_44570);
nor U47395 (N_47395,N_45135,N_44032);
nand U47396 (N_47396,N_44979,N_45026);
or U47397 (N_47397,N_44046,N_45267);
nand U47398 (N_47398,N_45422,N_45207);
xor U47399 (N_47399,N_44021,N_44735);
nor U47400 (N_47400,N_44998,N_45837);
and U47401 (N_47401,N_44087,N_45756);
nand U47402 (N_47402,N_45589,N_45216);
nand U47403 (N_47403,N_44141,N_44965);
or U47404 (N_47404,N_44364,N_44585);
nand U47405 (N_47405,N_45603,N_44130);
or U47406 (N_47406,N_45522,N_45700);
or U47407 (N_47407,N_44296,N_44559);
nor U47408 (N_47408,N_45127,N_45900);
nor U47409 (N_47409,N_44513,N_45877);
or U47410 (N_47410,N_45735,N_45730);
xor U47411 (N_47411,N_44433,N_45193);
nor U47412 (N_47412,N_44054,N_44351);
xor U47413 (N_47413,N_45189,N_44036);
xor U47414 (N_47414,N_45529,N_44864);
xnor U47415 (N_47415,N_44660,N_45435);
nand U47416 (N_47416,N_45205,N_44758);
xor U47417 (N_47417,N_45147,N_45605);
xnor U47418 (N_47418,N_44118,N_45024);
xnor U47419 (N_47419,N_45438,N_45527);
nand U47420 (N_47420,N_44769,N_45779);
xor U47421 (N_47421,N_45884,N_44493);
or U47422 (N_47422,N_44048,N_44726);
xor U47423 (N_47423,N_45234,N_44744);
and U47424 (N_47424,N_44547,N_44266);
nor U47425 (N_47425,N_44563,N_45080);
xnor U47426 (N_47426,N_44473,N_44718);
or U47427 (N_47427,N_45971,N_44241);
or U47428 (N_47428,N_45987,N_45570);
xor U47429 (N_47429,N_45232,N_45956);
nand U47430 (N_47430,N_44650,N_44805);
nand U47431 (N_47431,N_44595,N_45090);
nor U47432 (N_47432,N_45282,N_44962);
xnor U47433 (N_47433,N_45802,N_45711);
and U47434 (N_47434,N_44675,N_45662);
xor U47435 (N_47435,N_45726,N_44566);
xor U47436 (N_47436,N_45103,N_44612);
and U47437 (N_47437,N_44493,N_44731);
nand U47438 (N_47438,N_45771,N_45212);
nor U47439 (N_47439,N_44700,N_44418);
xnor U47440 (N_47440,N_44788,N_44139);
nor U47441 (N_47441,N_44838,N_44252);
nor U47442 (N_47442,N_44031,N_44511);
xnor U47443 (N_47443,N_45793,N_45298);
or U47444 (N_47444,N_45380,N_44284);
xnor U47445 (N_47445,N_44000,N_45008);
xor U47446 (N_47446,N_45888,N_45282);
nand U47447 (N_47447,N_45552,N_44226);
nand U47448 (N_47448,N_44581,N_45398);
xnor U47449 (N_47449,N_45022,N_44082);
nor U47450 (N_47450,N_44130,N_45977);
and U47451 (N_47451,N_45755,N_44070);
and U47452 (N_47452,N_44584,N_45720);
or U47453 (N_47453,N_45116,N_45538);
nor U47454 (N_47454,N_45542,N_45614);
and U47455 (N_47455,N_45654,N_44231);
xor U47456 (N_47456,N_44641,N_45989);
nand U47457 (N_47457,N_45398,N_44303);
nand U47458 (N_47458,N_44343,N_44615);
nor U47459 (N_47459,N_45709,N_45513);
nor U47460 (N_47460,N_45331,N_44842);
nand U47461 (N_47461,N_44563,N_44867);
xnor U47462 (N_47462,N_45493,N_44255);
or U47463 (N_47463,N_45367,N_44567);
nor U47464 (N_47464,N_44494,N_44113);
and U47465 (N_47465,N_44894,N_45066);
nor U47466 (N_47466,N_44085,N_45829);
xor U47467 (N_47467,N_45129,N_45956);
nand U47468 (N_47468,N_44497,N_45872);
and U47469 (N_47469,N_45666,N_45995);
or U47470 (N_47470,N_45954,N_44304);
nand U47471 (N_47471,N_45562,N_44561);
xnor U47472 (N_47472,N_45405,N_44267);
or U47473 (N_47473,N_44411,N_45707);
nand U47474 (N_47474,N_45146,N_44717);
nor U47475 (N_47475,N_45318,N_45243);
or U47476 (N_47476,N_45196,N_44541);
nand U47477 (N_47477,N_45732,N_44355);
nor U47478 (N_47478,N_44100,N_45087);
xor U47479 (N_47479,N_44421,N_45201);
xnor U47480 (N_47480,N_44434,N_44189);
xnor U47481 (N_47481,N_44055,N_45206);
nand U47482 (N_47482,N_44289,N_45350);
and U47483 (N_47483,N_44769,N_45686);
and U47484 (N_47484,N_45752,N_45216);
nand U47485 (N_47485,N_44881,N_44677);
and U47486 (N_47486,N_45317,N_44397);
nor U47487 (N_47487,N_45903,N_45846);
nor U47488 (N_47488,N_45017,N_45996);
and U47489 (N_47489,N_45570,N_45729);
nor U47490 (N_47490,N_45190,N_45691);
xnor U47491 (N_47491,N_45949,N_45487);
nand U47492 (N_47492,N_45702,N_44725);
nor U47493 (N_47493,N_45125,N_45247);
and U47494 (N_47494,N_45962,N_44287);
xor U47495 (N_47495,N_44932,N_44706);
and U47496 (N_47496,N_45588,N_44108);
and U47497 (N_47497,N_45714,N_45630);
nor U47498 (N_47498,N_45391,N_45925);
or U47499 (N_47499,N_45065,N_44695);
nand U47500 (N_47500,N_44570,N_44827);
nand U47501 (N_47501,N_45106,N_45285);
or U47502 (N_47502,N_44802,N_45728);
xnor U47503 (N_47503,N_44014,N_44725);
or U47504 (N_47504,N_44377,N_44513);
xnor U47505 (N_47505,N_45308,N_45416);
nor U47506 (N_47506,N_44062,N_44557);
or U47507 (N_47507,N_45159,N_45741);
or U47508 (N_47508,N_45116,N_44296);
nor U47509 (N_47509,N_45429,N_44456);
xor U47510 (N_47510,N_45672,N_45635);
or U47511 (N_47511,N_45662,N_45343);
nand U47512 (N_47512,N_45381,N_44969);
and U47513 (N_47513,N_44974,N_45050);
nand U47514 (N_47514,N_44338,N_45575);
or U47515 (N_47515,N_45531,N_45433);
nand U47516 (N_47516,N_44801,N_45234);
and U47517 (N_47517,N_44735,N_44073);
nor U47518 (N_47518,N_45917,N_44729);
and U47519 (N_47519,N_45417,N_44993);
xor U47520 (N_47520,N_45797,N_45308);
xnor U47521 (N_47521,N_44725,N_44885);
xnor U47522 (N_47522,N_45004,N_44959);
nor U47523 (N_47523,N_45754,N_45630);
xnor U47524 (N_47524,N_45291,N_44559);
and U47525 (N_47525,N_44182,N_44217);
and U47526 (N_47526,N_44478,N_44304);
or U47527 (N_47527,N_45945,N_45342);
and U47528 (N_47528,N_44679,N_44436);
nand U47529 (N_47529,N_45340,N_44922);
xor U47530 (N_47530,N_45121,N_44125);
nor U47531 (N_47531,N_44215,N_45364);
xor U47532 (N_47532,N_44978,N_44372);
nor U47533 (N_47533,N_45910,N_45188);
or U47534 (N_47534,N_45065,N_45110);
xnor U47535 (N_47535,N_44503,N_45827);
and U47536 (N_47536,N_44049,N_45573);
nor U47537 (N_47537,N_45987,N_45133);
or U47538 (N_47538,N_44884,N_44000);
nor U47539 (N_47539,N_44219,N_45055);
nand U47540 (N_47540,N_45051,N_44708);
and U47541 (N_47541,N_45249,N_44458);
and U47542 (N_47542,N_44987,N_44781);
nor U47543 (N_47543,N_44828,N_44939);
nand U47544 (N_47544,N_45169,N_45351);
nor U47545 (N_47545,N_44577,N_45634);
and U47546 (N_47546,N_44322,N_44203);
nand U47547 (N_47547,N_44245,N_45165);
and U47548 (N_47548,N_44965,N_45985);
nor U47549 (N_47549,N_45908,N_44158);
xnor U47550 (N_47550,N_45193,N_45653);
and U47551 (N_47551,N_44708,N_44754);
nor U47552 (N_47552,N_45878,N_45092);
nand U47553 (N_47553,N_45655,N_44242);
or U47554 (N_47554,N_44734,N_45821);
xor U47555 (N_47555,N_45000,N_44515);
and U47556 (N_47556,N_45248,N_44114);
and U47557 (N_47557,N_44737,N_45257);
nand U47558 (N_47558,N_45839,N_45964);
xnor U47559 (N_47559,N_45533,N_44524);
xnor U47560 (N_47560,N_45763,N_44025);
nand U47561 (N_47561,N_45391,N_45139);
or U47562 (N_47562,N_45520,N_45634);
and U47563 (N_47563,N_44431,N_44433);
nor U47564 (N_47564,N_44894,N_44938);
nor U47565 (N_47565,N_45315,N_45505);
nor U47566 (N_47566,N_44256,N_45950);
or U47567 (N_47567,N_44012,N_45470);
nor U47568 (N_47568,N_44999,N_44433);
nand U47569 (N_47569,N_45650,N_45427);
xnor U47570 (N_47570,N_44531,N_45998);
and U47571 (N_47571,N_45962,N_45546);
nor U47572 (N_47572,N_44491,N_44503);
nand U47573 (N_47573,N_44974,N_45888);
nor U47574 (N_47574,N_44202,N_45741);
nor U47575 (N_47575,N_44629,N_44942);
nor U47576 (N_47576,N_45598,N_45786);
nor U47577 (N_47577,N_45168,N_44275);
xor U47578 (N_47578,N_45993,N_45083);
nand U47579 (N_47579,N_45784,N_45347);
nor U47580 (N_47580,N_44768,N_44760);
xor U47581 (N_47581,N_45327,N_44555);
nor U47582 (N_47582,N_44788,N_45624);
xnor U47583 (N_47583,N_45210,N_45793);
and U47584 (N_47584,N_44099,N_45944);
or U47585 (N_47585,N_44025,N_45128);
nor U47586 (N_47586,N_45557,N_45329);
xor U47587 (N_47587,N_45459,N_44390);
or U47588 (N_47588,N_44209,N_45964);
nand U47589 (N_47589,N_45599,N_45722);
and U47590 (N_47590,N_45630,N_44267);
or U47591 (N_47591,N_45170,N_45844);
and U47592 (N_47592,N_45898,N_45009);
xor U47593 (N_47593,N_45766,N_45911);
xor U47594 (N_47594,N_44677,N_44940);
or U47595 (N_47595,N_44714,N_44160);
xor U47596 (N_47596,N_45697,N_44769);
xnor U47597 (N_47597,N_45119,N_45299);
nor U47598 (N_47598,N_45062,N_44774);
or U47599 (N_47599,N_45875,N_45118);
nand U47600 (N_47600,N_45590,N_44638);
or U47601 (N_47601,N_45257,N_44720);
xor U47602 (N_47602,N_45697,N_44526);
nor U47603 (N_47603,N_44799,N_45113);
xnor U47604 (N_47604,N_45748,N_45854);
xor U47605 (N_47605,N_44487,N_45672);
or U47606 (N_47606,N_44538,N_44274);
or U47607 (N_47607,N_45952,N_44986);
xnor U47608 (N_47608,N_44400,N_44819);
nand U47609 (N_47609,N_45338,N_44646);
or U47610 (N_47610,N_44904,N_44069);
nand U47611 (N_47611,N_44104,N_45814);
xor U47612 (N_47612,N_44329,N_44164);
and U47613 (N_47613,N_44996,N_44971);
and U47614 (N_47614,N_45146,N_44032);
nor U47615 (N_47615,N_44271,N_45500);
and U47616 (N_47616,N_44156,N_44941);
and U47617 (N_47617,N_45793,N_45829);
xnor U47618 (N_47618,N_45465,N_45178);
or U47619 (N_47619,N_44783,N_44926);
nand U47620 (N_47620,N_45772,N_45571);
nor U47621 (N_47621,N_44017,N_45615);
nand U47622 (N_47622,N_44807,N_45081);
and U47623 (N_47623,N_45800,N_45150);
nand U47624 (N_47624,N_45014,N_44552);
and U47625 (N_47625,N_45634,N_45540);
nand U47626 (N_47626,N_44667,N_44278);
nor U47627 (N_47627,N_44918,N_44496);
nand U47628 (N_47628,N_44777,N_45730);
and U47629 (N_47629,N_44905,N_44908);
and U47630 (N_47630,N_45011,N_44890);
and U47631 (N_47631,N_45784,N_45573);
and U47632 (N_47632,N_45812,N_45772);
nor U47633 (N_47633,N_45231,N_44205);
xor U47634 (N_47634,N_45628,N_44256);
xnor U47635 (N_47635,N_44203,N_45060);
nor U47636 (N_47636,N_44868,N_45135);
or U47637 (N_47637,N_44903,N_45710);
nand U47638 (N_47638,N_44544,N_45878);
nor U47639 (N_47639,N_45669,N_45880);
xnor U47640 (N_47640,N_44570,N_44065);
and U47641 (N_47641,N_44468,N_45713);
nand U47642 (N_47642,N_45915,N_44020);
nor U47643 (N_47643,N_45839,N_45065);
xnor U47644 (N_47644,N_45205,N_45938);
nor U47645 (N_47645,N_44017,N_44117);
nor U47646 (N_47646,N_45181,N_44422);
nor U47647 (N_47647,N_44318,N_45760);
nor U47648 (N_47648,N_45123,N_44091);
or U47649 (N_47649,N_45467,N_44312);
nand U47650 (N_47650,N_44379,N_44252);
nand U47651 (N_47651,N_45957,N_45302);
nand U47652 (N_47652,N_45613,N_45304);
nor U47653 (N_47653,N_45809,N_45401);
nor U47654 (N_47654,N_44897,N_44371);
xor U47655 (N_47655,N_44293,N_44763);
or U47656 (N_47656,N_44392,N_45124);
nor U47657 (N_47657,N_45179,N_45191);
xor U47658 (N_47658,N_45412,N_45258);
xnor U47659 (N_47659,N_45622,N_45007);
or U47660 (N_47660,N_45806,N_44371);
xnor U47661 (N_47661,N_44246,N_45981);
and U47662 (N_47662,N_44089,N_45949);
or U47663 (N_47663,N_45711,N_44581);
or U47664 (N_47664,N_44857,N_45817);
nand U47665 (N_47665,N_44831,N_44587);
xnor U47666 (N_47666,N_45262,N_45800);
or U47667 (N_47667,N_44399,N_45129);
xnor U47668 (N_47668,N_45035,N_44828);
or U47669 (N_47669,N_44995,N_44482);
xnor U47670 (N_47670,N_44827,N_45750);
or U47671 (N_47671,N_44794,N_45137);
nor U47672 (N_47672,N_44589,N_45667);
or U47673 (N_47673,N_44951,N_45326);
nor U47674 (N_47674,N_45347,N_44271);
and U47675 (N_47675,N_44497,N_45294);
nor U47676 (N_47676,N_44360,N_44831);
and U47677 (N_47677,N_44055,N_44767);
nor U47678 (N_47678,N_45673,N_45853);
xnor U47679 (N_47679,N_45555,N_44460);
nand U47680 (N_47680,N_45484,N_44548);
or U47681 (N_47681,N_45305,N_44438);
nand U47682 (N_47682,N_45606,N_45051);
xnor U47683 (N_47683,N_45299,N_45878);
and U47684 (N_47684,N_44936,N_44578);
nand U47685 (N_47685,N_44612,N_44089);
xor U47686 (N_47686,N_45543,N_44812);
or U47687 (N_47687,N_45267,N_45186);
nand U47688 (N_47688,N_45817,N_44496);
and U47689 (N_47689,N_44126,N_45239);
or U47690 (N_47690,N_44488,N_45518);
and U47691 (N_47691,N_45173,N_44640);
nand U47692 (N_47692,N_44223,N_45712);
or U47693 (N_47693,N_44842,N_45663);
xnor U47694 (N_47694,N_44251,N_45749);
xnor U47695 (N_47695,N_44090,N_45446);
nand U47696 (N_47696,N_44751,N_45962);
nand U47697 (N_47697,N_45115,N_44385);
nor U47698 (N_47698,N_44746,N_44394);
and U47699 (N_47699,N_44686,N_44284);
nor U47700 (N_47700,N_45408,N_45635);
nand U47701 (N_47701,N_45391,N_44217);
nor U47702 (N_47702,N_45600,N_44457);
and U47703 (N_47703,N_45053,N_44400);
xor U47704 (N_47704,N_44831,N_44270);
or U47705 (N_47705,N_45413,N_44882);
nor U47706 (N_47706,N_45233,N_44181);
and U47707 (N_47707,N_45545,N_45625);
nor U47708 (N_47708,N_45399,N_44948);
nor U47709 (N_47709,N_44304,N_45568);
and U47710 (N_47710,N_44684,N_44504);
nand U47711 (N_47711,N_45220,N_45676);
or U47712 (N_47712,N_45848,N_45783);
nand U47713 (N_47713,N_44073,N_44890);
and U47714 (N_47714,N_45002,N_45907);
nand U47715 (N_47715,N_45579,N_44652);
nand U47716 (N_47716,N_44634,N_45543);
or U47717 (N_47717,N_44211,N_44832);
xnor U47718 (N_47718,N_45405,N_45307);
nor U47719 (N_47719,N_45168,N_45259);
nor U47720 (N_47720,N_45423,N_44420);
and U47721 (N_47721,N_44461,N_44524);
xor U47722 (N_47722,N_45196,N_44157);
xnor U47723 (N_47723,N_44339,N_45423);
xnor U47724 (N_47724,N_45024,N_44380);
nand U47725 (N_47725,N_44158,N_45735);
or U47726 (N_47726,N_45442,N_45454);
xnor U47727 (N_47727,N_44253,N_45161);
xor U47728 (N_47728,N_45449,N_45708);
and U47729 (N_47729,N_45731,N_44878);
nor U47730 (N_47730,N_44138,N_44552);
xnor U47731 (N_47731,N_45534,N_45159);
and U47732 (N_47732,N_45656,N_45431);
and U47733 (N_47733,N_45123,N_45471);
xnor U47734 (N_47734,N_45646,N_45884);
xnor U47735 (N_47735,N_45587,N_45012);
nand U47736 (N_47736,N_44299,N_45385);
xor U47737 (N_47737,N_44064,N_44589);
xor U47738 (N_47738,N_45429,N_44954);
nand U47739 (N_47739,N_45755,N_44889);
or U47740 (N_47740,N_45412,N_44944);
and U47741 (N_47741,N_44211,N_45240);
or U47742 (N_47742,N_44163,N_44102);
nor U47743 (N_47743,N_45257,N_44226);
and U47744 (N_47744,N_44165,N_45502);
nor U47745 (N_47745,N_44396,N_44087);
nor U47746 (N_47746,N_45455,N_44552);
or U47747 (N_47747,N_45069,N_45785);
and U47748 (N_47748,N_45277,N_45150);
xor U47749 (N_47749,N_44866,N_44583);
nor U47750 (N_47750,N_44203,N_44838);
nor U47751 (N_47751,N_45107,N_44856);
xnor U47752 (N_47752,N_44954,N_44797);
and U47753 (N_47753,N_44422,N_44705);
nand U47754 (N_47754,N_44287,N_45099);
or U47755 (N_47755,N_44040,N_45927);
nand U47756 (N_47756,N_45141,N_45165);
nor U47757 (N_47757,N_44989,N_45752);
or U47758 (N_47758,N_44802,N_44329);
or U47759 (N_47759,N_45671,N_44536);
nand U47760 (N_47760,N_44211,N_45222);
nand U47761 (N_47761,N_44914,N_45795);
xor U47762 (N_47762,N_45672,N_45330);
and U47763 (N_47763,N_45418,N_44650);
and U47764 (N_47764,N_45717,N_44804);
or U47765 (N_47765,N_45632,N_45574);
and U47766 (N_47766,N_45492,N_44899);
nand U47767 (N_47767,N_45301,N_44060);
or U47768 (N_47768,N_45663,N_44807);
nor U47769 (N_47769,N_45261,N_45445);
or U47770 (N_47770,N_44431,N_45980);
xor U47771 (N_47771,N_44090,N_45876);
nand U47772 (N_47772,N_45351,N_44405);
nand U47773 (N_47773,N_45363,N_44299);
or U47774 (N_47774,N_45796,N_44336);
and U47775 (N_47775,N_45898,N_44897);
or U47776 (N_47776,N_44505,N_44720);
and U47777 (N_47777,N_44625,N_45635);
xor U47778 (N_47778,N_44522,N_45497);
or U47779 (N_47779,N_45670,N_45463);
and U47780 (N_47780,N_45182,N_44348);
or U47781 (N_47781,N_44036,N_44557);
xnor U47782 (N_47782,N_45150,N_44243);
xor U47783 (N_47783,N_44836,N_45345);
nand U47784 (N_47784,N_45439,N_44902);
and U47785 (N_47785,N_44791,N_44676);
or U47786 (N_47786,N_44100,N_45573);
and U47787 (N_47787,N_44879,N_45437);
nor U47788 (N_47788,N_45522,N_45606);
or U47789 (N_47789,N_44570,N_44413);
nor U47790 (N_47790,N_45704,N_45194);
or U47791 (N_47791,N_45593,N_44568);
nand U47792 (N_47792,N_44303,N_44441);
nor U47793 (N_47793,N_44924,N_45935);
nand U47794 (N_47794,N_45907,N_44535);
xor U47795 (N_47795,N_45649,N_45142);
xnor U47796 (N_47796,N_45390,N_44469);
or U47797 (N_47797,N_45528,N_45096);
nor U47798 (N_47798,N_45189,N_44504);
or U47799 (N_47799,N_45869,N_45751);
nand U47800 (N_47800,N_44839,N_45229);
xnor U47801 (N_47801,N_45565,N_44045);
and U47802 (N_47802,N_45201,N_45518);
nand U47803 (N_47803,N_45377,N_45994);
and U47804 (N_47804,N_44321,N_45136);
nor U47805 (N_47805,N_44736,N_44493);
nor U47806 (N_47806,N_44850,N_44129);
and U47807 (N_47807,N_45257,N_45287);
and U47808 (N_47808,N_45443,N_45957);
and U47809 (N_47809,N_45034,N_44999);
or U47810 (N_47810,N_44512,N_44406);
nand U47811 (N_47811,N_45104,N_45853);
xor U47812 (N_47812,N_44971,N_44617);
xor U47813 (N_47813,N_45973,N_45542);
xnor U47814 (N_47814,N_45006,N_44845);
xor U47815 (N_47815,N_45781,N_45244);
nor U47816 (N_47816,N_45677,N_44164);
or U47817 (N_47817,N_45031,N_44663);
nand U47818 (N_47818,N_44959,N_44592);
or U47819 (N_47819,N_45543,N_45925);
xnor U47820 (N_47820,N_44587,N_45902);
xnor U47821 (N_47821,N_44040,N_44141);
nor U47822 (N_47822,N_44978,N_45671);
and U47823 (N_47823,N_44332,N_45620);
and U47824 (N_47824,N_45607,N_45964);
nor U47825 (N_47825,N_45053,N_44928);
and U47826 (N_47826,N_45595,N_44152);
or U47827 (N_47827,N_44025,N_45666);
xnor U47828 (N_47828,N_45857,N_44608);
nand U47829 (N_47829,N_45834,N_44296);
xor U47830 (N_47830,N_44486,N_44938);
nand U47831 (N_47831,N_44927,N_45567);
nor U47832 (N_47832,N_44631,N_44328);
nor U47833 (N_47833,N_44807,N_44916);
nand U47834 (N_47834,N_45522,N_45326);
nand U47835 (N_47835,N_44377,N_45020);
nand U47836 (N_47836,N_44677,N_44859);
xor U47837 (N_47837,N_45970,N_45041);
nor U47838 (N_47838,N_45670,N_44397);
or U47839 (N_47839,N_44796,N_45248);
or U47840 (N_47840,N_44357,N_45730);
xor U47841 (N_47841,N_44071,N_45667);
nand U47842 (N_47842,N_45215,N_44995);
nor U47843 (N_47843,N_45210,N_44705);
nor U47844 (N_47844,N_44502,N_44111);
xnor U47845 (N_47845,N_44861,N_45986);
nand U47846 (N_47846,N_45481,N_44951);
and U47847 (N_47847,N_45303,N_45128);
and U47848 (N_47848,N_45293,N_45137);
or U47849 (N_47849,N_44347,N_44583);
and U47850 (N_47850,N_44841,N_44423);
xor U47851 (N_47851,N_45603,N_44806);
xor U47852 (N_47852,N_44938,N_45120);
xnor U47853 (N_47853,N_45547,N_45613);
and U47854 (N_47854,N_44996,N_44869);
nor U47855 (N_47855,N_44456,N_45821);
xnor U47856 (N_47856,N_45383,N_45343);
nor U47857 (N_47857,N_44130,N_45632);
and U47858 (N_47858,N_44832,N_44651);
xnor U47859 (N_47859,N_45465,N_44693);
nand U47860 (N_47860,N_45702,N_45562);
xnor U47861 (N_47861,N_44357,N_45837);
nor U47862 (N_47862,N_45124,N_45871);
xnor U47863 (N_47863,N_44461,N_45607);
and U47864 (N_47864,N_44921,N_45508);
and U47865 (N_47865,N_45078,N_45231);
or U47866 (N_47866,N_44089,N_44633);
nand U47867 (N_47867,N_45160,N_44902);
nor U47868 (N_47868,N_44237,N_44117);
and U47869 (N_47869,N_44486,N_45091);
xor U47870 (N_47870,N_44464,N_44233);
nor U47871 (N_47871,N_45615,N_45322);
or U47872 (N_47872,N_44759,N_44416);
nor U47873 (N_47873,N_44236,N_45267);
and U47874 (N_47874,N_44368,N_44959);
nand U47875 (N_47875,N_44091,N_44522);
or U47876 (N_47876,N_45048,N_44703);
and U47877 (N_47877,N_45251,N_44365);
xor U47878 (N_47878,N_45209,N_44723);
or U47879 (N_47879,N_44412,N_45695);
and U47880 (N_47880,N_44976,N_45389);
nand U47881 (N_47881,N_44665,N_44532);
and U47882 (N_47882,N_45215,N_45578);
xnor U47883 (N_47883,N_45057,N_45281);
nor U47884 (N_47884,N_45777,N_45730);
xor U47885 (N_47885,N_45778,N_44114);
xor U47886 (N_47886,N_45707,N_44636);
or U47887 (N_47887,N_45739,N_44124);
and U47888 (N_47888,N_44878,N_44101);
or U47889 (N_47889,N_45557,N_44131);
nand U47890 (N_47890,N_45221,N_45550);
nand U47891 (N_47891,N_44206,N_45205);
and U47892 (N_47892,N_45648,N_45221);
xnor U47893 (N_47893,N_45992,N_45726);
or U47894 (N_47894,N_44397,N_44189);
and U47895 (N_47895,N_45540,N_45716);
nand U47896 (N_47896,N_44963,N_44722);
nand U47897 (N_47897,N_45367,N_44903);
nand U47898 (N_47898,N_44605,N_45965);
nand U47899 (N_47899,N_45634,N_45037);
or U47900 (N_47900,N_45124,N_45819);
or U47901 (N_47901,N_44121,N_44697);
or U47902 (N_47902,N_45572,N_45313);
xnor U47903 (N_47903,N_45041,N_45693);
or U47904 (N_47904,N_45769,N_45319);
nand U47905 (N_47905,N_44661,N_44720);
and U47906 (N_47906,N_45844,N_45880);
and U47907 (N_47907,N_45260,N_45822);
nand U47908 (N_47908,N_45164,N_45751);
xnor U47909 (N_47909,N_45272,N_44197);
or U47910 (N_47910,N_45290,N_44427);
and U47911 (N_47911,N_44668,N_44697);
xnor U47912 (N_47912,N_44876,N_45437);
or U47913 (N_47913,N_44744,N_44128);
or U47914 (N_47914,N_45246,N_44364);
nor U47915 (N_47915,N_44178,N_44125);
xnor U47916 (N_47916,N_44649,N_45843);
or U47917 (N_47917,N_45710,N_45664);
or U47918 (N_47918,N_44938,N_44870);
nand U47919 (N_47919,N_45785,N_44073);
and U47920 (N_47920,N_45167,N_44901);
or U47921 (N_47921,N_44357,N_44659);
and U47922 (N_47922,N_45397,N_45544);
nand U47923 (N_47923,N_44915,N_44212);
xor U47924 (N_47924,N_45085,N_45180);
or U47925 (N_47925,N_45226,N_44192);
and U47926 (N_47926,N_44020,N_44688);
or U47927 (N_47927,N_44995,N_45784);
or U47928 (N_47928,N_44016,N_45923);
nor U47929 (N_47929,N_45189,N_44722);
nand U47930 (N_47930,N_44160,N_45749);
and U47931 (N_47931,N_44296,N_44246);
and U47932 (N_47932,N_45991,N_45294);
nand U47933 (N_47933,N_45471,N_45758);
xnor U47934 (N_47934,N_44578,N_45445);
xor U47935 (N_47935,N_45570,N_45141);
xor U47936 (N_47936,N_44904,N_45151);
and U47937 (N_47937,N_45366,N_44690);
nand U47938 (N_47938,N_44366,N_45446);
xnor U47939 (N_47939,N_45271,N_44093);
and U47940 (N_47940,N_45294,N_44682);
nor U47941 (N_47941,N_44563,N_45199);
or U47942 (N_47942,N_45142,N_44373);
or U47943 (N_47943,N_45302,N_44468);
xor U47944 (N_47944,N_44125,N_44048);
xor U47945 (N_47945,N_44309,N_45827);
and U47946 (N_47946,N_44626,N_45764);
xnor U47947 (N_47947,N_45809,N_44581);
nand U47948 (N_47948,N_45572,N_45061);
nand U47949 (N_47949,N_44847,N_44948);
and U47950 (N_47950,N_45826,N_44877);
and U47951 (N_47951,N_44095,N_44508);
nor U47952 (N_47952,N_44283,N_45710);
nand U47953 (N_47953,N_44191,N_44233);
nor U47954 (N_47954,N_44404,N_44045);
and U47955 (N_47955,N_45697,N_44562);
nor U47956 (N_47956,N_45770,N_45646);
nand U47957 (N_47957,N_44597,N_45488);
xor U47958 (N_47958,N_45101,N_45734);
and U47959 (N_47959,N_45027,N_44607);
or U47960 (N_47960,N_44419,N_44017);
nor U47961 (N_47961,N_44619,N_45294);
or U47962 (N_47962,N_45422,N_44510);
nor U47963 (N_47963,N_45208,N_45834);
or U47964 (N_47964,N_45039,N_44446);
xnor U47965 (N_47965,N_45269,N_45135);
nand U47966 (N_47966,N_44471,N_44111);
xor U47967 (N_47967,N_44874,N_44041);
xor U47968 (N_47968,N_45987,N_45490);
or U47969 (N_47969,N_45075,N_44353);
xor U47970 (N_47970,N_44113,N_45954);
and U47971 (N_47971,N_45796,N_45656);
xor U47972 (N_47972,N_45113,N_44335);
xor U47973 (N_47973,N_45604,N_44587);
or U47974 (N_47974,N_45980,N_45903);
xor U47975 (N_47975,N_44988,N_45270);
nand U47976 (N_47976,N_45898,N_44339);
nor U47977 (N_47977,N_45269,N_45600);
nor U47978 (N_47978,N_45084,N_45809);
nor U47979 (N_47979,N_45003,N_44181);
xnor U47980 (N_47980,N_44079,N_44304);
nand U47981 (N_47981,N_44955,N_45751);
xnor U47982 (N_47982,N_45836,N_45754);
nand U47983 (N_47983,N_45549,N_45735);
xor U47984 (N_47984,N_44768,N_45302);
nand U47985 (N_47985,N_44990,N_44332);
and U47986 (N_47986,N_45580,N_45755);
or U47987 (N_47987,N_45904,N_44075);
or U47988 (N_47988,N_45302,N_45627);
xor U47989 (N_47989,N_44645,N_45136);
nor U47990 (N_47990,N_45035,N_45928);
nand U47991 (N_47991,N_44837,N_45469);
or U47992 (N_47992,N_44545,N_45610);
nand U47993 (N_47993,N_45521,N_45700);
nand U47994 (N_47994,N_44655,N_44342);
and U47995 (N_47995,N_45256,N_45864);
or U47996 (N_47996,N_44698,N_44648);
or U47997 (N_47997,N_45500,N_44610);
nor U47998 (N_47998,N_44716,N_44419);
and U47999 (N_47999,N_44547,N_45643);
and U48000 (N_48000,N_47647,N_46816);
and U48001 (N_48001,N_47435,N_46843);
and U48002 (N_48002,N_47086,N_46564);
or U48003 (N_48003,N_47166,N_47518);
nor U48004 (N_48004,N_47207,N_47648);
nor U48005 (N_48005,N_47653,N_47246);
xnor U48006 (N_48006,N_47122,N_47358);
or U48007 (N_48007,N_47916,N_47157);
nor U48008 (N_48008,N_46881,N_47556);
xnor U48009 (N_48009,N_46479,N_46361);
xnor U48010 (N_48010,N_46658,N_47586);
xor U48011 (N_48011,N_47508,N_46462);
xor U48012 (N_48012,N_47046,N_47546);
xnor U48013 (N_48013,N_47231,N_47761);
nand U48014 (N_48014,N_46427,N_46923);
xor U48015 (N_48015,N_46886,N_47901);
or U48016 (N_48016,N_47198,N_47027);
and U48017 (N_48017,N_46268,N_46793);
xor U48018 (N_48018,N_46161,N_46039);
nand U48019 (N_48019,N_46720,N_46723);
and U48020 (N_48020,N_47377,N_46027);
and U48021 (N_48021,N_46790,N_47188);
and U48022 (N_48022,N_47737,N_47178);
or U48023 (N_48023,N_46120,N_46249);
nand U48024 (N_48024,N_46074,N_46111);
or U48025 (N_48025,N_46679,N_46169);
xor U48026 (N_48026,N_47095,N_46890);
and U48027 (N_48027,N_46256,N_47357);
xor U48028 (N_48028,N_46451,N_46885);
and U48029 (N_48029,N_46563,N_46367);
xor U48030 (N_48030,N_47999,N_47504);
nor U48031 (N_48031,N_46476,N_46138);
or U48032 (N_48032,N_46731,N_46434);
and U48033 (N_48033,N_46058,N_47200);
or U48034 (N_48034,N_47941,N_46013);
xor U48035 (N_48035,N_46714,N_47028);
nor U48036 (N_48036,N_47078,N_46783);
nor U48037 (N_48037,N_46412,N_47312);
and U48038 (N_48038,N_46985,N_46053);
and U48039 (N_48039,N_46078,N_46849);
nand U48040 (N_48040,N_47215,N_46568);
or U48041 (N_48041,N_46704,N_47505);
or U48042 (N_48042,N_46775,N_47488);
or U48043 (N_48043,N_47510,N_46520);
xor U48044 (N_48044,N_47446,N_46421);
nand U48045 (N_48045,N_46023,N_47611);
and U48046 (N_48046,N_46273,N_46917);
and U48047 (N_48047,N_46153,N_46506);
nor U48048 (N_48048,N_46175,N_46746);
and U48049 (N_48049,N_46713,N_47303);
nand U48050 (N_48050,N_47764,N_47381);
xnor U48051 (N_48051,N_46113,N_46542);
or U48052 (N_48052,N_46470,N_46229);
and U48053 (N_48053,N_47535,N_47110);
nor U48054 (N_48054,N_47282,N_46072);
or U48055 (N_48055,N_46370,N_47224);
nand U48056 (N_48056,N_46641,N_47242);
nand U48057 (N_48057,N_46937,N_46348);
and U48058 (N_48058,N_47197,N_47346);
nor U48059 (N_48059,N_46295,N_47663);
xor U48060 (N_48060,N_46057,N_47905);
or U48061 (N_48061,N_47530,N_47990);
xor U48062 (N_48062,N_46684,N_47772);
xnor U48063 (N_48063,N_46910,N_47688);
nor U48064 (N_48064,N_46149,N_47199);
and U48065 (N_48065,N_46029,N_47855);
xor U48066 (N_48066,N_47263,N_47895);
xor U48067 (N_48067,N_46776,N_47393);
and U48068 (N_48068,N_47472,N_46709);
xor U48069 (N_48069,N_46270,N_46635);
xnor U48070 (N_48070,N_47115,N_47871);
nor U48071 (N_48071,N_47707,N_46395);
or U48072 (N_48072,N_47991,N_46871);
or U48073 (N_48073,N_47969,N_46547);
nand U48074 (N_48074,N_46499,N_47770);
nand U48075 (N_48075,N_46305,N_47475);
xor U48076 (N_48076,N_46645,N_46947);
nand U48077 (N_48077,N_47238,N_46449);
xnor U48078 (N_48078,N_46255,N_47755);
nor U48079 (N_48079,N_46445,N_47018);
nor U48080 (N_48080,N_47699,N_47387);
or U48081 (N_48081,N_46541,N_46101);
nor U48082 (N_48082,N_47585,N_46204);
nor U48083 (N_48083,N_46328,N_46241);
nor U48084 (N_48084,N_46181,N_47296);
nor U48085 (N_48085,N_47172,N_46016);
nor U48086 (N_48086,N_47844,N_47070);
and U48087 (N_48087,N_47436,N_46948);
and U48088 (N_48088,N_46152,N_47645);
xnor U48089 (N_48089,N_47654,N_46815);
nor U48090 (N_48090,N_46488,N_46810);
nor U48091 (N_48091,N_47763,N_46595);
and U48092 (N_48092,N_46675,N_46480);
nor U48093 (N_48093,N_46493,N_47208);
and U48094 (N_48094,N_47592,N_46835);
nand U48095 (N_48095,N_46888,N_46509);
or U48096 (N_48096,N_47203,N_46222);
xnor U48097 (N_48097,N_47998,N_46104);
xor U48098 (N_48098,N_46077,N_47927);
nand U48099 (N_48099,N_46555,N_47361);
xor U48100 (N_48100,N_47971,N_47824);
nand U48101 (N_48101,N_47049,N_47039);
nand U48102 (N_48102,N_46093,N_47938);
nor U48103 (N_48103,N_46892,N_47751);
and U48104 (N_48104,N_46308,N_46096);
and U48105 (N_48105,N_47536,N_46654);
xor U48106 (N_48106,N_47730,N_47142);
nor U48107 (N_48107,N_46371,N_46114);
xor U48108 (N_48108,N_46409,N_46124);
or U48109 (N_48109,N_46549,N_47118);
and U48110 (N_48110,N_46267,N_47960);
or U48111 (N_48111,N_47913,N_47462);
nor U48112 (N_48112,N_47532,N_46396);
and U48113 (N_48113,N_46218,N_47635);
xnor U48114 (N_48114,N_47909,N_46807);
and U48115 (N_48115,N_47691,N_46192);
and U48116 (N_48116,N_47622,N_46208);
or U48117 (N_48117,N_47547,N_46014);
nor U48118 (N_48118,N_46426,N_46082);
xnor U48119 (N_48119,N_46213,N_47450);
nand U48120 (N_48120,N_46264,N_47310);
or U48121 (N_48121,N_47766,N_46227);
nand U48122 (N_48122,N_46177,N_47900);
nor U48123 (N_48123,N_47814,N_46770);
xnor U48124 (N_48124,N_47422,N_47050);
nor U48125 (N_48125,N_46316,N_47798);
xnor U48126 (N_48126,N_47390,N_47064);
xnor U48127 (N_48127,N_47352,N_46147);
or U48128 (N_48128,N_47785,N_47232);
nor U48129 (N_48129,N_47152,N_47126);
nor U48130 (N_48130,N_47201,N_46442);
xnor U48131 (N_48131,N_47407,N_46293);
nor U48132 (N_48132,N_46364,N_46719);
nand U48133 (N_48133,N_47348,N_47665);
xnor U48134 (N_48134,N_46696,N_46453);
nand U48135 (N_48135,N_47099,N_47526);
nor U48136 (N_48136,N_46360,N_46188);
or U48137 (N_48137,N_47401,N_47162);
nor U48138 (N_48138,N_47204,N_47805);
nor U48139 (N_48139,N_46613,N_46374);
nor U48140 (N_48140,N_46199,N_47290);
and U48141 (N_48141,N_47155,N_47255);
and U48142 (N_48142,N_46333,N_46610);
or U48143 (N_48143,N_47241,N_47173);
nor U48144 (N_48144,N_46601,N_47291);
xnor U48145 (N_48145,N_46182,N_46724);
and U48146 (N_48146,N_46909,N_47644);
nand U48147 (N_48147,N_46266,N_46365);
and U48148 (N_48148,N_47513,N_46605);
nor U48149 (N_48149,N_47331,N_46779);
nand U48150 (N_48150,N_47044,N_46748);
nor U48151 (N_48151,N_46945,N_47421);
or U48152 (N_48152,N_47794,N_46135);
and U48153 (N_48153,N_47870,N_47749);
and U48154 (N_48154,N_47013,N_47080);
and U48155 (N_48155,N_46042,N_46350);
xor U48156 (N_48156,N_47425,N_47946);
nor U48157 (N_48157,N_47087,N_46545);
and U48158 (N_48158,N_46800,N_47048);
nor U48159 (N_48159,N_47917,N_47906);
and U48160 (N_48160,N_46855,N_46358);
nand U48161 (N_48161,N_46336,N_47692);
xor U48162 (N_48162,N_47693,N_47497);
xnor U48163 (N_48163,N_46686,N_46926);
nand U48164 (N_48164,N_47477,N_47284);
nor U48165 (N_48165,N_47278,N_46059);
xnor U48166 (N_48166,N_47822,N_47955);
xnor U48167 (N_48167,N_47926,N_47759);
xnor U48168 (N_48168,N_46484,N_46047);
or U48169 (N_48169,N_46632,N_47340);
and U48170 (N_48170,N_46536,N_46763);
or U48171 (N_48171,N_47214,N_47796);
and U48172 (N_48172,N_47218,N_47182);
and U48173 (N_48173,N_47486,N_46738);
xnor U48174 (N_48174,N_46162,N_46463);
xor U48175 (N_48175,N_46244,N_47298);
and U48176 (N_48176,N_47561,N_47107);
or U48177 (N_48177,N_46651,N_46503);
nand U48178 (N_48178,N_46676,N_46340);
and U48179 (N_48179,N_47174,N_46502);
nand U48180 (N_48180,N_46750,N_47384);
and U48181 (N_48181,N_47285,N_46960);
or U48182 (N_48182,N_47803,N_47704);
and U48183 (N_48183,N_46403,N_47982);
and U48184 (N_48184,N_46845,N_46257);
nand U48185 (N_48185,N_46962,N_46544);
xor U48186 (N_48186,N_47079,N_47935);
nand U48187 (N_48187,N_47826,N_47575);
or U48188 (N_48188,N_47459,N_47410);
or U48189 (N_48189,N_47958,N_46311);
and U48190 (N_48190,N_47088,N_47524);
and U48191 (N_48191,N_46500,N_46225);
nand U48192 (N_48192,N_47499,N_47506);
xnor U48193 (N_48193,N_46160,N_47374);
nor U48194 (N_48194,N_46982,N_46010);
and U48195 (N_48195,N_47184,N_47360);
nand U48196 (N_48196,N_47633,N_47300);
and U48197 (N_48197,N_47891,N_47581);
nor U48198 (N_48198,N_46475,N_46315);
or U48199 (N_48199,N_47779,N_47394);
or U48200 (N_48200,N_46924,N_46325);
nand U48201 (N_48201,N_47863,N_46851);
and U48202 (N_48202,N_47453,N_46323);
and U48203 (N_48203,N_46247,N_47769);
and U48204 (N_48204,N_46408,N_46991);
xnor U48205 (N_48205,N_47601,N_47458);
and U48206 (N_48206,N_47503,N_46322);
and U48207 (N_48207,N_46183,N_47864);
nor U48208 (N_48208,N_46980,N_46394);
xor U48209 (N_48209,N_47321,N_47213);
nor U48210 (N_48210,N_47727,N_46879);
and U48211 (N_48211,N_47799,N_46377);
and U48212 (N_48212,N_46938,N_46884);
xor U48213 (N_48213,N_47343,N_47771);
nand U48214 (N_48214,N_47565,N_47065);
or U48215 (N_48215,N_47922,N_47783);
and U48216 (N_48216,N_46435,N_47041);
nand U48217 (N_48217,N_46265,N_47976);
or U48218 (N_48218,N_47075,N_46146);
and U48219 (N_48219,N_47484,N_46665);
or U48220 (N_48220,N_47131,N_47217);
nand U48221 (N_48221,N_47067,N_47409);
xnor U48222 (N_48222,N_46401,N_47090);
nand U48223 (N_48223,N_47137,N_46652);
or U48224 (N_48224,N_47161,N_47528);
or U48225 (N_48225,N_46179,N_47679);
xor U48226 (N_48226,N_47205,N_46575);
nor U48227 (N_48227,N_47550,N_46703);
and U48228 (N_48228,N_47167,N_46024);
or U48229 (N_48229,N_46596,N_46424);
nor U48230 (N_48230,N_47868,N_47420);
nand U48231 (N_48231,N_47010,N_46521);
nor U48232 (N_48232,N_47083,N_47689);
xor U48233 (N_48233,N_46519,N_46319);
nor U48234 (N_48234,N_47587,N_47825);
and U48235 (N_48235,N_47037,N_46341);
and U48236 (N_48236,N_47514,N_47397);
nor U48237 (N_48237,N_47379,N_47886);
and U48238 (N_48238,N_46172,N_46460);
xnor U48239 (N_48239,N_46697,N_47657);
nor U48240 (N_48240,N_46667,N_47280);
or U48241 (N_48241,N_46130,N_46232);
xor U48242 (N_48242,N_47024,N_46356);
xnor U48243 (N_48243,N_47627,N_46951);
or U48244 (N_48244,N_46105,N_46128);
nor U48245 (N_48245,N_47327,N_46646);
or U48246 (N_48246,N_47744,N_46876);
and U48247 (N_48247,N_46139,N_47681);
nand U48248 (N_48248,N_47521,N_47624);
nor U48249 (N_48249,N_47001,N_47711);
and U48250 (N_48250,N_47192,N_47671);
and U48251 (N_48251,N_47997,N_46718);
xnor U48252 (N_48252,N_47568,N_47372);
or U48253 (N_48253,N_46492,N_47845);
or U48254 (N_48254,N_46231,N_47442);
nor U48255 (N_48255,N_47406,N_46640);
nand U48256 (N_48256,N_46936,N_47884);
nor U48257 (N_48257,N_47936,N_46301);
and U48258 (N_48258,N_46122,N_47288);
nor U48259 (N_48259,N_47852,N_47376);
and U48260 (N_48260,N_47438,N_46622);
nand U48261 (N_48261,N_46051,N_47915);
nand U48262 (N_48262,N_46875,N_46739);
nor U48263 (N_48263,N_47823,N_47713);
xnor U48264 (N_48264,N_46907,N_46446);
nand U48265 (N_48265,N_47543,N_46604);
nor U48266 (N_48266,N_46136,N_46725);
and U48267 (N_48267,N_46398,N_46098);
nand U48268 (N_48268,N_47652,N_46469);
nor U48269 (N_48269,N_46045,N_46338);
and U48270 (N_48270,N_47403,N_46226);
nor U48271 (N_48271,N_47341,N_47818);
nand U48272 (N_48272,N_47967,N_46242);
nand U48273 (N_48273,N_47978,N_46209);
or U48274 (N_48274,N_46819,N_47029);
and U48275 (N_48275,N_46872,N_46869);
nor U48276 (N_48276,N_47591,N_46811);
xor U48277 (N_48277,N_46299,N_46882);
nor U48278 (N_48278,N_47778,N_47345);
xor U48279 (N_48279,N_46617,N_47252);
nand U48280 (N_48280,N_47792,N_47183);
and U48281 (N_48281,N_46863,N_46669);
xnor U48282 (N_48282,N_47856,N_47190);
xnor U48283 (N_48283,N_47795,N_46729);
and U48284 (N_48284,N_46964,N_46769);
nand U48285 (N_48285,N_46523,N_47800);
nand U48286 (N_48286,N_47669,N_47009);
xor U48287 (N_48287,N_47271,N_46473);
and U48288 (N_48288,N_47317,N_46543);
xor U48289 (N_48289,N_47593,N_47714);
or U48290 (N_48290,N_47431,N_47716);
or U48291 (N_48291,N_46334,N_47239);
nand U48292 (N_48292,N_47081,N_46223);
and U48293 (N_48293,N_46952,N_46789);
nand U48294 (N_48294,N_47718,N_46376);
nand U48295 (N_48295,N_47570,N_46198);
nand U48296 (N_48296,N_47059,N_47701);
or U48297 (N_48297,N_47983,N_47875);
nand U48298 (N_48298,N_47114,N_47194);
nor U48299 (N_48299,N_47094,N_47816);
nand U48300 (N_48300,N_46954,N_47482);
or U48301 (N_48301,N_47417,N_46711);
and U48302 (N_48302,N_47382,N_46785);
nand U48303 (N_48303,N_47077,N_47202);
xor U48304 (N_48304,N_47702,N_46466);
or U48305 (N_48305,N_47685,N_46387);
nand U48306 (N_48306,N_46764,N_47861);
nand U48307 (N_48307,N_47225,N_47897);
nor U48308 (N_48308,N_47996,N_46963);
or U48309 (N_48309,N_46620,N_46413);
or U48310 (N_48310,N_47159,N_47272);
nand U48311 (N_48311,N_47577,N_46933);
or U48312 (N_48312,N_46158,N_47835);
nand U48313 (N_48313,N_46832,N_46992);
xor U48314 (N_48314,N_47944,N_47270);
xor U48315 (N_48315,N_47196,N_46674);
and U48316 (N_48316,N_46321,N_46762);
nor U48317 (N_48317,N_47756,N_46196);
nor U48318 (N_48318,N_46312,N_47491);
xor U48319 (N_48319,N_46300,N_46379);
or U48320 (N_48320,N_47138,N_47353);
and U48321 (N_48321,N_46834,N_46178);
nor U48322 (N_48322,N_47493,N_47660);
nor U48323 (N_48323,N_47896,N_47834);
and U48324 (N_48324,N_46616,N_47878);
xor U48325 (N_48325,N_46317,N_46525);
xnor U48326 (N_48326,N_47618,N_46766);
and U48327 (N_48327,N_47790,N_47880);
or U48328 (N_48328,N_46671,N_46715);
xor U48329 (N_48329,N_47851,N_46489);
or U48330 (N_48330,N_47541,N_47650);
nand U48331 (N_48331,N_46737,N_46025);
or U48332 (N_48332,N_46979,N_46230);
or U48333 (N_48333,N_47175,N_47912);
nand U48334 (N_48334,N_47538,N_46778);
and U48335 (N_48335,N_46721,N_47918);
nand U48336 (N_48336,N_47854,N_47670);
xnor U48337 (N_48337,N_46971,N_46044);
nand U48338 (N_48338,N_46548,N_47914);
or U48339 (N_48339,N_47180,N_46274);
xnor U48340 (N_48340,N_47383,N_47899);
nand U48341 (N_48341,N_46538,N_46796);
nand U48342 (N_48342,N_46864,N_47148);
nand U48343 (N_48343,N_47664,N_46190);
and U48344 (N_48344,N_46609,N_46798);
and U48345 (N_48345,N_46611,N_46431);
xor U48346 (N_48346,N_46943,N_47682);
xor U48347 (N_48347,N_46858,N_46730);
xnor U48348 (N_48348,N_46438,N_46994);
xnor U48349 (N_48349,N_47646,N_47236);
nor U48350 (N_48350,N_46977,N_46692);
and U48351 (N_48351,N_47216,N_47125);
or U48352 (N_48352,N_47748,N_46399);
or U48353 (N_48353,N_47674,N_47698);
and U48354 (N_48354,N_47572,N_47108);
and U48355 (N_48355,N_47700,N_46187);
nand U48356 (N_48356,N_46452,N_47487);
nor U48357 (N_48357,N_47728,N_47637);
or U48358 (N_48358,N_47055,N_47832);
nand U48359 (N_48359,N_47153,N_46173);
nor U48360 (N_48360,N_47370,N_46801);
xnor U48361 (N_48361,N_47111,N_47500);
nand U48362 (N_48362,N_47023,N_46695);
nor U48363 (N_48363,N_47753,N_46700);
and U48364 (N_48364,N_46477,N_46397);
and U48365 (N_48365,N_47551,N_46517);
and U48366 (N_48366,N_46612,N_46151);
and U48367 (N_48367,N_46526,N_46369);
and U48368 (N_48368,N_47266,N_46782);
and U48369 (N_48369,N_47838,N_47143);
xor U48370 (N_48370,N_46245,N_47973);
nand U48371 (N_48371,N_46857,N_47021);
nand U48372 (N_48372,N_46436,N_46831);
nor U48373 (N_48373,N_46569,N_47668);
xor U48374 (N_48374,N_47939,N_47053);
nand U48375 (N_48375,N_46922,N_46974);
nand U48376 (N_48376,N_46942,N_46248);
nand U48377 (N_48377,N_47710,N_46593);
xor U48378 (N_48378,N_47995,N_47786);
xnor U48379 (N_48379,N_47877,N_47811);
and U48380 (N_48380,N_47449,N_46701);
and U48381 (N_48381,N_47502,N_46588);
xor U48382 (N_48382,N_46643,N_46707);
nand U48383 (N_48383,N_47599,N_46567);
nor U48384 (N_48384,N_47819,N_47355);
nand U48385 (N_48385,N_47015,N_47326);
nor U48386 (N_48386,N_47311,N_46243);
xnor U48387 (N_48387,N_46837,N_47429);
nor U48388 (N_48388,N_46799,N_46597);
or U48389 (N_48389,N_46156,N_46705);
and U48390 (N_48390,N_47620,N_47416);
or U48391 (N_48391,N_46608,N_47375);
xor U48392 (N_48392,N_47164,N_47365);
xnor U48393 (N_48393,N_46263,N_47469);
nand U48394 (N_48394,N_47519,N_47760);
and U48395 (N_48395,N_46824,N_46180);
nor U48396 (N_48396,N_46967,N_46165);
nand U48397 (N_48397,N_47349,N_47350);
nor U48398 (N_48398,N_46726,N_47402);
nor U48399 (N_48399,N_46986,N_46064);
nand U48400 (N_48400,N_46107,N_47413);
and U48401 (N_48401,N_46740,N_46405);
nand U48402 (N_48402,N_46690,N_46902);
xnor U48403 (N_48403,N_47068,N_46914);
and U48404 (N_48404,N_47130,N_46079);
or U48405 (N_48405,N_47304,N_46211);
nor U48406 (N_48406,N_47741,N_47097);
and U48407 (N_48407,N_46202,N_46870);
or U48408 (N_48408,N_47862,N_46224);
or U48409 (N_48409,N_47391,N_46972);
nand U48410 (N_48410,N_46068,N_46732);
or U48411 (N_48411,N_46866,N_47276);
and U48412 (N_48412,N_47940,N_47829);
nor U48413 (N_48413,N_47750,N_46468);
xnor U48414 (N_48414,N_46392,N_46556);
nand U48415 (N_48415,N_46335,N_46464);
nor U48416 (N_48416,N_47723,N_47545);
nand U48417 (N_48417,N_46736,N_47554);
or U48418 (N_48418,N_46550,N_46054);
or U48419 (N_48419,N_46653,N_47140);
nor U48420 (N_48420,N_47658,N_47583);
xor U48421 (N_48421,N_46303,N_47100);
nand U48422 (N_48422,N_47842,N_47150);
nor U48423 (N_48423,N_47533,N_47069);
xor U48424 (N_48424,N_46825,N_47734);
and U48425 (N_48425,N_46990,N_46031);
nor U48426 (N_48426,N_47222,N_46628);
and U48427 (N_48427,N_46167,N_47970);
nor U48428 (N_48428,N_46251,N_47929);
nor U48429 (N_48429,N_47961,N_47522);
or U48430 (N_48430,N_46580,N_47085);
nand U48431 (N_48431,N_47582,N_47705);
and U48432 (N_48432,N_46472,N_47243);
or U48433 (N_48433,N_46826,N_46874);
nand U48434 (N_48434,N_47223,N_47775);
and U48435 (N_48435,N_47736,N_46116);
nand U48436 (N_48436,N_46457,N_46794);
nor U48437 (N_48437,N_46275,N_46757);
and U48438 (N_48438,N_46347,N_46003);
nand U48439 (N_48439,N_47440,N_46561);
xnor U48440 (N_48440,N_47780,N_46282);
xor U48441 (N_48441,N_46049,N_47919);
and U48442 (N_48442,N_46889,N_47038);
xor U48443 (N_48443,N_47883,N_47517);
nand U48444 (N_48444,N_46817,N_47898);
nand U48445 (N_48445,N_46005,N_47724);
nand U48446 (N_48446,N_47812,N_46210);
and U48447 (N_48447,N_47256,N_46459);
nor U48448 (N_48448,N_46296,N_46461);
and U48449 (N_48449,N_46052,N_47557);
xnor U48450 (N_48450,N_46998,N_47604);
and U48451 (N_48451,N_47042,N_47481);
nand U48452 (N_48452,N_46214,N_47398);
nand U48453 (N_48453,N_47949,N_47220);
or U48454 (N_48454,N_46297,N_46913);
and U48455 (N_48455,N_47418,N_46966);
and U48456 (N_48456,N_47747,N_47793);
or U48457 (N_48457,N_47219,N_47866);
nor U48458 (N_48458,N_47496,N_47807);
nor U48459 (N_48459,N_46915,N_46505);
or U48460 (N_48460,N_46084,N_46219);
nand U48461 (N_48461,N_46946,N_46552);
or U48462 (N_48462,N_46754,N_47452);
or U48463 (N_48463,N_46761,N_46159);
xor U48464 (N_48464,N_46428,N_46513);
and U48465 (N_48465,N_47774,N_46423);
or U48466 (N_48466,N_46017,N_47316);
nand U48467 (N_48467,N_46877,N_47451);
and U48468 (N_48468,N_46823,N_47427);
xnor U48469 (N_48469,N_47739,N_47259);
or U48470 (N_48470,N_46033,N_46015);
nor U48471 (N_48471,N_47141,N_46481);
nor U48472 (N_48472,N_46501,N_46490);
nand U48473 (N_48473,N_47257,N_47709);
or U48474 (N_48474,N_46573,N_47292);
nor U48475 (N_48475,N_46742,N_47694);
or U48476 (N_48476,N_47732,N_47968);
nand U48477 (N_48477,N_46145,N_46846);
or U48478 (N_48478,N_47007,N_46931);
nor U48479 (N_48479,N_46125,N_46706);
or U48480 (N_48480,N_46166,N_46806);
nand U48481 (N_48481,N_47726,N_47512);
nor U48482 (N_48482,N_47116,N_47731);
nand U48483 (N_48483,N_47060,N_47328);
and U48484 (N_48484,N_47334,N_47621);
nor U48485 (N_48485,N_46018,N_47457);
xnor U48486 (N_48486,N_46661,N_47843);
xor U48487 (N_48487,N_46061,N_47539);
or U48488 (N_48488,N_46821,N_46558);
or U48489 (N_48489,N_46822,N_47247);
nand U48490 (N_48490,N_47531,N_47179);
or U48491 (N_48491,N_47076,N_47124);
xnor U48492 (N_48492,N_47945,N_46840);
xnor U48493 (N_48493,N_46383,N_46518);
xnor U48494 (N_48494,N_47537,N_46818);
nor U48495 (N_48495,N_46894,N_46735);
and U48496 (N_48496,N_46919,N_46615);
xor U48497 (N_48497,N_47789,N_47014);
or U48498 (N_48498,N_46932,N_47894);
xnor U48499 (N_48499,N_47563,N_46900);
and U48500 (N_48500,N_46326,N_46698);
xor U48501 (N_48501,N_46584,N_46486);
nor U48502 (N_48502,N_47281,N_47985);
nor U48503 (N_48503,N_47569,N_47359);
nor U48504 (N_48504,N_47089,N_46137);
and U48505 (N_48505,N_46485,N_46918);
nand U48506 (N_48506,N_46759,N_46659);
nor U48507 (N_48507,N_47672,N_47977);
nand U48508 (N_48508,N_47036,N_47265);
nor U48509 (N_48509,N_46318,N_47874);
nand U48510 (N_48510,N_46095,N_47342);
xnor U48511 (N_48511,N_46028,N_47149);
nor U48512 (N_48512,N_46030,N_46999);
nor U48513 (N_48513,N_46089,N_46433);
and U48514 (N_48514,N_46592,N_47302);
xnor U48515 (N_48515,N_46655,N_47466);
nand U48516 (N_48516,N_46099,N_47872);
nand U48517 (N_48517,N_47260,N_46443);
and U48518 (N_48518,N_46540,N_46551);
nor U48519 (N_48519,N_47687,N_47540);
and U48520 (N_48520,N_46498,N_46908);
nor U48521 (N_48521,N_46716,N_46389);
xnor U48522 (N_48522,N_47921,N_47598);
nor U48523 (N_48523,N_46533,N_47489);
nor U48524 (N_48524,N_47850,N_47109);
xor U48525 (N_48525,N_46903,N_47226);
or U48526 (N_48526,N_47721,N_46553);
nor U48527 (N_48527,N_46043,N_46528);
nand U48528 (N_48528,N_46752,N_46262);
or U48529 (N_48529,N_47762,N_46805);
or U48530 (N_48530,N_47636,N_47479);
and U48531 (N_48531,N_46133,N_46771);
nor U48532 (N_48532,N_46780,N_46184);
nor U48533 (N_48533,N_47640,N_47564);
and U48534 (N_48534,N_46949,N_46934);
nor U48535 (N_48535,N_46235,N_46880);
nand U48536 (N_48536,N_46193,N_47408);
nor U48537 (N_48537,N_47423,N_46978);
or U48538 (N_48538,N_46375,N_47767);
xor U48539 (N_48539,N_46055,N_46080);
nand U48540 (N_48540,N_46495,N_46140);
and U48541 (N_48541,N_47578,N_46100);
or U48542 (N_48542,N_47667,N_46062);
nand U48543 (N_48543,N_47662,N_46865);
or U48544 (N_48544,N_46280,N_46420);
nor U48545 (N_48545,N_46170,N_47320);
nor U48546 (N_48546,N_47993,N_46702);
or U48547 (N_48547,N_46812,N_47910);
nor U48548 (N_48548,N_47879,N_47857);
xnor U48549 (N_48549,N_46638,N_47040);
and U48550 (N_48550,N_47170,N_46893);
or U48551 (N_48551,N_46154,N_46119);
or U48552 (N_48552,N_46176,N_46647);
and U48553 (N_48553,N_46788,N_47073);
nor U48554 (N_48554,N_47474,N_47987);
and U48555 (N_48555,N_46272,N_46847);
nor U48556 (N_48556,N_46487,N_46637);
nor U48557 (N_48557,N_46745,N_46381);
and U48558 (N_48558,N_47523,N_47571);
or U48559 (N_48559,N_47613,N_46332);
nand U48560 (N_48560,N_46594,N_47378);
or U48561 (N_48561,N_47411,N_47160);
nand U48562 (N_48562,N_46688,N_46827);
nand U48563 (N_48563,N_46901,N_46662);
and U48564 (N_48564,N_46494,N_46400);
and U48565 (N_48565,N_46694,N_46032);
and U48566 (N_48566,N_46203,N_47924);
xor U48567 (N_48567,N_46474,N_47258);
xnor U48568 (N_48568,N_46970,N_47133);
and U48569 (N_48569,N_46510,N_46581);
xor U48570 (N_48570,N_46432,N_47956);
and U48571 (N_48571,N_47959,N_47555);
nor U48572 (N_48572,N_47347,N_46102);
xnor U48573 (N_48573,N_47279,N_47476);
nor U48574 (N_48574,N_46767,N_47781);
and U48575 (N_48575,N_46019,N_46511);
and U48576 (N_48576,N_46623,N_47952);
nor U48577 (N_48577,N_47098,N_46677);
or U48578 (N_48578,N_47974,N_47942);
and U48579 (N_48579,N_46777,N_47560);
or U48580 (N_48580,N_47132,N_46359);
nor U48581 (N_48581,N_47364,N_46406);
and U48582 (N_48582,N_47567,N_47101);
xor U48583 (N_48583,N_47703,N_47881);
xor U48584 (N_48584,N_46259,N_46691);
and U48585 (N_48585,N_47791,N_47117);
nor U48586 (N_48586,N_46414,N_46634);
xnor U48587 (N_48587,N_46021,N_47146);
or U48588 (N_48588,N_47030,N_47022);
nor U48589 (N_48589,N_47743,N_47465);
nand U48590 (N_48590,N_46346,N_46097);
nor U48591 (N_48591,N_47210,N_46228);
or U48592 (N_48592,N_46534,N_46284);
nand U48593 (N_48593,N_46129,N_47840);
or U48594 (N_48594,N_46532,N_47400);
xor U48595 (N_48595,N_46508,N_47579);
and U48596 (N_48596,N_47630,N_47815);
nand U48597 (N_48597,N_46828,N_46529);
nor U48598 (N_48598,N_46278,N_47492);
xnor U48599 (N_48599,N_47782,N_46802);
or U48600 (N_48600,N_46155,N_46388);
nand U48601 (N_48601,N_47831,N_47368);
nor U48602 (N_48602,N_46342,N_47957);
nor U48603 (N_48603,N_46384,N_46071);
nor U48604 (N_48604,N_46941,N_47254);
nor U48605 (N_48605,N_47082,N_46639);
nor U48606 (N_48606,N_46034,N_46753);
xor U48607 (N_48607,N_47443,N_47948);
nor U48608 (N_48608,N_46189,N_47562);
nand U48609 (N_48609,N_46276,N_47313);
and U48610 (N_48610,N_46144,N_46304);
xnor U48611 (N_48611,N_47000,N_46566);
nand U48612 (N_48612,N_47695,N_47610);
nor U48613 (N_48613,N_46562,N_46221);
nand U48614 (N_48614,N_46961,N_47168);
xnor U48615 (N_48615,N_47186,N_46565);
or U48616 (N_48616,N_46878,N_47947);
and U48617 (N_48617,N_46571,N_47461);
nand U48618 (N_48618,N_47019,N_46804);
nor U48619 (N_48619,N_47071,N_46269);
or U48620 (N_48620,N_46004,N_46314);
xnor U48621 (N_48621,N_47444,N_46354);
nand U48622 (N_48622,N_47385,N_46965);
nand U48623 (N_48623,N_46570,N_47833);
xor U48624 (N_48624,N_47433,N_46585);
or U48625 (N_48625,N_46657,N_47006);
nor U48626 (N_48626,N_47371,N_46624);
nand U48627 (N_48627,N_46087,N_46599);
or U48628 (N_48628,N_47363,N_47299);
or U48629 (N_48629,N_47185,N_46925);
nand U48630 (N_48630,N_47655,N_47447);
nor U48631 (N_48631,N_46040,N_47145);
nand U48632 (N_48632,N_47330,N_46717);
and U48633 (N_48633,N_46744,N_47626);
nor U48634 (N_48634,N_47642,N_47963);
and U48635 (N_48635,N_46625,N_46123);
nor U48636 (N_48636,N_46853,N_47483);
nand U48637 (N_48637,N_47337,N_47809);
and U48638 (N_48638,N_46239,N_46743);
and U48639 (N_48639,N_47264,N_46065);
nor U48640 (N_48640,N_46252,N_47776);
xor U48641 (N_48641,N_47629,N_46969);
and U48642 (N_48642,N_46554,N_47876);
nor U48643 (N_48643,N_46727,N_46514);
and U48644 (N_48644,N_46343,N_47392);
and U48645 (N_48645,N_46987,N_47156);
or U48646 (N_48646,N_47158,N_47511);
nand U48647 (N_48647,N_46791,N_47984);
nor U48648 (N_48648,N_46215,N_47490);
xnor U48649 (N_48649,N_46772,N_46349);
nor U48650 (N_48650,N_47841,N_47093);
xnor U48651 (N_48651,N_47839,N_47396);
or U48652 (N_48652,N_46357,N_47283);
nand U48653 (N_48653,N_47399,N_47596);
xnor U48654 (N_48654,N_46220,N_47603);
and U48655 (N_48655,N_47643,N_47057);
nand U48656 (N_48656,N_46171,N_47902);
or U48657 (N_48657,N_46663,N_46760);
and U48658 (N_48658,N_47020,N_47005);
and U48659 (N_48659,N_47553,N_46201);
or U48660 (N_48660,N_46046,N_47002);
nand U48661 (N_48661,N_46957,N_47889);
nor U48662 (N_48662,N_47043,N_47501);
nand U48663 (N_48663,N_46430,N_46680);
nand U48664 (N_48664,N_46868,N_46773);
and U48665 (N_48665,N_47892,N_46522);
and U48666 (N_48666,N_46236,N_47322);
nand U48667 (N_48667,N_47163,N_46483);
or U48668 (N_48668,N_46410,N_47930);
xor U48669 (N_48669,N_46309,N_46984);
nor U48670 (N_48670,N_47923,N_47003);
nor U48671 (N_48671,N_46512,N_46939);
xnor U48672 (N_48672,N_47103,N_47339);
nor U48673 (N_48673,N_47628,N_46530);
nor U48674 (N_48674,N_47297,N_47432);
or U48675 (N_48675,N_47980,N_46976);
xor U48676 (N_48676,N_47925,N_47638);
nor U48677 (N_48677,N_47250,N_47943);
and U48678 (N_48678,N_47719,N_46378);
xnor U48679 (N_48679,N_46076,N_47269);
and U48680 (N_48680,N_46036,N_46586);
and U48681 (N_48681,N_47460,N_47120);
nor U48682 (N_48682,N_47676,N_47262);
xor U48683 (N_48683,N_46656,N_47004);
nand U48684 (N_48684,N_47552,N_47456);
nand U48685 (N_48685,N_46163,N_46975);
and U48686 (N_48686,N_47908,N_46118);
or U48687 (N_48687,N_47666,N_47195);
nor U48688 (N_48688,N_47615,N_47445);
and U48689 (N_48689,N_47981,N_47244);
nor U48690 (N_48690,N_47434,N_47240);
nand U48691 (N_48691,N_46515,N_46393);
nor U48692 (N_48692,N_47380,N_46277);
and U48693 (N_48693,N_46233,N_47191);
nand U48694 (N_48694,N_47091,N_46895);
nand U48695 (N_48695,N_46829,N_47287);
and U48696 (N_48696,N_46687,N_46291);
or U48697 (N_48697,N_46904,N_47464);
and U48698 (N_48698,N_47858,N_47430);
xnor U48699 (N_48699,N_47335,N_46935);
and U48700 (N_48700,N_46996,N_46478);
nor U48701 (N_48701,N_46631,N_47605);
and U48702 (N_48702,N_47468,N_46168);
or U48703 (N_48703,N_47882,N_47931);
and U48704 (N_48704,N_47074,N_46150);
or U48705 (N_48705,N_47651,N_47752);
nor U48706 (N_48706,N_47966,N_47907);
and U48707 (N_48707,N_46758,N_46339);
and U48708 (N_48708,N_46607,N_47084);
and U48709 (N_48709,N_47454,N_47234);
nand U48710 (N_48710,N_47307,N_47301);
xor U48711 (N_48711,N_46626,N_46862);
or U48712 (N_48712,N_47412,N_46385);
or U48713 (N_48713,N_46418,N_47333);
and U48714 (N_48714,N_46271,N_47988);
nand U48715 (N_48715,N_47369,N_47305);
nand U48716 (N_48716,N_46813,N_47573);
nor U48717 (N_48717,N_47294,N_47773);
or U48718 (N_48718,N_46108,N_47594);
and U48719 (N_48719,N_46629,N_47574);
xnor U48720 (N_48720,N_46353,N_46591);
nand U48721 (N_48721,N_46854,N_46619);
nand U48722 (N_48722,N_46873,N_47837);
nor U48723 (N_48723,N_47309,N_47177);
and U48724 (N_48724,N_47758,N_46037);
and U48725 (N_48725,N_46708,N_47848);
nor U48726 (N_48726,N_47600,N_47306);
or U48727 (N_48727,N_47544,N_47631);
nor U48728 (N_48728,N_46983,N_46650);
xnor U48729 (N_48729,N_47515,N_47123);
and U48730 (N_48730,N_47106,N_47616);
nor U48731 (N_48731,N_47386,N_47697);
and U48732 (N_48732,N_47187,N_47063);
xor U48733 (N_48733,N_47139,N_47052);
or U48734 (N_48734,N_46134,N_47329);
and U48735 (N_48735,N_46286,N_46337);
nor U48736 (N_48736,N_47426,N_46491);
and U48737 (N_48737,N_46797,N_46559);
and U48738 (N_48738,N_46141,N_46411);
or U48739 (N_48739,N_46930,N_46995);
nand U48740 (N_48740,N_47012,N_47964);
and U48741 (N_48741,N_46524,N_46240);
nor U48742 (N_48742,N_47797,N_47171);
xor U48743 (N_48743,N_47405,N_46787);
nor U48744 (N_48744,N_46681,N_46795);
nand U48745 (N_48745,N_47548,N_47494);
nand U48746 (N_48746,N_47325,N_47725);
xor U48747 (N_48747,N_46666,N_46728);
xnor U48748 (N_48748,N_46440,N_46352);
nor U48749 (N_48749,N_46081,N_46417);
and U48750 (N_48750,N_46345,N_47275);
nor U48751 (N_48751,N_47828,N_46195);
and U48752 (N_48752,N_47846,N_47808);
nor U48753 (N_48753,N_46008,N_46216);
or U48754 (N_48754,N_46330,N_46649);
nor U48755 (N_48755,N_46368,N_47470);
nand U48756 (N_48756,N_46572,N_47542);
and U48757 (N_48757,N_46143,N_47612);
xnor U48758 (N_48758,N_46741,N_47338);
and U48759 (N_48759,N_47678,N_46212);
or U48760 (N_48760,N_46682,N_47641);
and U48761 (N_48761,N_46009,N_46002);
or U48762 (N_48762,N_46685,N_47181);
xor U48763 (N_48763,N_46131,N_47455);
nand U48764 (N_48764,N_47787,N_46366);
nor U48765 (N_48765,N_46774,N_47746);
nand U48766 (N_48766,N_47777,N_46852);
xnor U48767 (N_48767,N_46577,N_46668);
or U48768 (N_48768,N_46205,N_46644);
or U48769 (N_48769,N_46439,N_46407);
nand U48770 (N_48770,N_47606,N_47953);
or U48771 (N_48771,N_46006,N_47609);
xor U48772 (N_48772,N_47836,N_47267);
nor U48773 (N_48773,N_47729,N_46026);
nand U48774 (N_48774,N_47534,N_47209);
or U48775 (N_48775,N_47388,N_47448);
xor U48776 (N_48776,N_46290,N_47206);
or U48777 (N_48777,N_47169,N_47686);
xor U48778 (N_48778,N_47485,N_46576);
nand U48779 (N_48779,N_46261,N_47441);
xor U48780 (N_48780,N_46109,N_46419);
or U48781 (N_48781,N_47054,N_47308);
nand U48782 (N_48782,N_47979,N_47336);
nor U48783 (N_48783,N_47801,N_47011);
or U48784 (N_48784,N_47784,N_46063);
nor U48785 (N_48785,N_47608,N_46603);
nor U48786 (N_48786,N_46527,N_47367);
and U48787 (N_48787,N_46993,N_47415);
xor U48788 (N_48788,N_46246,N_46001);
and U48789 (N_48789,N_46912,N_46465);
nor U48790 (N_48790,N_46444,N_47025);
and U48791 (N_48791,N_47690,N_46441);
or U48792 (N_48792,N_47607,N_46539);
nor U48793 (N_48793,N_46683,N_47128);
or U48794 (N_48794,N_47887,N_47765);
nor U48795 (N_48795,N_47675,N_46557);
nand U48796 (N_48796,N_46546,N_46329);
and U48797 (N_48797,N_46088,N_46689);
nand U48798 (N_48798,N_46324,N_46038);
xnor U48799 (N_48799,N_46606,N_47165);
nand U48800 (N_48800,N_47677,N_46968);
nand U48801 (N_48801,N_46496,N_46836);
nand U48802 (N_48802,N_47176,N_47332);
nor U48803 (N_48803,N_46382,N_46362);
nand U48804 (N_48804,N_47389,N_47975);
nor U48805 (N_48805,N_47590,N_47885);
xnor U48806 (N_48806,N_46194,N_46916);
or U48807 (N_48807,N_46422,N_46755);
xor U48808 (N_48808,N_46911,N_47649);
xnor U48809 (N_48809,N_47529,N_47965);
nor U48810 (N_48810,N_46842,N_47031);
or U48811 (N_48811,N_46848,N_46174);
nor U48812 (N_48812,N_47193,N_47495);
nor U48813 (N_48813,N_47934,N_46699);
or U48814 (N_48814,N_47323,N_47096);
xor U48815 (N_48815,N_47659,N_47715);
or U48816 (N_48816,N_47439,N_47428);
xor U48817 (N_48817,N_47058,N_46973);
or U48818 (N_48818,N_47189,N_47516);
nand U48819 (N_48819,N_46958,N_46237);
nor U48820 (N_48820,N_46197,N_46020);
and U48821 (N_48821,N_47950,N_47634);
nor U48822 (N_48822,N_46664,N_46112);
and U48823 (N_48823,N_46633,N_46860);
and U48824 (N_48824,N_46844,N_46327);
and U48825 (N_48825,N_47813,N_47920);
or U48826 (N_48826,N_47989,N_46959);
xor U48827 (N_48827,N_47274,N_47147);
nor U48828 (N_48828,N_47768,N_46928);
or U48829 (N_48829,N_46404,N_47424);
nor U48830 (N_48830,N_47933,N_46035);
nand U48831 (N_48831,N_46940,N_46722);
and U48832 (N_48832,N_47008,N_46504);
nand U48833 (N_48833,N_47437,N_47419);
and U48834 (N_48834,N_47295,N_47827);
nand U48835 (N_48835,N_47471,N_47102);
xnor U48836 (N_48836,N_47558,N_46091);
nand U48837 (N_48837,N_47696,N_46598);
or U48838 (N_48838,N_47853,N_46455);
or U48839 (N_48839,N_46313,N_46814);
nand U48840 (N_48840,N_47757,N_46905);
and U48841 (N_48841,N_47903,N_46590);
or U48842 (N_48842,N_47992,N_46355);
and U48843 (N_48843,N_46363,N_46200);
nand U48844 (N_48844,N_47228,N_46989);
xor U48845 (N_48845,N_46830,N_47720);
or U48846 (N_48846,N_46956,N_47273);
xor U48847 (N_48847,N_46784,N_47810);
or U48848 (N_48848,N_47230,N_47994);
nor U48849 (N_48849,N_47351,N_46258);
nor U48850 (N_48850,N_47602,N_47344);
nor U48851 (N_48851,N_47414,N_46906);
nand U48852 (N_48852,N_47233,N_47830);
nand U48853 (N_48853,N_46285,N_47113);
xnor U48854 (N_48854,N_46578,N_47673);
nor U48855 (N_48855,N_47245,N_47154);
and U48856 (N_48856,N_47683,N_47467);
xor U48857 (N_48857,N_47356,N_46897);
and U48858 (N_48858,N_47806,N_46191);
xnor U48859 (N_48859,N_46614,N_47507);
nand U48860 (N_48860,N_46206,N_47869);
and U48861 (N_48861,N_47733,N_46458);
or U48862 (N_48862,N_46627,N_47362);
nor U48863 (N_48863,N_46238,N_46516);
or U48864 (N_48864,N_47227,N_46749);
or U48865 (N_48865,N_46820,N_46207);
xor U48866 (N_48866,N_46786,N_46217);
or U48867 (N_48867,N_46022,N_46756);
xnor U48868 (N_48868,N_46186,N_46450);
nand U48869 (N_48869,N_47549,N_47017);
nand U48870 (N_48870,N_46587,N_47016);
nand U48871 (N_48871,N_46073,N_47104);
or U48872 (N_48872,N_46537,N_46579);
nand U48873 (N_48873,N_47112,N_47249);
nor U48874 (N_48874,N_47849,N_47463);
and U48875 (N_48875,N_46106,N_47136);
nor U48876 (N_48876,N_47248,N_47821);
xor U48877 (N_48877,N_46747,N_46850);
or U48878 (N_48878,N_47121,N_46636);
or U48879 (N_48879,N_46254,N_46867);
nand U48880 (N_48880,N_46678,N_46298);
nor U48881 (N_48881,N_47589,N_46531);
nor U48882 (N_48882,N_46302,N_47754);
or U48883 (N_48883,N_46838,N_46898);
and U48884 (N_48884,N_46560,N_46927);
nor U48885 (N_48885,N_46351,N_46092);
xor U48886 (N_48886,N_46066,N_47473);
and U48887 (N_48887,N_46670,N_46660);
xor U48888 (N_48888,N_46497,N_46126);
nand U48889 (N_48889,N_46672,N_46693);
xor U48890 (N_48890,N_47525,N_46148);
or U48891 (N_48891,N_46164,N_46535);
or U48892 (N_48892,N_47395,N_46281);
or U48893 (N_48893,N_46283,N_47888);
nor U48894 (N_48894,N_47478,N_46582);
or U48895 (N_48895,N_46391,N_47237);
nor U48896 (N_48896,N_47527,N_46673);
xnor U48897 (N_48897,N_47597,N_46781);
and U48898 (N_48898,N_47354,N_46712);
xnor U48899 (N_48899,N_47802,N_46060);
or U48900 (N_48900,N_47135,N_46507);
and U48901 (N_48901,N_46768,N_47873);
and U48902 (N_48902,N_46482,N_46710);
and U48903 (N_48903,N_46921,N_47235);
or U48904 (N_48904,N_47268,N_47911);
or U48905 (N_48905,N_46260,N_46048);
and U48906 (N_48906,N_47289,N_47661);
nand U48907 (N_48907,N_46861,N_47625);
nand U48908 (N_48908,N_46310,N_46070);
and U48909 (N_48909,N_46086,N_47026);
or U48910 (N_48910,N_46765,N_46648);
nor U48911 (N_48911,N_47566,N_47066);
nor U48912 (N_48912,N_47035,N_46415);
xnor U48913 (N_48913,N_46067,N_46429);
or U48914 (N_48914,N_47286,N_46589);
nor U48915 (N_48915,N_46883,N_46751);
nor U48916 (N_48916,N_47859,N_47033);
nor U48917 (N_48917,N_47509,N_47293);
xor U48918 (N_48918,N_46618,N_46075);
nor U48919 (N_48919,N_47595,N_46621);
nand U48920 (N_48920,N_46402,N_46234);
nor U48921 (N_48921,N_46955,N_46253);
or U48922 (N_48922,N_46050,N_47045);
and U48923 (N_48923,N_46803,N_46792);
nor U48924 (N_48924,N_47277,N_47319);
xnor U48925 (N_48925,N_46839,N_46891);
nand U48926 (N_48926,N_46085,N_46859);
or U48927 (N_48927,N_46734,N_47817);
nand U48928 (N_48928,N_47614,N_47712);
nand U48929 (N_48929,N_47404,N_47788);
nand U48930 (N_48930,N_46467,N_47092);
or U48931 (N_48931,N_47324,N_46390);
nand U48932 (N_48932,N_47937,N_46437);
nand U48933 (N_48933,N_46320,N_46454);
nor U48934 (N_48934,N_47684,N_46920);
or U48935 (N_48935,N_47632,N_47498);
or U48936 (N_48936,N_47745,N_47584);
and U48937 (N_48937,N_46287,N_47211);
and U48938 (N_48938,N_46574,N_47708);
and U48939 (N_48939,N_47619,N_47735);
xor U48940 (N_48940,N_46953,N_47127);
nand U48941 (N_48941,N_46344,N_47480);
or U48942 (N_48942,N_47580,N_46157);
nor U48943 (N_48943,N_47738,N_47051);
nand U48944 (N_48944,N_47706,N_47032);
nor U48945 (N_48945,N_46630,N_47972);
and U48946 (N_48946,N_46833,N_47129);
nor U48947 (N_48947,N_47893,N_46887);
nand U48948 (N_48948,N_46110,N_47520);
and U48949 (N_48949,N_47576,N_47105);
and U48950 (N_48950,N_47904,N_47047);
nand U48951 (N_48951,N_46642,N_47056);
nor U48952 (N_48952,N_46447,N_47251);
and U48953 (N_48953,N_46386,N_47119);
nand U48954 (N_48954,N_46142,N_46307);
and U48955 (N_48955,N_46896,N_46121);
or U48956 (N_48956,N_47315,N_46841);
and U48957 (N_48957,N_47951,N_47962);
or U48958 (N_48958,N_46997,N_46809);
or U48959 (N_48959,N_46185,N_47559);
or U48960 (N_48960,N_46127,N_47932);
or U48961 (N_48961,N_46083,N_46331);
nor U48962 (N_48962,N_47820,N_47144);
nand U48963 (N_48963,N_46069,N_46471);
nor U48964 (N_48964,N_46425,N_47366);
or U48965 (N_48965,N_47072,N_47061);
and U48966 (N_48966,N_46380,N_46306);
xor U48967 (N_48967,N_46416,N_47860);
nand U48968 (N_48968,N_46000,N_47623);
or U48969 (N_48969,N_47261,N_47847);
and U48970 (N_48970,N_47740,N_46600);
xor U48971 (N_48971,N_46988,N_47314);
or U48972 (N_48972,N_47890,N_47253);
or U48973 (N_48973,N_47151,N_47954);
xnor U48974 (N_48974,N_47639,N_46856);
nand U48975 (N_48975,N_47034,N_46250);
xor U48976 (N_48976,N_46094,N_46041);
nand U48977 (N_48977,N_46929,N_47867);
xnor U48978 (N_48978,N_46372,N_46289);
nand U48979 (N_48979,N_47318,N_46090);
or U48980 (N_48980,N_46808,N_47221);
xnor U48981 (N_48981,N_46012,N_46944);
nand U48982 (N_48982,N_47865,N_46117);
nor U48983 (N_48983,N_46981,N_47229);
nand U48984 (N_48984,N_47680,N_46456);
and U48985 (N_48985,N_46448,N_46583);
nor U48986 (N_48986,N_46733,N_47134);
nand U48987 (N_48987,N_46602,N_46132);
or U48988 (N_48988,N_46011,N_47722);
and U48989 (N_48989,N_46292,N_46007);
and U48990 (N_48990,N_47717,N_47062);
nor U48991 (N_48991,N_47986,N_46103);
xnor U48992 (N_48992,N_47928,N_47742);
xor U48993 (N_48993,N_47373,N_47656);
and U48994 (N_48994,N_47804,N_46288);
xor U48995 (N_48995,N_46373,N_47588);
and U48996 (N_48996,N_46056,N_46899);
or U48997 (N_48997,N_47617,N_46950);
xnor U48998 (N_48998,N_46294,N_47212);
nor U48999 (N_48999,N_46279,N_46115);
or U49000 (N_49000,N_46605,N_46273);
and U49001 (N_49001,N_47945,N_47497);
nor U49002 (N_49002,N_46087,N_47593);
or U49003 (N_49003,N_47996,N_47541);
and U49004 (N_49004,N_47802,N_46258);
and U49005 (N_49005,N_46772,N_46873);
or U49006 (N_49006,N_47517,N_47290);
or U49007 (N_49007,N_46873,N_47472);
nor U49008 (N_49008,N_46047,N_47904);
and U49009 (N_49009,N_46703,N_47693);
nor U49010 (N_49010,N_46682,N_46141);
or U49011 (N_49011,N_46800,N_47420);
nor U49012 (N_49012,N_47916,N_46918);
nor U49013 (N_49013,N_46106,N_47509);
xor U49014 (N_49014,N_47037,N_47720);
nand U49015 (N_49015,N_46666,N_47883);
and U49016 (N_49016,N_47082,N_46077);
xor U49017 (N_49017,N_47078,N_47057);
nand U49018 (N_49018,N_47466,N_46958);
nor U49019 (N_49019,N_46356,N_47926);
and U49020 (N_49020,N_47250,N_47296);
or U49021 (N_49021,N_46005,N_47612);
xor U49022 (N_49022,N_47683,N_46451);
nor U49023 (N_49023,N_46980,N_47704);
nand U49024 (N_49024,N_46536,N_47399);
xnor U49025 (N_49025,N_47488,N_46310);
xor U49026 (N_49026,N_47472,N_46374);
or U49027 (N_49027,N_47995,N_47347);
nand U49028 (N_49028,N_47719,N_46988);
nand U49029 (N_49029,N_46754,N_47868);
or U49030 (N_49030,N_46985,N_46511);
xnor U49031 (N_49031,N_46149,N_46022);
nor U49032 (N_49032,N_46076,N_47608);
xnor U49033 (N_49033,N_46562,N_47325);
xnor U49034 (N_49034,N_46640,N_47454);
nor U49035 (N_49035,N_46423,N_46869);
and U49036 (N_49036,N_47116,N_47412);
nand U49037 (N_49037,N_46418,N_47517);
and U49038 (N_49038,N_46865,N_47572);
xnor U49039 (N_49039,N_47747,N_47827);
or U49040 (N_49040,N_47406,N_47405);
xnor U49041 (N_49041,N_47530,N_46935);
and U49042 (N_49042,N_47171,N_46234);
or U49043 (N_49043,N_46059,N_46255);
xor U49044 (N_49044,N_47270,N_46379);
xor U49045 (N_49045,N_47372,N_46368);
nor U49046 (N_49046,N_46669,N_47389);
xor U49047 (N_49047,N_46964,N_47581);
and U49048 (N_49048,N_46139,N_46061);
nor U49049 (N_49049,N_46648,N_47812);
or U49050 (N_49050,N_46440,N_47909);
xnor U49051 (N_49051,N_46537,N_47529);
xor U49052 (N_49052,N_47116,N_46387);
and U49053 (N_49053,N_46644,N_46167);
nor U49054 (N_49054,N_46240,N_47100);
and U49055 (N_49055,N_46515,N_47469);
nor U49056 (N_49056,N_47836,N_46695);
nand U49057 (N_49057,N_47330,N_47152);
or U49058 (N_49058,N_46256,N_46462);
nand U49059 (N_49059,N_46301,N_46916);
nor U49060 (N_49060,N_46293,N_47453);
xor U49061 (N_49061,N_47105,N_47052);
nand U49062 (N_49062,N_47838,N_47706);
xnor U49063 (N_49063,N_47983,N_46938);
xnor U49064 (N_49064,N_46974,N_47422);
and U49065 (N_49065,N_47467,N_46290);
nor U49066 (N_49066,N_47996,N_47547);
nor U49067 (N_49067,N_47179,N_46938);
xor U49068 (N_49068,N_47924,N_46348);
and U49069 (N_49069,N_47935,N_46182);
nand U49070 (N_49070,N_47770,N_46239);
or U49071 (N_49071,N_46910,N_46705);
nor U49072 (N_49072,N_46473,N_47070);
nor U49073 (N_49073,N_46659,N_46718);
and U49074 (N_49074,N_47213,N_47994);
nand U49075 (N_49075,N_46216,N_46502);
nand U49076 (N_49076,N_46457,N_46592);
or U49077 (N_49077,N_46635,N_46706);
or U49078 (N_49078,N_46521,N_46207);
xor U49079 (N_49079,N_46357,N_47877);
xnor U49080 (N_49080,N_47018,N_47839);
and U49081 (N_49081,N_46126,N_47418);
and U49082 (N_49082,N_46711,N_46255);
nand U49083 (N_49083,N_46210,N_46047);
nand U49084 (N_49084,N_47332,N_46987);
xnor U49085 (N_49085,N_47261,N_46677);
xnor U49086 (N_49086,N_46048,N_47998);
nor U49087 (N_49087,N_47416,N_47243);
and U49088 (N_49088,N_47365,N_46425);
and U49089 (N_49089,N_46593,N_46463);
and U49090 (N_49090,N_47785,N_47875);
nor U49091 (N_49091,N_47651,N_46297);
xor U49092 (N_49092,N_46256,N_47752);
nand U49093 (N_49093,N_46234,N_47658);
and U49094 (N_49094,N_46683,N_46989);
nand U49095 (N_49095,N_46337,N_46999);
and U49096 (N_49096,N_46691,N_47584);
or U49097 (N_49097,N_47916,N_47214);
xor U49098 (N_49098,N_46371,N_47387);
xor U49099 (N_49099,N_46811,N_46087);
xor U49100 (N_49100,N_46339,N_46162);
and U49101 (N_49101,N_47444,N_47308);
and U49102 (N_49102,N_47853,N_46740);
xnor U49103 (N_49103,N_47355,N_47145);
nand U49104 (N_49104,N_47234,N_47092);
nor U49105 (N_49105,N_46077,N_47809);
nand U49106 (N_49106,N_46161,N_47559);
xor U49107 (N_49107,N_47126,N_46193);
nand U49108 (N_49108,N_46589,N_47289);
and U49109 (N_49109,N_47443,N_46182);
nor U49110 (N_49110,N_47487,N_46139);
nor U49111 (N_49111,N_46753,N_47900);
and U49112 (N_49112,N_46547,N_46729);
nand U49113 (N_49113,N_46103,N_47033);
and U49114 (N_49114,N_47351,N_47886);
xor U49115 (N_49115,N_47650,N_47170);
xnor U49116 (N_49116,N_46412,N_47065);
nand U49117 (N_49117,N_46494,N_46764);
or U49118 (N_49118,N_46383,N_46961);
and U49119 (N_49119,N_46316,N_47701);
nor U49120 (N_49120,N_47746,N_47564);
or U49121 (N_49121,N_47492,N_47121);
and U49122 (N_49122,N_46567,N_46136);
xnor U49123 (N_49123,N_47213,N_46337);
and U49124 (N_49124,N_46416,N_46771);
and U49125 (N_49125,N_47032,N_46899);
xnor U49126 (N_49126,N_47415,N_47594);
or U49127 (N_49127,N_47021,N_46485);
nor U49128 (N_49128,N_47913,N_47960);
or U49129 (N_49129,N_46666,N_47424);
nand U49130 (N_49130,N_46318,N_47821);
nor U49131 (N_49131,N_46579,N_46680);
nand U49132 (N_49132,N_47264,N_46479);
or U49133 (N_49133,N_47809,N_47559);
and U49134 (N_49134,N_46257,N_47830);
xnor U49135 (N_49135,N_46932,N_47356);
xor U49136 (N_49136,N_46638,N_47020);
or U49137 (N_49137,N_47264,N_47137);
or U49138 (N_49138,N_47695,N_47467);
nand U49139 (N_49139,N_47960,N_46157);
or U49140 (N_49140,N_47011,N_46819);
nor U49141 (N_49141,N_47422,N_46902);
or U49142 (N_49142,N_46076,N_47475);
nand U49143 (N_49143,N_47781,N_47111);
nand U49144 (N_49144,N_47291,N_47266);
xor U49145 (N_49145,N_47783,N_46259);
xnor U49146 (N_49146,N_47405,N_46584);
and U49147 (N_49147,N_46705,N_46787);
xnor U49148 (N_49148,N_47007,N_47864);
xnor U49149 (N_49149,N_47619,N_46780);
xor U49150 (N_49150,N_47682,N_46454);
nor U49151 (N_49151,N_46842,N_47671);
nor U49152 (N_49152,N_47300,N_47826);
or U49153 (N_49153,N_46622,N_46250);
or U49154 (N_49154,N_46499,N_47483);
nor U49155 (N_49155,N_46673,N_47222);
nor U49156 (N_49156,N_46364,N_46739);
nand U49157 (N_49157,N_47162,N_47521);
nor U49158 (N_49158,N_47150,N_47537);
xor U49159 (N_49159,N_46518,N_47610);
xor U49160 (N_49160,N_46880,N_47968);
and U49161 (N_49161,N_47567,N_47995);
nand U49162 (N_49162,N_46847,N_47145);
or U49163 (N_49163,N_47254,N_46494);
nor U49164 (N_49164,N_46309,N_46748);
nor U49165 (N_49165,N_46837,N_47713);
or U49166 (N_49166,N_47126,N_46508);
nor U49167 (N_49167,N_47206,N_47672);
or U49168 (N_49168,N_46491,N_47132);
nor U49169 (N_49169,N_47931,N_46262);
or U49170 (N_49170,N_47612,N_46479);
and U49171 (N_49171,N_47211,N_47635);
xnor U49172 (N_49172,N_47029,N_46188);
and U49173 (N_49173,N_46221,N_46631);
nor U49174 (N_49174,N_47374,N_47109);
nand U49175 (N_49175,N_47427,N_46963);
and U49176 (N_49176,N_47723,N_46914);
and U49177 (N_49177,N_46464,N_47520);
nand U49178 (N_49178,N_46484,N_46439);
nand U49179 (N_49179,N_46469,N_47206);
and U49180 (N_49180,N_46993,N_46652);
nor U49181 (N_49181,N_47781,N_46491);
nor U49182 (N_49182,N_46375,N_46562);
xnor U49183 (N_49183,N_47184,N_47223);
nor U49184 (N_49184,N_47364,N_47170);
nor U49185 (N_49185,N_47086,N_46187);
and U49186 (N_49186,N_47553,N_47487);
and U49187 (N_49187,N_46046,N_47204);
nand U49188 (N_49188,N_46771,N_46177);
nand U49189 (N_49189,N_47351,N_46439);
xnor U49190 (N_49190,N_47021,N_46081);
nand U49191 (N_49191,N_46620,N_47865);
nor U49192 (N_49192,N_46467,N_46619);
or U49193 (N_49193,N_47689,N_47281);
xnor U49194 (N_49194,N_47190,N_47343);
xnor U49195 (N_49195,N_47843,N_47229);
xor U49196 (N_49196,N_47235,N_46053);
xor U49197 (N_49197,N_47613,N_47404);
xor U49198 (N_49198,N_46912,N_46520);
and U49199 (N_49199,N_46058,N_47174);
and U49200 (N_49200,N_46185,N_47675);
or U49201 (N_49201,N_47196,N_46698);
and U49202 (N_49202,N_47307,N_46503);
and U49203 (N_49203,N_47669,N_47611);
and U49204 (N_49204,N_46283,N_46912);
and U49205 (N_49205,N_47215,N_47609);
nand U49206 (N_49206,N_47842,N_46837);
and U49207 (N_49207,N_47697,N_46902);
nand U49208 (N_49208,N_47474,N_46406);
nor U49209 (N_49209,N_47267,N_46987);
or U49210 (N_49210,N_46040,N_46518);
or U49211 (N_49211,N_47084,N_46067);
or U49212 (N_49212,N_47418,N_46930);
nor U49213 (N_49213,N_47557,N_47034);
or U49214 (N_49214,N_47933,N_47553);
and U49215 (N_49215,N_47360,N_46829);
nor U49216 (N_49216,N_47016,N_46635);
nor U49217 (N_49217,N_47068,N_46618);
or U49218 (N_49218,N_46639,N_47498);
nor U49219 (N_49219,N_47565,N_46876);
or U49220 (N_49220,N_46802,N_46493);
or U49221 (N_49221,N_47205,N_46803);
nand U49222 (N_49222,N_47611,N_47591);
nand U49223 (N_49223,N_46076,N_46452);
and U49224 (N_49224,N_46475,N_46265);
nor U49225 (N_49225,N_46330,N_46940);
and U49226 (N_49226,N_46183,N_46802);
nor U49227 (N_49227,N_47712,N_47291);
or U49228 (N_49228,N_46470,N_47349);
and U49229 (N_49229,N_47689,N_47008);
nor U49230 (N_49230,N_46868,N_46842);
and U49231 (N_49231,N_47728,N_47249);
nor U49232 (N_49232,N_47084,N_46484);
nor U49233 (N_49233,N_46960,N_46062);
nor U49234 (N_49234,N_47314,N_47161);
or U49235 (N_49235,N_47086,N_47865);
nor U49236 (N_49236,N_47133,N_46394);
nand U49237 (N_49237,N_46864,N_46370);
nand U49238 (N_49238,N_46505,N_46515);
and U49239 (N_49239,N_47298,N_47682);
or U49240 (N_49240,N_46559,N_46015);
xnor U49241 (N_49241,N_46904,N_46365);
xor U49242 (N_49242,N_47009,N_46639);
or U49243 (N_49243,N_46187,N_47246);
xnor U49244 (N_49244,N_46837,N_47721);
nor U49245 (N_49245,N_47705,N_46856);
and U49246 (N_49246,N_46916,N_46832);
nand U49247 (N_49247,N_47540,N_47786);
and U49248 (N_49248,N_46785,N_46427);
nor U49249 (N_49249,N_47913,N_47235);
nor U49250 (N_49250,N_46117,N_46999);
or U49251 (N_49251,N_46637,N_46548);
xor U49252 (N_49252,N_47827,N_46825);
or U49253 (N_49253,N_46167,N_47685);
or U49254 (N_49254,N_46038,N_46188);
nor U49255 (N_49255,N_47527,N_47386);
or U49256 (N_49256,N_46388,N_47208);
and U49257 (N_49257,N_47264,N_47156);
nand U49258 (N_49258,N_46548,N_46873);
or U49259 (N_49259,N_46290,N_46829);
xor U49260 (N_49260,N_47209,N_47412);
or U49261 (N_49261,N_46762,N_47304);
or U49262 (N_49262,N_47736,N_46854);
nor U49263 (N_49263,N_46102,N_47501);
and U49264 (N_49264,N_47743,N_46635);
or U49265 (N_49265,N_46808,N_47934);
xnor U49266 (N_49266,N_47544,N_46688);
nor U49267 (N_49267,N_47869,N_47761);
nor U49268 (N_49268,N_46480,N_46082);
or U49269 (N_49269,N_47414,N_47969);
or U49270 (N_49270,N_47965,N_47611);
nor U49271 (N_49271,N_46967,N_46723);
and U49272 (N_49272,N_47962,N_46479);
xnor U49273 (N_49273,N_46323,N_47019);
or U49274 (N_49274,N_46688,N_46328);
or U49275 (N_49275,N_47198,N_47701);
nand U49276 (N_49276,N_46791,N_46821);
xnor U49277 (N_49277,N_47704,N_47192);
and U49278 (N_49278,N_47821,N_47665);
and U49279 (N_49279,N_46556,N_46350);
nand U49280 (N_49280,N_47776,N_47240);
or U49281 (N_49281,N_47374,N_46665);
xor U49282 (N_49282,N_46226,N_47994);
or U49283 (N_49283,N_46166,N_46370);
or U49284 (N_49284,N_46484,N_47147);
xor U49285 (N_49285,N_46761,N_46310);
xnor U49286 (N_49286,N_46790,N_47623);
and U49287 (N_49287,N_46289,N_47302);
or U49288 (N_49288,N_47362,N_47241);
or U49289 (N_49289,N_46301,N_47313);
nor U49290 (N_49290,N_46452,N_46763);
and U49291 (N_49291,N_46501,N_47756);
nor U49292 (N_49292,N_46938,N_47341);
and U49293 (N_49293,N_47777,N_46688);
xnor U49294 (N_49294,N_47108,N_47578);
nand U49295 (N_49295,N_47068,N_47733);
or U49296 (N_49296,N_47555,N_47991);
or U49297 (N_49297,N_47753,N_47456);
and U49298 (N_49298,N_47635,N_47456);
nor U49299 (N_49299,N_46683,N_47935);
xor U49300 (N_49300,N_46931,N_46128);
nor U49301 (N_49301,N_46318,N_47401);
and U49302 (N_49302,N_47866,N_47006);
and U49303 (N_49303,N_46336,N_47790);
and U49304 (N_49304,N_47338,N_47762);
or U49305 (N_49305,N_46176,N_47376);
nand U49306 (N_49306,N_47051,N_46502);
and U49307 (N_49307,N_47210,N_46346);
xor U49308 (N_49308,N_46511,N_46241);
xor U49309 (N_49309,N_46448,N_47176);
and U49310 (N_49310,N_46264,N_46959);
xnor U49311 (N_49311,N_46659,N_47756);
or U49312 (N_49312,N_46781,N_47443);
and U49313 (N_49313,N_47327,N_47776);
or U49314 (N_49314,N_46038,N_47248);
xor U49315 (N_49315,N_47993,N_47978);
xor U49316 (N_49316,N_47559,N_47881);
and U49317 (N_49317,N_47102,N_46061);
and U49318 (N_49318,N_47931,N_47638);
xnor U49319 (N_49319,N_47245,N_46306);
xnor U49320 (N_49320,N_46669,N_47970);
and U49321 (N_49321,N_46661,N_46458);
nand U49322 (N_49322,N_47400,N_47510);
or U49323 (N_49323,N_47628,N_46475);
nor U49324 (N_49324,N_46907,N_46280);
nand U49325 (N_49325,N_47854,N_47171);
and U49326 (N_49326,N_46829,N_47908);
and U49327 (N_49327,N_47782,N_46076);
or U49328 (N_49328,N_47666,N_46609);
nand U49329 (N_49329,N_47509,N_47078);
xnor U49330 (N_49330,N_47478,N_47937);
nand U49331 (N_49331,N_47018,N_46796);
and U49332 (N_49332,N_47337,N_47761);
nor U49333 (N_49333,N_46709,N_46573);
xor U49334 (N_49334,N_46086,N_46041);
nor U49335 (N_49335,N_46698,N_46457);
nand U49336 (N_49336,N_46429,N_46546);
and U49337 (N_49337,N_46491,N_47980);
xor U49338 (N_49338,N_47848,N_47282);
and U49339 (N_49339,N_46505,N_47010);
and U49340 (N_49340,N_46111,N_46653);
and U49341 (N_49341,N_47180,N_46242);
and U49342 (N_49342,N_46245,N_47316);
nor U49343 (N_49343,N_46267,N_46318);
nor U49344 (N_49344,N_46484,N_46821);
or U49345 (N_49345,N_46100,N_47632);
nand U49346 (N_49346,N_47165,N_46789);
and U49347 (N_49347,N_46117,N_47054);
nand U49348 (N_49348,N_46474,N_47527);
xor U49349 (N_49349,N_46416,N_46883);
xnor U49350 (N_49350,N_46823,N_47821);
nand U49351 (N_49351,N_47872,N_46884);
or U49352 (N_49352,N_46501,N_47359);
and U49353 (N_49353,N_46307,N_46972);
nor U49354 (N_49354,N_47464,N_47124);
nor U49355 (N_49355,N_46479,N_47756);
nor U49356 (N_49356,N_47681,N_46723);
xnor U49357 (N_49357,N_46951,N_46140);
nand U49358 (N_49358,N_47375,N_46401);
nor U49359 (N_49359,N_47746,N_46303);
or U49360 (N_49360,N_47480,N_47430);
and U49361 (N_49361,N_47446,N_46460);
xnor U49362 (N_49362,N_47752,N_46995);
or U49363 (N_49363,N_46974,N_46906);
or U49364 (N_49364,N_46779,N_46987);
nand U49365 (N_49365,N_47654,N_46333);
or U49366 (N_49366,N_46050,N_46180);
or U49367 (N_49367,N_46806,N_47194);
or U49368 (N_49368,N_46330,N_47397);
xor U49369 (N_49369,N_47650,N_46846);
or U49370 (N_49370,N_47979,N_46866);
and U49371 (N_49371,N_46485,N_47668);
or U49372 (N_49372,N_47492,N_46213);
nor U49373 (N_49373,N_47266,N_47591);
or U49374 (N_49374,N_46878,N_46555);
xor U49375 (N_49375,N_46043,N_47488);
and U49376 (N_49376,N_47220,N_47527);
xor U49377 (N_49377,N_46449,N_46822);
or U49378 (N_49378,N_47991,N_47112);
and U49379 (N_49379,N_47133,N_46146);
nand U49380 (N_49380,N_46838,N_46202);
and U49381 (N_49381,N_46522,N_47725);
nand U49382 (N_49382,N_47005,N_47826);
xor U49383 (N_49383,N_47284,N_46614);
or U49384 (N_49384,N_46771,N_46758);
and U49385 (N_49385,N_46584,N_46921);
nand U49386 (N_49386,N_46813,N_47537);
or U49387 (N_49387,N_47493,N_47229);
nor U49388 (N_49388,N_47000,N_47577);
xnor U49389 (N_49389,N_47148,N_47009);
xnor U49390 (N_49390,N_46767,N_46947);
or U49391 (N_49391,N_47935,N_47709);
and U49392 (N_49392,N_47586,N_47699);
nor U49393 (N_49393,N_47540,N_46673);
nor U49394 (N_49394,N_46933,N_47397);
xnor U49395 (N_49395,N_46598,N_47753);
and U49396 (N_49396,N_46078,N_46891);
or U49397 (N_49397,N_47824,N_47819);
xnor U49398 (N_49398,N_47708,N_47146);
nor U49399 (N_49399,N_46915,N_47070);
or U49400 (N_49400,N_46515,N_47085);
nor U49401 (N_49401,N_46711,N_46405);
and U49402 (N_49402,N_46195,N_47560);
nor U49403 (N_49403,N_46815,N_46027);
xnor U49404 (N_49404,N_47508,N_46880);
or U49405 (N_49405,N_47647,N_47325);
nor U49406 (N_49406,N_47794,N_47732);
nor U49407 (N_49407,N_46451,N_46567);
and U49408 (N_49408,N_47290,N_47223);
nor U49409 (N_49409,N_46929,N_47032);
nor U49410 (N_49410,N_46198,N_47985);
xor U49411 (N_49411,N_47898,N_47439);
or U49412 (N_49412,N_46645,N_46166);
nand U49413 (N_49413,N_46391,N_46635);
or U49414 (N_49414,N_46457,N_46147);
nand U49415 (N_49415,N_46928,N_46439);
nor U49416 (N_49416,N_47622,N_47310);
nand U49417 (N_49417,N_46015,N_46637);
and U49418 (N_49418,N_46073,N_47452);
nor U49419 (N_49419,N_47440,N_47457);
or U49420 (N_49420,N_46226,N_47525);
or U49421 (N_49421,N_47764,N_47319);
nand U49422 (N_49422,N_47819,N_46488);
nor U49423 (N_49423,N_47533,N_46601);
or U49424 (N_49424,N_47956,N_47265);
nand U49425 (N_49425,N_47066,N_47742);
xor U49426 (N_49426,N_46442,N_46059);
or U49427 (N_49427,N_46535,N_46324);
xnor U49428 (N_49428,N_47146,N_47650);
or U49429 (N_49429,N_47587,N_46415);
and U49430 (N_49430,N_47277,N_47290);
nand U49431 (N_49431,N_47285,N_47676);
nor U49432 (N_49432,N_46521,N_46876);
nor U49433 (N_49433,N_47736,N_46608);
nand U49434 (N_49434,N_47734,N_47283);
nand U49435 (N_49435,N_47197,N_46560);
or U49436 (N_49436,N_46204,N_47632);
and U49437 (N_49437,N_46159,N_46351);
nand U49438 (N_49438,N_47343,N_47242);
xnor U49439 (N_49439,N_46857,N_46063);
or U49440 (N_49440,N_47837,N_47710);
nor U49441 (N_49441,N_47683,N_47800);
and U49442 (N_49442,N_47104,N_46501);
xnor U49443 (N_49443,N_47065,N_46467);
nor U49444 (N_49444,N_46783,N_47940);
nand U49445 (N_49445,N_46467,N_46400);
and U49446 (N_49446,N_46640,N_46198);
nand U49447 (N_49447,N_46145,N_47243);
or U49448 (N_49448,N_47029,N_46841);
xnor U49449 (N_49449,N_46572,N_46019);
nor U49450 (N_49450,N_46374,N_47451);
nor U49451 (N_49451,N_46163,N_46878);
nand U49452 (N_49452,N_46472,N_47969);
and U49453 (N_49453,N_46475,N_46733);
nand U49454 (N_49454,N_46730,N_47309);
xor U49455 (N_49455,N_46087,N_46485);
and U49456 (N_49456,N_46407,N_46251);
xnor U49457 (N_49457,N_46247,N_46344);
or U49458 (N_49458,N_47410,N_47129);
nor U49459 (N_49459,N_46305,N_47900);
xnor U49460 (N_49460,N_46762,N_47521);
nand U49461 (N_49461,N_46665,N_47368);
and U49462 (N_49462,N_47948,N_46162);
nor U49463 (N_49463,N_47956,N_47075);
and U49464 (N_49464,N_47790,N_46727);
xor U49465 (N_49465,N_47974,N_47180);
nor U49466 (N_49466,N_46102,N_46250);
nand U49467 (N_49467,N_46491,N_46313);
nand U49468 (N_49468,N_46565,N_46653);
and U49469 (N_49469,N_46493,N_46422);
xnor U49470 (N_49470,N_46871,N_47097);
nand U49471 (N_49471,N_46961,N_46727);
and U49472 (N_49472,N_46491,N_46074);
xor U49473 (N_49473,N_46627,N_46962);
and U49474 (N_49474,N_47624,N_46898);
nor U49475 (N_49475,N_47479,N_46547);
nor U49476 (N_49476,N_47235,N_47664);
and U49477 (N_49477,N_47671,N_46278);
or U49478 (N_49478,N_47979,N_46060);
and U49479 (N_49479,N_46864,N_47755);
nor U49480 (N_49480,N_47454,N_46327);
and U49481 (N_49481,N_47471,N_46231);
and U49482 (N_49482,N_46503,N_46570);
and U49483 (N_49483,N_47947,N_46614);
and U49484 (N_49484,N_46875,N_46085);
nand U49485 (N_49485,N_47014,N_46394);
or U49486 (N_49486,N_46419,N_47106);
nand U49487 (N_49487,N_46108,N_47261);
xnor U49488 (N_49488,N_47910,N_47668);
and U49489 (N_49489,N_46921,N_47880);
and U49490 (N_49490,N_46194,N_47015);
nor U49491 (N_49491,N_46389,N_46831);
xnor U49492 (N_49492,N_47693,N_46951);
nand U49493 (N_49493,N_46424,N_46959);
or U49494 (N_49494,N_46017,N_47834);
xnor U49495 (N_49495,N_47084,N_47454);
nor U49496 (N_49496,N_47335,N_46884);
or U49497 (N_49497,N_47397,N_47361);
nand U49498 (N_49498,N_46603,N_46344);
xnor U49499 (N_49499,N_46465,N_47042);
nor U49500 (N_49500,N_47884,N_46040);
xnor U49501 (N_49501,N_46235,N_47669);
xnor U49502 (N_49502,N_46917,N_47381);
xor U49503 (N_49503,N_47573,N_47571);
nand U49504 (N_49504,N_46942,N_47572);
or U49505 (N_49505,N_47512,N_47845);
nor U49506 (N_49506,N_47509,N_46085);
nand U49507 (N_49507,N_47859,N_46162);
or U49508 (N_49508,N_47561,N_46777);
xnor U49509 (N_49509,N_47777,N_46931);
or U49510 (N_49510,N_47602,N_46929);
nor U49511 (N_49511,N_46039,N_46821);
xor U49512 (N_49512,N_46386,N_46112);
xnor U49513 (N_49513,N_47012,N_47638);
nor U49514 (N_49514,N_46504,N_46450);
or U49515 (N_49515,N_46115,N_46484);
and U49516 (N_49516,N_46267,N_46687);
nor U49517 (N_49517,N_47100,N_47959);
nand U49518 (N_49518,N_47073,N_46912);
and U49519 (N_49519,N_47500,N_47704);
nor U49520 (N_49520,N_47965,N_47399);
nand U49521 (N_49521,N_46254,N_47630);
nor U49522 (N_49522,N_46318,N_46365);
nor U49523 (N_49523,N_46817,N_46208);
and U49524 (N_49524,N_46237,N_47519);
nor U49525 (N_49525,N_46236,N_47567);
xnor U49526 (N_49526,N_46247,N_47873);
nor U49527 (N_49527,N_46872,N_46418);
or U49528 (N_49528,N_47923,N_46855);
nor U49529 (N_49529,N_47834,N_47332);
and U49530 (N_49530,N_46915,N_46561);
or U49531 (N_49531,N_46911,N_47908);
nor U49532 (N_49532,N_47001,N_47989);
nor U49533 (N_49533,N_46358,N_47719);
nand U49534 (N_49534,N_46363,N_47778);
or U49535 (N_49535,N_46811,N_47737);
or U49536 (N_49536,N_46481,N_47664);
and U49537 (N_49537,N_47549,N_47941);
xnor U49538 (N_49538,N_46674,N_46894);
nand U49539 (N_49539,N_47516,N_47828);
xor U49540 (N_49540,N_46849,N_46404);
xnor U49541 (N_49541,N_46732,N_46940);
and U49542 (N_49542,N_46404,N_46827);
nand U49543 (N_49543,N_47685,N_46709);
nor U49544 (N_49544,N_46456,N_46202);
and U49545 (N_49545,N_46282,N_46512);
nand U49546 (N_49546,N_47140,N_46005);
and U49547 (N_49547,N_46882,N_46015);
xnor U49548 (N_49548,N_46914,N_47416);
and U49549 (N_49549,N_46302,N_46446);
or U49550 (N_49550,N_47645,N_47779);
or U49551 (N_49551,N_47346,N_46854);
and U49552 (N_49552,N_47550,N_46362);
nor U49553 (N_49553,N_46990,N_46268);
nor U49554 (N_49554,N_47416,N_46814);
or U49555 (N_49555,N_46825,N_47656);
xnor U49556 (N_49556,N_47933,N_47475);
and U49557 (N_49557,N_46152,N_46400);
nand U49558 (N_49558,N_47451,N_46112);
or U49559 (N_49559,N_46793,N_46545);
or U49560 (N_49560,N_47456,N_47305);
or U49561 (N_49561,N_47042,N_46077);
nor U49562 (N_49562,N_47917,N_47754);
nor U49563 (N_49563,N_46459,N_46796);
or U49564 (N_49564,N_47434,N_46139);
xnor U49565 (N_49565,N_46337,N_46774);
nor U49566 (N_49566,N_46200,N_47837);
nor U49567 (N_49567,N_46732,N_47005);
and U49568 (N_49568,N_46045,N_46756);
or U49569 (N_49569,N_47271,N_46873);
or U49570 (N_49570,N_46857,N_47076);
or U49571 (N_49571,N_46189,N_46520);
or U49572 (N_49572,N_47186,N_47548);
and U49573 (N_49573,N_47984,N_47381);
xnor U49574 (N_49574,N_46213,N_46893);
nand U49575 (N_49575,N_46920,N_47228);
and U49576 (N_49576,N_47697,N_46849);
nor U49577 (N_49577,N_47831,N_47348);
and U49578 (N_49578,N_47843,N_46978);
and U49579 (N_49579,N_46828,N_47271);
nor U49580 (N_49580,N_46386,N_47725);
and U49581 (N_49581,N_46771,N_47711);
and U49582 (N_49582,N_46125,N_47073);
xor U49583 (N_49583,N_46431,N_47877);
nor U49584 (N_49584,N_46869,N_47924);
nor U49585 (N_49585,N_47781,N_46403);
nand U49586 (N_49586,N_46688,N_47379);
or U49587 (N_49587,N_47464,N_46446);
nand U49588 (N_49588,N_46852,N_47495);
or U49589 (N_49589,N_46940,N_47787);
or U49590 (N_49590,N_46498,N_46736);
xnor U49591 (N_49591,N_46332,N_47457);
xor U49592 (N_49592,N_46988,N_46417);
xnor U49593 (N_49593,N_47780,N_47058);
or U49594 (N_49594,N_47265,N_46911);
or U49595 (N_49595,N_46240,N_46521);
and U49596 (N_49596,N_47906,N_47501);
nor U49597 (N_49597,N_46274,N_46424);
or U49598 (N_49598,N_46502,N_46356);
nor U49599 (N_49599,N_47485,N_46406);
or U49600 (N_49600,N_46583,N_47144);
nor U49601 (N_49601,N_46118,N_47327);
or U49602 (N_49602,N_46572,N_47645);
xor U49603 (N_49603,N_47666,N_46250);
nand U49604 (N_49604,N_46711,N_47315);
nand U49605 (N_49605,N_47684,N_47094);
xnor U49606 (N_49606,N_46820,N_46146);
or U49607 (N_49607,N_46568,N_47186);
xor U49608 (N_49608,N_47900,N_46112);
and U49609 (N_49609,N_47390,N_47843);
and U49610 (N_49610,N_47005,N_47986);
or U49611 (N_49611,N_46964,N_47403);
nor U49612 (N_49612,N_47712,N_47552);
nor U49613 (N_49613,N_47466,N_46920);
or U49614 (N_49614,N_47085,N_47712);
and U49615 (N_49615,N_46744,N_47164);
nor U49616 (N_49616,N_47161,N_46695);
xor U49617 (N_49617,N_46826,N_46156);
xnor U49618 (N_49618,N_46821,N_46947);
and U49619 (N_49619,N_47443,N_47909);
nor U49620 (N_49620,N_46825,N_47567);
or U49621 (N_49621,N_47131,N_47390);
nand U49622 (N_49622,N_46225,N_46501);
or U49623 (N_49623,N_47624,N_46984);
xor U49624 (N_49624,N_46797,N_46963);
nand U49625 (N_49625,N_46000,N_47816);
nor U49626 (N_49626,N_46931,N_47138);
nand U49627 (N_49627,N_46079,N_47791);
nand U49628 (N_49628,N_46519,N_47452);
and U49629 (N_49629,N_46050,N_46859);
nand U49630 (N_49630,N_46647,N_47482);
nand U49631 (N_49631,N_46370,N_47384);
xnor U49632 (N_49632,N_47949,N_47335);
nor U49633 (N_49633,N_46322,N_47698);
or U49634 (N_49634,N_46856,N_46773);
xor U49635 (N_49635,N_46963,N_46695);
or U49636 (N_49636,N_46902,N_46709);
or U49637 (N_49637,N_47534,N_46378);
nand U49638 (N_49638,N_46297,N_47435);
and U49639 (N_49639,N_47154,N_47833);
xnor U49640 (N_49640,N_47331,N_46929);
nor U49641 (N_49641,N_47989,N_46669);
nand U49642 (N_49642,N_46398,N_46915);
nand U49643 (N_49643,N_46436,N_47808);
nand U49644 (N_49644,N_47166,N_47622);
nor U49645 (N_49645,N_46848,N_46119);
or U49646 (N_49646,N_46256,N_47467);
nor U49647 (N_49647,N_46382,N_46633);
xnor U49648 (N_49648,N_47145,N_47380);
nor U49649 (N_49649,N_46640,N_47082);
nor U49650 (N_49650,N_47159,N_47024);
nand U49651 (N_49651,N_47581,N_47120);
nor U49652 (N_49652,N_46818,N_47757);
xor U49653 (N_49653,N_47809,N_47212);
and U49654 (N_49654,N_46067,N_47763);
nand U49655 (N_49655,N_46827,N_47315);
xor U49656 (N_49656,N_46113,N_46062);
xor U49657 (N_49657,N_46127,N_47933);
xnor U49658 (N_49658,N_46071,N_47973);
nand U49659 (N_49659,N_46817,N_47621);
nor U49660 (N_49660,N_46790,N_47881);
nand U49661 (N_49661,N_46744,N_46314);
or U49662 (N_49662,N_47576,N_46298);
or U49663 (N_49663,N_47301,N_47165);
and U49664 (N_49664,N_47915,N_47288);
xor U49665 (N_49665,N_46740,N_46471);
nor U49666 (N_49666,N_47256,N_47671);
nand U49667 (N_49667,N_47827,N_47659);
nor U49668 (N_49668,N_47288,N_46306);
and U49669 (N_49669,N_47812,N_47758);
nand U49670 (N_49670,N_47249,N_46789);
xor U49671 (N_49671,N_47359,N_46188);
nor U49672 (N_49672,N_47233,N_47451);
xor U49673 (N_49673,N_47638,N_46625);
nand U49674 (N_49674,N_47617,N_46093);
xor U49675 (N_49675,N_47796,N_47538);
nand U49676 (N_49676,N_47376,N_46050);
xor U49677 (N_49677,N_47308,N_47692);
or U49678 (N_49678,N_46419,N_47660);
nor U49679 (N_49679,N_47711,N_47296);
nor U49680 (N_49680,N_46405,N_46862);
or U49681 (N_49681,N_46059,N_47520);
and U49682 (N_49682,N_47656,N_47813);
xor U49683 (N_49683,N_47641,N_46483);
and U49684 (N_49684,N_47671,N_47762);
nand U49685 (N_49685,N_47111,N_46457);
nand U49686 (N_49686,N_46812,N_47962);
or U49687 (N_49687,N_46023,N_46021);
xnor U49688 (N_49688,N_46184,N_46008);
nand U49689 (N_49689,N_46453,N_47260);
xor U49690 (N_49690,N_46870,N_47078);
nor U49691 (N_49691,N_47934,N_47741);
or U49692 (N_49692,N_47209,N_46184);
nor U49693 (N_49693,N_46086,N_47580);
and U49694 (N_49694,N_46910,N_47592);
xor U49695 (N_49695,N_47060,N_47468);
and U49696 (N_49696,N_46216,N_46550);
nor U49697 (N_49697,N_47681,N_46271);
nand U49698 (N_49698,N_46421,N_46527);
xnor U49699 (N_49699,N_47188,N_47019);
xnor U49700 (N_49700,N_46341,N_46375);
nand U49701 (N_49701,N_46324,N_47058);
or U49702 (N_49702,N_46885,N_47191);
xor U49703 (N_49703,N_47934,N_47170);
nor U49704 (N_49704,N_47347,N_46590);
nand U49705 (N_49705,N_46439,N_47911);
or U49706 (N_49706,N_46655,N_46259);
and U49707 (N_49707,N_47496,N_47284);
and U49708 (N_49708,N_47990,N_47847);
and U49709 (N_49709,N_46840,N_47874);
and U49710 (N_49710,N_46883,N_47393);
nor U49711 (N_49711,N_47643,N_47151);
nand U49712 (N_49712,N_46088,N_47783);
or U49713 (N_49713,N_46909,N_47906);
xor U49714 (N_49714,N_46927,N_47268);
and U49715 (N_49715,N_47077,N_46766);
and U49716 (N_49716,N_47676,N_47567);
nand U49717 (N_49717,N_46548,N_46292);
and U49718 (N_49718,N_47991,N_46179);
and U49719 (N_49719,N_47798,N_47285);
xor U49720 (N_49720,N_46011,N_47886);
and U49721 (N_49721,N_46525,N_46059);
or U49722 (N_49722,N_46767,N_46027);
nand U49723 (N_49723,N_46916,N_47731);
xor U49724 (N_49724,N_46192,N_47516);
nor U49725 (N_49725,N_46512,N_46926);
xnor U49726 (N_49726,N_47517,N_47097);
xnor U49727 (N_49727,N_47780,N_47672);
or U49728 (N_49728,N_46576,N_47608);
nor U49729 (N_49729,N_46439,N_47680);
nand U49730 (N_49730,N_46573,N_46863);
xnor U49731 (N_49731,N_46996,N_47681);
nor U49732 (N_49732,N_46624,N_46143);
nand U49733 (N_49733,N_47809,N_46506);
and U49734 (N_49734,N_46649,N_47406);
nand U49735 (N_49735,N_46726,N_46873);
or U49736 (N_49736,N_47774,N_47777);
and U49737 (N_49737,N_47936,N_47913);
and U49738 (N_49738,N_46829,N_46421);
or U49739 (N_49739,N_46530,N_47110);
and U49740 (N_49740,N_47405,N_46254);
xor U49741 (N_49741,N_47846,N_46752);
or U49742 (N_49742,N_46558,N_47168);
nand U49743 (N_49743,N_47354,N_47473);
xor U49744 (N_49744,N_46296,N_47413);
nor U49745 (N_49745,N_46365,N_46884);
nor U49746 (N_49746,N_46861,N_47664);
or U49747 (N_49747,N_47351,N_46061);
nor U49748 (N_49748,N_47007,N_47990);
and U49749 (N_49749,N_46560,N_47572);
nor U49750 (N_49750,N_46026,N_47434);
nor U49751 (N_49751,N_46887,N_46205);
nand U49752 (N_49752,N_47506,N_46791);
nor U49753 (N_49753,N_47276,N_46418);
nor U49754 (N_49754,N_46235,N_46529);
nor U49755 (N_49755,N_46092,N_46391);
and U49756 (N_49756,N_46331,N_46133);
and U49757 (N_49757,N_46871,N_47358);
nor U49758 (N_49758,N_47800,N_46184);
and U49759 (N_49759,N_47857,N_47450);
nand U49760 (N_49760,N_47387,N_47962);
or U49761 (N_49761,N_46934,N_47557);
xor U49762 (N_49762,N_46362,N_47064);
nand U49763 (N_49763,N_46596,N_47769);
xor U49764 (N_49764,N_47031,N_47966);
xnor U49765 (N_49765,N_47710,N_47841);
and U49766 (N_49766,N_47129,N_47151);
nand U49767 (N_49767,N_46428,N_46968);
nor U49768 (N_49768,N_47118,N_47180);
nor U49769 (N_49769,N_46821,N_46734);
nand U49770 (N_49770,N_46883,N_47893);
and U49771 (N_49771,N_47578,N_46714);
xor U49772 (N_49772,N_47224,N_46980);
nor U49773 (N_49773,N_46434,N_46867);
xor U49774 (N_49774,N_46720,N_47292);
or U49775 (N_49775,N_47876,N_47188);
nor U49776 (N_49776,N_47901,N_46306);
or U49777 (N_49777,N_46216,N_47761);
nand U49778 (N_49778,N_46385,N_47111);
xnor U49779 (N_49779,N_46302,N_47457);
nor U49780 (N_49780,N_46041,N_46234);
nand U49781 (N_49781,N_47331,N_46631);
nor U49782 (N_49782,N_46051,N_46103);
and U49783 (N_49783,N_47933,N_46596);
nand U49784 (N_49784,N_46786,N_47427);
xnor U49785 (N_49785,N_47122,N_46287);
xnor U49786 (N_49786,N_47082,N_46106);
and U49787 (N_49787,N_46823,N_46159);
and U49788 (N_49788,N_47144,N_47432);
nor U49789 (N_49789,N_47560,N_46147);
xor U49790 (N_49790,N_47815,N_47934);
nand U49791 (N_49791,N_46628,N_46675);
xnor U49792 (N_49792,N_46554,N_47608);
and U49793 (N_49793,N_47032,N_46478);
nor U49794 (N_49794,N_47208,N_46902);
and U49795 (N_49795,N_47537,N_46560);
nand U49796 (N_49796,N_46307,N_47930);
nand U49797 (N_49797,N_46337,N_46671);
and U49798 (N_49798,N_47019,N_46636);
or U49799 (N_49799,N_47806,N_46116);
nor U49800 (N_49800,N_46363,N_47375);
nand U49801 (N_49801,N_46660,N_46606);
nand U49802 (N_49802,N_46781,N_47927);
xnor U49803 (N_49803,N_46173,N_46217);
nand U49804 (N_49804,N_46448,N_46905);
nor U49805 (N_49805,N_46295,N_47584);
nor U49806 (N_49806,N_46444,N_47323);
xnor U49807 (N_49807,N_47233,N_46898);
nor U49808 (N_49808,N_47065,N_47859);
nor U49809 (N_49809,N_46742,N_47669);
nor U49810 (N_49810,N_46627,N_46206);
and U49811 (N_49811,N_47238,N_47061);
nor U49812 (N_49812,N_47417,N_47580);
and U49813 (N_49813,N_47181,N_46406);
or U49814 (N_49814,N_47628,N_47831);
and U49815 (N_49815,N_47066,N_47551);
or U49816 (N_49816,N_47053,N_47374);
nand U49817 (N_49817,N_47404,N_46060);
xnor U49818 (N_49818,N_47501,N_47296);
or U49819 (N_49819,N_47721,N_46253);
nor U49820 (N_49820,N_47465,N_46522);
nor U49821 (N_49821,N_46586,N_47545);
nand U49822 (N_49822,N_46765,N_47561);
and U49823 (N_49823,N_46377,N_46878);
nand U49824 (N_49824,N_47767,N_46037);
xnor U49825 (N_49825,N_47206,N_46565);
nand U49826 (N_49826,N_46856,N_46001);
nand U49827 (N_49827,N_46893,N_47993);
or U49828 (N_49828,N_46992,N_47706);
nor U49829 (N_49829,N_46227,N_47435);
nand U49830 (N_49830,N_47303,N_47564);
xor U49831 (N_49831,N_47076,N_46891);
xor U49832 (N_49832,N_47097,N_46045);
xnor U49833 (N_49833,N_47644,N_47422);
and U49834 (N_49834,N_46994,N_47958);
and U49835 (N_49835,N_47092,N_46776);
xnor U49836 (N_49836,N_47809,N_46056);
nor U49837 (N_49837,N_46510,N_46445);
and U49838 (N_49838,N_47769,N_47002);
nand U49839 (N_49839,N_46830,N_46376);
and U49840 (N_49840,N_46787,N_46856);
nor U49841 (N_49841,N_46500,N_47095);
nor U49842 (N_49842,N_47668,N_47789);
or U49843 (N_49843,N_47291,N_47955);
and U49844 (N_49844,N_46851,N_47709);
and U49845 (N_49845,N_47407,N_47201);
nand U49846 (N_49846,N_46773,N_47683);
and U49847 (N_49847,N_47308,N_46513);
or U49848 (N_49848,N_47265,N_46675);
and U49849 (N_49849,N_47405,N_46097);
nor U49850 (N_49850,N_46059,N_46698);
nor U49851 (N_49851,N_46381,N_46774);
and U49852 (N_49852,N_46404,N_47192);
or U49853 (N_49853,N_46955,N_46736);
nand U49854 (N_49854,N_47689,N_46357);
nand U49855 (N_49855,N_47202,N_47551);
nand U49856 (N_49856,N_46759,N_47688);
or U49857 (N_49857,N_47638,N_47884);
nand U49858 (N_49858,N_46005,N_46067);
nor U49859 (N_49859,N_46757,N_46753);
nor U49860 (N_49860,N_47249,N_47800);
and U49861 (N_49861,N_46417,N_46632);
nand U49862 (N_49862,N_47862,N_46105);
and U49863 (N_49863,N_47449,N_47792);
nor U49864 (N_49864,N_46249,N_46540);
nand U49865 (N_49865,N_46281,N_47641);
and U49866 (N_49866,N_47856,N_47640);
nor U49867 (N_49867,N_46518,N_47659);
nand U49868 (N_49868,N_46035,N_47990);
xor U49869 (N_49869,N_47994,N_46048);
xor U49870 (N_49870,N_47272,N_47837);
nand U49871 (N_49871,N_46690,N_46719);
nor U49872 (N_49872,N_46211,N_46831);
nand U49873 (N_49873,N_47918,N_47985);
xnor U49874 (N_49874,N_47528,N_46579);
xor U49875 (N_49875,N_47503,N_46758);
or U49876 (N_49876,N_47656,N_47881);
nor U49877 (N_49877,N_46996,N_46660);
and U49878 (N_49878,N_46605,N_46543);
nor U49879 (N_49879,N_47369,N_47131);
nor U49880 (N_49880,N_47543,N_47693);
xor U49881 (N_49881,N_47762,N_47324);
nand U49882 (N_49882,N_46498,N_47195);
nand U49883 (N_49883,N_47048,N_46523);
nor U49884 (N_49884,N_46239,N_47398);
xor U49885 (N_49885,N_47085,N_46202);
nor U49886 (N_49886,N_46667,N_47339);
or U49887 (N_49887,N_47602,N_46610);
nand U49888 (N_49888,N_47637,N_46452);
nor U49889 (N_49889,N_47366,N_47736);
nor U49890 (N_49890,N_46339,N_46282);
nor U49891 (N_49891,N_47381,N_46857);
xor U49892 (N_49892,N_46028,N_47590);
or U49893 (N_49893,N_47273,N_46715);
nor U49894 (N_49894,N_46427,N_47476);
nand U49895 (N_49895,N_46305,N_47043);
or U49896 (N_49896,N_47731,N_46905);
and U49897 (N_49897,N_47200,N_46797);
nor U49898 (N_49898,N_46505,N_46280);
nand U49899 (N_49899,N_46669,N_46475);
or U49900 (N_49900,N_46353,N_46379);
or U49901 (N_49901,N_46541,N_47127);
nor U49902 (N_49902,N_46717,N_47342);
nand U49903 (N_49903,N_46416,N_46381);
nor U49904 (N_49904,N_47127,N_47444);
or U49905 (N_49905,N_46201,N_46424);
xor U49906 (N_49906,N_47085,N_47313);
and U49907 (N_49907,N_46110,N_47560);
or U49908 (N_49908,N_47757,N_46747);
nand U49909 (N_49909,N_47630,N_47515);
xnor U49910 (N_49910,N_47667,N_47063);
xnor U49911 (N_49911,N_47433,N_47401);
and U49912 (N_49912,N_47673,N_46618);
or U49913 (N_49913,N_47405,N_46577);
nand U49914 (N_49914,N_47149,N_46947);
nand U49915 (N_49915,N_47230,N_47344);
xor U49916 (N_49916,N_46108,N_47809);
xor U49917 (N_49917,N_46987,N_46998);
nand U49918 (N_49918,N_47795,N_47947);
nand U49919 (N_49919,N_46019,N_47163);
nand U49920 (N_49920,N_46735,N_47325);
xor U49921 (N_49921,N_47856,N_47209);
or U49922 (N_49922,N_46639,N_47897);
and U49923 (N_49923,N_47702,N_47092);
nand U49924 (N_49924,N_47876,N_46866);
nand U49925 (N_49925,N_47972,N_47940);
xnor U49926 (N_49926,N_47855,N_47036);
nand U49927 (N_49927,N_46578,N_46346);
or U49928 (N_49928,N_47621,N_46122);
and U49929 (N_49929,N_47921,N_47448);
nand U49930 (N_49930,N_47687,N_46990);
or U49931 (N_49931,N_47622,N_46311);
nor U49932 (N_49932,N_47626,N_46398);
nand U49933 (N_49933,N_46270,N_47871);
nor U49934 (N_49934,N_47951,N_46635);
or U49935 (N_49935,N_46645,N_47544);
nand U49936 (N_49936,N_47751,N_46216);
nor U49937 (N_49937,N_46823,N_46184);
xor U49938 (N_49938,N_46370,N_46735);
and U49939 (N_49939,N_47280,N_46058);
nor U49940 (N_49940,N_46589,N_47033);
xor U49941 (N_49941,N_47037,N_46920);
and U49942 (N_49942,N_46573,N_46051);
or U49943 (N_49943,N_47770,N_47373);
and U49944 (N_49944,N_47961,N_47173);
nor U49945 (N_49945,N_46483,N_46567);
and U49946 (N_49946,N_46516,N_46518);
or U49947 (N_49947,N_47774,N_46732);
xor U49948 (N_49948,N_46219,N_46358);
nand U49949 (N_49949,N_47248,N_47986);
or U49950 (N_49950,N_47959,N_47026);
nand U49951 (N_49951,N_46316,N_46341);
and U49952 (N_49952,N_46403,N_47569);
xnor U49953 (N_49953,N_47704,N_47839);
nor U49954 (N_49954,N_47526,N_46409);
nor U49955 (N_49955,N_46944,N_47449);
and U49956 (N_49956,N_46167,N_47500);
or U49957 (N_49957,N_46094,N_46604);
nand U49958 (N_49958,N_47524,N_47560);
or U49959 (N_49959,N_46948,N_47012);
or U49960 (N_49960,N_47277,N_46059);
nand U49961 (N_49961,N_46388,N_46104);
xnor U49962 (N_49962,N_46591,N_46132);
or U49963 (N_49963,N_47973,N_47098);
xor U49964 (N_49964,N_46482,N_46551);
or U49965 (N_49965,N_46300,N_47930);
and U49966 (N_49966,N_47601,N_47382);
or U49967 (N_49967,N_47261,N_46495);
nor U49968 (N_49968,N_46876,N_46134);
nand U49969 (N_49969,N_47613,N_47243);
nor U49970 (N_49970,N_46137,N_46204);
or U49971 (N_49971,N_46736,N_47738);
nand U49972 (N_49972,N_47807,N_47440);
nor U49973 (N_49973,N_46642,N_47280);
nor U49974 (N_49974,N_46966,N_47486);
or U49975 (N_49975,N_47675,N_47493);
xor U49976 (N_49976,N_47833,N_47899);
nor U49977 (N_49977,N_46465,N_46707);
and U49978 (N_49978,N_46955,N_47608);
or U49979 (N_49979,N_46301,N_47743);
xor U49980 (N_49980,N_47124,N_46919);
and U49981 (N_49981,N_47628,N_47699);
nor U49982 (N_49982,N_47535,N_47508);
or U49983 (N_49983,N_46221,N_47214);
nor U49984 (N_49984,N_46719,N_47211);
xnor U49985 (N_49985,N_47793,N_47528);
xnor U49986 (N_49986,N_46798,N_46128);
nor U49987 (N_49987,N_47111,N_46152);
xnor U49988 (N_49988,N_46672,N_47094);
or U49989 (N_49989,N_46614,N_46852);
nand U49990 (N_49990,N_47508,N_46799);
nor U49991 (N_49991,N_47080,N_47156);
nand U49992 (N_49992,N_46840,N_47921);
or U49993 (N_49993,N_46806,N_46136);
and U49994 (N_49994,N_46036,N_46013);
or U49995 (N_49995,N_46621,N_47369);
xnor U49996 (N_49996,N_46302,N_47578);
nor U49997 (N_49997,N_46501,N_46604);
xnor U49998 (N_49998,N_46483,N_46078);
xnor U49999 (N_49999,N_46017,N_46726);
nor UO_0 (O_0,N_48977,N_48821);
xor UO_1 (O_1,N_49441,N_48965);
or UO_2 (O_2,N_48953,N_48131);
or UO_3 (O_3,N_48041,N_49796);
nor UO_4 (O_4,N_48088,N_49229);
nor UO_5 (O_5,N_48955,N_48391);
xor UO_6 (O_6,N_49766,N_49198);
xor UO_7 (O_7,N_49697,N_49500);
or UO_8 (O_8,N_49779,N_48360);
nor UO_9 (O_9,N_48229,N_48364);
xnor UO_10 (O_10,N_49768,N_48467);
and UO_11 (O_11,N_49345,N_49675);
xnor UO_12 (O_12,N_49221,N_48021);
xnor UO_13 (O_13,N_48835,N_49888);
or UO_14 (O_14,N_49076,N_49893);
xor UO_15 (O_15,N_48944,N_49609);
and UO_16 (O_16,N_49900,N_48848);
nor UO_17 (O_17,N_49445,N_48428);
and UO_18 (O_18,N_49048,N_48401);
and UO_19 (O_19,N_48878,N_49561);
nor UO_20 (O_20,N_48404,N_48441);
or UO_21 (O_21,N_48692,N_49167);
xor UO_22 (O_22,N_48800,N_48031);
nor UO_23 (O_23,N_49702,N_49460);
or UO_24 (O_24,N_48228,N_48054);
or UO_25 (O_25,N_49898,N_49645);
and UO_26 (O_26,N_49897,N_48497);
or UO_27 (O_27,N_49138,N_49406);
nand UO_28 (O_28,N_49479,N_48556);
or UO_29 (O_29,N_49189,N_48175);
nor UO_30 (O_30,N_48411,N_49588);
or UO_31 (O_31,N_49781,N_49709);
xnor UO_32 (O_32,N_48709,N_48924);
xor UO_33 (O_33,N_48792,N_49089);
nor UO_34 (O_34,N_49165,N_49295);
xor UO_35 (O_35,N_48765,N_49948);
nor UO_36 (O_36,N_49589,N_48998);
nand UO_37 (O_37,N_48094,N_48019);
nor UO_38 (O_38,N_49087,N_48827);
nor UO_39 (O_39,N_48331,N_49615);
and UO_40 (O_40,N_49947,N_48978);
and UO_41 (O_41,N_49598,N_48166);
nor UO_42 (O_42,N_49513,N_49554);
or UO_43 (O_43,N_49823,N_49602);
and UO_44 (O_44,N_48516,N_49862);
and UO_45 (O_45,N_48453,N_49582);
nand UO_46 (O_46,N_48513,N_48731);
or UO_47 (O_47,N_49223,N_49106);
or UO_48 (O_48,N_49631,N_49028);
and UO_49 (O_49,N_49543,N_48990);
xor UO_50 (O_50,N_48743,N_49827);
xnor UO_51 (O_51,N_49855,N_48046);
and UO_52 (O_52,N_49140,N_49724);
or UO_53 (O_53,N_49693,N_48890);
xor UO_54 (O_54,N_49309,N_49120);
or UO_55 (O_55,N_48334,N_49437);
nor UO_56 (O_56,N_48586,N_48185);
nor UO_57 (O_57,N_49293,N_48525);
xnor UO_58 (O_58,N_48281,N_48104);
nand UO_59 (O_59,N_48913,N_49245);
and UO_60 (O_60,N_49289,N_49253);
nor UO_61 (O_61,N_48011,N_49300);
nand UO_62 (O_62,N_49585,N_48072);
or UO_63 (O_63,N_49177,N_48947);
nor UO_64 (O_64,N_49705,N_49596);
xnor UO_65 (O_65,N_48674,N_48168);
xor UO_66 (O_66,N_49677,N_48015);
or UO_67 (O_67,N_48464,N_48442);
nor UO_68 (O_68,N_49938,N_49889);
and UO_69 (O_69,N_49986,N_49813);
nor UO_70 (O_70,N_49185,N_49394);
xnor UO_71 (O_71,N_49337,N_49110);
nand UO_72 (O_72,N_48730,N_48287);
or UO_73 (O_73,N_49679,N_49727);
and UO_74 (O_74,N_49451,N_48134);
xnor UO_75 (O_75,N_48213,N_48592);
xor UO_76 (O_76,N_48652,N_49269);
xnor UO_77 (O_77,N_49860,N_49924);
and UO_78 (O_78,N_49836,N_49504);
nor UO_79 (O_79,N_48257,N_48738);
or UO_80 (O_80,N_49945,N_48122);
nand UO_81 (O_81,N_48301,N_48209);
xor UO_82 (O_82,N_49321,N_48403);
and UO_83 (O_83,N_49549,N_49193);
or UO_84 (O_84,N_48968,N_48376);
nand UO_85 (O_85,N_48520,N_49388);
and UO_86 (O_86,N_48518,N_48959);
nor UO_87 (O_87,N_49204,N_49985);
or UO_88 (O_88,N_49787,N_49670);
nor UO_89 (O_89,N_48893,N_48010);
nand UO_90 (O_90,N_49051,N_48174);
and UO_91 (O_91,N_49100,N_48207);
nor UO_92 (O_92,N_49344,N_48811);
nand UO_93 (O_93,N_49919,N_48127);
nor UO_94 (O_94,N_48970,N_48636);
or UO_95 (O_95,N_49440,N_49876);
nor UO_96 (O_96,N_48877,N_49107);
or UO_97 (O_97,N_49625,N_49061);
nor UO_98 (O_98,N_48052,N_49079);
xnor UO_99 (O_99,N_49902,N_48384);
xnor UO_100 (O_100,N_48107,N_49516);
or UO_101 (O_101,N_48723,N_49009);
nor UO_102 (O_102,N_49085,N_48038);
nor UO_103 (O_103,N_48292,N_49978);
xor UO_104 (O_104,N_48123,N_48964);
nor UO_105 (O_105,N_48489,N_48142);
nand UO_106 (O_106,N_49043,N_48492);
nand UO_107 (O_107,N_48236,N_48533);
nor UO_108 (O_108,N_49010,N_48787);
xnor UO_109 (O_109,N_48728,N_49056);
xor UO_110 (O_110,N_48883,N_48853);
or UO_111 (O_111,N_48666,N_49314);
xnor UO_112 (O_112,N_48850,N_48387);
xor UO_113 (O_113,N_48300,N_48767);
and UO_114 (O_114,N_49179,N_49152);
and UO_115 (O_115,N_48690,N_48565);
nor UO_116 (O_116,N_48626,N_49077);
nor UO_117 (O_117,N_49470,N_49268);
and UO_118 (O_118,N_49852,N_48706);
nor UO_119 (O_119,N_48870,N_48033);
nor UO_120 (O_120,N_48218,N_49760);
nor UO_121 (O_121,N_49515,N_48354);
nand UO_122 (O_122,N_49023,N_48357);
nand UO_123 (O_123,N_48697,N_48476);
nor UO_124 (O_124,N_48825,N_49383);
xnor UO_125 (O_125,N_48058,N_49046);
xnor UO_126 (O_126,N_49001,N_49932);
xnor UO_127 (O_127,N_49686,N_49117);
and UO_128 (O_128,N_48223,N_49116);
nor UO_129 (O_129,N_48112,N_49415);
nand UO_130 (O_130,N_48269,N_48278);
and UO_131 (O_131,N_48725,N_49775);
nor UO_132 (O_132,N_49772,N_49570);
nand UO_133 (O_133,N_48539,N_48608);
xnor UO_134 (O_134,N_49328,N_48936);
or UO_135 (O_135,N_48527,N_48050);
and UO_136 (O_136,N_49567,N_48397);
or UO_137 (O_137,N_49886,N_49723);
nor UO_138 (O_138,N_49916,N_49499);
nor UO_139 (O_139,N_48258,N_48399);
xor UO_140 (O_140,N_48077,N_49658);
nor UO_141 (O_141,N_49143,N_49160);
or UO_142 (O_142,N_49127,N_48715);
nor UO_143 (O_143,N_48386,N_49867);
nand UO_144 (O_144,N_49937,N_49320);
xor UO_145 (O_145,N_49398,N_49111);
nor UO_146 (O_146,N_48108,N_48101);
and UO_147 (O_147,N_48275,N_48864);
xor UO_148 (O_148,N_49771,N_48147);
nand UO_149 (O_149,N_48845,N_49015);
and UO_150 (O_150,N_48405,N_48180);
and UO_151 (O_151,N_49839,N_49846);
and UO_152 (O_152,N_48995,N_48319);
and UO_153 (O_153,N_48896,N_48103);
and UO_154 (O_154,N_49962,N_48068);
and UO_155 (O_155,N_49339,N_48559);
or UO_156 (O_156,N_48008,N_48426);
or UO_157 (O_157,N_49424,N_48139);
and UO_158 (O_158,N_48456,N_48348);
nand UO_159 (O_159,N_49044,N_48819);
xnor UO_160 (O_160,N_49207,N_48691);
and UO_161 (O_161,N_49599,N_49864);
xor UO_162 (O_162,N_49035,N_48065);
or UO_163 (O_163,N_49792,N_49538);
xor UO_164 (O_164,N_49075,N_49374);
nor UO_165 (O_165,N_49361,N_49785);
nand UO_166 (O_166,N_49783,N_48244);
nor UO_167 (O_167,N_49804,N_49395);
nand UO_168 (O_168,N_49400,N_48501);
or UO_169 (O_169,N_49149,N_48627);
xnor UO_170 (O_170,N_48702,N_49283);
xnor UO_171 (O_171,N_48698,N_48190);
or UO_172 (O_172,N_48942,N_48764);
and UO_173 (O_173,N_49552,N_48832);
and UO_174 (O_174,N_49537,N_49491);
nand UO_175 (O_175,N_48198,N_49340);
and UO_176 (O_176,N_48443,N_49489);
or UO_177 (O_177,N_48111,N_48654);
xnor UO_178 (O_178,N_49141,N_49928);
nand UO_179 (O_179,N_49995,N_49795);
or UO_180 (O_180,N_49072,N_49030);
or UO_181 (O_181,N_49545,N_49966);
nand UO_182 (O_182,N_49096,N_48914);
xnor UO_183 (O_183,N_48162,N_48847);
and UO_184 (O_184,N_48161,N_48865);
or UO_185 (O_185,N_48570,N_49069);
nand UO_186 (O_186,N_49573,N_48581);
or UO_187 (O_187,N_49237,N_49331);
nand UO_188 (O_188,N_49422,N_49575);
nor UO_189 (O_189,N_48249,N_49977);
nand UO_190 (O_190,N_48812,N_49820);
or UO_191 (O_191,N_48621,N_48984);
and UO_192 (O_192,N_48340,N_48915);
and UO_193 (O_193,N_48553,N_49119);
nor UO_194 (O_194,N_49510,N_48176);
nand UO_195 (O_195,N_49074,N_48528);
and UO_196 (O_196,N_49358,N_48991);
and UO_197 (O_197,N_49904,N_48795);
xor UO_198 (O_198,N_49536,N_48826);
nor UO_199 (O_199,N_49905,N_48140);
or UO_200 (O_200,N_49416,N_49991);
nor UO_201 (O_201,N_48635,N_49381);
nor UO_202 (O_202,N_49668,N_48951);
or UO_203 (O_203,N_49999,N_49475);
nor UO_204 (O_204,N_49448,N_48773);
nand UO_205 (O_205,N_48557,N_48171);
nand UO_206 (O_206,N_48096,N_49874);
xor UO_207 (O_207,N_48284,N_48283);
or UO_208 (O_208,N_48071,N_48113);
nor UO_209 (O_209,N_49255,N_49742);
or UO_210 (O_210,N_49605,N_48552);
or UO_211 (O_211,N_49529,N_48461);
nor UO_212 (O_212,N_48925,N_48524);
or UO_213 (O_213,N_48866,N_48831);
nand UO_214 (O_214,N_49959,N_48933);
or UO_215 (O_215,N_49464,N_49154);
xor UO_216 (O_216,N_48941,N_48742);
nor UO_217 (O_217,N_49203,N_48745);
xnor UO_218 (O_218,N_48976,N_49814);
xor UO_219 (O_219,N_49369,N_49982);
nand UO_220 (O_220,N_49908,N_49829);
or UO_221 (O_221,N_49463,N_48145);
nor UO_222 (O_222,N_48963,N_49486);
xor UO_223 (O_223,N_49115,N_48860);
nand UO_224 (O_224,N_49591,N_48656);
nand UO_225 (O_225,N_49018,N_48682);
or UO_226 (O_226,N_49547,N_49711);
nand UO_227 (O_227,N_48798,N_48302);
or UO_228 (O_228,N_48027,N_48957);
or UO_229 (O_229,N_49581,N_48818);
nand UO_230 (O_230,N_48274,N_48546);
and UO_231 (O_231,N_49642,N_49050);
nand UO_232 (O_232,N_48637,N_48882);
nor UO_233 (O_233,N_49611,N_48529);
and UO_234 (O_234,N_48517,N_49216);
nor UO_235 (O_235,N_49348,N_49685);
or UO_236 (O_236,N_49740,N_48614);
or UO_237 (O_237,N_48593,N_48303);
xnor UO_238 (O_238,N_49758,N_48829);
nor UO_239 (O_239,N_49343,N_49389);
and UO_240 (O_240,N_49007,N_48807);
nand UO_241 (O_241,N_48153,N_49965);
and UO_242 (O_242,N_49482,N_48954);
nand UO_243 (O_243,N_49461,N_48922);
nor UO_244 (O_244,N_48396,N_48076);
or UO_245 (O_245,N_49435,N_48538);
xnor UO_246 (O_246,N_48962,N_49454);
xor UO_247 (O_247,N_48341,N_48353);
nand UO_248 (O_248,N_48260,N_48509);
xnor UO_249 (O_249,N_49147,N_48351);
and UO_250 (O_250,N_49202,N_49624);
nor UO_251 (O_251,N_49040,N_48500);
and UO_252 (O_252,N_49971,N_49614);
nand UO_253 (O_253,N_49559,N_48377);
xor UO_254 (O_254,N_49684,N_49788);
nand UO_255 (O_255,N_48155,N_49586);
xnor UO_256 (O_256,N_49092,N_49907);
nor UO_257 (O_257,N_49921,N_48439);
nand UO_258 (O_258,N_49218,N_49297);
nand UO_259 (O_259,N_48642,N_48215);
and UO_260 (O_260,N_48020,N_48633);
nor UO_261 (O_261,N_49024,N_48801);
and UO_262 (O_262,N_49811,N_48115);
nor UO_263 (O_263,N_48057,N_49634);
or UO_264 (O_264,N_48918,N_49146);
nand UO_265 (O_265,N_48810,N_49666);
nor UO_266 (O_266,N_48596,N_48632);
xnor UO_267 (O_267,N_48118,N_48321);
and UO_268 (O_268,N_48708,N_49161);
xor UO_269 (O_269,N_49312,N_48335);
nand UO_270 (O_270,N_48880,N_48061);
nand UO_271 (O_271,N_48043,N_48701);
nand UO_272 (O_272,N_49101,N_49041);
nand UO_273 (O_273,N_49952,N_48371);
or UO_274 (O_274,N_48651,N_48413);
xnor UO_275 (O_275,N_48078,N_49923);
and UO_276 (O_276,N_49249,N_49483);
nor UO_277 (O_277,N_48803,N_48887);
nor UO_278 (O_278,N_49228,N_49719);
xor UO_279 (O_279,N_48734,N_48521);
and UO_280 (O_280,N_48242,N_48082);
xnor UO_281 (O_281,N_48744,N_49122);
nand UO_282 (O_282,N_49818,N_49484);
or UO_283 (O_283,N_49850,N_49583);
xnor UO_284 (O_284,N_48432,N_48707);
or UO_285 (O_285,N_49251,N_49857);
or UO_286 (O_286,N_49946,N_48450);
nand UO_287 (O_287,N_49196,N_49191);
nand UO_288 (O_288,N_49663,N_48151);
xor UO_289 (O_289,N_48202,N_48774);
and UO_290 (O_290,N_49831,N_48366);
nand UO_291 (O_291,N_49821,N_48481);
nand UO_292 (O_292,N_49329,N_49825);
xor UO_293 (O_293,N_48062,N_49326);
or UO_294 (O_294,N_49129,N_48232);
nor UO_295 (O_295,N_48458,N_48132);
or UO_296 (O_296,N_48809,N_48844);
nand UO_297 (O_297,N_48294,N_49718);
or UO_298 (O_298,N_48645,N_48781);
and UO_299 (O_299,N_48583,N_48178);
xor UO_300 (O_300,N_49338,N_49540);
or UO_301 (O_301,N_48023,N_48634);
xor UO_302 (O_302,N_49450,N_49993);
nand UO_303 (O_303,N_49005,N_49014);
nand UO_304 (O_304,N_49108,N_48813);
xor UO_305 (O_305,N_49187,N_48230);
or UO_306 (O_306,N_49696,N_49220);
nand UO_307 (O_307,N_49401,N_49425);
and UO_308 (O_308,N_48536,N_48028);
or UO_309 (O_309,N_48729,N_49812);
or UO_310 (O_310,N_48163,N_48952);
nand UO_311 (O_311,N_48234,N_48159);
nor UO_312 (O_312,N_49590,N_48541);
and UO_313 (O_313,N_48237,N_49956);
and UO_314 (O_314,N_48506,N_48551);
and UO_315 (O_315,N_49789,N_48150);
xor UO_316 (O_316,N_49651,N_48452);
xor UO_317 (O_317,N_49842,N_49743);
nand UO_318 (O_318,N_48170,N_49080);
or UO_319 (O_319,N_49619,N_49987);
nand UO_320 (O_320,N_49194,N_49533);
xnor UO_321 (O_321,N_48472,N_49459);
and UO_322 (O_322,N_49502,N_49428);
nor UO_323 (O_323,N_48259,N_48119);
nor UO_324 (O_324,N_48638,N_48624);
xor UO_325 (O_325,N_49390,N_49773);
and UO_326 (O_326,N_48051,N_48099);
or UO_327 (O_327,N_48352,N_48736);
nor UO_328 (O_328,N_49099,N_49082);
xnor UO_329 (O_329,N_48224,N_49420);
or UO_330 (O_330,N_48045,N_48675);
and UO_331 (O_331,N_49815,N_49012);
xor UO_332 (O_332,N_48316,N_48587);
xor UO_333 (O_333,N_48898,N_49915);
nand UO_334 (O_334,N_48929,N_48036);
and UO_335 (O_335,N_48868,N_48554);
nand UO_336 (O_336,N_49299,N_49863);
nor UO_337 (O_337,N_49021,N_49168);
nor UO_338 (O_338,N_49016,N_49426);
nand UO_339 (O_339,N_49020,N_48225);
and UO_340 (O_340,N_49455,N_49319);
nor UO_341 (O_341,N_49501,N_49342);
or UO_342 (O_342,N_48372,N_49148);
or UO_343 (O_343,N_49994,N_49682);
and UO_344 (O_344,N_48620,N_48394);
and UO_345 (O_345,N_49066,N_49641);
nand UO_346 (O_346,N_49166,N_48063);
nor UO_347 (O_347,N_49749,N_48980);
and UO_348 (O_348,N_49438,N_48653);
or UO_349 (O_349,N_48245,N_49121);
and UO_350 (O_350,N_49210,N_48262);
xnor UO_351 (O_351,N_48985,N_49094);
xnor UO_352 (O_352,N_49770,N_49695);
nor UO_353 (O_353,N_49488,N_48479);
nor UO_354 (O_354,N_49182,N_48598);
or UO_355 (O_355,N_49837,N_48547);
nand UO_356 (O_356,N_48875,N_49112);
or UO_357 (O_357,N_49953,N_48746);
nand UO_358 (O_358,N_49026,N_48012);
nor UO_359 (O_359,N_49519,N_49070);
or UO_360 (O_360,N_48418,N_48474);
and UO_361 (O_361,N_49282,N_49764);
nor UO_362 (O_362,N_48885,N_49310);
and UO_363 (O_363,N_49364,N_48312);
or UO_364 (O_364,N_49560,N_49188);
nand UO_365 (O_365,N_49183,N_49909);
nand UO_366 (O_366,N_49354,N_48891);
xnor UO_367 (O_367,N_48618,N_49496);
nand UO_368 (O_368,N_48772,N_49225);
nor UO_369 (O_369,N_49175,N_49920);
nand UO_370 (O_370,N_49260,N_48704);
or UO_371 (O_371,N_49988,N_49073);
xnor UO_372 (O_372,N_49278,N_48266);
or UO_373 (O_373,N_49507,N_49861);
or UO_374 (O_374,N_48713,N_48879);
xor UO_375 (O_375,N_48267,N_49532);
or UO_376 (O_376,N_49490,N_49279);
nand UO_377 (O_377,N_48408,N_49530);
nor UO_378 (O_378,N_49726,N_48345);
nor UO_379 (O_379,N_48034,N_49034);
nor UO_380 (O_380,N_49646,N_48855);
nand UO_381 (O_381,N_48235,N_48610);
xnor UO_382 (O_382,N_48393,N_48109);
and UO_383 (O_383,N_49989,N_49674);
xor UO_384 (O_384,N_49431,N_48049);
and UO_385 (O_385,N_48992,N_49049);
nand UO_386 (O_386,N_49201,N_48623);
or UO_387 (O_387,N_48889,N_48678);
or UO_388 (O_388,N_49866,N_48695);
and UO_389 (O_389,N_49700,N_49801);
xnor UO_390 (O_390,N_49277,N_48102);
nand UO_391 (O_391,N_48342,N_48808);
nor UO_392 (O_392,N_49264,N_49118);
nand UO_393 (O_393,N_49308,N_48687);
nand UO_394 (O_394,N_49518,N_48960);
or UO_395 (O_395,N_49901,N_48999);
and UO_396 (O_396,N_49613,N_48966);
nor UO_397 (O_397,N_49974,N_49423);
xnor UO_398 (O_398,N_49865,N_48669);
xnor UO_399 (O_399,N_49180,N_48498);
xor UO_400 (O_400,N_49911,N_49712);
nand UO_401 (O_401,N_48040,N_49622);
xnor UO_402 (O_402,N_48007,N_49184);
and UO_403 (O_403,N_49055,N_48226);
nand UO_404 (O_404,N_48897,N_49457);
nand UO_405 (O_405,N_48194,N_48932);
or UO_406 (O_406,N_48415,N_48582);
xnor UO_407 (O_407,N_49209,N_49013);
xor UO_408 (O_408,N_48646,N_49535);
nor UO_409 (O_409,N_49735,N_48188);
and UO_410 (O_410,N_48814,N_48931);
nor UO_411 (O_411,N_49144,N_48323);
or UO_412 (O_412,N_48722,N_48937);
nor UO_413 (O_413,N_49155,N_49178);
nand UO_414 (O_414,N_48628,N_49826);
and UO_415 (O_415,N_49480,N_48688);
nand UO_416 (O_416,N_48785,N_49137);
xor UO_417 (O_417,N_48251,N_48158);
xnor UO_418 (O_418,N_48197,N_49317);
xnor UO_419 (O_419,N_48362,N_48895);
or UO_420 (O_420,N_48741,N_49350);
xor UO_421 (O_421,N_49794,N_48116);
xnor UO_422 (O_422,N_48327,N_49276);
or UO_423 (O_423,N_49380,N_48212);
nor UO_424 (O_424,N_48422,N_48575);
and UO_425 (O_425,N_48322,N_49476);
nand UO_426 (O_426,N_49405,N_48016);
and UO_427 (O_427,N_48920,N_49360);
and UO_428 (O_428,N_49159,N_48703);
nand UO_429 (O_429,N_48711,N_49617);
and UO_430 (O_430,N_49246,N_48462);
xnor UO_431 (O_431,N_48305,N_49647);
xnor UO_432 (O_432,N_49557,N_48768);
or UO_433 (O_433,N_48700,N_48205);
and UO_434 (O_434,N_49610,N_48948);
and UO_435 (O_435,N_49652,N_49305);
nand UO_436 (O_436,N_49714,N_49741);
or UO_437 (O_437,N_48757,N_48753);
xnor UO_438 (O_438,N_48272,N_49748);
or UO_439 (O_439,N_48378,N_48542);
nor UO_440 (O_440,N_48817,N_49678);
nor UO_441 (O_441,N_49270,N_48070);
nor UO_442 (O_442,N_48208,N_49856);
or UO_443 (O_443,N_49095,N_48361);
and UO_444 (O_444,N_49135,N_49471);
and UO_445 (O_445,N_48470,N_48749);
xor UO_446 (O_446,N_49481,N_49485);
and UO_447 (O_447,N_48059,N_48297);
and UO_448 (O_448,N_49835,N_49996);
nor UO_449 (O_449,N_48469,N_48606);
and UO_450 (O_450,N_48961,N_48935);
nor UO_451 (O_451,N_48095,N_48595);
or UO_452 (O_452,N_48605,N_48858);
xor UO_453 (O_453,N_49256,N_49884);
and UO_454 (O_454,N_49163,N_49434);
nor UO_455 (O_455,N_48973,N_48114);
nor UO_456 (O_456,N_49158,N_48755);
and UO_457 (O_457,N_48169,N_48429);
and UO_458 (O_458,N_49341,N_48664);
xnor UO_459 (O_459,N_49373,N_48504);
nor UO_460 (O_460,N_49720,N_49899);
or UO_461 (O_461,N_48804,N_48263);
or UO_462 (O_462,N_48579,N_48676);
and UO_463 (O_463,N_49151,N_49566);
or UO_464 (O_464,N_48958,N_49473);
and UO_465 (O_465,N_49150,N_49528);
xnor UO_466 (O_466,N_48466,N_49311);
nand UO_467 (O_467,N_49067,N_49042);
nor UO_468 (O_468,N_49799,N_49227);
nor UO_469 (O_469,N_49247,N_49970);
xnor UO_470 (O_470,N_48017,N_49630);
nor UO_471 (O_471,N_49452,N_49038);
nor UO_472 (O_472,N_49219,N_48268);
and UO_473 (O_473,N_48981,N_49396);
or UO_474 (O_474,N_48950,N_48480);
and UO_475 (O_475,N_48383,N_49673);
nand UO_476 (O_476,N_49877,N_48568);
and UO_477 (O_477,N_48318,N_48837);
xnor UO_478 (O_478,N_49142,N_48721);
and UO_479 (O_479,N_49493,N_48238);
nand UO_480 (O_480,N_48009,N_48747);
xnor UO_481 (O_481,N_49384,N_48346);
nor UO_482 (O_482,N_49292,N_48407);
and UO_483 (O_483,N_48836,N_49002);
and UO_484 (O_484,N_49478,N_48056);
and UO_485 (O_485,N_48400,N_49565);
nand UO_486 (O_486,N_49241,N_48577);
nor UO_487 (O_487,N_49632,N_48499);
nand UO_488 (O_488,N_48609,N_49542);
nor UO_489 (O_489,N_49199,N_49828);
nor UO_490 (O_490,N_48219,N_49332);
nand UO_491 (O_491,N_49895,N_48299);
or UO_492 (O_492,N_48838,N_48983);
nand UO_493 (O_493,N_49458,N_48004);
xnor UO_494 (O_494,N_49859,N_48816);
and UO_495 (O_495,N_48279,N_49556);
nor UO_496 (O_496,N_48295,N_48600);
or UO_497 (O_497,N_49913,N_48710);
nor UO_498 (O_498,N_49654,N_48211);
nor UO_499 (O_499,N_49362,N_48449);
nand UO_500 (O_500,N_48409,N_48683);
xor UO_501 (O_501,N_48763,N_48630);
nand UO_502 (O_502,N_49534,N_48091);
nand UO_503 (O_503,N_49233,N_49392);
and UO_504 (O_504,N_48681,N_48643);
or UO_505 (O_505,N_49032,N_48996);
nand UO_506 (O_506,N_49508,N_48833);
or UO_507 (O_507,N_48899,N_48558);
and UO_508 (O_508,N_49660,N_49676);
or UO_509 (O_509,N_49307,N_48549);
or UO_510 (O_510,N_48179,N_48421);
xor UO_511 (O_511,N_49097,N_49669);
nand UO_512 (O_512,N_49649,N_48358);
and UO_513 (O_513,N_49755,N_48884);
or UO_514 (O_514,N_48607,N_48121);
nand UO_515 (O_515,N_48217,N_48876);
nand UO_516 (O_516,N_49037,N_48647);
nand UO_517 (O_517,N_49824,N_48852);
nand UO_518 (O_518,N_49505,N_48148);
or UO_519 (O_519,N_49363,N_48906);
or UO_520 (O_520,N_48945,N_49128);
and UO_521 (O_521,N_48786,N_49964);
xor UO_522 (O_522,N_49782,N_48390);
xnor UO_523 (O_523,N_49506,N_49174);
nor UO_524 (O_524,N_48714,N_48849);
xnor UO_525 (O_525,N_49304,N_48699);
xnor UO_526 (O_526,N_48888,N_48907);
xnor UO_527 (O_527,N_49205,N_49230);
nand UO_528 (O_528,N_48144,N_48967);
and UO_529 (O_529,N_48074,N_49315);
nand UO_530 (O_530,N_49918,N_48337);
and UO_531 (O_531,N_49242,N_49621);
xor UO_532 (O_532,N_48164,N_49601);
nor UO_533 (O_533,N_48756,N_48022);
xor UO_534 (O_534,N_49661,N_49261);
or UO_535 (O_535,N_49468,N_49873);
xor UO_536 (O_536,N_49291,N_49453);
and UO_537 (O_537,N_48779,N_48444);
nor UO_538 (O_538,N_48802,N_48485);
nand UO_539 (O_539,N_49777,N_49088);
xnor UO_540 (O_540,N_48523,N_48307);
nand UO_541 (O_541,N_48815,N_49206);
nor UO_542 (O_542,N_48820,N_48726);
nor UO_543 (O_543,N_49756,N_49563);
or UO_544 (O_544,N_48672,N_49819);
and UO_545 (O_545,N_49550,N_49858);
nand UO_546 (O_546,N_48460,N_48092);
xor UO_547 (O_547,N_48374,N_48783);
and UO_548 (O_548,N_49410,N_48629);
nand UO_549 (O_549,N_49318,N_48356);
and UO_550 (O_550,N_48490,N_48846);
nand UO_551 (O_551,N_49541,N_49659);
nor UO_552 (O_552,N_49402,N_49776);
nand UO_553 (O_553,N_49644,N_49665);
nor UO_554 (O_554,N_48233,N_48157);
nand UO_555 (O_555,N_48203,N_48315);
or UO_556 (O_556,N_48032,N_49868);
and UO_557 (O_557,N_48154,N_48298);
or UO_558 (O_558,N_48684,N_49136);
nor UO_559 (O_559,N_49544,N_48333);
nor UO_560 (O_560,N_48256,N_49430);
nand UO_561 (O_561,N_49347,N_49841);
nand UO_562 (O_562,N_48425,N_48921);
nor UO_563 (O_563,N_48349,N_49885);
xnor UO_564 (O_564,N_49531,N_49262);
nand UO_565 (O_565,N_48916,N_49604);
and UO_566 (O_566,N_48473,N_49134);
and UO_567 (O_567,N_49954,N_48487);
nor UO_568 (O_568,N_48350,N_48576);
nor UO_569 (O_569,N_48083,N_48613);
xor UO_570 (O_570,N_48184,N_49477);
or UO_571 (O_571,N_49997,N_49791);
xor UO_572 (O_572,N_49629,N_49058);
or UO_573 (O_573,N_48839,N_49774);
or UO_574 (O_574,N_48571,N_49059);
nand UO_575 (O_575,N_48060,N_48975);
nand UO_576 (O_576,N_48130,N_48762);
xor UO_577 (O_577,N_48661,N_48495);
or UO_578 (O_578,N_49894,N_48903);
and UO_579 (O_579,N_49235,N_49732);
nand UO_580 (O_580,N_48309,N_49503);
xor UO_581 (O_581,N_48433,N_48373);
xnor UO_582 (O_582,N_49728,N_48018);
and UO_583 (O_583,N_49145,N_48160);
or UO_584 (O_584,N_49429,N_49972);
nor UO_585 (O_585,N_49125,N_48265);
or UO_586 (O_586,N_49883,N_49834);
and UO_587 (O_587,N_49153,N_49730);
nand UO_588 (O_588,N_48006,N_49940);
nor UO_589 (O_589,N_49683,N_49271);
xor UO_590 (O_590,N_49701,N_49881);
nor UO_591 (O_591,N_48398,N_48567);
or UO_592 (O_592,N_48718,N_48594);
xnor UO_593 (O_593,N_48573,N_49466);
or UO_594 (O_594,N_48511,N_49640);
nand UO_595 (O_595,N_48243,N_49608);
xor UO_596 (O_596,N_49680,N_48972);
nand UO_597 (O_597,N_48604,N_49068);
and UO_598 (O_598,N_49892,N_48325);
nand UO_599 (O_599,N_49546,N_49737);
nor UO_600 (O_600,N_48367,N_48328);
or UO_601 (O_601,N_49284,N_48181);
or UO_602 (O_602,N_49365,N_48067);
xor UO_603 (O_603,N_49487,N_49690);
and UO_604 (O_604,N_48380,N_49745);
nand UO_605 (O_605,N_49689,N_48857);
or UO_606 (O_606,N_48663,N_49060);
xor UO_607 (O_607,N_48840,N_48037);
xor UO_608 (O_608,N_49672,N_48569);
or UO_609 (O_609,N_48477,N_48097);
nor UO_610 (O_610,N_49215,N_49912);
and UO_611 (O_611,N_49404,N_48137);
or UO_612 (O_612,N_48183,N_48044);
or UO_613 (O_613,N_48639,N_49664);
xnor UO_614 (O_614,N_48754,N_49236);
nand UO_615 (O_615,N_49694,N_48438);
and UO_616 (O_616,N_48856,N_49407);
xor UO_617 (O_617,N_48724,N_49752);
nand UO_618 (O_618,N_48270,N_49890);
or UO_619 (O_619,N_49057,N_49744);
xnor UO_620 (O_620,N_48526,N_49102);
or UO_621 (O_621,N_48339,N_49662);
nor UO_622 (O_622,N_49382,N_49303);
nor UO_623 (O_623,N_49086,N_49104);
nand UO_624 (O_624,N_48619,N_49399);
xnor UO_625 (O_625,N_49969,N_49706);
and UO_626 (O_626,N_49725,N_49620);
and UO_627 (O_627,N_48974,N_48105);
xor UO_628 (O_628,N_48901,N_49462);
and UO_629 (O_629,N_48385,N_49934);
nand UO_630 (O_630,N_48679,N_48141);
and UO_631 (O_631,N_48611,N_48406);
nor UO_632 (O_632,N_48182,N_49698);
xor UO_633 (O_633,N_48530,N_48030);
xnor UO_634 (O_634,N_48510,N_49600);
nand UO_635 (O_635,N_48874,N_48979);
or UO_636 (O_636,N_48908,N_49612);
or UO_637 (O_637,N_49418,N_48986);
xor UO_638 (O_638,N_48987,N_49564);
nand UO_639 (O_639,N_48680,N_48454);
or UO_640 (O_640,N_49047,N_49103);
or UO_641 (O_641,N_48603,N_48081);
nand UO_642 (O_642,N_49713,N_49577);
nand UO_643 (O_643,N_48780,N_48085);
xor UO_644 (O_644,N_48670,N_48759);
xnor UO_645 (O_645,N_48370,N_49845);
nor UO_646 (O_646,N_48216,N_49523);
or UO_647 (O_647,N_48693,N_49707);
and UO_648 (O_648,N_48892,N_48069);
nand UO_649 (O_649,N_49960,N_48599);
xnor UO_650 (O_650,N_48423,N_48451);
and UO_651 (O_651,N_48534,N_49633);
nor UO_652 (O_652,N_49656,N_48537);
nand UO_653 (O_653,N_49169,N_48277);
or UO_654 (O_654,N_48640,N_49753);
and UO_655 (O_655,N_48435,N_48667);
nor UO_656 (O_656,N_49936,N_49109);
nand UO_657 (O_657,N_49958,N_49022);
and UO_658 (O_658,N_48843,N_48241);
xnor UO_659 (O_659,N_49930,N_48842);
nor UO_660 (O_660,N_49848,N_48336);
nor UO_661 (O_661,N_48285,N_49627);
and UO_662 (O_662,N_48375,N_48280);
and UO_663 (O_663,N_48253,N_49951);
xnor UO_664 (O_664,N_49716,N_48494);
or UO_665 (O_665,N_49807,N_48042);
nor UO_666 (O_666,N_48293,N_49643);
xor UO_667 (O_667,N_48574,N_48794);
xnor UO_668 (O_668,N_49618,N_49164);
and UO_669 (O_669,N_49551,N_49265);
nand UO_670 (O_670,N_48201,N_49306);
nand UO_671 (O_671,N_48410,N_48555);
or UO_672 (O_672,N_48079,N_49313);
nand UO_673 (O_673,N_48463,N_48047);
xnor UO_674 (O_674,N_49967,N_49492);
nor UO_675 (O_675,N_49738,N_49927);
or UO_676 (O_676,N_49671,N_48660);
xnor UO_677 (O_677,N_49054,N_48658);
nand UO_678 (O_678,N_48512,N_49250);
nand UO_679 (O_679,N_49579,N_49432);
xor UO_680 (O_680,N_48830,N_48940);
or UO_681 (O_681,N_48193,N_48912);
and UO_682 (O_682,N_48231,N_49950);
nand UO_683 (O_683,N_48982,N_48192);
or UO_684 (O_684,N_48503,N_49465);
or UO_685 (O_685,N_49562,N_49715);
or UO_686 (O_686,N_49816,N_49514);
nor UO_687 (O_687,N_48389,N_49062);
or UO_688 (O_688,N_49222,N_48117);
nand UO_689 (O_689,N_49335,N_48196);
nand UO_690 (O_690,N_49421,N_48250);
or UO_691 (O_691,N_49181,N_48900);
or UO_692 (O_692,N_49847,N_48430);
xor UO_693 (O_693,N_48881,N_48177);
xor UO_694 (O_694,N_49132,N_49346);
nor UO_695 (O_695,N_48689,N_49790);
nand UO_696 (O_696,N_48894,N_48310);
or UO_697 (O_697,N_49746,N_49006);
xor UO_698 (O_698,N_49497,N_48001);
nand UO_699 (O_699,N_49195,N_49922);
xnor UO_700 (O_700,N_49208,N_48904);
or UO_701 (O_701,N_48943,N_48872);
and UO_702 (O_702,N_48246,N_49467);
nand UO_703 (O_703,N_49553,N_49172);
nand UO_704 (O_704,N_48195,N_48448);
xnor UO_705 (O_705,N_49170,N_49449);
xnor UO_706 (O_706,N_48649,N_49926);
nand UO_707 (O_707,N_48355,N_48392);
and UO_708 (O_708,N_48505,N_48507);
and UO_709 (O_709,N_49992,N_48080);
nor UO_710 (O_710,N_49984,N_49592);
or UO_711 (O_711,N_49657,N_48758);
nor UO_712 (O_712,N_49157,N_49784);
or UO_713 (O_713,N_48644,N_49896);
nor UO_714 (O_714,N_49761,N_48748);
and UO_715 (O_715,N_49650,N_48191);
nor UO_716 (O_716,N_49213,N_48412);
and UO_717 (O_717,N_49780,N_48686);
or UO_718 (O_718,N_48617,N_48793);
or UO_719 (O_719,N_49525,N_48591);
nor UO_720 (O_720,N_49655,N_49123);
and UO_721 (O_721,N_48326,N_49248);
or UO_722 (O_722,N_49244,N_49809);
nand UO_723 (O_723,N_49257,N_49653);
nor UO_724 (O_724,N_49584,N_48014);
nand UO_725 (O_725,N_48465,N_49469);
or UO_726 (O_726,N_49139,N_49444);
nor UO_727 (O_727,N_49699,N_49870);
xnor UO_728 (O_728,N_49687,N_48560);
nand UO_729 (O_729,N_49763,N_48338);
nor UO_730 (O_730,N_49635,N_49708);
or UO_731 (O_731,N_49387,N_49555);
and UO_732 (O_732,N_49607,N_48344);
and UO_733 (O_733,N_49833,N_49372);
or UO_734 (O_734,N_49762,N_48752);
xnor UO_735 (O_735,N_48156,N_49393);
nor UO_736 (O_736,N_49286,N_49838);
or UO_737 (O_737,N_48612,N_48308);
and UO_738 (O_738,N_49330,N_48437);
or UO_739 (O_739,N_48424,N_49378);
or UO_740 (O_740,N_48550,N_49869);
nand UO_741 (O_741,N_48491,N_48716);
xor UO_742 (O_742,N_48317,N_49875);
nand UO_743 (O_743,N_49681,N_48622);
and UO_744 (O_744,N_49081,N_49793);
xor UO_745 (O_745,N_49301,N_48597);
nor UO_746 (O_746,N_49356,N_49456);
xnor UO_747 (O_747,N_49366,N_49093);
or UO_748 (O_748,N_49190,N_48905);
and UO_749 (O_749,N_49084,N_49322);
or UO_750 (O_750,N_49280,N_48531);
xnor UO_751 (O_751,N_48388,N_49786);
nand UO_752 (O_752,N_48075,N_48100);
nand UO_753 (O_753,N_49767,N_48093);
nor UO_754 (O_754,N_48311,N_49808);
nor UO_755 (O_755,N_48304,N_49302);
xor UO_756 (O_756,N_49721,N_49124);
and UO_757 (O_757,N_49000,N_49805);
or UO_758 (O_758,N_48431,N_49955);
xor UO_759 (O_759,N_49691,N_48589);
nand UO_760 (O_760,N_48005,N_48368);
xor UO_761 (O_761,N_49351,N_48329);
nand UO_762 (O_762,N_49281,N_49403);
xor UO_763 (O_763,N_48993,N_49368);
xor UO_764 (O_764,N_48543,N_48737);
and UO_765 (O_765,N_48578,N_49447);
xnor UO_766 (O_766,N_48126,N_48120);
nor UO_767 (O_767,N_48025,N_49512);
nor UO_768 (O_768,N_48732,N_49090);
and UO_769 (O_769,N_48347,N_48288);
and UO_770 (O_770,N_49105,N_48416);
nand UO_771 (O_771,N_49981,N_48939);
nand UO_772 (O_772,N_48615,N_49334);
xnor UO_773 (O_773,N_49949,N_49925);
xnor UO_774 (O_774,N_49980,N_49290);
xor UO_775 (O_775,N_48544,N_49446);
or UO_776 (O_776,N_49976,N_48359);
nor UO_777 (O_777,N_49439,N_48769);
xnor UO_778 (O_778,N_49990,N_48146);
and UO_779 (O_779,N_48616,N_48135);
xnor UO_780 (O_780,N_49272,N_49033);
xnor UO_781 (O_781,N_48247,N_48402);
nor UO_782 (O_782,N_48210,N_48761);
nand UO_783 (O_783,N_49910,N_49173);
nand UO_784 (O_784,N_48110,N_49433);
xor UO_785 (O_785,N_49628,N_48601);
or UO_786 (O_786,N_49323,N_48214);
xor UO_787 (O_787,N_48420,N_48419);
nand UO_788 (O_788,N_49568,N_48938);
xor UO_789 (O_789,N_48776,N_49212);
nor UO_790 (O_790,N_48035,N_48173);
nor UO_791 (O_791,N_49587,N_48414);
nor UO_792 (O_792,N_48306,N_48923);
and UO_793 (O_793,N_49769,N_48563);
and UO_794 (O_794,N_48276,N_48475);
xor UO_795 (O_795,N_48343,N_49597);
and UO_796 (O_796,N_49511,N_48720);
xor UO_797 (O_797,N_48221,N_49285);
xnor UO_798 (O_798,N_49065,N_48871);
or UO_799 (O_799,N_48282,N_49854);
or UO_800 (O_800,N_48861,N_49052);
nor UO_801 (O_801,N_49239,N_49667);
or UO_802 (O_802,N_49474,N_48564);
nor UO_803 (O_803,N_49259,N_49064);
nor UO_804 (O_804,N_48084,N_49810);
nor UO_805 (O_805,N_49045,N_49349);
and UO_806 (O_806,N_49526,N_48199);
and UO_807 (O_807,N_48822,N_49871);
or UO_808 (O_808,N_48971,N_48694);
xnor UO_809 (O_809,N_49234,N_49498);
and UO_810 (O_810,N_49797,N_48824);
nand UO_811 (O_811,N_48483,N_49998);
or UO_812 (O_812,N_49031,N_48227);
or UO_813 (O_813,N_49840,N_48048);
or UO_814 (O_814,N_48873,N_49638);
xor UO_815 (O_815,N_48482,N_49603);
nor UO_816 (O_816,N_48522,N_49025);
or UO_817 (O_817,N_48910,N_48189);
xor UO_818 (O_818,N_49806,N_48788);
xor UO_819 (O_819,N_49703,N_49114);
or UO_820 (O_820,N_48791,N_49539);
nand UO_821 (O_821,N_48417,N_49232);
or UO_822 (O_822,N_48187,N_48834);
nand UO_823 (O_823,N_49379,N_48705);
and UO_824 (O_824,N_48024,N_48073);
or UO_825 (O_825,N_48286,N_49412);
xnor UO_826 (O_826,N_49240,N_49238);
nor UO_827 (O_827,N_49750,N_48200);
xnor UO_828 (O_828,N_49802,N_49853);
or UO_829 (O_829,N_48806,N_49288);
and UO_830 (O_830,N_49759,N_49414);
xor UO_831 (O_831,N_49594,N_48427);
nand UO_832 (O_832,N_48434,N_48733);
nor UO_833 (O_833,N_48296,N_48446);
nor UO_834 (O_834,N_49409,N_48648);
and UO_835 (O_835,N_49830,N_49411);
xnor UO_836 (O_836,N_49494,N_49832);
or UO_837 (O_837,N_49844,N_48548);
xor UO_838 (O_838,N_49849,N_48911);
or UO_839 (O_839,N_48457,N_49327);
and UO_840 (O_840,N_49798,N_48851);
xnor UO_841 (O_841,N_48631,N_48994);
xor UO_842 (O_842,N_49942,N_49029);
and UO_843 (O_843,N_48445,N_49524);
and UO_844 (O_844,N_49126,N_49355);
and UO_845 (O_845,N_48222,N_48775);
nor UO_846 (O_846,N_49472,N_49580);
or UO_847 (O_847,N_48590,N_49083);
nand UO_848 (O_848,N_48668,N_48382);
xnor UO_849 (O_849,N_49595,N_49757);
xnor UO_850 (O_850,N_48459,N_48930);
and UO_851 (O_851,N_49397,N_49296);
or UO_852 (O_852,N_49039,N_49882);
xnor UO_853 (O_853,N_49214,N_49294);
and UO_854 (O_854,N_48488,N_49071);
nor UO_855 (O_855,N_48314,N_48771);
xor UO_856 (O_856,N_48540,N_49287);
nor UO_857 (O_857,N_48515,N_48496);
and UO_858 (O_858,N_49091,N_49961);
or UO_859 (O_859,N_48089,N_48138);
or UO_860 (O_860,N_49509,N_49019);
and UO_861 (O_861,N_49263,N_49975);
nand UO_862 (O_862,N_48248,N_49521);
or UO_863 (O_863,N_48902,N_49803);
xnor UO_864 (O_864,N_48740,N_48365);
nand UO_865 (O_865,N_49224,N_48029);
nand UO_866 (O_866,N_48919,N_48098);
or UO_867 (O_867,N_49729,N_49800);
and UO_868 (O_868,N_48324,N_49367);
xnor UO_869 (O_869,N_48867,N_48502);
nor UO_870 (O_870,N_49593,N_49275);
and UO_871 (O_871,N_49822,N_48254);
and UO_872 (O_872,N_48671,N_48395);
xnor UO_873 (O_873,N_49851,N_49872);
nor UO_874 (O_874,N_49011,N_49747);
nor UO_875 (O_875,N_49903,N_49098);
or UO_876 (O_876,N_49217,N_48625);
or UO_877 (O_877,N_48588,N_49419);
and UO_878 (O_878,N_48514,N_48363);
nor UO_879 (O_879,N_49944,N_49391);
and UO_880 (O_880,N_48997,N_49231);
nand UO_881 (O_881,N_49324,N_49688);
xnor UO_882 (O_882,N_48436,N_48519);
nor UO_883 (O_883,N_48369,N_49186);
or UO_884 (O_884,N_48330,N_48719);
xor UO_885 (O_885,N_48805,N_49626);
xnor UO_886 (O_886,N_48869,N_49443);
xnor UO_887 (O_887,N_49113,N_49200);
nand UO_888 (O_888,N_48641,N_49983);
xor UO_889 (O_889,N_48255,N_48440);
and UO_890 (O_890,N_49717,N_48064);
nor UO_891 (O_891,N_49008,N_48125);
xnor UO_892 (O_892,N_49266,N_48717);
nor UO_893 (O_893,N_49336,N_48750);
xor UO_894 (O_894,N_48739,N_48662);
xnor UO_895 (O_895,N_49375,N_49891);
or UO_896 (O_896,N_48149,N_48136);
and UO_897 (O_897,N_49385,N_48956);
and UO_898 (O_898,N_48471,N_49003);
and UO_899 (O_899,N_48204,N_48790);
nand UO_900 (O_900,N_49692,N_49436);
or UO_901 (O_901,N_48859,N_48789);
xor UO_902 (O_902,N_48909,N_48013);
xor UO_903 (O_903,N_48828,N_48261);
xnor UO_904 (O_904,N_49371,N_49751);
or UO_905 (O_905,N_49765,N_48129);
or UO_906 (O_906,N_49517,N_48381);
nand UO_907 (O_907,N_48778,N_49352);
or UO_908 (O_908,N_49778,N_48585);
and UO_909 (O_909,N_48508,N_49258);
xor UO_910 (O_910,N_48264,N_48039);
nor UO_911 (O_911,N_48003,N_49131);
xnor UO_912 (O_912,N_48677,N_49574);
xnor UO_913 (O_913,N_48055,N_49520);
xnor UO_914 (O_914,N_49442,N_49623);
xor UO_915 (O_915,N_49817,N_49171);
nand UO_916 (O_916,N_49941,N_48240);
or UO_917 (O_917,N_48455,N_48657);
and UO_918 (O_918,N_49427,N_48580);
nor UO_919 (O_919,N_48000,N_49130);
and UO_920 (O_920,N_49176,N_48186);
nand UO_921 (O_921,N_49935,N_48650);
xnor UO_922 (O_922,N_49252,N_48447);
nand UO_923 (O_923,N_49576,N_49353);
or UO_924 (O_924,N_49906,N_49736);
and UO_925 (O_925,N_49017,N_49754);
nand UO_926 (O_926,N_49843,N_48797);
nand UO_927 (O_927,N_49929,N_49522);
nand UO_928 (O_928,N_48379,N_49914);
and UO_929 (O_929,N_49731,N_49548);
xnor UO_930 (O_930,N_48167,N_49192);
or UO_931 (O_931,N_48659,N_49917);
nor UO_932 (O_932,N_48561,N_49933);
nor UO_933 (O_933,N_48320,N_49370);
nand UO_934 (O_934,N_48572,N_48841);
nand UO_935 (O_935,N_49162,N_48584);
and UO_936 (O_936,N_48562,N_49156);
and UO_937 (O_937,N_49133,N_49957);
nand UO_938 (O_938,N_49878,N_48665);
nor UO_939 (O_939,N_49880,N_49243);
nor UO_940 (O_940,N_48969,N_48770);
nand UO_941 (O_941,N_49578,N_48796);
nor UO_942 (O_942,N_49036,N_49704);
or UO_943 (O_943,N_49887,N_49325);
nand UO_944 (O_944,N_48133,N_49413);
nand UO_945 (O_945,N_49639,N_48493);
and UO_946 (O_946,N_48917,N_49254);
nor UO_947 (O_947,N_48239,N_49734);
nand UO_948 (O_948,N_48566,N_48777);
and UO_949 (O_949,N_48766,N_48799);
xnor UO_950 (O_950,N_48106,N_49298);
and UO_951 (O_951,N_48545,N_49572);
nand UO_952 (O_952,N_48751,N_49027);
nand UO_953 (O_953,N_49316,N_48478);
nor UO_954 (O_954,N_48782,N_49357);
xor UO_955 (O_955,N_49571,N_48886);
or UO_956 (O_956,N_48927,N_49376);
or UO_957 (O_957,N_48271,N_48484);
nand UO_958 (O_958,N_49939,N_49078);
nor UO_959 (O_959,N_49943,N_48165);
nor UO_960 (O_960,N_48735,N_48128);
and UO_961 (O_961,N_48090,N_49527);
and UO_962 (O_962,N_48290,N_48696);
or UO_963 (O_963,N_49963,N_48273);
or UO_964 (O_964,N_48252,N_49274);
and UO_965 (O_965,N_49973,N_48934);
nand UO_966 (O_966,N_48291,N_49636);
and UO_967 (O_967,N_49637,N_48989);
nand UO_968 (O_968,N_49616,N_49879);
xor UO_969 (O_969,N_48332,N_49979);
and UO_970 (O_970,N_49053,N_49004);
xnor UO_971 (O_971,N_48532,N_48673);
nand UO_972 (O_972,N_49733,N_49359);
xnor UO_973 (O_973,N_48053,N_48712);
nor UO_974 (O_974,N_49408,N_49648);
nand UO_975 (O_975,N_48926,N_48988);
nand UO_976 (O_976,N_48602,N_48066);
and UO_977 (O_977,N_48220,N_49273);
or UO_978 (O_978,N_49569,N_49226);
and UO_979 (O_979,N_49267,N_48468);
nand UO_980 (O_980,N_48784,N_49710);
nor UO_981 (O_981,N_49558,N_48863);
xnor UO_982 (O_982,N_49377,N_48862);
and UO_983 (O_983,N_49063,N_48143);
nand UO_984 (O_984,N_48124,N_48823);
nand UO_985 (O_985,N_48172,N_48655);
or UO_986 (O_986,N_48949,N_48206);
and UO_987 (O_987,N_48002,N_48152);
or UO_988 (O_988,N_49606,N_49197);
xnor UO_989 (O_989,N_49333,N_48685);
or UO_990 (O_990,N_48289,N_48535);
and UO_991 (O_991,N_48486,N_49417);
nand UO_992 (O_992,N_48928,N_48026);
xor UO_993 (O_993,N_48086,N_49211);
nand UO_994 (O_994,N_49739,N_49722);
nand UO_995 (O_995,N_48946,N_48313);
or UO_996 (O_996,N_48727,N_48760);
or UO_997 (O_997,N_48854,N_49968);
xnor UO_998 (O_998,N_49495,N_48087);
and UO_999 (O_999,N_49931,N_49386);
or UO_1000 (O_1000,N_49423,N_49379);
xor UO_1001 (O_1001,N_49193,N_48318);
nand UO_1002 (O_1002,N_48871,N_49627);
nor UO_1003 (O_1003,N_48146,N_48151);
xnor UO_1004 (O_1004,N_49942,N_48891);
and UO_1005 (O_1005,N_48009,N_48578);
nand UO_1006 (O_1006,N_48625,N_48145);
and UO_1007 (O_1007,N_49240,N_49389);
and UO_1008 (O_1008,N_48227,N_49605);
or UO_1009 (O_1009,N_49937,N_49500);
nor UO_1010 (O_1010,N_48801,N_48867);
xor UO_1011 (O_1011,N_49966,N_49864);
xnor UO_1012 (O_1012,N_48461,N_49230);
nor UO_1013 (O_1013,N_48120,N_49974);
or UO_1014 (O_1014,N_49649,N_49328);
nor UO_1015 (O_1015,N_48074,N_49400);
nor UO_1016 (O_1016,N_49011,N_48767);
and UO_1017 (O_1017,N_48383,N_49008);
and UO_1018 (O_1018,N_49576,N_49931);
xor UO_1019 (O_1019,N_49008,N_49025);
and UO_1020 (O_1020,N_48201,N_48496);
nand UO_1021 (O_1021,N_49264,N_49939);
nand UO_1022 (O_1022,N_49970,N_48920);
and UO_1023 (O_1023,N_48662,N_49095);
xor UO_1024 (O_1024,N_48445,N_48205);
nor UO_1025 (O_1025,N_49038,N_49145);
nand UO_1026 (O_1026,N_48669,N_48411);
xnor UO_1027 (O_1027,N_49640,N_48895);
nor UO_1028 (O_1028,N_48769,N_49582);
nor UO_1029 (O_1029,N_49898,N_48798);
xor UO_1030 (O_1030,N_49801,N_49943);
and UO_1031 (O_1031,N_49741,N_48188);
and UO_1032 (O_1032,N_49935,N_49614);
nor UO_1033 (O_1033,N_48539,N_49804);
or UO_1034 (O_1034,N_49700,N_49083);
and UO_1035 (O_1035,N_48222,N_49189);
and UO_1036 (O_1036,N_49298,N_49747);
and UO_1037 (O_1037,N_48827,N_48293);
xnor UO_1038 (O_1038,N_49217,N_48589);
nand UO_1039 (O_1039,N_48222,N_49034);
or UO_1040 (O_1040,N_48021,N_49027);
xnor UO_1041 (O_1041,N_49967,N_49447);
nor UO_1042 (O_1042,N_48721,N_48093);
nand UO_1043 (O_1043,N_48252,N_49358);
or UO_1044 (O_1044,N_48317,N_49939);
nand UO_1045 (O_1045,N_49500,N_49310);
and UO_1046 (O_1046,N_49627,N_49006);
or UO_1047 (O_1047,N_48051,N_49535);
or UO_1048 (O_1048,N_48425,N_49861);
or UO_1049 (O_1049,N_49697,N_48307);
nand UO_1050 (O_1050,N_49145,N_49720);
or UO_1051 (O_1051,N_48338,N_49319);
nor UO_1052 (O_1052,N_49581,N_48003);
nor UO_1053 (O_1053,N_49396,N_48356);
nor UO_1054 (O_1054,N_48558,N_48970);
xor UO_1055 (O_1055,N_49460,N_48624);
nand UO_1056 (O_1056,N_49442,N_49183);
xor UO_1057 (O_1057,N_48675,N_49511);
nand UO_1058 (O_1058,N_48345,N_49036);
nor UO_1059 (O_1059,N_49959,N_48645);
or UO_1060 (O_1060,N_48462,N_49546);
xnor UO_1061 (O_1061,N_48961,N_48331);
or UO_1062 (O_1062,N_49490,N_48589);
and UO_1063 (O_1063,N_48428,N_49421);
or UO_1064 (O_1064,N_49381,N_48527);
xor UO_1065 (O_1065,N_49729,N_49533);
or UO_1066 (O_1066,N_48974,N_49000);
and UO_1067 (O_1067,N_49766,N_48489);
nor UO_1068 (O_1068,N_48372,N_48414);
nor UO_1069 (O_1069,N_49759,N_49337);
and UO_1070 (O_1070,N_48770,N_49341);
or UO_1071 (O_1071,N_48853,N_49229);
xnor UO_1072 (O_1072,N_48689,N_48423);
xnor UO_1073 (O_1073,N_48103,N_48413);
xor UO_1074 (O_1074,N_48616,N_48923);
or UO_1075 (O_1075,N_48215,N_48557);
nor UO_1076 (O_1076,N_49895,N_49814);
nand UO_1077 (O_1077,N_49140,N_49865);
or UO_1078 (O_1078,N_48264,N_48012);
and UO_1079 (O_1079,N_49228,N_49849);
and UO_1080 (O_1080,N_48670,N_48225);
or UO_1081 (O_1081,N_49050,N_48210);
and UO_1082 (O_1082,N_48559,N_49020);
and UO_1083 (O_1083,N_49096,N_48174);
nand UO_1084 (O_1084,N_49867,N_48391);
nor UO_1085 (O_1085,N_48449,N_49431);
and UO_1086 (O_1086,N_48529,N_48831);
or UO_1087 (O_1087,N_49584,N_49206);
nand UO_1088 (O_1088,N_49789,N_49856);
xor UO_1089 (O_1089,N_48847,N_48457);
or UO_1090 (O_1090,N_48785,N_49449);
and UO_1091 (O_1091,N_48123,N_48790);
nand UO_1092 (O_1092,N_49248,N_49166);
and UO_1093 (O_1093,N_49505,N_48674);
or UO_1094 (O_1094,N_48679,N_49726);
and UO_1095 (O_1095,N_48694,N_49490);
and UO_1096 (O_1096,N_49522,N_48495);
or UO_1097 (O_1097,N_48498,N_49100);
nand UO_1098 (O_1098,N_48952,N_48854);
or UO_1099 (O_1099,N_48539,N_49615);
and UO_1100 (O_1100,N_48044,N_48473);
nand UO_1101 (O_1101,N_48702,N_49547);
or UO_1102 (O_1102,N_48894,N_48948);
nor UO_1103 (O_1103,N_48103,N_48010);
nand UO_1104 (O_1104,N_49793,N_49726);
or UO_1105 (O_1105,N_49022,N_49324);
nor UO_1106 (O_1106,N_49221,N_48154);
nor UO_1107 (O_1107,N_48624,N_49239);
nor UO_1108 (O_1108,N_49577,N_48112);
and UO_1109 (O_1109,N_48438,N_49965);
and UO_1110 (O_1110,N_49938,N_48295);
and UO_1111 (O_1111,N_48692,N_49270);
or UO_1112 (O_1112,N_49921,N_49753);
xor UO_1113 (O_1113,N_48637,N_49878);
and UO_1114 (O_1114,N_48675,N_49650);
nor UO_1115 (O_1115,N_48128,N_49744);
or UO_1116 (O_1116,N_49393,N_49873);
and UO_1117 (O_1117,N_48328,N_48237);
nand UO_1118 (O_1118,N_49640,N_49427);
xnor UO_1119 (O_1119,N_48421,N_48865);
and UO_1120 (O_1120,N_48929,N_48623);
or UO_1121 (O_1121,N_48132,N_49821);
or UO_1122 (O_1122,N_49857,N_49189);
or UO_1123 (O_1123,N_49836,N_48499);
nand UO_1124 (O_1124,N_48228,N_49006);
nor UO_1125 (O_1125,N_49466,N_48333);
or UO_1126 (O_1126,N_48860,N_48286);
and UO_1127 (O_1127,N_49154,N_48816);
nand UO_1128 (O_1128,N_49979,N_48962);
and UO_1129 (O_1129,N_49178,N_49277);
or UO_1130 (O_1130,N_48546,N_48666);
xnor UO_1131 (O_1131,N_48788,N_48936);
nor UO_1132 (O_1132,N_49609,N_48620);
nor UO_1133 (O_1133,N_49320,N_48925);
and UO_1134 (O_1134,N_49946,N_48683);
nor UO_1135 (O_1135,N_49240,N_48642);
and UO_1136 (O_1136,N_49338,N_49025);
xor UO_1137 (O_1137,N_48861,N_49948);
nor UO_1138 (O_1138,N_49763,N_48439);
and UO_1139 (O_1139,N_48739,N_48187);
nor UO_1140 (O_1140,N_48334,N_48887);
and UO_1141 (O_1141,N_48105,N_48072);
or UO_1142 (O_1142,N_49332,N_49900);
nor UO_1143 (O_1143,N_48319,N_49797);
nand UO_1144 (O_1144,N_49990,N_48751);
or UO_1145 (O_1145,N_49567,N_48536);
nor UO_1146 (O_1146,N_49413,N_48046);
or UO_1147 (O_1147,N_48350,N_49502);
nand UO_1148 (O_1148,N_48648,N_48360);
xnor UO_1149 (O_1149,N_48816,N_48106);
nor UO_1150 (O_1150,N_48472,N_49224);
or UO_1151 (O_1151,N_48613,N_48022);
or UO_1152 (O_1152,N_48836,N_49875);
or UO_1153 (O_1153,N_48098,N_48130);
and UO_1154 (O_1154,N_49320,N_49050);
nor UO_1155 (O_1155,N_49197,N_49115);
nand UO_1156 (O_1156,N_48769,N_49724);
xor UO_1157 (O_1157,N_48095,N_48305);
or UO_1158 (O_1158,N_49859,N_49289);
or UO_1159 (O_1159,N_49401,N_48554);
and UO_1160 (O_1160,N_49475,N_49817);
nor UO_1161 (O_1161,N_49030,N_49683);
nor UO_1162 (O_1162,N_49611,N_48169);
and UO_1163 (O_1163,N_48272,N_49205);
xor UO_1164 (O_1164,N_48280,N_48552);
and UO_1165 (O_1165,N_49900,N_48719);
nor UO_1166 (O_1166,N_49969,N_49574);
nand UO_1167 (O_1167,N_49806,N_49135);
and UO_1168 (O_1168,N_48955,N_48608);
nand UO_1169 (O_1169,N_49707,N_49579);
nand UO_1170 (O_1170,N_48080,N_48189);
nand UO_1171 (O_1171,N_49535,N_49608);
nand UO_1172 (O_1172,N_48528,N_48681);
nand UO_1173 (O_1173,N_49162,N_48763);
or UO_1174 (O_1174,N_48682,N_49388);
and UO_1175 (O_1175,N_49356,N_48311);
or UO_1176 (O_1176,N_48313,N_48602);
or UO_1177 (O_1177,N_49412,N_49947);
nand UO_1178 (O_1178,N_49774,N_48791);
nor UO_1179 (O_1179,N_49338,N_49670);
xor UO_1180 (O_1180,N_49690,N_49683);
nand UO_1181 (O_1181,N_49541,N_49610);
or UO_1182 (O_1182,N_49869,N_48478);
nor UO_1183 (O_1183,N_48011,N_49317);
and UO_1184 (O_1184,N_48831,N_48004);
nand UO_1185 (O_1185,N_49162,N_48851);
nor UO_1186 (O_1186,N_49091,N_49441);
nor UO_1187 (O_1187,N_48522,N_48032);
xnor UO_1188 (O_1188,N_48581,N_49872);
nor UO_1189 (O_1189,N_49316,N_48981);
xor UO_1190 (O_1190,N_48312,N_48326);
or UO_1191 (O_1191,N_48310,N_48758);
nor UO_1192 (O_1192,N_49794,N_49107);
or UO_1193 (O_1193,N_49025,N_48840);
nand UO_1194 (O_1194,N_48805,N_48407);
xor UO_1195 (O_1195,N_48665,N_49612);
xor UO_1196 (O_1196,N_49279,N_48886);
and UO_1197 (O_1197,N_48817,N_48738);
or UO_1198 (O_1198,N_48785,N_49434);
and UO_1199 (O_1199,N_48194,N_48460);
or UO_1200 (O_1200,N_48543,N_49406);
and UO_1201 (O_1201,N_49485,N_48629);
nor UO_1202 (O_1202,N_49789,N_49874);
nor UO_1203 (O_1203,N_49105,N_49009);
nand UO_1204 (O_1204,N_49918,N_48263);
and UO_1205 (O_1205,N_49708,N_48333);
nor UO_1206 (O_1206,N_49565,N_48179);
xor UO_1207 (O_1207,N_49072,N_49247);
nor UO_1208 (O_1208,N_49664,N_48381);
nor UO_1209 (O_1209,N_48338,N_48896);
nand UO_1210 (O_1210,N_49565,N_48504);
xor UO_1211 (O_1211,N_49768,N_49263);
nand UO_1212 (O_1212,N_49975,N_48817);
nor UO_1213 (O_1213,N_49323,N_48112);
and UO_1214 (O_1214,N_49449,N_49341);
or UO_1215 (O_1215,N_49879,N_49519);
or UO_1216 (O_1216,N_48622,N_48852);
or UO_1217 (O_1217,N_49381,N_49217);
nor UO_1218 (O_1218,N_48973,N_49383);
xor UO_1219 (O_1219,N_49552,N_49523);
nand UO_1220 (O_1220,N_49439,N_49317);
nand UO_1221 (O_1221,N_49604,N_48949);
and UO_1222 (O_1222,N_48298,N_49694);
and UO_1223 (O_1223,N_49160,N_49981);
nand UO_1224 (O_1224,N_48211,N_49238);
xnor UO_1225 (O_1225,N_48362,N_49562);
and UO_1226 (O_1226,N_49278,N_48976);
and UO_1227 (O_1227,N_49993,N_48534);
or UO_1228 (O_1228,N_49636,N_48045);
nand UO_1229 (O_1229,N_48063,N_48164);
xnor UO_1230 (O_1230,N_49997,N_49086);
nand UO_1231 (O_1231,N_48364,N_49985);
nand UO_1232 (O_1232,N_49509,N_49285);
nor UO_1233 (O_1233,N_49835,N_48790);
xnor UO_1234 (O_1234,N_49539,N_49237);
and UO_1235 (O_1235,N_48414,N_49231);
xnor UO_1236 (O_1236,N_49765,N_49992);
nand UO_1237 (O_1237,N_48971,N_49390);
or UO_1238 (O_1238,N_49360,N_48577);
and UO_1239 (O_1239,N_49296,N_48752);
nand UO_1240 (O_1240,N_48698,N_48407);
xnor UO_1241 (O_1241,N_48725,N_49456);
or UO_1242 (O_1242,N_49839,N_49126);
xor UO_1243 (O_1243,N_48325,N_48784);
nor UO_1244 (O_1244,N_49231,N_48394);
nor UO_1245 (O_1245,N_49627,N_49346);
xor UO_1246 (O_1246,N_48619,N_48961);
nand UO_1247 (O_1247,N_49616,N_48386);
xor UO_1248 (O_1248,N_48730,N_49667);
nand UO_1249 (O_1249,N_49525,N_49816);
nand UO_1250 (O_1250,N_49173,N_49647);
xnor UO_1251 (O_1251,N_49130,N_49443);
and UO_1252 (O_1252,N_48049,N_49581);
nand UO_1253 (O_1253,N_48414,N_49248);
nor UO_1254 (O_1254,N_49660,N_49566);
nor UO_1255 (O_1255,N_48631,N_49560);
nor UO_1256 (O_1256,N_48281,N_49670);
nor UO_1257 (O_1257,N_49258,N_49215);
nand UO_1258 (O_1258,N_49575,N_48959);
nor UO_1259 (O_1259,N_48837,N_49501);
and UO_1260 (O_1260,N_49967,N_48709);
nand UO_1261 (O_1261,N_49080,N_48549);
nand UO_1262 (O_1262,N_48955,N_48749);
xnor UO_1263 (O_1263,N_49193,N_49228);
and UO_1264 (O_1264,N_49048,N_49604);
and UO_1265 (O_1265,N_49043,N_48135);
or UO_1266 (O_1266,N_48939,N_48885);
nand UO_1267 (O_1267,N_48111,N_49714);
or UO_1268 (O_1268,N_49656,N_49828);
nand UO_1269 (O_1269,N_48156,N_48678);
and UO_1270 (O_1270,N_49009,N_49067);
xor UO_1271 (O_1271,N_48003,N_49453);
or UO_1272 (O_1272,N_48392,N_49241);
xnor UO_1273 (O_1273,N_48271,N_49225);
or UO_1274 (O_1274,N_49257,N_48141);
xor UO_1275 (O_1275,N_48997,N_49814);
xor UO_1276 (O_1276,N_49802,N_49817);
nand UO_1277 (O_1277,N_49743,N_48189);
nor UO_1278 (O_1278,N_49130,N_48388);
nand UO_1279 (O_1279,N_48076,N_49028);
nand UO_1280 (O_1280,N_49860,N_48869);
nor UO_1281 (O_1281,N_49707,N_48391);
nor UO_1282 (O_1282,N_48528,N_48914);
nor UO_1283 (O_1283,N_49201,N_48183);
nand UO_1284 (O_1284,N_49063,N_49433);
nor UO_1285 (O_1285,N_48762,N_48553);
and UO_1286 (O_1286,N_48001,N_49182);
nand UO_1287 (O_1287,N_48494,N_48396);
and UO_1288 (O_1288,N_49712,N_49777);
and UO_1289 (O_1289,N_49445,N_48449);
or UO_1290 (O_1290,N_49426,N_49456);
xor UO_1291 (O_1291,N_48963,N_49768);
nand UO_1292 (O_1292,N_48064,N_48931);
xor UO_1293 (O_1293,N_48638,N_49762);
or UO_1294 (O_1294,N_49935,N_49615);
xor UO_1295 (O_1295,N_49327,N_49433);
or UO_1296 (O_1296,N_48132,N_48981);
nor UO_1297 (O_1297,N_48588,N_49660);
nor UO_1298 (O_1298,N_49737,N_48290);
or UO_1299 (O_1299,N_49702,N_48022);
or UO_1300 (O_1300,N_49185,N_48675);
xor UO_1301 (O_1301,N_48371,N_49561);
xor UO_1302 (O_1302,N_49670,N_49281);
or UO_1303 (O_1303,N_48372,N_48200);
and UO_1304 (O_1304,N_49595,N_48689);
nor UO_1305 (O_1305,N_48391,N_48011);
and UO_1306 (O_1306,N_48256,N_48762);
xor UO_1307 (O_1307,N_49862,N_48793);
nor UO_1308 (O_1308,N_48288,N_49292);
or UO_1309 (O_1309,N_49377,N_49298);
or UO_1310 (O_1310,N_49543,N_48657);
nor UO_1311 (O_1311,N_48597,N_48860);
or UO_1312 (O_1312,N_49389,N_48710);
or UO_1313 (O_1313,N_49848,N_49364);
nand UO_1314 (O_1314,N_48904,N_48481);
xnor UO_1315 (O_1315,N_49431,N_49784);
nor UO_1316 (O_1316,N_49712,N_49702);
or UO_1317 (O_1317,N_48357,N_49365);
xor UO_1318 (O_1318,N_48102,N_48141);
nor UO_1319 (O_1319,N_49211,N_48973);
and UO_1320 (O_1320,N_48038,N_48123);
nand UO_1321 (O_1321,N_49780,N_49266);
nand UO_1322 (O_1322,N_48607,N_49928);
xor UO_1323 (O_1323,N_49900,N_48918);
nand UO_1324 (O_1324,N_49557,N_48784);
or UO_1325 (O_1325,N_48368,N_48594);
or UO_1326 (O_1326,N_48183,N_48746);
nor UO_1327 (O_1327,N_49917,N_49420);
nand UO_1328 (O_1328,N_49037,N_48573);
and UO_1329 (O_1329,N_48637,N_49488);
nand UO_1330 (O_1330,N_49582,N_48192);
nor UO_1331 (O_1331,N_48012,N_49963);
xor UO_1332 (O_1332,N_49705,N_48606);
xor UO_1333 (O_1333,N_49718,N_48188);
nand UO_1334 (O_1334,N_49545,N_49994);
nand UO_1335 (O_1335,N_48961,N_49864);
or UO_1336 (O_1336,N_48405,N_49382);
xor UO_1337 (O_1337,N_49150,N_49179);
nor UO_1338 (O_1338,N_49781,N_49552);
and UO_1339 (O_1339,N_48649,N_48563);
nor UO_1340 (O_1340,N_49101,N_49608);
nor UO_1341 (O_1341,N_49148,N_48951);
nor UO_1342 (O_1342,N_49437,N_49026);
and UO_1343 (O_1343,N_48129,N_49132);
or UO_1344 (O_1344,N_49903,N_48291);
nand UO_1345 (O_1345,N_48518,N_49894);
nor UO_1346 (O_1346,N_49291,N_49421);
nand UO_1347 (O_1347,N_48621,N_48518);
nor UO_1348 (O_1348,N_48836,N_48984);
nor UO_1349 (O_1349,N_48811,N_48026);
nor UO_1350 (O_1350,N_48310,N_48468);
nand UO_1351 (O_1351,N_49949,N_49070);
xnor UO_1352 (O_1352,N_48842,N_48246);
nand UO_1353 (O_1353,N_48048,N_48476);
nor UO_1354 (O_1354,N_49164,N_48769);
nand UO_1355 (O_1355,N_49128,N_49615);
nor UO_1356 (O_1356,N_48019,N_49511);
nand UO_1357 (O_1357,N_49988,N_48534);
xor UO_1358 (O_1358,N_49239,N_48297);
or UO_1359 (O_1359,N_48946,N_49373);
or UO_1360 (O_1360,N_48541,N_48103);
nor UO_1361 (O_1361,N_48900,N_49747);
or UO_1362 (O_1362,N_48659,N_49942);
and UO_1363 (O_1363,N_48418,N_48912);
and UO_1364 (O_1364,N_49161,N_49972);
or UO_1365 (O_1365,N_49835,N_48140);
xor UO_1366 (O_1366,N_48020,N_48663);
xnor UO_1367 (O_1367,N_49932,N_49964);
or UO_1368 (O_1368,N_49504,N_49440);
or UO_1369 (O_1369,N_48069,N_49359);
xnor UO_1370 (O_1370,N_48720,N_49748);
xnor UO_1371 (O_1371,N_49565,N_49377);
nand UO_1372 (O_1372,N_49069,N_48742);
nand UO_1373 (O_1373,N_49210,N_48335);
and UO_1374 (O_1374,N_49898,N_49273);
xor UO_1375 (O_1375,N_48291,N_48916);
or UO_1376 (O_1376,N_49831,N_48680);
or UO_1377 (O_1377,N_48928,N_49068);
nand UO_1378 (O_1378,N_49286,N_49888);
xnor UO_1379 (O_1379,N_49367,N_49918);
nand UO_1380 (O_1380,N_48523,N_49311);
nand UO_1381 (O_1381,N_48174,N_48842);
or UO_1382 (O_1382,N_49461,N_48831);
and UO_1383 (O_1383,N_49651,N_48395);
nand UO_1384 (O_1384,N_49069,N_49770);
nand UO_1385 (O_1385,N_48032,N_48324);
and UO_1386 (O_1386,N_48440,N_48628);
and UO_1387 (O_1387,N_49749,N_49860);
or UO_1388 (O_1388,N_49276,N_48075);
or UO_1389 (O_1389,N_48306,N_49914);
nand UO_1390 (O_1390,N_49548,N_48711);
or UO_1391 (O_1391,N_48894,N_48029);
nor UO_1392 (O_1392,N_49353,N_48638);
or UO_1393 (O_1393,N_49244,N_48039);
xnor UO_1394 (O_1394,N_49827,N_49981);
nor UO_1395 (O_1395,N_49972,N_48383);
nand UO_1396 (O_1396,N_48869,N_49671);
nand UO_1397 (O_1397,N_48220,N_48624);
nand UO_1398 (O_1398,N_49056,N_49550);
xnor UO_1399 (O_1399,N_48686,N_48486);
nor UO_1400 (O_1400,N_49397,N_49546);
or UO_1401 (O_1401,N_49690,N_48900);
nor UO_1402 (O_1402,N_49131,N_49229);
xnor UO_1403 (O_1403,N_49123,N_49662);
xnor UO_1404 (O_1404,N_48869,N_48878);
nor UO_1405 (O_1405,N_48822,N_49873);
nand UO_1406 (O_1406,N_49545,N_49142);
or UO_1407 (O_1407,N_48905,N_48461);
nand UO_1408 (O_1408,N_49220,N_48051);
nand UO_1409 (O_1409,N_48455,N_49774);
nor UO_1410 (O_1410,N_49754,N_49771);
xor UO_1411 (O_1411,N_49140,N_49230);
nor UO_1412 (O_1412,N_49642,N_48643);
xnor UO_1413 (O_1413,N_48024,N_49435);
xor UO_1414 (O_1414,N_48193,N_48221);
or UO_1415 (O_1415,N_48365,N_49567);
nor UO_1416 (O_1416,N_48944,N_49248);
and UO_1417 (O_1417,N_49660,N_49563);
or UO_1418 (O_1418,N_49540,N_49911);
nand UO_1419 (O_1419,N_48742,N_48898);
nor UO_1420 (O_1420,N_49106,N_48428);
and UO_1421 (O_1421,N_48252,N_49557);
or UO_1422 (O_1422,N_48821,N_48259);
xnor UO_1423 (O_1423,N_48305,N_49736);
or UO_1424 (O_1424,N_48341,N_49748);
nor UO_1425 (O_1425,N_48844,N_49701);
or UO_1426 (O_1426,N_48761,N_48943);
and UO_1427 (O_1427,N_48760,N_48890);
and UO_1428 (O_1428,N_49233,N_49188);
xor UO_1429 (O_1429,N_49914,N_48830);
or UO_1430 (O_1430,N_48460,N_49804);
or UO_1431 (O_1431,N_49384,N_49908);
or UO_1432 (O_1432,N_49384,N_49653);
or UO_1433 (O_1433,N_49871,N_48776);
and UO_1434 (O_1434,N_49031,N_49102);
nor UO_1435 (O_1435,N_49186,N_48241);
nor UO_1436 (O_1436,N_49525,N_49362);
nand UO_1437 (O_1437,N_49447,N_48134);
nor UO_1438 (O_1438,N_49006,N_49361);
xor UO_1439 (O_1439,N_49974,N_49259);
and UO_1440 (O_1440,N_48357,N_48758);
or UO_1441 (O_1441,N_48326,N_49574);
nor UO_1442 (O_1442,N_49125,N_49755);
and UO_1443 (O_1443,N_48980,N_49351);
or UO_1444 (O_1444,N_48612,N_48750);
or UO_1445 (O_1445,N_49422,N_48001);
and UO_1446 (O_1446,N_49535,N_48071);
xor UO_1447 (O_1447,N_49441,N_48123);
or UO_1448 (O_1448,N_48365,N_49386);
xor UO_1449 (O_1449,N_49524,N_49314);
nor UO_1450 (O_1450,N_49028,N_48921);
xor UO_1451 (O_1451,N_49154,N_48088);
or UO_1452 (O_1452,N_48450,N_49623);
nor UO_1453 (O_1453,N_48603,N_48916);
nand UO_1454 (O_1454,N_48213,N_49313);
xnor UO_1455 (O_1455,N_49158,N_48096);
nand UO_1456 (O_1456,N_48357,N_49521);
or UO_1457 (O_1457,N_49358,N_49877);
xor UO_1458 (O_1458,N_48388,N_48871);
xor UO_1459 (O_1459,N_48680,N_49780);
and UO_1460 (O_1460,N_48425,N_48924);
or UO_1461 (O_1461,N_49195,N_48396);
nor UO_1462 (O_1462,N_49885,N_48458);
or UO_1463 (O_1463,N_48920,N_48864);
and UO_1464 (O_1464,N_48331,N_48395);
xnor UO_1465 (O_1465,N_49125,N_48376);
nand UO_1466 (O_1466,N_49905,N_49104);
and UO_1467 (O_1467,N_49110,N_48678);
xnor UO_1468 (O_1468,N_49543,N_49863);
xnor UO_1469 (O_1469,N_49152,N_48470);
and UO_1470 (O_1470,N_48559,N_48522);
nand UO_1471 (O_1471,N_48672,N_48415);
xor UO_1472 (O_1472,N_49621,N_48979);
nand UO_1473 (O_1473,N_48175,N_49252);
nor UO_1474 (O_1474,N_49811,N_48758);
nand UO_1475 (O_1475,N_48669,N_49635);
and UO_1476 (O_1476,N_48087,N_49819);
nor UO_1477 (O_1477,N_49425,N_48416);
xnor UO_1478 (O_1478,N_49351,N_49348);
or UO_1479 (O_1479,N_49965,N_48367);
nor UO_1480 (O_1480,N_49581,N_49218);
and UO_1481 (O_1481,N_48761,N_49995);
or UO_1482 (O_1482,N_48814,N_49536);
nand UO_1483 (O_1483,N_49232,N_48735);
and UO_1484 (O_1484,N_49862,N_48103);
or UO_1485 (O_1485,N_48918,N_49480);
nand UO_1486 (O_1486,N_48303,N_49366);
and UO_1487 (O_1487,N_48726,N_48365);
nor UO_1488 (O_1488,N_49623,N_49242);
nor UO_1489 (O_1489,N_49825,N_48057);
nor UO_1490 (O_1490,N_48160,N_48871);
nor UO_1491 (O_1491,N_49262,N_48470);
and UO_1492 (O_1492,N_48491,N_48849);
nand UO_1493 (O_1493,N_48713,N_48021);
nand UO_1494 (O_1494,N_49326,N_49671);
and UO_1495 (O_1495,N_49942,N_48131);
nor UO_1496 (O_1496,N_48688,N_48955);
nor UO_1497 (O_1497,N_48041,N_48395);
or UO_1498 (O_1498,N_49016,N_49907);
or UO_1499 (O_1499,N_49434,N_49031);
xnor UO_1500 (O_1500,N_49561,N_49229);
or UO_1501 (O_1501,N_49532,N_49707);
nor UO_1502 (O_1502,N_48259,N_48373);
xor UO_1503 (O_1503,N_49605,N_48901);
nor UO_1504 (O_1504,N_49031,N_48016);
nand UO_1505 (O_1505,N_48167,N_49966);
and UO_1506 (O_1506,N_49617,N_49331);
nor UO_1507 (O_1507,N_48429,N_48811);
and UO_1508 (O_1508,N_48057,N_49440);
and UO_1509 (O_1509,N_48175,N_49685);
and UO_1510 (O_1510,N_49271,N_48495);
nand UO_1511 (O_1511,N_48381,N_48727);
nor UO_1512 (O_1512,N_49278,N_49336);
nand UO_1513 (O_1513,N_49399,N_48154);
or UO_1514 (O_1514,N_49231,N_48480);
or UO_1515 (O_1515,N_49763,N_48897);
nand UO_1516 (O_1516,N_48232,N_48582);
nand UO_1517 (O_1517,N_48401,N_48530);
nand UO_1518 (O_1518,N_48248,N_48000);
nor UO_1519 (O_1519,N_48272,N_49275);
nand UO_1520 (O_1520,N_49886,N_49793);
or UO_1521 (O_1521,N_48504,N_49697);
and UO_1522 (O_1522,N_49951,N_48351);
or UO_1523 (O_1523,N_49959,N_48055);
nand UO_1524 (O_1524,N_48012,N_48000);
and UO_1525 (O_1525,N_48120,N_48543);
nand UO_1526 (O_1526,N_49353,N_48804);
nor UO_1527 (O_1527,N_48839,N_48966);
and UO_1528 (O_1528,N_49644,N_49654);
nor UO_1529 (O_1529,N_48001,N_49065);
and UO_1530 (O_1530,N_49646,N_49200);
and UO_1531 (O_1531,N_48492,N_48655);
xnor UO_1532 (O_1532,N_49639,N_49737);
and UO_1533 (O_1533,N_49596,N_48463);
nand UO_1534 (O_1534,N_49398,N_49818);
nand UO_1535 (O_1535,N_49987,N_48687);
or UO_1536 (O_1536,N_49438,N_49331);
or UO_1537 (O_1537,N_48544,N_49239);
nand UO_1538 (O_1538,N_48414,N_48991);
and UO_1539 (O_1539,N_49532,N_49381);
or UO_1540 (O_1540,N_48303,N_49657);
xor UO_1541 (O_1541,N_49121,N_48836);
and UO_1542 (O_1542,N_48247,N_48422);
and UO_1543 (O_1543,N_49685,N_48319);
or UO_1544 (O_1544,N_49340,N_48985);
nor UO_1545 (O_1545,N_48280,N_49000);
xor UO_1546 (O_1546,N_48234,N_49694);
or UO_1547 (O_1547,N_48279,N_49021);
nor UO_1548 (O_1548,N_49404,N_49029);
nand UO_1549 (O_1549,N_48743,N_48390);
or UO_1550 (O_1550,N_48343,N_48066);
nor UO_1551 (O_1551,N_49238,N_49138);
nor UO_1552 (O_1552,N_48707,N_48433);
nand UO_1553 (O_1553,N_48799,N_49583);
xnor UO_1554 (O_1554,N_49232,N_49268);
xnor UO_1555 (O_1555,N_48688,N_49007);
or UO_1556 (O_1556,N_49225,N_48034);
or UO_1557 (O_1557,N_49777,N_48806);
nor UO_1558 (O_1558,N_48610,N_48537);
xnor UO_1559 (O_1559,N_48594,N_48801);
xnor UO_1560 (O_1560,N_49734,N_48933);
xor UO_1561 (O_1561,N_48721,N_48868);
nor UO_1562 (O_1562,N_49377,N_49363);
nand UO_1563 (O_1563,N_49522,N_49894);
and UO_1564 (O_1564,N_48749,N_49430);
xnor UO_1565 (O_1565,N_48312,N_49256);
and UO_1566 (O_1566,N_49657,N_49587);
or UO_1567 (O_1567,N_48262,N_48689);
nand UO_1568 (O_1568,N_49758,N_48439);
or UO_1569 (O_1569,N_48719,N_49842);
and UO_1570 (O_1570,N_48126,N_49896);
and UO_1571 (O_1571,N_49713,N_48104);
or UO_1572 (O_1572,N_49051,N_48811);
nand UO_1573 (O_1573,N_48886,N_49312);
or UO_1574 (O_1574,N_49767,N_49676);
xor UO_1575 (O_1575,N_49800,N_48257);
nor UO_1576 (O_1576,N_49909,N_48399);
and UO_1577 (O_1577,N_48792,N_48965);
nand UO_1578 (O_1578,N_48499,N_48820);
nor UO_1579 (O_1579,N_48384,N_49163);
nor UO_1580 (O_1580,N_48945,N_48355);
xor UO_1581 (O_1581,N_49277,N_48920);
and UO_1582 (O_1582,N_48841,N_48455);
nand UO_1583 (O_1583,N_48626,N_48851);
nand UO_1584 (O_1584,N_49585,N_48041);
xor UO_1585 (O_1585,N_49688,N_48211);
nand UO_1586 (O_1586,N_49738,N_48778);
xnor UO_1587 (O_1587,N_49620,N_48500);
and UO_1588 (O_1588,N_48697,N_49542);
and UO_1589 (O_1589,N_48764,N_48258);
xor UO_1590 (O_1590,N_49604,N_48513);
or UO_1591 (O_1591,N_49742,N_48386);
xnor UO_1592 (O_1592,N_49982,N_48750);
or UO_1593 (O_1593,N_49089,N_49330);
nand UO_1594 (O_1594,N_48017,N_48203);
nand UO_1595 (O_1595,N_48868,N_48475);
nor UO_1596 (O_1596,N_49610,N_48535);
nand UO_1597 (O_1597,N_49465,N_48556);
and UO_1598 (O_1598,N_49598,N_49237);
nor UO_1599 (O_1599,N_48191,N_48711);
or UO_1600 (O_1600,N_48051,N_49698);
xnor UO_1601 (O_1601,N_49105,N_49194);
or UO_1602 (O_1602,N_48660,N_48747);
nor UO_1603 (O_1603,N_49855,N_49335);
xor UO_1604 (O_1604,N_48632,N_48683);
or UO_1605 (O_1605,N_48919,N_49620);
or UO_1606 (O_1606,N_49406,N_48939);
nand UO_1607 (O_1607,N_48845,N_49625);
or UO_1608 (O_1608,N_48803,N_48024);
and UO_1609 (O_1609,N_48970,N_48381);
and UO_1610 (O_1610,N_49123,N_48733);
nand UO_1611 (O_1611,N_48735,N_48066);
or UO_1612 (O_1612,N_49478,N_49887);
xnor UO_1613 (O_1613,N_48898,N_49210);
nand UO_1614 (O_1614,N_49790,N_48065);
xor UO_1615 (O_1615,N_48373,N_49461);
xor UO_1616 (O_1616,N_49000,N_48250);
and UO_1617 (O_1617,N_49567,N_49929);
xnor UO_1618 (O_1618,N_49507,N_49266);
nand UO_1619 (O_1619,N_48108,N_49158);
xnor UO_1620 (O_1620,N_48993,N_48885);
nand UO_1621 (O_1621,N_49590,N_48520);
nand UO_1622 (O_1622,N_48264,N_49203);
and UO_1623 (O_1623,N_49356,N_48924);
nor UO_1624 (O_1624,N_49900,N_49238);
xnor UO_1625 (O_1625,N_49224,N_49135);
and UO_1626 (O_1626,N_49245,N_49801);
and UO_1627 (O_1627,N_48779,N_48923);
or UO_1628 (O_1628,N_48549,N_48515);
xor UO_1629 (O_1629,N_49779,N_49089);
nor UO_1630 (O_1630,N_48491,N_49332);
nand UO_1631 (O_1631,N_48563,N_49517);
nand UO_1632 (O_1632,N_49702,N_49687);
xnor UO_1633 (O_1633,N_49400,N_48727);
and UO_1634 (O_1634,N_49494,N_48401);
and UO_1635 (O_1635,N_49227,N_49981);
and UO_1636 (O_1636,N_49830,N_48083);
xor UO_1637 (O_1637,N_48245,N_49536);
nand UO_1638 (O_1638,N_48148,N_48726);
nor UO_1639 (O_1639,N_49246,N_48182);
nor UO_1640 (O_1640,N_48064,N_49042);
nor UO_1641 (O_1641,N_48691,N_49563);
or UO_1642 (O_1642,N_49564,N_48582);
and UO_1643 (O_1643,N_49156,N_49727);
nor UO_1644 (O_1644,N_49533,N_49485);
or UO_1645 (O_1645,N_48128,N_48075);
nor UO_1646 (O_1646,N_48210,N_49173);
nand UO_1647 (O_1647,N_49655,N_48059);
or UO_1648 (O_1648,N_49681,N_49839);
xor UO_1649 (O_1649,N_49817,N_48932);
and UO_1650 (O_1650,N_49546,N_49673);
and UO_1651 (O_1651,N_49376,N_48486);
xnor UO_1652 (O_1652,N_49042,N_49810);
and UO_1653 (O_1653,N_48991,N_49252);
or UO_1654 (O_1654,N_48606,N_49340);
nand UO_1655 (O_1655,N_49142,N_49252);
and UO_1656 (O_1656,N_48565,N_49265);
nand UO_1657 (O_1657,N_48926,N_48521);
nor UO_1658 (O_1658,N_48939,N_49230);
and UO_1659 (O_1659,N_48516,N_48773);
nor UO_1660 (O_1660,N_49076,N_49355);
nand UO_1661 (O_1661,N_48271,N_48427);
or UO_1662 (O_1662,N_48524,N_48101);
and UO_1663 (O_1663,N_49705,N_48970);
nor UO_1664 (O_1664,N_49949,N_48841);
nand UO_1665 (O_1665,N_49510,N_48847);
xor UO_1666 (O_1666,N_48564,N_49437);
nand UO_1667 (O_1667,N_49116,N_49208);
nand UO_1668 (O_1668,N_48296,N_48674);
and UO_1669 (O_1669,N_48428,N_49025);
nand UO_1670 (O_1670,N_48429,N_49105);
nand UO_1671 (O_1671,N_48938,N_49814);
or UO_1672 (O_1672,N_48458,N_49152);
or UO_1673 (O_1673,N_49927,N_49849);
nand UO_1674 (O_1674,N_49070,N_49227);
and UO_1675 (O_1675,N_49861,N_48056);
or UO_1676 (O_1676,N_49755,N_48877);
nand UO_1677 (O_1677,N_48789,N_48838);
xnor UO_1678 (O_1678,N_49460,N_49768);
nor UO_1679 (O_1679,N_49617,N_48224);
or UO_1680 (O_1680,N_49853,N_49404);
and UO_1681 (O_1681,N_48010,N_48095);
nor UO_1682 (O_1682,N_49594,N_49434);
and UO_1683 (O_1683,N_48036,N_49570);
nor UO_1684 (O_1684,N_49139,N_48684);
nor UO_1685 (O_1685,N_49925,N_49363);
or UO_1686 (O_1686,N_48653,N_48085);
xnor UO_1687 (O_1687,N_49571,N_49136);
and UO_1688 (O_1688,N_49880,N_49703);
or UO_1689 (O_1689,N_48528,N_49177);
xor UO_1690 (O_1690,N_48505,N_49272);
nor UO_1691 (O_1691,N_48643,N_49420);
nor UO_1692 (O_1692,N_49242,N_48629);
and UO_1693 (O_1693,N_48738,N_49206);
nand UO_1694 (O_1694,N_48102,N_49455);
xor UO_1695 (O_1695,N_49243,N_49335);
nor UO_1696 (O_1696,N_49522,N_49663);
xor UO_1697 (O_1697,N_48870,N_48741);
xnor UO_1698 (O_1698,N_49863,N_48765);
or UO_1699 (O_1699,N_49602,N_48433);
nand UO_1700 (O_1700,N_49183,N_48061);
or UO_1701 (O_1701,N_48468,N_49734);
or UO_1702 (O_1702,N_49919,N_49285);
nor UO_1703 (O_1703,N_48298,N_49932);
and UO_1704 (O_1704,N_49903,N_49630);
nor UO_1705 (O_1705,N_48956,N_48208);
or UO_1706 (O_1706,N_48949,N_49869);
nor UO_1707 (O_1707,N_49565,N_48173);
xor UO_1708 (O_1708,N_48052,N_49893);
nand UO_1709 (O_1709,N_48874,N_48701);
and UO_1710 (O_1710,N_49258,N_48922);
or UO_1711 (O_1711,N_48890,N_48449);
or UO_1712 (O_1712,N_49915,N_49740);
nor UO_1713 (O_1713,N_49150,N_48603);
nor UO_1714 (O_1714,N_49989,N_48762);
or UO_1715 (O_1715,N_49141,N_48591);
nor UO_1716 (O_1716,N_49108,N_48925);
or UO_1717 (O_1717,N_48146,N_49382);
xor UO_1718 (O_1718,N_49582,N_49098);
nor UO_1719 (O_1719,N_48055,N_48390);
xnor UO_1720 (O_1720,N_49320,N_48510);
xnor UO_1721 (O_1721,N_48261,N_48766);
nand UO_1722 (O_1722,N_48400,N_49002);
nor UO_1723 (O_1723,N_49005,N_49635);
nor UO_1724 (O_1724,N_49836,N_49626);
nor UO_1725 (O_1725,N_49097,N_49768);
xnor UO_1726 (O_1726,N_48599,N_49016);
nor UO_1727 (O_1727,N_49204,N_48194);
and UO_1728 (O_1728,N_49340,N_48143);
and UO_1729 (O_1729,N_48017,N_49509);
nor UO_1730 (O_1730,N_49370,N_48522);
xnor UO_1731 (O_1731,N_48395,N_48945);
nor UO_1732 (O_1732,N_49005,N_49855);
and UO_1733 (O_1733,N_48567,N_48968);
nand UO_1734 (O_1734,N_49867,N_48700);
nor UO_1735 (O_1735,N_49701,N_49009);
nand UO_1736 (O_1736,N_48292,N_49065);
nor UO_1737 (O_1737,N_49254,N_49256);
or UO_1738 (O_1738,N_49811,N_49312);
nor UO_1739 (O_1739,N_48925,N_48124);
xor UO_1740 (O_1740,N_48279,N_48406);
nand UO_1741 (O_1741,N_49104,N_49517);
xnor UO_1742 (O_1742,N_49664,N_49061);
or UO_1743 (O_1743,N_49189,N_49981);
nand UO_1744 (O_1744,N_49348,N_49942);
nor UO_1745 (O_1745,N_49599,N_48533);
nor UO_1746 (O_1746,N_49230,N_49869);
nor UO_1747 (O_1747,N_49468,N_49347);
and UO_1748 (O_1748,N_48880,N_48553);
and UO_1749 (O_1749,N_49001,N_48865);
xnor UO_1750 (O_1750,N_48739,N_48090);
nand UO_1751 (O_1751,N_48281,N_48463);
nand UO_1752 (O_1752,N_49647,N_49007);
and UO_1753 (O_1753,N_49404,N_49539);
xnor UO_1754 (O_1754,N_49534,N_49142);
and UO_1755 (O_1755,N_48876,N_49348);
xnor UO_1756 (O_1756,N_49619,N_48466);
and UO_1757 (O_1757,N_48171,N_49191);
nand UO_1758 (O_1758,N_49352,N_48943);
xnor UO_1759 (O_1759,N_49284,N_48043);
or UO_1760 (O_1760,N_48284,N_48075);
xor UO_1761 (O_1761,N_49710,N_48579);
nand UO_1762 (O_1762,N_49342,N_49365);
nor UO_1763 (O_1763,N_48295,N_49763);
nand UO_1764 (O_1764,N_48117,N_48732);
and UO_1765 (O_1765,N_48882,N_49936);
xor UO_1766 (O_1766,N_49005,N_49364);
xor UO_1767 (O_1767,N_48065,N_49272);
and UO_1768 (O_1768,N_48444,N_49929);
or UO_1769 (O_1769,N_49564,N_49192);
xnor UO_1770 (O_1770,N_49723,N_48967);
xor UO_1771 (O_1771,N_49043,N_49010);
nand UO_1772 (O_1772,N_49180,N_48045);
xnor UO_1773 (O_1773,N_48266,N_49650);
or UO_1774 (O_1774,N_49923,N_48960);
nand UO_1775 (O_1775,N_49594,N_48682);
xnor UO_1776 (O_1776,N_48767,N_49951);
or UO_1777 (O_1777,N_48625,N_48992);
and UO_1778 (O_1778,N_48677,N_48718);
and UO_1779 (O_1779,N_48115,N_48952);
or UO_1780 (O_1780,N_49927,N_48181);
and UO_1781 (O_1781,N_48724,N_48149);
and UO_1782 (O_1782,N_48321,N_49227);
xor UO_1783 (O_1783,N_49443,N_48024);
nand UO_1784 (O_1784,N_49834,N_49266);
nor UO_1785 (O_1785,N_49892,N_49477);
nor UO_1786 (O_1786,N_48092,N_49559);
xnor UO_1787 (O_1787,N_49612,N_49778);
and UO_1788 (O_1788,N_49752,N_48519);
xnor UO_1789 (O_1789,N_48451,N_49025);
and UO_1790 (O_1790,N_49787,N_48295);
xnor UO_1791 (O_1791,N_48000,N_49504);
nand UO_1792 (O_1792,N_49737,N_48785);
nor UO_1793 (O_1793,N_48011,N_48739);
or UO_1794 (O_1794,N_49398,N_48406);
and UO_1795 (O_1795,N_48949,N_49467);
nand UO_1796 (O_1796,N_49725,N_48007);
and UO_1797 (O_1797,N_49211,N_49624);
or UO_1798 (O_1798,N_49311,N_49988);
nand UO_1799 (O_1799,N_48289,N_48216);
nand UO_1800 (O_1800,N_48303,N_48048);
and UO_1801 (O_1801,N_48023,N_49383);
xnor UO_1802 (O_1802,N_49333,N_49493);
nand UO_1803 (O_1803,N_48303,N_48639);
xor UO_1804 (O_1804,N_49651,N_48925);
and UO_1805 (O_1805,N_48210,N_49454);
and UO_1806 (O_1806,N_48545,N_48757);
and UO_1807 (O_1807,N_48366,N_48228);
or UO_1808 (O_1808,N_48989,N_49373);
xnor UO_1809 (O_1809,N_49896,N_48100);
nand UO_1810 (O_1810,N_49452,N_48649);
and UO_1811 (O_1811,N_49431,N_49697);
xnor UO_1812 (O_1812,N_49283,N_49694);
xor UO_1813 (O_1813,N_49325,N_48392);
nor UO_1814 (O_1814,N_48549,N_49195);
xnor UO_1815 (O_1815,N_49495,N_49050);
xnor UO_1816 (O_1816,N_48384,N_49632);
or UO_1817 (O_1817,N_48501,N_48942);
and UO_1818 (O_1818,N_48720,N_49964);
nand UO_1819 (O_1819,N_48723,N_49798);
nor UO_1820 (O_1820,N_48776,N_48552);
nand UO_1821 (O_1821,N_49176,N_48143);
xor UO_1822 (O_1822,N_49320,N_48554);
and UO_1823 (O_1823,N_49624,N_48239);
and UO_1824 (O_1824,N_48801,N_48896);
nor UO_1825 (O_1825,N_49997,N_49910);
xnor UO_1826 (O_1826,N_49869,N_48042);
nor UO_1827 (O_1827,N_48440,N_48124);
and UO_1828 (O_1828,N_49989,N_49924);
or UO_1829 (O_1829,N_48672,N_48297);
nor UO_1830 (O_1830,N_49850,N_49935);
xnor UO_1831 (O_1831,N_48654,N_49407);
nand UO_1832 (O_1832,N_48107,N_48596);
and UO_1833 (O_1833,N_48249,N_49808);
or UO_1834 (O_1834,N_49174,N_49863);
xor UO_1835 (O_1835,N_48825,N_48628);
nor UO_1836 (O_1836,N_49246,N_49344);
xnor UO_1837 (O_1837,N_48313,N_49971);
or UO_1838 (O_1838,N_48783,N_48316);
nand UO_1839 (O_1839,N_49701,N_49404);
or UO_1840 (O_1840,N_48664,N_48227);
nand UO_1841 (O_1841,N_49061,N_49711);
xor UO_1842 (O_1842,N_49446,N_49459);
nor UO_1843 (O_1843,N_48412,N_48204);
and UO_1844 (O_1844,N_48219,N_49306);
or UO_1845 (O_1845,N_48318,N_49394);
or UO_1846 (O_1846,N_49882,N_49250);
nand UO_1847 (O_1847,N_48826,N_49195);
nor UO_1848 (O_1848,N_49105,N_49098);
and UO_1849 (O_1849,N_48054,N_48827);
nor UO_1850 (O_1850,N_49479,N_49436);
nand UO_1851 (O_1851,N_49047,N_49418);
nand UO_1852 (O_1852,N_48492,N_49771);
or UO_1853 (O_1853,N_48055,N_48981);
nand UO_1854 (O_1854,N_49838,N_49056);
or UO_1855 (O_1855,N_48461,N_48376);
nor UO_1856 (O_1856,N_48573,N_48349);
and UO_1857 (O_1857,N_48512,N_48016);
nand UO_1858 (O_1858,N_49690,N_48902);
xnor UO_1859 (O_1859,N_48015,N_48244);
or UO_1860 (O_1860,N_48410,N_49102);
or UO_1861 (O_1861,N_49511,N_49394);
or UO_1862 (O_1862,N_49833,N_48793);
or UO_1863 (O_1863,N_48353,N_48557);
nand UO_1864 (O_1864,N_48990,N_49670);
nor UO_1865 (O_1865,N_49689,N_49859);
nand UO_1866 (O_1866,N_48500,N_48343);
or UO_1867 (O_1867,N_48031,N_49860);
nor UO_1868 (O_1868,N_49691,N_48356);
nor UO_1869 (O_1869,N_48930,N_48102);
and UO_1870 (O_1870,N_48992,N_48153);
xnor UO_1871 (O_1871,N_48014,N_48334);
nor UO_1872 (O_1872,N_49579,N_48853);
or UO_1873 (O_1873,N_48772,N_49176);
nand UO_1874 (O_1874,N_49996,N_48501);
nand UO_1875 (O_1875,N_49232,N_48460);
or UO_1876 (O_1876,N_49480,N_48037);
or UO_1877 (O_1877,N_49158,N_49151);
xnor UO_1878 (O_1878,N_49976,N_49112);
nand UO_1879 (O_1879,N_48107,N_48849);
nand UO_1880 (O_1880,N_49271,N_48729);
xnor UO_1881 (O_1881,N_48218,N_48259);
and UO_1882 (O_1882,N_48376,N_48031);
xor UO_1883 (O_1883,N_48865,N_49238);
xor UO_1884 (O_1884,N_49027,N_48098);
nand UO_1885 (O_1885,N_48712,N_49734);
nor UO_1886 (O_1886,N_49053,N_49760);
and UO_1887 (O_1887,N_49604,N_48369);
or UO_1888 (O_1888,N_49518,N_49308);
nor UO_1889 (O_1889,N_48655,N_49869);
nand UO_1890 (O_1890,N_48806,N_48430);
xnor UO_1891 (O_1891,N_48290,N_49136);
and UO_1892 (O_1892,N_48213,N_49209);
xnor UO_1893 (O_1893,N_49142,N_48860);
nor UO_1894 (O_1894,N_48623,N_48618);
and UO_1895 (O_1895,N_49471,N_49220);
nand UO_1896 (O_1896,N_48578,N_49051);
xor UO_1897 (O_1897,N_48063,N_49095);
and UO_1898 (O_1898,N_49887,N_48639);
or UO_1899 (O_1899,N_48553,N_48722);
and UO_1900 (O_1900,N_49409,N_48412);
nand UO_1901 (O_1901,N_48176,N_48057);
nand UO_1902 (O_1902,N_49448,N_48285);
and UO_1903 (O_1903,N_49264,N_49970);
and UO_1904 (O_1904,N_48916,N_49338);
nor UO_1905 (O_1905,N_48407,N_48976);
and UO_1906 (O_1906,N_48733,N_49035);
nor UO_1907 (O_1907,N_48050,N_48828);
nand UO_1908 (O_1908,N_49031,N_48798);
nand UO_1909 (O_1909,N_48514,N_48287);
nand UO_1910 (O_1910,N_49679,N_48773);
nor UO_1911 (O_1911,N_49821,N_48087);
or UO_1912 (O_1912,N_48197,N_49790);
nand UO_1913 (O_1913,N_49377,N_49811);
and UO_1914 (O_1914,N_48796,N_49952);
xnor UO_1915 (O_1915,N_48242,N_48775);
xnor UO_1916 (O_1916,N_48573,N_48094);
nor UO_1917 (O_1917,N_48184,N_49592);
xor UO_1918 (O_1918,N_48104,N_49416);
and UO_1919 (O_1919,N_49264,N_48556);
nand UO_1920 (O_1920,N_49375,N_48109);
nor UO_1921 (O_1921,N_48222,N_48326);
or UO_1922 (O_1922,N_48992,N_48423);
and UO_1923 (O_1923,N_49174,N_48891);
and UO_1924 (O_1924,N_48313,N_48578);
xnor UO_1925 (O_1925,N_48140,N_49918);
nor UO_1926 (O_1926,N_49430,N_49796);
and UO_1927 (O_1927,N_49833,N_48087);
xnor UO_1928 (O_1928,N_48310,N_49714);
xnor UO_1929 (O_1929,N_49495,N_48395);
xor UO_1930 (O_1930,N_48032,N_49919);
xnor UO_1931 (O_1931,N_49833,N_48968);
and UO_1932 (O_1932,N_48971,N_48980);
and UO_1933 (O_1933,N_48733,N_49763);
nor UO_1934 (O_1934,N_49989,N_48203);
or UO_1935 (O_1935,N_48049,N_48370);
nand UO_1936 (O_1936,N_48966,N_48750);
nand UO_1937 (O_1937,N_49553,N_48061);
or UO_1938 (O_1938,N_48455,N_49922);
or UO_1939 (O_1939,N_49942,N_48996);
and UO_1940 (O_1940,N_49244,N_48283);
nor UO_1941 (O_1941,N_49033,N_49884);
nand UO_1942 (O_1942,N_49358,N_49031);
nand UO_1943 (O_1943,N_49873,N_48765);
nand UO_1944 (O_1944,N_49752,N_48007);
nor UO_1945 (O_1945,N_48411,N_49147);
nor UO_1946 (O_1946,N_49291,N_48419);
or UO_1947 (O_1947,N_48246,N_49081);
nor UO_1948 (O_1948,N_49094,N_48218);
nor UO_1949 (O_1949,N_49409,N_49170);
nor UO_1950 (O_1950,N_48561,N_49412);
xnor UO_1951 (O_1951,N_49608,N_49856);
and UO_1952 (O_1952,N_48800,N_49982);
nor UO_1953 (O_1953,N_48955,N_48339);
nand UO_1954 (O_1954,N_48213,N_48285);
and UO_1955 (O_1955,N_49048,N_48177);
and UO_1956 (O_1956,N_49702,N_49784);
and UO_1957 (O_1957,N_49104,N_49202);
xor UO_1958 (O_1958,N_48011,N_49333);
nor UO_1959 (O_1959,N_48744,N_49295);
xor UO_1960 (O_1960,N_48965,N_48009);
and UO_1961 (O_1961,N_49703,N_49732);
or UO_1962 (O_1962,N_48481,N_49543);
nor UO_1963 (O_1963,N_49168,N_49439);
nor UO_1964 (O_1964,N_49257,N_48329);
nand UO_1965 (O_1965,N_48056,N_49234);
nor UO_1966 (O_1966,N_48006,N_49731);
nor UO_1967 (O_1967,N_49211,N_48998);
and UO_1968 (O_1968,N_48101,N_49748);
and UO_1969 (O_1969,N_49031,N_48646);
nand UO_1970 (O_1970,N_48725,N_48123);
or UO_1971 (O_1971,N_48170,N_49727);
or UO_1972 (O_1972,N_49389,N_48676);
or UO_1973 (O_1973,N_48217,N_49342);
and UO_1974 (O_1974,N_49243,N_49122);
xnor UO_1975 (O_1975,N_49919,N_49543);
nor UO_1976 (O_1976,N_49992,N_49736);
or UO_1977 (O_1977,N_48470,N_49878);
nand UO_1978 (O_1978,N_49225,N_49437);
nand UO_1979 (O_1979,N_49534,N_48731);
and UO_1980 (O_1980,N_48429,N_48029);
or UO_1981 (O_1981,N_49148,N_49182);
nor UO_1982 (O_1982,N_49490,N_49859);
or UO_1983 (O_1983,N_49131,N_48639);
or UO_1984 (O_1984,N_48928,N_48948);
nand UO_1985 (O_1985,N_49226,N_48335);
nand UO_1986 (O_1986,N_48289,N_49314);
xnor UO_1987 (O_1987,N_49021,N_49050);
nor UO_1988 (O_1988,N_49227,N_48553);
and UO_1989 (O_1989,N_48281,N_48075);
or UO_1990 (O_1990,N_48926,N_49986);
and UO_1991 (O_1991,N_48036,N_48979);
nor UO_1992 (O_1992,N_48289,N_49089);
or UO_1993 (O_1993,N_48233,N_48466);
or UO_1994 (O_1994,N_48707,N_49482);
and UO_1995 (O_1995,N_48885,N_48642);
and UO_1996 (O_1996,N_49011,N_49665);
nor UO_1997 (O_1997,N_48458,N_49133);
nor UO_1998 (O_1998,N_48254,N_49723);
nor UO_1999 (O_1999,N_48804,N_48582);
nor UO_2000 (O_2000,N_49545,N_48906);
or UO_2001 (O_2001,N_49942,N_48979);
or UO_2002 (O_2002,N_49468,N_48540);
or UO_2003 (O_2003,N_48267,N_48114);
nand UO_2004 (O_2004,N_49281,N_48025);
or UO_2005 (O_2005,N_49792,N_49213);
nand UO_2006 (O_2006,N_48867,N_49067);
nand UO_2007 (O_2007,N_48674,N_49736);
or UO_2008 (O_2008,N_48277,N_48972);
nor UO_2009 (O_2009,N_48795,N_49388);
xor UO_2010 (O_2010,N_48488,N_49919);
xnor UO_2011 (O_2011,N_48065,N_49705);
and UO_2012 (O_2012,N_49311,N_49352);
xnor UO_2013 (O_2013,N_49702,N_49139);
and UO_2014 (O_2014,N_49518,N_48328);
or UO_2015 (O_2015,N_48641,N_49124);
or UO_2016 (O_2016,N_48744,N_49608);
nor UO_2017 (O_2017,N_48153,N_48470);
nand UO_2018 (O_2018,N_49901,N_48005);
and UO_2019 (O_2019,N_48059,N_49821);
and UO_2020 (O_2020,N_49504,N_49935);
nand UO_2021 (O_2021,N_49107,N_49054);
or UO_2022 (O_2022,N_48942,N_48013);
and UO_2023 (O_2023,N_49556,N_48743);
nand UO_2024 (O_2024,N_49717,N_48947);
nand UO_2025 (O_2025,N_48148,N_49181);
and UO_2026 (O_2026,N_48655,N_48480);
nand UO_2027 (O_2027,N_48151,N_48900);
nand UO_2028 (O_2028,N_49689,N_48206);
nand UO_2029 (O_2029,N_49285,N_48830);
nor UO_2030 (O_2030,N_49420,N_49640);
or UO_2031 (O_2031,N_49010,N_48855);
nor UO_2032 (O_2032,N_48514,N_48719);
or UO_2033 (O_2033,N_48282,N_48570);
nand UO_2034 (O_2034,N_48125,N_48168);
or UO_2035 (O_2035,N_49808,N_48198);
or UO_2036 (O_2036,N_49838,N_48420);
nor UO_2037 (O_2037,N_48859,N_48215);
and UO_2038 (O_2038,N_49384,N_48045);
or UO_2039 (O_2039,N_49425,N_49661);
nor UO_2040 (O_2040,N_49759,N_48870);
or UO_2041 (O_2041,N_48284,N_48484);
and UO_2042 (O_2042,N_48460,N_49299);
xnor UO_2043 (O_2043,N_48164,N_49677);
xnor UO_2044 (O_2044,N_48034,N_49489);
or UO_2045 (O_2045,N_49158,N_49164);
or UO_2046 (O_2046,N_49537,N_49752);
or UO_2047 (O_2047,N_48693,N_48627);
or UO_2048 (O_2048,N_48832,N_48050);
xor UO_2049 (O_2049,N_49837,N_49140);
nor UO_2050 (O_2050,N_48007,N_48448);
and UO_2051 (O_2051,N_48746,N_48934);
nand UO_2052 (O_2052,N_49836,N_49253);
xor UO_2053 (O_2053,N_49268,N_49734);
nor UO_2054 (O_2054,N_48097,N_48231);
nand UO_2055 (O_2055,N_48541,N_49526);
nor UO_2056 (O_2056,N_49575,N_49271);
and UO_2057 (O_2057,N_48965,N_49653);
and UO_2058 (O_2058,N_48442,N_49607);
and UO_2059 (O_2059,N_49693,N_48079);
or UO_2060 (O_2060,N_48041,N_48163);
and UO_2061 (O_2061,N_48819,N_48226);
nor UO_2062 (O_2062,N_48188,N_49443);
nand UO_2063 (O_2063,N_48774,N_49099);
nor UO_2064 (O_2064,N_48394,N_49443);
or UO_2065 (O_2065,N_48518,N_49492);
nand UO_2066 (O_2066,N_48737,N_48740);
xnor UO_2067 (O_2067,N_48607,N_49484);
and UO_2068 (O_2068,N_49702,N_48842);
or UO_2069 (O_2069,N_48017,N_48942);
nor UO_2070 (O_2070,N_49456,N_49828);
xnor UO_2071 (O_2071,N_48233,N_48048);
xnor UO_2072 (O_2072,N_49992,N_49751);
or UO_2073 (O_2073,N_49053,N_49761);
and UO_2074 (O_2074,N_48645,N_48431);
and UO_2075 (O_2075,N_49031,N_49025);
or UO_2076 (O_2076,N_49676,N_48617);
nand UO_2077 (O_2077,N_49491,N_48711);
and UO_2078 (O_2078,N_48000,N_48592);
xor UO_2079 (O_2079,N_48243,N_49291);
or UO_2080 (O_2080,N_49092,N_49093);
nor UO_2081 (O_2081,N_48425,N_48910);
or UO_2082 (O_2082,N_49526,N_48948);
and UO_2083 (O_2083,N_49389,N_49078);
xor UO_2084 (O_2084,N_48635,N_48720);
nor UO_2085 (O_2085,N_48601,N_48913);
and UO_2086 (O_2086,N_49101,N_48693);
nor UO_2087 (O_2087,N_49820,N_49380);
nand UO_2088 (O_2088,N_48604,N_48299);
or UO_2089 (O_2089,N_48922,N_48597);
nor UO_2090 (O_2090,N_49106,N_48427);
nand UO_2091 (O_2091,N_48531,N_48508);
and UO_2092 (O_2092,N_48159,N_48632);
xor UO_2093 (O_2093,N_49990,N_48953);
or UO_2094 (O_2094,N_49639,N_48506);
xor UO_2095 (O_2095,N_48720,N_48992);
nor UO_2096 (O_2096,N_48903,N_49485);
xnor UO_2097 (O_2097,N_48072,N_48592);
and UO_2098 (O_2098,N_49980,N_48521);
or UO_2099 (O_2099,N_49180,N_48093);
nor UO_2100 (O_2100,N_48482,N_48904);
or UO_2101 (O_2101,N_49599,N_48687);
or UO_2102 (O_2102,N_48564,N_49633);
nand UO_2103 (O_2103,N_48184,N_49665);
nand UO_2104 (O_2104,N_48823,N_48143);
or UO_2105 (O_2105,N_49695,N_49440);
xnor UO_2106 (O_2106,N_49716,N_48540);
and UO_2107 (O_2107,N_49417,N_48684);
and UO_2108 (O_2108,N_48494,N_49189);
xor UO_2109 (O_2109,N_49088,N_49940);
and UO_2110 (O_2110,N_49482,N_49742);
xor UO_2111 (O_2111,N_49292,N_49557);
and UO_2112 (O_2112,N_49611,N_49502);
nand UO_2113 (O_2113,N_48161,N_49121);
and UO_2114 (O_2114,N_49444,N_48108);
and UO_2115 (O_2115,N_49317,N_49719);
and UO_2116 (O_2116,N_48846,N_49645);
nor UO_2117 (O_2117,N_48270,N_48936);
nor UO_2118 (O_2118,N_48663,N_48824);
or UO_2119 (O_2119,N_48088,N_49236);
nor UO_2120 (O_2120,N_49197,N_48749);
or UO_2121 (O_2121,N_49880,N_49072);
nor UO_2122 (O_2122,N_48721,N_49427);
or UO_2123 (O_2123,N_48478,N_48483);
nor UO_2124 (O_2124,N_48799,N_49808);
xor UO_2125 (O_2125,N_48944,N_48146);
nor UO_2126 (O_2126,N_48468,N_48734);
or UO_2127 (O_2127,N_49786,N_48566);
xor UO_2128 (O_2128,N_48893,N_48667);
nand UO_2129 (O_2129,N_48676,N_48509);
nor UO_2130 (O_2130,N_49814,N_49338);
xnor UO_2131 (O_2131,N_49262,N_48389);
nor UO_2132 (O_2132,N_48565,N_49035);
and UO_2133 (O_2133,N_48398,N_48301);
nand UO_2134 (O_2134,N_49898,N_48694);
xor UO_2135 (O_2135,N_48225,N_49704);
nand UO_2136 (O_2136,N_49983,N_48912);
and UO_2137 (O_2137,N_48015,N_48534);
nand UO_2138 (O_2138,N_49157,N_49571);
xnor UO_2139 (O_2139,N_48455,N_49429);
and UO_2140 (O_2140,N_49575,N_49800);
or UO_2141 (O_2141,N_49470,N_49485);
nand UO_2142 (O_2142,N_49056,N_49476);
or UO_2143 (O_2143,N_48618,N_49079);
nand UO_2144 (O_2144,N_49935,N_49709);
or UO_2145 (O_2145,N_48482,N_48839);
xor UO_2146 (O_2146,N_49825,N_49928);
xor UO_2147 (O_2147,N_49377,N_49073);
or UO_2148 (O_2148,N_49322,N_49297);
or UO_2149 (O_2149,N_49632,N_49340);
nand UO_2150 (O_2150,N_48362,N_49886);
xor UO_2151 (O_2151,N_48629,N_49327);
nor UO_2152 (O_2152,N_48282,N_49698);
nor UO_2153 (O_2153,N_49302,N_49939);
nand UO_2154 (O_2154,N_48800,N_48179);
xor UO_2155 (O_2155,N_49216,N_49220);
nand UO_2156 (O_2156,N_48825,N_49602);
xor UO_2157 (O_2157,N_49765,N_48458);
xnor UO_2158 (O_2158,N_49077,N_49608);
and UO_2159 (O_2159,N_48077,N_48089);
or UO_2160 (O_2160,N_48405,N_49454);
or UO_2161 (O_2161,N_48975,N_48618);
or UO_2162 (O_2162,N_48912,N_48110);
or UO_2163 (O_2163,N_49562,N_49502);
nand UO_2164 (O_2164,N_49394,N_48593);
nand UO_2165 (O_2165,N_49049,N_49910);
nand UO_2166 (O_2166,N_49364,N_48965);
nor UO_2167 (O_2167,N_48725,N_49306);
or UO_2168 (O_2168,N_49405,N_48655);
nand UO_2169 (O_2169,N_49399,N_49696);
nand UO_2170 (O_2170,N_49575,N_49571);
and UO_2171 (O_2171,N_48501,N_49982);
nor UO_2172 (O_2172,N_49580,N_48898);
xnor UO_2173 (O_2173,N_49381,N_49220);
or UO_2174 (O_2174,N_49865,N_48712);
and UO_2175 (O_2175,N_49839,N_49739);
xor UO_2176 (O_2176,N_48707,N_48269);
or UO_2177 (O_2177,N_48178,N_49867);
nand UO_2178 (O_2178,N_48669,N_48638);
xnor UO_2179 (O_2179,N_48748,N_48931);
and UO_2180 (O_2180,N_49577,N_48597);
and UO_2181 (O_2181,N_48753,N_49902);
xnor UO_2182 (O_2182,N_49051,N_49361);
and UO_2183 (O_2183,N_49756,N_48478);
or UO_2184 (O_2184,N_49382,N_49875);
nand UO_2185 (O_2185,N_49695,N_48400);
xor UO_2186 (O_2186,N_49689,N_49483);
xnor UO_2187 (O_2187,N_49655,N_48765);
xor UO_2188 (O_2188,N_49423,N_49003);
xnor UO_2189 (O_2189,N_49584,N_48286);
xor UO_2190 (O_2190,N_48178,N_49577);
nor UO_2191 (O_2191,N_48071,N_48519);
xor UO_2192 (O_2192,N_49976,N_48558);
nand UO_2193 (O_2193,N_48096,N_48289);
or UO_2194 (O_2194,N_48827,N_48905);
or UO_2195 (O_2195,N_49775,N_48984);
nand UO_2196 (O_2196,N_49266,N_49112);
and UO_2197 (O_2197,N_48567,N_49252);
or UO_2198 (O_2198,N_49560,N_48123);
or UO_2199 (O_2199,N_48682,N_48425);
xor UO_2200 (O_2200,N_49799,N_49628);
nor UO_2201 (O_2201,N_49295,N_49851);
xnor UO_2202 (O_2202,N_48949,N_49211);
nand UO_2203 (O_2203,N_49017,N_49382);
nand UO_2204 (O_2204,N_48444,N_49275);
and UO_2205 (O_2205,N_49469,N_49619);
and UO_2206 (O_2206,N_48013,N_48168);
nor UO_2207 (O_2207,N_49561,N_48778);
nor UO_2208 (O_2208,N_48807,N_49819);
and UO_2209 (O_2209,N_48723,N_48114);
and UO_2210 (O_2210,N_48596,N_48839);
nor UO_2211 (O_2211,N_48989,N_48121);
xnor UO_2212 (O_2212,N_48991,N_48887);
xor UO_2213 (O_2213,N_49947,N_49904);
xnor UO_2214 (O_2214,N_49575,N_49407);
xnor UO_2215 (O_2215,N_48426,N_49405);
xor UO_2216 (O_2216,N_48591,N_49280);
nor UO_2217 (O_2217,N_49458,N_49411);
and UO_2218 (O_2218,N_49682,N_48078);
or UO_2219 (O_2219,N_49534,N_49797);
or UO_2220 (O_2220,N_48525,N_49910);
nand UO_2221 (O_2221,N_49864,N_48354);
nand UO_2222 (O_2222,N_48296,N_48222);
nor UO_2223 (O_2223,N_49237,N_48456);
and UO_2224 (O_2224,N_49993,N_49181);
or UO_2225 (O_2225,N_48911,N_48124);
and UO_2226 (O_2226,N_49324,N_49099);
or UO_2227 (O_2227,N_48015,N_49311);
xnor UO_2228 (O_2228,N_49228,N_48188);
and UO_2229 (O_2229,N_49528,N_48783);
or UO_2230 (O_2230,N_49290,N_48233);
xnor UO_2231 (O_2231,N_49336,N_48490);
and UO_2232 (O_2232,N_48027,N_49088);
xnor UO_2233 (O_2233,N_48461,N_49135);
or UO_2234 (O_2234,N_48124,N_49642);
and UO_2235 (O_2235,N_48120,N_48641);
xnor UO_2236 (O_2236,N_48043,N_48843);
xnor UO_2237 (O_2237,N_49823,N_49189);
or UO_2238 (O_2238,N_49573,N_48468);
xnor UO_2239 (O_2239,N_48814,N_48234);
nand UO_2240 (O_2240,N_48100,N_48944);
nor UO_2241 (O_2241,N_49497,N_49841);
nor UO_2242 (O_2242,N_48007,N_48270);
nand UO_2243 (O_2243,N_48567,N_48487);
nand UO_2244 (O_2244,N_48808,N_49353);
nor UO_2245 (O_2245,N_49544,N_49983);
or UO_2246 (O_2246,N_49636,N_48392);
and UO_2247 (O_2247,N_48618,N_48031);
or UO_2248 (O_2248,N_49984,N_48549);
and UO_2249 (O_2249,N_48542,N_49536);
nand UO_2250 (O_2250,N_48393,N_48890);
nor UO_2251 (O_2251,N_49450,N_49368);
nand UO_2252 (O_2252,N_49979,N_49628);
nor UO_2253 (O_2253,N_49769,N_49519);
and UO_2254 (O_2254,N_49603,N_48531);
and UO_2255 (O_2255,N_48651,N_48616);
nand UO_2256 (O_2256,N_49360,N_48306);
nand UO_2257 (O_2257,N_48291,N_49175);
nand UO_2258 (O_2258,N_48329,N_49400);
or UO_2259 (O_2259,N_48740,N_49180);
or UO_2260 (O_2260,N_48225,N_48764);
or UO_2261 (O_2261,N_49638,N_49380);
nor UO_2262 (O_2262,N_49979,N_48935);
nor UO_2263 (O_2263,N_48136,N_48280);
xor UO_2264 (O_2264,N_49649,N_49199);
nand UO_2265 (O_2265,N_48141,N_49436);
xnor UO_2266 (O_2266,N_48978,N_48340);
or UO_2267 (O_2267,N_49410,N_48726);
and UO_2268 (O_2268,N_48605,N_49365);
nor UO_2269 (O_2269,N_48452,N_48077);
xnor UO_2270 (O_2270,N_49035,N_48875);
xor UO_2271 (O_2271,N_49953,N_48844);
or UO_2272 (O_2272,N_49796,N_49213);
xnor UO_2273 (O_2273,N_49727,N_49314);
nand UO_2274 (O_2274,N_48635,N_49834);
nand UO_2275 (O_2275,N_48227,N_48594);
nand UO_2276 (O_2276,N_48225,N_49883);
nor UO_2277 (O_2277,N_49500,N_48678);
and UO_2278 (O_2278,N_48317,N_49464);
xnor UO_2279 (O_2279,N_48262,N_49638);
or UO_2280 (O_2280,N_48080,N_48110);
xor UO_2281 (O_2281,N_49430,N_48430);
xor UO_2282 (O_2282,N_49868,N_49018);
nor UO_2283 (O_2283,N_49010,N_48279);
or UO_2284 (O_2284,N_48295,N_49845);
nor UO_2285 (O_2285,N_48686,N_48623);
xor UO_2286 (O_2286,N_48860,N_49206);
nand UO_2287 (O_2287,N_49226,N_48370);
and UO_2288 (O_2288,N_48083,N_49525);
xor UO_2289 (O_2289,N_48706,N_49134);
nor UO_2290 (O_2290,N_48784,N_49601);
and UO_2291 (O_2291,N_48400,N_49266);
nor UO_2292 (O_2292,N_49280,N_48661);
and UO_2293 (O_2293,N_48080,N_48481);
nand UO_2294 (O_2294,N_49903,N_48121);
and UO_2295 (O_2295,N_49552,N_49561);
or UO_2296 (O_2296,N_49943,N_49812);
nand UO_2297 (O_2297,N_49193,N_48018);
or UO_2298 (O_2298,N_48411,N_48634);
nor UO_2299 (O_2299,N_49844,N_48863);
nor UO_2300 (O_2300,N_49798,N_49791);
nand UO_2301 (O_2301,N_48346,N_48352);
nand UO_2302 (O_2302,N_49190,N_48117);
nor UO_2303 (O_2303,N_49892,N_49472);
or UO_2304 (O_2304,N_49941,N_48618);
nor UO_2305 (O_2305,N_49123,N_48600);
or UO_2306 (O_2306,N_49807,N_48183);
nor UO_2307 (O_2307,N_49561,N_49964);
or UO_2308 (O_2308,N_48388,N_49153);
nand UO_2309 (O_2309,N_48533,N_49878);
or UO_2310 (O_2310,N_48288,N_49454);
xnor UO_2311 (O_2311,N_49506,N_48863);
nor UO_2312 (O_2312,N_48729,N_49315);
nor UO_2313 (O_2313,N_49323,N_48670);
and UO_2314 (O_2314,N_48864,N_49100);
nand UO_2315 (O_2315,N_48048,N_49764);
or UO_2316 (O_2316,N_48240,N_48780);
and UO_2317 (O_2317,N_48296,N_48522);
nor UO_2318 (O_2318,N_48843,N_48946);
and UO_2319 (O_2319,N_48214,N_49438);
or UO_2320 (O_2320,N_49131,N_48467);
or UO_2321 (O_2321,N_48098,N_49864);
and UO_2322 (O_2322,N_48147,N_48211);
or UO_2323 (O_2323,N_49420,N_49199);
nand UO_2324 (O_2324,N_48216,N_49091);
and UO_2325 (O_2325,N_48648,N_49646);
nand UO_2326 (O_2326,N_48259,N_48212);
nand UO_2327 (O_2327,N_48553,N_49907);
or UO_2328 (O_2328,N_49414,N_48760);
nand UO_2329 (O_2329,N_48717,N_49783);
or UO_2330 (O_2330,N_49140,N_49184);
and UO_2331 (O_2331,N_49648,N_49054);
nor UO_2332 (O_2332,N_48354,N_49671);
xor UO_2333 (O_2333,N_49626,N_49741);
nor UO_2334 (O_2334,N_48471,N_48522);
or UO_2335 (O_2335,N_49467,N_48791);
nor UO_2336 (O_2336,N_49850,N_49824);
xnor UO_2337 (O_2337,N_48757,N_49460);
nor UO_2338 (O_2338,N_49181,N_48190);
and UO_2339 (O_2339,N_48598,N_48498);
nor UO_2340 (O_2340,N_48418,N_48997);
or UO_2341 (O_2341,N_48268,N_48121);
nand UO_2342 (O_2342,N_49669,N_48410);
and UO_2343 (O_2343,N_49334,N_48180);
xor UO_2344 (O_2344,N_48886,N_48644);
or UO_2345 (O_2345,N_49030,N_48260);
and UO_2346 (O_2346,N_48495,N_48647);
and UO_2347 (O_2347,N_48045,N_49100);
nor UO_2348 (O_2348,N_49933,N_49504);
or UO_2349 (O_2349,N_49546,N_48944);
or UO_2350 (O_2350,N_49064,N_48778);
or UO_2351 (O_2351,N_48710,N_49813);
nor UO_2352 (O_2352,N_48875,N_48456);
or UO_2353 (O_2353,N_48524,N_49187);
or UO_2354 (O_2354,N_48647,N_48955);
and UO_2355 (O_2355,N_48472,N_49468);
xnor UO_2356 (O_2356,N_48156,N_48539);
and UO_2357 (O_2357,N_48104,N_49922);
and UO_2358 (O_2358,N_48792,N_48526);
and UO_2359 (O_2359,N_49939,N_48208);
or UO_2360 (O_2360,N_48561,N_48102);
nor UO_2361 (O_2361,N_49484,N_49627);
or UO_2362 (O_2362,N_48568,N_48675);
xor UO_2363 (O_2363,N_48918,N_48049);
xor UO_2364 (O_2364,N_48242,N_49562);
or UO_2365 (O_2365,N_48249,N_49545);
and UO_2366 (O_2366,N_49484,N_49549);
nand UO_2367 (O_2367,N_49741,N_48110);
and UO_2368 (O_2368,N_49401,N_48912);
and UO_2369 (O_2369,N_48550,N_48806);
or UO_2370 (O_2370,N_49038,N_48242);
and UO_2371 (O_2371,N_48820,N_49896);
xnor UO_2372 (O_2372,N_49664,N_49053);
and UO_2373 (O_2373,N_48896,N_48114);
xor UO_2374 (O_2374,N_49008,N_49780);
nand UO_2375 (O_2375,N_48912,N_48335);
nand UO_2376 (O_2376,N_48619,N_49682);
or UO_2377 (O_2377,N_48783,N_49470);
and UO_2378 (O_2378,N_49826,N_49226);
xnor UO_2379 (O_2379,N_48976,N_49588);
nor UO_2380 (O_2380,N_49068,N_48210);
nand UO_2381 (O_2381,N_49316,N_48379);
xnor UO_2382 (O_2382,N_48866,N_48356);
nand UO_2383 (O_2383,N_48730,N_49747);
nor UO_2384 (O_2384,N_48875,N_49664);
or UO_2385 (O_2385,N_48184,N_49911);
xor UO_2386 (O_2386,N_48497,N_49972);
xor UO_2387 (O_2387,N_48230,N_49588);
nor UO_2388 (O_2388,N_48626,N_49668);
xor UO_2389 (O_2389,N_48802,N_49021);
xnor UO_2390 (O_2390,N_48233,N_49505);
xnor UO_2391 (O_2391,N_49158,N_48456);
xnor UO_2392 (O_2392,N_49075,N_49888);
or UO_2393 (O_2393,N_48480,N_49465);
nor UO_2394 (O_2394,N_48460,N_48608);
and UO_2395 (O_2395,N_49143,N_49741);
and UO_2396 (O_2396,N_48783,N_48286);
and UO_2397 (O_2397,N_48138,N_49490);
nand UO_2398 (O_2398,N_48060,N_49533);
nor UO_2399 (O_2399,N_48723,N_49939);
and UO_2400 (O_2400,N_49673,N_49242);
xnor UO_2401 (O_2401,N_48915,N_49537);
or UO_2402 (O_2402,N_48146,N_49056);
nand UO_2403 (O_2403,N_48596,N_48057);
or UO_2404 (O_2404,N_48055,N_49193);
and UO_2405 (O_2405,N_49812,N_49058);
nor UO_2406 (O_2406,N_49092,N_49710);
or UO_2407 (O_2407,N_49526,N_48074);
or UO_2408 (O_2408,N_49958,N_49583);
xor UO_2409 (O_2409,N_48178,N_49888);
nand UO_2410 (O_2410,N_48947,N_48961);
or UO_2411 (O_2411,N_49244,N_49482);
nor UO_2412 (O_2412,N_48006,N_48945);
nor UO_2413 (O_2413,N_49725,N_49624);
nand UO_2414 (O_2414,N_49100,N_49121);
nand UO_2415 (O_2415,N_49454,N_48540);
xnor UO_2416 (O_2416,N_49174,N_48750);
nand UO_2417 (O_2417,N_48658,N_49431);
and UO_2418 (O_2418,N_49824,N_49175);
nand UO_2419 (O_2419,N_48992,N_49412);
xnor UO_2420 (O_2420,N_48444,N_49597);
and UO_2421 (O_2421,N_48052,N_48822);
xnor UO_2422 (O_2422,N_49977,N_49683);
or UO_2423 (O_2423,N_48094,N_49331);
nor UO_2424 (O_2424,N_49439,N_49283);
nor UO_2425 (O_2425,N_48354,N_49761);
nor UO_2426 (O_2426,N_48102,N_49742);
xnor UO_2427 (O_2427,N_48480,N_49269);
or UO_2428 (O_2428,N_49331,N_49306);
nand UO_2429 (O_2429,N_49787,N_48382);
or UO_2430 (O_2430,N_48051,N_48125);
xnor UO_2431 (O_2431,N_48523,N_48338);
nand UO_2432 (O_2432,N_49751,N_48012);
nand UO_2433 (O_2433,N_49814,N_49361);
nand UO_2434 (O_2434,N_49660,N_48409);
nand UO_2435 (O_2435,N_49431,N_48059);
nor UO_2436 (O_2436,N_48651,N_48218);
xnor UO_2437 (O_2437,N_48531,N_49764);
xor UO_2438 (O_2438,N_49863,N_48393);
nand UO_2439 (O_2439,N_48280,N_49862);
xor UO_2440 (O_2440,N_49870,N_49091);
and UO_2441 (O_2441,N_49455,N_48610);
nand UO_2442 (O_2442,N_49906,N_48924);
xnor UO_2443 (O_2443,N_48194,N_48383);
xnor UO_2444 (O_2444,N_48286,N_49142);
or UO_2445 (O_2445,N_49219,N_48930);
or UO_2446 (O_2446,N_48611,N_49372);
nand UO_2447 (O_2447,N_49215,N_49256);
nor UO_2448 (O_2448,N_49148,N_48906);
nor UO_2449 (O_2449,N_48526,N_48219);
nor UO_2450 (O_2450,N_48529,N_49161);
xnor UO_2451 (O_2451,N_48577,N_48765);
or UO_2452 (O_2452,N_49955,N_48190);
nand UO_2453 (O_2453,N_48536,N_49142);
xor UO_2454 (O_2454,N_49222,N_48913);
and UO_2455 (O_2455,N_49053,N_48898);
xnor UO_2456 (O_2456,N_48454,N_49802);
xnor UO_2457 (O_2457,N_48905,N_48791);
xor UO_2458 (O_2458,N_49171,N_49170);
or UO_2459 (O_2459,N_48798,N_49446);
or UO_2460 (O_2460,N_48850,N_48413);
and UO_2461 (O_2461,N_48243,N_48823);
nor UO_2462 (O_2462,N_49807,N_49537);
and UO_2463 (O_2463,N_48593,N_49234);
xnor UO_2464 (O_2464,N_48880,N_49489);
and UO_2465 (O_2465,N_48777,N_49303);
or UO_2466 (O_2466,N_48156,N_49321);
or UO_2467 (O_2467,N_48346,N_48900);
nand UO_2468 (O_2468,N_49507,N_49886);
xnor UO_2469 (O_2469,N_49339,N_49540);
xnor UO_2470 (O_2470,N_49165,N_48772);
nor UO_2471 (O_2471,N_48690,N_48095);
xnor UO_2472 (O_2472,N_49460,N_48059);
or UO_2473 (O_2473,N_49178,N_48352);
or UO_2474 (O_2474,N_48811,N_49753);
or UO_2475 (O_2475,N_48374,N_48144);
or UO_2476 (O_2476,N_48713,N_48656);
or UO_2477 (O_2477,N_48191,N_48434);
and UO_2478 (O_2478,N_48278,N_48317);
or UO_2479 (O_2479,N_49337,N_49543);
and UO_2480 (O_2480,N_48030,N_49275);
nand UO_2481 (O_2481,N_49392,N_48070);
nand UO_2482 (O_2482,N_49728,N_49343);
xor UO_2483 (O_2483,N_48191,N_49829);
xor UO_2484 (O_2484,N_49225,N_48628);
nor UO_2485 (O_2485,N_48049,N_49478);
xnor UO_2486 (O_2486,N_49011,N_48495);
xor UO_2487 (O_2487,N_48186,N_48254);
xnor UO_2488 (O_2488,N_49807,N_48800);
and UO_2489 (O_2489,N_48034,N_48598);
nor UO_2490 (O_2490,N_48210,N_48213);
nor UO_2491 (O_2491,N_49831,N_48023);
xor UO_2492 (O_2492,N_49699,N_49350);
nand UO_2493 (O_2493,N_48513,N_49256);
nand UO_2494 (O_2494,N_49463,N_49451);
nor UO_2495 (O_2495,N_48496,N_49031);
nor UO_2496 (O_2496,N_48215,N_48226);
nand UO_2497 (O_2497,N_49916,N_48761);
and UO_2498 (O_2498,N_49135,N_48938);
and UO_2499 (O_2499,N_49742,N_48709);
nand UO_2500 (O_2500,N_49160,N_48154);
xor UO_2501 (O_2501,N_49416,N_49066);
and UO_2502 (O_2502,N_48542,N_48081);
nand UO_2503 (O_2503,N_48493,N_48074);
and UO_2504 (O_2504,N_48854,N_49254);
and UO_2505 (O_2505,N_49779,N_48253);
nor UO_2506 (O_2506,N_48728,N_48056);
and UO_2507 (O_2507,N_49105,N_48149);
nor UO_2508 (O_2508,N_49600,N_48347);
nand UO_2509 (O_2509,N_48752,N_49460);
xor UO_2510 (O_2510,N_49161,N_48763);
and UO_2511 (O_2511,N_48691,N_48260);
xor UO_2512 (O_2512,N_49458,N_48764);
or UO_2513 (O_2513,N_48665,N_49033);
nor UO_2514 (O_2514,N_48595,N_48793);
nand UO_2515 (O_2515,N_49852,N_49885);
nor UO_2516 (O_2516,N_48997,N_49731);
xor UO_2517 (O_2517,N_49178,N_48908);
xnor UO_2518 (O_2518,N_49634,N_48051);
xnor UO_2519 (O_2519,N_49588,N_49177);
xor UO_2520 (O_2520,N_49240,N_48233);
nor UO_2521 (O_2521,N_49930,N_48010);
nor UO_2522 (O_2522,N_49027,N_48747);
or UO_2523 (O_2523,N_49382,N_48052);
or UO_2524 (O_2524,N_49165,N_48185);
and UO_2525 (O_2525,N_49082,N_49071);
and UO_2526 (O_2526,N_49235,N_48737);
xnor UO_2527 (O_2527,N_48247,N_49423);
xor UO_2528 (O_2528,N_49005,N_49777);
and UO_2529 (O_2529,N_49514,N_48275);
nand UO_2530 (O_2530,N_48446,N_48541);
nor UO_2531 (O_2531,N_49950,N_49924);
nand UO_2532 (O_2532,N_48557,N_49317);
nor UO_2533 (O_2533,N_49942,N_48950);
nand UO_2534 (O_2534,N_49828,N_49689);
xnor UO_2535 (O_2535,N_49120,N_49931);
nor UO_2536 (O_2536,N_49677,N_49784);
nor UO_2537 (O_2537,N_49539,N_48658);
and UO_2538 (O_2538,N_49765,N_49796);
nor UO_2539 (O_2539,N_48707,N_49777);
xor UO_2540 (O_2540,N_49412,N_49411);
nand UO_2541 (O_2541,N_48525,N_48132);
nor UO_2542 (O_2542,N_49555,N_49917);
nand UO_2543 (O_2543,N_49653,N_48448);
nor UO_2544 (O_2544,N_48502,N_48303);
nand UO_2545 (O_2545,N_48312,N_49888);
and UO_2546 (O_2546,N_48502,N_49882);
xor UO_2547 (O_2547,N_49000,N_48325);
nor UO_2548 (O_2548,N_49903,N_49433);
nand UO_2549 (O_2549,N_48069,N_48735);
and UO_2550 (O_2550,N_49958,N_48161);
xnor UO_2551 (O_2551,N_49225,N_48828);
or UO_2552 (O_2552,N_49199,N_49860);
and UO_2553 (O_2553,N_48985,N_49638);
or UO_2554 (O_2554,N_48910,N_48751);
xor UO_2555 (O_2555,N_49224,N_48440);
nor UO_2556 (O_2556,N_49200,N_48841);
and UO_2557 (O_2557,N_48632,N_49716);
xor UO_2558 (O_2558,N_48983,N_49746);
and UO_2559 (O_2559,N_48655,N_49630);
nor UO_2560 (O_2560,N_49308,N_48570);
xor UO_2561 (O_2561,N_48516,N_49463);
xnor UO_2562 (O_2562,N_48513,N_48170);
xnor UO_2563 (O_2563,N_48574,N_49974);
nor UO_2564 (O_2564,N_49709,N_49953);
or UO_2565 (O_2565,N_48567,N_48207);
or UO_2566 (O_2566,N_48635,N_48203);
nor UO_2567 (O_2567,N_48162,N_49628);
and UO_2568 (O_2568,N_48444,N_48987);
and UO_2569 (O_2569,N_49973,N_48736);
nor UO_2570 (O_2570,N_48753,N_49855);
nand UO_2571 (O_2571,N_48914,N_49469);
xnor UO_2572 (O_2572,N_49071,N_49602);
nor UO_2573 (O_2573,N_49877,N_49635);
nor UO_2574 (O_2574,N_49869,N_49887);
or UO_2575 (O_2575,N_48552,N_48236);
xnor UO_2576 (O_2576,N_49477,N_48894);
nor UO_2577 (O_2577,N_49576,N_48850);
nand UO_2578 (O_2578,N_49802,N_49424);
nand UO_2579 (O_2579,N_48790,N_48570);
xnor UO_2580 (O_2580,N_48733,N_49066);
nor UO_2581 (O_2581,N_49876,N_48691);
nand UO_2582 (O_2582,N_48725,N_49270);
and UO_2583 (O_2583,N_48428,N_48300);
and UO_2584 (O_2584,N_48686,N_49319);
or UO_2585 (O_2585,N_48600,N_48936);
nand UO_2586 (O_2586,N_48966,N_49851);
xor UO_2587 (O_2587,N_49604,N_48830);
xor UO_2588 (O_2588,N_48906,N_48625);
and UO_2589 (O_2589,N_49813,N_48681);
nor UO_2590 (O_2590,N_48103,N_48828);
nor UO_2591 (O_2591,N_49827,N_49714);
or UO_2592 (O_2592,N_48045,N_48631);
xor UO_2593 (O_2593,N_49493,N_49216);
and UO_2594 (O_2594,N_49832,N_49243);
and UO_2595 (O_2595,N_49610,N_48730);
nand UO_2596 (O_2596,N_48731,N_48543);
or UO_2597 (O_2597,N_48884,N_48145);
or UO_2598 (O_2598,N_48617,N_48998);
or UO_2599 (O_2599,N_48999,N_49567);
nor UO_2600 (O_2600,N_48776,N_49441);
nand UO_2601 (O_2601,N_48463,N_49285);
nor UO_2602 (O_2602,N_49242,N_48524);
and UO_2603 (O_2603,N_49922,N_48345);
nand UO_2604 (O_2604,N_48123,N_48868);
xor UO_2605 (O_2605,N_48557,N_48454);
xor UO_2606 (O_2606,N_48160,N_49079);
and UO_2607 (O_2607,N_49198,N_48142);
or UO_2608 (O_2608,N_49927,N_49823);
and UO_2609 (O_2609,N_48190,N_48875);
or UO_2610 (O_2610,N_49005,N_49199);
xnor UO_2611 (O_2611,N_48514,N_49361);
and UO_2612 (O_2612,N_48618,N_49827);
xnor UO_2613 (O_2613,N_49567,N_48230);
nand UO_2614 (O_2614,N_48791,N_49452);
nor UO_2615 (O_2615,N_48695,N_49529);
nand UO_2616 (O_2616,N_48135,N_49277);
nor UO_2617 (O_2617,N_48851,N_49155);
or UO_2618 (O_2618,N_49956,N_49327);
nand UO_2619 (O_2619,N_49277,N_48701);
nand UO_2620 (O_2620,N_49451,N_48199);
and UO_2621 (O_2621,N_48023,N_48324);
xnor UO_2622 (O_2622,N_48970,N_48287);
and UO_2623 (O_2623,N_48002,N_48117);
or UO_2624 (O_2624,N_48887,N_48819);
nor UO_2625 (O_2625,N_49566,N_48845);
nand UO_2626 (O_2626,N_49262,N_48406);
or UO_2627 (O_2627,N_48298,N_49975);
xor UO_2628 (O_2628,N_49473,N_48088);
nand UO_2629 (O_2629,N_48148,N_49199);
and UO_2630 (O_2630,N_49655,N_48792);
or UO_2631 (O_2631,N_49782,N_48846);
nand UO_2632 (O_2632,N_48807,N_49186);
nand UO_2633 (O_2633,N_49473,N_49346);
nor UO_2634 (O_2634,N_49158,N_49531);
or UO_2635 (O_2635,N_48305,N_48387);
nand UO_2636 (O_2636,N_49938,N_48871);
or UO_2637 (O_2637,N_49797,N_48538);
xnor UO_2638 (O_2638,N_49039,N_48602);
nor UO_2639 (O_2639,N_48247,N_48047);
or UO_2640 (O_2640,N_49057,N_48067);
nor UO_2641 (O_2641,N_49517,N_48219);
nand UO_2642 (O_2642,N_48251,N_48868);
nand UO_2643 (O_2643,N_48084,N_49913);
nor UO_2644 (O_2644,N_49758,N_49776);
nor UO_2645 (O_2645,N_48852,N_48882);
nor UO_2646 (O_2646,N_49808,N_49074);
xnor UO_2647 (O_2647,N_49639,N_48540);
and UO_2648 (O_2648,N_49942,N_49613);
and UO_2649 (O_2649,N_48271,N_49178);
and UO_2650 (O_2650,N_48266,N_48345);
nor UO_2651 (O_2651,N_48538,N_48047);
xor UO_2652 (O_2652,N_49076,N_49059);
and UO_2653 (O_2653,N_48983,N_49853);
or UO_2654 (O_2654,N_49295,N_48144);
nand UO_2655 (O_2655,N_49727,N_48670);
xnor UO_2656 (O_2656,N_48680,N_48535);
nor UO_2657 (O_2657,N_49011,N_48778);
xnor UO_2658 (O_2658,N_49976,N_48764);
nand UO_2659 (O_2659,N_48578,N_48763);
nor UO_2660 (O_2660,N_49571,N_48725);
nor UO_2661 (O_2661,N_48078,N_49522);
nand UO_2662 (O_2662,N_48196,N_48858);
nand UO_2663 (O_2663,N_48540,N_48065);
or UO_2664 (O_2664,N_48288,N_48784);
nand UO_2665 (O_2665,N_49203,N_48802);
nor UO_2666 (O_2666,N_49707,N_48199);
nand UO_2667 (O_2667,N_49734,N_48555);
nor UO_2668 (O_2668,N_49476,N_48852);
nor UO_2669 (O_2669,N_49740,N_49824);
nor UO_2670 (O_2670,N_49391,N_48032);
or UO_2671 (O_2671,N_49354,N_49560);
or UO_2672 (O_2672,N_48611,N_49098);
xnor UO_2673 (O_2673,N_48863,N_48639);
or UO_2674 (O_2674,N_49168,N_49089);
or UO_2675 (O_2675,N_49398,N_48863);
xor UO_2676 (O_2676,N_49520,N_48307);
and UO_2677 (O_2677,N_49565,N_48899);
nor UO_2678 (O_2678,N_49583,N_49989);
and UO_2679 (O_2679,N_49120,N_49438);
or UO_2680 (O_2680,N_48355,N_49661);
or UO_2681 (O_2681,N_49998,N_48354);
xor UO_2682 (O_2682,N_49838,N_49438);
nand UO_2683 (O_2683,N_49937,N_49579);
xor UO_2684 (O_2684,N_48049,N_48755);
xnor UO_2685 (O_2685,N_49588,N_48311);
or UO_2686 (O_2686,N_48620,N_48012);
nand UO_2687 (O_2687,N_49737,N_48867);
nand UO_2688 (O_2688,N_48411,N_49810);
and UO_2689 (O_2689,N_49293,N_49610);
or UO_2690 (O_2690,N_49403,N_48049);
or UO_2691 (O_2691,N_49178,N_48486);
nand UO_2692 (O_2692,N_48244,N_48544);
or UO_2693 (O_2693,N_48307,N_48363);
xor UO_2694 (O_2694,N_49479,N_49028);
xnor UO_2695 (O_2695,N_49140,N_49268);
or UO_2696 (O_2696,N_49237,N_48149);
nand UO_2697 (O_2697,N_48510,N_48080);
xnor UO_2698 (O_2698,N_49117,N_49935);
nor UO_2699 (O_2699,N_49842,N_48372);
or UO_2700 (O_2700,N_49146,N_49559);
and UO_2701 (O_2701,N_49299,N_48520);
xor UO_2702 (O_2702,N_48296,N_49974);
nor UO_2703 (O_2703,N_48569,N_49998);
or UO_2704 (O_2704,N_48196,N_48500);
nand UO_2705 (O_2705,N_49691,N_49121);
xor UO_2706 (O_2706,N_49578,N_48771);
xnor UO_2707 (O_2707,N_49688,N_49511);
or UO_2708 (O_2708,N_49385,N_48895);
xor UO_2709 (O_2709,N_49278,N_49873);
and UO_2710 (O_2710,N_48108,N_49935);
nand UO_2711 (O_2711,N_49888,N_49975);
and UO_2712 (O_2712,N_48994,N_49563);
or UO_2713 (O_2713,N_49965,N_49815);
xor UO_2714 (O_2714,N_48413,N_49350);
nand UO_2715 (O_2715,N_49112,N_48894);
and UO_2716 (O_2716,N_48000,N_48840);
xor UO_2717 (O_2717,N_48255,N_49800);
nor UO_2718 (O_2718,N_49188,N_48522);
or UO_2719 (O_2719,N_48308,N_49812);
or UO_2720 (O_2720,N_49629,N_49328);
and UO_2721 (O_2721,N_49877,N_49206);
or UO_2722 (O_2722,N_49253,N_49281);
and UO_2723 (O_2723,N_49944,N_49654);
or UO_2724 (O_2724,N_49081,N_49088);
nor UO_2725 (O_2725,N_49790,N_48959);
and UO_2726 (O_2726,N_49650,N_48918);
or UO_2727 (O_2727,N_48583,N_48281);
nor UO_2728 (O_2728,N_49321,N_48794);
xnor UO_2729 (O_2729,N_49389,N_49287);
or UO_2730 (O_2730,N_48724,N_49462);
nand UO_2731 (O_2731,N_48192,N_48071);
or UO_2732 (O_2732,N_49232,N_48158);
or UO_2733 (O_2733,N_49798,N_48206);
or UO_2734 (O_2734,N_48333,N_49802);
nor UO_2735 (O_2735,N_49857,N_49120);
nor UO_2736 (O_2736,N_48706,N_49918);
and UO_2737 (O_2737,N_48737,N_48008);
and UO_2738 (O_2738,N_49207,N_49810);
and UO_2739 (O_2739,N_48531,N_48592);
nand UO_2740 (O_2740,N_48873,N_48046);
or UO_2741 (O_2741,N_48039,N_49562);
nand UO_2742 (O_2742,N_48581,N_48787);
and UO_2743 (O_2743,N_49029,N_48454);
or UO_2744 (O_2744,N_49451,N_49023);
xor UO_2745 (O_2745,N_49479,N_48779);
xnor UO_2746 (O_2746,N_49200,N_49350);
and UO_2747 (O_2747,N_49667,N_48004);
and UO_2748 (O_2748,N_49251,N_48007);
and UO_2749 (O_2749,N_49354,N_49428);
nor UO_2750 (O_2750,N_49823,N_49402);
or UO_2751 (O_2751,N_49168,N_48672);
xor UO_2752 (O_2752,N_49176,N_48063);
or UO_2753 (O_2753,N_49624,N_48222);
xor UO_2754 (O_2754,N_48665,N_49838);
and UO_2755 (O_2755,N_49287,N_49827);
nand UO_2756 (O_2756,N_49371,N_49467);
xor UO_2757 (O_2757,N_48843,N_49029);
or UO_2758 (O_2758,N_49210,N_49241);
and UO_2759 (O_2759,N_49094,N_48125);
and UO_2760 (O_2760,N_49324,N_49962);
nand UO_2761 (O_2761,N_49555,N_49436);
nand UO_2762 (O_2762,N_48272,N_48640);
nand UO_2763 (O_2763,N_49237,N_49650);
nor UO_2764 (O_2764,N_48309,N_49463);
and UO_2765 (O_2765,N_48798,N_48793);
nand UO_2766 (O_2766,N_48738,N_48106);
and UO_2767 (O_2767,N_49885,N_49609);
nand UO_2768 (O_2768,N_49320,N_48535);
and UO_2769 (O_2769,N_48637,N_49481);
nand UO_2770 (O_2770,N_49644,N_48529);
or UO_2771 (O_2771,N_49546,N_48946);
xnor UO_2772 (O_2772,N_48184,N_49557);
nand UO_2773 (O_2773,N_49233,N_49141);
xor UO_2774 (O_2774,N_48906,N_48825);
nor UO_2775 (O_2775,N_48763,N_49899);
nand UO_2776 (O_2776,N_49798,N_49079);
nand UO_2777 (O_2777,N_49136,N_48314);
xor UO_2778 (O_2778,N_48905,N_49124);
nand UO_2779 (O_2779,N_48296,N_49665);
or UO_2780 (O_2780,N_48938,N_49314);
and UO_2781 (O_2781,N_48531,N_49238);
nand UO_2782 (O_2782,N_49530,N_48694);
and UO_2783 (O_2783,N_48243,N_49875);
or UO_2784 (O_2784,N_49101,N_49030);
nand UO_2785 (O_2785,N_48714,N_49416);
and UO_2786 (O_2786,N_49864,N_48408);
and UO_2787 (O_2787,N_48706,N_48522);
xnor UO_2788 (O_2788,N_49439,N_49649);
xor UO_2789 (O_2789,N_49597,N_49245);
xnor UO_2790 (O_2790,N_48722,N_49029);
nand UO_2791 (O_2791,N_49142,N_49020);
and UO_2792 (O_2792,N_49983,N_49324);
or UO_2793 (O_2793,N_48247,N_48007);
or UO_2794 (O_2794,N_48759,N_48765);
nor UO_2795 (O_2795,N_48454,N_49273);
xnor UO_2796 (O_2796,N_49569,N_49131);
or UO_2797 (O_2797,N_48306,N_48626);
and UO_2798 (O_2798,N_48926,N_49130);
or UO_2799 (O_2799,N_48873,N_48017);
nor UO_2800 (O_2800,N_49349,N_49933);
nor UO_2801 (O_2801,N_49243,N_49284);
and UO_2802 (O_2802,N_49937,N_48659);
nand UO_2803 (O_2803,N_49497,N_48387);
nor UO_2804 (O_2804,N_49199,N_49100);
or UO_2805 (O_2805,N_49154,N_49077);
and UO_2806 (O_2806,N_48707,N_48390);
or UO_2807 (O_2807,N_49631,N_48677);
or UO_2808 (O_2808,N_49267,N_49531);
or UO_2809 (O_2809,N_48978,N_49237);
nand UO_2810 (O_2810,N_48309,N_49360);
xor UO_2811 (O_2811,N_49958,N_48937);
and UO_2812 (O_2812,N_49365,N_49967);
nand UO_2813 (O_2813,N_49086,N_49931);
and UO_2814 (O_2814,N_48753,N_49495);
nand UO_2815 (O_2815,N_48459,N_48454);
xor UO_2816 (O_2816,N_48710,N_48906);
or UO_2817 (O_2817,N_48066,N_48781);
nor UO_2818 (O_2818,N_49376,N_48013);
nor UO_2819 (O_2819,N_49871,N_49648);
xnor UO_2820 (O_2820,N_48410,N_49872);
and UO_2821 (O_2821,N_49501,N_49224);
nor UO_2822 (O_2822,N_48071,N_49134);
nor UO_2823 (O_2823,N_48586,N_48072);
or UO_2824 (O_2824,N_48689,N_49270);
xnor UO_2825 (O_2825,N_49388,N_49135);
xor UO_2826 (O_2826,N_49771,N_49707);
nor UO_2827 (O_2827,N_49581,N_48799);
xor UO_2828 (O_2828,N_48453,N_49268);
or UO_2829 (O_2829,N_48347,N_49900);
or UO_2830 (O_2830,N_49076,N_48789);
or UO_2831 (O_2831,N_48305,N_48710);
xnor UO_2832 (O_2832,N_49994,N_49262);
and UO_2833 (O_2833,N_49567,N_48649);
nor UO_2834 (O_2834,N_48449,N_48216);
or UO_2835 (O_2835,N_49225,N_49664);
and UO_2836 (O_2836,N_49307,N_48316);
and UO_2837 (O_2837,N_48339,N_49075);
nand UO_2838 (O_2838,N_48900,N_48561);
nor UO_2839 (O_2839,N_49592,N_48702);
and UO_2840 (O_2840,N_48649,N_48688);
xnor UO_2841 (O_2841,N_49750,N_48618);
or UO_2842 (O_2842,N_49344,N_49006);
xor UO_2843 (O_2843,N_48769,N_48690);
nand UO_2844 (O_2844,N_48458,N_48816);
or UO_2845 (O_2845,N_48094,N_48659);
xnor UO_2846 (O_2846,N_49475,N_48464);
nor UO_2847 (O_2847,N_49827,N_49797);
and UO_2848 (O_2848,N_48913,N_49478);
nor UO_2849 (O_2849,N_49297,N_48715);
nand UO_2850 (O_2850,N_48144,N_48352);
or UO_2851 (O_2851,N_49938,N_49836);
or UO_2852 (O_2852,N_49818,N_48602);
nor UO_2853 (O_2853,N_49037,N_49168);
nor UO_2854 (O_2854,N_49918,N_49686);
or UO_2855 (O_2855,N_49827,N_48041);
nand UO_2856 (O_2856,N_49906,N_48225);
nand UO_2857 (O_2857,N_48214,N_49331);
nand UO_2858 (O_2858,N_48495,N_49608);
nor UO_2859 (O_2859,N_49464,N_48962);
and UO_2860 (O_2860,N_48261,N_49079);
and UO_2861 (O_2861,N_49707,N_48333);
or UO_2862 (O_2862,N_49103,N_48131);
or UO_2863 (O_2863,N_49703,N_48749);
nand UO_2864 (O_2864,N_48377,N_48339);
and UO_2865 (O_2865,N_49163,N_49077);
xnor UO_2866 (O_2866,N_48849,N_48794);
xor UO_2867 (O_2867,N_48449,N_48306);
nand UO_2868 (O_2868,N_48854,N_48996);
xor UO_2869 (O_2869,N_48765,N_48649);
or UO_2870 (O_2870,N_48574,N_49229);
nand UO_2871 (O_2871,N_48207,N_48536);
nand UO_2872 (O_2872,N_48931,N_48321);
nand UO_2873 (O_2873,N_49521,N_49405);
xnor UO_2874 (O_2874,N_48833,N_48165);
or UO_2875 (O_2875,N_49010,N_49269);
or UO_2876 (O_2876,N_48876,N_49053);
nand UO_2877 (O_2877,N_48445,N_49330);
nor UO_2878 (O_2878,N_48855,N_49964);
and UO_2879 (O_2879,N_48144,N_49049);
nor UO_2880 (O_2880,N_48560,N_49194);
and UO_2881 (O_2881,N_49804,N_49425);
or UO_2882 (O_2882,N_49621,N_49092);
and UO_2883 (O_2883,N_49259,N_48619);
and UO_2884 (O_2884,N_48676,N_48431);
or UO_2885 (O_2885,N_49629,N_49756);
xnor UO_2886 (O_2886,N_48084,N_48614);
and UO_2887 (O_2887,N_49366,N_48200);
nor UO_2888 (O_2888,N_48226,N_48361);
xnor UO_2889 (O_2889,N_49654,N_48189);
or UO_2890 (O_2890,N_49304,N_49493);
nand UO_2891 (O_2891,N_48154,N_49333);
nor UO_2892 (O_2892,N_48612,N_49966);
nor UO_2893 (O_2893,N_48671,N_48980);
or UO_2894 (O_2894,N_48401,N_49561);
nand UO_2895 (O_2895,N_49591,N_48387);
nand UO_2896 (O_2896,N_49319,N_49992);
nor UO_2897 (O_2897,N_48894,N_48977);
nor UO_2898 (O_2898,N_48792,N_48487);
xnor UO_2899 (O_2899,N_48380,N_48125);
nand UO_2900 (O_2900,N_49818,N_48888);
xnor UO_2901 (O_2901,N_48669,N_48169);
and UO_2902 (O_2902,N_48643,N_49554);
xnor UO_2903 (O_2903,N_48370,N_48569);
and UO_2904 (O_2904,N_49099,N_48266);
xnor UO_2905 (O_2905,N_48124,N_48323);
or UO_2906 (O_2906,N_48137,N_48671);
or UO_2907 (O_2907,N_49825,N_48870);
nor UO_2908 (O_2908,N_48667,N_49505);
nor UO_2909 (O_2909,N_49528,N_49430);
or UO_2910 (O_2910,N_48527,N_48981);
and UO_2911 (O_2911,N_49870,N_48341);
or UO_2912 (O_2912,N_49545,N_48082);
nor UO_2913 (O_2913,N_49366,N_48274);
nand UO_2914 (O_2914,N_48149,N_48833);
nor UO_2915 (O_2915,N_48414,N_48158);
or UO_2916 (O_2916,N_48685,N_49329);
and UO_2917 (O_2917,N_48891,N_48138);
or UO_2918 (O_2918,N_48711,N_48222);
or UO_2919 (O_2919,N_48641,N_49661);
or UO_2920 (O_2920,N_49924,N_48741);
nand UO_2921 (O_2921,N_48586,N_48404);
and UO_2922 (O_2922,N_48622,N_48743);
and UO_2923 (O_2923,N_49255,N_48842);
or UO_2924 (O_2924,N_48094,N_49905);
and UO_2925 (O_2925,N_48923,N_48886);
and UO_2926 (O_2926,N_48198,N_49324);
nand UO_2927 (O_2927,N_48809,N_49698);
nor UO_2928 (O_2928,N_49507,N_48514);
and UO_2929 (O_2929,N_49494,N_49834);
nand UO_2930 (O_2930,N_48204,N_48311);
and UO_2931 (O_2931,N_49634,N_48938);
xnor UO_2932 (O_2932,N_48189,N_48951);
nor UO_2933 (O_2933,N_48274,N_49859);
nor UO_2934 (O_2934,N_49694,N_49385);
nor UO_2935 (O_2935,N_48533,N_48421);
nand UO_2936 (O_2936,N_48984,N_48534);
xnor UO_2937 (O_2937,N_49007,N_48966);
nand UO_2938 (O_2938,N_48513,N_49088);
or UO_2939 (O_2939,N_49992,N_49430);
nand UO_2940 (O_2940,N_49221,N_49893);
xnor UO_2941 (O_2941,N_48508,N_49157);
or UO_2942 (O_2942,N_49044,N_49266);
nand UO_2943 (O_2943,N_49757,N_49133);
nor UO_2944 (O_2944,N_49169,N_49308);
and UO_2945 (O_2945,N_49710,N_48938);
nand UO_2946 (O_2946,N_49825,N_49613);
nand UO_2947 (O_2947,N_49263,N_49386);
nand UO_2948 (O_2948,N_49945,N_48260);
xor UO_2949 (O_2949,N_48527,N_49896);
nand UO_2950 (O_2950,N_49580,N_48631);
and UO_2951 (O_2951,N_48130,N_49770);
xnor UO_2952 (O_2952,N_48775,N_48379);
and UO_2953 (O_2953,N_48504,N_49588);
and UO_2954 (O_2954,N_48673,N_48408);
and UO_2955 (O_2955,N_49230,N_48419);
and UO_2956 (O_2956,N_48289,N_48655);
xor UO_2957 (O_2957,N_49499,N_48673);
and UO_2958 (O_2958,N_49853,N_49529);
nand UO_2959 (O_2959,N_49700,N_49306);
or UO_2960 (O_2960,N_49248,N_49640);
and UO_2961 (O_2961,N_49416,N_49145);
xnor UO_2962 (O_2962,N_49867,N_48534);
xnor UO_2963 (O_2963,N_48969,N_48629);
or UO_2964 (O_2964,N_49220,N_49865);
nor UO_2965 (O_2965,N_48473,N_49751);
nor UO_2966 (O_2966,N_48931,N_48339);
or UO_2967 (O_2967,N_49791,N_49251);
nor UO_2968 (O_2968,N_48769,N_48101);
xor UO_2969 (O_2969,N_48461,N_49152);
or UO_2970 (O_2970,N_49582,N_48789);
xnor UO_2971 (O_2971,N_49344,N_48646);
xor UO_2972 (O_2972,N_48948,N_48848);
nor UO_2973 (O_2973,N_49745,N_48832);
xor UO_2974 (O_2974,N_49630,N_48797);
and UO_2975 (O_2975,N_48204,N_48401);
nand UO_2976 (O_2976,N_49989,N_49682);
nand UO_2977 (O_2977,N_48594,N_48772);
xor UO_2978 (O_2978,N_49282,N_48535);
or UO_2979 (O_2979,N_49212,N_48383);
or UO_2980 (O_2980,N_49341,N_48419);
xor UO_2981 (O_2981,N_49621,N_49982);
nand UO_2982 (O_2982,N_49892,N_49854);
and UO_2983 (O_2983,N_49743,N_48782);
nand UO_2984 (O_2984,N_49853,N_49889);
nor UO_2985 (O_2985,N_49516,N_49176);
and UO_2986 (O_2986,N_48777,N_48509);
xnor UO_2987 (O_2987,N_49520,N_49901);
or UO_2988 (O_2988,N_49074,N_49741);
or UO_2989 (O_2989,N_48293,N_49729);
nor UO_2990 (O_2990,N_49798,N_48655);
and UO_2991 (O_2991,N_49593,N_48072);
and UO_2992 (O_2992,N_49795,N_49810);
or UO_2993 (O_2993,N_49311,N_48235);
and UO_2994 (O_2994,N_49864,N_48042);
nor UO_2995 (O_2995,N_48678,N_48433);
xnor UO_2996 (O_2996,N_48868,N_49826);
nor UO_2997 (O_2997,N_49354,N_48839);
or UO_2998 (O_2998,N_49747,N_48647);
or UO_2999 (O_2999,N_48346,N_48948);
or UO_3000 (O_3000,N_49244,N_48666);
nand UO_3001 (O_3001,N_48534,N_49054);
nand UO_3002 (O_3002,N_49597,N_48376);
nand UO_3003 (O_3003,N_49995,N_49078);
nand UO_3004 (O_3004,N_49931,N_48372);
xor UO_3005 (O_3005,N_49174,N_49032);
and UO_3006 (O_3006,N_48236,N_49993);
and UO_3007 (O_3007,N_49068,N_48057);
xnor UO_3008 (O_3008,N_48112,N_48722);
xnor UO_3009 (O_3009,N_48929,N_48157);
or UO_3010 (O_3010,N_49787,N_49437);
xor UO_3011 (O_3011,N_49060,N_49597);
or UO_3012 (O_3012,N_49029,N_48247);
or UO_3013 (O_3013,N_48515,N_49729);
and UO_3014 (O_3014,N_49087,N_48043);
nand UO_3015 (O_3015,N_49041,N_49233);
nand UO_3016 (O_3016,N_48926,N_48420);
and UO_3017 (O_3017,N_49317,N_48478);
or UO_3018 (O_3018,N_49095,N_49871);
and UO_3019 (O_3019,N_49918,N_49436);
and UO_3020 (O_3020,N_48361,N_49623);
or UO_3021 (O_3021,N_49293,N_48597);
xnor UO_3022 (O_3022,N_48662,N_48963);
nand UO_3023 (O_3023,N_48065,N_48551);
nor UO_3024 (O_3024,N_49872,N_48533);
nand UO_3025 (O_3025,N_49846,N_49528);
and UO_3026 (O_3026,N_49291,N_49727);
or UO_3027 (O_3027,N_49091,N_48945);
nor UO_3028 (O_3028,N_49792,N_49512);
or UO_3029 (O_3029,N_48366,N_49564);
nand UO_3030 (O_3030,N_48726,N_48126);
nand UO_3031 (O_3031,N_48692,N_49208);
xor UO_3032 (O_3032,N_48596,N_48062);
or UO_3033 (O_3033,N_49285,N_49071);
nor UO_3034 (O_3034,N_49187,N_48146);
and UO_3035 (O_3035,N_48663,N_49281);
xnor UO_3036 (O_3036,N_48720,N_49895);
nor UO_3037 (O_3037,N_49608,N_48612);
nand UO_3038 (O_3038,N_49509,N_49867);
or UO_3039 (O_3039,N_48082,N_49300);
nand UO_3040 (O_3040,N_49175,N_48083);
and UO_3041 (O_3041,N_49029,N_49694);
nand UO_3042 (O_3042,N_48274,N_49545);
and UO_3043 (O_3043,N_49129,N_48258);
nor UO_3044 (O_3044,N_48666,N_49367);
and UO_3045 (O_3045,N_48236,N_48276);
nand UO_3046 (O_3046,N_48384,N_48873);
nand UO_3047 (O_3047,N_48166,N_48545);
nor UO_3048 (O_3048,N_49866,N_48608);
or UO_3049 (O_3049,N_48667,N_49301);
xnor UO_3050 (O_3050,N_48478,N_49183);
or UO_3051 (O_3051,N_48495,N_49793);
and UO_3052 (O_3052,N_48156,N_48600);
or UO_3053 (O_3053,N_49520,N_49602);
nand UO_3054 (O_3054,N_49055,N_48146);
or UO_3055 (O_3055,N_49877,N_48006);
nand UO_3056 (O_3056,N_48722,N_48399);
and UO_3057 (O_3057,N_48721,N_48675);
or UO_3058 (O_3058,N_49344,N_48213);
or UO_3059 (O_3059,N_48414,N_49212);
or UO_3060 (O_3060,N_48146,N_48026);
or UO_3061 (O_3061,N_49835,N_48144);
xor UO_3062 (O_3062,N_48448,N_49844);
xor UO_3063 (O_3063,N_48522,N_49108);
nand UO_3064 (O_3064,N_48859,N_49564);
and UO_3065 (O_3065,N_48104,N_48350);
or UO_3066 (O_3066,N_49053,N_48996);
nand UO_3067 (O_3067,N_49397,N_49393);
xor UO_3068 (O_3068,N_49082,N_48565);
nor UO_3069 (O_3069,N_49358,N_49059);
and UO_3070 (O_3070,N_48057,N_49961);
nand UO_3071 (O_3071,N_48358,N_48242);
nand UO_3072 (O_3072,N_49159,N_48155);
nand UO_3073 (O_3073,N_49795,N_49752);
or UO_3074 (O_3074,N_49011,N_48936);
or UO_3075 (O_3075,N_49904,N_49623);
nor UO_3076 (O_3076,N_48374,N_49098);
nor UO_3077 (O_3077,N_48190,N_48904);
or UO_3078 (O_3078,N_49200,N_48083);
or UO_3079 (O_3079,N_48467,N_49234);
and UO_3080 (O_3080,N_49938,N_48988);
nand UO_3081 (O_3081,N_49299,N_48967);
xor UO_3082 (O_3082,N_49811,N_49993);
nor UO_3083 (O_3083,N_49511,N_49334);
xnor UO_3084 (O_3084,N_49208,N_49997);
nor UO_3085 (O_3085,N_48970,N_49144);
and UO_3086 (O_3086,N_49777,N_49603);
or UO_3087 (O_3087,N_48376,N_48705);
and UO_3088 (O_3088,N_49699,N_49976);
nand UO_3089 (O_3089,N_48608,N_48411);
xor UO_3090 (O_3090,N_48861,N_48003);
xnor UO_3091 (O_3091,N_48046,N_49817);
xnor UO_3092 (O_3092,N_49813,N_49644);
or UO_3093 (O_3093,N_48309,N_49982);
or UO_3094 (O_3094,N_48847,N_48222);
nor UO_3095 (O_3095,N_49005,N_49484);
nand UO_3096 (O_3096,N_48871,N_48276);
xor UO_3097 (O_3097,N_49162,N_49337);
xnor UO_3098 (O_3098,N_49587,N_48411);
xor UO_3099 (O_3099,N_49016,N_48362);
and UO_3100 (O_3100,N_49762,N_49032);
nor UO_3101 (O_3101,N_49909,N_49371);
xor UO_3102 (O_3102,N_49924,N_49976);
nand UO_3103 (O_3103,N_48907,N_49807);
nor UO_3104 (O_3104,N_49675,N_48729);
xor UO_3105 (O_3105,N_48307,N_49762);
and UO_3106 (O_3106,N_48707,N_49121);
xnor UO_3107 (O_3107,N_49948,N_49321);
xor UO_3108 (O_3108,N_49327,N_49724);
or UO_3109 (O_3109,N_49005,N_49867);
or UO_3110 (O_3110,N_48566,N_49606);
nand UO_3111 (O_3111,N_49806,N_48643);
xor UO_3112 (O_3112,N_49948,N_49628);
or UO_3113 (O_3113,N_49054,N_48624);
nor UO_3114 (O_3114,N_48686,N_49052);
nand UO_3115 (O_3115,N_49087,N_49907);
nand UO_3116 (O_3116,N_49274,N_48922);
and UO_3117 (O_3117,N_49696,N_49636);
and UO_3118 (O_3118,N_48203,N_48367);
nand UO_3119 (O_3119,N_49366,N_49396);
nand UO_3120 (O_3120,N_48328,N_49718);
nand UO_3121 (O_3121,N_49054,N_49676);
xnor UO_3122 (O_3122,N_49206,N_49285);
and UO_3123 (O_3123,N_49651,N_48635);
xor UO_3124 (O_3124,N_48010,N_48742);
nand UO_3125 (O_3125,N_49840,N_48837);
xor UO_3126 (O_3126,N_48098,N_49043);
and UO_3127 (O_3127,N_48225,N_49496);
nor UO_3128 (O_3128,N_48154,N_48204);
nor UO_3129 (O_3129,N_48339,N_49550);
and UO_3130 (O_3130,N_49953,N_48102);
and UO_3131 (O_3131,N_48483,N_49593);
nor UO_3132 (O_3132,N_49018,N_49109);
or UO_3133 (O_3133,N_48373,N_49480);
xor UO_3134 (O_3134,N_48512,N_48723);
nand UO_3135 (O_3135,N_48584,N_49273);
nor UO_3136 (O_3136,N_49034,N_49727);
nor UO_3137 (O_3137,N_49169,N_48145);
xor UO_3138 (O_3138,N_48377,N_49441);
nor UO_3139 (O_3139,N_49114,N_48482);
nor UO_3140 (O_3140,N_48469,N_48296);
nor UO_3141 (O_3141,N_49169,N_49024);
nand UO_3142 (O_3142,N_48286,N_48015);
nor UO_3143 (O_3143,N_49430,N_48751);
or UO_3144 (O_3144,N_49622,N_49336);
xnor UO_3145 (O_3145,N_49856,N_48650);
nor UO_3146 (O_3146,N_49401,N_49065);
or UO_3147 (O_3147,N_49106,N_48462);
nor UO_3148 (O_3148,N_48843,N_48051);
or UO_3149 (O_3149,N_49131,N_48323);
and UO_3150 (O_3150,N_49490,N_49887);
or UO_3151 (O_3151,N_49060,N_49668);
or UO_3152 (O_3152,N_48988,N_48754);
nand UO_3153 (O_3153,N_48381,N_49071);
nor UO_3154 (O_3154,N_48348,N_49507);
and UO_3155 (O_3155,N_49982,N_49228);
xor UO_3156 (O_3156,N_48019,N_49311);
or UO_3157 (O_3157,N_48261,N_49956);
and UO_3158 (O_3158,N_49707,N_49651);
nor UO_3159 (O_3159,N_48434,N_48950);
and UO_3160 (O_3160,N_49621,N_48498);
xnor UO_3161 (O_3161,N_48964,N_49822);
nor UO_3162 (O_3162,N_48077,N_49361);
or UO_3163 (O_3163,N_49056,N_48697);
nor UO_3164 (O_3164,N_49509,N_48327);
and UO_3165 (O_3165,N_49016,N_49608);
nand UO_3166 (O_3166,N_49000,N_48432);
and UO_3167 (O_3167,N_48124,N_49593);
or UO_3168 (O_3168,N_48994,N_48871);
nand UO_3169 (O_3169,N_49263,N_49147);
and UO_3170 (O_3170,N_49802,N_48932);
or UO_3171 (O_3171,N_49360,N_48248);
nor UO_3172 (O_3172,N_48664,N_49158);
xor UO_3173 (O_3173,N_49741,N_49981);
and UO_3174 (O_3174,N_48043,N_48001);
nor UO_3175 (O_3175,N_48956,N_49787);
nand UO_3176 (O_3176,N_48557,N_48264);
xor UO_3177 (O_3177,N_49398,N_49003);
nor UO_3178 (O_3178,N_48187,N_49873);
nor UO_3179 (O_3179,N_48916,N_48492);
and UO_3180 (O_3180,N_49101,N_48734);
and UO_3181 (O_3181,N_49183,N_49220);
and UO_3182 (O_3182,N_49196,N_48552);
xnor UO_3183 (O_3183,N_48424,N_48430);
xnor UO_3184 (O_3184,N_48917,N_48887);
and UO_3185 (O_3185,N_49264,N_49385);
nand UO_3186 (O_3186,N_48647,N_49263);
nor UO_3187 (O_3187,N_49312,N_49654);
or UO_3188 (O_3188,N_49176,N_49055);
and UO_3189 (O_3189,N_49523,N_48360);
or UO_3190 (O_3190,N_49522,N_48095);
nor UO_3191 (O_3191,N_48753,N_49319);
nand UO_3192 (O_3192,N_48152,N_48219);
nand UO_3193 (O_3193,N_49460,N_48563);
nor UO_3194 (O_3194,N_49257,N_48384);
or UO_3195 (O_3195,N_49290,N_49125);
or UO_3196 (O_3196,N_49292,N_49025);
or UO_3197 (O_3197,N_48334,N_48761);
nand UO_3198 (O_3198,N_48698,N_49313);
xnor UO_3199 (O_3199,N_48867,N_49905);
nor UO_3200 (O_3200,N_49101,N_48051);
and UO_3201 (O_3201,N_48796,N_48882);
and UO_3202 (O_3202,N_48349,N_49817);
nand UO_3203 (O_3203,N_48834,N_49651);
and UO_3204 (O_3204,N_49190,N_48593);
or UO_3205 (O_3205,N_48132,N_49260);
xor UO_3206 (O_3206,N_48865,N_49302);
xnor UO_3207 (O_3207,N_49909,N_49975);
nor UO_3208 (O_3208,N_48964,N_48738);
or UO_3209 (O_3209,N_49675,N_49116);
and UO_3210 (O_3210,N_49053,N_49460);
nor UO_3211 (O_3211,N_49082,N_48835);
xor UO_3212 (O_3212,N_49751,N_48984);
or UO_3213 (O_3213,N_49757,N_48861);
nand UO_3214 (O_3214,N_48332,N_49444);
nor UO_3215 (O_3215,N_48132,N_49578);
or UO_3216 (O_3216,N_49633,N_49148);
or UO_3217 (O_3217,N_48275,N_48761);
xor UO_3218 (O_3218,N_49667,N_48148);
or UO_3219 (O_3219,N_48659,N_48565);
xnor UO_3220 (O_3220,N_49201,N_48752);
and UO_3221 (O_3221,N_49936,N_48790);
and UO_3222 (O_3222,N_49638,N_49711);
or UO_3223 (O_3223,N_48757,N_49714);
or UO_3224 (O_3224,N_49712,N_49716);
and UO_3225 (O_3225,N_48084,N_49029);
and UO_3226 (O_3226,N_49827,N_48284);
nand UO_3227 (O_3227,N_49993,N_49632);
nand UO_3228 (O_3228,N_48696,N_49661);
and UO_3229 (O_3229,N_48881,N_48068);
nor UO_3230 (O_3230,N_49355,N_49227);
nor UO_3231 (O_3231,N_49633,N_48640);
or UO_3232 (O_3232,N_49920,N_48113);
nor UO_3233 (O_3233,N_49507,N_48350);
nand UO_3234 (O_3234,N_48972,N_49731);
and UO_3235 (O_3235,N_49188,N_48496);
xor UO_3236 (O_3236,N_49479,N_49991);
nand UO_3237 (O_3237,N_48970,N_49584);
and UO_3238 (O_3238,N_49989,N_48412);
or UO_3239 (O_3239,N_48833,N_49978);
and UO_3240 (O_3240,N_48306,N_49269);
xnor UO_3241 (O_3241,N_48393,N_48651);
and UO_3242 (O_3242,N_48419,N_48308);
nor UO_3243 (O_3243,N_49561,N_49076);
or UO_3244 (O_3244,N_49363,N_48573);
and UO_3245 (O_3245,N_48950,N_48517);
and UO_3246 (O_3246,N_48570,N_49085);
and UO_3247 (O_3247,N_48822,N_49362);
and UO_3248 (O_3248,N_48956,N_49403);
xor UO_3249 (O_3249,N_49059,N_48330);
or UO_3250 (O_3250,N_49341,N_49281);
nand UO_3251 (O_3251,N_48776,N_48794);
or UO_3252 (O_3252,N_49350,N_49615);
nand UO_3253 (O_3253,N_48805,N_48488);
and UO_3254 (O_3254,N_49842,N_49111);
nand UO_3255 (O_3255,N_49386,N_48751);
nor UO_3256 (O_3256,N_49963,N_48902);
xnor UO_3257 (O_3257,N_48283,N_49434);
or UO_3258 (O_3258,N_48457,N_48659);
or UO_3259 (O_3259,N_49461,N_49420);
nand UO_3260 (O_3260,N_48818,N_48711);
and UO_3261 (O_3261,N_48357,N_48603);
nor UO_3262 (O_3262,N_48747,N_48089);
xor UO_3263 (O_3263,N_48549,N_48945);
xnor UO_3264 (O_3264,N_49506,N_48080);
and UO_3265 (O_3265,N_48585,N_49715);
and UO_3266 (O_3266,N_49136,N_48559);
and UO_3267 (O_3267,N_49201,N_48605);
xnor UO_3268 (O_3268,N_49495,N_49750);
nor UO_3269 (O_3269,N_48057,N_49768);
or UO_3270 (O_3270,N_48046,N_49894);
and UO_3271 (O_3271,N_49140,N_48224);
or UO_3272 (O_3272,N_48325,N_48711);
nand UO_3273 (O_3273,N_49009,N_49869);
nand UO_3274 (O_3274,N_48426,N_49888);
nand UO_3275 (O_3275,N_48151,N_49385);
or UO_3276 (O_3276,N_48969,N_49585);
and UO_3277 (O_3277,N_48106,N_48802);
nor UO_3278 (O_3278,N_49390,N_48276);
nor UO_3279 (O_3279,N_49111,N_48110);
and UO_3280 (O_3280,N_49665,N_49994);
or UO_3281 (O_3281,N_49010,N_48169);
or UO_3282 (O_3282,N_49941,N_48032);
xnor UO_3283 (O_3283,N_48181,N_49052);
nor UO_3284 (O_3284,N_49183,N_49619);
or UO_3285 (O_3285,N_49539,N_48104);
nand UO_3286 (O_3286,N_49014,N_48909);
and UO_3287 (O_3287,N_49995,N_49644);
and UO_3288 (O_3288,N_48889,N_49696);
or UO_3289 (O_3289,N_48180,N_48522);
nand UO_3290 (O_3290,N_48103,N_48629);
and UO_3291 (O_3291,N_48746,N_48340);
xor UO_3292 (O_3292,N_49361,N_48211);
nand UO_3293 (O_3293,N_48838,N_48877);
nor UO_3294 (O_3294,N_49338,N_48561);
nand UO_3295 (O_3295,N_48576,N_49206);
nand UO_3296 (O_3296,N_49957,N_48118);
nand UO_3297 (O_3297,N_49462,N_49818);
nor UO_3298 (O_3298,N_48221,N_49098);
nor UO_3299 (O_3299,N_48748,N_49994);
nand UO_3300 (O_3300,N_48982,N_49695);
and UO_3301 (O_3301,N_48833,N_48720);
nor UO_3302 (O_3302,N_48747,N_49526);
or UO_3303 (O_3303,N_49941,N_48223);
xnor UO_3304 (O_3304,N_49568,N_48287);
xor UO_3305 (O_3305,N_48694,N_49849);
or UO_3306 (O_3306,N_49933,N_49597);
and UO_3307 (O_3307,N_48420,N_48265);
xor UO_3308 (O_3308,N_49926,N_49922);
nor UO_3309 (O_3309,N_49907,N_49580);
nand UO_3310 (O_3310,N_49377,N_48964);
nand UO_3311 (O_3311,N_49687,N_49422);
nand UO_3312 (O_3312,N_49152,N_49574);
nor UO_3313 (O_3313,N_49370,N_49496);
or UO_3314 (O_3314,N_49286,N_48407);
and UO_3315 (O_3315,N_48333,N_49886);
nor UO_3316 (O_3316,N_48357,N_49404);
or UO_3317 (O_3317,N_49410,N_49053);
and UO_3318 (O_3318,N_49737,N_48418);
nand UO_3319 (O_3319,N_49115,N_49411);
nand UO_3320 (O_3320,N_49606,N_49435);
and UO_3321 (O_3321,N_49142,N_49433);
nor UO_3322 (O_3322,N_49952,N_48657);
or UO_3323 (O_3323,N_49307,N_48083);
xnor UO_3324 (O_3324,N_48725,N_49272);
and UO_3325 (O_3325,N_49166,N_48073);
xor UO_3326 (O_3326,N_49780,N_48800);
nor UO_3327 (O_3327,N_49245,N_48496);
and UO_3328 (O_3328,N_48310,N_48969);
and UO_3329 (O_3329,N_49196,N_49877);
nand UO_3330 (O_3330,N_48751,N_49407);
xor UO_3331 (O_3331,N_49892,N_48176);
nand UO_3332 (O_3332,N_48010,N_49184);
nor UO_3333 (O_3333,N_49561,N_48333);
xnor UO_3334 (O_3334,N_49576,N_49929);
nor UO_3335 (O_3335,N_49995,N_49533);
xor UO_3336 (O_3336,N_49565,N_48637);
and UO_3337 (O_3337,N_48491,N_49208);
xnor UO_3338 (O_3338,N_48057,N_48694);
or UO_3339 (O_3339,N_49219,N_49697);
xnor UO_3340 (O_3340,N_49853,N_48964);
nor UO_3341 (O_3341,N_48145,N_48887);
nor UO_3342 (O_3342,N_49443,N_48425);
and UO_3343 (O_3343,N_48357,N_49206);
xnor UO_3344 (O_3344,N_48978,N_49991);
or UO_3345 (O_3345,N_48591,N_49320);
xnor UO_3346 (O_3346,N_48455,N_49545);
or UO_3347 (O_3347,N_48159,N_49289);
or UO_3348 (O_3348,N_49555,N_48303);
xnor UO_3349 (O_3349,N_49442,N_48674);
or UO_3350 (O_3350,N_49402,N_48780);
nor UO_3351 (O_3351,N_48687,N_48717);
xnor UO_3352 (O_3352,N_48833,N_49899);
xor UO_3353 (O_3353,N_48509,N_49562);
nor UO_3354 (O_3354,N_48628,N_48070);
nand UO_3355 (O_3355,N_49522,N_49282);
nand UO_3356 (O_3356,N_48188,N_48906);
nand UO_3357 (O_3357,N_49467,N_49697);
nor UO_3358 (O_3358,N_48649,N_48913);
nor UO_3359 (O_3359,N_48306,N_49079);
or UO_3360 (O_3360,N_48959,N_48225);
nand UO_3361 (O_3361,N_48583,N_49532);
and UO_3362 (O_3362,N_48419,N_48275);
nor UO_3363 (O_3363,N_48408,N_48188);
xor UO_3364 (O_3364,N_49862,N_49215);
nor UO_3365 (O_3365,N_48040,N_49469);
and UO_3366 (O_3366,N_49260,N_48080);
xor UO_3367 (O_3367,N_48042,N_49070);
and UO_3368 (O_3368,N_49908,N_49406);
and UO_3369 (O_3369,N_49460,N_48098);
or UO_3370 (O_3370,N_48837,N_48967);
nor UO_3371 (O_3371,N_49139,N_49720);
or UO_3372 (O_3372,N_49834,N_48512);
nor UO_3373 (O_3373,N_49193,N_48781);
or UO_3374 (O_3374,N_49168,N_49297);
nor UO_3375 (O_3375,N_49704,N_48402);
xnor UO_3376 (O_3376,N_49478,N_48271);
or UO_3377 (O_3377,N_48933,N_48602);
xor UO_3378 (O_3378,N_48769,N_48973);
nor UO_3379 (O_3379,N_48693,N_48650);
nor UO_3380 (O_3380,N_49546,N_48827);
and UO_3381 (O_3381,N_48017,N_48711);
or UO_3382 (O_3382,N_49376,N_49377);
or UO_3383 (O_3383,N_49382,N_48460);
xnor UO_3384 (O_3384,N_49531,N_48604);
nand UO_3385 (O_3385,N_49112,N_49111);
xor UO_3386 (O_3386,N_48682,N_49327);
nand UO_3387 (O_3387,N_48090,N_48610);
or UO_3388 (O_3388,N_48969,N_49761);
and UO_3389 (O_3389,N_48204,N_49685);
or UO_3390 (O_3390,N_48692,N_49039);
xnor UO_3391 (O_3391,N_48355,N_49212);
or UO_3392 (O_3392,N_49150,N_48513);
or UO_3393 (O_3393,N_48587,N_48847);
nand UO_3394 (O_3394,N_48222,N_48018);
or UO_3395 (O_3395,N_48846,N_49161);
nor UO_3396 (O_3396,N_48422,N_48155);
and UO_3397 (O_3397,N_48425,N_48108);
xor UO_3398 (O_3398,N_49385,N_49073);
xnor UO_3399 (O_3399,N_48281,N_48087);
and UO_3400 (O_3400,N_48402,N_48989);
xor UO_3401 (O_3401,N_48697,N_49800);
and UO_3402 (O_3402,N_48805,N_48386);
xnor UO_3403 (O_3403,N_48592,N_49803);
or UO_3404 (O_3404,N_49595,N_49819);
nor UO_3405 (O_3405,N_48347,N_48343);
or UO_3406 (O_3406,N_49696,N_48745);
nand UO_3407 (O_3407,N_49536,N_49747);
or UO_3408 (O_3408,N_49068,N_49574);
and UO_3409 (O_3409,N_48387,N_49104);
and UO_3410 (O_3410,N_49771,N_48498);
xnor UO_3411 (O_3411,N_48779,N_49514);
xnor UO_3412 (O_3412,N_48689,N_48647);
nor UO_3413 (O_3413,N_49194,N_49657);
nor UO_3414 (O_3414,N_48926,N_49733);
or UO_3415 (O_3415,N_48019,N_49645);
xor UO_3416 (O_3416,N_48571,N_48517);
and UO_3417 (O_3417,N_48073,N_49014);
nor UO_3418 (O_3418,N_49334,N_49895);
nor UO_3419 (O_3419,N_49430,N_48177);
and UO_3420 (O_3420,N_48262,N_49585);
nor UO_3421 (O_3421,N_49219,N_49277);
or UO_3422 (O_3422,N_48125,N_48592);
and UO_3423 (O_3423,N_49033,N_49028);
xnor UO_3424 (O_3424,N_48170,N_48251);
and UO_3425 (O_3425,N_48552,N_48472);
and UO_3426 (O_3426,N_48612,N_48624);
or UO_3427 (O_3427,N_48665,N_48316);
or UO_3428 (O_3428,N_48577,N_49629);
xor UO_3429 (O_3429,N_48564,N_48347);
or UO_3430 (O_3430,N_49483,N_49059);
and UO_3431 (O_3431,N_49202,N_49714);
xor UO_3432 (O_3432,N_48674,N_49042);
nand UO_3433 (O_3433,N_49903,N_48487);
nand UO_3434 (O_3434,N_48028,N_49822);
and UO_3435 (O_3435,N_48583,N_48669);
and UO_3436 (O_3436,N_48787,N_48234);
nor UO_3437 (O_3437,N_49443,N_49163);
xor UO_3438 (O_3438,N_49702,N_49945);
nand UO_3439 (O_3439,N_49213,N_49635);
nand UO_3440 (O_3440,N_48772,N_49072);
xnor UO_3441 (O_3441,N_48271,N_48905);
nor UO_3442 (O_3442,N_49042,N_49138);
and UO_3443 (O_3443,N_49503,N_48156);
and UO_3444 (O_3444,N_49066,N_49532);
and UO_3445 (O_3445,N_48637,N_48908);
and UO_3446 (O_3446,N_49542,N_48746);
and UO_3447 (O_3447,N_48775,N_48073);
and UO_3448 (O_3448,N_48724,N_49121);
nand UO_3449 (O_3449,N_49294,N_48876);
xnor UO_3450 (O_3450,N_48774,N_48300);
or UO_3451 (O_3451,N_48643,N_49617);
nand UO_3452 (O_3452,N_48510,N_49767);
nand UO_3453 (O_3453,N_48069,N_48468);
xnor UO_3454 (O_3454,N_49778,N_48043);
nand UO_3455 (O_3455,N_48560,N_49372);
and UO_3456 (O_3456,N_49237,N_49218);
or UO_3457 (O_3457,N_49683,N_49531);
xor UO_3458 (O_3458,N_49358,N_48452);
nor UO_3459 (O_3459,N_48909,N_49504);
nand UO_3460 (O_3460,N_48996,N_49330);
nand UO_3461 (O_3461,N_48357,N_48657);
nand UO_3462 (O_3462,N_49079,N_49178);
or UO_3463 (O_3463,N_49271,N_48809);
xor UO_3464 (O_3464,N_49443,N_48798);
xnor UO_3465 (O_3465,N_49377,N_48788);
and UO_3466 (O_3466,N_48411,N_49286);
xor UO_3467 (O_3467,N_49912,N_48280);
and UO_3468 (O_3468,N_49566,N_48782);
or UO_3469 (O_3469,N_49389,N_49010);
and UO_3470 (O_3470,N_49375,N_49519);
xnor UO_3471 (O_3471,N_48244,N_49274);
nand UO_3472 (O_3472,N_48730,N_48057);
nor UO_3473 (O_3473,N_48525,N_49059);
nor UO_3474 (O_3474,N_48732,N_49862);
and UO_3475 (O_3475,N_48492,N_49825);
nor UO_3476 (O_3476,N_48544,N_48481);
and UO_3477 (O_3477,N_48963,N_49259);
nor UO_3478 (O_3478,N_49767,N_48578);
or UO_3479 (O_3479,N_49896,N_48710);
and UO_3480 (O_3480,N_48740,N_49300);
xnor UO_3481 (O_3481,N_48990,N_49261);
nor UO_3482 (O_3482,N_48962,N_49295);
and UO_3483 (O_3483,N_48225,N_49275);
xnor UO_3484 (O_3484,N_48855,N_49892);
xnor UO_3485 (O_3485,N_48179,N_49398);
nor UO_3486 (O_3486,N_49644,N_48472);
or UO_3487 (O_3487,N_49193,N_48197);
nand UO_3488 (O_3488,N_48264,N_49162);
nor UO_3489 (O_3489,N_48663,N_49758);
or UO_3490 (O_3490,N_48248,N_49742);
nand UO_3491 (O_3491,N_48949,N_48002);
xor UO_3492 (O_3492,N_49201,N_49641);
or UO_3493 (O_3493,N_49360,N_49444);
xor UO_3494 (O_3494,N_48933,N_48913);
and UO_3495 (O_3495,N_48429,N_48427);
or UO_3496 (O_3496,N_48193,N_48903);
nand UO_3497 (O_3497,N_48954,N_48519);
and UO_3498 (O_3498,N_48181,N_48815);
nor UO_3499 (O_3499,N_49555,N_49305);
or UO_3500 (O_3500,N_48932,N_49598);
and UO_3501 (O_3501,N_49042,N_49725);
xor UO_3502 (O_3502,N_48998,N_48623);
xor UO_3503 (O_3503,N_49437,N_49669);
or UO_3504 (O_3504,N_48913,N_48854);
and UO_3505 (O_3505,N_48058,N_48755);
nor UO_3506 (O_3506,N_49978,N_48077);
xor UO_3507 (O_3507,N_48733,N_48749);
and UO_3508 (O_3508,N_49488,N_48382);
nand UO_3509 (O_3509,N_49249,N_48907);
and UO_3510 (O_3510,N_48181,N_49364);
and UO_3511 (O_3511,N_49301,N_48666);
xnor UO_3512 (O_3512,N_48929,N_49851);
xnor UO_3513 (O_3513,N_49330,N_48878);
and UO_3514 (O_3514,N_48420,N_48523);
and UO_3515 (O_3515,N_48572,N_49766);
nand UO_3516 (O_3516,N_49905,N_49698);
nor UO_3517 (O_3517,N_49335,N_48933);
and UO_3518 (O_3518,N_49235,N_49055);
and UO_3519 (O_3519,N_48770,N_48054);
nand UO_3520 (O_3520,N_48687,N_48763);
xnor UO_3521 (O_3521,N_49626,N_48698);
and UO_3522 (O_3522,N_49731,N_48984);
nor UO_3523 (O_3523,N_48176,N_48281);
and UO_3524 (O_3524,N_49461,N_48379);
nand UO_3525 (O_3525,N_49157,N_49076);
nor UO_3526 (O_3526,N_49432,N_48193);
and UO_3527 (O_3527,N_49987,N_48112);
and UO_3528 (O_3528,N_48726,N_49705);
nand UO_3529 (O_3529,N_48756,N_48119);
nand UO_3530 (O_3530,N_48925,N_49948);
xor UO_3531 (O_3531,N_48721,N_48541);
nor UO_3532 (O_3532,N_49370,N_48397);
xnor UO_3533 (O_3533,N_48028,N_49802);
or UO_3534 (O_3534,N_49103,N_49859);
nand UO_3535 (O_3535,N_48425,N_49337);
nand UO_3536 (O_3536,N_48910,N_48029);
or UO_3537 (O_3537,N_49760,N_48683);
nor UO_3538 (O_3538,N_49252,N_49911);
and UO_3539 (O_3539,N_49030,N_49209);
xnor UO_3540 (O_3540,N_48944,N_48942);
nand UO_3541 (O_3541,N_48444,N_49681);
or UO_3542 (O_3542,N_49985,N_48829);
and UO_3543 (O_3543,N_49027,N_48307);
xor UO_3544 (O_3544,N_48146,N_48050);
or UO_3545 (O_3545,N_48273,N_49131);
nand UO_3546 (O_3546,N_49010,N_49921);
or UO_3547 (O_3547,N_48089,N_49478);
nor UO_3548 (O_3548,N_48492,N_48924);
and UO_3549 (O_3549,N_49054,N_49581);
nor UO_3550 (O_3550,N_49153,N_49147);
or UO_3551 (O_3551,N_49009,N_48963);
or UO_3552 (O_3552,N_49803,N_49341);
or UO_3553 (O_3553,N_48905,N_48087);
nand UO_3554 (O_3554,N_49314,N_48438);
or UO_3555 (O_3555,N_49213,N_48092);
and UO_3556 (O_3556,N_49082,N_48317);
xor UO_3557 (O_3557,N_48748,N_49876);
nand UO_3558 (O_3558,N_49025,N_48071);
nor UO_3559 (O_3559,N_49953,N_49730);
xor UO_3560 (O_3560,N_48225,N_48087);
nand UO_3561 (O_3561,N_48390,N_49546);
xor UO_3562 (O_3562,N_48569,N_49938);
nor UO_3563 (O_3563,N_49310,N_49803);
nand UO_3564 (O_3564,N_48001,N_49062);
and UO_3565 (O_3565,N_48185,N_49078);
or UO_3566 (O_3566,N_49933,N_49904);
nand UO_3567 (O_3567,N_48611,N_49254);
and UO_3568 (O_3568,N_48091,N_49180);
xor UO_3569 (O_3569,N_49661,N_49796);
xnor UO_3570 (O_3570,N_49493,N_48991);
nor UO_3571 (O_3571,N_48580,N_48965);
nor UO_3572 (O_3572,N_49195,N_48776);
nand UO_3573 (O_3573,N_48587,N_48882);
nand UO_3574 (O_3574,N_48032,N_49291);
nand UO_3575 (O_3575,N_49385,N_48709);
and UO_3576 (O_3576,N_49087,N_48968);
nand UO_3577 (O_3577,N_48445,N_49430);
xor UO_3578 (O_3578,N_48435,N_49147);
xnor UO_3579 (O_3579,N_48032,N_48588);
and UO_3580 (O_3580,N_49080,N_49809);
and UO_3581 (O_3581,N_49779,N_48846);
or UO_3582 (O_3582,N_49678,N_48991);
and UO_3583 (O_3583,N_49535,N_49285);
and UO_3584 (O_3584,N_49067,N_49010);
or UO_3585 (O_3585,N_49995,N_48900);
and UO_3586 (O_3586,N_49318,N_49294);
xnor UO_3587 (O_3587,N_48853,N_48166);
nand UO_3588 (O_3588,N_49438,N_48829);
nand UO_3589 (O_3589,N_48822,N_48223);
or UO_3590 (O_3590,N_48363,N_49504);
nor UO_3591 (O_3591,N_48987,N_48132);
and UO_3592 (O_3592,N_49634,N_48254);
or UO_3593 (O_3593,N_49065,N_48745);
xnor UO_3594 (O_3594,N_49708,N_49970);
nor UO_3595 (O_3595,N_48551,N_48493);
nand UO_3596 (O_3596,N_48420,N_49816);
nor UO_3597 (O_3597,N_48622,N_48000);
nand UO_3598 (O_3598,N_48097,N_49460);
nand UO_3599 (O_3599,N_49210,N_48707);
nor UO_3600 (O_3600,N_48232,N_49175);
nor UO_3601 (O_3601,N_48435,N_49647);
nand UO_3602 (O_3602,N_49215,N_49403);
or UO_3603 (O_3603,N_49691,N_48197);
nand UO_3604 (O_3604,N_48815,N_48905);
and UO_3605 (O_3605,N_49932,N_48400);
xnor UO_3606 (O_3606,N_48676,N_49742);
or UO_3607 (O_3607,N_49250,N_49145);
xnor UO_3608 (O_3608,N_49166,N_48405);
nand UO_3609 (O_3609,N_48821,N_48019);
nor UO_3610 (O_3610,N_48960,N_49429);
xor UO_3611 (O_3611,N_49218,N_49229);
and UO_3612 (O_3612,N_48087,N_49231);
and UO_3613 (O_3613,N_49814,N_48244);
xnor UO_3614 (O_3614,N_48937,N_49508);
xor UO_3615 (O_3615,N_49352,N_48763);
nand UO_3616 (O_3616,N_48506,N_49627);
and UO_3617 (O_3617,N_48861,N_49189);
xnor UO_3618 (O_3618,N_49857,N_48308);
nor UO_3619 (O_3619,N_48423,N_49246);
xnor UO_3620 (O_3620,N_49155,N_49848);
and UO_3621 (O_3621,N_49395,N_49854);
nand UO_3622 (O_3622,N_48588,N_48506);
nand UO_3623 (O_3623,N_48459,N_48728);
nor UO_3624 (O_3624,N_48718,N_48531);
xor UO_3625 (O_3625,N_49169,N_49952);
nand UO_3626 (O_3626,N_48963,N_49360);
and UO_3627 (O_3627,N_49529,N_48113);
or UO_3628 (O_3628,N_49049,N_48896);
xnor UO_3629 (O_3629,N_49483,N_49167);
or UO_3630 (O_3630,N_48707,N_48077);
nor UO_3631 (O_3631,N_49977,N_48749);
or UO_3632 (O_3632,N_49519,N_49142);
nand UO_3633 (O_3633,N_49909,N_49586);
nor UO_3634 (O_3634,N_48421,N_48181);
nor UO_3635 (O_3635,N_48167,N_48033);
or UO_3636 (O_3636,N_48117,N_49478);
nand UO_3637 (O_3637,N_48583,N_49277);
nor UO_3638 (O_3638,N_48294,N_48257);
and UO_3639 (O_3639,N_49844,N_49288);
and UO_3640 (O_3640,N_48087,N_49568);
nand UO_3641 (O_3641,N_48849,N_49010);
nand UO_3642 (O_3642,N_49654,N_48333);
nor UO_3643 (O_3643,N_48703,N_49235);
nand UO_3644 (O_3644,N_49615,N_48261);
xor UO_3645 (O_3645,N_48097,N_49428);
or UO_3646 (O_3646,N_49345,N_49566);
or UO_3647 (O_3647,N_49907,N_48108);
nor UO_3648 (O_3648,N_48782,N_48069);
or UO_3649 (O_3649,N_49896,N_49964);
nand UO_3650 (O_3650,N_49554,N_48017);
and UO_3651 (O_3651,N_49571,N_48000);
or UO_3652 (O_3652,N_48734,N_49095);
or UO_3653 (O_3653,N_48233,N_48843);
or UO_3654 (O_3654,N_48425,N_48381);
nor UO_3655 (O_3655,N_49025,N_49740);
or UO_3656 (O_3656,N_49828,N_48527);
nor UO_3657 (O_3657,N_48945,N_49225);
nand UO_3658 (O_3658,N_48146,N_48680);
and UO_3659 (O_3659,N_49016,N_49978);
nor UO_3660 (O_3660,N_48910,N_48917);
and UO_3661 (O_3661,N_48184,N_49518);
nor UO_3662 (O_3662,N_48315,N_49750);
and UO_3663 (O_3663,N_49058,N_49653);
nor UO_3664 (O_3664,N_49715,N_49839);
xnor UO_3665 (O_3665,N_49824,N_49388);
and UO_3666 (O_3666,N_48728,N_48826);
or UO_3667 (O_3667,N_48245,N_48082);
xnor UO_3668 (O_3668,N_48821,N_49732);
nor UO_3669 (O_3669,N_48638,N_48046);
or UO_3670 (O_3670,N_48611,N_49338);
and UO_3671 (O_3671,N_49350,N_48437);
nand UO_3672 (O_3672,N_48793,N_49873);
xnor UO_3673 (O_3673,N_49542,N_49017);
nor UO_3674 (O_3674,N_48818,N_49774);
nor UO_3675 (O_3675,N_49922,N_49271);
nor UO_3676 (O_3676,N_48896,N_49590);
nor UO_3677 (O_3677,N_49898,N_48511);
nor UO_3678 (O_3678,N_49618,N_49843);
and UO_3679 (O_3679,N_48223,N_48163);
nand UO_3680 (O_3680,N_49132,N_49163);
or UO_3681 (O_3681,N_48397,N_49058);
nor UO_3682 (O_3682,N_49394,N_49320);
nand UO_3683 (O_3683,N_49212,N_49096);
or UO_3684 (O_3684,N_49112,N_48846);
and UO_3685 (O_3685,N_49247,N_49824);
or UO_3686 (O_3686,N_48128,N_48680);
or UO_3687 (O_3687,N_48933,N_49210);
or UO_3688 (O_3688,N_48312,N_48609);
xnor UO_3689 (O_3689,N_48282,N_48169);
and UO_3690 (O_3690,N_48669,N_48006);
nor UO_3691 (O_3691,N_49550,N_48983);
xnor UO_3692 (O_3692,N_48263,N_49206);
nand UO_3693 (O_3693,N_48846,N_48211);
and UO_3694 (O_3694,N_48033,N_49219);
nand UO_3695 (O_3695,N_49641,N_49757);
or UO_3696 (O_3696,N_48373,N_49672);
and UO_3697 (O_3697,N_49732,N_49425);
xnor UO_3698 (O_3698,N_48077,N_49076);
and UO_3699 (O_3699,N_49565,N_49593);
and UO_3700 (O_3700,N_48800,N_49603);
nor UO_3701 (O_3701,N_48113,N_48000);
and UO_3702 (O_3702,N_49219,N_49003);
xnor UO_3703 (O_3703,N_49379,N_49984);
nor UO_3704 (O_3704,N_48763,N_48641);
nor UO_3705 (O_3705,N_49446,N_49684);
and UO_3706 (O_3706,N_48007,N_49450);
and UO_3707 (O_3707,N_48331,N_48051);
or UO_3708 (O_3708,N_49976,N_48440);
or UO_3709 (O_3709,N_49995,N_48139);
and UO_3710 (O_3710,N_49817,N_49440);
and UO_3711 (O_3711,N_49244,N_49677);
or UO_3712 (O_3712,N_48823,N_49103);
or UO_3713 (O_3713,N_49771,N_49737);
and UO_3714 (O_3714,N_49544,N_49786);
xor UO_3715 (O_3715,N_48086,N_48889);
nor UO_3716 (O_3716,N_48019,N_49892);
xor UO_3717 (O_3717,N_48571,N_48455);
nand UO_3718 (O_3718,N_49857,N_48959);
xnor UO_3719 (O_3719,N_48462,N_48858);
and UO_3720 (O_3720,N_48243,N_49240);
nor UO_3721 (O_3721,N_49092,N_48163);
and UO_3722 (O_3722,N_49712,N_49387);
nand UO_3723 (O_3723,N_49245,N_48802);
and UO_3724 (O_3724,N_49045,N_49432);
or UO_3725 (O_3725,N_49029,N_48303);
nand UO_3726 (O_3726,N_49810,N_48023);
nor UO_3727 (O_3727,N_49319,N_48051);
and UO_3728 (O_3728,N_49071,N_48563);
xnor UO_3729 (O_3729,N_49874,N_49812);
and UO_3730 (O_3730,N_49028,N_48840);
nor UO_3731 (O_3731,N_49983,N_48696);
xnor UO_3732 (O_3732,N_49271,N_48417);
or UO_3733 (O_3733,N_48038,N_48780);
or UO_3734 (O_3734,N_49921,N_48657);
nor UO_3735 (O_3735,N_49416,N_49382);
nand UO_3736 (O_3736,N_48870,N_48641);
nor UO_3737 (O_3737,N_49149,N_49438);
nand UO_3738 (O_3738,N_49062,N_49567);
nand UO_3739 (O_3739,N_49367,N_48204);
or UO_3740 (O_3740,N_48844,N_48217);
nand UO_3741 (O_3741,N_49139,N_49381);
or UO_3742 (O_3742,N_49671,N_48942);
nand UO_3743 (O_3743,N_49910,N_48604);
nor UO_3744 (O_3744,N_48317,N_49891);
xnor UO_3745 (O_3745,N_49961,N_49599);
or UO_3746 (O_3746,N_48907,N_49131);
xor UO_3747 (O_3747,N_48874,N_48966);
nor UO_3748 (O_3748,N_48901,N_48607);
or UO_3749 (O_3749,N_49953,N_48438);
xnor UO_3750 (O_3750,N_48255,N_49161);
xor UO_3751 (O_3751,N_48516,N_49922);
xnor UO_3752 (O_3752,N_48380,N_48065);
nand UO_3753 (O_3753,N_49076,N_48731);
or UO_3754 (O_3754,N_48825,N_48244);
xor UO_3755 (O_3755,N_49914,N_49972);
xnor UO_3756 (O_3756,N_48879,N_48840);
and UO_3757 (O_3757,N_49736,N_49252);
nor UO_3758 (O_3758,N_48257,N_48442);
xnor UO_3759 (O_3759,N_48427,N_49902);
or UO_3760 (O_3760,N_49019,N_49251);
or UO_3761 (O_3761,N_49634,N_48020);
or UO_3762 (O_3762,N_49248,N_49836);
xnor UO_3763 (O_3763,N_48611,N_49240);
xnor UO_3764 (O_3764,N_48080,N_49946);
or UO_3765 (O_3765,N_49760,N_48977);
and UO_3766 (O_3766,N_49112,N_48423);
nor UO_3767 (O_3767,N_49222,N_49006);
and UO_3768 (O_3768,N_49395,N_48360);
and UO_3769 (O_3769,N_48553,N_48175);
xnor UO_3770 (O_3770,N_49093,N_49290);
xor UO_3771 (O_3771,N_48934,N_48950);
nand UO_3772 (O_3772,N_49626,N_49038);
or UO_3773 (O_3773,N_49848,N_49367);
and UO_3774 (O_3774,N_48773,N_49838);
xnor UO_3775 (O_3775,N_49481,N_48793);
xor UO_3776 (O_3776,N_49858,N_49034);
nand UO_3777 (O_3777,N_48303,N_48237);
xor UO_3778 (O_3778,N_49533,N_49747);
and UO_3779 (O_3779,N_49593,N_48559);
and UO_3780 (O_3780,N_48677,N_48146);
xor UO_3781 (O_3781,N_49313,N_48668);
xnor UO_3782 (O_3782,N_48602,N_49034);
nor UO_3783 (O_3783,N_49484,N_49871);
nand UO_3784 (O_3784,N_48839,N_49000);
and UO_3785 (O_3785,N_49182,N_48570);
nor UO_3786 (O_3786,N_49023,N_49280);
nand UO_3787 (O_3787,N_49014,N_48022);
nor UO_3788 (O_3788,N_49077,N_49622);
and UO_3789 (O_3789,N_49162,N_49287);
or UO_3790 (O_3790,N_49377,N_49331);
xnor UO_3791 (O_3791,N_49562,N_48064);
and UO_3792 (O_3792,N_48910,N_49469);
or UO_3793 (O_3793,N_49972,N_49813);
or UO_3794 (O_3794,N_48694,N_49859);
xor UO_3795 (O_3795,N_49776,N_48704);
nand UO_3796 (O_3796,N_48747,N_49899);
nand UO_3797 (O_3797,N_48066,N_49138);
or UO_3798 (O_3798,N_49154,N_49165);
nand UO_3799 (O_3799,N_49591,N_49910);
nor UO_3800 (O_3800,N_48578,N_48623);
nor UO_3801 (O_3801,N_49328,N_49300);
or UO_3802 (O_3802,N_49318,N_48590);
nand UO_3803 (O_3803,N_49356,N_48048);
or UO_3804 (O_3804,N_49621,N_48109);
xnor UO_3805 (O_3805,N_48668,N_49607);
nand UO_3806 (O_3806,N_48986,N_49488);
xnor UO_3807 (O_3807,N_48449,N_49764);
nor UO_3808 (O_3808,N_48499,N_49521);
and UO_3809 (O_3809,N_49225,N_49527);
or UO_3810 (O_3810,N_48785,N_48723);
nand UO_3811 (O_3811,N_49799,N_49117);
xnor UO_3812 (O_3812,N_49101,N_48811);
nor UO_3813 (O_3813,N_48011,N_49481);
xnor UO_3814 (O_3814,N_48054,N_49487);
xnor UO_3815 (O_3815,N_49412,N_49850);
nand UO_3816 (O_3816,N_48796,N_49292);
xor UO_3817 (O_3817,N_49047,N_49900);
xor UO_3818 (O_3818,N_48946,N_49335);
or UO_3819 (O_3819,N_49545,N_49847);
xnor UO_3820 (O_3820,N_49309,N_48256);
or UO_3821 (O_3821,N_49592,N_49387);
xor UO_3822 (O_3822,N_48112,N_49119);
and UO_3823 (O_3823,N_48025,N_49407);
nand UO_3824 (O_3824,N_48031,N_48843);
or UO_3825 (O_3825,N_49135,N_49834);
or UO_3826 (O_3826,N_49457,N_49259);
or UO_3827 (O_3827,N_48494,N_49702);
xor UO_3828 (O_3828,N_49907,N_49751);
xnor UO_3829 (O_3829,N_49700,N_49660);
nand UO_3830 (O_3830,N_48753,N_49295);
nand UO_3831 (O_3831,N_48375,N_48940);
xor UO_3832 (O_3832,N_48769,N_49438);
and UO_3833 (O_3833,N_48072,N_48343);
xor UO_3834 (O_3834,N_48708,N_48992);
or UO_3835 (O_3835,N_48252,N_48655);
nand UO_3836 (O_3836,N_49352,N_48386);
nor UO_3837 (O_3837,N_49155,N_48811);
nor UO_3838 (O_3838,N_49028,N_48606);
xnor UO_3839 (O_3839,N_49940,N_49347);
nor UO_3840 (O_3840,N_49467,N_48148);
or UO_3841 (O_3841,N_48706,N_48192);
xnor UO_3842 (O_3842,N_48270,N_49240);
or UO_3843 (O_3843,N_48962,N_48433);
and UO_3844 (O_3844,N_48032,N_49060);
xor UO_3845 (O_3845,N_49373,N_48084);
and UO_3846 (O_3846,N_49383,N_48011);
or UO_3847 (O_3847,N_49023,N_49733);
and UO_3848 (O_3848,N_48481,N_48784);
nor UO_3849 (O_3849,N_49636,N_48071);
xor UO_3850 (O_3850,N_49919,N_48204);
and UO_3851 (O_3851,N_49885,N_49084);
or UO_3852 (O_3852,N_48371,N_48422);
and UO_3853 (O_3853,N_49422,N_49567);
or UO_3854 (O_3854,N_49757,N_48860);
nand UO_3855 (O_3855,N_49423,N_48699);
and UO_3856 (O_3856,N_48182,N_49937);
nor UO_3857 (O_3857,N_49137,N_48539);
or UO_3858 (O_3858,N_48412,N_49402);
nand UO_3859 (O_3859,N_48088,N_49331);
or UO_3860 (O_3860,N_49765,N_49560);
and UO_3861 (O_3861,N_48285,N_49757);
or UO_3862 (O_3862,N_49418,N_49824);
and UO_3863 (O_3863,N_49386,N_48429);
nand UO_3864 (O_3864,N_49991,N_49965);
nor UO_3865 (O_3865,N_48305,N_49084);
nand UO_3866 (O_3866,N_49090,N_48910);
nor UO_3867 (O_3867,N_48676,N_48386);
nand UO_3868 (O_3868,N_48322,N_48104);
or UO_3869 (O_3869,N_49864,N_49544);
or UO_3870 (O_3870,N_49067,N_48362);
or UO_3871 (O_3871,N_48919,N_48865);
nor UO_3872 (O_3872,N_48565,N_48033);
nand UO_3873 (O_3873,N_49504,N_49491);
nor UO_3874 (O_3874,N_49051,N_49276);
xor UO_3875 (O_3875,N_48629,N_48286);
or UO_3876 (O_3876,N_49300,N_48436);
nor UO_3877 (O_3877,N_48653,N_48604);
or UO_3878 (O_3878,N_49068,N_48313);
and UO_3879 (O_3879,N_48860,N_48610);
nand UO_3880 (O_3880,N_48065,N_48995);
or UO_3881 (O_3881,N_48798,N_48669);
xor UO_3882 (O_3882,N_48315,N_48575);
nor UO_3883 (O_3883,N_49963,N_48472);
xor UO_3884 (O_3884,N_48340,N_49990);
or UO_3885 (O_3885,N_48064,N_48600);
nor UO_3886 (O_3886,N_48413,N_48035);
nand UO_3887 (O_3887,N_48706,N_48266);
xor UO_3888 (O_3888,N_48954,N_48568);
nor UO_3889 (O_3889,N_49036,N_48870);
or UO_3890 (O_3890,N_48674,N_48816);
nand UO_3891 (O_3891,N_49214,N_49132);
or UO_3892 (O_3892,N_48778,N_49079);
and UO_3893 (O_3893,N_49444,N_49953);
nor UO_3894 (O_3894,N_49905,N_48107);
nor UO_3895 (O_3895,N_48182,N_48110);
and UO_3896 (O_3896,N_48536,N_49933);
xor UO_3897 (O_3897,N_49914,N_48382);
nand UO_3898 (O_3898,N_49535,N_48553);
xnor UO_3899 (O_3899,N_48518,N_49489);
and UO_3900 (O_3900,N_48095,N_49313);
xor UO_3901 (O_3901,N_48980,N_49105);
xor UO_3902 (O_3902,N_48955,N_48027);
nand UO_3903 (O_3903,N_48847,N_48483);
xor UO_3904 (O_3904,N_49187,N_49735);
or UO_3905 (O_3905,N_48951,N_49447);
or UO_3906 (O_3906,N_48441,N_49631);
xnor UO_3907 (O_3907,N_48776,N_48522);
nor UO_3908 (O_3908,N_48076,N_48793);
nor UO_3909 (O_3909,N_49497,N_48068);
and UO_3910 (O_3910,N_48723,N_49933);
nor UO_3911 (O_3911,N_48045,N_49930);
nor UO_3912 (O_3912,N_48311,N_49063);
or UO_3913 (O_3913,N_49789,N_49524);
or UO_3914 (O_3914,N_49895,N_49532);
xnor UO_3915 (O_3915,N_49688,N_48271);
and UO_3916 (O_3916,N_48451,N_49428);
nand UO_3917 (O_3917,N_48358,N_48447);
nor UO_3918 (O_3918,N_49289,N_48469);
nand UO_3919 (O_3919,N_49374,N_49615);
xnor UO_3920 (O_3920,N_49476,N_48593);
or UO_3921 (O_3921,N_48738,N_48807);
xor UO_3922 (O_3922,N_48916,N_49894);
and UO_3923 (O_3923,N_48194,N_49364);
xor UO_3924 (O_3924,N_49377,N_48138);
or UO_3925 (O_3925,N_49238,N_49380);
xor UO_3926 (O_3926,N_49015,N_48086);
and UO_3927 (O_3927,N_48199,N_49489);
or UO_3928 (O_3928,N_49067,N_49323);
nand UO_3929 (O_3929,N_49119,N_49323);
and UO_3930 (O_3930,N_48138,N_49320);
and UO_3931 (O_3931,N_48829,N_48878);
or UO_3932 (O_3932,N_49603,N_48602);
xor UO_3933 (O_3933,N_48791,N_48566);
nor UO_3934 (O_3934,N_48433,N_48773);
or UO_3935 (O_3935,N_48817,N_49358);
and UO_3936 (O_3936,N_48876,N_49716);
nand UO_3937 (O_3937,N_49764,N_48912);
xor UO_3938 (O_3938,N_49453,N_48676);
xor UO_3939 (O_3939,N_49610,N_49893);
nor UO_3940 (O_3940,N_49779,N_49163);
xnor UO_3941 (O_3941,N_48524,N_48515);
xnor UO_3942 (O_3942,N_48204,N_48775);
and UO_3943 (O_3943,N_49602,N_49471);
or UO_3944 (O_3944,N_48355,N_48193);
xor UO_3945 (O_3945,N_49692,N_49754);
and UO_3946 (O_3946,N_49496,N_49536);
and UO_3947 (O_3947,N_48542,N_49879);
or UO_3948 (O_3948,N_48106,N_49663);
nor UO_3949 (O_3949,N_48984,N_49918);
nand UO_3950 (O_3950,N_49875,N_49571);
nor UO_3951 (O_3951,N_49093,N_49964);
nor UO_3952 (O_3952,N_48805,N_49548);
nor UO_3953 (O_3953,N_49925,N_49094);
or UO_3954 (O_3954,N_49440,N_48151);
xnor UO_3955 (O_3955,N_48877,N_48504);
and UO_3956 (O_3956,N_48248,N_48499);
nor UO_3957 (O_3957,N_48906,N_49045);
or UO_3958 (O_3958,N_49431,N_48609);
nand UO_3959 (O_3959,N_48470,N_48985);
xor UO_3960 (O_3960,N_49568,N_49545);
xnor UO_3961 (O_3961,N_48161,N_49985);
nor UO_3962 (O_3962,N_49590,N_49662);
or UO_3963 (O_3963,N_49277,N_49643);
or UO_3964 (O_3964,N_49544,N_48356);
or UO_3965 (O_3965,N_49301,N_49594);
and UO_3966 (O_3966,N_49537,N_48638);
nand UO_3967 (O_3967,N_48073,N_48435);
nand UO_3968 (O_3968,N_48210,N_48559);
xor UO_3969 (O_3969,N_48980,N_49379);
nor UO_3970 (O_3970,N_48285,N_48156);
nand UO_3971 (O_3971,N_49202,N_49641);
nor UO_3972 (O_3972,N_48807,N_49751);
xor UO_3973 (O_3973,N_48711,N_48111);
nor UO_3974 (O_3974,N_49897,N_48027);
or UO_3975 (O_3975,N_49888,N_49905);
and UO_3976 (O_3976,N_49055,N_48338);
or UO_3977 (O_3977,N_48960,N_48646);
nor UO_3978 (O_3978,N_48757,N_48273);
xnor UO_3979 (O_3979,N_48659,N_48884);
or UO_3980 (O_3980,N_48453,N_48062);
or UO_3981 (O_3981,N_49188,N_49787);
and UO_3982 (O_3982,N_49892,N_48921);
nor UO_3983 (O_3983,N_48856,N_49631);
and UO_3984 (O_3984,N_49452,N_48015);
nor UO_3985 (O_3985,N_48946,N_49367);
and UO_3986 (O_3986,N_49002,N_48330);
or UO_3987 (O_3987,N_48562,N_48833);
xor UO_3988 (O_3988,N_49168,N_49513);
xor UO_3989 (O_3989,N_49380,N_49938);
or UO_3990 (O_3990,N_48392,N_49419);
nand UO_3991 (O_3991,N_49042,N_48178);
and UO_3992 (O_3992,N_48556,N_48630);
xnor UO_3993 (O_3993,N_48406,N_48507);
xnor UO_3994 (O_3994,N_49772,N_49371);
nand UO_3995 (O_3995,N_48774,N_49694);
nor UO_3996 (O_3996,N_49729,N_48597);
or UO_3997 (O_3997,N_49694,N_49998);
nand UO_3998 (O_3998,N_48751,N_49038);
or UO_3999 (O_3999,N_48110,N_48716);
or UO_4000 (O_4000,N_49480,N_48692);
or UO_4001 (O_4001,N_48179,N_48202);
and UO_4002 (O_4002,N_49654,N_48032);
nor UO_4003 (O_4003,N_48644,N_49440);
or UO_4004 (O_4004,N_48473,N_49090);
and UO_4005 (O_4005,N_48184,N_49478);
xor UO_4006 (O_4006,N_49103,N_48779);
xnor UO_4007 (O_4007,N_48017,N_48468);
xor UO_4008 (O_4008,N_48164,N_48528);
nor UO_4009 (O_4009,N_48532,N_48045);
or UO_4010 (O_4010,N_48521,N_48532);
nor UO_4011 (O_4011,N_48402,N_49349);
nand UO_4012 (O_4012,N_48630,N_48688);
xor UO_4013 (O_4013,N_49840,N_48392);
and UO_4014 (O_4014,N_48509,N_48377);
and UO_4015 (O_4015,N_49170,N_49937);
or UO_4016 (O_4016,N_49723,N_49292);
nor UO_4017 (O_4017,N_48618,N_49463);
or UO_4018 (O_4018,N_49138,N_49448);
nand UO_4019 (O_4019,N_48346,N_49244);
xor UO_4020 (O_4020,N_48912,N_48578);
nand UO_4021 (O_4021,N_49989,N_49502);
nor UO_4022 (O_4022,N_49335,N_48661);
or UO_4023 (O_4023,N_48908,N_48423);
and UO_4024 (O_4024,N_48320,N_48184);
nand UO_4025 (O_4025,N_49216,N_48627);
nand UO_4026 (O_4026,N_48941,N_49253);
nor UO_4027 (O_4027,N_48305,N_48466);
nor UO_4028 (O_4028,N_48381,N_49040);
xor UO_4029 (O_4029,N_48636,N_48280);
or UO_4030 (O_4030,N_49168,N_48469);
nand UO_4031 (O_4031,N_49173,N_49304);
xnor UO_4032 (O_4032,N_49294,N_49456);
nor UO_4033 (O_4033,N_49552,N_48793);
nand UO_4034 (O_4034,N_49355,N_48444);
and UO_4035 (O_4035,N_49900,N_48966);
and UO_4036 (O_4036,N_48887,N_48983);
xor UO_4037 (O_4037,N_49490,N_49777);
and UO_4038 (O_4038,N_49761,N_49005);
xor UO_4039 (O_4039,N_48434,N_49468);
or UO_4040 (O_4040,N_49551,N_49315);
nor UO_4041 (O_4041,N_48217,N_49515);
and UO_4042 (O_4042,N_49224,N_48606);
nand UO_4043 (O_4043,N_49249,N_48517);
and UO_4044 (O_4044,N_48767,N_48804);
nand UO_4045 (O_4045,N_48661,N_49799);
and UO_4046 (O_4046,N_49755,N_48048);
or UO_4047 (O_4047,N_49194,N_48096);
and UO_4048 (O_4048,N_48824,N_48305);
nor UO_4049 (O_4049,N_48180,N_48195);
and UO_4050 (O_4050,N_49586,N_49807);
nand UO_4051 (O_4051,N_49376,N_48181);
nor UO_4052 (O_4052,N_48925,N_49858);
nor UO_4053 (O_4053,N_49885,N_49703);
and UO_4054 (O_4054,N_49903,N_48519);
or UO_4055 (O_4055,N_48521,N_48207);
nand UO_4056 (O_4056,N_49286,N_48510);
and UO_4057 (O_4057,N_49826,N_49867);
nor UO_4058 (O_4058,N_48006,N_49765);
nor UO_4059 (O_4059,N_48827,N_48762);
xnor UO_4060 (O_4060,N_48311,N_49933);
xor UO_4061 (O_4061,N_49012,N_48229);
nand UO_4062 (O_4062,N_49923,N_49163);
or UO_4063 (O_4063,N_48864,N_49095);
or UO_4064 (O_4064,N_49160,N_49901);
or UO_4065 (O_4065,N_49918,N_48735);
nand UO_4066 (O_4066,N_48751,N_48522);
or UO_4067 (O_4067,N_49260,N_49661);
nor UO_4068 (O_4068,N_49520,N_48415);
and UO_4069 (O_4069,N_48910,N_48182);
or UO_4070 (O_4070,N_49361,N_49924);
nor UO_4071 (O_4071,N_48103,N_49267);
xnor UO_4072 (O_4072,N_48684,N_49153);
and UO_4073 (O_4073,N_48612,N_48095);
nor UO_4074 (O_4074,N_49955,N_49681);
nand UO_4075 (O_4075,N_48487,N_49991);
nor UO_4076 (O_4076,N_48361,N_48995);
nand UO_4077 (O_4077,N_49957,N_48551);
and UO_4078 (O_4078,N_49358,N_49414);
or UO_4079 (O_4079,N_48032,N_49007);
nor UO_4080 (O_4080,N_48720,N_49232);
nor UO_4081 (O_4081,N_48560,N_49144);
nand UO_4082 (O_4082,N_49254,N_49248);
nand UO_4083 (O_4083,N_48629,N_49559);
nand UO_4084 (O_4084,N_49743,N_49383);
xor UO_4085 (O_4085,N_48436,N_48562);
xnor UO_4086 (O_4086,N_49901,N_48801);
and UO_4087 (O_4087,N_48869,N_48236);
or UO_4088 (O_4088,N_49326,N_48690);
or UO_4089 (O_4089,N_48110,N_48063);
or UO_4090 (O_4090,N_49808,N_49912);
or UO_4091 (O_4091,N_49777,N_49896);
nand UO_4092 (O_4092,N_49383,N_48231);
nor UO_4093 (O_4093,N_48764,N_49047);
or UO_4094 (O_4094,N_49606,N_48051);
xnor UO_4095 (O_4095,N_49769,N_48271);
nor UO_4096 (O_4096,N_49037,N_48639);
or UO_4097 (O_4097,N_48046,N_48266);
xnor UO_4098 (O_4098,N_49595,N_48577);
or UO_4099 (O_4099,N_48052,N_48800);
xnor UO_4100 (O_4100,N_49684,N_49500);
xor UO_4101 (O_4101,N_49513,N_48622);
nor UO_4102 (O_4102,N_49492,N_49305);
xnor UO_4103 (O_4103,N_49951,N_49753);
nand UO_4104 (O_4104,N_49064,N_48248);
or UO_4105 (O_4105,N_49313,N_48183);
and UO_4106 (O_4106,N_49013,N_48568);
xnor UO_4107 (O_4107,N_48878,N_49135);
and UO_4108 (O_4108,N_48869,N_48811);
nand UO_4109 (O_4109,N_49311,N_49394);
xnor UO_4110 (O_4110,N_48862,N_48647);
nand UO_4111 (O_4111,N_49561,N_49109);
nor UO_4112 (O_4112,N_48321,N_49561);
xor UO_4113 (O_4113,N_48684,N_48959);
nand UO_4114 (O_4114,N_49272,N_49156);
nand UO_4115 (O_4115,N_48916,N_49441);
and UO_4116 (O_4116,N_48224,N_48894);
nor UO_4117 (O_4117,N_49348,N_48705);
and UO_4118 (O_4118,N_48470,N_48870);
xnor UO_4119 (O_4119,N_48653,N_48881);
xor UO_4120 (O_4120,N_49376,N_48418);
or UO_4121 (O_4121,N_48261,N_48182);
or UO_4122 (O_4122,N_49380,N_48131);
nor UO_4123 (O_4123,N_49017,N_49487);
xnor UO_4124 (O_4124,N_49795,N_49332);
nor UO_4125 (O_4125,N_49490,N_49963);
or UO_4126 (O_4126,N_49241,N_48325);
nand UO_4127 (O_4127,N_49643,N_49728);
xor UO_4128 (O_4128,N_48087,N_48945);
and UO_4129 (O_4129,N_48603,N_49512);
nand UO_4130 (O_4130,N_49302,N_48435);
xnor UO_4131 (O_4131,N_49057,N_48769);
nand UO_4132 (O_4132,N_48674,N_48070);
nor UO_4133 (O_4133,N_48737,N_48529);
nor UO_4134 (O_4134,N_49894,N_48412);
or UO_4135 (O_4135,N_48626,N_49655);
nand UO_4136 (O_4136,N_48844,N_48725);
nand UO_4137 (O_4137,N_48789,N_49980);
xnor UO_4138 (O_4138,N_48398,N_48796);
xor UO_4139 (O_4139,N_48065,N_48996);
and UO_4140 (O_4140,N_49120,N_48978);
or UO_4141 (O_4141,N_48405,N_49522);
xor UO_4142 (O_4142,N_49724,N_48498);
or UO_4143 (O_4143,N_49827,N_49780);
nand UO_4144 (O_4144,N_48692,N_49097);
or UO_4145 (O_4145,N_49178,N_48014);
and UO_4146 (O_4146,N_48871,N_49368);
or UO_4147 (O_4147,N_49723,N_48651);
or UO_4148 (O_4148,N_48608,N_48162);
or UO_4149 (O_4149,N_48724,N_48861);
or UO_4150 (O_4150,N_49216,N_49855);
xor UO_4151 (O_4151,N_48957,N_48831);
and UO_4152 (O_4152,N_48969,N_48412);
nor UO_4153 (O_4153,N_49150,N_48669);
and UO_4154 (O_4154,N_48022,N_49695);
nor UO_4155 (O_4155,N_49525,N_49747);
and UO_4156 (O_4156,N_49635,N_48286);
and UO_4157 (O_4157,N_49604,N_49384);
xor UO_4158 (O_4158,N_49253,N_48598);
xnor UO_4159 (O_4159,N_48689,N_48709);
xnor UO_4160 (O_4160,N_49767,N_48967);
and UO_4161 (O_4161,N_49302,N_49645);
xor UO_4162 (O_4162,N_48038,N_49021);
or UO_4163 (O_4163,N_48217,N_48605);
and UO_4164 (O_4164,N_48319,N_48371);
nand UO_4165 (O_4165,N_49646,N_48238);
or UO_4166 (O_4166,N_48401,N_49013);
or UO_4167 (O_4167,N_49461,N_49793);
or UO_4168 (O_4168,N_49235,N_49814);
nand UO_4169 (O_4169,N_49411,N_49726);
or UO_4170 (O_4170,N_49026,N_49522);
or UO_4171 (O_4171,N_49505,N_48746);
nand UO_4172 (O_4172,N_48211,N_49278);
xnor UO_4173 (O_4173,N_48331,N_48465);
or UO_4174 (O_4174,N_48079,N_49120);
nand UO_4175 (O_4175,N_48731,N_48889);
nand UO_4176 (O_4176,N_48071,N_49596);
or UO_4177 (O_4177,N_49215,N_48728);
and UO_4178 (O_4178,N_49911,N_48928);
nor UO_4179 (O_4179,N_48742,N_48330);
nand UO_4180 (O_4180,N_49829,N_49841);
xor UO_4181 (O_4181,N_49716,N_49785);
or UO_4182 (O_4182,N_48770,N_49122);
or UO_4183 (O_4183,N_48505,N_48646);
nor UO_4184 (O_4184,N_49863,N_48877);
nand UO_4185 (O_4185,N_49101,N_48847);
nor UO_4186 (O_4186,N_48034,N_48746);
xnor UO_4187 (O_4187,N_49681,N_48814);
xor UO_4188 (O_4188,N_48344,N_48782);
xor UO_4189 (O_4189,N_49780,N_49578);
xor UO_4190 (O_4190,N_49198,N_48783);
nor UO_4191 (O_4191,N_48820,N_48585);
and UO_4192 (O_4192,N_48196,N_48557);
nor UO_4193 (O_4193,N_49220,N_49070);
nor UO_4194 (O_4194,N_49389,N_49630);
xnor UO_4195 (O_4195,N_49102,N_49295);
nor UO_4196 (O_4196,N_49083,N_49056);
xor UO_4197 (O_4197,N_48223,N_49813);
or UO_4198 (O_4198,N_49725,N_48254);
nand UO_4199 (O_4199,N_48880,N_48541);
nor UO_4200 (O_4200,N_49641,N_48584);
nor UO_4201 (O_4201,N_48027,N_48638);
xnor UO_4202 (O_4202,N_49021,N_49113);
or UO_4203 (O_4203,N_48254,N_49359);
nand UO_4204 (O_4204,N_48992,N_49839);
nor UO_4205 (O_4205,N_49207,N_48939);
or UO_4206 (O_4206,N_49013,N_49452);
nand UO_4207 (O_4207,N_48518,N_48858);
nor UO_4208 (O_4208,N_49118,N_49029);
xor UO_4209 (O_4209,N_49895,N_49129);
nor UO_4210 (O_4210,N_49909,N_48923);
nor UO_4211 (O_4211,N_48875,N_49871);
nand UO_4212 (O_4212,N_49452,N_48004);
or UO_4213 (O_4213,N_48890,N_49276);
nand UO_4214 (O_4214,N_48893,N_48450);
xor UO_4215 (O_4215,N_48747,N_48180);
or UO_4216 (O_4216,N_48081,N_49472);
and UO_4217 (O_4217,N_48314,N_49289);
or UO_4218 (O_4218,N_49656,N_49025);
or UO_4219 (O_4219,N_48173,N_49461);
and UO_4220 (O_4220,N_48380,N_49835);
nand UO_4221 (O_4221,N_49418,N_48445);
nor UO_4222 (O_4222,N_48686,N_48542);
xnor UO_4223 (O_4223,N_49704,N_49864);
nor UO_4224 (O_4224,N_48933,N_48127);
or UO_4225 (O_4225,N_49891,N_49101);
nand UO_4226 (O_4226,N_48757,N_48694);
and UO_4227 (O_4227,N_49628,N_48637);
nor UO_4228 (O_4228,N_49593,N_49010);
and UO_4229 (O_4229,N_48651,N_49104);
xor UO_4230 (O_4230,N_48980,N_48933);
xor UO_4231 (O_4231,N_48183,N_48239);
or UO_4232 (O_4232,N_49740,N_49475);
or UO_4233 (O_4233,N_49721,N_48819);
nand UO_4234 (O_4234,N_48540,N_48589);
nor UO_4235 (O_4235,N_48558,N_48274);
or UO_4236 (O_4236,N_48234,N_49671);
nor UO_4237 (O_4237,N_48807,N_48872);
or UO_4238 (O_4238,N_49850,N_49121);
nor UO_4239 (O_4239,N_49744,N_49206);
or UO_4240 (O_4240,N_48279,N_49921);
nor UO_4241 (O_4241,N_48220,N_48581);
and UO_4242 (O_4242,N_49872,N_49732);
nor UO_4243 (O_4243,N_48274,N_48245);
nand UO_4244 (O_4244,N_49541,N_48772);
nor UO_4245 (O_4245,N_48633,N_49640);
and UO_4246 (O_4246,N_49204,N_48904);
nor UO_4247 (O_4247,N_48047,N_48675);
or UO_4248 (O_4248,N_49564,N_48287);
nor UO_4249 (O_4249,N_48137,N_49329);
and UO_4250 (O_4250,N_49084,N_48704);
xnor UO_4251 (O_4251,N_48140,N_49205);
nor UO_4252 (O_4252,N_49546,N_48831);
nor UO_4253 (O_4253,N_48619,N_48457);
xor UO_4254 (O_4254,N_48480,N_49370);
or UO_4255 (O_4255,N_48977,N_49200);
and UO_4256 (O_4256,N_49410,N_49447);
nor UO_4257 (O_4257,N_49462,N_49854);
or UO_4258 (O_4258,N_49011,N_49727);
nand UO_4259 (O_4259,N_49903,N_49346);
or UO_4260 (O_4260,N_48262,N_49136);
nor UO_4261 (O_4261,N_49857,N_48865);
nand UO_4262 (O_4262,N_48150,N_49375);
nand UO_4263 (O_4263,N_48398,N_49126);
xnor UO_4264 (O_4264,N_49332,N_48755);
xnor UO_4265 (O_4265,N_49098,N_49055);
xnor UO_4266 (O_4266,N_48797,N_48003);
nor UO_4267 (O_4267,N_48922,N_48099);
xor UO_4268 (O_4268,N_49566,N_49301);
xor UO_4269 (O_4269,N_49087,N_49050);
or UO_4270 (O_4270,N_49199,N_49647);
nand UO_4271 (O_4271,N_48778,N_49344);
nor UO_4272 (O_4272,N_49751,N_48181);
xnor UO_4273 (O_4273,N_48884,N_48203);
nand UO_4274 (O_4274,N_49101,N_49563);
and UO_4275 (O_4275,N_48600,N_48584);
and UO_4276 (O_4276,N_49456,N_48119);
nor UO_4277 (O_4277,N_49906,N_49631);
or UO_4278 (O_4278,N_48270,N_48194);
nor UO_4279 (O_4279,N_48317,N_49025);
nand UO_4280 (O_4280,N_49772,N_48288);
nor UO_4281 (O_4281,N_49643,N_49832);
or UO_4282 (O_4282,N_48938,N_49654);
xnor UO_4283 (O_4283,N_48163,N_49101);
and UO_4284 (O_4284,N_48129,N_49102);
or UO_4285 (O_4285,N_49153,N_48036);
xor UO_4286 (O_4286,N_48548,N_49396);
xor UO_4287 (O_4287,N_48576,N_49773);
xnor UO_4288 (O_4288,N_49811,N_48044);
or UO_4289 (O_4289,N_49483,N_49375);
and UO_4290 (O_4290,N_48639,N_48393);
xnor UO_4291 (O_4291,N_48627,N_48326);
nand UO_4292 (O_4292,N_48473,N_49834);
xor UO_4293 (O_4293,N_48748,N_49137);
and UO_4294 (O_4294,N_49809,N_48605);
nor UO_4295 (O_4295,N_49656,N_49499);
or UO_4296 (O_4296,N_48093,N_48919);
nand UO_4297 (O_4297,N_49579,N_49418);
xor UO_4298 (O_4298,N_49905,N_49436);
xnor UO_4299 (O_4299,N_48117,N_48874);
nand UO_4300 (O_4300,N_49574,N_48822);
and UO_4301 (O_4301,N_48241,N_48783);
nand UO_4302 (O_4302,N_48568,N_49947);
or UO_4303 (O_4303,N_49383,N_48983);
nor UO_4304 (O_4304,N_49730,N_49633);
nor UO_4305 (O_4305,N_48160,N_49826);
nor UO_4306 (O_4306,N_49423,N_49737);
or UO_4307 (O_4307,N_49567,N_49722);
and UO_4308 (O_4308,N_48174,N_48460);
and UO_4309 (O_4309,N_49673,N_49973);
nor UO_4310 (O_4310,N_49161,N_48744);
xor UO_4311 (O_4311,N_48548,N_48925);
xor UO_4312 (O_4312,N_49358,N_49452);
or UO_4313 (O_4313,N_48111,N_49836);
or UO_4314 (O_4314,N_48079,N_48086);
and UO_4315 (O_4315,N_48304,N_48987);
nor UO_4316 (O_4316,N_49716,N_49768);
nor UO_4317 (O_4317,N_48827,N_49263);
or UO_4318 (O_4318,N_49094,N_48783);
and UO_4319 (O_4319,N_49643,N_49492);
nor UO_4320 (O_4320,N_49521,N_48676);
and UO_4321 (O_4321,N_48127,N_48107);
or UO_4322 (O_4322,N_49524,N_49890);
nor UO_4323 (O_4323,N_49124,N_49634);
xnor UO_4324 (O_4324,N_48108,N_48209);
xnor UO_4325 (O_4325,N_49881,N_49879);
nand UO_4326 (O_4326,N_49106,N_48531);
nor UO_4327 (O_4327,N_49532,N_48023);
and UO_4328 (O_4328,N_49305,N_49726);
or UO_4329 (O_4329,N_49869,N_49167);
and UO_4330 (O_4330,N_49702,N_48203);
and UO_4331 (O_4331,N_49970,N_49113);
or UO_4332 (O_4332,N_49380,N_49589);
and UO_4333 (O_4333,N_48327,N_48126);
or UO_4334 (O_4334,N_48557,N_48764);
nand UO_4335 (O_4335,N_48992,N_49540);
nand UO_4336 (O_4336,N_48083,N_49400);
nand UO_4337 (O_4337,N_48273,N_48268);
and UO_4338 (O_4338,N_49286,N_48211);
nand UO_4339 (O_4339,N_49313,N_49835);
nor UO_4340 (O_4340,N_49629,N_49800);
or UO_4341 (O_4341,N_49121,N_49006);
nor UO_4342 (O_4342,N_48812,N_48316);
and UO_4343 (O_4343,N_48787,N_49617);
nor UO_4344 (O_4344,N_48720,N_48465);
xnor UO_4345 (O_4345,N_48952,N_49999);
or UO_4346 (O_4346,N_48767,N_48187);
nand UO_4347 (O_4347,N_48054,N_49738);
xnor UO_4348 (O_4348,N_48144,N_49412);
and UO_4349 (O_4349,N_49871,N_48228);
nand UO_4350 (O_4350,N_48173,N_48322);
xor UO_4351 (O_4351,N_48055,N_48315);
nand UO_4352 (O_4352,N_49351,N_48868);
nand UO_4353 (O_4353,N_48301,N_48056);
nor UO_4354 (O_4354,N_48108,N_49644);
and UO_4355 (O_4355,N_48365,N_49427);
nand UO_4356 (O_4356,N_48092,N_49930);
and UO_4357 (O_4357,N_49063,N_48099);
nand UO_4358 (O_4358,N_49266,N_49836);
or UO_4359 (O_4359,N_49405,N_48728);
xnor UO_4360 (O_4360,N_49921,N_49125);
and UO_4361 (O_4361,N_48011,N_49414);
nand UO_4362 (O_4362,N_49779,N_48572);
xor UO_4363 (O_4363,N_48911,N_48899);
xor UO_4364 (O_4364,N_48059,N_49900);
nand UO_4365 (O_4365,N_48341,N_48997);
xnor UO_4366 (O_4366,N_49271,N_49213);
and UO_4367 (O_4367,N_49268,N_49883);
and UO_4368 (O_4368,N_49505,N_48514);
nor UO_4369 (O_4369,N_48855,N_48723);
or UO_4370 (O_4370,N_49240,N_48372);
nand UO_4371 (O_4371,N_48249,N_49413);
nand UO_4372 (O_4372,N_48589,N_48709);
nor UO_4373 (O_4373,N_49447,N_48650);
and UO_4374 (O_4374,N_48498,N_48216);
or UO_4375 (O_4375,N_49361,N_49650);
nor UO_4376 (O_4376,N_48680,N_48309);
nor UO_4377 (O_4377,N_48535,N_48254);
nor UO_4378 (O_4378,N_48051,N_48599);
xor UO_4379 (O_4379,N_49424,N_48755);
nor UO_4380 (O_4380,N_48625,N_48414);
xnor UO_4381 (O_4381,N_49934,N_49993);
or UO_4382 (O_4382,N_49838,N_49722);
or UO_4383 (O_4383,N_48198,N_49140);
and UO_4384 (O_4384,N_49888,N_48429);
or UO_4385 (O_4385,N_49586,N_49034);
or UO_4386 (O_4386,N_49646,N_48973);
nor UO_4387 (O_4387,N_48557,N_49347);
xor UO_4388 (O_4388,N_49826,N_48216);
or UO_4389 (O_4389,N_49397,N_48306);
nand UO_4390 (O_4390,N_49063,N_48032);
nand UO_4391 (O_4391,N_49569,N_48015);
or UO_4392 (O_4392,N_49541,N_48731);
nand UO_4393 (O_4393,N_49119,N_49898);
or UO_4394 (O_4394,N_49858,N_48348);
nand UO_4395 (O_4395,N_49741,N_49630);
and UO_4396 (O_4396,N_48102,N_48610);
nand UO_4397 (O_4397,N_48675,N_48447);
nor UO_4398 (O_4398,N_49952,N_48463);
nor UO_4399 (O_4399,N_49229,N_49283);
or UO_4400 (O_4400,N_49483,N_49236);
and UO_4401 (O_4401,N_49725,N_49312);
nand UO_4402 (O_4402,N_49597,N_48371);
nor UO_4403 (O_4403,N_49788,N_48814);
xnor UO_4404 (O_4404,N_48954,N_48413);
and UO_4405 (O_4405,N_49154,N_49083);
nand UO_4406 (O_4406,N_48138,N_48083);
and UO_4407 (O_4407,N_49409,N_49401);
nor UO_4408 (O_4408,N_49642,N_49400);
and UO_4409 (O_4409,N_49505,N_48697);
nand UO_4410 (O_4410,N_49198,N_48911);
nor UO_4411 (O_4411,N_49123,N_49357);
nor UO_4412 (O_4412,N_48266,N_49885);
and UO_4413 (O_4413,N_49489,N_49339);
nand UO_4414 (O_4414,N_48018,N_49259);
nor UO_4415 (O_4415,N_48712,N_48861);
and UO_4416 (O_4416,N_49533,N_49120);
nand UO_4417 (O_4417,N_49507,N_49727);
xor UO_4418 (O_4418,N_49869,N_48317);
nor UO_4419 (O_4419,N_49281,N_49225);
nand UO_4420 (O_4420,N_48461,N_48873);
nand UO_4421 (O_4421,N_48030,N_49531);
nand UO_4422 (O_4422,N_48308,N_49505);
nand UO_4423 (O_4423,N_49267,N_48906);
nand UO_4424 (O_4424,N_49822,N_49472);
xnor UO_4425 (O_4425,N_48384,N_49655);
nand UO_4426 (O_4426,N_48252,N_49801);
or UO_4427 (O_4427,N_49714,N_49126);
and UO_4428 (O_4428,N_48671,N_49074);
nand UO_4429 (O_4429,N_48453,N_49319);
xor UO_4430 (O_4430,N_49559,N_49987);
xnor UO_4431 (O_4431,N_48347,N_49917);
or UO_4432 (O_4432,N_48310,N_48270);
xnor UO_4433 (O_4433,N_48540,N_48877);
nor UO_4434 (O_4434,N_48269,N_48535);
or UO_4435 (O_4435,N_48083,N_49815);
or UO_4436 (O_4436,N_49880,N_49020);
and UO_4437 (O_4437,N_49547,N_49895);
or UO_4438 (O_4438,N_49260,N_48151);
or UO_4439 (O_4439,N_49564,N_48629);
nand UO_4440 (O_4440,N_49645,N_48368);
xnor UO_4441 (O_4441,N_48396,N_49089);
nor UO_4442 (O_4442,N_49124,N_48476);
xnor UO_4443 (O_4443,N_49222,N_48437);
or UO_4444 (O_4444,N_48159,N_49596);
nor UO_4445 (O_4445,N_49653,N_48420);
nand UO_4446 (O_4446,N_48103,N_48124);
xor UO_4447 (O_4447,N_49010,N_49196);
nor UO_4448 (O_4448,N_48164,N_48532);
or UO_4449 (O_4449,N_48110,N_49455);
nor UO_4450 (O_4450,N_49488,N_49859);
nand UO_4451 (O_4451,N_49906,N_48094);
nand UO_4452 (O_4452,N_48750,N_49545);
nand UO_4453 (O_4453,N_48120,N_48622);
xnor UO_4454 (O_4454,N_49507,N_48015);
nor UO_4455 (O_4455,N_48572,N_49996);
nand UO_4456 (O_4456,N_49088,N_49649);
nor UO_4457 (O_4457,N_49989,N_49065);
and UO_4458 (O_4458,N_48774,N_48012);
and UO_4459 (O_4459,N_49444,N_49140);
or UO_4460 (O_4460,N_48192,N_48513);
xor UO_4461 (O_4461,N_48665,N_49164);
nand UO_4462 (O_4462,N_48854,N_48797);
or UO_4463 (O_4463,N_48461,N_49353);
nor UO_4464 (O_4464,N_48465,N_49746);
or UO_4465 (O_4465,N_49496,N_49763);
nor UO_4466 (O_4466,N_48830,N_48309);
nor UO_4467 (O_4467,N_48343,N_48400);
xnor UO_4468 (O_4468,N_49090,N_49190);
nor UO_4469 (O_4469,N_48349,N_49539);
nand UO_4470 (O_4470,N_48697,N_48620);
nor UO_4471 (O_4471,N_48891,N_48448);
xor UO_4472 (O_4472,N_49185,N_49854);
xnor UO_4473 (O_4473,N_49653,N_49899);
nor UO_4474 (O_4474,N_48347,N_49427);
or UO_4475 (O_4475,N_48465,N_48017);
nand UO_4476 (O_4476,N_49958,N_48309);
xor UO_4477 (O_4477,N_48801,N_48129);
nor UO_4478 (O_4478,N_49790,N_49065);
nand UO_4479 (O_4479,N_48059,N_48610);
or UO_4480 (O_4480,N_49866,N_49766);
xnor UO_4481 (O_4481,N_48427,N_48180);
or UO_4482 (O_4482,N_48663,N_48397);
xnor UO_4483 (O_4483,N_48866,N_48746);
xnor UO_4484 (O_4484,N_48517,N_48614);
or UO_4485 (O_4485,N_48432,N_49518);
or UO_4486 (O_4486,N_48293,N_49626);
xor UO_4487 (O_4487,N_48811,N_49724);
or UO_4488 (O_4488,N_49196,N_49676);
and UO_4489 (O_4489,N_48196,N_48681);
and UO_4490 (O_4490,N_48406,N_48653);
and UO_4491 (O_4491,N_49389,N_49243);
xor UO_4492 (O_4492,N_48403,N_49580);
and UO_4493 (O_4493,N_48421,N_48853);
and UO_4494 (O_4494,N_48647,N_49844);
or UO_4495 (O_4495,N_48002,N_48450);
xor UO_4496 (O_4496,N_48837,N_49662);
nand UO_4497 (O_4497,N_49144,N_49609);
xnor UO_4498 (O_4498,N_49014,N_49870);
nand UO_4499 (O_4499,N_49740,N_48182);
and UO_4500 (O_4500,N_49264,N_48966);
xnor UO_4501 (O_4501,N_49861,N_48166);
and UO_4502 (O_4502,N_48645,N_49856);
xor UO_4503 (O_4503,N_48313,N_49822);
and UO_4504 (O_4504,N_49447,N_49840);
and UO_4505 (O_4505,N_49527,N_48305);
and UO_4506 (O_4506,N_49009,N_49390);
nand UO_4507 (O_4507,N_48711,N_48141);
or UO_4508 (O_4508,N_48996,N_48240);
and UO_4509 (O_4509,N_49112,N_49923);
and UO_4510 (O_4510,N_48509,N_48966);
nor UO_4511 (O_4511,N_48628,N_49328);
nand UO_4512 (O_4512,N_48305,N_48756);
nand UO_4513 (O_4513,N_48495,N_48351);
xor UO_4514 (O_4514,N_48797,N_48264);
nand UO_4515 (O_4515,N_48527,N_49535);
xor UO_4516 (O_4516,N_49234,N_49322);
nor UO_4517 (O_4517,N_49382,N_48631);
and UO_4518 (O_4518,N_49363,N_48954);
nand UO_4519 (O_4519,N_49857,N_48183);
and UO_4520 (O_4520,N_49307,N_49958);
xor UO_4521 (O_4521,N_49044,N_49049);
xor UO_4522 (O_4522,N_48586,N_48798);
and UO_4523 (O_4523,N_49714,N_49363);
xor UO_4524 (O_4524,N_48483,N_49963);
nand UO_4525 (O_4525,N_48103,N_48718);
nor UO_4526 (O_4526,N_48758,N_49776);
xnor UO_4527 (O_4527,N_48081,N_49390);
nor UO_4528 (O_4528,N_49715,N_49892);
nor UO_4529 (O_4529,N_49224,N_48398);
xnor UO_4530 (O_4530,N_49734,N_49618);
nor UO_4531 (O_4531,N_48564,N_48549);
and UO_4532 (O_4532,N_48293,N_48546);
nand UO_4533 (O_4533,N_49450,N_49688);
or UO_4534 (O_4534,N_48815,N_48611);
or UO_4535 (O_4535,N_48073,N_48557);
or UO_4536 (O_4536,N_49972,N_49663);
nand UO_4537 (O_4537,N_48180,N_48616);
nor UO_4538 (O_4538,N_49524,N_49903);
or UO_4539 (O_4539,N_49553,N_49175);
nand UO_4540 (O_4540,N_48649,N_49017);
or UO_4541 (O_4541,N_49060,N_49204);
nand UO_4542 (O_4542,N_48222,N_48792);
and UO_4543 (O_4543,N_48661,N_48293);
or UO_4544 (O_4544,N_49365,N_49594);
xor UO_4545 (O_4545,N_48126,N_48363);
nand UO_4546 (O_4546,N_49121,N_48909);
nor UO_4547 (O_4547,N_49428,N_48553);
and UO_4548 (O_4548,N_49393,N_49271);
and UO_4549 (O_4549,N_48332,N_48642);
or UO_4550 (O_4550,N_49857,N_48814);
or UO_4551 (O_4551,N_48177,N_48933);
xnor UO_4552 (O_4552,N_49464,N_48465);
and UO_4553 (O_4553,N_49275,N_49673);
and UO_4554 (O_4554,N_49229,N_49637);
xor UO_4555 (O_4555,N_48752,N_48293);
xor UO_4556 (O_4556,N_48194,N_49896);
nand UO_4557 (O_4557,N_48097,N_49997);
xor UO_4558 (O_4558,N_48785,N_49265);
xnor UO_4559 (O_4559,N_49573,N_49905);
xor UO_4560 (O_4560,N_48268,N_49737);
xnor UO_4561 (O_4561,N_48077,N_48400);
nand UO_4562 (O_4562,N_49990,N_48029);
xor UO_4563 (O_4563,N_48653,N_48129);
and UO_4564 (O_4564,N_49451,N_49237);
and UO_4565 (O_4565,N_48335,N_48954);
xnor UO_4566 (O_4566,N_49716,N_48965);
or UO_4567 (O_4567,N_48359,N_49505);
xnor UO_4568 (O_4568,N_48791,N_49934);
and UO_4569 (O_4569,N_49040,N_48019);
or UO_4570 (O_4570,N_49715,N_49236);
xnor UO_4571 (O_4571,N_48613,N_49836);
nor UO_4572 (O_4572,N_48042,N_49694);
xor UO_4573 (O_4573,N_48157,N_49953);
and UO_4574 (O_4574,N_49552,N_49029);
nor UO_4575 (O_4575,N_48477,N_49509);
nor UO_4576 (O_4576,N_48576,N_48186);
xnor UO_4577 (O_4577,N_48787,N_49747);
or UO_4578 (O_4578,N_49694,N_49738);
nor UO_4579 (O_4579,N_49085,N_48533);
nor UO_4580 (O_4580,N_49549,N_49080);
or UO_4581 (O_4581,N_48942,N_48867);
nor UO_4582 (O_4582,N_48619,N_48662);
and UO_4583 (O_4583,N_48738,N_49540);
nand UO_4584 (O_4584,N_49326,N_48596);
or UO_4585 (O_4585,N_48855,N_48934);
nor UO_4586 (O_4586,N_48962,N_48998);
and UO_4587 (O_4587,N_48378,N_48158);
nand UO_4588 (O_4588,N_48282,N_48696);
and UO_4589 (O_4589,N_49675,N_48961);
nand UO_4590 (O_4590,N_48659,N_49318);
or UO_4591 (O_4591,N_48235,N_48334);
xor UO_4592 (O_4592,N_48104,N_48466);
or UO_4593 (O_4593,N_49304,N_49513);
xnor UO_4594 (O_4594,N_48837,N_49096);
nand UO_4595 (O_4595,N_49308,N_49213);
nand UO_4596 (O_4596,N_49369,N_48357);
xnor UO_4597 (O_4597,N_48343,N_49858);
nor UO_4598 (O_4598,N_49269,N_49238);
nand UO_4599 (O_4599,N_48568,N_48086);
xnor UO_4600 (O_4600,N_48839,N_49401);
nor UO_4601 (O_4601,N_48865,N_48033);
nor UO_4602 (O_4602,N_49410,N_48242);
nor UO_4603 (O_4603,N_49493,N_48017);
xor UO_4604 (O_4604,N_48701,N_48371);
xnor UO_4605 (O_4605,N_49350,N_48328);
nor UO_4606 (O_4606,N_49391,N_48153);
and UO_4607 (O_4607,N_49400,N_48716);
or UO_4608 (O_4608,N_49350,N_49818);
nand UO_4609 (O_4609,N_49601,N_49702);
nor UO_4610 (O_4610,N_49282,N_48886);
nor UO_4611 (O_4611,N_49107,N_48397);
xnor UO_4612 (O_4612,N_48171,N_48380);
xnor UO_4613 (O_4613,N_49885,N_48327);
or UO_4614 (O_4614,N_48339,N_49025);
nand UO_4615 (O_4615,N_48034,N_48228);
and UO_4616 (O_4616,N_48432,N_48679);
nor UO_4617 (O_4617,N_48884,N_49839);
nand UO_4618 (O_4618,N_48250,N_48689);
nand UO_4619 (O_4619,N_48071,N_49494);
nand UO_4620 (O_4620,N_49277,N_48278);
or UO_4621 (O_4621,N_48366,N_49133);
and UO_4622 (O_4622,N_49876,N_48027);
nand UO_4623 (O_4623,N_48104,N_48723);
and UO_4624 (O_4624,N_48432,N_48845);
nor UO_4625 (O_4625,N_48981,N_48403);
or UO_4626 (O_4626,N_49283,N_48891);
nor UO_4627 (O_4627,N_49171,N_48187);
nand UO_4628 (O_4628,N_49194,N_49501);
xor UO_4629 (O_4629,N_48139,N_49370);
xnor UO_4630 (O_4630,N_48178,N_49359);
or UO_4631 (O_4631,N_48936,N_48709);
or UO_4632 (O_4632,N_49411,N_49175);
nand UO_4633 (O_4633,N_49250,N_48200);
or UO_4634 (O_4634,N_48949,N_48390);
nand UO_4635 (O_4635,N_48062,N_48697);
and UO_4636 (O_4636,N_49870,N_49015);
nor UO_4637 (O_4637,N_48781,N_48271);
or UO_4638 (O_4638,N_49960,N_48701);
nand UO_4639 (O_4639,N_48045,N_49667);
nor UO_4640 (O_4640,N_49562,N_49958);
and UO_4641 (O_4641,N_48898,N_49537);
or UO_4642 (O_4642,N_49922,N_49337);
nand UO_4643 (O_4643,N_49181,N_48463);
and UO_4644 (O_4644,N_49505,N_48957);
nor UO_4645 (O_4645,N_48314,N_48328);
nand UO_4646 (O_4646,N_48338,N_48053);
nor UO_4647 (O_4647,N_49508,N_48270);
and UO_4648 (O_4648,N_48769,N_48776);
or UO_4649 (O_4649,N_48922,N_48712);
and UO_4650 (O_4650,N_48438,N_48843);
nand UO_4651 (O_4651,N_49951,N_49427);
or UO_4652 (O_4652,N_48766,N_49269);
xor UO_4653 (O_4653,N_49531,N_49634);
or UO_4654 (O_4654,N_49682,N_48959);
nand UO_4655 (O_4655,N_49011,N_48327);
and UO_4656 (O_4656,N_49309,N_49799);
nand UO_4657 (O_4657,N_49953,N_49576);
or UO_4658 (O_4658,N_48771,N_49245);
or UO_4659 (O_4659,N_48160,N_49880);
nand UO_4660 (O_4660,N_48275,N_48794);
xnor UO_4661 (O_4661,N_48095,N_48230);
nand UO_4662 (O_4662,N_48595,N_48088);
nor UO_4663 (O_4663,N_49134,N_49816);
nor UO_4664 (O_4664,N_48293,N_49593);
nand UO_4665 (O_4665,N_48313,N_48580);
xor UO_4666 (O_4666,N_49393,N_48427);
xor UO_4667 (O_4667,N_48175,N_49749);
or UO_4668 (O_4668,N_49744,N_48374);
or UO_4669 (O_4669,N_48838,N_49790);
xnor UO_4670 (O_4670,N_49061,N_48789);
nor UO_4671 (O_4671,N_48759,N_48383);
nand UO_4672 (O_4672,N_49187,N_49414);
xnor UO_4673 (O_4673,N_48660,N_48156);
or UO_4674 (O_4674,N_49435,N_48522);
xnor UO_4675 (O_4675,N_49546,N_49030);
nor UO_4676 (O_4676,N_48494,N_48955);
or UO_4677 (O_4677,N_49778,N_49278);
xor UO_4678 (O_4678,N_49596,N_48622);
and UO_4679 (O_4679,N_48494,N_49946);
or UO_4680 (O_4680,N_48061,N_48346);
xnor UO_4681 (O_4681,N_48760,N_49558);
nand UO_4682 (O_4682,N_48656,N_49666);
nand UO_4683 (O_4683,N_49637,N_48806);
nand UO_4684 (O_4684,N_48585,N_48587);
nor UO_4685 (O_4685,N_49482,N_48832);
nand UO_4686 (O_4686,N_49000,N_48005);
xor UO_4687 (O_4687,N_49129,N_49136);
nand UO_4688 (O_4688,N_49079,N_49909);
nand UO_4689 (O_4689,N_48653,N_48592);
nand UO_4690 (O_4690,N_48162,N_48278);
nor UO_4691 (O_4691,N_49215,N_48715);
nand UO_4692 (O_4692,N_49459,N_49902);
or UO_4693 (O_4693,N_48422,N_49758);
or UO_4694 (O_4694,N_49789,N_48982);
nor UO_4695 (O_4695,N_48225,N_49416);
and UO_4696 (O_4696,N_49211,N_48606);
xnor UO_4697 (O_4697,N_48872,N_49877);
xnor UO_4698 (O_4698,N_49204,N_49170);
and UO_4699 (O_4699,N_48020,N_48855);
nand UO_4700 (O_4700,N_48300,N_49260);
xnor UO_4701 (O_4701,N_49642,N_49075);
and UO_4702 (O_4702,N_49973,N_49912);
xnor UO_4703 (O_4703,N_49599,N_49689);
xnor UO_4704 (O_4704,N_48097,N_49303);
nand UO_4705 (O_4705,N_48414,N_49325);
nand UO_4706 (O_4706,N_49827,N_48466);
or UO_4707 (O_4707,N_49496,N_48076);
nand UO_4708 (O_4708,N_49010,N_49978);
nand UO_4709 (O_4709,N_48037,N_48117);
nand UO_4710 (O_4710,N_48081,N_48870);
xor UO_4711 (O_4711,N_49910,N_48490);
and UO_4712 (O_4712,N_48099,N_49257);
nor UO_4713 (O_4713,N_49944,N_48453);
xor UO_4714 (O_4714,N_49316,N_48873);
nand UO_4715 (O_4715,N_48661,N_48714);
and UO_4716 (O_4716,N_48951,N_49745);
xor UO_4717 (O_4717,N_49840,N_49759);
xnor UO_4718 (O_4718,N_48668,N_48436);
xnor UO_4719 (O_4719,N_49604,N_49564);
xnor UO_4720 (O_4720,N_48147,N_49169);
and UO_4721 (O_4721,N_48898,N_48651);
xnor UO_4722 (O_4722,N_48886,N_49488);
and UO_4723 (O_4723,N_48517,N_48860);
nor UO_4724 (O_4724,N_49466,N_49189);
nand UO_4725 (O_4725,N_49128,N_48413);
nor UO_4726 (O_4726,N_48684,N_49387);
and UO_4727 (O_4727,N_49820,N_49276);
and UO_4728 (O_4728,N_48167,N_48315);
nor UO_4729 (O_4729,N_49161,N_49758);
nor UO_4730 (O_4730,N_49124,N_48068);
and UO_4731 (O_4731,N_48835,N_49843);
and UO_4732 (O_4732,N_49285,N_48307);
xor UO_4733 (O_4733,N_48455,N_48315);
and UO_4734 (O_4734,N_48361,N_48686);
nand UO_4735 (O_4735,N_49955,N_48000);
nor UO_4736 (O_4736,N_48717,N_48912);
and UO_4737 (O_4737,N_49837,N_49603);
xnor UO_4738 (O_4738,N_49554,N_49220);
xnor UO_4739 (O_4739,N_48320,N_49573);
nand UO_4740 (O_4740,N_49919,N_49407);
nand UO_4741 (O_4741,N_49383,N_49718);
xor UO_4742 (O_4742,N_48817,N_49605);
xnor UO_4743 (O_4743,N_49582,N_49472);
nor UO_4744 (O_4744,N_48756,N_49083);
or UO_4745 (O_4745,N_48779,N_49008);
or UO_4746 (O_4746,N_48148,N_49824);
nor UO_4747 (O_4747,N_48330,N_49266);
xor UO_4748 (O_4748,N_48493,N_48534);
nand UO_4749 (O_4749,N_49203,N_48584);
and UO_4750 (O_4750,N_48753,N_49946);
and UO_4751 (O_4751,N_49379,N_49180);
xnor UO_4752 (O_4752,N_49052,N_49194);
xor UO_4753 (O_4753,N_48173,N_49297);
xor UO_4754 (O_4754,N_48701,N_48772);
nor UO_4755 (O_4755,N_49471,N_48594);
xnor UO_4756 (O_4756,N_48439,N_49464);
nand UO_4757 (O_4757,N_49540,N_49435);
and UO_4758 (O_4758,N_49810,N_49314);
nand UO_4759 (O_4759,N_48008,N_48558);
nor UO_4760 (O_4760,N_49388,N_48287);
nand UO_4761 (O_4761,N_49990,N_49389);
and UO_4762 (O_4762,N_48735,N_49377);
xnor UO_4763 (O_4763,N_48151,N_49677);
nand UO_4764 (O_4764,N_48550,N_48390);
and UO_4765 (O_4765,N_48636,N_48863);
nand UO_4766 (O_4766,N_48275,N_49550);
and UO_4767 (O_4767,N_48338,N_49500);
or UO_4768 (O_4768,N_49264,N_48276);
xor UO_4769 (O_4769,N_48761,N_49663);
xnor UO_4770 (O_4770,N_48202,N_49354);
or UO_4771 (O_4771,N_49637,N_48710);
and UO_4772 (O_4772,N_48081,N_48622);
or UO_4773 (O_4773,N_49498,N_48237);
xor UO_4774 (O_4774,N_49460,N_49529);
and UO_4775 (O_4775,N_49746,N_48216);
nor UO_4776 (O_4776,N_49396,N_48970);
nand UO_4777 (O_4777,N_49396,N_49955);
nand UO_4778 (O_4778,N_48904,N_49266);
and UO_4779 (O_4779,N_49553,N_48807);
and UO_4780 (O_4780,N_49493,N_49715);
xor UO_4781 (O_4781,N_49381,N_49638);
xor UO_4782 (O_4782,N_49519,N_48885);
xnor UO_4783 (O_4783,N_48732,N_48772);
or UO_4784 (O_4784,N_48635,N_48661);
nand UO_4785 (O_4785,N_48022,N_49442);
and UO_4786 (O_4786,N_49153,N_49479);
xnor UO_4787 (O_4787,N_49246,N_49319);
and UO_4788 (O_4788,N_48467,N_48456);
nor UO_4789 (O_4789,N_48083,N_49802);
or UO_4790 (O_4790,N_49861,N_49993);
or UO_4791 (O_4791,N_49326,N_49502);
or UO_4792 (O_4792,N_49244,N_49027);
and UO_4793 (O_4793,N_49527,N_48007);
and UO_4794 (O_4794,N_49014,N_48883);
nor UO_4795 (O_4795,N_48426,N_49963);
nand UO_4796 (O_4796,N_48367,N_48005);
nor UO_4797 (O_4797,N_49404,N_48820);
nor UO_4798 (O_4798,N_49339,N_48643);
nor UO_4799 (O_4799,N_48588,N_49969);
nand UO_4800 (O_4800,N_49510,N_48175);
nor UO_4801 (O_4801,N_48384,N_48708);
nand UO_4802 (O_4802,N_48836,N_49316);
nor UO_4803 (O_4803,N_48555,N_48046);
xor UO_4804 (O_4804,N_49510,N_48115);
or UO_4805 (O_4805,N_48699,N_49983);
nor UO_4806 (O_4806,N_48925,N_49522);
nor UO_4807 (O_4807,N_48745,N_49465);
and UO_4808 (O_4808,N_48814,N_49507);
nor UO_4809 (O_4809,N_49756,N_49095);
or UO_4810 (O_4810,N_49459,N_49043);
nand UO_4811 (O_4811,N_48438,N_48141);
nor UO_4812 (O_4812,N_48766,N_48560);
nor UO_4813 (O_4813,N_48035,N_49693);
nand UO_4814 (O_4814,N_49124,N_49288);
xnor UO_4815 (O_4815,N_49282,N_49965);
xor UO_4816 (O_4816,N_48821,N_49017);
or UO_4817 (O_4817,N_49563,N_49375);
xor UO_4818 (O_4818,N_49578,N_48171);
nand UO_4819 (O_4819,N_48170,N_48381);
or UO_4820 (O_4820,N_49417,N_49669);
and UO_4821 (O_4821,N_48039,N_49088);
nand UO_4822 (O_4822,N_48611,N_49550);
or UO_4823 (O_4823,N_49862,N_48397);
or UO_4824 (O_4824,N_49716,N_48377);
xor UO_4825 (O_4825,N_49949,N_48421);
and UO_4826 (O_4826,N_48451,N_48706);
nor UO_4827 (O_4827,N_49712,N_48349);
xnor UO_4828 (O_4828,N_49289,N_48341);
nand UO_4829 (O_4829,N_48378,N_48154);
and UO_4830 (O_4830,N_49860,N_49783);
xor UO_4831 (O_4831,N_49263,N_48453);
or UO_4832 (O_4832,N_48066,N_49135);
and UO_4833 (O_4833,N_48836,N_48645);
nor UO_4834 (O_4834,N_48857,N_48885);
and UO_4835 (O_4835,N_49241,N_49714);
and UO_4836 (O_4836,N_49598,N_49363);
xor UO_4837 (O_4837,N_48850,N_49690);
xnor UO_4838 (O_4838,N_48985,N_48285);
xor UO_4839 (O_4839,N_48184,N_49623);
nand UO_4840 (O_4840,N_48658,N_48474);
and UO_4841 (O_4841,N_49235,N_48598);
nor UO_4842 (O_4842,N_49582,N_49854);
and UO_4843 (O_4843,N_48684,N_49407);
nand UO_4844 (O_4844,N_49579,N_48934);
and UO_4845 (O_4845,N_48936,N_48367);
and UO_4846 (O_4846,N_48561,N_49581);
nor UO_4847 (O_4847,N_48612,N_49501);
and UO_4848 (O_4848,N_48155,N_49566);
and UO_4849 (O_4849,N_49397,N_49558);
or UO_4850 (O_4850,N_49486,N_49999);
nand UO_4851 (O_4851,N_48797,N_49267);
and UO_4852 (O_4852,N_48982,N_49854);
nor UO_4853 (O_4853,N_48891,N_49385);
xor UO_4854 (O_4854,N_49625,N_49496);
xnor UO_4855 (O_4855,N_48631,N_49371);
nor UO_4856 (O_4856,N_49702,N_49241);
or UO_4857 (O_4857,N_49030,N_48627);
and UO_4858 (O_4858,N_49691,N_49652);
or UO_4859 (O_4859,N_49165,N_48538);
xor UO_4860 (O_4860,N_49905,N_48137);
nand UO_4861 (O_4861,N_48767,N_49865);
nand UO_4862 (O_4862,N_49115,N_49639);
nand UO_4863 (O_4863,N_48847,N_49813);
and UO_4864 (O_4864,N_48235,N_49875);
and UO_4865 (O_4865,N_48698,N_48143);
and UO_4866 (O_4866,N_49765,N_48822);
xor UO_4867 (O_4867,N_49005,N_48071);
nor UO_4868 (O_4868,N_48889,N_48586);
nor UO_4869 (O_4869,N_49276,N_48540);
or UO_4870 (O_4870,N_49326,N_48499);
xor UO_4871 (O_4871,N_48772,N_49261);
and UO_4872 (O_4872,N_49338,N_49053);
xor UO_4873 (O_4873,N_49701,N_48824);
nor UO_4874 (O_4874,N_48209,N_49252);
or UO_4875 (O_4875,N_49710,N_49363);
nor UO_4876 (O_4876,N_48045,N_48605);
xor UO_4877 (O_4877,N_48412,N_48209);
nor UO_4878 (O_4878,N_49591,N_49899);
or UO_4879 (O_4879,N_49499,N_49921);
xor UO_4880 (O_4880,N_49976,N_49927);
xnor UO_4881 (O_4881,N_49381,N_49344);
nand UO_4882 (O_4882,N_49289,N_48833);
and UO_4883 (O_4883,N_49093,N_49108);
and UO_4884 (O_4884,N_49537,N_48109);
or UO_4885 (O_4885,N_49475,N_49147);
nand UO_4886 (O_4886,N_49244,N_49127);
nor UO_4887 (O_4887,N_48373,N_48358);
xnor UO_4888 (O_4888,N_49983,N_48966);
nor UO_4889 (O_4889,N_49199,N_48844);
or UO_4890 (O_4890,N_48843,N_48207);
xnor UO_4891 (O_4891,N_48102,N_48749);
or UO_4892 (O_4892,N_48441,N_49685);
nand UO_4893 (O_4893,N_48367,N_49194);
xnor UO_4894 (O_4894,N_48312,N_49567);
nor UO_4895 (O_4895,N_49404,N_48753);
nor UO_4896 (O_4896,N_48663,N_49726);
nand UO_4897 (O_4897,N_49903,N_49829);
nand UO_4898 (O_4898,N_49913,N_49696);
xor UO_4899 (O_4899,N_48175,N_49505);
and UO_4900 (O_4900,N_49497,N_48616);
xnor UO_4901 (O_4901,N_48617,N_49753);
nand UO_4902 (O_4902,N_49980,N_48730);
xnor UO_4903 (O_4903,N_48737,N_48321);
nor UO_4904 (O_4904,N_48451,N_49914);
nand UO_4905 (O_4905,N_49397,N_48608);
or UO_4906 (O_4906,N_48272,N_48183);
nand UO_4907 (O_4907,N_49935,N_48220);
nor UO_4908 (O_4908,N_49631,N_49597);
and UO_4909 (O_4909,N_49313,N_49469);
and UO_4910 (O_4910,N_49949,N_49247);
or UO_4911 (O_4911,N_48747,N_48452);
and UO_4912 (O_4912,N_48081,N_48348);
and UO_4913 (O_4913,N_48043,N_49506);
xor UO_4914 (O_4914,N_49171,N_49799);
or UO_4915 (O_4915,N_49700,N_48273);
or UO_4916 (O_4916,N_49877,N_49719);
xnor UO_4917 (O_4917,N_48818,N_48794);
nand UO_4918 (O_4918,N_49991,N_49262);
nor UO_4919 (O_4919,N_49438,N_49304);
and UO_4920 (O_4920,N_49956,N_48564);
nand UO_4921 (O_4921,N_48264,N_49557);
xor UO_4922 (O_4922,N_49070,N_49550);
and UO_4923 (O_4923,N_49960,N_49232);
nand UO_4924 (O_4924,N_48933,N_48019);
xor UO_4925 (O_4925,N_49618,N_48259);
nor UO_4926 (O_4926,N_49112,N_49788);
or UO_4927 (O_4927,N_49019,N_49336);
nor UO_4928 (O_4928,N_49906,N_48442);
or UO_4929 (O_4929,N_48683,N_48719);
nor UO_4930 (O_4930,N_49610,N_48142);
or UO_4931 (O_4931,N_48059,N_49284);
xnor UO_4932 (O_4932,N_49678,N_49343);
or UO_4933 (O_4933,N_48538,N_49796);
and UO_4934 (O_4934,N_49390,N_49094);
or UO_4935 (O_4935,N_48895,N_49630);
nand UO_4936 (O_4936,N_48769,N_48016);
xnor UO_4937 (O_4937,N_48206,N_49967);
nor UO_4938 (O_4938,N_49032,N_48310);
nor UO_4939 (O_4939,N_48508,N_49454);
or UO_4940 (O_4940,N_48402,N_48896);
nor UO_4941 (O_4941,N_48913,N_48562);
and UO_4942 (O_4942,N_49856,N_49812);
or UO_4943 (O_4943,N_48760,N_49367);
or UO_4944 (O_4944,N_49940,N_49696);
xor UO_4945 (O_4945,N_49387,N_48447);
nand UO_4946 (O_4946,N_48171,N_49484);
and UO_4947 (O_4947,N_49457,N_49400);
and UO_4948 (O_4948,N_49859,N_48503);
and UO_4949 (O_4949,N_49248,N_49463);
xor UO_4950 (O_4950,N_49876,N_48516);
or UO_4951 (O_4951,N_48825,N_49045);
xnor UO_4952 (O_4952,N_48973,N_49652);
xor UO_4953 (O_4953,N_48025,N_49090);
or UO_4954 (O_4954,N_48762,N_48875);
xor UO_4955 (O_4955,N_48984,N_49589);
nand UO_4956 (O_4956,N_48577,N_48415);
xnor UO_4957 (O_4957,N_48940,N_49255);
or UO_4958 (O_4958,N_49328,N_48098);
xnor UO_4959 (O_4959,N_49949,N_49665);
and UO_4960 (O_4960,N_48679,N_49841);
nand UO_4961 (O_4961,N_49492,N_49683);
nand UO_4962 (O_4962,N_48948,N_49993);
and UO_4963 (O_4963,N_49206,N_48899);
or UO_4964 (O_4964,N_48641,N_49649);
xor UO_4965 (O_4965,N_48366,N_48216);
or UO_4966 (O_4966,N_49659,N_49918);
or UO_4967 (O_4967,N_48350,N_48886);
nor UO_4968 (O_4968,N_49256,N_49738);
nand UO_4969 (O_4969,N_48073,N_48077);
xor UO_4970 (O_4970,N_48818,N_49038);
xnor UO_4971 (O_4971,N_49926,N_49657);
or UO_4972 (O_4972,N_48426,N_49010);
and UO_4973 (O_4973,N_48000,N_49309);
nand UO_4974 (O_4974,N_49838,N_49992);
and UO_4975 (O_4975,N_49836,N_49591);
nor UO_4976 (O_4976,N_48878,N_49734);
nor UO_4977 (O_4977,N_49267,N_48717);
nor UO_4978 (O_4978,N_49508,N_49351);
nand UO_4979 (O_4979,N_48832,N_49349);
or UO_4980 (O_4980,N_48870,N_48208);
and UO_4981 (O_4981,N_48801,N_48367);
nand UO_4982 (O_4982,N_49113,N_48602);
xnor UO_4983 (O_4983,N_48206,N_49897);
xor UO_4984 (O_4984,N_49895,N_48362);
or UO_4985 (O_4985,N_49295,N_49427);
nand UO_4986 (O_4986,N_48524,N_49915);
nand UO_4987 (O_4987,N_49826,N_48798);
or UO_4988 (O_4988,N_48666,N_48612);
nor UO_4989 (O_4989,N_48956,N_48999);
nor UO_4990 (O_4990,N_48924,N_48072);
nand UO_4991 (O_4991,N_48561,N_48744);
nor UO_4992 (O_4992,N_49067,N_48534);
xnor UO_4993 (O_4993,N_48293,N_49970);
nor UO_4994 (O_4994,N_48647,N_48891);
nor UO_4995 (O_4995,N_48697,N_48189);
nand UO_4996 (O_4996,N_48351,N_48547);
or UO_4997 (O_4997,N_49565,N_48645);
or UO_4998 (O_4998,N_48819,N_48189);
or UO_4999 (O_4999,N_49149,N_49480);
endmodule