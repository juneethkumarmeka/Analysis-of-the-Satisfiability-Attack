module basic_3000_30000_3500_100_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2626,In_1315);
xnor U1 (N_1,In_1220,In_30);
nand U2 (N_2,In_2174,In_1474);
nor U3 (N_3,In_606,In_462);
or U4 (N_4,In_2314,In_552);
or U5 (N_5,In_1496,In_169);
and U6 (N_6,In_1292,In_446);
or U7 (N_7,In_961,In_2076);
and U8 (N_8,In_198,In_866);
and U9 (N_9,In_2553,In_484);
nand U10 (N_10,In_2638,In_2729);
xnor U11 (N_11,In_1020,In_2029);
nor U12 (N_12,In_1097,In_2505);
and U13 (N_13,In_831,In_2120);
and U14 (N_14,In_527,In_1074);
nand U15 (N_15,In_878,In_1549);
nor U16 (N_16,In_792,In_1890);
and U17 (N_17,In_740,In_620);
or U18 (N_18,In_2479,In_787);
and U19 (N_19,In_767,In_2504);
and U20 (N_20,In_2933,In_144);
or U21 (N_21,In_1221,In_1499);
nand U22 (N_22,In_337,In_1889);
nand U23 (N_23,In_2861,In_2579);
and U24 (N_24,In_773,In_38);
xnor U25 (N_25,In_2750,In_966);
nor U26 (N_26,In_1516,In_2113);
and U27 (N_27,In_1631,In_1079);
nor U28 (N_28,In_1766,In_1666);
nor U29 (N_29,In_2222,In_2136);
xor U30 (N_30,In_1385,In_1783);
nand U31 (N_31,In_475,In_1787);
and U32 (N_32,In_1651,In_960);
or U33 (N_33,In_1392,In_2610);
and U34 (N_34,In_2059,In_2129);
and U35 (N_35,In_2480,In_2071);
nor U36 (N_36,In_2958,In_2023);
xnor U37 (N_37,In_2318,In_724);
nor U38 (N_38,In_2332,In_575);
or U39 (N_39,In_503,In_2909);
nand U40 (N_40,In_11,In_2527);
nand U41 (N_41,In_1540,In_2162);
or U42 (N_42,In_447,In_2916);
and U43 (N_43,In_2712,In_2485);
nand U44 (N_44,In_2284,In_1551);
and U45 (N_45,In_2664,In_2628);
nor U46 (N_46,In_2675,In_1722);
and U47 (N_47,In_612,In_406);
and U48 (N_48,In_304,In_2082);
or U49 (N_49,In_1948,In_886);
and U50 (N_50,In_303,In_1242);
xor U51 (N_51,In_892,In_2459);
nor U52 (N_52,In_1015,In_2022);
nor U53 (N_53,In_1086,In_1535);
nor U54 (N_54,In_2808,In_922);
and U55 (N_55,In_784,In_1665);
nor U56 (N_56,In_121,In_1262);
or U57 (N_57,In_2942,In_1753);
xor U58 (N_58,In_1974,In_432);
or U59 (N_59,In_2697,In_1260);
nor U60 (N_60,In_841,In_2234);
or U61 (N_61,In_1085,In_2379);
nor U62 (N_62,In_2900,In_893);
and U63 (N_63,In_2233,In_322);
xor U64 (N_64,In_1969,In_542);
xnor U65 (N_65,In_1923,In_1866);
nor U66 (N_66,In_1492,In_1489);
and U67 (N_67,In_1917,In_1700);
nand U68 (N_68,In_1579,In_2213);
and U69 (N_69,In_1448,In_2403);
nand U70 (N_70,In_1180,In_1121);
xor U71 (N_71,In_701,In_2524);
nor U72 (N_72,In_1172,In_857);
nand U73 (N_73,In_890,In_2765);
and U74 (N_74,In_572,In_327);
or U75 (N_75,In_2689,In_847);
nor U76 (N_76,In_2782,In_270);
nor U77 (N_77,In_654,In_1790);
or U78 (N_78,In_1911,In_342);
nor U79 (N_79,In_36,In_1184);
nor U80 (N_80,In_362,In_430);
nor U81 (N_81,In_2606,In_418);
and U82 (N_82,In_419,In_1028);
xnor U83 (N_83,In_1275,In_1487);
xor U84 (N_84,In_1583,In_1880);
or U85 (N_85,In_228,In_158);
and U86 (N_86,In_2425,In_1855);
nor U87 (N_87,In_648,In_1950);
xnor U88 (N_88,In_423,In_994);
and U89 (N_89,In_2793,In_436);
and U90 (N_90,In_1146,In_2354);
nand U91 (N_91,In_2047,In_167);
xor U92 (N_92,In_108,In_1286);
and U93 (N_93,In_443,In_1681);
nand U94 (N_94,In_309,In_1649);
and U95 (N_95,In_1368,In_1189);
nand U96 (N_96,In_904,In_725);
xnor U97 (N_97,In_2173,In_2776);
nor U98 (N_98,In_1192,In_1104);
or U99 (N_99,In_481,In_830);
nand U100 (N_100,In_1826,In_1591);
and U101 (N_101,In_1282,In_2096);
and U102 (N_102,In_2005,In_1329);
nor U103 (N_103,In_1747,In_1570);
nor U104 (N_104,In_1853,In_496);
and U105 (N_105,In_452,In_2061);
nor U106 (N_106,In_989,In_429);
and U107 (N_107,In_433,In_1862);
nor U108 (N_108,In_279,In_398);
and U109 (N_109,In_1979,In_2310);
or U110 (N_110,In_1542,In_1793);
nor U111 (N_111,In_2367,In_2705);
or U112 (N_112,In_906,In_2164);
or U113 (N_113,In_2516,In_2418);
nor U114 (N_114,In_427,In_827);
or U115 (N_115,In_1264,In_2848);
nor U116 (N_116,In_1530,In_2271);
or U117 (N_117,In_313,In_2017);
nand U118 (N_118,In_995,In_2454);
and U119 (N_119,In_2435,In_1557);
or U120 (N_120,In_1791,In_464);
nand U121 (N_121,In_1566,In_134);
nand U122 (N_122,In_2856,In_1961);
xnor U123 (N_123,In_289,In_1908);
nand U124 (N_124,In_128,In_1378);
or U125 (N_125,In_2919,In_405);
xnor U126 (N_126,In_1204,In_2789);
nand U127 (N_127,In_1161,In_1049);
nand U128 (N_128,In_2122,In_2883);
nand U129 (N_129,In_2088,In_2167);
and U130 (N_130,In_78,In_1254);
or U131 (N_131,In_448,In_1091);
nor U132 (N_132,In_71,In_1439);
and U133 (N_133,In_569,In_1431);
and U134 (N_134,In_455,In_412);
or U135 (N_135,In_2615,In_2405);
xor U136 (N_136,In_2652,In_488);
nor U137 (N_137,In_1182,In_2401);
and U138 (N_138,In_772,In_1323);
nor U139 (N_139,In_2008,In_958);
or U140 (N_140,In_400,In_2482);
and U141 (N_141,In_663,In_1854);
or U142 (N_142,In_1026,In_145);
nor U143 (N_143,In_1462,In_1812);
xnor U144 (N_144,In_340,In_1076);
or U145 (N_145,In_2000,In_2428);
or U146 (N_146,In_2016,In_2571);
nor U147 (N_147,In_1706,In_2097);
or U148 (N_148,In_2278,In_288);
and U149 (N_149,In_2833,In_2903);
nand U150 (N_150,In_335,In_68);
xor U151 (N_151,In_684,In_1864);
or U152 (N_152,In_576,In_2394);
and U153 (N_153,In_1522,In_2834);
and U154 (N_154,In_823,In_245);
nand U155 (N_155,In_1336,In_1699);
nor U156 (N_156,In_1475,In_1018);
nand U157 (N_157,In_929,In_903);
nor U158 (N_158,In_1650,In_1498);
nand U159 (N_159,In_162,In_2198);
and U160 (N_160,In_720,In_1830);
nor U161 (N_161,In_2941,In_1445);
xor U162 (N_162,In_1620,In_2749);
nand U163 (N_163,In_2984,In_763);
nor U164 (N_164,In_1767,In_2436);
or U165 (N_165,In_1678,In_2257);
and U166 (N_166,In_113,In_2921);
nor U167 (N_167,In_1344,In_1563);
nor U168 (N_168,In_1125,In_1723);
nand U169 (N_169,In_2528,In_1003);
or U170 (N_170,In_550,In_662);
xor U171 (N_171,In_1879,In_1034);
and U172 (N_172,In_1605,In_1256);
and U173 (N_173,In_482,In_1546);
nand U174 (N_174,In_2533,In_1603);
nand U175 (N_175,In_345,In_17);
nor U176 (N_176,In_2503,In_1395);
xor U177 (N_177,In_921,In_2562);
nand U178 (N_178,In_2719,In_840);
nand U179 (N_179,In_579,In_2975);
nand U180 (N_180,In_2678,In_949);
nor U181 (N_181,In_696,In_101);
xnor U182 (N_182,In_1046,In_616);
xnor U183 (N_183,In_1607,In_1343);
xnor U184 (N_184,In_1179,In_1616);
or U185 (N_185,In_2741,In_1960);
nand U186 (N_186,In_2980,In_1435);
nand U187 (N_187,In_514,In_421);
and U188 (N_188,In_199,In_79);
nor U189 (N_189,In_1981,In_1803);
nand U190 (N_190,In_1840,In_2429);
or U191 (N_191,In_2590,In_2823);
or U192 (N_192,In_2352,In_2398);
nand U193 (N_193,In_1721,In_1545);
and U194 (N_194,In_2778,In_2118);
or U195 (N_195,In_1623,In_96);
and U196 (N_196,In_672,In_1946);
nand U197 (N_197,In_2918,In_2602);
nand U198 (N_198,In_1446,In_2733);
nor U199 (N_199,In_1967,In_2825);
xnor U200 (N_200,In_1560,In_1165);
or U201 (N_201,In_1571,In_856);
xor U202 (N_202,In_1815,In_2668);
nand U203 (N_203,In_94,In_1027);
or U204 (N_204,In_875,In_1138);
nor U205 (N_205,In_846,In_1088);
and U206 (N_206,In_1502,In_204);
xnor U207 (N_207,In_1597,In_28);
and U208 (N_208,In_2341,In_2117);
nand U209 (N_209,In_2221,In_1784);
or U210 (N_210,In_839,In_1274);
nor U211 (N_211,In_1763,In_1328);
nand U212 (N_212,In_250,In_750);
or U213 (N_213,In_2507,In_1453);
xnor U214 (N_214,In_2681,In_986);
nor U215 (N_215,In_155,In_213);
nand U216 (N_216,In_1166,In_2779);
nor U217 (N_217,In_858,In_721);
xnor U218 (N_218,In_1910,In_2715);
xnor U219 (N_219,In_2100,In_2598);
xor U220 (N_220,In_2753,In_1170);
or U221 (N_221,In_853,In_291);
xnor U222 (N_222,In_2756,In_714);
and U223 (N_223,In_844,In_2423);
xnor U224 (N_224,In_388,In_2754);
or U225 (N_225,In_2214,In_2334);
and U226 (N_226,In_883,In_2366);
nand U227 (N_227,In_2333,In_221);
and U228 (N_228,In_717,In_2589);
nand U229 (N_229,In_190,In_642);
xnor U230 (N_230,In_2265,In_1541);
or U231 (N_231,In_2069,In_1949);
xor U232 (N_232,In_2619,In_2688);
xor U233 (N_233,In_1847,In_865);
and U234 (N_234,In_2669,In_2327);
or U235 (N_235,In_618,In_2349);
nand U236 (N_236,In_2850,In_2094);
and U237 (N_237,In_1482,In_2440);
or U238 (N_238,In_2841,In_2704);
nand U239 (N_239,In_330,In_2250);
and U240 (N_240,In_1430,In_2653);
or U241 (N_241,In_44,In_66);
xnor U242 (N_242,In_2330,In_1568);
nand U243 (N_243,In_1355,In_1929);
nand U244 (N_244,In_1313,In_2303);
or U245 (N_245,In_2104,In_2926);
nor U246 (N_246,In_2677,In_2790);
nor U247 (N_247,In_1209,In_235);
nand U248 (N_248,In_2720,In_163);
and U249 (N_249,In_31,In_237);
or U250 (N_250,In_2402,In_1225);
and U251 (N_251,In_461,In_1555);
or U252 (N_252,In_457,In_869);
xnor U253 (N_253,In_1127,In_2362);
nor U254 (N_254,In_105,In_1627);
nand U255 (N_255,In_563,In_231);
and U256 (N_256,In_2489,In_2228);
xor U257 (N_257,In_442,In_1525);
nor U258 (N_258,In_1765,In_2506);
xor U259 (N_259,In_440,In_1009);
xor U260 (N_260,In_272,In_668);
and U261 (N_261,In_2892,In_349);
xor U262 (N_262,In_782,In_2891);
or U263 (N_263,In_88,In_617);
or U264 (N_264,In_394,In_296);
and U265 (N_265,In_1108,In_1459);
nor U266 (N_266,In_2899,In_165);
and U267 (N_267,In_1068,In_2966);
nand U268 (N_268,In_943,In_69);
nand U269 (N_269,In_2988,In_803);
and U270 (N_270,In_545,In_2078);
or U271 (N_271,In_1695,In_339);
or U272 (N_272,In_1116,In_2177);
nand U273 (N_273,In_1234,In_381);
or U274 (N_274,In_1423,In_1188);
nand U275 (N_275,In_581,In_2180);
and U276 (N_276,In_2018,In_1450);
and U277 (N_277,In_657,In_506);
nand U278 (N_278,In_1661,In_1987);
xor U279 (N_279,In_1219,In_1001);
nor U280 (N_280,In_1303,In_346);
and U281 (N_281,In_1374,In_2817);
nand U282 (N_282,In_1604,In_1884);
and U283 (N_283,In_182,In_894);
or U284 (N_284,In_248,In_2744);
and U285 (N_285,In_534,In_2742);
or U286 (N_286,In_981,In_107);
xnor U287 (N_287,In_1071,In_202);
and U288 (N_288,In_794,In_2747);
or U289 (N_289,In_1141,In_1080);
or U290 (N_290,In_262,In_2380);
or U291 (N_291,In_467,In_806);
nor U292 (N_292,In_1696,In_2969);
and U293 (N_293,In_89,In_2316);
xnor U294 (N_294,In_927,In_1726);
nor U295 (N_295,In_781,In_1955);
nor U296 (N_296,In_1117,In_996);
nor U297 (N_297,In_2868,In_2137);
nand U298 (N_298,In_1066,In_1490);
nand U299 (N_299,In_1384,In_320);
nor U300 (N_300,In_765,In_1684);
nand U301 (N_301,In_2329,In_2205);
xnor U302 (N_302,In_1133,In_897);
nor U303 (N_303,In_2761,N_170);
xnor U304 (N_304,In_512,In_2940);
xnor U305 (N_305,N_220,In_2927);
or U306 (N_306,In_1156,In_473);
nand U307 (N_307,In_373,In_969);
nand U308 (N_308,In_1741,In_1750);
and U309 (N_309,In_716,In_679);
nor U310 (N_310,In_1801,In_1364);
or U311 (N_311,N_245,In_2549);
or U312 (N_312,In_32,In_1594);
nand U313 (N_313,N_253,N_24);
nand U314 (N_314,N_229,In_2857);
or U315 (N_315,In_465,In_2434);
nor U316 (N_316,In_1107,In_605);
nor U317 (N_317,In_2703,In_2027);
nor U318 (N_318,In_1007,N_231);
or U319 (N_319,In_546,In_2378);
xor U320 (N_320,In_1333,In_597);
and U321 (N_321,In_450,In_1858);
nand U322 (N_322,N_219,In_1366);
and U323 (N_323,N_159,In_1207);
nand U324 (N_324,In_2740,In_985);
xnor U325 (N_325,In_741,In_812);
nor U326 (N_326,In_12,In_1304);
and U327 (N_327,In_2110,In_212);
xnor U328 (N_328,In_305,In_417);
nor U329 (N_329,In_2643,In_2152);
xnor U330 (N_330,In_2490,In_21);
nand U331 (N_331,In_2475,N_279);
nor U332 (N_332,In_6,In_1472);
and U333 (N_333,In_562,In_116);
nand U334 (N_334,In_1521,In_602);
nand U335 (N_335,In_2014,In_2873);
or U336 (N_336,In_2932,In_907);
or U337 (N_337,In_81,In_1985);
and U338 (N_338,N_278,In_1720);
xnor U339 (N_339,In_141,In_2344);
xor U340 (N_340,N_50,N_124);
xor U341 (N_341,N_5,N_185);
nor U342 (N_342,In_468,In_926);
and U343 (N_343,In_2124,In_2599);
nor U344 (N_344,In_249,In_2649);
nor U345 (N_345,In_2295,In_637);
and U346 (N_346,In_1638,In_2994);
or U347 (N_347,In_2930,In_1802);
nor U348 (N_348,In_828,In_2182);
xnor U349 (N_349,In_1913,In_656);
or U350 (N_350,N_273,In_1301);
or U351 (N_351,In_1269,In_2869);
xnor U352 (N_352,N_108,In_178);
nand U353 (N_353,In_592,In_2391);
and U354 (N_354,In_1201,In_1589);
xor U355 (N_355,In_1732,N_134);
xor U356 (N_356,In_205,In_2557);
or U357 (N_357,In_2542,In_863);
or U358 (N_358,In_1824,In_2215);
nand U359 (N_359,N_286,In_2368);
and U360 (N_360,In_232,In_1794);
nor U361 (N_361,In_2300,N_44);
or U362 (N_362,In_1342,In_601);
nor U363 (N_363,In_83,In_2365);
nor U364 (N_364,In_1514,In_2737);
and U365 (N_365,In_770,In_1373);
or U366 (N_366,In_2632,In_1317);
or U367 (N_367,In_2207,In_2627);
xnor U368 (N_368,In_2457,In_323);
or U369 (N_369,In_1224,In_2311);
and U370 (N_370,In_1193,In_664);
or U371 (N_371,In_62,In_2383);
and U372 (N_372,In_1572,In_2563);
nand U373 (N_373,In_363,In_1994);
and U374 (N_374,In_476,N_299);
nand U375 (N_375,In_2235,In_2218);
xor U376 (N_376,In_1401,In_74);
or U377 (N_377,In_454,In_2583);
or U378 (N_378,In_1672,In_2758);
or U379 (N_379,In_1289,In_1992);
or U380 (N_380,In_1140,In_1771);
xnor U381 (N_381,In_1302,In_1503);
xnor U382 (N_382,N_131,In_1692);
nor U383 (N_383,In_2544,In_2057);
nor U384 (N_384,In_755,In_1040);
and U385 (N_385,In_1965,In_1162);
nand U386 (N_386,In_2496,N_140);
or U387 (N_387,In_416,In_1659);
nor U388 (N_388,In_2395,N_7);
and U389 (N_389,In_1154,In_2777);
xnor U390 (N_390,In_2993,In_1668);
xnor U391 (N_391,N_76,In_2847);
xnor U392 (N_392,In_2738,In_1479);
nor U393 (N_393,In_877,In_1279);
nand U394 (N_394,In_1137,In_1874);
nand U395 (N_395,In_491,N_175);
and U396 (N_396,In_2784,N_48);
nor U397 (N_397,In_1215,In_1083);
nand U398 (N_398,In_2343,In_520);
and U399 (N_399,In_1978,In_1327);
xnor U400 (N_400,In_1804,In_938);
nor U401 (N_401,In_1270,In_466);
or U402 (N_402,N_230,In_46);
nand U403 (N_403,In_1443,In_2531);
xnor U404 (N_404,In_709,In_676);
nor U405 (N_405,In_1740,N_258);
nand U406 (N_406,In_1465,In_2093);
or U407 (N_407,In_2252,In_1419);
or U408 (N_408,In_1466,In_885);
xnor U409 (N_409,In_1069,In_1197);
and U410 (N_410,In_365,In_1675);
nand U411 (N_411,In_126,In_1926);
nand U412 (N_412,In_1959,In_1314);
or U413 (N_413,In_2077,In_2955);
nand U414 (N_414,In_2063,In_2293);
or U415 (N_415,In_789,In_414);
nor U416 (N_416,In_2947,In_2141);
and U417 (N_417,In_1507,In_729);
nor U418 (N_418,In_1513,In_2863);
nor U419 (N_419,In_1782,In_2229);
xnor U420 (N_420,In_2159,In_2112);
nand U421 (N_421,In_2055,In_1781);
and U422 (N_422,In_1101,In_2671);
and U423 (N_423,In_1425,N_88);
nand U424 (N_424,In_407,In_2201);
nand U425 (N_425,In_2534,In_1236);
or U426 (N_426,In_1996,In_312);
xnor U427 (N_427,In_1089,In_510);
and U428 (N_428,In_855,In_2396);
nand U429 (N_429,N_142,In_1537);
nand U430 (N_430,In_2983,N_31);
and U431 (N_431,In_364,In_1047);
or U432 (N_432,In_2843,In_193);
and U433 (N_433,In_2769,In_2655);
nor U434 (N_434,In_396,In_2683);
nand U435 (N_435,In_973,In_1982);
or U436 (N_436,In_804,In_1473);
nand U437 (N_437,In_1126,In_426);
and U438 (N_438,In_2363,N_254);
or U439 (N_439,In_1506,In_1434);
and U440 (N_440,In_2154,In_859);
and U441 (N_441,In_1887,In_2725);
xor U442 (N_442,In_186,In_1451);
and U443 (N_443,N_298,In_2304);
xor U444 (N_444,In_2509,In_1072);
xnor U445 (N_445,In_762,In_2775);
nor U446 (N_446,In_633,In_422);
nand U447 (N_447,In_1893,In_1021);
xnor U448 (N_448,N_52,In_1426);
and U449 (N_449,In_2997,In_2624);
nand U450 (N_450,N_106,In_1956);
nand U451 (N_451,In_1206,In_2670);
xor U452 (N_452,In_1837,In_593);
nor U453 (N_453,In_950,In_2746);
xnor U454 (N_454,In_1878,In_2080);
nor U455 (N_455,In_882,In_1660);
or U456 (N_456,In_399,In_2034);
and U457 (N_457,In_528,In_2290);
and U458 (N_458,N_32,In_2537);
xnor U459 (N_459,In_114,In_2636);
xnor U460 (N_460,In_2259,In_1005);
or U461 (N_461,In_2170,In_2);
and U462 (N_462,In_707,In_880);
nand U463 (N_463,N_152,In_1060);
or U464 (N_464,In_1511,N_42);
nor U465 (N_465,In_776,In_2672);
and U466 (N_466,In_1142,In_1694);
and U467 (N_467,N_213,In_142);
and U468 (N_468,In_2433,In_811);
nand U469 (N_469,In_207,In_2511);
xor U470 (N_470,In_1531,N_72);
nor U471 (N_471,In_1115,In_1023);
nor U472 (N_472,In_2153,In_2826);
or U473 (N_473,In_522,In_185);
nand U474 (N_474,In_594,In_2908);
xor U475 (N_475,In_1135,In_1230);
or U476 (N_476,In_824,N_54);
nor U477 (N_477,In_2225,N_73);
or U478 (N_478,In_752,In_1458);
nor U479 (N_479,In_93,In_571);
nor U480 (N_480,In_2830,In_490);
or U481 (N_481,In_1476,In_2595);
or U482 (N_482,In_1724,In_2949);
and U483 (N_483,In_529,In_2532);
and U484 (N_484,In_5,In_172);
or U485 (N_485,In_1202,In_2565);
nand U486 (N_486,In_1057,In_2852);
nand U487 (N_487,In_497,In_896);
and U488 (N_488,In_393,In_53);
or U489 (N_489,In_2190,In_867);
xor U490 (N_490,In_1173,In_1587);
or U491 (N_491,In_1346,In_377);
and U492 (N_492,In_1169,In_1658);
or U493 (N_493,In_2945,In_180);
xnor U494 (N_494,In_745,In_775);
or U495 (N_495,In_1986,N_241);
xnor U496 (N_496,In_1504,In_1679);
or U497 (N_497,N_181,In_2044);
xnor U498 (N_498,In_1970,In_1575);
nand U499 (N_499,In_136,In_1110);
nor U500 (N_500,In_631,In_2592);
or U501 (N_501,In_1934,In_2498);
and U502 (N_502,In_1573,In_2249);
nor U503 (N_503,In_1370,In_146);
or U504 (N_504,In_671,In_1687);
or U505 (N_505,In_2197,In_2443);
and U506 (N_506,In_2256,In_1857);
nor U507 (N_507,In_901,In_2359);
xor U508 (N_508,In_2128,In_2060);
xnor U509 (N_509,In_646,N_111);
and U510 (N_510,In_615,In_1191);
nand U511 (N_511,In_166,N_125);
xnor U512 (N_512,In_240,In_2886);
nor U513 (N_513,In_2846,In_8);
xnor U514 (N_514,N_135,In_1280);
nand U515 (N_515,In_2317,In_1734);
xnor U516 (N_516,In_940,N_289);
and U517 (N_517,In_1227,In_1118);
nor U518 (N_518,In_386,In_227);
xor U519 (N_519,In_526,In_1628);
nor U520 (N_520,In_1014,In_1640);
or U521 (N_521,In_2600,In_598);
xnor U522 (N_522,N_129,In_1241);
nand U523 (N_523,In_1429,In_1098);
or U524 (N_524,In_328,In_2139);
nor U525 (N_525,In_1084,In_214);
nor U526 (N_526,In_106,N_293);
xor U527 (N_527,In_1697,In_1331);
xor U528 (N_528,In_2748,In_2601);
and U529 (N_529,In_1998,In_2065);
nor U530 (N_530,In_843,In_1744);
and U531 (N_531,In_273,N_237);
xor U532 (N_532,In_2192,N_86);
nor U533 (N_533,In_2347,In_1932);
nand U534 (N_534,In_911,In_793);
and U535 (N_535,In_1856,In_1367);
or U536 (N_536,N_58,N_64);
or U537 (N_537,In_9,In_1653);
nor U538 (N_538,In_2787,In_1927);
xnor U539 (N_539,In_97,N_126);
xor U540 (N_540,In_2477,In_1159);
and U541 (N_541,In_1712,In_1013);
nand U542 (N_542,In_2404,N_146);
or U543 (N_543,In_1593,In_1768);
and U544 (N_544,In_1937,In_2370);
nand U545 (N_545,In_1158,In_1848);
and U546 (N_546,N_112,In_744);
xor U547 (N_547,N_239,In_1349);
or U548 (N_548,In_29,N_1);
or U549 (N_549,In_125,In_2231);
or U550 (N_550,In_1606,In_891);
nor U551 (N_551,In_1065,In_1778);
and U552 (N_552,N_82,In_2119);
nor U553 (N_553,In_627,In_343);
and U554 (N_554,In_67,In_1916);
xnor U555 (N_555,In_682,In_688);
and U556 (N_556,In_1444,In_523);
nand U557 (N_557,In_873,In_181);
nor U558 (N_558,In_285,In_445);
or U559 (N_559,In_2373,In_224);
nand U560 (N_560,In_2555,In_1823);
nand U561 (N_561,In_2635,In_2138);
or U562 (N_562,In_2642,In_2513);
nand U563 (N_563,In_1397,In_292);
xor U564 (N_564,In_2280,In_2357);
and U565 (N_565,In_1850,In_2085);
and U566 (N_566,In_2559,In_1405);
or U567 (N_567,In_1727,In_519);
nor U568 (N_568,In_1052,In_1585);
or U569 (N_569,In_761,In_2039);
xor U570 (N_570,In_915,In_2204);
xnor U571 (N_571,In_1309,In_1111);
or U572 (N_572,In_1371,In_2824);
xor U573 (N_573,In_413,N_218);
and U574 (N_574,In_77,In_551);
nand U575 (N_575,In_1407,In_2665);
nor U576 (N_576,In_2931,In_194);
nor U577 (N_577,In_909,In_1664);
nand U578 (N_578,In_2613,In_1497);
xor U579 (N_579,In_1656,In_694);
or U580 (N_580,In_257,In_2133);
nand U581 (N_581,N_30,In_947);
and U582 (N_582,In_1231,In_2147);
or U583 (N_583,In_531,In_478);
or U584 (N_584,In_1035,In_1144);
nand U585 (N_585,N_204,In_2536);
and U586 (N_586,N_173,In_1155);
nand U587 (N_587,In_1307,N_211);
and U588 (N_588,In_639,In_1109);
nor U589 (N_589,In_972,In_2717);
xnor U590 (N_590,In_524,In_919);
xor U591 (N_591,In_152,In_815);
nand U592 (N_592,In_1276,In_2788);
xor U593 (N_593,In_1272,In_2126);
nor U594 (N_594,In_1210,In_1318);
xnor U595 (N_595,In_600,N_203);
or U596 (N_596,N_167,In_608);
or U597 (N_597,N_196,In_956);
xnor U598 (N_598,In_590,In_2268);
nor U599 (N_599,In_1352,In_2646);
xnor U600 (N_600,In_25,N_475);
xor U601 (N_601,In_2522,In_1106);
and U602 (N_602,In_1629,In_1024);
nand U603 (N_603,N_115,N_190);
xnor U604 (N_604,N_120,In_1050);
and U605 (N_605,N_468,In_102);
and U606 (N_606,N_574,In_652);
and U607 (N_607,In_2011,N_25);
and U608 (N_608,N_331,In_1552);
or U609 (N_609,In_999,In_2397);
and U610 (N_610,In_2466,In_233);
nor U611 (N_611,In_1652,In_86);
or U612 (N_612,In_2580,In_1056);
xor U613 (N_613,N_478,In_2202);
and U614 (N_614,In_802,In_1811);
nor U615 (N_615,N_2,In_1176);
nor U616 (N_616,In_2828,N_592);
and U617 (N_617,In_1160,In_2448);
and U618 (N_618,In_1123,In_2183);
nand U619 (N_619,In_1785,In_2538);
and U620 (N_620,In_640,In_1524);
nand U621 (N_621,N_366,In_870);
and U622 (N_622,N_572,In_300);
or U623 (N_623,In_2471,In_2101);
xor U624 (N_624,In_1381,N_197);
xnor U625 (N_625,In_764,In_2803);
nand U626 (N_626,In_980,In_1518);
xor U627 (N_627,N_518,In_2420);
xnor U628 (N_628,N_515,In_1590);
and U629 (N_629,In_2131,In_1719);
xor U630 (N_630,In_861,In_2422);
xnor U631 (N_631,In_2973,In_521);
nand U632 (N_632,N_520,In_1361);
and U633 (N_633,N_236,In_780);
xor U634 (N_634,In_372,N_153);
and U635 (N_635,In_1806,In_771);
xnor U636 (N_636,In_1051,N_410);
nand U637 (N_637,N_375,N_122);
and U638 (N_638,N_3,In_1625);
or U639 (N_639,N_311,In_820);
and U640 (N_640,In_129,In_2792);
and U641 (N_641,N_327,N_316);
nor U642 (N_642,In_1612,In_807);
or U643 (N_643,In_1636,N_70);
and U644 (N_644,In_945,N_455);
and U645 (N_645,In_2241,In_1877);
nor U646 (N_646,N_587,In_884);
nand U647 (N_647,In_1860,In_715);
and U648 (N_648,In_1409,N_416);
xor U649 (N_649,In_702,In_1639);
and U650 (N_650,In_2232,In_568);
xor U651 (N_651,In_2695,N_536);
xnor U652 (N_652,N_47,In_1898);
xor U653 (N_653,N_55,In_555);
and U654 (N_654,In_2321,In_347);
and U655 (N_655,In_210,In_1251);
or U656 (N_656,In_1822,In_2691);
or U657 (N_657,In_2814,In_2292);
nand U658 (N_658,In_1742,In_2878);
nand U659 (N_659,In_2680,In_1845);
nand U660 (N_660,In_2262,In_333);
nor U661 (N_661,N_309,In_1253);
xnor U662 (N_662,In_2301,In_1022);
xor U663 (N_663,N_95,In_1032);
nor U664 (N_664,In_1760,N_492);
or U665 (N_665,N_578,In_1470);
xor U666 (N_666,In_1413,In_2774);
and U667 (N_667,In_1990,N_75);
and U668 (N_668,In_2384,N_391);
and U669 (N_669,N_354,In_1164);
nand U670 (N_670,In_974,In_1477);
xnor U671 (N_671,In_541,In_15);
and U672 (N_672,In_623,N_502);
and U673 (N_673,In_61,In_1968);
or U674 (N_674,In_2326,In_1143);
nand U675 (N_675,In_1174,In_253);
or U676 (N_676,In_2074,In_55);
or U677 (N_677,In_2979,In_2109);
or U678 (N_678,In_2247,In_916);
nor U679 (N_679,N_144,In_2272);
and U680 (N_680,N_582,In_2185);
xor U681 (N_681,In_1054,In_2910);
and U682 (N_682,In_281,N_534);
xor U683 (N_683,In_87,N_481);
or U684 (N_684,N_406,In_987);
or U685 (N_685,In_112,In_1181);
nand U686 (N_686,In_2157,In_2560);
and U687 (N_687,In_2007,N_325);
nand U688 (N_688,N_418,In_1360);
or U689 (N_689,N_319,In_1515);
nor U690 (N_690,In_1059,N_247);
and U691 (N_691,In_1752,In_821);
nand U692 (N_692,In_2604,In_301);
or U693 (N_693,In_1412,In_583);
or U694 (N_694,In_2844,In_2586);
or U695 (N_695,In_704,In_645);
nand U696 (N_696,In_661,N_43);
xor U697 (N_697,In_2356,In_747);
and U698 (N_698,In_1063,N_97);
or U699 (N_699,In_2258,In_2075);
or U700 (N_700,In_1246,In_307);
xnor U701 (N_701,N_379,In_1237);
and U702 (N_702,In_2277,N_504);
nand U703 (N_703,N_36,In_266);
and U704 (N_704,In_1449,In_1);
xnor U705 (N_705,In_2102,N_506);
nor U706 (N_706,In_2961,In_1296);
nand U707 (N_707,In_2419,N_318);
xor U708 (N_708,N_399,N_491);
and U709 (N_709,In_314,In_1369);
or U710 (N_710,In_564,In_1320);
nor U711 (N_711,In_610,N_276);
nor U712 (N_712,In_2888,In_2603);
nor U713 (N_713,In_1859,N_113);
nor U714 (N_714,In_2230,In_2409);
nor U715 (N_715,In_0,In_160);
nor U716 (N_716,In_1427,In_2572);
nand U717 (N_717,In_2853,N_87);
nand U718 (N_718,In_2211,In_124);
or U719 (N_719,In_2884,In_267);
or U720 (N_720,In_970,In_946);
and U721 (N_721,In_294,In_1759);
nand U722 (N_722,In_1713,In_2943);
nor U723 (N_723,In_463,In_1690);
xnor U724 (N_724,In_284,N_377);
or U725 (N_725,In_504,In_2013);
nand U726 (N_726,N_498,In_1553);
or U727 (N_727,N_450,In_1936);
nand U728 (N_728,In_2442,In_2149);
and U729 (N_729,N_266,In_424);
nor U730 (N_730,In_1461,In_1493);
nand U731 (N_731,N_110,N_420);
nand U732 (N_732,In_395,In_2839);
nor U733 (N_733,In_2693,In_1907);
and U734 (N_734,In_998,In_2541);
nor U735 (N_735,In_100,N_100);
nor U736 (N_736,In_2188,In_1484);
nand U737 (N_737,In_1403,In_1087);
xor U738 (N_738,N_489,In_170);
or U739 (N_739,In_2010,In_1924);
nor U740 (N_740,In_982,In_1743);
xnor U741 (N_741,N_382,N_22);
or U742 (N_742,N_347,In_1471);
nor U743 (N_743,In_539,In_923);
xnor U744 (N_744,N_198,In_263);
or U745 (N_745,In_1648,N_249);
nor U746 (N_746,In_324,In_1464);
and U747 (N_747,N_500,In_1134);
nand U748 (N_748,In_1548,N_556);
or U749 (N_749,In_2686,In_1168);
nand U750 (N_750,In_1749,In_942);
xnor U751 (N_751,In_220,N_89);
or U752 (N_752,In_2340,In_1745);
xor U753 (N_753,N_361,In_1534);
and U754 (N_754,N_488,N_158);
xor U755 (N_755,In_1480,In_850);
or U756 (N_756,In_2882,In_2650);
nor U757 (N_757,In_2086,In_2621);
nand U758 (N_758,In_2577,N_162);
or U759 (N_759,In_387,In_585);
or U760 (N_760,In_350,N_314);
and U761 (N_761,N_501,In_1339);
and U762 (N_762,In_2493,N_105);
xnor U763 (N_763,In_2116,In_2091);
nand U764 (N_764,In_1306,In_1733);
xnor U765 (N_765,In_727,N_541);
or U766 (N_766,N_18,In_2467);
xnor U767 (N_767,In_1199,In_1728);
nand U768 (N_768,In_2859,N_51);
and U769 (N_769,N_529,In_1147);
and U770 (N_770,In_2307,In_2608);
or U771 (N_771,N_164,In_836);
or U772 (N_772,In_137,In_1061);
xnor U773 (N_773,In_887,In_2449);
nor U774 (N_774,In_695,In_1394);
nor U775 (N_775,In_1599,In_1294);
xor U776 (N_776,N_242,In_2582);
or U777 (N_777,In_1421,N_251);
nor U778 (N_778,In_1365,In_1151);
nand U779 (N_779,In_2829,In_122);
xor U780 (N_780,In_174,In_599);
and U781 (N_781,N_169,In_2514);
and U782 (N_782,In_1729,In_1356);
or U783 (N_783,In_1841,In_208);
or U784 (N_784,In_24,In_1963);
nand U785 (N_785,N_421,In_1821);
and U786 (N_786,In_2651,In_2306);
nor U787 (N_787,N_323,In_2025);
nand U788 (N_788,In_2417,In_1265);
and U789 (N_789,In_1554,In_2220);
and U790 (N_790,In_2896,In_778);
nor U791 (N_791,N_401,In_1010);
xnor U792 (N_792,N_404,N_244);
xnor U793 (N_793,N_365,In_474);
xor U794 (N_794,N_186,In_201);
nand U795 (N_795,In_1835,In_494);
nand U796 (N_796,In_2807,In_2911);
and U797 (N_797,In_1731,In_532);
xor U798 (N_798,In_2982,In_2193);
or U799 (N_799,In_732,In_489);
or U800 (N_800,N_41,N_372);
and U801 (N_801,N_99,In_1730);
xor U802 (N_802,In_1988,In_1748);
or U803 (N_803,In_2083,In_1977);
nor U804 (N_804,N_283,In_103);
xnor U805 (N_805,In_1577,In_1829);
nor U806 (N_806,In_1810,In_1341);
nand U807 (N_807,In_110,In_33);
xnor U808 (N_808,In_1223,N_4);
or U809 (N_809,In_1637,In_1200);
or U810 (N_810,In_513,In_316);
nor U811 (N_811,In_1912,In_2261);
nor U812 (N_812,In_516,N_147);
or U813 (N_813,In_1171,In_1340);
and U814 (N_814,In_1645,In_2305);
and U815 (N_815,In_609,In_1195);
or U816 (N_816,In_777,N_338);
nor U817 (N_817,In_1953,In_1528);
and U818 (N_818,In_1576,In_2458);
or U819 (N_819,N_364,In_2388);
nor U820 (N_820,In_2976,In_2390);
xor U821 (N_821,In_1019,In_879);
or U822 (N_822,In_2090,In_2981);
and U823 (N_823,In_2836,N_69);
xor U824 (N_824,In_151,In_2707);
and U825 (N_825,N_412,In_2521);
and U826 (N_826,In_1351,In_276);
and U827 (N_827,In_2038,In_1764);
nand U828 (N_828,In_1332,In_2647);
and U829 (N_829,In_56,In_1233);
xor U830 (N_830,In_183,N_426);
and U831 (N_831,In_2445,N_439);
nand U832 (N_832,In_726,In_1311);
nand U833 (N_833,In_971,In_509);
nor U834 (N_834,In_297,In_1558);
nor U835 (N_835,In_2243,N_136);
nor U836 (N_836,In_2809,N_558);
and U837 (N_837,N_21,In_358);
nor U838 (N_838,In_2639,In_2605);
or U839 (N_839,In_582,N_374);
nand U840 (N_840,In_359,N_539);
and U841 (N_841,N_270,In_1582);
nor U842 (N_842,N_60,In_2794);
nor U843 (N_843,In_1348,In_2804);
nor U844 (N_844,In_2889,In_1619);
or U845 (N_845,In_1773,In_2385);
xor U846 (N_846,N_551,In_2438);
nor U847 (N_847,In_2700,In_370);
nor U848 (N_848,In_1520,In_1437);
nor U849 (N_849,In_1222,In_91);
or U850 (N_850,In_2210,N_324);
xnor U851 (N_851,In_659,In_1457);
nor U852 (N_852,N_215,In_1252);
or U853 (N_853,In_1300,N_322);
or U854 (N_854,N_546,In_2121);
nand U855 (N_855,N_313,N_535);
and U856 (N_856,In_2564,N_66);
nand U857 (N_857,In_2622,N_476);
and U858 (N_858,In_2629,In_1762);
and U859 (N_859,In_2009,In_1839);
nand U860 (N_860,N_191,N_201);
nor U861 (N_861,In_2674,In_2996);
nor U862 (N_862,In_834,In_439);
nand U863 (N_863,In_2407,N_172);
xor U864 (N_864,N_560,In_728);
nand U865 (N_865,In_2142,In_2508);
nand U866 (N_866,In_2223,In_2135);
and U867 (N_867,In_1325,In_2245);
and U868 (N_868,N_559,In_2410);
xor U869 (N_869,N_553,N_444);
nor U870 (N_870,In_1902,N_415);
nor U871 (N_871,N_337,In_2614);
nor U872 (N_872,In_2386,In_2872);
and U873 (N_873,In_1682,In_578);
xor U874 (N_874,N_228,N_267);
nor U875 (N_875,In_700,In_930);
nor U876 (N_876,In_2281,N_573);
nand U877 (N_877,N_297,N_212);
or U878 (N_878,N_594,In_2348);
or U879 (N_879,N_177,N_261);
or U880 (N_880,In_153,In_1238);
nor U881 (N_881,In_2335,In_1776);
xnor U882 (N_882,In_1226,In_2546);
nor U883 (N_883,In_2282,N_459);
nand U884 (N_884,In_2336,In_357);
or U885 (N_885,In_2339,In_2762);
nor U886 (N_886,N_479,In_1819);
xor U887 (N_887,In_2660,N_373);
xor U888 (N_888,In_329,In_1131);
or U889 (N_889,In_2581,In_1739);
nor U890 (N_890,In_553,In_1081);
and U891 (N_891,In_1129,In_634);
or U892 (N_892,In_864,In_2985);
and U893 (N_893,In_2591,In_2160);
and U894 (N_894,In_2832,In_1250);
and U895 (N_895,N_287,In_1562);
xnor U896 (N_896,N_284,N_143);
or U897 (N_897,N_310,N_524);
xnor U898 (N_898,In_2736,In_1428);
nor U899 (N_899,In_2937,N_317);
nand U900 (N_900,N_769,N_383);
or U901 (N_901,In_1725,In_2929);
nor U902 (N_902,In_2001,In_1030);
xnor U903 (N_903,N_400,In_647);
nor U904 (N_904,In_409,In_1283);
xnor U905 (N_905,N_505,In_1881);
nor U906 (N_906,N_477,N_225);
nor U907 (N_907,In_1901,In_1505);
nand U908 (N_908,N_77,N_480);
nand U909 (N_909,In_1362,In_1053);
and U910 (N_910,In_2430,In_2690);
nor U911 (N_911,In_1406,N_78);
nor U912 (N_912,In_2702,In_783);
nand U913 (N_913,In_660,In_176);
and U914 (N_914,N_35,N_768);
and U915 (N_915,N_224,N_447);
and U916 (N_916,In_2875,N_831);
nor U917 (N_917,N_395,N_453);
nand U918 (N_918,In_75,In_2561);
nand U919 (N_919,In_547,In_1478);
xor U920 (N_920,N_511,In_1920);
and U921 (N_921,In_268,N_509);
nor U922 (N_922,N_694,In_1433);
nor U923 (N_923,N_868,N_92);
nand U924 (N_924,In_2260,N_429);
nand U925 (N_925,N_840,In_816);
or U926 (N_926,N_431,In_1239);
xnor U927 (N_927,In_1940,In_1096);
nand U928 (N_928,In_1240,In_2481);
nor U929 (N_929,In_2369,In_1693);
or U930 (N_930,In_1680,N_708);
and U931 (N_931,In_384,In_458);
or U932 (N_932,In_1295,In_392);
or U933 (N_933,In_111,In_1543);
nor U934 (N_934,In_1900,N_625);
xor U935 (N_935,In_1975,N_703);
nor U936 (N_936,In_2355,In_1468);
nor U937 (N_937,In_937,In_2666);
nand U938 (N_938,In_1248,In_825);
nor U939 (N_939,N_891,In_2634);
nand U940 (N_940,In_1828,N_790);
nand U941 (N_941,N_484,In_1036);
or U942 (N_942,N_121,In_2353);
nor U943 (N_943,In_334,In_1769);
nor U944 (N_944,N_654,In_2024);
or U945 (N_945,In_2813,In_1064);
and U946 (N_946,In_979,In_931);
nand U947 (N_947,In_271,In_1921);
or U948 (N_948,In_1102,In_769);
nand U949 (N_949,N_79,N_823);
and U950 (N_950,In_2716,N_351);
nor U951 (N_951,N_613,In_1564);
nor U952 (N_952,In_951,In_1337);
xor U953 (N_953,In_2837,N_295);
or U954 (N_954,N_802,In_1257);
or U955 (N_955,N_789,N_666);
nor U956 (N_956,N_260,N_893);
and U957 (N_957,In_1441,In_2845);
nand U958 (N_958,In_1467,N_850);
nand U959 (N_959,In_2068,In_200);
nor U960 (N_960,In_1622,In_2319);
nor U961 (N_961,In_2838,In_1305);
and U962 (N_962,N_405,N_819);
xnor U963 (N_963,In_197,N_606);
or U964 (N_964,N_208,In_2342);
xor U965 (N_965,N_233,In_222);
nor U966 (N_966,In_2724,In_2726);
and U967 (N_967,N_889,In_786);
and U968 (N_968,In_2288,In_1042);
nor U969 (N_969,In_2963,In_603);
nor U970 (N_970,In_1869,In_308);
nand U971 (N_971,In_415,N_446);
nand U972 (N_972,In_2212,N_302);
xnor U973 (N_973,In_2713,In_1673);
xor U974 (N_974,In_948,N_715);
xor U975 (N_975,In_1941,In_2840);
and U976 (N_976,In_881,In_2759);
or U977 (N_977,In_2492,In_2915);
xor U978 (N_978,N_248,In_390);
xnor U979 (N_979,In_1655,In_1885);
xnor U980 (N_980,In_1136,N_684);
nor U981 (N_981,In_746,In_2168);
or U982 (N_982,N_788,N_305);
and U983 (N_983,In_1529,In_2447);
and U984 (N_984,In_1358,N_853);
xor U985 (N_985,N_423,In_408);
or U986 (N_986,N_628,N_332);
or U987 (N_987,In_1297,In_1359);
and U988 (N_988,N_371,In_368);
nand U989 (N_989,In_2658,In_150);
and U990 (N_990,In_1701,In_2216);
and U991 (N_991,In_2178,In_2461);
and U992 (N_992,In_2456,In_2654);
nand U993 (N_993,N_860,N_430);
xnor U994 (N_994,N_639,N_839);
nor U995 (N_995,N_306,In_2520);
xnor U996 (N_996,N_892,N_693);
xnor U997 (N_997,In_1838,In_2338);
and U998 (N_998,In_964,In_1676);
xnor U999 (N_999,In_1186,In_968);
and U1000 (N_1000,N_223,N_243);
nand U1001 (N_1001,N_691,In_2372);
nand U1002 (N_1002,In_2952,In_1547);
nand U1003 (N_1003,In_1004,In_379);
and U1004 (N_1004,In_2181,In_411);
xor U1005 (N_1005,In_2236,In_2568);
nor U1006 (N_1006,In_40,N_549);
or U1007 (N_1007,In_321,In_2270);
xnor U1008 (N_1008,N_188,N_595);
or U1009 (N_1009,In_686,N_847);
nor U1010 (N_1010,In_1261,In_385);
and U1011 (N_1011,N_760,In_2052);
and U1012 (N_1012,In_2144,N_630);
nand U1013 (N_1013,N_820,In_933);
or U1014 (N_1014,In_2818,In_2767);
nor U1015 (N_1015,In_1183,In_711);
nor U1016 (N_1016,In_2974,N_680);
nor U1017 (N_1017,N_866,In_1055);
nand U1018 (N_1018,In_130,In_621);
nand U1019 (N_1019,In_810,In_2661);
nand U1020 (N_1020,N_192,N_897);
xor U1021 (N_1021,In_1942,In_459);
and U1022 (N_1022,In_2607,In_471);
or U1023 (N_1023,In_2637,In_1800);
and U1024 (N_1024,N_116,In_543);
nand U1025 (N_1025,In_1737,In_1805);
xnor U1026 (N_1026,In_845,In_353);
or U1027 (N_1027,N_754,In_2079);
or U1028 (N_1028,In_2800,N_470);
and U1029 (N_1029,In_1044,In_1062);
xnor U1030 (N_1030,In_1871,In_1814);
xor U1031 (N_1031,In_52,In_1232);
xor U1032 (N_1032,In_420,In_1922);
and U1033 (N_1033,N_861,In_2898);
and U1034 (N_1034,N_217,N_161);
nor U1035 (N_1035,In_2662,In_2358);
nand U1036 (N_1036,In_1017,N_852);
xor U1037 (N_1037,In_1266,In_1809);
or U1038 (N_1038,In_2012,In_2566);
nor U1039 (N_1039,In_1383,In_1067);
nand U1040 (N_1040,In_1377,In_2593);
and U1041 (N_1041,N_575,In_1396);
xor U1042 (N_1042,In_2968,In_641);
nand U1043 (N_1043,In_2312,In_41);
and U1044 (N_1044,N_114,In_518);
or U1045 (N_1045,In_26,N_646);
nand U1046 (N_1046,In_1408,In_1735);
nand U1047 (N_1047,N_880,In_2594);
nor U1048 (N_1048,In_1928,In_766);
nor U1049 (N_1049,N_508,In_655);
or U1050 (N_1050,In_540,In_2917);
nand U1051 (N_1051,In_658,In_1284);
and U1052 (N_1052,N_109,In_2951);
xnor U1053 (N_1053,N_568,N_490);
nand U1054 (N_1054,In_719,N_59);
xor U1055 (N_1055,N_707,In_483);
and U1056 (N_1056,In_2186,In_65);
or U1057 (N_1057,In_57,N_733);
and U1058 (N_1058,In_1379,In_809);
and U1059 (N_1059,N_156,N_829);
xor U1060 (N_1060,N_528,In_932);
nand U1061 (N_1061,In_1925,In_693);
nand U1062 (N_1062,In_544,In_2751);
and U1063 (N_1063,In_2095,In_2200);
or U1064 (N_1064,In_1757,In_1517);
and U1065 (N_1065,In_710,In_1626);
xor U1066 (N_1066,In_2028,In_2150);
xnor U1067 (N_1067,N_321,N_638);
nand U1068 (N_1068,N_397,In_1758);
nand U1069 (N_1069,N_84,In_589);
nor U1070 (N_1070,N_485,In_2415);
and U1071 (N_1071,In_2299,In_862);
and U1072 (N_1072,In_2209,In_1345);
or U1073 (N_1073,N_329,N_497);
and U1074 (N_1074,In_1657,In_939);
xnor U1075 (N_1075,In_120,N_333);
xnor U1076 (N_1076,In_2977,In_118);
xor U1077 (N_1077,N_53,In_239);
nor U1078 (N_1078,N_235,N_28);
or U1079 (N_1079,In_2289,N_487);
or U1080 (N_1080,In_2273,In_2757);
nand U1081 (N_1081,In_1039,In_2037);
xor U1082 (N_1082,In_1933,N_620);
or U1083 (N_1083,In_2203,N_8);
nand U1084 (N_1084,N_895,N_803);
nand U1085 (N_1085,N_658,N_640);
nand U1086 (N_1086,In_2350,In_244);
and U1087 (N_1087,In_1382,In_2644);
and U1088 (N_1088,In_2161,In_2584);
xor U1089 (N_1089,N_163,In_1662);
and U1090 (N_1090,N_685,In_431);
nor U1091 (N_1091,In_47,In_2337);
xor U1092 (N_1092,N_380,N_711);
nor U1093 (N_1093,N_645,In_669);
and U1094 (N_1094,In_1574,In_790);
nand U1095 (N_1095,In_2957,In_470);
or U1096 (N_1096,In_1268,In_1689);
or U1097 (N_1097,In_1644,In_177);
xor U1098 (N_1098,In_1031,N_597);
xnor U1099 (N_1099,In_833,N_813);
nor U1100 (N_1100,In_1707,N_778);
nor U1101 (N_1101,N_585,In_402);
xnor U1102 (N_1102,In_835,N_782);
xnor U1103 (N_1103,In_1586,In_336);
and U1104 (N_1104,N_890,In_1588);
and U1105 (N_1105,In_2679,In_2320);
nand U1106 (N_1106,In_2098,In_7);
nor U1107 (N_1107,In_1611,In_818);
and U1108 (N_1108,In_255,In_2708);
xor U1109 (N_1109,In_1872,In_1962);
and U1110 (N_1110,In_768,In_2529);
nand U1111 (N_1111,N_644,In_115);
xor U1112 (N_1112,In_733,In_2374);
nand U1113 (N_1113,N_815,In_1353);
nand U1114 (N_1114,In_2224,In_2264);
and U1115 (N_1115,In_1113,In_1938);
and U1116 (N_1116,N_150,In_760);
nand U1117 (N_1117,N_748,N_403);
and U1118 (N_1118,In_2694,In_2239);
xor U1119 (N_1119,N_221,N_653);
and U1120 (N_1120,N_83,In_173);
xnor U1121 (N_1121,In_706,In_369);
xnor U1122 (N_1122,In_1980,In_990);
nand U1123 (N_1123,In_917,N_101);
xor U1124 (N_1124,In_1393,In_1843);
xnor U1125 (N_1125,In_2867,In_871);
and U1126 (N_1126,N_824,In_2575);
and U1127 (N_1127,In_801,N_346);
and U1128 (N_1128,In_1875,In_282);
xnor U1129 (N_1129,In_1438,N_687);
xnor U1130 (N_1130,In_595,In_1249);
nor U1131 (N_1131,N_465,In_242);
nand U1132 (N_1132,In_2042,N_238);
or U1133 (N_1133,In_1633,N_837);
nand U1134 (N_1134,In_577,In_280);
and U1135 (N_1135,In_2953,In_2483);
nand U1136 (N_1136,In_1533,In_1820);
xor U1137 (N_1137,In_1212,N_626);
xor U1138 (N_1138,In_1945,In_2478);
nand U1139 (N_1139,In_2525,In_161);
nor U1140 (N_1140,N_751,In_2950);
or U1141 (N_1141,N_449,In_2003);
xor U1142 (N_1142,In_808,In_876);
or U1143 (N_1143,N_525,N_442);
and U1144 (N_1144,N_608,N_0);
and U1145 (N_1145,In_1536,In_517);
or U1146 (N_1146,In_2811,In_2283);
nand U1147 (N_1147,N_647,In_1834);
and U1148 (N_1148,N_189,In_1825);
nand U1149 (N_1149,N_672,In_944);
nor U1150 (N_1150,In_1099,In_230);
xnor U1151 (N_1151,In_351,In_1972);
and U1152 (N_1152,In_2323,In_722);
and U1153 (N_1153,N_616,N_178);
and U1154 (N_1154,In_192,N_352);
xor U1155 (N_1155,In_456,In_1460);
xnor U1156 (N_1156,In_1635,In_1519);
nand U1157 (N_1157,N_74,In_814);
or U1158 (N_1158,In_2556,N_6);
nand U1159 (N_1159,N_682,N_166);
nor U1160 (N_1160,N_141,In_1324);
xor U1161 (N_1161,In_849,In_2587);
nor U1162 (N_1162,In_2421,In_277);
and U1163 (N_1163,In_82,In_156);
nand U1164 (N_1164,In_757,In_138);
nand U1165 (N_1165,In_2081,In_561);
nor U1166 (N_1166,In_1436,In_441);
nor U1167 (N_1167,In_2002,N_117);
xor U1168 (N_1168,N_818,In_1455);
nor U1169 (N_1169,N_149,In_748);
nor U1170 (N_1170,N_272,N_214);
xor U1171 (N_1171,In_2936,N_210);
or U1172 (N_1172,N_884,In_1846);
nor U1173 (N_1173,In_2050,In_1216);
nand U1174 (N_1174,N_734,In_383);
and U1175 (N_1175,In_1196,In_2488);
xnor U1176 (N_1176,N_554,In_1746);
and U1177 (N_1177,N_776,In_64);
nand U1178 (N_1178,N_530,N_801);
nor U1179 (N_1179,In_1958,N_544);
nor U1180 (N_1180,N_737,N_826);
nand U1181 (N_1181,N_304,N_845);
nand U1182 (N_1182,In_1454,N_552);
xor U1183 (N_1183,N_567,In_1674);
nor U1184 (N_1184,In_2512,In_43);
xnor U1185 (N_1185,N_130,In_2431);
xor U1186 (N_1186,In_2389,In_1581);
nor U1187 (N_1187,In_278,N_424);
nand U1188 (N_1188,In_1578,In_203);
nor U1189 (N_1189,In_1892,In_1432);
xor U1190 (N_1190,In_953,N_798);
nor U1191 (N_1191,In_2427,In_2698);
nand U1192 (N_1192,In_1947,In_2735);
or U1193 (N_1193,In_1354,N_63);
and U1194 (N_1194,In_1119,In_168);
or U1195 (N_1195,In_1194,In_1614);
or U1196 (N_1196,In_2165,N_673);
nand U1197 (N_1197,In_2827,N_200);
xor U1198 (N_1198,N_34,In_962);
nand U1199 (N_1199,In_1418,In_261);
or U1200 (N_1200,N_1048,N_588);
nand U1201 (N_1201,N_665,In_2865);
xnor U1202 (N_1202,N_80,In_2539);
and U1203 (N_1203,N_978,In_189);
xor U1204 (N_1204,In_188,In_1795);
and U1205 (N_1205,In_1999,In_2912);
nor U1206 (N_1206,In_2444,N_259);
or U1207 (N_1207,N_686,N_727);
xor U1208 (N_1208,In_2965,In_2049);
or U1209 (N_1209,N_435,N_1178);
xor U1210 (N_1210,In_2452,In_1844);
nor U1211 (N_1211,In_2739,N_1181);
nor U1212 (N_1212,N_636,N_633);
nand U1213 (N_1213,In_705,N_519);
and U1214 (N_1214,In_259,In_2752);
nand U1215 (N_1215,In_1190,In_1705);
or U1216 (N_1216,In_505,N_357);
nor U1217 (N_1217,In_1350,N_1108);
xor U1218 (N_1218,N_454,In_997);
nand U1219 (N_1219,In_187,In_298);
or U1220 (N_1220,In_1891,N_605);
and U1221 (N_1221,N_637,N_1028);
xor U1222 (N_1222,In_290,N_512);
nor U1223 (N_1223,N_94,In_1817);
or U1224 (N_1224,In_1070,In_1299);
or U1225 (N_1225,N_874,In_1424);
or U1226 (N_1226,In_2146,N_10);
nor U1227 (N_1227,In_98,In_2313);
or U1228 (N_1228,N_894,In_195);
xnor U1229 (N_1229,N_951,N_859);
or U1230 (N_1230,N_303,In_2939);
and U1231 (N_1231,In_1243,In_1288);
nor U1232 (N_1232,N_486,In_1245);
nand U1233 (N_1233,N_877,In_2935);
nand U1234 (N_1234,In_1456,In_319);
and U1235 (N_1235,In_978,N_791);
nor U1236 (N_1236,N_12,N_483);
xnor U1237 (N_1237,N_1087,In_311);
nand U1238 (N_1238,In_2053,N_696);
and U1239 (N_1239,N_879,N_849);
nand U1240 (N_1240,In_2728,N_467);
nand U1241 (N_1241,In_1613,N_1094);
xnor U1242 (N_1242,In_147,In_713);
nor U1243 (N_1243,N_1060,N_729);
and U1244 (N_1244,In_16,In_2412);
xor U1245 (N_1245,In_211,N_1013);
xor U1246 (N_1246,N_596,In_2640);
xnor U1247 (N_1247,In_1816,In_1976);
or U1248 (N_1248,In_1122,In_2495);
nand U1249 (N_1249,In_2502,In_2325);
xor U1250 (N_1250,N_958,In_1905);
xor U1251 (N_1251,N_906,In_238);
or U1252 (N_1252,N_1192,In_326);
nand U1253 (N_1253,In_2822,In_899);
nand U1254 (N_1254,N_205,N_763);
and U1255 (N_1255,In_1000,N_443);
and U1256 (N_1256,N_1129,In_1338);
nand U1257 (N_1257,In_2842,N_947);
xnor U1258 (N_1258,In_2254,In_1789);
and U1259 (N_1259,In_1702,In_2194);
nor U1260 (N_1260,In_2783,In_797);
or U1261 (N_1261,N_1024,In_2597);
nand U1262 (N_1262,N_842,In_269);
nand U1263 (N_1263,N_335,N_974);
xor U1264 (N_1264,N_67,In_683);
nor U1265 (N_1265,N_1172,N_1164);
nor U1266 (N_1266,N_246,N_876);
xor U1267 (N_1267,In_2734,In_76);
xnor U1268 (N_1268,N_902,In_2199);
nand U1269 (N_1269,N_780,In_1995);
nor U1270 (N_1270,In_678,N_655);
xor U1271 (N_1271,N_627,In_685);
nor U1272 (N_1272,N_517,N_937);
nand U1273 (N_1273,In_1285,N_216);
and U1274 (N_1274,In_2519,In_206);
nor U1275 (N_1275,In_14,In_1770);
nor U1276 (N_1276,In_2105,In_2805);
or U1277 (N_1277,In_912,N_1075);
or U1278 (N_1278,In_1964,In_2956);
xnor U1279 (N_1279,In_1561,In_779);
or U1280 (N_1280,In_50,In_1736);
and U1281 (N_1281,N_1134,In_1255);
nand U1282 (N_1282,N_670,In_1984);
nand U1283 (N_1283,In_908,In_626);
nand U1284 (N_1284,N_744,In_1501);
or U1285 (N_1285,N_376,N_138);
and U1286 (N_1286,In_1671,N_288);
or U1287 (N_1287,In_341,N_643);
nand U1288 (N_1288,N_1147,In_670);
or U1289 (N_1289,N_956,In_1670);
and U1290 (N_1290,N_29,In_1310);
nor U1291 (N_1291,N_368,N_792);
and U1292 (N_1292,In_1075,N_973);
and U1293 (N_1293,N_1090,In_1569);
nand U1294 (N_1294,N_770,N_721);
nand U1295 (N_1295,N_773,In_2573);
and U1296 (N_1296,In_2219,In_35);
or U1297 (N_1297,N_783,In_2004);
and U1298 (N_1298,N_521,N_699);
nand U1299 (N_1299,In_1918,In_2266);
nor U1300 (N_1300,In_2115,N_1143);
nor U1301 (N_1301,In_1526,In_619);
nand U1302 (N_1302,In_889,In_2554);
and U1303 (N_1303,N_701,N_262);
xor U1304 (N_1304,In_902,N_918);
nor U1305 (N_1305,N_878,N_983);
nor U1306 (N_1306,N_864,In_2631);
and U1307 (N_1307,In_1711,In_2711);
nand U1308 (N_1308,N_724,N_772);
and U1309 (N_1309,N_274,In_1716);
nand U1310 (N_1310,In_2015,N_690);
xor U1311 (N_1311,N_1041,In_2172);
and U1312 (N_1312,N_875,N_320);
nand U1313 (N_1313,In_171,N_1165);
nand U1314 (N_1314,N_920,N_398);
xnor U1315 (N_1315,N_1023,N_564);
nor U1316 (N_1316,N_604,In_1211);
xnor U1317 (N_1317,In_2072,In_2545);
nand U1318 (N_1318,N_330,In_632);
or U1319 (N_1319,In_2324,N_623);
and U1320 (N_1320,In_260,N_787);
nand U1321 (N_1321,In_910,In_1128);
xor U1322 (N_1322,In_1897,N_960);
and U1323 (N_1323,N_33,N_635);
or U1324 (N_1324,N_547,N_939);
nand U1325 (N_1325,N_46,N_954);
or U1326 (N_1326,N_433,N_1115);
nand U1327 (N_1327,In_425,N_735);
or U1328 (N_1328,In_638,N_1195);
or U1329 (N_1329,In_1411,N_1007);
nor U1330 (N_1330,In_1414,N_1082);
nand U1331 (N_1331,N_422,N_1183);
nor U1332 (N_1332,In_1836,N_1176);
and U1333 (N_1333,In_1509,N_901);
xnor U1334 (N_1334,N_496,In_723);
nand U1335 (N_1335,In_2125,N_1074);
and U1336 (N_1336,N_1059,N_615);
and U1337 (N_1337,N_39,In_2970);
nand U1338 (N_1338,In_2771,In_1002);
and U1339 (N_1339,In_84,In_2184);
nand U1340 (N_1340,In_1646,N_1029);
xnor U1341 (N_1341,N_1015,In_2460);
and U1342 (N_1342,In_2802,N_903);
or U1343 (N_1343,In_1796,In_584);
and U1344 (N_1344,In_913,In_236);
and U1345 (N_1345,In_635,In_1584);
nor U1346 (N_1346,In_1873,N_107);
and U1347 (N_1347,N_1070,N_93);
and U1348 (N_1348,In_629,N_1117);
and U1349 (N_1349,In_1082,N_1104);
and U1350 (N_1350,N_576,In_2515);
xor U1351 (N_1351,N_132,In_554);
or U1352 (N_1352,N_752,In_2361);
nor U1353 (N_1353,In_2296,N_339);
or U1354 (N_1354,In_374,In_2451);
or U1355 (N_1355,N_793,In_2244);
and U1356 (N_1356,N_301,In_674);
nor U1357 (N_1357,N_848,In_127);
xnor U1358 (N_1358,N_1006,In_73);
and U1359 (N_1359,In_2714,In_936);
nand U1360 (N_1360,In_1483,In_1957);
xnor U1361 (N_1361,N_1020,N_953);
xnor U1362 (N_1362,N_38,N_1168);
nand U1363 (N_1363,In_2727,N_292);
xor U1364 (N_1364,In_2494,In_1632);
and U1365 (N_1365,In_375,In_1647);
nor U1366 (N_1366,N_904,N_1145);
nand U1367 (N_1367,In_378,N_1003);
nand U1368 (N_1368,N_702,In_1775);
and U1369 (N_1369,In_1389,N_65);
and U1370 (N_1370,In_159,N_1047);
nor U1371 (N_1371,N_464,In_2967);
nand U1372 (N_1372,N_976,In_2806);
xnor U1373 (N_1373,In_1322,N_1190);
nor U1374 (N_1374,N_312,In_588);
or U1375 (N_1375,N_57,In_148);
and U1376 (N_1376,N_621,In_788);
xnor U1377 (N_1377,N_590,N_503);
xnor U1378 (N_1378,In_1527,In_283);
or U1379 (N_1379,In_2902,N_1066);
xor U1380 (N_1380,In_1761,N_825);
xnor U1381 (N_1381,In_1714,In_2550);
nand U1382 (N_1382,In_2934,In_591);
and U1383 (N_1383,N_821,In_2641);
xnor U1384 (N_1384,N_614,In_254);
or U1385 (N_1385,In_2978,N_786);
and U1386 (N_1386,In_2242,N_1163);
and U1387 (N_1387,In_1376,N_602);
xor U1388 (N_1388,N_1130,In_251);
nand U1389 (N_1389,N_264,N_624);
or U1390 (N_1390,In_354,N_674);
or U1391 (N_1391,In_217,N_1174);
and U1392 (N_1392,N_168,In_1148);
xor U1393 (N_1393,N_1053,N_899);
and U1394 (N_1394,In_2171,In_1952);
or U1395 (N_1395,N_277,N_118);
nor U1396 (N_1396,In_868,In_607);
and U1397 (N_1397,In_1213,N_870);
or U1398 (N_1398,N_678,N_1105);
nor U1399 (N_1399,In_243,In_2946);
and U1400 (N_1400,In_1600,N_1162);
or U1401 (N_1401,N_256,In_2099);
nor U1402 (N_1402,N_955,In_2030);
nand U1403 (N_1403,N_240,In_611);
or U1404 (N_1404,In_1609,N_651);
xor U1405 (N_1405,In_2021,In_734);
nor U1406 (N_1406,N_671,In_1095);
nor U1407 (N_1407,N_617,In_920);
xnor U1408 (N_1408,In_673,In_2816);
nand U1409 (N_1409,In_2772,In_692);
or U1410 (N_1410,In_738,N_1169);
xor U1411 (N_1411,N_669,In_1906);
nor U1412 (N_1412,N_814,In_587);
nand U1413 (N_1413,In_1717,N_1067);
and U1414 (N_1414,N_1144,In_2413);
and U1415 (N_1415,In_1715,N_1131);
and U1416 (N_1416,N_731,In_2255);
nand U1417 (N_1417,In_888,In_2392);
xor U1418 (N_1418,In_2588,In_2928);
or U1419 (N_1419,In_397,N_532);
nand U1420 (N_1420,N_1045,N_182);
xor U1421 (N_1421,N_473,N_1055);
and U1422 (N_1422,In_2441,In_2893);
nand U1423 (N_1423,N_545,N_387);
and U1424 (N_1424,In_2574,In_1290);
or U1425 (N_1425,In_2709,In_1882);
and U1426 (N_1426,In_2127,N_747);
and U1427 (N_1427,In_2633,In_538);
or U1428 (N_1428,In_1708,In_2114);
nor U1429 (N_1429,N_531,In_1567);
xor U1430 (N_1430,In_2920,N_856);
xnor U1431 (N_1431,In_1849,N_362);
nor U1432 (N_1432,N_1199,N_982);
nand U1433 (N_1433,In_1011,In_247);
nand U1434 (N_1434,N_928,In_60);
or U1435 (N_1435,N_1138,In_1326);
and U1436 (N_1436,N_432,In_1388);
nor U1437 (N_1437,In_1780,In_133);
nor U1438 (N_1438,N_367,N_1170);
xor U1439 (N_1439,In_410,N_171);
and U1440 (N_1440,In_1888,In_558);
nand U1441 (N_1441,N_1078,N_315);
or U1442 (N_1442,N_96,In_822);
nand U1443 (N_1443,In_2155,N_607);
and U1444 (N_1444,N_151,N_589);
or U1445 (N_1445,In_2437,In_2450);
nand U1446 (N_1446,In_965,N_940);
and U1447 (N_1447,In_1951,In_225);
xor U1448 (N_1448,N_1193,In_1217);
and U1449 (N_1449,In_287,N_300);
xnor U1450 (N_1450,In_2986,In_2487);
and U1451 (N_1451,In_2795,N_1046);
nand U1452 (N_1452,N_445,In_179);
and U1453 (N_1453,N_740,In_508);
nor U1454 (N_1454,In_525,In_2819);
and U1455 (N_1455,In_1685,In_1271);
nor U1456 (N_1456,In_2346,In_2862);
nor U1457 (N_1457,In_1391,N_1180);
xnor U1458 (N_1458,In_1703,N_91);
xnor U1459 (N_1459,N_809,In_1416);
nor U1460 (N_1460,N_562,N_611);
nor U1461 (N_1461,N_1069,In_1751);
xnor U1462 (N_1462,In_154,In_332);
nor U1463 (N_1463,N_194,N_157);
nor U1464 (N_1464,N_386,In_1025);
xnor U1465 (N_1465,In_2770,In_1258);
nand U1466 (N_1466,N_882,In_1334);
xnor U1467 (N_1467,In_485,In_23);
and U1468 (N_1468,In_1863,N_1103);
nand U1469 (N_1469,In_2971,N_1014);
nor U1470 (N_1470,In_2999,In_736);
xor U1471 (N_1471,N_863,In_265);
or U1472 (N_1472,N_913,N_550);
and U1473 (N_1473,In_2468,In_1048);
nand U1474 (N_1474,In_1943,In_2684);
xor U1475 (N_1475,In_548,In_1813);
and U1476 (N_1476,N_764,In_2630);
and U1477 (N_1477,In_2815,N_438);
xor U1478 (N_1478,N_966,In_2851);
xnor U1479 (N_1479,In_1944,N_428);
or U1480 (N_1480,N_975,N_828);
xor U1481 (N_1481,N_334,N_13);
nand U1482 (N_1482,In_2237,N_499);
xnor U1483 (N_1483,N_948,N_1177);
nand U1484 (N_1484,In_10,In_2810);
xnor U1485 (N_1485,In_2158,N_336);
xnor U1486 (N_1486,In_759,N_1051);
and U1487 (N_1487,In_1993,In_1939);
nand U1488 (N_1488,In_2377,In_1495);
nor U1489 (N_1489,In_1228,N_448);
or U1490 (N_1490,In_653,N_206);
nor U1491 (N_1491,In_2287,In_2944);
or U1492 (N_1492,In_2111,In_1105);
xnor U1493 (N_1493,N_698,N_1123);
and U1494 (N_1494,In_2274,N_1175);
and U1495 (N_1495,N_1196,In_2530);
or U1496 (N_1496,N_1001,In_832);
or U1497 (N_1497,N_970,N_563);
xnor U1498 (N_1498,In_500,In_758);
nor U1499 (N_1499,In_690,In_800);
and U1500 (N_1500,N_1152,In_306);
xnor U1501 (N_1501,In_371,In_2491);
xor U1502 (N_1502,In_215,N_413);
and U1503 (N_1503,N_961,In_1738);
xor U1504 (N_1504,In_560,In_1842);
xnor U1505 (N_1505,N_1118,N_1073);
and U1506 (N_1506,N_579,In_1754);
or U1507 (N_1507,N_618,In_703);
or U1508 (N_1508,In_149,N_1121);
nand U1509 (N_1509,In_898,N_527);
xnor U1510 (N_1510,In_1608,N_1448);
or U1511 (N_1511,N_1217,N_1189);
nand U1512 (N_1512,In_2510,N_758);
nand U1513 (N_1513,In_1667,In_1565);
xor U1514 (N_1514,In_2474,N_660);
nor U1515 (N_1515,In_2959,N_1461);
or U1516 (N_1516,In_751,In_2701);
and U1517 (N_1517,N_1287,N_836);
and U1518 (N_1518,In_842,In_2400);
xor U1519 (N_1519,N_601,N_1468);
xnor U1520 (N_1520,In_1008,N_1339);
nand U1521 (N_1521,N_998,N_1246);
or U1522 (N_1522,In_143,In_1991);
and U1523 (N_1523,In_469,N_1000);
nor U1524 (N_1524,In_2187,N_469);
nand U1525 (N_1525,N_1083,N_49);
nand U1526 (N_1526,N_723,In_2710);
and U1527 (N_1527,N_629,In_51);
nand U1528 (N_1528,N_1351,In_391);
xor U1529 (N_1529,N_943,In_1833);
nor U1530 (N_1530,N_1459,N_681);
xnor U1531 (N_1531,N_85,N_1248);
nor U1532 (N_1532,N_1283,In_229);
and U1533 (N_1533,N_1438,In_854);
and U1534 (N_1534,N_165,N_999);
and U1535 (N_1535,N_806,N_1101);
and U1536 (N_1536,N_381,N_1457);
nor U1537 (N_1537,N_98,N_1489);
xnor U1538 (N_1538,In_2625,N_179);
xnor U1539 (N_1539,In_1208,N_972);
and U1540 (N_1540,N_810,In_837);
nor U1541 (N_1541,N_984,N_1188);
or U1542 (N_1542,N_466,In_1177);
and U1543 (N_1543,N_1484,In_874);
or U1544 (N_1544,N_268,N_1379);
nand U1545 (N_1545,In_1380,N_1295);
nand U1546 (N_1546,N_855,N_533);
nand U1547 (N_1547,In_628,N_1424);
or U1548 (N_1548,In_2140,In_310);
or U1549 (N_1549,In_1185,N_1497);
xor U1550 (N_1550,In_2322,In_1831);
or U1551 (N_1551,N_857,N_1308);
nand U1552 (N_1552,N_1470,N_1280);
or U1553 (N_1553,In_712,In_580);
or U1554 (N_1554,N_931,In_27);
nand U1555 (N_1555,In_132,N_648);
or U1556 (N_1556,In_2786,N_676);
and U1557 (N_1557,In_895,N_944);
or U1558 (N_1558,In_2914,In_2432);
xor U1559 (N_1559,N_1453,N_1112);
xor U1560 (N_1560,N_718,In_2706);
or U1561 (N_1561,N_160,N_1033);
or U1562 (N_1562,N_1396,In_851);
nor U1563 (N_1563,N_742,In_2820);
or U1564 (N_1564,In_2453,In_2880);
or U1565 (N_1565,N_832,In_2667);
xor U1566 (N_1566,In_643,In_1205);
or U1567 (N_1567,In_718,In_1704);
nand U1568 (N_1568,In_434,N_474);
nor U1569 (N_1569,In_2371,N_1186);
and U1570 (N_1570,N_1194,N_1464);
xor U1571 (N_1571,N_1088,N_1392);
xnor U1572 (N_1572,N_1210,N_437);
xor U1573 (N_1573,N_349,N_139);
or U1574 (N_1574,N_1360,N_872);
nor U1575 (N_1575,N_1458,In_2897);
or U1576 (N_1576,In_2548,In_157);
and U1577 (N_1577,N_1364,N_1316);
nand U1578 (N_1578,In_2089,N_290);
and U1579 (N_1579,In_1092,N_1229);
or U1580 (N_1580,In_1643,N_932);
nand U1581 (N_1581,N_593,N_207);
nor U1582 (N_1582,N_979,N_909);
or U1583 (N_1583,N_102,In_1321);
and U1584 (N_1584,In_735,N_1494);
nor U1585 (N_1585,N_1010,N_68);
or U1586 (N_1586,In_1308,In_1641);
or U1587 (N_1587,N_1357,In_2189);
nand U1588 (N_1588,N_1161,N_1441);
or U1589 (N_1589,In_1966,N_414);
nor U1590 (N_1590,N_1142,In_2924);
nand U1591 (N_1591,In_487,In_530);
nand U1592 (N_1592,N_282,N_494);
xnor U1593 (N_1593,N_378,N_695);
xor U1594 (N_1594,N_1260,N_762);
and U1595 (N_1595,N_1207,N_1369);
xor U1596 (N_1596,N_804,N_1405);
nand U1597 (N_1597,N_1202,N_799);
or U1598 (N_1598,In_2798,In_2298);
nand U1599 (N_1599,N_209,N_555);
and U1600 (N_1600,N_1340,N_993);
and U1601 (N_1601,In_1293,N_1040);
and U1602 (N_1602,N_919,In_2179);
nor U1603 (N_1603,In_344,In_567);
or U1604 (N_1604,N_1433,In_104);
or U1605 (N_1605,N_1098,N_1333);
nand U1606 (N_1606,N_1081,In_1316);
nand U1607 (N_1607,In_451,N_1404);
nand U1608 (N_1608,In_838,N_1124);
nor U1609 (N_1609,N_1491,N_817);
xnor U1610 (N_1610,N_683,N_1456);
or U1611 (N_1611,In_2499,In_1663);
xor U1612 (N_1612,N_649,N_394);
nor U1613 (N_1613,N_1284,In_2987);
nand U1614 (N_1614,In_1363,N_493);
nand U1615 (N_1615,N_1402,In_2858);
or U1616 (N_1616,In_1045,N_1111);
xnor U1617 (N_1617,In_2462,N_1166);
xnor U1618 (N_1618,N_1109,N_193);
nor U1619 (N_1619,N_732,In_1491);
xor U1620 (N_1620,In_1012,N_1274);
xor U1621 (N_1621,N_1122,N_1107);
nand U1622 (N_1622,In_2387,In_1997);
or U1623 (N_1623,In_737,N_1324);
or U1624 (N_1624,In_689,N_1390);
or U1625 (N_1625,N_1052,In_928);
nand U1626 (N_1626,In_1774,N_1228);
nand U1627 (N_1627,N_390,N_1454);
nand U1628 (N_1628,In_479,In_1090);
nand U1629 (N_1629,In_2439,In_1601);
nor U1630 (N_1630,N_667,In_2612);
nor U1631 (N_1631,In_977,N_195);
and U1632 (N_1632,In_95,In_650);
nand U1633 (N_1633,N_1410,N_1097);
xnor U1634 (N_1634,In_2276,N_1206);
nor U1635 (N_1635,N_1146,In_2033);
and U1636 (N_1636,In_140,In_2195);
nor U1637 (N_1637,In_498,N_1345);
nand U1638 (N_1638,N_1139,N_712);
and U1639 (N_1639,In_449,N_1317);
and U1640 (N_1640,N_1325,N_456);
nand U1641 (N_1641,In_2890,N_1395);
or U1642 (N_1642,N_950,N_1235);
nor U1643 (N_1643,In_164,N_1423);
or U1644 (N_1644,In_1876,N_726);
and U1645 (N_1645,N_441,In_1909);
xnor U1646 (N_1646,N_411,N_56);
and U1647 (N_1647,In_1273,In_1402);
and U1648 (N_1648,In_817,N_610);
and U1649 (N_1649,In_649,N_1328);
or U1650 (N_1650,N_350,In_955);
or U1651 (N_1651,N_741,N_1211);
nor U1652 (N_1652,In_295,In_109);
nor U1653 (N_1653,N_1227,In_2552);
and U1654 (N_1654,In_1094,N_1417);
nor U1655 (N_1655,In_1398,N_1442);
and U1656 (N_1656,N_1200,N_1300);
and U1657 (N_1657,In_1319,In_438);
or U1658 (N_1658,In_1808,In_1481);
nand U1659 (N_1659,In_1915,N_27);
or U1660 (N_1660,N_344,N_1126);
nor U1661 (N_1661,N_226,In_2107);
and U1662 (N_1662,In_63,In_1041);
nand U1663 (N_1663,In_42,In_501);
nand U1664 (N_1664,N_255,In_2870);
xor U1665 (N_1665,N_822,In_1167);
and U1666 (N_1666,In_1973,In_2835);
nand U1667 (N_1667,N_1371,N_834);
nand U1668 (N_1668,N_1077,In_2745);
nand U1669 (N_1669,In_666,In_984);
or U1670 (N_1670,N_176,N_308);
nor U1671 (N_1671,N_516,N_16);
nand U1672 (N_1672,N_1322,N_1239);
and U1673 (N_1673,N_757,In_1263);
xnor U1674 (N_1674,In_651,N_1269);
xor U1675 (N_1675,In_2964,In_753);
nand U1676 (N_1676,In_2051,In_2864);
or U1677 (N_1677,N_1290,In_1602);
nand U1678 (N_1678,In_1404,In_1175);
xor U1679 (N_1679,N_753,In_2881);
and U1680 (N_1680,N_1439,In_2925);
nand U1681 (N_1681,In_135,N_566);
nand U1682 (N_1682,N_1398,N_795);
or U1683 (N_1683,N_1263,In_697);
or U1684 (N_1684,In_2269,In_2990);
and U1685 (N_1685,In_2877,N_1412);
nor U1686 (N_1686,N_965,N_1044);
nor U1687 (N_1687,N_523,N_1155);
nor U1688 (N_1688,In_624,In_2041);
or U1689 (N_1689,N_697,In_2145);
nand U1690 (N_1690,In_2036,N_622);
nor U1691 (N_1691,N_1080,In_813);
nand U1692 (N_1692,N_981,In_2801);
xnor U1693 (N_1693,In_2812,N_1485);
and U1694 (N_1694,N_1311,N_1446);
or U1695 (N_1695,In_1463,In_223);
xor U1696 (N_1696,N_1259,N_360);
nand U1697 (N_1697,In_1452,In_2895);
and U1698 (N_1698,In_325,N_358);
or U1699 (N_1699,N_1363,N_1110);
nand U1700 (N_1700,N_1219,In_1642);
nand U1701 (N_1701,N_1270,In_2217);
or U1702 (N_1702,In_2543,N_584);
and U1703 (N_1703,N_1359,N_755);
nand U1704 (N_1704,N_1406,In_403);
or U1705 (N_1705,In_905,In_2416);
and U1706 (N_1706,N_510,N_995);
nand U1707 (N_1707,N_340,In_742);
nand U1708 (N_1708,In_1688,In_1058);
nand U1709 (N_1709,N_540,N_1285);
nand U1710 (N_1710,In_934,In_1710);
xor U1711 (N_1711,N_841,N_17);
xnor U1712 (N_1712,N_427,In_355);
and U1713 (N_1713,N_1231,N_1466);
or U1714 (N_1714,N_174,In_1037);
xor U1715 (N_1715,In_1132,N_1085);
nand U1716 (N_1716,N_816,In_54);
xor U1717 (N_1717,In_852,In_2331);
nand U1718 (N_1718,In_1532,In_2687);
or U1719 (N_1719,In_819,N_785);
or U1720 (N_1720,N_571,N_720);
nand U1721 (N_1721,N_1383,N_1303);
xor U1722 (N_1722,N_766,N_1370);
or U1723 (N_1723,In_2854,In_19);
or U1724 (N_1724,N_1156,In_502);
xnor U1725 (N_1725,N_1477,In_991);
and U1726 (N_1726,N_348,In_2723);
xor U1727 (N_1727,N_1355,N_127);
and U1728 (N_1728,N_811,In_596);
nor U1729 (N_1729,In_2163,N_103);
nor U1730 (N_1730,In_2585,N_659);
nand U1731 (N_1731,In_18,In_2473);
and U1732 (N_1732,In_739,In_2623);
xnor U1733 (N_1733,In_2992,N_1481);
and U1734 (N_1734,N_1474,In_1038);
and U1735 (N_1735,N_234,In_731);
nand U1736 (N_1736,N_1276,In_677);
xnor U1737 (N_1737,N_187,In_2535);
nor U1738 (N_1738,In_1150,N_949);
nor U1739 (N_1739,In_460,N_1264);
xor U1740 (N_1740,In_2676,In_2084);
xor U1741 (N_1741,N_1071,N_989);
nor U1742 (N_1742,In_535,In_754);
xor U1743 (N_1743,In_1931,In_2699);
or U1744 (N_1744,In_1420,In_191);
and U1745 (N_1745,In_1124,In_2894);
and U1746 (N_1746,In_2730,In_1621);
and U1747 (N_1747,N_914,In_2497);
xor U1748 (N_1748,N_1465,In_1935);
nand U1749 (N_1749,N_20,N_1391);
nor U1750 (N_1750,In_860,N_1148);
and U1751 (N_1751,N_363,In_2406);
nand U1752 (N_1752,In_80,N_968);
nor U1753 (N_1753,In_2375,In_1786);
nand U1754 (N_1754,In_1868,In_286);
nand U1755 (N_1755,In_1618,N_749);
nor U1756 (N_1756,N_1305,In_302);
xor U1757 (N_1757,N_779,In_184);
nand U1758 (N_1758,N_800,In_2648);
and U1759 (N_1759,N_717,N_714);
and U1760 (N_1760,In_2874,In_2755);
nand U1761 (N_1761,In_1595,In_1709);
xor U1762 (N_1762,N_807,N_1063);
or U1763 (N_1763,N_986,In_1139);
nor U1764 (N_1764,N_1354,In_493);
xnor U1765 (N_1765,N_1419,N_997);
or U1766 (N_1766,N_1018,In_798);
or U1767 (N_1767,N_959,N_765);
xnor U1768 (N_1768,N_1366,In_2611);
nor U1769 (N_1769,N_1365,In_665);
xnor U1770 (N_1770,N_370,N_1062);
and U1771 (N_1771,In_975,In_1375);
or U1772 (N_1772,In_2780,In_1797);
nor U1773 (N_1773,In_1914,N_461);
nand U1774 (N_1774,In_1989,N_1149);
and U1775 (N_1775,N_827,N_1230);
or U1776 (N_1776,N_1216,In_2718);
nor U1777 (N_1777,N_557,N_1171);
and U1778 (N_1778,In_1203,N_1197);
nor U1779 (N_1779,N_963,In_2821);
xor U1780 (N_1780,N_934,N_1184);
and U1781 (N_1781,In_2134,In_533);
or U1782 (N_1782,N_1241,N_1358);
xnor U1783 (N_1783,In_2328,N_1495);
and U1784 (N_1784,N_1102,N_1286);
xor U1785 (N_1785,N_1384,N_37);
nor U1786 (N_1786,N_759,N_941);
nor U1787 (N_1787,In_1235,N_705);
nor U1788 (N_1788,N_996,N_1249);
nand U1789 (N_1789,N_992,In_2609);
xnor U1790 (N_1790,N_767,In_428);
xor U1791 (N_1791,In_13,In_258);
and U1792 (N_1792,In_2054,In_2426);
or U1793 (N_1793,N_936,N_471);
xnor U1794 (N_1794,In_2799,N_700);
nor U1795 (N_1795,In_1153,In_2020);
and U1796 (N_1796,N_472,N_1220);
xnor U1797 (N_1797,N_90,N_1209);
and U1798 (N_1798,N_1030,N_1086);
xor U1799 (N_1799,In_401,N_1301);
xnor U1800 (N_1800,In_2766,N_1353);
nor U1801 (N_1801,N_1798,In_708);
xnor U1802 (N_1802,In_799,N_269);
nand U1803 (N_1803,N_1728,N_634);
and U1804 (N_1804,In_1617,N_1179);
xor U1805 (N_1805,In_667,In_1485);
and U1806 (N_1806,N_1686,In_1422);
nor U1807 (N_1807,N_1492,In_48);
and U1808 (N_1808,N_1332,N_706);
xnor U1809 (N_1809,In_829,N_1685);
nor U1810 (N_1810,N_1606,N_1725);
xnor U1811 (N_1811,N_1376,In_1073);
and U1812 (N_1812,In_2056,N_275);
or U1813 (N_1813,N_1361,N_1488);
nor U1814 (N_1814,N_514,In_2279);
xor U1815 (N_1815,In_2954,N_1515);
nor U1816 (N_1816,N_1413,N_1597);
nor U1817 (N_1817,N_1411,N_1582);
xnor U1818 (N_1818,In_2446,In_630);
or U1819 (N_1819,N_356,N_1645);
and U1820 (N_1820,In_2731,N_1699);
or U1821 (N_1821,N_1002,N_148);
or U1822 (N_1822,N_1695,N_1380);
and U1823 (N_1823,N_457,N_1266);
and U1824 (N_1824,N_1037,In_1077);
xnor U1825 (N_1825,N_1564,In_234);
xnor U1826 (N_1826,N_869,N_871);
nand U1827 (N_1827,In_3,In_1178);
nor U1828 (N_1828,N_1614,N_1426);
nand U1829 (N_1829,In_2685,N_679);
and U1830 (N_1830,N_1601,N_1298);
or U1831 (N_1831,In_1187,In_2616);
nor U1832 (N_1832,In_492,N_1604);
nor U1833 (N_1833,N_565,In_1610);
or U1834 (N_1834,N_1518,N_812);
xor U1835 (N_1835,In_2046,In_1500);
or U1836 (N_1836,N_1659,N_689);
and U1837 (N_1837,In_2130,N_396);
and U1838 (N_1838,N_1783,N_725);
nand U1839 (N_1839,N_451,N_1674);
and U1840 (N_1840,N_409,N_452);
or U1841 (N_1841,In_99,In_515);
and U1842 (N_1842,N_1224,N_1517);
nor U1843 (N_1843,In_39,N_910);
and U1844 (N_1844,N_1372,N_307);
and U1845 (N_1845,N_1032,In_2064);
nor U1846 (N_1846,N_1649,In_2092);
or U1847 (N_1847,In_2860,In_241);
nand U1848 (N_1848,N_1034,N_1708);
xor U1849 (N_1849,N_1525,N_586);
or U1850 (N_1850,In_2251,N_1640);
or U1851 (N_1851,N_728,In_90);
and U1852 (N_1852,In_2849,N_1566);
nand U1853 (N_1853,N_1613,N_1524);
and U1854 (N_1854,N_1455,N_1389);
nor U1855 (N_1855,In_954,N_45);
and U1856 (N_1856,N_1619,N_1723);
and U1857 (N_1857,In_976,N_569);
nand U1858 (N_1858,N_1403,N_1562);
xor U1859 (N_1859,N_581,In_2297);
nor U1860 (N_1860,In_85,N_1378);
nor U1861 (N_1861,N_1042,N_1559);
nand U1862 (N_1862,N_1460,N_328);
nor U1863 (N_1863,N_1510,N_1782);
nand U1864 (N_1864,N_460,In_2176);
nand U1865 (N_1865,In_536,N_1791);
and U1866 (N_1866,N_1746,In_1886);
nand U1867 (N_1867,N_1626,In_1683);
xnor U1868 (N_1868,N_1752,N_952);
nand U1869 (N_1869,N_1580,In_2285);
or U1870 (N_1870,In_1867,N_71);
or U1871 (N_1871,N_1749,N_1314);
nand U1872 (N_1872,In_2238,N_796);
nor U1873 (N_1873,In_2518,In_1399);
xor U1874 (N_1874,N_985,N_1735);
nand U1875 (N_1875,N_1012,N_1479);
xnor U1876 (N_1876,N_1701,N_1400);
nor U1877 (N_1877,N_1570,N_1486);
or U1878 (N_1878,N_1766,In_2923);
nor U1879 (N_1879,N_1336,N_942);
xnor U1880 (N_1880,N_1530,N_1440);
and U1881 (N_1881,In_1799,N_1634);
nor U1882 (N_1882,In_796,In_1093);
and U1883 (N_1883,In_952,In_848);
and U1884 (N_1884,N_1651,In_2732);
and U1885 (N_1885,N_180,N_1240);
xnor U1886 (N_1886,N_1622,In_2673);
nand U1887 (N_1887,N_1450,N_1128);
nand U1888 (N_1888,N_1534,N_1150);
or U1889 (N_1889,In_2657,N_1551);
nand U1890 (N_1890,In_1387,N_1427);
nand U1891 (N_1891,N_1234,In_2424);
xor U1892 (N_1892,N_1277,N_994);
xnor U1893 (N_1893,In_2043,In_2208);
xnor U1894 (N_1894,N_908,In_293);
nor U1895 (N_1895,In_805,In_918);
nand U1896 (N_1896,N_1679,N_867);
nand U1897 (N_1897,N_1135,In_2248);
nor U1898 (N_1898,N_1348,N_1793);
xnor U1899 (N_1899,N_145,In_1971);
or U1900 (N_1900,N_1624,N_1552);
xnor U1901 (N_1901,In_1335,N_1420);
nand U1902 (N_1902,N_1764,In_2617);
or U1903 (N_1903,N_609,In_1488);
nand U1904 (N_1904,In_2831,In_2768);
nand U1905 (N_1905,In_226,N_1496);
and U1906 (N_1906,N_873,N_341);
nor U1907 (N_1907,N_1675,In_382);
nor U1908 (N_1908,In_367,In_131);
and U1909 (N_1909,N_1668,In_2408);
nor U1910 (N_1910,In_1580,N_1019);
and U1911 (N_1911,N_1538,N_1713);
and U1912 (N_1912,N_883,N_1106);
or U1913 (N_1913,N_1099,In_1298);
and U1914 (N_1914,N_1256,N_342);
nor U1915 (N_1915,N_1662,In_1756);
or U1916 (N_1916,N_988,In_2558);
xnor U1917 (N_1917,N_1546,In_435);
or U1918 (N_1918,N_771,N_1346);
xor U1919 (N_1919,N_1508,N_1789);
nor U1920 (N_1920,N_962,N_1212);
xnor U1921 (N_1921,N_1254,N_1321);
nand U1922 (N_1922,N_1531,N_1609);
nand U1923 (N_1923,N_777,N_1215);
xnor U1924 (N_1924,In_196,N_990);
or U1925 (N_1925,N_1382,In_1029);
nand U1926 (N_1926,N_1368,N_1498);
nor U1927 (N_1927,In_45,In_119);
or U1928 (N_1928,In_2760,In_1669);
xnor U1929 (N_1929,N_1205,N_1637);
or U1930 (N_1930,In_2019,In_2175);
xor U1931 (N_1931,In_556,N_1133);
and U1932 (N_1932,N_1535,In_573);
or U1933 (N_1933,N_1593,N_1630);
nor U1934 (N_1934,In_20,N_1615);
nand U1935 (N_1935,N_713,N_1792);
nor U1936 (N_1936,N_1532,N_561);
nor U1937 (N_1937,N_750,N_62);
nor U1938 (N_1938,In_2905,N_1596);
xnor U1939 (N_1939,N_1157,In_1895);
xor U1940 (N_1940,In_1120,N_1678);
nand U1941 (N_1941,In_2663,In_1016);
and U1942 (N_1942,N_1765,In_2570);
or U1943 (N_1943,N_1093,N_1540);
or U1944 (N_1944,N_1475,N_907);
or U1945 (N_1945,N_1289,N_1120);
nand U1946 (N_1946,N_774,In_70);
nor U1947 (N_1947,N_1393,In_2308);
xor U1948 (N_1948,N_1550,N_11);
and U1949 (N_1949,In_2376,In_4);
xor U1950 (N_1950,N_1425,N_905);
xor U1951 (N_1951,N_1501,In_2540);
and U1952 (N_1952,N_911,In_924);
xnor U1953 (N_1953,N_745,N_843);
nand U1954 (N_1954,N_1648,N_1153);
xnor U1955 (N_1955,N_1610,In_2414);
and U1956 (N_1956,N_1586,In_2143);
nand U1957 (N_1957,N_19,N_1304);
nand U1958 (N_1958,N_1247,N_1611);
nor U1959 (N_1959,N_580,N_1483);
nand U1960 (N_1960,N_1035,N_761);
nand U1961 (N_1961,In_2364,In_574);
or U1962 (N_1962,In_2796,N_921);
xnor U1963 (N_1963,N_967,In_2692);
nor U1964 (N_1964,N_1711,N_1302);
nand U1965 (N_1965,N_1536,N_1435);
nor U1966 (N_1966,N_1167,N_1140);
or U1967 (N_1967,In_49,N_1539);
nor U1968 (N_1968,N_1653,In_1852);
nand U1969 (N_1969,N_652,N_980);
xor U1970 (N_1970,In_1006,N_1719);
or U1971 (N_1971,N_1594,In_1145);
xor U1972 (N_1972,In_2773,N_933);
and U1973 (N_1973,N_1650,In_730);
nand U1974 (N_1974,N_1409,N_1265);
and U1975 (N_1975,In_2696,In_1415);
xnor U1976 (N_1976,N_1262,N_1421);
xor U1977 (N_1977,N_917,N_1236);
xnor U1978 (N_1978,N_1521,In_2070);
and U1979 (N_1979,N_1696,N_650);
nor U1980 (N_1980,N_1469,In_318);
and U1981 (N_1981,N_1431,In_687);
xor U1982 (N_1982,In_967,N_1554);
xnor U1983 (N_1983,N_526,N_1452);
or U1984 (N_1984,N_1774,In_1883);
and U1985 (N_1985,N_436,N_1091);
xor U1986 (N_1986,N_1499,N_1733);
nor U1987 (N_1987,In_2913,N_1603);
or U1988 (N_1988,N_1557,N_1141);
or U1989 (N_1989,In_2547,In_2040);
and U1990 (N_1990,In_675,In_774);
nor U1991 (N_1991,N_1664,In_1903);
nor U1992 (N_1992,N_1401,In_2067);
or U1993 (N_1993,In_2472,N_1437);
nand U1994 (N_1994,In_1510,N_1587);
xor U1995 (N_1995,N_1279,In_1861);
xor U1996 (N_1996,N_964,In_1149);
nor U1997 (N_1997,N_1573,N_1436);
or U1998 (N_1998,In_2048,N_1068);
xnor U1999 (N_1999,N_1770,In_2156);
nand U2000 (N_2000,In_1624,In_404);
and U2001 (N_2001,In_1130,In_2501);
nor U2002 (N_2002,N_1616,N_1718);
xor U2003 (N_2003,N_1503,N_1267);
nand U2004 (N_2004,N_402,In_2169);
xor U2005 (N_2005,N_227,In_1865);
xnor U2006 (N_2006,N_137,In_1870);
or U2007 (N_2007,In_1494,N_1772);
nor U2008 (N_2008,N_1272,N_280);
xor U2009 (N_2009,In_477,In_2659);
or U2010 (N_2010,N_507,N_1797);
xnor U2011 (N_2011,In_380,N_1744);
or U2012 (N_2012,In_1818,N_1756);
and U2013 (N_2013,In_2464,N_663);
nor U2014 (N_2014,In_1556,N_1799);
and U2015 (N_2015,N_1154,N_1136);
nand U2016 (N_2016,In_1954,In_2315);
and U2017 (N_2017,N_1683,In_264);
or U2018 (N_2018,N_1487,N_662);
nand U2019 (N_2019,N_916,In_2907);
nand U2020 (N_2020,N_1592,In_1851);
nor U2021 (N_2021,N_522,N_1638);
nand U2022 (N_2022,N_1337,In_2995);
and U2023 (N_2023,In_2576,N_887);
xor U2024 (N_2024,In_1596,N_1244);
nor U2025 (N_2025,N_600,N_1553);
or U2026 (N_2026,In_444,N_1467);
nand U2027 (N_2027,In_1896,N_719);
or U2028 (N_2028,N_1598,In_1277);
xnor U2029 (N_2029,N_1631,N_641);
and U2030 (N_2030,In_2523,N_1738);
xor U2031 (N_2031,N_1089,N_513);
or U2032 (N_2032,N_797,In_356);
nand U2033 (N_2033,In_331,In_2166);
nor U2034 (N_2034,In_376,N_577);
nor U2035 (N_2035,N_1079,N_1250);
or U2036 (N_2036,In_2035,In_566);
nor U2037 (N_2037,N_1347,N_709);
or U2038 (N_2038,In_2743,N_1422);
xnor U2039 (N_2039,In_92,N_389);
nor U2040 (N_2040,N_1721,In_2108);
nor U2041 (N_2041,N_1061,N_1299);
and U2042 (N_2042,N_1323,N_408);
or U2043 (N_2043,N_1444,N_1137);
nor U2044 (N_2044,N_1692,N_1710);
xor U2045 (N_2045,N_1237,N_1057);
nor U2046 (N_2046,N_1743,N_1445);
or U2047 (N_2047,N_1676,N_1790);
or U2048 (N_2048,N_252,N_1769);
and U2049 (N_2049,In_2887,N_1581);
and U2050 (N_2050,N_1527,In_1686);
or U2051 (N_2051,N_1687,N_1753);
nor U2052 (N_2052,N_1387,N_730);
or U2053 (N_2053,N_1778,In_495);
or U2054 (N_2054,N_1636,N_656);
nor U2055 (N_2055,N_1751,N_1318);
nand U2056 (N_2056,N_1297,N_1548);
and U2057 (N_2057,In_1792,N_1654);
nand U2058 (N_2058,N_1602,N_1709);
nor U2059 (N_2059,N_1716,N_977);
nor U2060 (N_2060,N_1341,N_1771);
nor U2061 (N_2061,N_1261,N_987);
xor U2062 (N_2062,N_1434,In_644);
nor U2063 (N_2063,N_1667,In_614);
or U2064 (N_2064,N_1595,N_40);
or U2065 (N_2065,N_851,N_271);
xnor U2066 (N_2066,N_915,In_1103);
nor U2067 (N_2067,N_858,N_1541);
or U2068 (N_2068,In_586,N_1065);
and U2069 (N_2069,In_2103,N_1724);
xor U2070 (N_2070,N_1350,N_23);
nor U2071 (N_2071,In_117,N_710);
nor U2072 (N_2072,In_72,N_1522);
xor U2073 (N_2073,N_1173,In_698);
xnor U2074 (N_2074,N_250,In_1259);
and U2075 (N_2075,N_1584,N_642);
nor U2076 (N_2076,In_1827,In_22);
nor U2077 (N_2077,N_1690,N_688);
or U2078 (N_2078,In_209,N_888);
nand U2079 (N_2079,N_1480,N_1607);
xnor U2080 (N_2080,N_1232,N_1663);
nor U2081 (N_2081,N_1747,In_613);
or U2082 (N_2082,In_791,N_862);
nand U2083 (N_2083,N_1050,In_1832);
and U2084 (N_2084,N_1697,N_1127);
and U2085 (N_2085,N_425,N_1571);
xor U2086 (N_2086,In_1152,N_570);
nor U2087 (N_2087,In_1417,N_9);
or U2088 (N_2088,N_1576,N_291);
xor U2089 (N_2089,N_969,N_1191);
nor U2090 (N_2090,In_1508,N_756);
xor U2091 (N_2091,N_1208,N_1385);
nor U2092 (N_2092,N_1773,N_677);
nor U2093 (N_2093,In_2781,In_2855);
or U2094 (N_2094,N_1054,N_1428);
and U2095 (N_2095,In_2567,N_808);
and U2096 (N_2096,N_784,In_699);
xnor U2097 (N_2097,N_1386,N_61);
and U2098 (N_2098,In_2291,N_1315);
or U2099 (N_2099,N_1038,N_1443);
nor U2100 (N_2100,In_2106,N_1556);
or U2101 (N_2101,N_1856,N_1027);
and U2102 (N_2102,N_1933,N_119);
nor U2103 (N_2103,N_2084,N_1867);
and U2104 (N_2104,N_2095,In_1615);
and U2105 (N_2105,N_1021,N_2003);
and U2106 (N_2106,N_1731,In_2206);
or U2107 (N_2107,N_925,N_1957);
xor U2108 (N_2108,N_265,In_1755);
nor U2109 (N_2109,In_2294,N_1968);
and U2110 (N_2110,N_1352,In_2682);
and U2111 (N_2111,N_2005,N_1449);
nor U2112 (N_2112,N_1414,N_1971);
or U2113 (N_2113,N_1954,In_2031);
nor U2114 (N_2114,N_1213,N_1320);
or U2115 (N_2115,N_1919,In_1229);
xor U2116 (N_2116,In_1440,N_1451);
nor U2117 (N_2117,N_805,In_219);
nor U2118 (N_2118,N_1853,N_1991);
nor U2119 (N_2119,N_2022,N_1914);
nor U2120 (N_2120,N_1418,N_1514);
or U2121 (N_2121,N_1819,N_1563);
xnor U2122 (N_2122,N_1666,N_1011);
nor U2123 (N_2123,In_2645,In_2764);
xnor U2124 (N_2124,In_1163,In_988);
nor U2125 (N_2125,In_622,N_1574);
nand U2126 (N_2126,N_1921,N_1430);
and U2127 (N_2127,In_2132,N_704);
or U2128 (N_2128,N_1688,N_1447);
nor U2129 (N_2129,N_1704,N_343);
or U2130 (N_2130,N_1408,N_1226);
and U2131 (N_2131,N_1815,N_2060);
xor U2132 (N_2132,In_175,N_417);
nor U2133 (N_2133,N_1567,N_155);
nand U2134 (N_2134,In_1390,In_2302);
or U2135 (N_2135,N_1820,N_1113);
xnor U2136 (N_2136,N_1942,N_830);
nor U2137 (N_2137,N_1838,N_1292);
xor U2138 (N_2138,In_2351,N_353);
and U2139 (N_2139,N_1907,N_1777);
or U2140 (N_2140,N_1750,In_2345);
xnor U2141 (N_2141,N_1367,N_583);
nor U2142 (N_2142,N_1837,N_1281);
or U2143 (N_2143,N_1343,N_1204);
nand U2144 (N_2144,N_632,In_1486);
nor U2145 (N_2145,N_1201,N_2048);
or U2146 (N_2146,N_2039,N_2031);
nor U2147 (N_2147,N_2019,In_914);
nand U2148 (N_2148,N_1888,N_2089);
nand U2149 (N_2149,N_1862,N_2059);
nand U2150 (N_2150,In_565,N_1880);
xor U2151 (N_2151,In_2191,N_1100);
or U2152 (N_2152,N_1644,N_1817);
xor U2153 (N_2153,N_2017,N_1970);
xnor U2154 (N_2154,N_2061,In_1386);
and U2155 (N_2155,In_2393,N_1472);
nand U2156 (N_2156,N_1739,N_2002);
nor U2157 (N_2157,N_2036,N_1748);
nand U2158 (N_2158,N_1927,N_1974);
and U2159 (N_2159,In_2226,N_1076);
and U2160 (N_2160,N_1572,N_844);
xor U2161 (N_2161,N_1657,In_486);
and U2162 (N_2162,N_1056,N_2015);
nand U2163 (N_2163,N_1956,N_407);
nor U2164 (N_2164,N_1775,N_1892);
or U2165 (N_2165,N_1840,N_1834);
or U2166 (N_2166,N_2075,N_1767);
nand U2167 (N_2167,In_2876,N_1160);
and U2168 (N_2168,N_598,N_1841);
and U2169 (N_2169,In_389,N_1884);
or U2170 (N_2170,N_1646,N_1017);
xor U2171 (N_2171,N_1349,In_317);
nand U2172 (N_2172,N_2018,N_1964);
xor U2173 (N_2173,In_274,N_232);
and U2174 (N_2174,N_1291,N_668);
nand U2175 (N_2175,N_1362,N_1677);
or U2176 (N_2176,N_1890,N_1661);
nand U2177 (N_2177,In_2551,N_1658);
or U2178 (N_2178,N_1903,N_1132);
or U2179 (N_2179,In_557,N_1578);
nand U2180 (N_2180,In_2962,In_2797);
or U2181 (N_2181,N_1873,In_2596);
and U2182 (N_2182,N_1647,N_2069);
or U2183 (N_2183,N_1901,In_2578);
xnor U2184 (N_2184,N_1036,N_1910);
nor U2185 (N_2185,N_1920,In_1112);
nand U2186 (N_2186,N_1504,In_1400);
nand U2187 (N_2187,N_2014,In_1538);
nor U2188 (N_2188,N_1811,N_1294);
nand U2189 (N_2189,In_299,N_1730);
nor U2190 (N_2190,N_1736,N_393);
nand U2191 (N_2191,N_2070,In_1281);
and U2192 (N_2192,N_1705,N_1740);
and U2193 (N_2193,N_1712,N_1072);
or U2194 (N_2194,N_1992,N_1810);
nor U2195 (N_2195,N_1781,In_2904);
nand U2196 (N_2196,N_2024,N_1951);
xnor U2197 (N_2197,N_2090,In_2151);
xor U2198 (N_2198,N_619,N_739);
and U2199 (N_2199,N_1839,In_256);
xnor U2200 (N_2200,N_462,N_1976);
or U2201 (N_2201,N_1660,N_2038);
or U2202 (N_2202,N_2093,N_388);
and U2203 (N_2203,N_794,N_1876);
xor U2204 (N_2204,N_1929,N_81);
nand U2205 (N_2205,N_1776,In_480);
nor U2206 (N_2206,N_1327,N_2088);
and U2207 (N_2207,N_1008,N_971);
or U2208 (N_2208,In_570,N_1275);
nand U2209 (N_2209,N_1643,In_941);
xnor U2210 (N_2210,In_2411,N_15);
and U2211 (N_2211,N_1043,N_1282);
xnor U2212 (N_2212,N_1516,N_1482);
or U2213 (N_2213,N_664,N_2065);
nand U2214 (N_2214,N_2092,N_736);
xor U2215 (N_2215,N_1732,In_2901);
and U2216 (N_2216,N_1828,N_935);
or U2217 (N_2217,N_1543,In_59);
or U2218 (N_2218,N_1243,N_1801);
nor U2219 (N_2219,In_2484,N_1513);
or U2220 (N_2220,In_935,In_1983);
nand U2221 (N_2221,N_1906,In_2721);
and U2222 (N_2222,N_1618,N_1943);
and U2223 (N_2223,N_1625,N_1983);
xor U2224 (N_2224,N_1338,N_1788);
or U2225 (N_2225,N_1979,In_2922);
and U2226 (N_2226,In_1410,In_352);
nand U2227 (N_2227,N_2098,N_419);
xnor U2228 (N_2228,N_1569,In_360);
xnor U2229 (N_2229,N_1394,N_1855);
or U2230 (N_2230,N_1984,In_2989);
nor U2231 (N_2231,N_1680,In_2785);
nand U2232 (N_2232,In_1442,N_2077);
or U2233 (N_2233,N_1116,In_2948);
nand U2234 (N_2234,N_1377,N_1872);
and U2235 (N_2235,N_495,N_1096);
nor U2236 (N_2236,N_1848,N_2076);
nor U2237 (N_2237,N_1588,N_1397);
nand U2238 (N_2238,In_1330,N_1900);
nand U2239 (N_2239,N_2023,N_2080);
or U2240 (N_2240,In_1598,N_1831);
nor U2241 (N_2241,In_2032,N_1507);
or U2242 (N_2242,N_722,In_604);
xnor U2243 (N_2243,In_2618,N_1560);
or U2244 (N_2244,In_1919,N_1542);
xor U2245 (N_2245,N_359,N_1998);
and U2246 (N_2246,N_1879,N_1847);
nand U2247 (N_2247,N_1432,N_2055);
or U2248 (N_2248,N_1805,N_912);
or U2249 (N_2249,N_1824,N_2074);
nor U2250 (N_2250,N_1883,N_1905);
nand U2251 (N_2251,N_1982,N_104);
and U2252 (N_2252,In_366,In_2148);
nor U2253 (N_2253,N_1203,N_1722);
xor U2254 (N_2254,N_1633,N_1939);
or U2255 (N_2255,N_1671,In_636);
and U2256 (N_2256,N_1986,N_2025);
xor U2257 (N_2257,N_1825,N_1693);
nor U2258 (N_2258,N_1490,N_1415);
nor U2259 (N_2259,N_926,N_345);
nand U2260 (N_2260,N_929,N_537);
and U2261 (N_2261,N_128,N_1821);
nor U2262 (N_2262,N_1568,N_1198);
and U2263 (N_2263,N_1934,In_1078);
or U2264 (N_2264,In_1218,N_2066);
or U2265 (N_2265,N_1923,N_1273);
xor U2266 (N_2266,N_1945,N_1960);
nand U2267 (N_2267,In_2240,N_2099);
and U2268 (N_2268,In_2885,N_854);
nor U2269 (N_2269,N_2011,N_1865);
and U2270 (N_2270,N_199,In_1592);
nor U2271 (N_2271,N_1319,N_924);
nand U2272 (N_2272,In_348,N_1941);
or U2273 (N_2273,N_1375,N_1575);
xnor U2274 (N_2274,N_1787,N_631);
and U2275 (N_2275,N_1955,N_1895);
nand U2276 (N_2276,In_1512,In_252);
and U2277 (N_2277,N_1009,N_1656);
nand U2278 (N_2278,In_681,N_1698);
nor U2279 (N_2279,In_925,N_1547);
nand U2280 (N_2280,N_1223,In_1291);
or U2281 (N_2281,N_1720,N_1612);
xnor U2282 (N_2282,In_1214,N_1670);
or U2283 (N_2283,In_507,N_384);
xor U2284 (N_2284,N_1278,N_896);
and U2285 (N_2285,N_1785,N_2013);
and U2286 (N_2286,In_2938,N_1882);
and U2287 (N_2287,N_1628,N_326);
xor U2288 (N_2288,N_1288,N_1928);
nand U2289 (N_2289,N_1930,N_2037);
and U2290 (N_2290,In_963,In_1691);
or U2291 (N_2291,N_1993,N_1940);
nand U2292 (N_2292,In_2381,In_2476);
nor U2293 (N_2293,N_2047,In_2906);
or U2294 (N_2294,N_1707,N_2063);
xnor U2295 (N_2295,N_1478,N_1963);
and U2296 (N_2296,N_1737,N_1870);
nand U2297 (N_2297,N_1996,In_2463);
xnor U2298 (N_2298,N_1715,N_355);
xor U2299 (N_2299,N_1509,In_2722);
and U2300 (N_2300,N_1092,N_1965);
and U2301 (N_2301,N_1589,N_2028);
and U2302 (N_2302,N_1990,N_1058);
nand U2303 (N_2303,N_1706,N_1462);
nand U2304 (N_2304,N_1512,N_1932);
and U2305 (N_2305,N_2027,N_1049);
and U2306 (N_2306,N_1691,N_1904);
nand U2307 (N_2307,N_1185,N_154);
and U2308 (N_2308,N_1463,N_1717);
nor U2309 (N_2309,N_1897,N_1926);
or U2310 (N_2310,N_1829,N_922);
or U2311 (N_2311,N_183,In_1544);
or U2312 (N_2312,N_1026,N_133);
xnor U2313 (N_2313,N_1918,N_434);
nand U2314 (N_2314,N_781,N_1700);
xnor U2315 (N_2315,N_1617,N_1757);
nand U2316 (N_2316,In_2871,N_1159);
or U2317 (N_2317,N_2052,N_938);
nor U2318 (N_2318,N_1754,N_1898);
nor U2319 (N_2319,N_1632,N_1125);
nor U2320 (N_2320,In_1114,N_1858);
xor U2321 (N_2321,N_1891,N_1889);
xnor U2322 (N_2322,N_1331,N_1095);
or U2323 (N_2323,N_2030,N_1953);
nand U2324 (N_2324,In_756,N_1832);
or U2325 (N_2325,In_2062,In_1718);
xor U2326 (N_2326,N_1836,N_543);
nor U2327 (N_2327,N_1961,N_1812);
nand U2328 (N_2328,N_1344,N_222);
or U2329 (N_2329,In_1347,N_1850);
nand U2330 (N_2330,N_661,N_1064);
xnor U2331 (N_2331,N_1293,N_1800);
and U2332 (N_2332,N_1727,In_1447);
and U2333 (N_2333,In_1798,N_1307);
or U2334 (N_2334,N_1528,N_1635);
nand U2335 (N_2335,N_1995,In_2263);
or U2336 (N_2336,N_1313,In_957);
and U2337 (N_2337,In_1807,N_1608);
or U2338 (N_2338,In_2998,N_1952);
xor U2339 (N_2339,N_838,N_2091);
xnor U2340 (N_2340,N_1672,N_1681);
xnor U2341 (N_2341,In_1630,N_1877);
or U2342 (N_2342,N_1689,In_2066);
nor U2343 (N_2343,N_1816,N_1988);
nor U2344 (N_2344,N_2096,In_1287);
nand U2345 (N_2345,In_511,N_1973);
xnor U2346 (N_2346,N_2064,N_2068);
xor U2347 (N_2347,N_1729,N_1225);
xor U2348 (N_2348,In_2526,N_1669);
nor U2349 (N_2349,In_1930,N_1673);
xor U2350 (N_2350,N_2009,N_1583);
or U2351 (N_2351,N_1599,N_1909);
xnor U2352 (N_2352,N_865,N_1641);
or U2353 (N_2353,N_885,In_625);
and U2354 (N_2354,N_1502,In_2275);
xor U2355 (N_2355,N_1585,N_1823);
nor U2356 (N_2356,N_1843,In_472);
nor U2357 (N_2357,In_58,N_599);
xor U2358 (N_2358,In_2879,N_1949);
nor U2359 (N_2359,N_1947,In_1469);
nor U2360 (N_2360,N_1857,N_1875);
nor U2361 (N_2361,N_1255,N_1874);
xnor U2362 (N_2362,N_1182,In_959);
nor U2363 (N_2363,N_1561,N_1005);
nand U2364 (N_2364,N_2073,In_2399);
xor U2365 (N_2365,N_1795,N_1306);
or U2366 (N_2366,N_2029,N_1814);
xor U2367 (N_2367,N_1925,N_1271);
and U2368 (N_2368,N_538,N_2045);
nand U2369 (N_2369,In_1198,In_2286);
xnor U2370 (N_2370,N_1655,N_1780);
xnor U2371 (N_2371,N_1859,In_1634);
nor U2372 (N_2372,N_716,N_692);
or U2373 (N_2373,In_1312,N_2083);
nand U2374 (N_2374,N_1989,N_2033);
or U2375 (N_2375,In_216,N_202);
xnor U2376 (N_2376,N_1158,N_1549);
nor U2377 (N_2377,N_1627,In_275);
or U2378 (N_2378,N_991,N_846);
nand U2379 (N_2379,N_1533,In_2763);
or U2380 (N_2380,N_1476,N_1966);
nand U2381 (N_2381,N_945,N_1962);
nor U2382 (N_2382,In_2058,N_1335);
nor U2383 (N_2383,N_1869,N_463);
and U2384 (N_2384,N_1257,N_1822);
or U2385 (N_2385,In_1788,In_743);
or U2386 (N_2386,N_1652,N_392);
xnor U2387 (N_2387,N_1218,N_1565);
and U2388 (N_2388,N_1734,In_499);
and U2389 (N_2389,In_2960,N_1894);
xnor U2390 (N_2390,N_1296,N_1911);
or U2391 (N_2391,N_1827,In_992);
nor U2392 (N_2392,N_1374,N_281);
nand U2393 (N_2393,N_542,N_1980);
xor U2394 (N_2394,In_2253,N_1899);
nand U2395 (N_2395,N_1537,N_1642);
nor U2396 (N_2396,N_886,N_1022);
xnor U2397 (N_2397,In_338,In_2465);
xnor U2398 (N_2398,N_2006,N_1591);
xnor U2399 (N_2399,N_1913,N_482);
xnor U2400 (N_2400,N_2233,N_2150);
nand U2401 (N_2401,In_2500,N_2086);
and U2402 (N_2402,N_1326,N_2187);
or U2403 (N_2403,N_2276,N_1763);
xnor U2404 (N_2404,N_2308,N_675);
xor U2405 (N_2405,N_2269,N_2324);
or U2406 (N_2406,N_1334,N_1826);
nor U2407 (N_2407,N_2032,N_2266);
nand U2408 (N_2408,N_2000,In_795);
and U2409 (N_2409,N_2216,N_2280);
xor U2410 (N_2410,N_2338,N_2120);
nand U2411 (N_2411,N_2369,N_2116);
or U2412 (N_2412,N_1605,N_1759);
xor U2413 (N_2413,N_2328,N_1500);
xor U2414 (N_2414,In_749,N_2012);
nand U2415 (N_2415,N_2316,N_2288);
or U2416 (N_2416,In_2569,In_559);
xnor U2417 (N_2417,N_1806,N_1977);
or U2418 (N_2418,N_1999,N_2218);
xnor U2419 (N_2419,N_2361,N_2339);
and U2420 (N_2420,N_1885,N_2345);
or U2421 (N_2421,N_1755,N_2365);
or U2422 (N_2422,N_1356,N_2142);
nand U2423 (N_2423,N_2278,N_1959);
nand U2424 (N_2424,N_458,N_1760);
xor U2425 (N_2425,N_2176,N_2222);
and U2426 (N_2426,N_1222,N_2366);
and U2427 (N_2427,N_1851,N_2165);
and U2428 (N_2428,N_2202,In_1157);
or U2429 (N_2429,N_2136,N_1579);
and U2430 (N_2430,N_2109,N_2110);
xnor U2431 (N_2431,N_2138,N_2199);
xor U2432 (N_2432,N_1373,N_2362);
xnor U2433 (N_2433,N_603,N_2287);
nand U2434 (N_2434,N_2240,N_2160);
nand U2435 (N_2435,N_2169,N_2331);
nor U2436 (N_2436,N_2113,N_2167);
nor U2437 (N_2437,N_2179,N_2340);
nor U2438 (N_2438,N_2396,N_1908);
nand U2439 (N_2439,N_1329,N_2154);
or U2440 (N_2440,N_2200,N_2292);
or U2441 (N_2441,N_1342,N_2388);
nor U2442 (N_2442,In_680,N_1682);
or U2443 (N_2443,N_2351,In_2866);
or U2444 (N_2444,N_2209,N_1871);
nor U2445 (N_2445,N_2051,N_184);
nor U2446 (N_2446,N_2035,In_1372);
xor U2447 (N_2447,In_993,N_2156);
nand U2448 (N_2448,In_2991,N_1808);
nor U2449 (N_2449,N_2188,In_1899);
and U2450 (N_2450,N_2105,In_2227);
xnor U2451 (N_2451,N_2231,N_14);
and U2452 (N_2452,N_2008,N_2082);
or U2453 (N_2453,In_246,N_2359);
and U2454 (N_2454,N_2270,N_2397);
and U2455 (N_2455,N_2230,N_1804);
xnor U2456 (N_2456,N_294,N_2117);
nand U2457 (N_2457,N_2321,N_2325);
nor U2458 (N_2458,N_1852,N_1505);
nor U2459 (N_2459,N_2279,N_2215);
nand U2460 (N_2460,N_1802,N_2146);
nor U2461 (N_2461,N_1818,N_2050);
nor U2462 (N_2462,N_2391,N_2301);
nand U2463 (N_2463,N_2399,N_2390);
xnor U2464 (N_2464,N_2078,N_2285);
xor U2465 (N_2465,N_2244,N_2021);
nor U2466 (N_2466,N_1114,N_2384);
nor U2467 (N_2467,In_2620,N_1887);
xnor U2468 (N_2468,N_1944,N_2041);
and U2469 (N_2469,N_1555,N_1969);
nor U2470 (N_2470,N_2198,N_2344);
and U2471 (N_2471,N_2326,N_738);
xor U2472 (N_2472,N_1846,N_2224);
xor U2473 (N_2473,N_2260,In_1267);
nand U2474 (N_2474,N_2327,N_2049);
or U2475 (N_2475,N_2272,N_1762);
nor U2476 (N_2476,N_1978,N_2255);
nand U2477 (N_2477,N_2001,N_2275);
nand U2478 (N_2478,N_2346,N_1526);
nor U2479 (N_2479,N_2081,N_2332);
xor U2480 (N_2480,N_1084,N_1714);
nand U2481 (N_2481,N_2371,N_2124);
or U2482 (N_2482,In_2087,N_1784);
nor U2483 (N_2483,N_385,N_1544);
nor U2484 (N_2484,N_900,N_1511);
or U2485 (N_2485,N_2297,In_2045);
nand U2486 (N_2486,N_2236,N_2294);
or U2487 (N_2487,N_2262,N_881);
or U2488 (N_2488,N_1916,N_1854);
xnor U2489 (N_2489,N_1520,N_1987);
nor U2490 (N_2490,N_2042,N_2172);
and U2491 (N_2491,N_1258,In_1100);
nor U2492 (N_2492,In_537,In_691);
nor U2493 (N_2493,N_1742,N_1972);
nor U2494 (N_2494,N_2170,N_2389);
xor U2495 (N_2495,N_1833,In_123);
xnor U2496 (N_2496,N_2249,N_2356);
nand U2497 (N_2497,In_2972,N_1221);
nand U2498 (N_2498,N_2135,N_2128);
or U2499 (N_2499,N_2134,N_1975);
nand U2500 (N_2500,In_37,N_2313);
nor U2501 (N_2501,N_2237,N_591);
xor U2502 (N_2502,In_826,N_2058);
and U2503 (N_2503,N_2234,N_1842);
xnor U2504 (N_2504,N_2214,In_1247);
nand U2505 (N_2505,N_2319,N_1621);
nor U2506 (N_2506,N_2072,N_2291);
or U2507 (N_2507,N_2374,In_2360);
xnor U2508 (N_2508,N_1924,N_1726);
nand U2509 (N_2509,N_2296,N_1506);
xnor U2510 (N_2510,N_2158,N_1935);
and U2511 (N_2511,N_2302,N_2191);
or U2512 (N_2512,N_2251,N_775);
or U2513 (N_2513,N_1694,N_2228);
or U2514 (N_2514,In_1677,N_1830);
xor U2515 (N_2515,N_2310,In_2382);
nor U2516 (N_2516,N_2175,N_2114);
nand U2517 (N_2517,N_2283,N_2194);
nor U2518 (N_2518,N_2201,N_2119);
xnor U2519 (N_2519,N_2273,N_1242);
nor U2520 (N_2520,In_2267,N_2108);
or U2521 (N_2521,N_1878,In_2455);
nand U2522 (N_2522,In_1777,In_2656);
and U2523 (N_2523,N_2349,N_2281);
nor U2524 (N_2524,N_2323,In_1033);
or U2525 (N_2525,N_2358,N_2149);
xor U2526 (N_2526,N_2239,N_2254);
or U2527 (N_2527,N_2380,N_2147);
nand U2528 (N_2528,N_2309,N_2372);
xor U2529 (N_2529,N_2122,N_1866);
nand U2530 (N_2530,N_1119,N_2219);
nand U2531 (N_2531,N_2243,N_1233);
xnor U2532 (N_2532,In_2469,N_1558);
nand U2533 (N_2533,N_2087,N_2261);
or U2534 (N_2534,N_2227,N_2333);
xor U2535 (N_2535,N_1620,N_26);
or U2536 (N_2536,N_2101,N_1946);
or U2537 (N_2537,N_1407,N_2067);
and U2538 (N_2538,N_2386,N_2159);
and U2539 (N_2539,N_2043,N_1786);
nand U2540 (N_2540,N_2343,N_1845);
and U2541 (N_2541,N_2181,N_1950);
or U2542 (N_2542,N_1702,N_2127);
and U2543 (N_2543,N_2232,N_2054);
nor U2544 (N_2544,N_1629,In_2246);
nor U2545 (N_2545,N_1917,N_2094);
xnor U2546 (N_2546,In_1244,N_2189);
nor U2547 (N_2547,N_2171,N_2263);
nand U2548 (N_2548,N_1994,In_1779);
and U2549 (N_2549,N_548,N_1238);
nand U2550 (N_2550,N_2378,N_2111);
nand U2551 (N_2551,N_2342,In_549);
xnor U2552 (N_2552,N_2207,N_2151);
or U2553 (N_2553,N_743,N_2129);
nand U2554 (N_2554,N_1807,N_296);
xnor U2555 (N_2555,N_2197,In_2517);
xnor U2556 (N_2556,N_1016,N_1844);
xnor U2557 (N_2557,N_2341,N_2007);
xnor U2558 (N_2558,N_2387,N_1330);
or U2559 (N_2559,N_2206,N_2367);
and U2560 (N_2560,N_2180,In_1559);
nand U2561 (N_2561,N_1931,N_2284);
or U2562 (N_2562,N_2026,N_1388);
nand U2563 (N_2563,N_1912,N_612);
nor U2564 (N_2564,N_2317,N_263);
nor U2565 (N_2565,N_2190,N_2290);
nand U2566 (N_2566,N_1623,N_2370);
nor U2567 (N_2567,In_139,N_1886);
xnor U2568 (N_2568,N_1529,N_2379);
or U2569 (N_2569,N_1577,N_2140);
nor U2570 (N_2570,N_1863,In_2006);
or U2571 (N_2571,N_2353,N_2226);
and U2572 (N_2572,In_1550,N_2155);
and U2573 (N_2573,N_1813,N_2335);
nand U2574 (N_2574,In_2486,N_1981);
nor U2575 (N_2575,N_2139,N_2256);
or U2576 (N_2576,N_2046,N_2364);
nor U2577 (N_2577,N_2271,N_2274);
or U2578 (N_2578,N_1493,N_2010);
nand U2579 (N_2579,N_2252,N_2257);
nand U2580 (N_2580,In_34,N_1985);
xnor U2581 (N_2581,N_2217,N_2100);
nor U2582 (N_2582,N_1893,N_835);
or U2583 (N_2583,N_123,N_2166);
nor U2584 (N_2584,N_2016,N_1741);
nand U2585 (N_2585,N_2314,In_1539);
or U2586 (N_2586,N_2195,N_2352);
xor U2587 (N_2587,N_1915,N_2210);
nand U2588 (N_2588,N_1399,N_2130);
and U2589 (N_2589,N_1902,N_1429);
nor U2590 (N_2590,N_2293,N_1471);
and U2591 (N_2591,N_2211,N_2363);
and U2592 (N_2592,N_2242,N_2137);
nor U2593 (N_2593,N_2268,N_2203);
and U2594 (N_2594,N_1809,N_2298);
and U2595 (N_2595,N_1590,N_1025);
and U2596 (N_2596,N_369,N_2148);
and U2597 (N_2597,N_2177,N_2107);
xor U2598 (N_2598,N_2220,N_2162);
xnor U2599 (N_2599,N_1031,N_2192);
nand U2600 (N_2600,N_2183,N_2004);
nand U2601 (N_2601,N_2395,N_2221);
and U2602 (N_2602,N_2398,N_2357);
nor U2603 (N_2603,In_2309,N_1768);
or U2604 (N_2604,N_2044,N_1896);
nand U2605 (N_2605,In_2470,N_1381);
or U2606 (N_2606,N_1794,N_2322);
or U2607 (N_2607,In_1523,N_2097);
nor U2608 (N_2608,N_1881,N_2174);
xnor U2609 (N_2609,N_2394,N_1835);
nand U2610 (N_2610,N_2212,N_2131);
xnor U2611 (N_2611,N_2377,In_361);
nand U2612 (N_2612,N_2141,N_2196);
nor U2613 (N_2613,N_898,N_1523);
nand U2614 (N_2614,N_1251,N_2373);
or U2615 (N_2615,N_2295,N_2168);
and U2616 (N_2616,N_1684,N_2121);
xnor U2617 (N_2617,N_2071,N_746);
nand U2618 (N_2618,N_2330,N_1779);
nand U2619 (N_2619,N_1997,N_2305);
and U2620 (N_2620,N_833,In_785);
xor U2621 (N_2621,In_1278,In_218);
nand U2622 (N_2622,N_957,N_2143);
nor U2623 (N_2623,N_1922,N_2182);
nand U2624 (N_2624,N_2277,N_2193);
xnor U2625 (N_2625,N_2383,In_437);
and U2626 (N_2626,N_1803,N_2112);
nand U2627 (N_2627,N_2115,N_2118);
xor U2628 (N_2628,N_1253,N_2354);
nor U2629 (N_2629,N_2153,N_1416);
xnor U2630 (N_2630,N_1936,N_2347);
nor U2631 (N_2631,In_1357,N_2248);
or U2632 (N_2632,N_2225,N_2145);
nor U2633 (N_2633,N_923,In_1772);
xnor U2634 (N_2634,N_2247,N_2161);
nand U2635 (N_2635,In_900,N_2238);
xor U2636 (N_2636,N_946,N_2385);
xnor U2637 (N_2637,N_1310,N_1004);
nor U2638 (N_2638,N_2157,N_440);
nand U2639 (N_2639,N_2208,N_2304);
nand U2640 (N_2640,N_1849,In_1043);
nand U2641 (N_2641,N_2376,N_1761);
nand U2642 (N_2642,N_1948,In_2026);
or U2643 (N_2643,In_453,N_2103);
nor U2644 (N_2644,N_1639,N_2334);
nand U2645 (N_2645,N_2375,N_1703);
or U2646 (N_2646,N_2125,N_2282);
nor U2647 (N_2647,N_2185,In_1904);
or U2648 (N_2648,N_2265,In_983);
nor U2649 (N_2649,N_2126,N_1860);
nor U2650 (N_2650,N_2329,N_1861);
or U2651 (N_2651,N_930,N_2348);
or U2652 (N_2652,N_2133,N_2062);
nor U2653 (N_2653,In_872,In_1894);
xnor U2654 (N_2654,N_2355,N_1868);
and U2655 (N_2655,N_2079,N_2104);
or U2656 (N_2656,N_2350,N_927);
nor U2657 (N_2657,N_2235,N_2020);
xor U2658 (N_2658,N_2102,N_2264);
nor U2659 (N_2659,N_1796,N_1214);
xnor U2660 (N_2660,N_2312,N_1519);
and U2661 (N_2661,N_2250,N_1252);
nor U2662 (N_2662,N_2163,N_2320);
and U2663 (N_2663,N_2306,N_2213);
and U2664 (N_2664,N_1473,N_2106);
or U2665 (N_2665,N_285,N_2034);
or U2666 (N_2666,N_2299,N_2382);
nor U2667 (N_2667,N_1758,N_2360);
or U2668 (N_2668,N_2368,N_2286);
or U2669 (N_2669,N_1151,N_2303);
xnor U2670 (N_2670,N_1039,N_2392);
nor U2671 (N_2671,N_1967,N_2259);
xor U2672 (N_2672,In_2791,N_2123);
xnor U2673 (N_2673,N_2040,N_2315);
or U2674 (N_2674,N_657,In_2073);
or U2675 (N_2675,N_2241,N_2267);
nand U2676 (N_2676,In_1654,N_2053);
nor U2677 (N_2677,N_1268,N_2246);
nand U2678 (N_2678,N_2132,N_2205);
and U2679 (N_2679,N_2337,N_2173);
xnor U2680 (N_2680,N_2307,N_2186);
nor U2681 (N_2681,N_1309,N_257);
or U2682 (N_2682,N_2336,N_2178);
nor U2683 (N_2683,N_2085,N_2164);
xor U2684 (N_2684,In_315,N_2318);
nand U2685 (N_2685,N_2311,N_2381);
and U2686 (N_2686,N_2229,N_1245);
and U2687 (N_2687,In_1698,N_1665);
nor U2688 (N_2688,N_2057,N_2204);
xnor U2689 (N_2689,N_2223,N_1958);
nor U2690 (N_2690,N_1545,N_2258);
nor U2691 (N_2691,N_2253,N_2056);
and U2692 (N_2692,N_1312,N_2152);
xnor U2693 (N_2693,N_1600,N_2289);
xnor U2694 (N_2694,N_1745,N_2144);
nand U2695 (N_2695,In_2123,N_1937);
nand U2696 (N_2696,N_1187,N_2393);
nor U2697 (N_2697,N_2300,N_2184);
xor U2698 (N_2698,In_2196,N_2245);
or U2699 (N_2699,N_1938,N_1864);
nor U2700 (N_2700,N_2625,N_2426);
nor U2701 (N_2701,N_2540,N_2425);
nand U2702 (N_2702,N_2594,N_2534);
or U2703 (N_2703,N_2404,N_2526);
or U2704 (N_2704,N_2627,N_2545);
xnor U2705 (N_2705,N_2610,N_2412);
and U2706 (N_2706,N_2600,N_2662);
nand U2707 (N_2707,N_2471,N_2570);
nand U2708 (N_2708,N_2410,N_2539);
or U2709 (N_2709,N_2485,N_2497);
nand U2710 (N_2710,N_2464,N_2628);
and U2711 (N_2711,N_2558,N_2634);
xnor U2712 (N_2712,N_2618,N_2605);
xor U2713 (N_2713,N_2688,N_2546);
or U2714 (N_2714,N_2595,N_2566);
or U2715 (N_2715,N_2599,N_2476);
nor U2716 (N_2716,N_2490,N_2661);
or U2717 (N_2717,N_2643,N_2547);
and U2718 (N_2718,N_2541,N_2665);
xor U2719 (N_2719,N_2685,N_2409);
or U2720 (N_2720,N_2427,N_2690);
and U2721 (N_2721,N_2517,N_2606);
xor U2722 (N_2722,N_2515,N_2576);
nor U2723 (N_2723,N_2639,N_2482);
nand U2724 (N_2724,N_2492,N_2486);
xor U2725 (N_2725,N_2556,N_2604);
xor U2726 (N_2726,N_2697,N_2520);
or U2727 (N_2727,N_2521,N_2589);
or U2728 (N_2728,N_2613,N_2455);
nor U2729 (N_2729,N_2419,N_2571);
nor U2730 (N_2730,N_2696,N_2569);
or U2731 (N_2731,N_2544,N_2514);
or U2732 (N_2732,N_2659,N_2684);
and U2733 (N_2733,N_2692,N_2417);
nor U2734 (N_2734,N_2565,N_2648);
and U2735 (N_2735,N_2585,N_2654);
and U2736 (N_2736,N_2527,N_2491);
and U2737 (N_2737,N_2531,N_2522);
or U2738 (N_2738,N_2577,N_2550);
xor U2739 (N_2739,N_2588,N_2602);
nor U2740 (N_2740,N_2532,N_2467);
nor U2741 (N_2741,N_2607,N_2411);
nand U2742 (N_2742,N_2584,N_2587);
or U2743 (N_2743,N_2528,N_2626);
nor U2744 (N_2744,N_2683,N_2500);
and U2745 (N_2745,N_2524,N_2611);
xnor U2746 (N_2746,N_2578,N_2616);
nand U2747 (N_2747,N_2601,N_2575);
nand U2748 (N_2748,N_2538,N_2449);
nand U2749 (N_2749,N_2580,N_2478);
xnor U2750 (N_2750,N_2676,N_2430);
nor U2751 (N_2751,N_2452,N_2622);
and U2752 (N_2752,N_2420,N_2621);
nor U2753 (N_2753,N_2504,N_2590);
xnor U2754 (N_2754,N_2433,N_2529);
nor U2755 (N_2755,N_2472,N_2615);
xor U2756 (N_2756,N_2463,N_2623);
or U2757 (N_2757,N_2651,N_2415);
and U2758 (N_2758,N_2592,N_2416);
nand U2759 (N_2759,N_2542,N_2630);
and U2760 (N_2760,N_2436,N_2445);
xor U2761 (N_2761,N_2653,N_2496);
nor U2762 (N_2762,N_2675,N_2687);
nand U2763 (N_2763,N_2477,N_2493);
xor U2764 (N_2764,N_2509,N_2406);
xor U2765 (N_2765,N_2667,N_2564);
xnor U2766 (N_2766,N_2466,N_2402);
or U2767 (N_2767,N_2439,N_2462);
and U2768 (N_2768,N_2597,N_2465);
or U2769 (N_2769,N_2553,N_2640);
nor U2770 (N_2770,N_2682,N_2423);
and U2771 (N_2771,N_2457,N_2518);
nor U2772 (N_2772,N_2668,N_2473);
nand U2773 (N_2773,N_2647,N_2519);
xnor U2774 (N_2774,N_2499,N_2428);
xor U2775 (N_2775,N_2503,N_2620);
and U2776 (N_2776,N_2549,N_2579);
and U2777 (N_2777,N_2679,N_2699);
and U2778 (N_2778,N_2638,N_2502);
nand U2779 (N_2779,N_2645,N_2568);
or U2780 (N_2780,N_2695,N_2669);
or U2781 (N_2781,N_2637,N_2484);
nand U2782 (N_2782,N_2450,N_2586);
xor U2783 (N_2783,N_2552,N_2469);
or U2784 (N_2784,N_2510,N_2663);
xnor U2785 (N_2785,N_2437,N_2656);
nand U2786 (N_2786,N_2421,N_2442);
nor U2787 (N_2787,N_2678,N_2448);
or U2788 (N_2788,N_2480,N_2596);
and U2789 (N_2789,N_2516,N_2495);
xor U2790 (N_2790,N_2631,N_2508);
or U2791 (N_2791,N_2536,N_2635);
nand U2792 (N_2792,N_2475,N_2543);
nand U2793 (N_2793,N_2481,N_2693);
nor U2794 (N_2794,N_2501,N_2424);
xor U2795 (N_2795,N_2657,N_2435);
xnor U2796 (N_2796,N_2672,N_2468);
nor U2797 (N_2797,N_2649,N_2507);
or U2798 (N_2798,N_2574,N_2664);
and U2799 (N_2799,N_2670,N_2535);
or U2800 (N_2800,N_2513,N_2418);
xor U2801 (N_2801,N_2660,N_2689);
nor U2802 (N_2802,N_2608,N_2461);
nor U2803 (N_2803,N_2488,N_2573);
xor U2804 (N_2804,N_2459,N_2686);
and U2805 (N_2805,N_2642,N_2698);
nand U2806 (N_2806,N_2505,N_2438);
or U2807 (N_2807,N_2440,N_2431);
and U2808 (N_2808,N_2453,N_2629);
and U2809 (N_2809,N_2633,N_2456);
nand U2810 (N_2810,N_2454,N_2644);
nor U2811 (N_2811,N_2562,N_2636);
nand U2812 (N_2812,N_2498,N_2460);
or U2813 (N_2813,N_2603,N_2474);
nor U2814 (N_2814,N_2494,N_2432);
nor U2815 (N_2815,N_2677,N_2487);
and U2816 (N_2816,N_2674,N_2646);
nand U2817 (N_2817,N_2658,N_2408);
nand U2818 (N_2818,N_2523,N_2512);
xnor U2819 (N_2819,N_2407,N_2612);
xor U2820 (N_2820,N_2561,N_2444);
nand U2821 (N_2821,N_2403,N_2655);
nand U2822 (N_2822,N_2548,N_2614);
or U2823 (N_2823,N_2434,N_2650);
or U2824 (N_2824,N_2429,N_2506);
nor U2825 (N_2825,N_2593,N_2447);
nor U2826 (N_2826,N_2400,N_2422);
nand U2827 (N_2827,N_2591,N_2563);
xnor U2828 (N_2828,N_2572,N_2557);
or U2829 (N_2829,N_2666,N_2441);
xor U2830 (N_2830,N_2559,N_2483);
nand U2831 (N_2831,N_2533,N_2555);
or U2832 (N_2832,N_2583,N_2673);
or U2833 (N_2833,N_2458,N_2598);
xnor U2834 (N_2834,N_2619,N_2641);
nand U2835 (N_2835,N_2405,N_2581);
nor U2836 (N_2836,N_2681,N_2671);
and U2837 (N_2837,N_2554,N_2652);
and U2838 (N_2838,N_2413,N_2451);
or U2839 (N_2839,N_2525,N_2530);
nor U2840 (N_2840,N_2551,N_2511);
xnor U2841 (N_2841,N_2489,N_2691);
or U2842 (N_2842,N_2609,N_2582);
and U2843 (N_2843,N_2479,N_2414);
or U2844 (N_2844,N_2680,N_2632);
xor U2845 (N_2845,N_2617,N_2446);
nand U2846 (N_2846,N_2537,N_2694);
xnor U2847 (N_2847,N_2567,N_2470);
and U2848 (N_2848,N_2560,N_2624);
xnor U2849 (N_2849,N_2443,N_2401);
and U2850 (N_2850,N_2568,N_2674);
nand U2851 (N_2851,N_2570,N_2468);
xor U2852 (N_2852,N_2405,N_2639);
and U2853 (N_2853,N_2559,N_2496);
nor U2854 (N_2854,N_2522,N_2463);
and U2855 (N_2855,N_2448,N_2514);
and U2856 (N_2856,N_2463,N_2433);
xnor U2857 (N_2857,N_2609,N_2573);
or U2858 (N_2858,N_2436,N_2437);
xnor U2859 (N_2859,N_2517,N_2662);
nand U2860 (N_2860,N_2443,N_2457);
nor U2861 (N_2861,N_2556,N_2593);
nor U2862 (N_2862,N_2592,N_2461);
xnor U2863 (N_2863,N_2655,N_2540);
nand U2864 (N_2864,N_2508,N_2412);
or U2865 (N_2865,N_2616,N_2418);
nor U2866 (N_2866,N_2606,N_2643);
nor U2867 (N_2867,N_2569,N_2606);
nor U2868 (N_2868,N_2421,N_2449);
nand U2869 (N_2869,N_2628,N_2692);
and U2870 (N_2870,N_2513,N_2423);
nand U2871 (N_2871,N_2551,N_2536);
or U2872 (N_2872,N_2593,N_2650);
nor U2873 (N_2873,N_2479,N_2692);
or U2874 (N_2874,N_2695,N_2575);
nand U2875 (N_2875,N_2515,N_2540);
nor U2876 (N_2876,N_2604,N_2653);
and U2877 (N_2877,N_2650,N_2568);
nor U2878 (N_2878,N_2489,N_2403);
nand U2879 (N_2879,N_2696,N_2639);
or U2880 (N_2880,N_2434,N_2548);
xor U2881 (N_2881,N_2528,N_2436);
and U2882 (N_2882,N_2647,N_2601);
nor U2883 (N_2883,N_2529,N_2631);
or U2884 (N_2884,N_2411,N_2483);
or U2885 (N_2885,N_2677,N_2434);
nor U2886 (N_2886,N_2635,N_2628);
nand U2887 (N_2887,N_2663,N_2557);
or U2888 (N_2888,N_2478,N_2626);
nor U2889 (N_2889,N_2502,N_2467);
and U2890 (N_2890,N_2437,N_2508);
and U2891 (N_2891,N_2451,N_2545);
and U2892 (N_2892,N_2480,N_2643);
xnor U2893 (N_2893,N_2578,N_2696);
and U2894 (N_2894,N_2412,N_2524);
nor U2895 (N_2895,N_2639,N_2535);
and U2896 (N_2896,N_2479,N_2554);
and U2897 (N_2897,N_2648,N_2470);
nand U2898 (N_2898,N_2580,N_2518);
and U2899 (N_2899,N_2417,N_2473);
and U2900 (N_2900,N_2411,N_2462);
and U2901 (N_2901,N_2676,N_2465);
xnor U2902 (N_2902,N_2530,N_2521);
nand U2903 (N_2903,N_2445,N_2419);
and U2904 (N_2904,N_2535,N_2573);
or U2905 (N_2905,N_2665,N_2624);
or U2906 (N_2906,N_2542,N_2469);
nand U2907 (N_2907,N_2520,N_2474);
xnor U2908 (N_2908,N_2630,N_2430);
nor U2909 (N_2909,N_2416,N_2470);
xor U2910 (N_2910,N_2403,N_2552);
nor U2911 (N_2911,N_2571,N_2432);
xor U2912 (N_2912,N_2617,N_2451);
and U2913 (N_2913,N_2566,N_2416);
nor U2914 (N_2914,N_2640,N_2683);
and U2915 (N_2915,N_2692,N_2606);
and U2916 (N_2916,N_2487,N_2631);
nand U2917 (N_2917,N_2669,N_2687);
and U2918 (N_2918,N_2675,N_2654);
or U2919 (N_2919,N_2634,N_2654);
nor U2920 (N_2920,N_2697,N_2588);
and U2921 (N_2921,N_2578,N_2638);
nor U2922 (N_2922,N_2402,N_2462);
and U2923 (N_2923,N_2472,N_2466);
nand U2924 (N_2924,N_2597,N_2622);
and U2925 (N_2925,N_2552,N_2451);
and U2926 (N_2926,N_2696,N_2447);
and U2927 (N_2927,N_2498,N_2579);
or U2928 (N_2928,N_2588,N_2505);
nor U2929 (N_2929,N_2584,N_2422);
nand U2930 (N_2930,N_2535,N_2617);
or U2931 (N_2931,N_2600,N_2556);
nor U2932 (N_2932,N_2575,N_2480);
or U2933 (N_2933,N_2572,N_2542);
nand U2934 (N_2934,N_2519,N_2585);
or U2935 (N_2935,N_2636,N_2662);
and U2936 (N_2936,N_2697,N_2639);
or U2937 (N_2937,N_2699,N_2504);
nor U2938 (N_2938,N_2545,N_2435);
nand U2939 (N_2939,N_2576,N_2567);
or U2940 (N_2940,N_2522,N_2659);
nand U2941 (N_2941,N_2447,N_2515);
or U2942 (N_2942,N_2553,N_2670);
or U2943 (N_2943,N_2615,N_2508);
or U2944 (N_2944,N_2630,N_2446);
or U2945 (N_2945,N_2684,N_2667);
and U2946 (N_2946,N_2492,N_2526);
or U2947 (N_2947,N_2508,N_2683);
nor U2948 (N_2948,N_2535,N_2471);
nor U2949 (N_2949,N_2607,N_2591);
xor U2950 (N_2950,N_2505,N_2611);
nor U2951 (N_2951,N_2478,N_2441);
and U2952 (N_2952,N_2515,N_2626);
xor U2953 (N_2953,N_2642,N_2471);
and U2954 (N_2954,N_2543,N_2608);
and U2955 (N_2955,N_2648,N_2409);
and U2956 (N_2956,N_2427,N_2590);
and U2957 (N_2957,N_2644,N_2565);
and U2958 (N_2958,N_2675,N_2663);
nor U2959 (N_2959,N_2653,N_2590);
and U2960 (N_2960,N_2404,N_2685);
or U2961 (N_2961,N_2474,N_2680);
nand U2962 (N_2962,N_2427,N_2462);
nand U2963 (N_2963,N_2539,N_2486);
and U2964 (N_2964,N_2467,N_2493);
xnor U2965 (N_2965,N_2517,N_2410);
or U2966 (N_2966,N_2573,N_2611);
nand U2967 (N_2967,N_2632,N_2449);
or U2968 (N_2968,N_2463,N_2487);
xor U2969 (N_2969,N_2484,N_2505);
xor U2970 (N_2970,N_2679,N_2665);
nand U2971 (N_2971,N_2523,N_2522);
nor U2972 (N_2972,N_2471,N_2671);
xor U2973 (N_2973,N_2501,N_2667);
nand U2974 (N_2974,N_2588,N_2535);
and U2975 (N_2975,N_2479,N_2453);
nor U2976 (N_2976,N_2460,N_2461);
nand U2977 (N_2977,N_2400,N_2416);
nor U2978 (N_2978,N_2612,N_2586);
xor U2979 (N_2979,N_2547,N_2505);
or U2980 (N_2980,N_2653,N_2699);
xor U2981 (N_2981,N_2665,N_2657);
nor U2982 (N_2982,N_2522,N_2687);
xnor U2983 (N_2983,N_2482,N_2574);
or U2984 (N_2984,N_2511,N_2476);
nor U2985 (N_2985,N_2486,N_2490);
nor U2986 (N_2986,N_2622,N_2431);
and U2987 (N_2987,N_2560,N_2469);
or U2988 (N_2988,N_2605,N_2580);
xor U2989 (N_2989,N_2402,N_2681);
or U2990 (N_2990,N_2494,N_2599);
or U2991 (N_2991,N_2655,N_2678);
xor U2992 (N_2992,N_2448,N_2645);
xnor U2993 (N_2993,N_2439,N_2405);
or U2994 (N_2994,N_2689,N_2620);
nand U2995 (N_2995,N_2581,N_2570);
nand U2996 (N_2996,N_2616,N_2456);
xnor U2997 (N_2997,N_2492,N_2400);
and U2998 (N_2998,N_2482,N_2648);
xor U2999 (N_2999,N_2670,N_2421);
or U3000 (N_3000,N_2838,N_2785);
xnor U3001 (N_3001,N_2819,N_2750);
nand U3002 (N_3002,N_2742,N_2964);
nor U3003 (N_3003,N_2725,N_2765);
nor U3004 (N_3004,N_2884,N_2780);
and U3005 (N_3005,N_2961,N_2745);
nor U3006 (N_3006,N_2933,N_2887);
nand U3007 (N_3007,N_2763,N_2712);
nor U3008 (N_3008,N_2892,N_2918);
nor U3009 (N_3009,N_2867,N_2718);
xnor U3010 (N_3010,N_2928,N_2782);
xor U3011 (N_3011,N_2898,N_2743);
nand U3012 (N_3012,N_2760,N_2879);
xnor U3013 (N_3013,N_2902,N_2793);
xor U3014 (N_3014,N_2886,N_2787);
nor U3015 (N_3015,N_2876,N_2901);
or U3016 (N_3016,N_2741,N_2940);
and U3017 (N_3017,N_2754,N_2791);
or U3018 (N_3018,N_2894,N_2783);
or U3019 (N_3019,N_2929,N_2857);
nor U3020 (N_3020,N_2922,N_2915);
or U3021 (N_3021,N_2871,N_2828);
nor U3022 (N_3022,N_2948,N_2988);
nor U3023 (N_3023,N_2885,N_2727);
nand U3024 (N_3024,N_2989,N_2888);
nor U3025 (N_3025,N_2721,N_2708);
xnor U3026 (N_3026,N_2702,N_2821);
nand U3027 (N_3027,N_2811,N_2963);
xnor U3028 (N_3028,N_2706,N_2805);
or U3029 (N_3029,N_2955,N_2970);
xor U3030 (N_3030,N_2959,N_2749);
nor U3031 (N_3031,N_2790,N_2996);
nand U3032 (N_3032,N_2992,N_2858);
and U3033 (N_3033,N_2766,N_2893);
xnor U3034 (N_3034,N_2987,N_2936);
nor U3035 (N_3035,N_2939,N_2736);
nand U3036 (N_3036,N_2903,N_2951);
nand U3037 (N_3037,N_2907,N_2826);
nor U3038 (N_3038,N_2817,N_2729);
nand U3039 (N_3039,N_2853,N_2877);
nor U3040 (N_3040,N_2966,N_2920);
or U3041 (N_3041,N_2769,N_2701);
or U3042 (N_3042,N_2971,N_2883);
nand U3043 (N_3043,N_2809,N_2734);
xnor U3044 (N_3044,N_2849,N_2968);
nor U3045 (N_3045,N_2947,N_2975);
nor U3046 (N_3046,N_2825,N_2764);
or U3047 (N_3047,N_2820,N_2722);
xnor U3048 (N_3048,N_2895,N_2733);
or U3049 (N_3049,N_2823,N_2812);
xnor U3050 (N_3050,N_2717,N_2934);
or U3051 (N_3051,N_2753,N_2930);
or U3052 (N_3052,N_2716,N_2709);
and U3053 (N_3053,N_2735,N_2796);
nand U3054 (N_3054,N_2831,N_2911);
nand U3055 (N_3055,N_2932,N_2843);
nor U3056 (N_3056,N_2899,N_2771);
or U3057 (N_3057,N_2962,N_2788);
nor U3058 (N_3058,N_2748,N_2967);
and U3059 (N_3059,N_2778,N_2839);
nor U3060 (N_3060,N_2744,N_2710);
xnor U3061 (N_3061,N_2739,N_2792);
xnor U3062 (N_3062,N_2991,N_2881);
and U3063 (N_3063,N_2943,N_2824);
nor U3064 (N_3064,N_2714,N_2807);
or U3065 (N_3065,N_2946,N_2995);
and U3066 (N_3066,N_2910,N_2762);
nor U3067 (N_3067,N_2954,N_2861);
nand U3068 (N_3068,N_2751,N_2784);
nand U3069 (N_3069,N_2836,N_2972);
and U3070 (N_3070,N_2850,N_2869);
nand U3071 (N_3071,N_2925,N_2866);
and U3072 (N_3072,N_2982,N_2956);
nor U3073 (N_3073,N_2700,N_2795);
or U3074 (N_3074,N_2832,N_2728);
and U3075 (N_3075,N_2957,N_2880);
nor U3076 (N_3076,N_2834,N_2985);
and U3077 (N_3077,N_2798,N_2874);
xnor U3078 (N_3078,N_2757,N_2814);
or U3079 (N_3079,N_2747,N_2740);
xnor U3080 (N_3080,N_2916,N_2865);
and U3081 (N_3081,N_2859,N_2997);
xnor U3082 (N_3082,N_2862,N_2905);
xnor U3083 (N_3083,N_2958,N_2801);
xnor U3084 (N_3084,N_2789,N_2837);
or U3085 (N_3085,N_2984,N_2856);
nor U3086 (N_3086,N_2917,N_2949);
nor U3087 (N_3087,N_2923,N_2974);
nor U3088 (N_3088,N_2841,N_2931);
xor U3089 (N_3089,N_2908,N_2794);
nand U3090 (N_3090,N_2707,N_2830);
and U3091 (N_3091,N_2950,N_2761);
nand U3092 (N_3092,N_2829,N_2840);
and U3093 (N_3093,N_2803,N_2855);
and U3094 (N_3094,N_2779,N_2800);
or U3095 (N_3095,N_2965,N_2758);
nor U3096 (N_3096,N_2797,N_2810);
xnor U3097 (N_3097,N_2873,N_2815);
nor U3098 (N_3098,N_2937,N_2724);
and U3099 (N_3099,N_2924,N_2777);
and U3100 (N_3100,N_2852,N_2711);
or U3101 (N_3101,N_2868,N_2896);
or U3102 (N_3102,N_2994,N_2851);
and U3103 (N_3103,N_2926,N_2914);
xnor U3104 (N_3104,N_2993,N_2770);
xnor U3105 (N_3105,N_2715,N_2818);
nand U3106 (N_3106,N_2941,N_2882);
and U3107 (N_3107,N_2842,N_2808);
xor U3108 (N_3108,N_2844,N_2909);
and U3109 (N_3109,N_2775,N_2953);
nand U3110 (N_3110,N_2904,N_2723);
or U3111 (N_3111,N_2768,N_2872);
nor U3112 (N_3112,N_2713,N_2816);
nor U3113 (N_3113,N_2860,N_2813);
nor U3114 (N_3114,N_2935,N_2774);
nor U3115 (N_3115,N_2978,N_2833);
xnor U3116 (N_3116,N_2878,N_2731);
and U3117 (N_3117,N_2705,N_2952);
nand U3118 (N_3118,N_2786,N_2848);
nor U3119 (N_3119,N_2979,N_2846);
xor U3120 (N_3120,N_2980,N_2983);
and U3121 (N_3121,N_2890,N_2863);
xnor U3122 (N_3122,N_2960,N_2942);
nand U3123 (N_3123,N_2938,N_2776);
nand U3124 (N_3124,N_2921,N_2737);
xor U3125 (N_3125,N_2976,N_2755);
xnor U3126 (N_3126,N_2719,N_2998);
or U3127 (N_3127,N_2802,N_2977);
and U3128 (N_3128,N_2759,N_2772);
nor U3129 (N_3129,N_2870,N_2704);
or U3130 (N_3130,N_2720,N_2875);
and U3131 (N_3131,N_2900,N_2756);
or U3132 (N_3132,N_2944,N_2973);
nor U3133 (N_3133,N_2945,N_2703);
xor U3134 (N_3134,N_2773,N_2746);
and U3135 (N_3135,N_2847,N_2889);
nand U3136 (N_3136,N_2897,N_2822);
xor U3137 (N_3137,N_2913,N_2799);
and U3138 (N_3138,N_2969,N_2912);
xnor U3139 (N_3139,N_2919,N_2864);
nor U3140 (N_3140,N_2835,N_2804);
or U3141 (N_3141,N_2891,N_2827);
nand U3142 (N_3142,N_2732,N_2726);
xor U3143 (N_3143,N_2845,N_2767);
nor U3144 (N_3144,N_2854,N_2981);
nor U3145 (N_3145,N_2927,N_2806);
nor U3146 (N_3146,N_2738,N_2990);
nor U3147 (N_3147,N_2986,N_2730);
and U3148 (N_3148,N_2906,N_2781);
or U3149 (N_3149,N_2752,N_2999);
and U3150 (N_3150,N_2982,N_2996);
nor U3151 (N_3151,N_2986,N_2900);
nor U3152 (N_3152,N_2921,N_2760);
and U3153 (N_3153,N_2801,N_2758);
or U3154 (N_3154,N_2958,N_2821);
nor U3155 (N_3155,N_2882,N_2710);
xor U3156 (N_3156,N_2983,N_2886);
nor U3157 (N_3157,N_2720,N_2974);
nor U3158 (N_3158,N_2734,N_2703);
and U3159 (N_3159,N_2947,N_2712);
nand U3160 (N_3160,N_2927,N_2739);
or U3161 (N_3161,N_2975,N_2984);
or U3162 (N_3162,N_2932,N_2884);
nand U3163 (N_3163,N_2947,N_2768);
nand U3164 (N_3164,N_2837,N_2987);
nor U3165 (N_3165,N_2892,N_2941);
xor U3166 (N_3166,N_2811,N_2761);
nand U3167 (N_3167,N_2822,N_2730);
or U3168 (N_3168,N_2716,N_2787);
nand U3169 (N_3169,N_2835,N_2926);
nor U3170 (N_3170,N_2738,N_2719);
or U3171 (N_3171,N_2926,N_2742);
nand U3172 (N_3172,N_2854,N_2732);
nand U3173 (N_3173,N_2999,N_2898);
nor U3174 (N_3174,N_2750,N_2996);
nor U3175 (N_3175,N_2974,N_2911);
nand U3176 (N_3176,N_2760,N_2882);
xnor U3177 (N_3177,N_2843,N_2817);
xnor U3178 (N_3178,N_2886,N_2793);
or U3179 (N_3179,N_2956,N_2746);
nand U3180 (N_3180,N_2894,N_2909);
nor U3181 (N_3181,N_2883,N_2776);
and U3182 (N_3182,N_2856,N_2783);
and U3183 (N_3183,N_2760,N_2864);
nor U3184 (N_3184,N_2992,N_2750);
or U3185 (N_3185,N_2718,N_2893);
or U3186 (N_3186,N_2824,N_2718);
nand U3187 (N_3187,N_2832,N_2815);
nand U3188 (N_3188,N_2777,N_2810);
xor U3189 (N_3189,N_2798,N_2820);
or U3190 (N_3190,N_2757,N_2967);
nor U3191 (N_3191,N_2741,N_2914);
nand U3192 (N_3192,N_2724,N_2885);
nand U3193 (N_3193,N_2869,N_2959);
or U3194 (N_3194,N_2843,N_2791);
nor U3195 (N_3195,N_2960,N_2775);
nand U3196 (N_3196,N_2966,N_2766);
or U3197 (N_3197,N_2852,N_2710);
xnor U3198 (N_3198,N_2792,N_2896);
nor U3199 (N_3199,N_2708,N_2975);
nand U3200 (N_3200,N_2800,N_2907);
nor U3201 (N_3201,N_2726,N_2829);
and U3202 (N_3202,N_2799,N_2895);
or U3203 (N_3203,N_2884,N_2981);
nor U3204 (N_3204,N_2716,N_2711);
nand U3205 (N_3205,N_2822,N_2923);
or U3206 (N_3206,N_2911,N_2988);
and U3207 (N_3207,N_2949,N_2970);
and U3208 (N_3208,N_2849,N_2777);
nor U3209 (N_3209,N_2970,N_2902);
and U3210 (N_3210,N_2991,N_2811);
or U3211 (N_3211,N_2919,N_2958);
or U3212 (N_3212,N_2732,N_2842);
or U3213 (N_3213,N_2766,N_2722);
or U3214 (N_3214,N_2820,N_2909);
and U3215 (N_3215,N_2878,N_2784);
or U3216 (N_3216,N_2839,N_2972);
xor U3217 (N_3217,N_2799,N_2995);
or U3218 (N_3218,N_2955,N_2974);
xnor U3219 (N_3219,N_2708,N_2967);
nand U3220 (N_3220,N_2808,N_2927);
xnor U3221 (N_3221,N_2934,N_2782);
nand U3222 (N_3222,N_2709,N_2957);
xor U3223 (N_3223,N_2773,N_2936);
and U3224 (N_3224,N_2939,N_2848);
nand U3225 (N_3225,N_2862,N_2837);
and U3226 (N_3226,N_2804,N_2719);
or U3227 (N_3227,N_2716,N_2931);
xor U3228 (N_3228,N_2910,N_2765);
nor U3229 (N_3229,N_2745,N_2756);
and U3230 (N_3230,N_2841,N_2718);
xnor U3231 (N_3231,N_2929,N_2999);
and U3232 (N_3232,N_2857,N_2935);
and U3233 (N_3233,N_2763,N_2914);
and U3234 (N_3234,N_2931,N_2975);
xnor U3235 (N_3235,N_2825,N_2750);
nand U3236 (N_3236,N_2894,N_2792);
and U3237 (N_3237,N_2884,N_2963);
nor U3238 (N_3238,N_2889,N_2757);
or U3239 (N_3239,N_2975,N_2953);
and U3240 (N_3240,N_2942,N_2989);
and U3241 (N_3241,N_2947,N_2800);
nor U3242 (N_3242,N_2856,N_2723);
xnor U3243 (N_3243,N_2920,N_2802);
nand U3244 (N_3244,N_2983,N_2844);
xnor U3245 (N_3245,N_2857,N_2819);
nand U3246 (N_3246,N_2881,N_2841);
nand U3247 (N_3247,N_2827,N_2849);
nand U3248 (N_3248,N_2994,N_2929);
xor U3249 (N_3249,N_2756,N_2888);
nand U3250 (N_3250,N_2701,N_2720);
and U3251 (N_3251,N_2893,N_2861);
nand U3252 (N_3252,N_2998,N_2840);
nand U3253 (N_3253,N_2936,N_2721);
nor U3254 (N_3254,N_2822,N_2885);
xor U3255 (N_3255,N_2871,N_2757);
nor U3256 (N_3256,N_2726,N_2866);
xnor U3257 (N_3257,N_2988,N_2719);
xor U3258 (N_3258,N_2927,N_2822);
nand U3259 (N_3259,N_2853,N_2712);
xnor U3260 (N_3260,N_2898,N_2782);
nand U3261 (N_3261,N_2898,N_2908);
nor U3262 (N_3262,N_2908,N_2779);
nand U3263 (N_3263,N_2752,N_2846);
and U3264 (N_3264,N_2715,N_2780);
xnor U3265 (N_3265,N_2887,N_2870);
xnor U3266 (N_3266,N_2830,N_2826);
nor U3267 (N_3267,N_2868,N_2848);
nor U3268 (N_3268,N_2966,N_2931);
xnor U3269 (N_3269,N_2823,N_2878);
or U3270 (N_3270,N_2910,N_2866);
xnor U3271 (N_3271,N_2868,N_2736);
nand U3272 (N_3272,N_2901,N_2729);
xor U3273 (N_3273,N_2978,N_2731);
or U3274 (N_3274,N_2842,N_2848);
nand U3275 (N_3275,N_2950,N_2749);
nor U3276 (N_3276,N_2844,N_2928);
nand U3277 (N_3277,N_2841,N_2732);
and U3278 (N_3278,N_2965,N_2721);
nand U3279 (N_3279,N_2846,N_2899);
nand U3280 (N_3280,N_2750,N_2735);
and U3281 (N_3281,N_2830,N_2778);
nor U3282 (N_3282,N_2948,N_2989);
nand U3283 (N_3283,N_2714,N_2850);
and U3284 (N_3284,N_2750,N_2803);
nand U3285 (N_3285,N_2766,N_2937);
and U3286 (N_3286,N_2790,N_2743);
nand U3287 (N_3287,N_2876,N_2976);
nor U3288 (N_3288,N_2855,N_2851);
nor U3289 (N_3289,N_2817,N_2815);
xnor U3290 (N_3290,N_2829,N_2856);
or U3291 (N_3291,N_2985,N_2780);
xor U3292 (N_3292,N_2880,N_2830);
xor U3293 (N_3293,N_2771,N_2873);
nor U3294 (N_3294,N_2981,N_2751);
xor U3295 (N_3295,N_2908,N_2920);
xor U3296 (N_3296,N_2947,N_2700);
nor U3297 (N_3297,N_2930,N_2747);
nor U3298 (N_3298,N_2929,N_2806);
xnor U3299 (N_3299,N_2941,N_2944);
xor U3300 (N_3300,N_3038,N_3209);
nand U3301 (N_3301,N_3231,N_3261);
xnor U3302 (N_3302,N_3126,N_3274);
xor U3303 (N_3303,N_3064,N_3028);
xor U3304 (N_3304,N_3153,N_3152);
nor U3305 (N_3305,N_3251,N_3241);
and U3306 (N_3306,N_3063,N_3086);
xor U3307 (N_3307,N_3098,N_3256);
or U3308 (N_3308,N_3083,N_3096);
nand U3309 (N_3309,N_3283,N_3151);
nor U3310 (N_3310,N_3087,N_3026);
or U3311 (N_3311,N_3162,N_3191);
nor U3312 (N_3312,N_3154,N_3131);
or U3313 (N_3313,N_3127,N_3246);
nor U3314 (N_3314,N_3088,N_3085);
xor U3315 (N_3315,N_3168,N_3189);
nand U3316 (N_3316,N_3128,N_3023);
xor U3317 (N_3317,N_3116,N_3198);
nand U3318 (N_3318,N_3172,N_3039);
nand U3319 (N_3319,N_3106,N_3067);
or U3320 (N_3320,N_3125,N_3214);
nor U3321 (N_3321,N_3091,N_3270);
and U3322 (N_3322,N_3148,N_3130);
and U3323 (N_3323,N_3236,N_3139);
nor U3324 (N_3324,N_3275,N_3069);
nand U3325 (N_3325,N_3277,N_3167);
or U3326 (N_3326,N_3158,N_3043);
xnor U3327 (N_3327,N_3239,N_3147);
xnor U3328 (N_3328,N_3273,N_3247);
or U3329 (N_3329,N_3201,N_3216);
or U3330 (N_3330,N_3193,N_3218);
and U3331 (N_3331,N_3264,N_3225);
xnor U3332 (N_3332,N_3245,N_3030);
xnor U3333 (N_3333,N_3047,N_3029);
nand U3334 (N_3334,N_3068,N_3137);
nor U3335 (N_3335,N_3017,N_3081);
and U3336 (N_3336,N_3119,N_3159);
nor U3337 (N_3337,N_3000,N_3296);
nor U3338 (N_3338,N_3242,N_3123);
nor U3339 (N_3339,N_3093,N_3124);
nand U3340 (N_3340,N_3019,N_3141);
nor U3341 (N_3341,N_3110,N_3161);
nand U3342 (N_3342,N_3072,N_3033);
nand U3343 (N_3343,N_3184,N_3135);
xnor U3344 (N_3344,N_3053,N_3260);
and U3345 (N_3345,N_3226,N_3004);
xor U3346 (N_3346,N_3206,N_3292);
xnor U3347 (N_3347,N_3012,N_3205);
xnor U3348 (N_3348,N_3133,N_3221);
nand U3349 (N_3349,N_3213,N_3006);
and U3350 (N_3350,N_3284,N_3257);
or U3351 (N_3351,N_3009,N_3014);
nor U3352 (N_3352,N_3254,N_3203);
xor U3353 (N_3353,N_3046,N_3145);
nor U3354 (N_3354,N_3049,N_3109);
xnor U3355 (N_3355,N_3045,N_3041);
xor U3356 (N_3356,N_3121,N_3117);
nor U3357 (N_3357,N_3266,N_3240);
and U3358 (N_3358,N_3015,N_3196);
nor U3359 (N_3359,N_3229,N_3078);
xnor U3360 (N_3360,N_3291,N_3056);
or U3361 (N_3361,N_3286,N_3287);
and U3362 (N_3362,N_3003,N_3020);
and U3363 (N_3363,N_3011,N_3071);
or U3364 (N_3364,N_3155,N_3080);
xnor U3365 (N_3365,N_3183,N_3024);
nand U3366 (N_3366,N_3174,N_3002);
or U3367 (N_3367,N_3101,N_3077);
and U3368 (N_3368,N_3188,N_3180);
and U3369 (N_3369,N_3212,N_3181);
nor U3370 (N_3370,N_3089,N_3007);
or U3371 (N_3371,N_3022,N_3170);
or U3372 (N_3372,N_3272,N_3095);
nand U3373 (N_3373,N_3136,N_3262);
xnor U3374 (N_3374,N_3243,N_3248);
or U3375 (N_3375,N_3237,N_3255);
and U3376 (N_3376,N_3177,N_3165);
nand U3377 (N_3377,N_3164,N_3061);
nor U3378 (N_3378,N_3105,N_3288);
xnor U3379 (N_3379,N_3271,N_3252);
and U3380 (N_3380,N_3143,N_3113);
and U3381 (N_3381,N_3142,N_3036);
xor U3382 (N_3382,N_3114,N_3025);
nor U3383 (N_3383,N_3233,N_3104);
xor U3384 (N_3384,N_3057,N_3010);
nand U3385 (N_3385,N_3055,N_3146);
nand U3386 (N_3386,N_3207,N_3235);
or U3387 (N_3387,N_3269,N_3129);
xor U3388 (N_3388,N_3250,N_3018);
nand U3389 (N_3389,N_3079,N_3108);
xor U3390 (N_3390,N_3285,N_3169);
and U3391 (N_3391,N_3008,N_3034);
nor U3392 (N_3392,N_3197,N_3279);
and U3393 (N_3393,N_3173,N_3115);
and U3394 (N_3394,N_3163,N_3199);
xnor U3395 (N_3395,N_3202,N_3032);
or U3396 (N_3396,N_3065,N_3040);
and U3397 (N_3397,N_3244,N_3132);
xnor U3398 (N_3398,N_3090,N_3060);
xnor U3399 (N_3399,N_3253,N_3295);
nand U3400 (N_3400,N_3210,N_3094);
nand U3401 (N_3401,N_3001,N_3082);
xnor U3402 (N_3402,N_3249,N_3228);
or U3403 (N_3403,N_3185,N_3016);
and U3404 (N_3404,N_3048,N_3192);
nor U3405 (N_3405,N_3186,N_3050);
or U3406 (N_3406,N_3294,N_3297);
nand U3407 (N_3407,N_3179,N_3111);
or U3408 (N_3408,N_3258,N_3289);
and U3409 (N_3409,N_3005,N_3176);
or U3410 (N_3410,N_3290,N_3182);
nor U3411 (N_3411,N_3070,N_3013);
and U3412 (N_3412,N_3021,N_3102);
nor U3413 (N_3413,N_3044,N_3073);
or U3414 (N_3414,N_3100,N_3160);
or U3415 (N_3415,N_3037,N_3149);
and U3416 (N_3416,N_3150,N_3280);
xor U3417 (N_3417,N_3076,N_3118);
nand U3418 (N_3418,N_3299,N_3267);
nor U3419 (N_3419,N_3276,N_3230);
and U3420 (N_3420,N_3175,N_3195);
nand U3421 (N_3421,N_3031,N_3238);
xnor U3422 (N_3422,N_3075,N_3120);
and U3423 (N_3423,N_3107,N_3092);
or U3424 (N_3424,N_3215,N_3062);
nor U3425 (N_3425,N_3122,N_3268);
and U3426 (N_3426,N_3227,N_3194);
xnor U3427 (N_3427,N_3265,N_3035);
xnor U3428 (N_3428,N_3051,N_3208);
xor U3429 (N_3429,N_3219,N_3281);
xor U3430 (N_3430,N_3222,N_3282);
xnor U3431 (N_3431,N_3099,N_3112);
or U3432 (N_3432,N_3058,N_3084);
or U3433 (N_3433,N_3259,N_3156);
nand U3434 (N_3434,N_3187,N_3144);
and U3435 (N_3435,N_3042,N_3190);
xnor U3436 (N_3436,N_3052,N_3097);
nand U3437 (N_3437,N_3074,N_3138);
xnor U3438 (N_3438,N_3298,N_3066);
and U3439 (N_3439,N_3178,N_3232);
and U3440 (N_3440,N_3140,N_3171);
nand U3441 (N_3441,N_3157,N_3200);
and U3442 (N_3442,N_3166,N_3027);
nand U3443 (N_3443,N_3059,N_3234);
nand U3444 (N_3444,N_3293,N_3103);
nand U3445 (N_3445,N_3278,N_3211);
nand U3446 (N_3446,N_3224,N_3217);
and U3447 (N_3447,N_3134,N_3220);
nand U3448 (N_3448,N_3223,N_3054);
or U3449 (N_3449,N_3204,N_3263);
or U3450 (N_3450,N_3212,N_3135);
or U3451 (N_3451,N_3187,N_3218);
or U3452 (N_3452,N_3029,N_3042);
nand U3453 (N_3453,N_3292,N_3101);
nand U3454 (N_3454,N_3004,N_3092);
and U3455 (N_3455,N_3168,N_3218);
and U3456 (N_3456,N_3175,N_3016);
xnor U3457 (N_3457,N_3035,N_3266);
nand U3458 (N_3458,N_3227,N_3196);
and U3459 (N_3459,N_3176,N_3298);
and U3460 (N_3460,N_3124,N_3062);
nor U3461 (N_3461,N_3232,N_3179);
or U3462 (N_3462,N_3073,N_3088);
xnor U3463 (N_3463,N_3080,N_3109);
nor U3464 (N_3464,N_3212,N_3017);
or U3465 (N_3465,N_3205,N_3230);
nand U3466 (N_3466,N_3002,N_3230);
or U3467 (N_3467,N_3078,N_3077);
and U3468 (N_3468,N_3161,N_3025);
and U3469 (N_3469,N_3002,N_3265);
xor U3470 (N_3470,N_3222,N_3174);
or U3471 (N_3471,N_3139,N_3009);
nand U3472 (N_3472,N_3270,N_3079);
nand U3473 (N_3473,N_3012,N_3126);
xnor U3474 (N_3474,N_3293,N_3202);
xor U3475 (N_3475,N_3255,N_3232);
nand U3476 (N_3476,N_3112,N_3294);
or U3477 (N_3477,N_3077,N_3082);
nor U3478 (N_3478,N_3290,N_3233);
or U3479 (N_3479,N_3242,N_3159);
or U3480 (N_3480,N_3007,N_3220);
nand U3481 (N_3481,N_3136,N_3207);
xor U3482 (N_3482,N_3077,N_3170);
nand U3483 (N_3483,N_3250,N_3131);
nand U3484 (N_3484,N_3178,N_3121);
or U3485 (N_3485,N_3293,N_3121);
nor U3486 (N_3486,N_3177,N_3291);
nor U3487 (N_3487,N_3255,N_3101);
nand U3488 (N_3488,N_3174,N_3061);
xnor U3489 (N_3489,N_3152,N_3276);
xor U3490 (N_3490,N_3043,N_3207);
xnor U3491 (N_3491,N_3163,N_3190);
xor U3492 (N_3492,N_3252,N_3161);
nor U3493 (N_3493,N_3070,N_3063);
nor U3494 (N_3494,N_3003,N_3083);
xor U3495 (N_3495,N_3119,N_3079);
xnor U3496 (N_3496,N_3274,N_3089);
xor U3497 (N_3497,N_3013,N_3050);
and U3498 (N_3498,N_3182,N_3239);
nand U3499 (N_3499,N_3266,N_3019);
nand U3500 (N_3500,N_3239,N_3144);
or U3501 (N_3501,N_3185,N_3106);
nor U3502 (N_3502,N_3073,N_3100);
or U3503 (N_3503,N_3174,N_3256);
and U3504 (N_3504,N_3097,N_3185);
xor U3505 (N_3505,N_3035,N_3074);
nand U3506 (N_3506,N_3163,N_3242);
or U3507 (N_3507,N_3166,N_3002);
or U3508 (N_3508,N_3031,N_3272);
nand U3509 (N_3509,N_3055,N_3014);
or U3510 (N_3510,N_3254,N_3182);
xnor U3511 (N_3511,N_3226,N_3202);
xor U3512 (N_3512,N_3224,N_3004);
or U3513 (N_3513,N_3267,N_3068);
and U3514 (N_3514,N_3222,N_3163);
or U3515 (N_3515,N_3015,N_3089);
xnor U3516 (N_3516,N_3163,N_3179);
and U3517 (N_3517,N_3294,N_3064);
or U3518 (N_3518,N_3204,N_3032);
or U3519 (N_3519,N_3256,N_3094);
nor U3520 (N_3520,N_3119,N_3284);
and U3521 (N_3521,N_3137,N_3005);
xnor U3522 (N_3522,N_3283,N_3231);
and U3523 (N_3523,N_3002,N_3226);
or U3524 (N_3524,N_3284,N_3295);
or U3525 (N_3525,N_3147,N_3201);
and U3526 (N_3526,N_3074,N_3077);
xnor U3527 (N_3527,N_3017,N_3214);
nor U3528 (N_3528,N_3274,N_3125);
and U3529 (N_3529,N_3175,N_3226);
nand U3530 (N_3530,N_3244,N_3136);
or U3531 (N_3531,N_3236,N_3073);
nand U3532 (N_3532,N_3286,N_3075);
and U3533 (N_3533,N_3280,N_3040);
and U3534 (N_3534,N_3213,N_3128);
and U3535 (N_3535,N_3105,N_3219);
or U3536 (N_3536,N_3023,N_3246);
nand U3537 (N_3537,N_3235,N_3164);
xnor U3538 (N_3538,N_3168,N_3222);
nor U3539 (N_3539,N_3037,N_3029);
and U3540 (N_3540,N_3084,N_3153);
or U3541 (N_3541,N_3293,N_3109);
nand U3542 (N_3542,N_3293,N_3033);
nor U3543 (N_3543,N_3289,N_3089);
xor U3544 (N_3544,N_3212,N_3188);
nor U3545 (N_3545,N_3285,N_3127);
or U3546 (N_3546,N_3192,N_3171);
nand U3547 (N_3547,N_3125,N_3041);
or U3548 (N_3548,N_3298,N_3160);
nand U3549 (N_3549,N_3283,N_3104);
xnor U3550 (N_3550,N_3076,N_3131);
xnor U3551 (N_3551,N_3193,N_3034);
nand U3552 (N_3552,N_3138,N_3082);
or U3553 (N_3553,N_3208,N_3297);
nand U3554 (N_3554,N_3110,N_3051);
or U3555 (N_3555,N_3169,N_3238);
nand U3556 (N_3556,N_3096,N_3200);
nor U3557 (N_3557,N_3280,N_3060);
xnor U3558 (N_3558,N_3179,N_3204);
and U3559 (N_3559,N_3159,N_3125);
nor U3560 (N_3560,N_3168,N_3166);
xor U3561 (N_3561,N_3079,N_3002);
nor U3562 (N_3562,N_3228,N_3242);
or U3563 (N_3563,N_3284,N_3168);
xor U3564 (N_3564,N_3294,N_3065);
or U3565 (N_3565,N_3164,N_3085);
nand U3566 (N_3566,N_3009,N_3164);
nor U3567 (N_3567,N_3008,N_3078);
xnor U3568 (N_3568,N_3135,N_3015);
and U3569 (N_3569,N_3058,N_3221);
nor U3570 (N_3570,N_3113,N_3204);
nor U3571 (N_3571,N_3254,N_3019);
nand U3572 (N_3572,N_3232,N_3080);
or U3573 (N_3573,N_3227,N_3035);
xnor U3574 (N_3574,N_3261,N_3001);
or U3575 (N_3575,N_3223,N_3073);
nor U3576 (N_3576,N_3282,N_3263);
or U3577 (N_3577,N_3021,N_3200);
and U3578 (N_3578,N_3249,N_3008);
nand U3579 (N_3579,N_3132,N_3198);
nand U3580 (N_3580,N_3153,N_3183);
nand U3581 (N_3581,N_3174,N_3121);
nand U3582 (N_3582,N_3142,N_3226);
xor U3583 (N_3583,N_3014,N_3181);
xnor U3584 (N_3584,N_3258,N_3150);
and U3585 (N_3585,N_3047,N_3158);
or U3586 (N_3586,N_3152,N_3216);
and U3587 (N_3587,N_3090,N_3267);
nand U3588 (N_3588,N_3223,N_3282);
nand U3589 (N_3589,N_3286,N_3294);
and U3590 (N_3590,N_3084,N_3193);
or U3591 (N_3591,N_3283,N_3278);
xnor U3592 (N_3592,N_3015,N_3295);
xor U3593 (N_3593,N_3045,N_3297);
nor U3594 (N_3594,N_3284,N_3189);
nor U3595 (N_3595,N_3125,N_3209);
and U3596 (N_3596,N_3100,N_3121);
nand U3597 (N_3597,N_3274,N_3206);
and U3598 (N_3598,N_3124,N_3180);
or U3599 (N_3599,N_3183,N_3294);
xnor U3600 (N_3600,N_3324,N_3585);
nor U3601 (N_3601,N_3539,N_3534);
or U3602 (N_3602,N_3571,N_3419);
or U3603 (N_3603,N_3498,N_3420);
nor U3604 (N_3604,N_3589,N_3303);
and U3605 (N_3605,N_3310,N_3400);
nand U3606 (N_3606,N_3432,N_3413);
and U3607 (N_3607,N_3320,N_3455);
xnor U3608 (N_3608,N_3450,N_3583);
or U3609 (N_3609,N_3325,N_3574);
xnor U3610 (N_3610,N_3406,N_3399);
or U3611 (N_3611,N_3497,N_3540);
or U3612 (N_3612,N_3304,N_3343);
nand U3613 (N_3613,N_3536,N_3597);
nand U3614 (N_3614,N_3469,N_3440);
xnor U3615 (N_3615,N_3431,N_3409);
xnor U3616 (N_3616,N_3551,N_3475);
and U3617 (N_3617,N_3547,N_3416);
nand U3618 (N_3618,N_3300,N_3573);
and U3619 (N_3619,N_3488,N_3356);
nand U3620 (N_3620,N_3441,N_3374);
nor U3621 (N_3621,N_3508,N_3368);
nor U3622 (N_3622,N_3372,N_3563);
xnor U3623 (N_3623,N_3579,N_3459);
nand U3624 (N_3624,N_3396,N_3433);
nor U3625 (N_3625,N_3347,N_3593);
or U3626 (N_3626,N_3595,N_3338);
nor U3627 (N_3627,N_3448,N_3403);
nand U3628 (N_3628,N_3430,N_3560);
nor U3629 (N_3629,N_3385,N_3355);
nand U3630 (N_3630,N_3516,N_3517);
xor U3631 (N_3631,N_3496,N_3504);
or U3632 (N_3632,N_3389,N_3468);
nand U3633 (N_3633,N_3442,N_3522);
nor U3634 (N_3634,N_3492,N_3477);
nand U3635 (N_3635,N_3580,N_3562);
nand U3636 (N_3636,N_3495,N_3466);
or U3637 (N_3637,N_3533,N_3371);
and U3638 (N_3638,N_3483,N_3568);
nor U3639 (N_3639,N_3353,N_3417);
and U3640 (N_3640,N_3337,N_3456);
nand U3641 (N_3641,N_3439,N_3557);
and U3642 (N_3642,N_3514,N_3546);
xnor U3643 (N_3643,N_3519,N_3373);
or U3644 (N_3644,N_3548,N_3341);
xnor U3645 (N_3645,N_3367,N_3476);
and U3646 (N_3646,N_3408,N_3532);
or U3647 (N_3647,N_3542,N_3463);
nor U3648 (N_3648,N_3319,N_3535);
nand U3649 (N_3649,N_3344,N_3305);
and U3650 (N_3650,N_3565,N_3596);
nor U3651 (N_3651,N_3474,N_3333);
xor U3652 (N_3652,N_3387,N_3379);
xor U3653 (N_3653,N_3415,N_3449);
nand U3654 (N_3654,N_3531,N_3435);
nor U3655 (N_3655,N_3552,N_3451);
xnor U3656 (N_3656,N_3566,N_3361);
and U3657 (N_3657,N_3308,N_3370);
xnor U3658 (N_3658,N_3545,N_3352);
nor U3659 (N_3659,N_3425,N_3484);
nor U3660 (N_3660,N_3502,N_3467);
nand U3661 (N_3661,N_3520,N_3453);
nand U3662 (N_3662,N_3349,N_3458);
nand U3663 (N_3663,N_3381,N_3365);
xnor U3664 (N_3664,N_3354,N_3318);
and U3665 (N_3665,N_3404,N_3598);
nand U3666 (N_3666,N_3340,N_3506);
or U3667 (N_3667,N_3584,N_3312);
and U3668 (N_3668,N_3588,N_3315);
xnor U3669 (N_3669,N_3587,N_3452);
and U3670 (N_3670,N_3329,N_3383);
nor U3671 (N_3671,N_3530,N_3541);
nor U3672 (N_3672,N_3364,N_3307);
nor U3673 (N_3673,N_3357,N_3544);
and U3674 (N_3674,N_3313,N_3422);
and U3675 (N_3675,N_3480,N_3558);
nand U3676 (N_3676,N_3369,N_3323);
and U3677 (N_3677,N_3412,N_3454);
nor U3678 (N_3678,N_3334,N_3493);
or U3679 (N_3679,N_3363,N_3576);
and U3680 (N_3680,N_3397,N_3479);
or U3681 (N_3681,N_3500,N_3486);
and U3682 (N_3682,N_3386,N_3457);
xnor U3683 (N_3683,N_3460,N_3436);
xnor U3684 (N_3684,N_3564,N_3376);
and U3685 (N_3685,N_3524,N_3342);
and U3686 (N_3686,N_3592,N_3426);
xnor U3687 (N_3687,N_3351,N_3473);
or U3688 (N_3688,N_3567,N_3366);
or U3689 (N_3689,N_3550,N_3301);
xor U3690 (N_3690,N_3393,N_3336);
nor U3691 (N_3691,N_3330,N_3461);
nand U3692 (N_3692,N_3447,N_3501);
or U3693 (N_3693,N_3377,N_3314);
nor U3694 (N_3694,N_3398,N_3311);
nor U3695 (N_3695,N_3405,N_3418);
and U3696 (N_3696,N_3316,N_3509);
nor U3697 (N_3697,N_3464,N_3481);
nand U3698 (N_3698,N_3328,N_3485);
or U3699 (N_3699,N_3554,N_3348);
nor U3700 (N_3700,N_3528,N_3331);
xnor U3701 (N_3701,N_3437,N_3309);
or U3702 (N_3702,N_3424,N_3359);
and U3703 (N_3703,N_3411,N_3339);
and U3704 (N_3704,N_3306,N_3438);
nand U3705 (N_3705,N_3443,N_3421);
nand U3706 (N_3706,N_3358,N_3378);
nand U3707 (N_3707,N_3526,N_3512);
or U3708 (N_3708,N_3577,N_3561);
or U3709 (N_3709,N_3499,N_3302);
xor U3710 (N_3710,N_3549,N_3462);
xnor U3711 (N_3711,N_3332,N_3513);
or U3712 (N_3712,N_3586,N_3382);
nand U3713 (N_3713,N_3482,N_3503);
or U3714 (N_3714,N_3578,N_3427);
nor U3715 (N_3715,N_3465,N_3472);
and U3716 (N_3716,N_3570,N_3401);
and U3717 (N_3717,N_3327,N_3591);
nand U3718 (N_3718,N_3407,N_3470);
nor U3719 (N_3719,N_3515,N_3434);
and U3720 (N_3720,N_3410,N_3525);
or U3721 (N_3721,N_3390,N_3444);
nand U3722 (N_3722,N_3599,N_3350);
or U3723 (N_3723,N_3394,N_3375);
xor U3724 (N_3724,N_3388,N_3487);
or U3725 (N_3725,N_3384,N_3537);
nor U3726 (N_3726,N_3362,N_3471);
nand U3727 (N_3727,N_3478,N_3569);
or U3728 (N_3728,N_3521,N_3490);
xor U3729 (N_3729,N_3518,N_3556);
or U3730 (N_3730,N_3360,N_3572);
nand U3731 (N_3731,N_3335,N_3529);
or U3732 (N_3732,N_3326,N_3345);
nand U3733 (N_3733,N_3380,N_3581);
xor U3734 (N_3734,N_3392,N_3505);
and U3735 (N_3735,N_3391,N_3346);
xnor U3736 (N_3736,N_3491,N_3322);
xnor U3737 (N_3737,N_3582,N_3321);
xor U3738 (N_3738,N_3445,N_3446);
nand U3739 (N_3739,N_3428,N_3510);
xnor U3740 (N_3740,N_3395,N_3429);
nand U3741 (N_3741,N_3543,N_3527);
or U3742 (N_3742,N_3414,N_3402);
nor U3743 (N_3743,N_3523,N_3317);
xor U3744 (N_3744,N_3511,N_3590);
nor U3745 (N_3745,N_3555,N_3538);
nand U3746 (N_3746,N_3553,N_3575);
nor U3747 (N_3747,N_3594,N_3489);
and U3748 (N_3748,N_3507,N_3494);
xor U3749 (N_3749,N_3423,N_3559);
xor U3750 (N_3750,N_3357,N_3343);
and U3751 (N_3751,N_3300,N_3361);
or U3752 (N_3752,N_3368,N_3421);
xor U3753 (N_3753,N_3576,N_3588);
and U3754 (N_3754,N_3484,N_3368);
nor U3755 (N_3755,N_3590,N_3380);
and U3756 (N_3756,N_3571,N_3397);
or U3757 (N_3757,N_3348,N_3514);
nand U3758 (N_3758,N_3397,N_3529);
nor U3759 (N_3759,N_3329,N_3481);
nand U3760 (N_3760,N_3403,N_3419);
nor U3761 (N_3761,N_3556,N_3584);
or U3762 (N_3762,N_3313,N_3331);
xnor U3763 (N_3763,N_3406,N_3544);
and U3764 (N_3764,N_3374,N_3426);
nor U3765 (N_3765,N_3490,N_3354);
xnor U3766 (N_3766,N_3314,N_3365);
xnor U3767 (N_3767,N_3402,N_3328);
nand U3768 (N_3768,N_3409,N_3402);
nand U3769 (N_3769,N_3553,N_3493);
and U3770 (N_3770,N_3469,N_3527);
nand U3771 (N_3771,N_3472,N_3332);
or U3772 (N_3772,N_3554,N_3498);
nor U3773 (N_3773,N_3391,N_3547);
and U3774 (N_3774,N_3313,N_3405);
nand U3775 (N_3775,N_3331,N_3556);
and U3776 (N_3776,N_3367,N_3526);
nor U3777 (N_3777,N_3540,N_3495);
nand U3778 (N_3778,N_3593,N_3541);
nand U3779 (N_3779,N_3386,N_3327);
and U3780 (N_3780,N_3306,N_3321);
or U3781 (N_3781,N_3379,N_3562);
xor U3782 (N_3782,N_3417,N_3423);
nand U3783 (N_3783,N_3349,N_3528);
and U3784 (N_3784,N_3473,N_3302);
xnor U3785 (N_3785,N_3571,N_3317);
and U3786 (N_3786,N_3318,N_3382);
or U3787 (N_3787,N_3427,N_3384);
nor U3788 (N_3788,N_3358,N_3508);
or U3789 (N_3789,N_3527,N_3319);
xor U3790 (N_3790,N_3375,N_3448);
and U3791 (N_3791,N_3487,N_3456);
nor U3792 (N_3792,N_3429,N_3368);
xor U3793 (N_3793,N_3456,N_3543);
xnor U3794 (N_3794,N_3468,N_3395);
and U3795 (N_3795,N_3508,N_3371);
and U3796 (N_3796,N_3491,N_3487);
and U3797 (N_3797,N_3453,N_3467);
nor U3798 (N_3798,N_3542,N_3584);
or U3799 (N_3799,N_3572,N_3521);
nand U3800 (N_3800,N_3428,N_3589);
xor U3801 (N_3801,N_3483,N_3599);
nand U3802 (N_3802,N_3587,N_3528);
and U3803 (N_3803,N_3520,N_3523);
and U3804 (N_3804,N_3405,N_3351);
nand U3805 (N_3805,N_3508,N_3370);
nor U3806 (N_3806,N_3585,N_3358);
nand U3807 (N_3807,N_3451,N_3456);
nand U3808 (N_3808,N_3580,N_3482);
nand U3809 (N_3809,N_3556,N_3551);
or U3810 (N_3810,N_3574,N_3489);
and U3811 (N_3811,N_3514,N_3326);
or U3812 (N_3812,N_3543,N_3391);
and U3813 (N_3813,N_3429,N_3454);
and U3814 (N_3814,N_3418,N_3489);
or U3815 (N_3815,N_3515,N_3591);
nor U3816 (N_3816,N_3469,N_3304);
nand U3817 (N_3817,N_3394,N_3537);
nand U3818 (N_3818,N_3311,N_3326);
and U3819 (N_3819,N_3339,N_3493);
and U3820 (N_3820,N_3568,N_3554);
xor U3821 (N_3821,N_3513,N_3599);
xor U3822 (N_3822,N_3501,N_3399);
or U3823 (N_3823,N_3411,N_3440);
nand U3824 (N_3824,N_3521,N_3492);
nor U3825 (N_3825,N_3593,N_3448);
and U3826 (N_3826,N_3484,N_3393);
nor U3827 (N_3827,N_3331,N_3500);
nor U3828 (N_3828,N_3569,N_3347);
xor U3829 (N_3829,N_3410,N_3309);
xor U3830 (N_3830,N_3304,N_3531);
xnor U3831 (N_3831,N_3391,N_3337);
nor U3832 (N_3832,N_3334,N_3302);
nor U3833 (N_3833,N_3562,N_3384);
and U3834 (N_3834,N_3581,N_3321);
xnor U3835 (N_3835,N_3414,N_3532);
or U3836 (N_3836,N_3442,N_3416);
nand U3837 (N_3837,N_3437,N_3399);
nor U3838 (N_3838,N_3535,N_3388);
nand U3839 (N_3839,N_3365,N_3322);
and U3840 (N_3840,N_3359,N_3380);
or U3841 (N_3841,N_3408,N_3457);
and U3842 (N_3842,N_3473,N_3408);
and U3843 (N_3843,N_3463,N_3578);
and U3844 (N_3844,N_3438,N_3416);
nor U3845 (N_3845,N_3448,N_3350);
xnor U3846 (N_3846,N_3566,N_3369);
nand U3847 (N_3847,N_3526,N_3330);
xor U3848 (N_3848,N_3432,N_3550);
nand U3849 (N_3849,N_3567,N_3305);
nand U3850 (N_3850,N_3512,N_3448);
nor U3851 (N_3851,N_3505,N_3414);
nor U3852 (N_3852,N_3552,N_3438);
or U3853 (N_3853,N_3404,N_3495);
xor U3854 (N_3854,N_3597,N_3490);
nor U3855 (N_3855,N_3377,N_3322);
and U3856 (N_3856,N_3473,N_3519);
or U3857 (N_3857,N_3519,N_3417);
xnor U3858 (N_3858,N_3407,N_3335);
and U3859 (N_3859,N_3338,N_3507);
nand U3860 (N_3860,N_3452,N_3524);
and U3861 (N_3861,N_3525,N_3363);
nand U3862 (N_3862,N_3514,N_3458);
xor U3863 (N_3863,N_3322,N_3383);
or U3864 (N_3864,N_3488,N_3307);
xnor U3865 (N_3865,N_3451,N_3538);
nand U3866 (N_3866,N_3437,N_3413);
nor U3867 (N_3867,N_3522,N_3366);
and U3868 (N_3868,N_3591,N_3522);
xnor U3869 (N_3869,N_3331,N_3515);
xnor U3870 (N_3870,N_3587,N_3325);
nand U3871 (N_3871,N_3405,N_3503);
nor U3872 (N_3872,N_3425,N_3396);
nand U3873 (N_3873,N_3432,N_3475);
and U3874 (N_3874,N_3352,N_3529);
nand U3875 (N_3875,N_3343,N_3445);
or U3876 (N_3876,N_3456,N_3533);
xnor U3877 (N_3877,N_3443,N_3307);
and U3878 (N_3878,N_3590,N_3491);
nor U3879 (N_3879,N_3405,N_3435);
or U3880 (N_3880,N_3396,N_3321);
nand U3881 (N_3881,N_3340,N_3574);
and U3882 (N_3882,N_3492,N_3404);
nor U3883 (N_3883,N_3527,N_3314);
xnor U3884 (N_3884,N_3447,N_3569);
or U3885 (N_3885,N_3537,N_3310);
or U3886 (N_3886,N_3491,N_3526);
nor U3887 (N_3887,N_3445,N_3439);
nand U3888 (N_3888,N_3440,N_3482);
or U3889 (N_3889,N_3395,N_3444);
nor U3890 (N_3890,N_3541,N_3584);
or U3891 (N_3891,N_3420,N_3590);
or U3892 (N_3892,N_3499,N_3465);
nand U3893 (N_3893,N_3386,N_3371);
and U3894 (N_3894,N_3550,N_3588);
or U3895 (N_3895,N_3311,N_3315);
or U3896 (N_3896,N_3406,N_3328);
xor U3897 (N_3897,N_3504,N_3445);
xnor U3898 (N_3898,N_3300,N_3473);
nor U3899 (N_3899,N_3303,N_3320);
nor U3900 (N_3900,N_3688,N_3789);
and U3901 (N_3901,N_3729,N_3808);
nor U3902 (N_3902,N_3692,N_3604);
and U3903 (N_3903,N_3700,N_3682);
and U3904 (N_3904,N_3823,N_3809);
and U3905 (N_3905,N_3785,N_3765);
and U3906 (N_3906,N_3690,N_3827);
or U3907 (N_3907,N_3640,N_3898);
and U3908 (N_3908,N_3782,N_3891);
xnor U3909 (N_3909,N_3818,N_3728);
xnor U3910 (N_3910,N_3780,N_3821);
or U3911 (N_3911,N_3753,N_3719);
and U3912 (N_3912,N_3831,N_3835);
xnor U3913 (N_3913,N_3703,N_3722);
nor U3914 (N_3914,N_3801,N_3767);
nand U3915 (N_3915,N_3881,N_3899);
nand U3916 (N_3916,N_3736,N_3664);
xnor U3917 (N_3917,N_3704,N_3768);
nor U3918 (N_3918,N_3607,N_3802);
or U3919 (N_3919,N_3796,N_3605);
nor U3920 (N_3920,N_3836,N_3739);
and U3921 (N_3921,N_3819,N_3868);
xnor U3922 (N_3922,N_3877,N_3636);
and U3923 (N_3923,N_3677,N_3631);
and U3924 (N_3924,N_3873,N_3681);
nand U3925 (N_3925,N_3769,N_3861);
or U3926 (N_3926,N_3807,N_3684);
nand U3927 (N_3927,N_3890,N_3689);
nand U3928 (N_3928,N_3754,N_3674);
nand U3929 (N_3929,N_3610,N_3755);
and U3930 (N_3930,N_3752,N_3647);
xnor U3931 (N_3931,N_3745,N_3805);
nor U3932 (N_3932,N_3852,N_3672);
or U3933 (N_3933,N_3601,N_3848);
nand U3934 (N_3934,N_3643,N_3649);
or U3935 (N_3935,N_3683,N_3866);
nor U3936 (N_3936,N_3756,N_3856);
nand U3937 (N_3937,N_3676,N_3661);
or U3938 (N_3938,N_3795,N_3693);
nor U3939 (N_3939,N_3716,N_3616);
and U3940 (N_3940,N_3845,N_3760);
nand U3941 (N_3941,N_3655,N_3670);
or U3942 (N_3942,N_3717,N_3726);
nand U3943 (N_3943,N_3800,N_3824);
nand U3944 (N_3944,N_3849,N_3713);
nand U3945 (N_3945,N_3699,N_3675);
or U3946 (N_3946,N_3758,N_3878);
nand U3947 (N_3947,N_3623,N_3749);
or U3948 (N_3948,N_3740,N_3705);
nor U3949 (N_3949,N_3656,N_3839);
nor U3950 (N_3950,N_3696,N_3666);
nand U3951 (N_3951,N_3872,N_3687);
and U3952 (N_3952,N_3630,N_3641);
nand U3953 (N_3953,N_3686,N_3888);
nand U3954 (N_3954,N_3741,N_3678);
or U3955 (N_3955,N_3615,N_3706);
nand U3956 (N_3956,N_3775,N_3727);
or U3957 (N_3957,N_3709,N_3799);
xnor U3958 (N_3958,N_3712,N_3685);
and U3959 (N_3959,N_3635,N_3810);
nand U3960 (N_3960,N_3762,N_3816);
and U3961 (N_3961,N_3869,N_3733);
or U3962 (N_3962,N_3885,N_3707);
nand U3963 (N_3963,N_3669,N_3847);
or U3964 (N_3964,N_3732,N_3628);
and U3965 (N_3965,N_3642,N_3798);
or U3966 (N_3966,N_3751,N_3659);
nor U3967 (N_3967,N_3855,N_3710);
nor U3968 (N_3968,N_3794,N_3771);
and U3969 (N_3969,N_3668,N_3750);
nand U3970 (N_3970,N_3725,N_3634);
nor U3971 (N_3971,N_3737,N_3608);
xor U3972 (N_3972,N_3777,N_3724);
nand U3973 (N_3973,N_3738,N_3870);
or U3974 (N_3974,N_3862,N_3770);
xor U3975 (N_3975,N_3679,N_3702);
or U3976 (N_3976,N_3886,N_3874);
xnor U3977 (N_3977,N_3639,N_3618);
or U3978 (N_3978,N_3882,N_3804);
nor U3979 (N_3979,N_3781,N_3680);
nor U3980 (N_3980,N_3791,N_3622);
and U3981 (N_3981,N_3654,N_3650);
nand U3982 (N_3982,N_3894,N_3833);
and U3983 (N_3983,N_3746,N_3883);
nor U3984 (N_3984,N_3662,N_3665);
nor U3985 (N_3985,N_3763,N_3853);
xnor U3986 (N_3986,N_3627,N_3834);
nor U3987 (N_3987,N_3837,N_3897);
nand U3988 (N_3988,N_3612,N_3600);
xor U3989 (N_3989,N_3708,N_3730);
nand U3990 (N_3990,N_3854,N_3633);
or U3991 (N_3991,N_3764,N_3875);
xor U3992 (N_3992,N_3609,N_3843);
nand U3993 (N_3993,N_3602,N_3813);
nor U3994 (N_3994,N_3863,N_3851);
xor U3995 (N_3995,N_3896,N_3718);
nand U3996 (N_3996,N_3698,N_3625);
and U3997 (N_3997,N_3773,N_3658);
or U3998 (N_3998,N_3761,N_3820);
or U3999 (N_3999,N_3644,N_3613);
and U4000 (N_4000,N_3734,N_3829);
nor U4001 (N_4001,N_3742,N_3857);
and U4002 (N_4002,N_3695,N_3614);
nand U4003 (N_4003,N_3766,N_3621);
or U4004 (N_4004,N_3840,N_3889);
or U4005 (N_4005,N_3691,N_3606);
and U4006 (N_4006,N_3826,N_3774);
xnor U4007 (N_4007,N_3701,N_3841);
nand U4008 (N_4008,N_3865,N_3822);
or U4009 (N_4009,N_3611,N_3697);
xnor U4010 (N_4010,N_3790,N_3830);
or U4011 (N_4011,N_3792,N_3788);
nand U4012 (N_4012,N_3815,N_3838);
nand U4013 (N_4013,N_3783,N_3757);
nand U4014 (N_4014,N_3603,N_3721);
xnor U4015 (N_4015,N_3620,N_3629);
xor U4016 (N_4016,N_3772,N_3651);
and U4017 (N_4017,N_3787,N_3842);
nand U4018 (N_4018,N_3663,N_3731);
nor U4019 (N_4019,N_3879,N_3779);
nand U4020 (N_4020,N_3653,N_3892);
nor U4021 (N_4021,N_3648,N_3871);
nand U4022 (N_4022,N_3803,N_3652);
or U4023 (N_4023,N_3895,N_3784);
nand U4024 (N_4024,N_3714,N_3844);
nor U4025 (N_4025,N_3748,N_3715);
and U4026 (N_4026,N_3637,N_3846);
or U4027 (N_4027,N_3632,N_3638);
or U4028 (N_4028,N_3832,N_3864);
xnor U4029 (N_4029,N_3626,N_3880);
or U4030 (N_4030,N_3720,N_3850);
nand U4031 (N_4031,N_3776,N_3797);
xnor U4032 (N_4032,N_3884,N_3793);
xor U4033 (N_4033,N_3806,N_3876);
and U4034 (N_4034,N_3747,N_3817);
or U4035 (N_4035,N_3660,N_3811);
or U4036 (N_4036,N_3860,N_3671);
nor U4037 (N_4037,N_3867,N_3858);
nand U4038 (N_4038,N_3859,N_3667);
nor U4039 (N_4039,N_3711,N_3657);
or U4040 (N_4040,N_3619,N_3887);
nor U4041 (N_4041,N_3735,N_3646);
nor U4042 (N_4042,N_3759,N_3778);
or U4043 (N_4043,N_3744,N_3694);
and U4044 (N_4044,N_3673,N_3743);
and U4045 (N_4045,N_3645,N_3825);
nor U4046 (N_4046,N_3814,N_3812);
xnor U4047 (N_4047,N_3624,N_3617);
and U4048 (N_4048,N_3786,N_3828);
nand U4049 (N_4049,N_3723,N_3893);
or U4050 (N_4050,N_3871,N_3686);
and U4051 (N_4051,N_3896,N_3877);
nand U4052 (N_4052,N_3718,N_3684);
nor U4053 (N_4053,N_3630,N_3619);
xnor U4054 (N_4054,N_3823,N_3786);
xor U4055 (N_4055,N_3671,N_3819);
or U4056 (N_4056,N_3707,N_3896);
xor U4057 (N_4057,N_3779,N_3807);
and U4058 (N_4058,N_3838,N_3629);
or U4059 (N_4059,N_3757,N_3606);
nand U4060 (N_4060,N_3757,N_3822);
xnor U4061 (N_4061,N_3713,N_3828);
nand U4062 (N_4062,N_3827,N_3741);
nand U4063 (N_4063,N_3680,N_3630);
xnor U4064 (N_4064,N_3717,N_3631);
nand U4065 (N_4065,N_3811,N_3894);
or U4066 (N_4066,N_3651,N_3773);
and U4067 (N_4067,N_3745,N_3602);
or U4068 (N_4068,N_3727,N_3897);
or U4069 (N_4069,N_3839,N_3604);
nor U4070 (N_4070,N_3840,N_3729);
xnor U4071 (N_4071,N_3818,N_3698);
xnor U4072 (N_4072,N_3730,N_3697);
or U4073 (N_4073,N_3604,N_3695);
and U4074 (N_4074,N_3737,N_3889);
nor U4075 (N_4075,N_3677,N_3862);
or U4076 (N_4076,N_3715,N_3710);
or U4077 (N_4077,N_3836,N_3817);
nand U4078 (N_4078,N_3862,N_3805);
nor U4079 (N_4079,N_3773,N_3638);
and U4080 (N_4080,N_3736,N_3743);
or U4081 (N_4081,N_3683,N_3637);
nand U4082 (N_4082,N_3843,N_3776);
nand U4083 (N_4083,N_3631,N_3655);
xor U4084 (N_4084,N_3699,N_3739);
nor U4085 (N_4085,N_3835,N_3781);
and U4086 (N_4086,N_3709,N_3801);
and U4087 (N_4087,N_3715,N_3786);
or U4088 (N_4088,N_3750,N_3858);
and U4089 (N_4089,N_3812,N_3826);
nor U4090 (N_4090,N_3656,N_3810);
or U4091 (N_4091,N_3600,N_3701);
xnor U4092 (N_4092,N_3760,N_3727);
xnor U4093 (N_4093,N_3887,N_3800);
and U4094 (N_4094,N_3855,N_3870);
nand U4095 (N_4095,N_3618,N_3700);
xor U4096 (N_4096,N_3605,N_3857);
xnor U4097 (N_4097,N_3671,N_3667);
nand U4098 (N_4098,N_3869,N_3710);
or U4099 (N_4099,N_3883,N_3676);
nor U4100 (N_4100,N_3796,N_3839);
nand U4101 (N_4101,N_3778,N_3729);
nor U4102 (N_4102,N_3707,N_3631);
and U4103 (N_4103,N_3864,N_3604);
xnor U4104 (N_4104,N_3656,N_3859);
xnor U4105 (N_4105,N_3772,N_3791);
nor U4106 (N_4106,N_3828,N_3659);
nand U4107 (N_4107,N_3746,N_3608);
and U4108 (N_4108,N_3728,N_3636);
and U4109 (N_4109,N_3810,N_3791);
nand U4110 (N_4110,N_3710,N_3674);
or U4111 (N_4111,N_3682,N_3727);
or U4112 (N_4112,N_3862,N_3606);
and U4113 (N_4113,N_3672,N_3761);
nand U4114 (N_4114,N_3830,N_3677);
nand U4115 (N_4115,N_3736,N_3831);
nor U4116 (N_4116,N_3694,N_3658);
nand U4117 (N_4117,N_3603,N_3606);
and U4118 (N_4118,N_3815,N_3858);
nand U4119 (N_4119,N_3690,N_3720);
nor U4120 (N_4120,N_3619,N_3792);
or U4121 (N_4121,N_3875,N_3892);
nor U4122 (N_4122,N_3870,N_3785);
and U4123 (N_4123,N_3687,N_3885);
nand U4124 (N_4124,N_3638,N_3791);
xor U4125 (N_4125,N_3773,N_3852);
or U4126 (N_4126,N_3746,N_3838);
or U4127 (N_4127,N_3717,N_3708);
nor U4128 (N_4128,N_3725,N_3637);
nor U4129 (N_4129,N_3618,N_3656);
xnor U4130 (N_4130,N_3616,N_3612);
or U4131 (N_4131,N_3643,N_3777);
nor U4132 (N_4132,N_3810,N_3737);
nor U4133 (N_4133,N_3628,N_3830);
nand U4134 (N_4134,N_3881,N_3880);
nor U4135 (N_4135,N_3623,N_3607);
or U4136 (N_4136,N_3777,N_3877);
or U4137 (N_4137,N_3791,N_3876);
and U4138 (N_4138,N_3615,N_3760);
or U4139 (N_4139,N_3757,N_3713);
xor U4140 (N_4140,N_3896,N_3674);
nand U4141 (N_4141,N_3676,N_3644);
nand U4142 (N_4142,N_3812,N_3868);
xnor U4143 (N_4143,N_3680,N_3642);
and U4144 (N_4144,N_3601,N_3807);
and U4145 (N_4145,N_3829,N_3816);
and U4146 (N_4146,N_3643,N_3884);
nand U4147 (N_4147,N_3818,N_3766);
or U4148 (N_4148,N_3704,N_3627);
nand U4149 (N_4149,N_3794,N_3686);
xor U4150 (N_4150,N_3747,N_3664);
nand U4151 (N_4151,N_3798,N_3646);
nor U4152 (N_4152,N_3872,N_3714);
and U4153 (N_4153,N_3820,N_3610);
and U4154 (N_4154,N_3639,N_3854);
xor U4155 (N_4155,N_3612,N_3640);
or U4156 (N_4156,N_3627,N_3774);
xnor U4157 (N_4157,N_3765,N_3767);
xor U4158 (N_4158,N_3717,N_3636);
xnor U4159 (N_4159,N_3753,N_3846);
xor U4160 (N_4160,N_3633,N_3756);
xnor U4161 (N_4161,N_3698,N_3844);
or U4162 (N_4162,N_3616,N_3831);
xnor U4163 (N_4163,N_3814,N_3716);
or U4164 (N_4164,N_3863,N_3797);
or U4165 (N_4165,N_3746,N_3784);
xor U4166 (N_4166,N_3643,N_3754);
and U4167 (N_4167,N_3872,N_3729);
nand U4168 (N_4168,N_3690,N_3751);
and U4169 (N_4169,N_3732,N_3690);
xnor U4170 (N_4170,N_3805,N_3815);
or U4171 (N_4171,N_3689,N_3869);
nor U4172 (N_4172,N_3689,N_3785);
nor U4173 (N_4173,N_3875,N_3773);
or U4174 (N_4174,N_3662,N_3890);
and U4175 (N_4175,N_3703,N_3602);
and U4176 (N_4176,N_3722,N_3606);
or U4177 (N_4177,N_3778,N_3754);
nor U4178 (N_4178,N_3857,N_3712);
nor U4179 (N_4179,N_3825,N_3799);
and U4180 (N_4180,N_3618,N_3657);
xor U4181 (N_4181,N_3794,N_3692);
nor U4182 (N_4182,N_3665,N_3848);
or U4183 (N_4183,N_3763,N_3816);
and U4184 (N_4184,N_3757,N_3726);
xnor U4185 (N_4185,N_3852,N_3848);
or U4186 (N_4186,N_3745,N_3831);
nand U4187 (N_4187,N_3626,N_3887);
or U4188 (N_4188,N_3637,N_3771);
nand U4189 (N_4189,N_3776,N_3702);
or U4190 (N_4190,N_3622,N_3893);
xor U4191 (N_4191,N_3774,N_3789);
xor U4192 (N_4192,N_3693,N_3629);
nor U4193 (N_4193,N_3757,N_3861);
or U4194 (N_4194,N_3639,N_3667);
xnor U4195 (N_4195,N_3682,N_3694);
nand U4196 (N_4196,N_3715,N_3881);
nand U4197 (N_4197,N_3642,N_3723);
and U4198 (N_4198,N_3703,N_3823);
and U4199 (N_4199,N_3811,N_3879);
or U4200 (N_4200,N_4189,N_3900);
and U4201 (N_4201,N_3960,N_3905);
nand U4202 (N_4202,N_3970,N_3926);
nand U4203 (N_4203,N_4067,N_4044);
xor U4204 (N_4204,N_4159,N_3990);
nand U4205 (N_4205,N_4151,N_4045);
nor U4206 (N_4206,N_4177,N_4007);
nor U4207 (N_4207,N_3993,N_4180);
and U4208 (N_4208,N_4173,N_4131);
xnor U4209 (N_4209,N_3918,N_4136);
and U4210 (N_4210,N_4008,N_4005);
nor U4211 (N_4211,N_4119,N_4124);
or U4212 (N_4212,N_3951,N_4167);
nor U4213 (N_4213,N_4192,N_3985);
xnor U4214 (N_4214,N_4006,N_4101);
xnor U4215 (N_4215,N_4077,N_4087);
and U4216 (N_4216,N_3991,N_4036);
nand U4217 (N_4217,N_3929,N_4175);
nor U4218 (N_4218,N_4051,N_4010);
nand U4219 (N_4219,N_3923,N_3925);
xnor U4220 (N_4220,N_4085,N_4161);
nand U4221 (N_4221,N_4066,N_4086);
xor U4222 (N_4222,N_4137,N_4133);
nor U4223 (N_4223,N_4164,N_3975);
nor U4224 (N_4224,N_4171,N_4011);
or U4225 (N_4225,N_3984,N_3971);
nand U4226 (N_4226,N_4021,N_4163);
xnor U4227 (N_4227,N_3955,N_3999);
xor U4228 (N_4228,N_4039,N_4146);
or U4229 (N_4229,N_3921,N_4110);
nor U4230 (N_4230,N_4182,N_4153);
nor U4231 (N_4231,N_4156,N_3964);
and U4232 (N_4232,N_4083,N_4048);
nand U4233 (N_4233,N_3978,N_3908);
nor U4234 (N_4234,N_4114,N_4075);
nor U4235 (N_4235,N_3930,N_4185);
nand U4236 (N_4236,N_4025,N_4097);
xor U4237 (N_4237,N_4014,N_4070);
or U4238 (N_4238,N_4040,N_4091);
nor U4239 (N_4239,N_3915,N_4043);
nor U4240 (N_4240,N_4191,N_3924);
nor U4241 (N_4241,N_4009,N_4024);
or U4242 (N_4242,N_4084,N_3947);
nand U4243 (N_4243,N_4176,N_4018);
or U4244 (N_4244,N_4138,N_4093);
and U4245 (N_4245,N_4130,N_4116);
or U4246 (N_4246,N_4169,N_3974);
xnor U4247 (N_4247,N_3997,N_4035);
xnor U4248 (N_4248,N_4029,N_3953);
and U4249 (N_4249,N_3934,N_4172);
and U4250 (N_4250,N_4057,N_3945);
nand U4251 (N_4251,N_3994,N_4072);
xor U4252 (N_4252,N_3901,N_4170);
nor U4253 (N_4253,N_4198,N_4199);
nand U4254 (N_4254,N_4019,N_4115);
and U4255 (N_4255,N_4060,N_4111);
xor U4256 (N_4256,N_4068,N_3943);
or U4257 (N_4257,N_4183,N_3907);
nor U4258 (N_4258,N_4184,N_4129);
xnor U4259 (N_4259,N_3961,N_4113);
and U4260 (N_4260,N_4100,N_4122);
and U4261 (N_4261,N_4166,N_3942);
nor U4262 (N_4262,N_4046,N_3928);
or U4263 (N_4263,N_4152,N_3957);
or U4264 (N_4264,N_3962,N_4052);
xnor U4265 (N_4265,N_3988,N_3948);
or U4266 (N_4266,N_4094,N_4090);
nand U4267 (N_4267,N_3940,N_4076);
xor U4268 (N_4268,N_4160,N_3956);
nand U4269 (N_4269,N_3916,N_3912);
nor U4270 (N_4270,N_3932,N_4098);
nor U4271 (N_4271,N_3949,N_4117);
or U4272 (N_4272,N_4125,N_4031);
xnor U4273 (N_4273,N_4079,N_3938);
or U4274 (N_4274,N_4030,N_4142);
nand U4275 (N_4275,N_4178,N_4012);
or U4276 (N_4276,N_3914,N_4132);
nor U4277 (N_4277,N_3910,N_4179);
xor U4278 (N_4278,N_3906,N_4104);
nor U4279 (N_4279,N_4108,N_3936);
nand U4280 (N_4280,N_3981,N_4181);
nand U4281 (N_4281,N_3941,N_4069);
xnor U4282 (N_4282,N_4154,N_3950);
nor U4283 (N_4283,N_4095,N_4054);
nand U4284 (N_4284,N_4073,N_4121);
xnor U4285 (N_4285,N_4027,N_3902);
nor U4286 (N_4286,N_3920,N_3944);
nor U4287 (N_4287,N_4033,N_4127);
or U4288 (N_4288,N_4001,N_4059);
nand U4289 (N_4289,N_4174,N_4107);
and U4290 (N_4290,N_3927,N_3986);
nor U4291 (N_4291,N_3967,N_3989);
xnor U4292 (N_4292,N_4096,N_4034);
xnor U4293 (N_4293,N_4081,N_3939);
or U4294 (N_4294,N_3954,N_4058);
xnor U4295 (N_4295,N_4015,N_4193);
nand U4296 (N_4296,N_4080,N_4135);
or U4297 (N_4297,N_4053,N_4150);
nand U4298 (N_4298,N_4112,N_4020);
nor U4299 (N_4299,N_4162,N_4141);
nand U4300 (N_4300,N_4158,N_4186);
and U4301 (N_4301,N_3996,N_4064);
nand U4302 (N_4302,N_3913,N_4194);
nor U4303 (N_4303,N_4013,N_3917);
nor U4304 (N_4304,N_3968,N_4140);
nor U4305 (N_4305,N_4099,N_4088);
and U4306 (N_4306,N_3937,N_4197);
and U4307 (N_4307,N_3965,N_3980);
nand U4308 (N_4308,N_4055,N_4061);
or U4309 (N_4309,N_4089,N_4165);
nand U4310 (N_4310,N_4139,N_4118);
or U4311 (N_4311,N_4004,N_3979);
nor U4312 (N_4312,N_3909,N_4047);
or U4313 (N_4313,N_3977,N_4023);
nor U4314 (N_4314,N_3966,N_4003);
and U4315 (N_4315,N_4128,N_4032);
and U4316 (N_4316,N_3987,N_4126);
and U4317 (N_4317,N_4105,N_4196);
or U4318 (N_4318,N_4148,N_4078);
nor U4319 (N_4319,N_4149,N_4017);
or U4320 (N_4320,N_3998,N_4016);
xor U4321 (N_4321,N_3976,N_3933);
xor U4322 (N_4322,N_4155,N_4050);
or U4323 (N_4323,N_4049,N_4103);
nand U4324 (N_4324,N_3952,N_3922);
and U4325 (N_4325,N_4071,N_4028);
nor U4326 (N_4326,N_4145,N_4062);
nand U4327 (N_4327,N_4092,N_3946);
or U4328 (N_4328,N_3982,N_4123);
xor U4329 (N_4329,N_4022,N_4134);
nand U4330 (N_4330,N_3983,N_4026);
and U4331 (N_4331,N_4109,N_4037);
and U4332 (N_4332,N_4065,N_4002);
or U4333 (N_4333,N_4144,N_3919);
xnor U4334 (N_4334,N_4195,N_3903);
nand U4335 (N_4335,N_3931,N_3958);
or U4336 (N_4336,N_3959,N_4102);
and U4337 (N_4337,N_4190,N_4168);
xnor U4338 (N_4338,N_4038,N_3969);
xnor U4339 (N_4339,N_4147,N_4120);
and U4340 (N_4340,N_3992,N_4143);
nand U4341 (N_4341,N_4000,N_3904);
nor U4342 (N_4342,N_4056,N_4042);
xor U4343 (N_4343,N_4188,N_4074);
nor U4344 (N_4344,N_3911,N_4106);
or U4345 (N_4345,N_4187,N_3973);
and U4346 (N_4346,N_4082,N_4063);
nand U4347 (N_4347,N_3935,N_3972);
and U4348 (N_4348,N_4157,N_3995);
xnor U4349 (N_4349,N_3963,N_4041);
nand U4350 (N_4350,N_4092,N_4041);
nor U4351 (N_4351,N_4025,N_4006);
nand U4352 (N_4352,N_3949,N_3933);
or U4353 (N_4353,N_3963,N_3980);
and U4354 (N_4354,N_4046,N_4111);
nor U4355 (N_4355,N_4124,N_3997);
and U4356 (N_4356,N_4081,N_4009);
or U4357 (N_4357,N_4033,N_4195);
nor U4358 (N_4358,N_3945,N_4101);
nor U4359 (N_4359,N_4092,N_3990);
xnor U4360 (N_4360,N_4103,N_3968);
xor U4361 (N_4361,N_4009,N_4069);
nand U4362 (N_4362,N_4154,N_4195);
or U4363 (N_4363,N_4028,N_3977);
nand U4364 (N_4364,N_4125,N_4091);
or U4365 (N_4365,N_3940,N_4117);
and U4366 (N_4366,N_3979,N_3971);
xor U4367 (N_4367,N_4046,N_4162);
nor U4368 (N_4368,N_4046,N_3923);
nand U4369 (N_4369,N_4153,N_3955);
xnor U4370 (N_4370,N_3970,N_4199);
or U4371 (N_4371,N_4059,N_4149);
nand U4372 (N_4372,N_4047,N_4016);
or U4373 (N_4373,N_3950,N_4158);
nor U4374 (N_4374,N_3900,N_4033);
nand U4375 (N_4375,N_4019,N_3926);
and U4376 (N_4376,N_3902,N_4034);
or U4377 (N_4377,N_4021,N_3900);
and U4378 (N_4378,N_4033,N_4091);
and U4379 (N_4379,N_3953,N_3986);
and U4380 (N_4380,N_4131,N_4137);
xor U4381 (N_4381,N_4155,N_3950);
or U4382 (N_4382,N_3973,N_4106);
or U4383 (N_4383,N_3945,N_4082);
or U4384 (N_4384,N_4119,N_4170);
nand U4385 (N_4385,N_3908,N_4173);
nand U4386 (N_4386,N_3969,N_4152);
xor U4387 (N_4387,N_4121,N_4174);
and U4388 (N_4388,N_4123,N_4139);
xnor U4389 (N_4389,N_4068,N_4120);
or U4390 (N_4390,N_3951,N_4189);
or U4391 (N_4391,N_4053,N_3977);
and U4392 (N_4392,N_4025,N_4041);
nand U4393 (N_4393,N_4193,N_4104);
or U4394 (N_4394,N_3998,N_4061);
or U4395 (N_4395,N_4056,N_4069);
xnor U4396 (N_4396,N_4115,N_4042);
or U4397 (N_4397,N_4120,N_4054);
xor U4398 (N_4398,N_4144,N_4149);
and U4399 (N_4399,N_4114,N_4006);
nand U4400 (N_4400,N_3949,N_4052);
and U4401 (N_4401,N_4068,N_4114);
or U4402 (N_4402,N_3980,N_4167);
or U4403 (N_4403,N_4084,N_4116);
or U4404 (N_4404,N_4098,N_3921);
nor U4405 (N_4405,N_4048,N_4187);
nand U4406 (N_4406,N_4074,N_4133);
nand U4407 (N_4407,N_3930,N_4039);
xor U4408 (N_4408,N_4151,N_3982);
or U4409 (N_4409,N_4067,N_4121);
xnor U4410 (N_4410,N_4169,N_3952);
nor U4411 (N_4411,N_4199,N_3919);
xor U4412 (N_4412,N_4147,N_3999);
nor U4413 (N_4413,N_4135,N_4057);
or U4414 (N_4414,N_3901,N_3903);
xor U4415 (N_4415,N_4054,N_4145);
nand U4416 (N_4416,N_4000,N_4135);
nor U4417 (N_4417,N_4023,N_4160);
and U4418 (N_4418,N_3990,N_3968);
xor U4419 (N_4419,N_4044,N_4003);
nand U4420 (N_4420,N_4076,N_4182);
xnor U4421 (N_4421,N_4153,N_4058);
or U4422 (N_4422,N_4133,N_4145);
nand U4423 (N_4423,N_3916,N_3933);
or U4424 (N_4424,N_4068,N_4184);
and U4425 (N_4425,N_4049,N_4151);
xnor U4426 (N_4426,N_3946,N_4082);
nor U4427 (N_4427,N_4019,N_4180);
xor U4428 (N_4428,N_3960,N_3943);
nor U4429 (N_4429,N_4089,N_4030);
or U4430 (N_4430,N_3952,N_3962);
or U4431 (N_4431,N_4054,N_4169);
and U4432 (N_4432,N_4162,N_3970);
nand U4433 (N_4433,N_3959,N_4004);
and U4434 (N_4434,N_4047,N_4072);
and U4435 (N_4435,N_4123,N_4017);
nor U4436 (N_4436,N_4146,N_4157);
xnor U4437 (N_4437,N_4058,N_3961);
nor U4438 (N_4438,N_3969,N_4079);
or U4439 (N_4439,N_3919,N_4074);
xnor U4440 (N_4440,N_3956,N_4019);
or U4441 (N_4441,N_4128,N_3901);
nand U4442 (N_4442,N_4048,N_4060);
nor U4443 (N_4443,N_4032,N_3909);
xnor U4444 (N_4444,N_4110,N_4003);
or U4445 (N_4445,N_4007,N_3976);
and U4446 (N_4446,N_3970,N_4025);
nand U4447 (N_4447,N_4077,N_4076);
nand U4448 (N_4448,N_4141,N_3992);
nand U4449 (N_4449,N_3939,N_4097);
or U4450 (N_4450,N_4131,N_3963);
or U4451 (N_4451,N_3946,N_4149);
nor U4452 (N_4452,N_4064,N_4103);
xor U4453 (N_4453,N_4105,N_4143);
xnor U4454 (N_4454,N_4017,N_3966);
nand U4455 (N_4455,N_3920,N_4062);
xor U4456 (N_4456,N_4176,N_4024);
nand U4457 (N_4457,N_3996,N_3995);
nor U4458 (N_4458,N_4051,N_4060);
nor U4459 (N_4459,N_4026,N_3959);
nand U4460 (N_4460,N_4073,N_4134);
or U4461 (N_4461,N_4029,N_4062);
nand U4462 (N_4462,N_3907,N_3979);
nor U4463 (N_4463,N_4159,N_4181);
or U4464 (N_4464,N_4127,N_4134);
or U4465 (N_4465,N_3984,N_3995);
or U4466 (N_4466,N_4118,N_4147);
nand U4467 (N_4467,N_4177,N_3950);
or U4468 (N_4468,N_4094,N_3918);
xnor U4469 (N_4469,N_4069,N_4187);
or U4470 (N_4470,N_3932,N_4095);
nor U4471 (N_4471,N_4191,N_3916);
or U4472 (N_4472,N_4042,N_4118);
or U4473 (N_4473,N_4123,N_3948);
nor U4474 (N_4474,N_4063,N_4118);
xnor U4475 (N_4475,N_3912,N_4175);
xor U4476 (N_4476,N_3996,N_4008);
xnor U4477 (N_4477,N_4070,N_3900);
xor U4478 (N_4478,N_4078,N_4015);
nor U4479 (N_4479,N_3909,N_4173);
xnor U4480 (N_4480,N_4008,N_3990);
nor U4481 (N_4481,N_4000,N_4078);
nand U4482 (N_4482,N_4138,N_3977);
and U4483 (N_4483,N_4051,N_4077);
or U4484 (N_4484,N_4032,N_4077);
nor U4485 (N_4485,N_3996,N_4146);
or U4486 (N_4486,N_4193,N_4108);
and U4487 (N_4487,N_4161,N_4142);
or U4488 (N_4488,N_3983,N_4123);
nor U4489 (N_4489,N_4116,N_4128);
or U4490 (N_4490,N_4096,N_4036);
and U4491 (N_4491,N_4152,N_4120);
xor U4492 (N_4492,N_4138,N_3900);
xor U4493 (N_4493,N_4110,N_3962);
and U4494 (N_4494,N_4138,N_3948);
and U4495 (N_4495,N_4128,N_4167);
xor U4496 (N_4496,N_4039,N_4153);
and U4497 (N_4497,N_3931,N_3992);
nor U4498 (N_4498,N_4170,N_4116);
or U4499 (N_4499,N_4045,N_4009);
and U4500 (N_4500,N_4349,N_4317);
nand U4501 (N_4501,N_4210,N_4437);
nand U4502 (N_4502,N_4448,N_4270);
or U4503 (N_4503,N_4353,N_4362);
xor U4504 (N_4504,N_4346,N_4465);
or U4505 (N_4505,N_4286,N_4466);
nor U4506 (N_4506,N_4388,N_4406);
xnor U4507 (N_4507,N_4201,N_4408);
nand U4508 (N_4508,N_4397,N_4398);
xnor U4509 (N_4509,N_4477,N_4416);
or U4510 (N_4510,N_4499,N_4381);
or U4511 (N_4511,N_4288,N_4219);
nor U4512 (N_4512,N_4402,N_4314);
xor U4513 (N_4513,N_4495,N_4231);
nand U4514 (N_4514,N_4269,N_4470);
or U4515 (N_4515,N_4464,N_4217);
and U4516 (N_4516,N_4278,N_4358);
or U4517 (N_4517,N_4438,N_4232);
xnor U4518 (N_4518,N_4257,N_4453);
nor U4519 (N_4519,N_4379,N_4469);
nand U4520 (N_4520,N_4423,N_4338);
and U4521 (N_4521,N_4372,N_4213);
or U4522 (N_4522,N_4235,N_4376);
nand U4523 (N_4523,N_4445,N_4229);
nor U4524 (N_4524,N_4485,N_4432);
and U4525 (N_4525,N_4289,N_4369);
xnor U4526 (N_4526,N_4242,N_4394);
and U4527 (N_4527,N_4295,N_4204);
xor U4528 (N_4528,N_4370,N_4413);
nand U4529 (N_4529,N_4458,N_4220);
nand U4530 (N_4530,N_4391,N_4202);
xor U4531 (N_4531,N_4247,N_4396);
xnor U4532 (N_4532,N_4365,N_4233);
xor U4533 (N_4533,N_4375,N_4313);
xor U4534 (N_4534,N_4225,N_4491);
or U4535 (N_4535,N_4303,N_4252);
or U4536 (N_4536,N_4393,N_4296);
xor U4537 (N_4537,N_4319,N_4431);
or U4538 (N_4538,N_4290,N_4246);
or U4539 (N_4539,N_4266,N_4254);
nand U4540 (N_4540,N_4449,N_4251);
nor U4541 (N_4541,N_4417,N_4294);
and U4542 (N_4542,N_4366,N_4447);
nor U4543 (N_4543,N_4227,N_4320);
nor U4544 (N_4544,N_4335,N_4304);
nand U4545 (N_4545,N_4498,N_4253);
or U4546 (N_4546,N_4436,N_4331);
nand U4547 (N_4547,N_4236,N_4421);
or U4548 (N_4548,N_4307,N_4308);
xnor U4549 (N_4549,N_4218,N_4324);
or U4550 (N_4550,N_4214,N_4390);
nor U4551 (N_4551,N_4336,N_4240);
nor U4552 (N_4552,N_4250,N_4378);
nand U4553 (N_4553,N_4333,N_4420);
xnor U4554 (N_4554,N_4260,N_4476);
and U4555 (N_4555,N_4442,N_4279);
nand U4556 (N_4556,N_4244,N_4483);
nand U4557 (N_4557,N_4482,N_4262);
nor U4558 (N_4558,N_4481,N_4435);
or U4559 (N_4559,N_4332,N_4454);
nand U4560 (N_4560,N_4385,N_4387);
xor U4561 (N_4561,N_4404,N_4328);
and U4562 (N_4562,N_4441,N_4329);
nor U4563 (N_4563,N_4216,N_4321);
nand U4564 (N_4564,N_4439,N_4340);
nand U4565 (N_4565,N_4489,N_4215);
or U4566 (N_4566,N_4367,N_4249);
nor U4567 (N_4567,N_4209,N_4348);
nand U4568 (N_4568,N_4461,N_4486);
nand U4569 (N_4569,N_4228,N_4463);
nor U4570 (N_4570,N_4323,N_4274);
and U4571 (N_4571,N_4206,N_4357);
nand U4572 (N_4572,N_4405,N_4356);
nor U4573 (N_4573,N_4468,N_4427);
nor U4574 (N_4574,N_4273,N_4345);
xor U4575 (N_4575,N_4203,N_4230);
xnor U4576 (N_4576,N_4237,N_4277);
or U4577 (N_4577,N_4309,N_4223);
and U4578 (N_4578,N_4315,N_4351);
nand U4579 (N_4579,N_4280,N_4239);
nand U4580 (N_4580,N_4424,N_4205);
nand U4581 (N_4581,N_4272,N_4327);
and U4582 (N_4582,N_4440,N_4342);
nand U4583 (N_4583,N_4292,N_4462);
nor U4584 (N_4584,N_4455,N_4467);
or U4585 (N_4585,N_4271,N_4374);
or U4586 (N_4586,N_4222,N_4316);
nand U4587 (N_4587,N_4446,N_4281);
and U4588 (N_4588,N_4415,N_4389);
nor U4589 (N_4589,N_4382,N_4259);
or U4590 (N_4590,N_4429,N_4474);
and U4591 (N_4591,N_4419,N_4494);
nand U4592 (N_4592,N_4359,N_4282);
xor U4593 (N_4593,N_4291,N_4268);
xnor U4594 (N_4594,N_4301,N_4409);
or U4595 (N_4595,N_4311,N_4361);
or U4596 (N_4596,N_4243,N_4487);
nand U4597 (N_4597,N_4241,N_4371);
nand U4598 (N_4598,N_4302,N_4380);
nand U4599 (N_4599,N_4444,N_4299);
and U4600 (N_4600,N_4399,N_4245);
nand U4601 (N_4601,N_4330,N_4403);
and U4602 (N_4602,N_4414,N_4347);
xor U4603 (N_4603,N_4322,N_4407);
and U4604 (N_4604,N_4212,N_4395);
nor U4605 (N_4605,N_4377,N_4422);
nor U4606 (N_4606,N_4451,N_4276);
nand U4607 (N_4607,N_4488,N_4472);
or U4608 (N_4608,N_4256,N_4460);
nor U4609 (N_4609,N_4425,N_4350);
or U4610 (N_4610,N_4384,N_4200);
xnor U4611 (N_4611,N_4298,N_4392);
or U4612 (N_4612,N_4263,N_4265);
or U4613 (N_4613,N_4343,N_4261);
xor U4614 (N_4614,N_4368,N_4471);
or U4615 (N_4615,N_4312,N_4211);
xnor U4616 (N_4616,N_4300,N_4339);
nor U4617 (N_4617,N_4267,N_4492);
nor U4618 (N_4618,N_4479,N_4293);
or U4619 (N_4619,N_4373,N_4264);
nor U4620 (N_4620,N_4360,N_4484);
nor U4621 (N_4621,N_4310,N_4426);
xnor U4622 (N_4622,N_4341,N_4475);
nand U4623 (N_4623,N_4285,N_4283);
or U4624 (N_4624,N_4412,N_4255);
nand U4625 (N_4625,N_4354,N_4430);
xor U4626 (N_4626,N_4355,N_4496);
or U4627 (N_4627,N_4208,N_4493);
and U4628 (N_4628,N_4364,N_4410);
and U4629 (N_4629,N_4411,N_4337);
nand U4630 (N_4630,N_4401,N_4480);
and U4631 (N_4631,N_4287,N_4248);
nor U4632 (N_4632,N_4318,N_4306);
nor U4633 (N_4633,N_4418,N_4234);
nand U4634 (N_4634,N_4383,N_4326);
nand U4635 (N_4635,N_4325,N_4497);
and U4636 (N_4636,N_4452,N_4443);
or U4637 (N_4637,N_4352,N_4297);
nand U4638 (N_4638,N_4457,N_4226);
nand U4639 (N_4639,N_4275,N_4478);
xnor U4640 (N_4640,N_4428,N_4334);
and U4641 (N_4641,N_4459,N_4386);
xnor U4642 (N_4642,N_4434,N_4433);
or U4643 (N_4643,N_4258,N_4284);
nor U4644 (N_4644,N_4238,N_4473);
nor U4645 (N_4645,N_4456,N_4344);
xor U4646 (N_4646,N_4224,N_4207);
or U4647 (N_4647,N_4490,N_4450);
nand U4648 (N_4648,N_4363,N_4221);
xnor U4649 (N_4649,N_4305,N_4400);
or U4650 (N_4650,N_4272,N_4353);
nand U4651 (N_4651,N_4487,N_4278);
and U4652 (N_4652,N_4485,N_4203);
nor U4653 (N_4653,N_4251,N_4398);
nor U4654 (N_4654,N_4484,N_4393);
nand U4655 (N_4655,N_4321,N_4247);
or U4656 (N_4656,N_4482,N_4236);
or U4657 (N_4657,N_4493,N_4235);
nor U4658 (N_4658,N_4288,N_4313);
nor U4659 (N_4659,N_4325,N_4248);
or U4660 (N_4660,N_4245,N_4230);
and U4661 (N_4661,N_4277,N_4391);
and U4662 (N_4662,N_4276,N_4490);
xnor U4663 (N_4663,N_4449,N_4294);
nor U4664 (N_4664,N_4401,N_4263);
nor U4665 (N_4665,N_4246,N_4237);
xnor U4666 (N_4666,N_4338,N_4389);
or U4667 (N_4667,N_4356,N_4439);
xnor U4668 (N_4668,N_4363,N_4436);
xor U4669 (N_4669,N_4408,N_4245);
nor U4670 (N_4670,N_4457,N_4246);
xor U4671 (N_4671,N_4209,N_4358);
nand U4672 (N_4672,N_4249,N_4486);
or U4673 (N_4673,N_4490,N_4473);
and U4674 (N_4674,N_4478,N_4394);
or U4675 (N_4675,N_4271,N_4203);
or U4676 (N_4676,N_4338,N_4473);
and U4677 (N_4677,N_4400,N_4231);
xnor U4678 (N_4678,N_4370,N_4215);
nand U4679 (N_4679,N_4381,N_4403);
and U4680 (N_4680,N_4350,N_4479);
nor U4681 (N_4681,N_4321,N_4463);
xor U4682 (N_4682,N_4407,N_4221);
xor U4683 (N_4683,N_4379,N_4344);
and U4684 (N_4684,N_4295,N_4480);
nand U4685 (N_4685,N_4431,N_4497);
nor U4686 (N_4686,N_4437,N_4263);
nor U4687 (N_4687,N_4436,N_4361);
xnor U4688 (N_4688,N_4496,N_4464);
nand U4689 (N_4689,N_4206,N_4398);
xor U4690 (N_4690,N_4227,N_4375);
nand U4691 (N_4691,N_4342,N_4470);
nor U4692 (N_4692,N_4344,N_4349);
nand U4693 (N_4693,N_4479,N_4307);
nor U4694 (N_4694,N_4285,N_4493);
nand U4695 (N_4695,N_4449,N_4205);
and U4696 (N_4696,N_4463,N_4279);
and U4697 (N_4697,N_4205,N_4277);
and U4698 (N_4698,N_4203,N_4293);
xor U4699 (N_4699,N_4363,N_4451);
xor U4700 (N_4700,N_4496,N_4330);
nand U4701 (N_4701,N_4452,N_4471);
nand U4702 (N_4702,N_4461,N_4237);
nand U4703 (N_4703,N_4220,N_4474);
xor U4704 (N_4704,N_4478,N_4241);
or U4705 (N_4705,N_4367,N_4498);
and U4706 (N_4706,N_4269,N_4396);
xnor U4707 (N_4707,N_4392,N_4289);
nand U4708 (N_4708,N_4230,N_4249);
nand U4709 (N_4709,N_4339,N_4465);
xor U4710 (N_4710,N_4491,N_4299);
and U4711 (N_4711,N_4278,N_4415);
and U4712 (N_4712,N_4429,N_4257);
nand U4713 (N_4713,N_4236,N_4386);
and U4714 (N_4714,N_4228,N_4222);
xor U4715 (N_4715,N_4495,N_4403);
or U4716 (N_4716,N_4281,N_4375);
and U4717 (N_4717,N_4357,N_4236);
or U4718 (N_4718,N_4282,N_4294);
nand U4719 (N_4719,N_4320,N_4455);
nor U4720 (N_4720,N_4222,N_4342);
nand U4721 (N_4721,N_4253,N_4370);
or U4722 (N_4722,N_4208,N_4443);
or U4723 (N_4723,N_4331,N_4429);
nand U4724 (N_4724,N_4382,N_4294);
and U4725 (N_4725,N_4439,N_4278);
xor U4726 (N_4726,N_4474,N_4418);
nand U4727 (N_4727,N_4393,N_4357);
nor U4728 (N_4728,N_4313,N_4404);
and U4729 (N_4729,N_4240,N_4241);
and U4730 (N_4730,N_4427,N_4444);
and U4731 (N_4731,N_4246,N_4247);
and U4732 (N_4732,N_4362,N_4324);
xor U4733 (N_4733,N_4296,N_4276);
nand U4734 (N_4734,N_4432,N_4311);
xor U4735 (N_4735,N_4487,N_4234);
or U4736 (N_4736,N_4258,N_4260);
and U4737 (N_4737,N_4220,N_4330);
and U4738 (N_4738,N_4346,N_4432);
and U4739 (N_4739,N_4354,N_4480);
nand U4740 (N_4740,N_4477,N_4439);
nor U4741 (N_4741,N_4344,N_4263);
xnor U4742 (N_4742,N_4496,N_4221);
or U4743 (N_4743,N_4237,N_4422);
nand U4744 (N_4744,N_4366,N_4443);
nor U4745 (N_4745,N_4286,N_4460);
or U4746 (N_4746,N_4443,N_4285);
and U4747 (N_4747,N_4247,N_4371);
or U4748 (N_4748,N_4324,N_4225);
and U4749 (N_4749,N_4427,N_4275);
nand U4750 (N_4750,N_4474,N_4416);
and U4751 (N_4751,N_4368,N_4230);
nor U4752 (N_4752,N_4381,N_4249);
xor U4753 (N_4753,N_4367,N_4362);
or U4754 (N_4754,N_4250,N_4302);
nor U4755 (N_4755,N_4267,N_4461);
or U4756 (N_4756,N_4301,N_4237);
or U4757 (N_4757,N_4304,N_4440);
xnor U4758 (N_4758,N_4479,N_4418);
nor U4759 (N_4759,N_4480,N_4344);
and U4760 (N_4760,N_4443,N_4453);
nand U4761 (N_4761,N_4450,N_4424);
and U4762 (N_4762,N_4237,N_4211);
or U4763 (N_4763,N_4355,N_4480);
nand U4764 (N_4764,N_4380,N_4404);
or U4765 (N_4765,N_4324,N_4455);
xnor U4766 (N_4766,N_4352,N_4426);
nand U4767 (N_4767,N_4477,N_4497);
or U4768 (N_4768,N_4378,N_4295);
and U4769 (N_4769,N_4498,N_4350);
nor U4770 (N_4770,N_4304,N_4413);
nand U4771 (N_4771,N_4387,N_4273);
xor U4772 (N_4772,N_4366,N_4376);
or U4773 (N_4773,N_4452,N_4281);
xor U4774 (N_4774,N_4486,N_4449);
xor U4775 (N_4775,N_4264,N_4329);
and U4776 (N_4776,N_4423,N_4444);
nor U4777 (N_4777,N_4363,N_4490);
nand U4778 (N_4778,N_4374,N_4303);
nand U4779 (N_4779,N_4436,N_4283);
nor U4780 (N_4780,N_4396,N_4394);
and U4781 (N_4781,N_4494,N_4303);
xnor U4782 (N_4782,N_4438,N_4362);
nor U4783 (N_4783,N_4222,N_4459);
and U4784 (N_4784,N_4202,N_4453);
nor U4785 (N_4785,N_4241,N_4403);
nor U4786 (N_4786,N_4299,N_4280);
xor U4787 (N_4787,N_4464,N_4263);
nor U4788 (N_4788,N_4243,N_4307);
and U4789 (N_4789,N_4254,N_4429);
or U4790 (N_4790,N_4488,N_4217);
or U4791 (N_4791,N_4351,N_4440);
or U4792 (N_4792,N_4423,N_4319);
nor U4793 (N_4793,N_4437,N_4236);
nand U4794 (N_4794,N_4388,N_4445);
and U4795 (N_4795,N_4455,N_4295);
nand U4796 (N_4796,N_4322,N_4279);
nand U4797 (N_4797,N_4374,N_4423);
xnor U4798 (N_4798,N_4246,N_4240);
xor U4799 (N_4799,N_4345,N_4263);
nor U4800 (N_4800,N_4646,N_4717);
and U4801 (N_4801,N_4612,N_4541);
or U4802 (N_4802,N_4573,N_4524);
xor U4803 (N_4803,N_4533,N_4571);
nand U4804 (N_4804,N_4553,N_4597);
xor U4805 (N_4805,N_4509,N_4770);
and U4806 (N_4806,N_4511,N_4599);
nor U4807 (N_4807,N_4631,N_4659);
nor U4808 (N_4808,N_4766,N_4591);
nor U4809 (N_4809,N_4572,N_4680);
or U4810 (N_4810,N_4633,N_4795);
and U4811 (N_4811,N_4764,N_4503);
xnor U4812 (N_4812,N_4748,N_4549);
or U4813 (N_4813,N_4784,N_4514);
nand U4814 (N_4814,N_4551,N_4502);
and U4815 (N_4815,N_4582,N_4506);
nor U4816 (N_4816,N_4647,N_4530);
nor U4817 (N_4817,N_4756,N_4793);
nor U4818 (N_4818,N_4746,N_4730);
nand U4819 (N_4819,N_4671,N_4713);
xor U4820 (N_4820,N_4562,N_4518);
nor U4821 (N_4821,N_4574,N_4508);
or U4822 (N_4822,N_4542,N_4564);
xor U4823 (N_4823,N_4517,N_4663);
nor U4824 (N_4824,N_4681,N_4648);
nand U4825 (N_4825,N_4735,N_4726);
nand U4826 (N_4826,N_4654,N_4622);
nor U4827 (N_4827,N_4516,N_4707);
nor U4828 (N_4828,N_4632,N_4783);
nand U4829 (N_4829,N_4585,N_4604);
nand U4830 (N_4830,N_4611,N_4566);
and U4831 (N_4831,N_4556,N_4652);
xor U4832 (N_4832,N_4769,N_4676);
xor U4833 (N_4833,N_4721,N_4620);
and U4834 (N_4834,N_4501,N_4704);
nand U4835 (N_4835,N_4512,N_4520);
xor U4836 (N_4836,N_4665,N_4535);
and U4837 (N_4837,N_4775,N_4757);
nor U4838 (N_4838,N_4525,N_4618);
xnor U4839 (N_4839,N_4710,N_4600);
and U4840 (N_4840,N_4615,N_4666);
or U4841 (N_4841,N_4588,N_4651);
xor U4842 (N_4842,N_4567,N_4658);
and U4843 (N_4843,N_4569,N_4732);
or U4844 (N_4844,N_4763,N_4543);
and U4845 (N_4845,N_4580,N_4609);
and U4846 (N_4846,N_4657,N_4772);
or U4847 (N_4847,N_4711,N_4690);
xor U4848 (N_4848,N_4660,N_4529);
nor U4849 (N_4849,N_4758,N_4694);
and U4850 (N_4850,N_4649,N_4547);
nand U4851 (N_4851,N_4742,N_4722);
xnor U4852 (N_4852,N_4797,N_4677);
nand U4853 (N_4853,N_4697,N_4531);
and U4854 (N_4854,N_4627,N_4598);
or U4855 (N_4855,N_4526,N_4593);
nor U4856 (N_4856,N_4767,N_4641);
nand U4857 (N_4857,N_4750,N_4522);
nor U4858 (N_4858,N_4555,N_4689);
or U4859 (N_4859,N_4774,N_4755);
xor U4860 (N_4860,N_4539,N_4575);
or U4861 (N_4861,N_4678,N_4528);
and U4862 (N_4862,N_4579,N_4560);
nor U4863 (N_4863,N_4623,N_4634);
nand U4864 (N_4864,N_4637,N_4776);
nand U4865 (N_4865,N_4673,N_4740);
xor U4866 (N_4866,N_4703,N_4626);
and U4867 (N_4867,N_4798,N_4590);
or U4868 (N_4868,N_4504,N_4781);
nor U4869 (N_4869,N_4702,N_4670);
and U4870 (N_4870,N_4794,N_4563);
xnor U4871 (N_4871,N_4537,N_4616);
nor U4872 (N_4872,N_4698,N_4692);
nand U4873 (N_4873,N_4765,N_4521);
nand U4874 (N_4874,N_4624,N_4577);
xnor U4875 (N_4875,N_4736,N_4583);
xor U4876 (N_4876,N_4589,N_4605);
nor U4877 (N_4877,N_4548,N_4661);
or U4878 (N_4878,N_4595,N_4630);
nand U4879 (N_4879,N_4761,N_4510);
nand U4880 (N_4880,N_4554,N_4723);
or U4881 (N_4881,N_4545,N_4636);
xnor U4882 (N_4882,N_4675,N_4603);
nor U4883 (N_4883,N_4714,N_4558);
xnor U4884 (N_4884,N_4662,N_4557);
nand U4885 (N_4885,N_4762,N_4515);
xor U4886 (N_4886,N_4706,N_4638);
xnor U4887 (N_4887,N_4570,N_4602);
nand U4888 (N_4888,N_4741,N_4733);
and U4889 (N_4889,N_4725,N_4619);
nand U4890 (N_4890,N_4792,N_4527);
nor U4891 (N_4891,N_4596,N_4607);
and U4892 (N_4892,N_4534,N_4639);
nand U4893 (N_4893,N_4644,N_4745);
xor U4894 (N_4894,N_4718,N_4532);
xnor U4895 (N_4895,N_4613,N_4601);
or U4896 (N_4896,N_4731,N_4779);
xor U4897 (N_4897,N_4688,N_4789);
and U4898 (N_4898,N_4716,N_4787);
or U4899 (N_4899,N_4561,N_4693);
or U4900 (N_4900,N_4751,N_4610);
nand U4901 (N_4901,N_4581,N_4559);
nand U4902 (N_4902,N_4507,N_4635);
nand U4903 (N_4903,N_4729,N_4513);
xor U4904 (N_4904,N_4696,N_4768);
and U4905 (N_4905,N_4782,N_4739);
nand U4906 (N_4906,N_4686,N_4540);
nand U4907 (N_4907,N_4544,N_4777);
and U4908 (N_4908,N_4674,N_4773);
nor U4909 (N_4909,N_4724,N_4753);
and U4910 (N_4910,N_4550,N_4536);
nor U4911 (N_4911,N_4645,N_4747);
or U4912 (N_4912,N_4606,N_4500);
nor U4913 (N_4913,N_4683,N_4655);
xor U4914 (N_4914,N_4628,N_4640);
xor U4915 (N_4915,N_4780,N_4584);
and U4916 (N_4916,N_4656,N_4653);
xor U4917 (N_4917,N_4738,N_4796);
xnor U4918 (N_4918,N_4728,N_4719);
or U4919 (N_4919,N_4752,N_4715);
nand U4920 (N_4920,N_4771,N_4749);
nor U4921 (N_4921,N_4691,N_4523);
or U4922 (N_4922,N_4621,N_4617);
or U4923 (N_4923,N_4608,N_4701);
nand U4924 (N_4924,N_4642,N_4625);
nor U4925 (N_4925,N_4519,N_4594);
xor U4926 (N_4926,N_4709,N_4759);
nor U4927 (N_4927,N_4705,N_4695);
nand U4928 (N_4928,N_4568,N_4708);
or U4929 (N_4929,N_4682,N_4785);
nor U4930 (N_4930,N_4743,N_4679);
and U4931 (N_4931,N_4667,N_4592);
nand U4932 (N_4932,N_4578,N_4788);
or U4933 (N_4933,N_4700,N_4720);
and U4934 (N_4934,N_4552,N_4643);
xor U4935 (N_4935,N_4754,N_4791);
nand U4936 (N_4936,N_4505,N_4699);
and U4937 (N_4937,N_4799,N_4760);
or U4938 (N_4938,N_4538,N_4687);
or U4939 (N_4939,N_4664,N_4744);
and U4940 (N_4940,N_4672,N_4669);
or U4941 (N_4941,N_4565,N_4786);
and U4942 (N_4942,N_4576,N_4778);
nor U4943 (N_4943,N_4587,N_4684);
xor U4944 (N_4944,N_4790,N_4727);
and U4945 (N_4945,N_4546,N_4737);
nand U4946 (N_4946,N_4734,N_4586);
or U4947 (N_4947,N_4629,N_4650);
xor U4948 (N_4948,N_4712,N_4668);
and U4949 (N_4949,N_4685,N_4614);
nor U4950 (N_4950,N_4552,N_4668);
and U4951 (N_4951,N_4559,N_4505);
or U4952 (N_4952,N_4768,N_4757);
nand U4953 (N_4953,N_4684,N_4715);
and U4954 (N_4954,N_4530,N_4532);
and U4955 (N_4955,N_4561,N_4793);
or U4956 (N_4956,N_4520,N_4613);
and U4957 (N_4957,N_4572,N_4530);
or U4958 (N_4958,N_4517,N_4511);
nand U4959 (N_4959,N_4687,N_4791);
and U4960 (N_4960,N_4628,N_4674);
xor U4961 (N_4961,N_4710,N_4627);
nand U4962 (N_4962,N_4636,N_4512);
xnor U4963 (N_4963,N_4712,N_4641);
and U4964 (N_4964,N_4688,N_4529);
nand U4965 (N_4965,N_4676,N_4507);
or U4966 (N_4966,N_4673,N_4666);
nor U4967 (N_4967,N_4664,N_4582);
and U4968 (N_4968,N_4608,N_4686);
nor U4969 (N_4969,N_4738,N_4781);
nand U4970 (N_4970,N_4546,N_4512);
nor U4971 (N_4971,N_4655,N_4661);
xor U4972 (N_4972,N_4672,N_4562);
and U4973 (N_4973,N_4687,N_4603);
and U4974 (N_4974,N_4513,N_4789);
xor U4975 (N_4975,N_4683,N_4608);
or U4976 (N_4976,N_4758,N_4542);
or U4977 (N_4977,N_4659,N_4530);
nand U4978 (N_4978,N_4757,N_4778);
xnor U4979 (N_4979,N_4528,N_4792);
or U4980 (N_4980,N_4552,N_4631);
nand U4981 (N_4981,N_4767,N_4604);
or U4982 (N_4982,N_4715,N_4699);
xor U4983 (N_4983,N_4719,N_4582);
nand U4984 (N_4984,N_4588,N_4677);
xor U4985 (N_4985,N_4679,N_4688);
nand U4986 (N_4986,N_4737,N_4731);
nand U4987 (N_4987,N_4511,N_4562);
xor U4988 (N_4988,N_4677,N_4638);
or U4989 (N_4989,N_4748,N_4622);
and U4990 (N_4990,N_4732,N_4682);
or U4991 (N_4991,N_4674,N_4614);
xor U4992 (N_4992,N_4720,N_4634);
nor U4993 (N_4993,N_4655,N_4518);
nor U4994 (N_4994,N_4758,N_4650);
xor U4995 (N_4995,N_4504,N_4585);
and U4996 (N_4996,N_4672,N_4544);
nand U4997 (N_4997,N_4690,N_4651);
and U4998 (N_4998,N_4743,N_4662);
xor U4999 (N_4999,N_4543,N_4639);
nor U5000 (N_5000,N_4708,N_4764);
nand U5001 (N_5001,N_4721,N_4573);
nor U5002 (N_5002,N_4555,N_4531);
and U5003 (N_5003,N_4756,N_4669);
xnor U5004 (N_5004,N_4519,N_4630);
nor U5005 (N_5005,N_4589,N_4623);
nand U5006 (N_5006,N_4708,N_4637);
and U5007 (N_5007,N_4752,N_4784);
nor U5008 (N_5008,N_4659,N_4632);
nor U5009 (N_5009,N_4681,N_4676);
nand U5010 (N_5010,N_4762,N_4537);
or U5011 (N_5011,N_4673,N_4560);
xnor U5012 (N_5012,N_4537,N_4632);
and U5013 (N_5013,N_4683,N_4589);
xor U5014 (N_5014,N_4619,N_4631);
or U5015 (N_5015,N_4634,N_4569);
or U5016 (N_5016,N_4699,N_4616);
nand U5017 (N_5017,N_4618,N_4580);
or U5018 (N_5018,N_4751,N_4591);
nor U5019 (N_5019,N_4549,N_4543);
nor U5020 (N_5020,N_4778,N_4747);
and U5021 (N_5021,N_4799,N_4576);
and U5022 (N_5022,N_4762,N_4760);
nand U5023 (N_5023,N_4648,N_4738);
xor U5024 (N_5024,N_4730,N_4609);
and U5025 (N_5025,N_4723,N_4592);
nand U5026 (N_5026,N_4646,N_4626);
or U5027 (N_5027,N_4702,N_4503);
xnor U5028 (N_5028,N_4692,N_4537);
and U5029 (N_5029,N_4643,N_4553);
xnor U5030 (N_5030,N_4780,N_4791);
or U5031 (N_5031,N_4691,N_4563);
and U5032 (N_5032,N_4707,N_4692);
and U5033 (N_5033,N_4512,N_4766);
nand U5034 (N_5034,N_4502,N_4625);
xnor U5035 (N_5035,N_4598,N_4507);
nor U5036 (N_5036,N_4591,N_4572);
and U5037 (N_5037,N_4667,N_4795);
nand U5038 (N_5038,N_4753,N_4750);
xor U5039 (N_5039,N_4534,N_4797);
xor U5040 (N_5040,N_4638,N_4503);
xor U5041 (N_5041,N_4646,N_4698);
or U5042 (N_5042,N_4535,N_4633);
xor U5043 (N_5043,N_4517,N_4736);
nand U5044 (N_5044,N_4623,N_4633);
or U5045 (N_5045,N_4657,N_4787);
and U5046 (N_5046,N_4637,N_4647);
nor U5047 (N_5047,N_4765,N_4709);
and U5048 (N_5048,N_4683,N_4682);
and U5049 (N_5049,N_4582,N_4786);
nor U5050 (N_5050,N_4536,N_4697);
and U5051 (N_5051,N_4796,N_4723);
or U5052 (N_5052,N_4715,N_4505);
nor U5053 (N_5053,N_4726,N_4765);
or U5054 (N_5054,N_4611,N_4762);
nand U5055 (N_5055,N_4544,N_4669);
or U5056 (N_5056,N_4713,N_4586);
and U5057 (N_5057,N_4622,N_4722);
nand U5058 (N_5058,N_4582,N_4731);
nand U5059 (N_5059,N_4732,N_4711);
nor U5060 (N_5060,N_4505,N_4606);
xnor U5061 (N_5061,N_4545,N_4544);
or U5062 (N_5062,N_4744,N_4609);
or U5063 (N_5063,N_4665,N_4546);
nor U5064 (N_5064,N_4798,N_4785);
nand U5065 (N_5065,N_4575,N_4584);
or U5066 (N_5066,N_4551,N_4675);
nand U5067 (N_5067,N_4692,N_4678);
nand U5068 (N_5068,N_4609,N_4556);
or U5069 (N_5069,N_4530,N_4521);
nand U5070 (N_5070,N_4568,N_4671);
nor U5071 (N_5071,N_4516,N_4729);
and U5072 (N_5072,N_4698,N_4667);
nor U5073 (N_5073,N_4782,N_4766);
and U5074 (N_5074,N_4692,N_4741);
xor U5075 (N_5075,N_4780,N_4573);
nor U5076 (N_5076,N_4648,N_4745);
and U5077 (N_5077,N_4604,N_4594);
nor U5078 (N_5078,N_4725,N_4709);
nor U5079 (N_5079,N_4705,N_4749);
nand U5080 (N_5080,N_4704,N_4503);
or U5081 (N_5081,N_4628,N_4581);
nand U5082 (N_5082,N_4589,N_4788);
and U5083 (N_5083,N_4506,N_4515);
and U5084 (N_5084,N_4543,N_4501);
xor U5085 (N_5085,N_4783,N_4663);
nor U5086 (N_5086,N_4608,N_4786);
nand U5087 (N_5087,N_4762,N_4782);
nand U5088 (N_5088,N_4683,N_4726);
and U5089 (N_5089,N_4556,N_4747);
nand U5090 (N_5090,N_4632,N_4669);
and U5091 (N_5091,N_4761,N_4540);
xor U5092 (N_5092,N_4749,N_4723);
and U5093 (N_5093,N_4633,N_4797);
xor U5094 (N_5094,N_4620,N_4508);
and U5095 (N_5095,N_4656,N_4556);
nor U5096 (N_5096,N_4721,N_4532);
nor U5097 (N_5097,N_4625,N_4628);
nor U5098 (N_5098,N_4713,N_4527);
xor U5099 (N_5099,N_4740,N_4570);
nand U5100 (N_5100,N_4955,N_5083);
or U5101 (N_5101,N_4928,N_5088);
and U5102 (N_5102,N_4936,N_4802);
xnor U5103 (N_5103,N_5010,N_5022);
nor U5104 (N_5104,N_4856,N_4912);
and U5105 (N_5105,N_4888,N_4875);
nor U5106 (N_5106,N_5078,N_4845);
nand U5107 (N_5107,N_5030,N_4833);
nor U5108 (N_5108,N_5042,N_4852);
and U5109 (N_5109,N_4886,N_5023);
or U5110 (N_5110,N_4935,N_5048);
and U5111 (N_5111,N_5082,N_4868);
or U5112 (N_5112,N_4987,N_4997);
xor U5113 (N_5113,N_4887,N_5089);
nand U5114 (N_5114,N_4860,N_5000);
nand U5115 (N_5115,N_4971,N_4885);
nor U5116 (N_5116,N_4942,N_4815);
and U5117 (N_5117,N_5097,N_5081);
and U5118 (N_5118,N_4873,N_4882);
nor U5119 (N_5119,N_4854,N_4900);
and U5120 (N_5120,N_4953,N_4991);
nand U5121 (N_5121,N_4908,N_4847);
xor U5122 (N_5122,N_4965,N_4807);
and U5123 (N_5123,N_4903,N_4956);
xor U5124 (N_5124,N_5001,N_4839);
or U5125 (N_5125,N_5084,N_5064);
or U5126 (N_5126,N_4977,N_4995);
nor U5127 (N_5127,N_5043,N_4867);
or U5128 (N_5128,N_5005,N_4906);
xor U5129 (N_5129,N_5062,N_4950);
nand U5130 (N_5130,N_4840,N_4913);
or U5131 (N_5131,N_4941,N_5057);
or U5132 (N_5132,N_4930,N_5099);
nor U5133 (N_5133,N_4907,N_4921);
or U5134 (N_5134,N_5036,N_5006);
and U5135 (N_5135,N_4872,N_5046);
nor U5136 (N_5136,N_4957,N_5017);
xor U5137 (N_5137,N_4880,N_5066);
or U5138 (N_5138,N_4989,N_4855);
nand U5139 (N_5139,N_5014,N_5059);
and U5140 (N_5140,N_4976,N_5018);
xnor U5141 (N_5141,N_5039,N_5074);
or U5142 (N_5142,N_5052,N_4831);
xnor U5143 (N_5143,N_4915,N_4862);
nand U5144 (N_5144,N_4984,N_4938);
xnor U5145 (N_5145,N_4983,N_4843);
and U5146 (N_5146,N_4877,N_5007);
and U5147 (N_5147,N_5056,N_4925);
nor U5148 (N_5148,N_5061,N_4901);
or U5149 (N_5149,N_4892,N_4810);
and U5150 (N_5150,N_5055,N_4943);
xnor U5151 (N_5151,N_5025,N_4905);
xor U5152 (N_5152,N_5034,N_4904);
and U5153 (N_5153,N_5086,N_5011);
nand U5154 (N_5154,N_4825,N_4902);
or U5155 (N_5155,N_4881,N_5054);
xor U5156 (N_5156,N_4974,N_5033);
nand U5157 (N_5157,N_5047,N_4927);
or U5158 (N_5158,N_4924,N_4806);
xnor U5159 (N_5159,N_4961,N_4919);
nor U5160 (N_5160,N_5076,N_4865);
xor U5161 (N_5161,N_5096,N_5035);
or U5162 (N_5162,N_4822,N_4849);
nor U5163 (N_5163,N_4914,N_4846);
or U5164 (N_5164,N_4805,N_5080);
and U5165 (N_5165,N_5002,N_4834);
xnor U5166 (N_5166,N_4883,N_4830);
nand U5167 (N_5167,N_4884,N_4985);
nand U5168 (N_5168,N_5098,N_4945);
or U5169 (N_5169,N_4922,N_4863);
and U5170 (N_5170,N_4981,N_5065);
or U5171 (N_5171,N_4842,N_4951);
or U5172 (N_5172,N_4896,N_4870);
nor U5173 (N_5173,N_5045,N_4968);
and U5174 (N_5174,N_4832,N_5027);
and U5175 (N_5175,N_4821,N_4923);
nor U5176 (N_5176,N_4948,N_5031);
nand U5177 (N_5177,N_4858,N_4857);
nor U5178 (N_5178,N_4836,N_5094);
xnor U5179 (N_5179,N_5040,N_4897);
or U5180 (N_5180,N_4871,N_4859);
xor U5181 (N_5181,N_4978,N_4917);
nand U5182 (N_5182,N_4851,N_5049);
or U5183 (N_5183,N_5038,N_4828);
xnor U5184 (N_5184,N_4979,N_4878);
xnor U5185 (N_5185,N_4894,N_5058);
or U5186 (N_5186,N_5016,N_4804);
nand U5187 (N_5187,N_4920,N_4876);
nand U5188 (N_5188,N_5085,N_5029);
nor U5189 (N_5189,N_4916,N_4931);
nor U5190 (N_5190,N_4823,N_4850);
nor U5191 (N_5191,N_4959,N_5013);
or U5192 (N_5192,N_4835,N_4944);
and U5193 (N_5193,N_4869,N_5024);
and U5194 (N_5194,N_4895,N_4972);
xnor U5195 (N_5195,N_5093,N_4861);
xnor U5196 (N_5196,N_4929,N_4949);
and U5197 (N_5197,N_4980,N_4864);
or U5198 (N_5198,N_4969,N_4937);
and U5199 (N_5199,N_4801,N_4812);
or U5200 (N_5200,N_5051,N_4874);
or U5201 (N_5201,N_4973,N_5026);
and U5202 (N_5202,N_4964,N_5077);
or U5203 (N_5203,N_5032,N_4932);
or U5204 (N_5204,N_4898,N_5087);
nand U5205 (N_5205,N_4866,N_4803);
or U5206 (N_5206,N_4967,N_4813);
and U5207 (N_5207,N_4975,N_4819);
nor U5208 (N_5208,N_5069,N_5037);
nand U5209 (N_5209,N_4818,N_4954);
and U5210 (N_5210,N_4946,N_4811);
or U5211 (N_5211,N_4958,N_4963);
nand U5212 (N_5212,N_4910,N_5067);
xor U5213 (N_5213,N_5050,N_4890);
nor U5214 (N_5214,N_4808,N_4999);
and U5215 (N_5215,N_4933,N_4814);
nand U5216 (N_5216,N_4817,N_4990);
xor U5217 (N_5217,N_4824,N_4829);
nand U5218 (N_5218,N_4992,N_4838);
nand U5219 (N_5219,N_5041,N_4816);
nand U5220 (N_5220,N_5072,N_4826);
xor U5221 (N_5221,N_4986,N_5091);
or U5222 (N_5222,N_5075,N_4891);
nor U5223 (N_5223,N_4988,N_4940);
nand U5224 (N_5224,N_5015,N_5071);
nor U5225 (N_5225,N_4800,N_4827);
or U5226 (N_5226,N_4952,N_5008);
or U5227 (N_5227,N_5090,N_5079);
and U5228 (N_5228,N_4947,N_5020);
nand U5229 (N_5229,N_4909,N_4960);
nor U5230 (N_5230,N_5009,N_5063);
nor U5231 (N_5231,N_5068,N_4926);
xnor U5232 (N_5232,N_4809,N_5021);
xnor U5233 (N_5233,N_4848,N_4918);
nor U5234 (N_5234,N_5028,N_5053);
nor U5235 (N_5235,N_5044,N_5060);
or U5236 (N_5236,N_5012,N_4982);
nand U5237 (N_5237,N_4934,N_5003);
xor U5238 (N_5238,N_4993,N_5070);
nand U5239 (N_5239,N_4966,N_4962);
xor U5240 (N_5240,N_5073,N_5095);
nor U5241 (N_5241,N_4844,N_4893);
nor U5242 (N_5242,N_4889,N_4970);
xor U5243 (N_5243,N_4820,N_4837);
nor U5244 (N_5244,N_4879,N_4939);
and U5245 (N_5245,N_5004,N_4853);
or U5246 (N_5246,N_5092,N_4911);
xor U5247 (N_5247,N_4899,N_4996);
xnor U5248 (N_5248,N_4994,N_5019);
nand U5249 (N_5249,N_4841,N_4998);
and U5250 (N_5250,N_5016,N_4999);
xor U5251 (N_5251,N_5082,N_5016);
nand U5252 (N_5252,N_4992,N_5066);
or U5253 (N_5253,N_5025,N_4934);
xnor U5254 (N_5254,N_4942,N_4928);
xnor U5255 (N_5255,N_5058,N_4960);
and U5256 (N_5256,N_4843,N_4908);
nand U5257 (N_5257,N_5013,N_4945);
or U5258 (N_5258,N_4876,N_5065);
and U5259 (N_5259,N_4866,N_4830);
nor U5260 (N_5260,N_4907,N_5075);
or U5261 (N_5261,N_4824,N_4822);
nand U5262 (N_5262,N_4873,N_5069);
or U5263 (N_5263,N_5076,N_4940);
xnor U5264 (N_5264,N_5009,N_4986);
and U5265 (N_5265,N_4852,N_4961);
and U5266 (N_5266,N_5005,N_5028);
xor U5267 (N_5267,N_4883,N_5086);
nand U5268 (N_5268,N_5054,N_5074);
and U5269 (N_5269,N_4906,N_4923);
nand U5270 (N_5270,N_4907,N_4974);
nand U5271 (N_5271,N_5002,N_4826);
nor U5272 (N_5272,N_5075,N_4844);
or U5273 (N_5273,N_4923,N_4930);
and U5274 (N_5274,N_5093,N_4880);
xnor U5275 (N_5275,N_4936,N_4873);
and U5276 (N_5276,N_5069,N_5011);
xor U5277 (N_5277,N_4839,N_4974);
xnor U5278 (N_5278,N_4997,N_4875);
or U5279 (N_5279,N_4931,N_4907);
or U5280 (N_5280,N_5086,N_4828);
nand U5281 (N_5281,N_4974,N_4991);
and U5282 (N_5282,N_4961,N_4973);
and U5283 (N_5283,N_4824,N_5019);
xnor U5284 (N_5284,N_4869,N_4823);
nand U5285 (N_5285,N_4839,N_5057);
nor U5286 (N_5286,N_4979,N_4970);
or U5287 (N_5287,N_5059,N_5058);
or U5288 (N_5288,N_5098,N_5072);
nor U5289 (N_5289,N_4932,N_5020);
nor U5290 (N_5290,N_4867,N_5067);
and U5291 (N_5291,N_5083,N_4881);
nor U5292 (N_5292,N_4827,N_4971);
and U5293 (N_5293,N_4907,N_4925);
and U5294 (N_5294,N_4955,N_4974);
nor U5295 (N_5295,N_5029,N_5048);
nand U5296 (N_5296,N_5061,N_4948);
or U5297 (N_5297,N_5094,N_4854);
nand U5298 (N_5298,N_4846,N_5061);
or U5299 (N_5299,N_4984,N_4819);
nand U5300 (N_5300,N_4863,N_4954);
xnor U5301 (N_5301,N_4955,N_4826);
or U5302 (N_5302,N_5060,N_5082);
nand U5303 (N_5303,N_5093,N_4826);
nand U5304 (N_5304,N_4913,N_4948);
xor U5305 (N_5305,N_4861,N_4884);
nor U5306 (N_5306,N_4866,N_4991);
nor U5307 (N_5307,N_4890,N_4989);
or U5308 (N_5308,N_5026,N_5074);
or U5309 (N_5309,N_4950,N_4903);
nor U5310 (N_5310,N_4844,N_4837);
nand U5311 (N_5311,N_4814,N_4856);
nor U5312 (N_5312,N_5044,N_4960);
nor U5313 (N_5313,N_4905,N_4900);
xnor U5314 (N_5314,N_5041,N_5082);
xor U5315 (N_5315,N_5013,N_5005);
or U5316 (N_5316,N_5070,N_5026);
nor U5317 (N_5317,N_4899,N_4864);
xnor U5318 (N_5318,N_4957,N_4835);
nand U5319 (N_5319,N_5029,N_4954);
nor U5320 (N_5320,N_4890,N_4997);
and U5321 (N_5321,N_4873,N_4892);
xor U5322 (N_5322,N_4987,N_4900);
or U5323 (N_5323,N_5082,N_4884);
nand U5324 (N_5324,N_4883,N_5099);
nand U5325 (N_5325,N_4877,N_5062);
nand U5326 (N_5326,N_4957,N_4825);
or U5327 (N_5327,N_5068,N_5023);
nor U5328 (N_5328,N_4947,N_4919);
xnor U5329 (N_5329,N_4875,N_5032);
and U5330 (N_5330,N_4967,N_5032);
and U5331 (N_5331,N_5006,N_4865);
and U5332 (N_5332,N_4812,N_4974);
nor U5333 (N_5333,N_4852,N_5054);
nand U5334 (N_5334,N_4953,N_4900);
and U5335 (N_5335,N_5093,N_4882);
xnor U5336 (N_5336,N_4842,N_4992);
nand U5337 (N_5337,N_5005,N_4841);
and U5338 (N_5338,N_4923,N_4881);
and U5339 (N_5339,N_5059,N_5060);
xor U5340 (N_5340,N_4967,N_5018);
nor U5341 (N_5341,N_5071,N_4905);
nor U5342 (N_5342,N_5033,N_4839);
or U5343 (N_5343,N_4876,N_4925);
xor U5344 (N_5344,N_5017,N_5011);
xor U5345 (N_5345,N_5073,N_4813);
nor U5346 (N_5346,N_4919,N_4965);
xor U5347 (N_5347,N_5001,N_4836);
or U5348 (N_5348,N_4977,N_4820);
and U5349 (N_5349,N_4832,N_4813);
nand U5350 (N_5350,N_5066,N_5016);
or U5351 (N_5351,N_5074,N_5069);
xor U5352 (N_5352,N_4906,N_4913);
nor U5353 (N_5353,N_4968,N_4943);
nand U5354 (N_5354,N_5096,N_4886);
nor U5355 (N_5355,N_5050,N_5017);
nand U5356 (N_5356,N_4838,N_4963);
xor U5357 (N_5357,N_4912,N_5092);
nand U5358 (N_5358,N_4906,N_4879);
nand U5359 (N_5359,N_5083,N_4919);
and U5360 (N_5360,N_4907,N_5008);
and U5361 (N_5361,N_4941,N_5004);
and U5362 (N_5362,N_4945,N_5010);
and U5363 (N_5363,N_5007,N_4811);
and U5364 (N_5364,N_5027,N_4965);
nand U5365 (N_5365,N_4908,N_5083);
nor U5366 (N_5366,N_5030,N_5067);
nor U5367 (N_5367,N_5058,N_4995);
nor U5368 (N_5368,N_4956,N_5096);
nor U5369 (N_5369,N_5035,N_5039);
or U5370 (N_5370,N_4994,N_4938);
nor U5371 (N_5371,N_4917,N_5076);
or U5372 (N_5372,N_4921,N_5042);
xnor U5373 (N_5373,N_4860,N_4826);
xnor U5374 (N_5374,N_4836,N_4800);
and U5375 (N_5375,N_4972,N_4843);
xor U5376 (N_5376,N_4858,N_4948);
nand U5377 (N_5377,N_4939,N_5085);
nor U5378 (N_5378,N_4832,N_4991);
and U5379 (N_5379,N_4917,N_4941);
xnor U5380 (N_5380,N_5088,N_4995);
nor U5381 (N_5381,N_5097,N_4930);
nand U5382 (N_5382,N_4924,N_5011);
xnor U5383 (N_5383,N_4917,N_5092);
xnor U5384 (N_5384,N_4928,N_4804);
nand U5385 (N_5385,N_4975,N_4957);
nor U5386 (N_5386,N_4821,N_4842);
and U5387 (N_5387,N_4889,N_4972);
and U5388 (N_5388,N_4878,N_4972);
xnor U5389 (N_5389,N_4942,N_5059);
xnor U5390 (N_5390,N_4915,N_5038);
and U5391 (N_5391,N_5005,N_4806);
and U5392 (N_5392,N_5012,N_5038);
nor U5393 (N_5393,N_4993,N_4877);
or U5394 (N_5394,N_5026,N_4918);
nor U5395 (N_5395,N_4912,N_4900);
or U5396 (N_5396,N_5053,N_4910);
nand U5397 (N_5397,N_5057,N_5045);
or U5398 (N_5398,N_4945,N_4888);
or U5399 (N_5399,N_5093,N_4968);
or U5400 (N_5400,N_5169,N_5235);
nor U5401 (N_5401,N_5393,N_5314);
nand U5402 (N_5402,N_5373,N_5369);
xnor U5403 (N_5403,N_5328,N_5221);
nand U5404 (N_5404,N_5307,N_5321);
nor U5405 (N_5405,N_5339,N_5318);
nor U5406 (N_5406,N_5262,N_5316);
and U5407 (N_5407,N_5120,N_5124);
xnor U5408 (N_5408,N_5215,N_5313);
and U5409 (N_5409,N_5255,N_5128);
or U5410 (N_5410,N_5150,N_5299);
or U5411 (N_5411,N_5140,N_5312);
or U5412 (N_5412,N_5164,N_5325);
nor U5413 (N_5413,N_5268,N_5345);
nand U5414 (N_5414,N_5204,N_5118);
nor U5415 (N_5415,N_5319,N_5352);
or U5416 (N_5416,N_5155,N_5288);
and U5417 (N_5417,N_5217,N_5156);
or U5418 (N_5418,N_5210,N_5361);
and U5419 (N_5419,N_5233,N_5119);
or U5420 (N_5420,N_5182,N_5368);
xnor U5421 (N_5421,N_5161,N_5175);
or U5422 (N_5422,N_5212,N_5218);
nand U5423 (N_5423,N_5146,N_5323);
nand U5424 (N_5424,N_5263,N_5102);
or U5425 (N_5425,N_5278,N_5335);
and U5426 (N_5426,N_5224,N_5272);
nand U5427 (N_5427,N_5162,N_5103);
xor U5428 (N_5428,N_5214,N_5107);
or U5429 (N_5429,N_5294,N_5139);
nor U5430 (N_5430,N_5179,N_5227);
nor U5431 (N_5431,N_5201,N_5358);
xor U5432 (N_5432,N_5160,N_5327);
and U5433 (N_5433,N_5283,N_5194);
nand U5434 (N_5434,N_5117,N_5289);
or U5435 (N_5435,N_5153,N_5122);
and U5436 (N_5436,N_5159,N_5396);
nand U5437 (N_5437,N_5306,N_5209);
nor U5438 (N_5438,N_5116,N_5362);
nor U5439 (N_5439,N_5195,N_5129);
or U5440 (N_5440,N_5101,N_5273);
or U5441 (N_5441,N_5338,N_5347);
nand U5442 (N_5442,N_5275,N_5183);
or U5443 (N_5443,N_5106,N_5178);
nand U5444 (N_5444,N_5348,N_5186);
nand U5445 (N_5445,N_5144,N_5320);
xor U5446 (N_5446,N_5308,N_5193);
nand U5447 (N_5447,N_5246,N_5104);
and U5448 (N_5448,N_5271,N_5398);
nor U5449 (N_5449,N_5211,N_5170);
or U5450 (N_5450,N_5105,N_5282);
nand U5451 (N_5451,N_5114,N_5166);
nand U5452 (N_5452,N_5324,N_5390);
xor U5453 (N_5453,N_5163,N_5229);
nor U5454 (N_5454,N_5252,N_5350);
or U5455 (N_5455,N_5364,N_5142);
or U5456 (N_5456,N_5113,N_5340);
or U5457 (N_5457,N_5250,N_5191);
nand U5458 (N_5458,N_5219,N_5213);
or U5459 (N_5459,N_5109,N_5165);
and U5460 (N_5460,N_5147,N_5239);
xor U5461 (N_5461,N_5137,N_5344);
nor U5462 (N_5462,N_5203,N_5134);
nand U5463 (N_5463,N_5216,N_5395);
xnor U5464 (N_5464,N_5130,N_5279);
and U5465 (N_5465,N_5176,N_5258);
nand U5466 (N_5466,N_5293,N_5208);
nor U5467 (N_5467,N_5322,N_5357);
nand U5468 (N_5468,N_5192,N_5317);
or U5469 (N_5469,N_5280,N_5135);
or U5470 (N_5470,N_5110,N_5173);
xnor U5471 (N_5471,N_5197,N_5123);
nor U5472 (N_5472,N_5355,N_5247);
nand U5473 (N_5473,N_5363,N_5349);
and U5474 (N_5474,N_5277,N_5200);
nand U5475 (N_5475,N_5380,N_5154);
nand U5476 (N_5476,N_5222,N_5291);
nand U5477 (N_5477,N_5240,N_5254);
and U5478 (N_5478,N_5196,N_5223);
and U5479 (N_5479,N_5133,N_5292);
nand U5480 (N_5480,N_5243,N_5365);
xor U5481 (N_5481,N_5285,N_5331);
nor U5482 (N_5482,N_5371,N_5187);
nor U5483 (N_5483,N_5377,N_5394);
and U5484 (N_5484,N_5310,N_5112);
nand U5485 (N_5485,N_5346,N_5351);
nor U5486 (N_5486,N_5256,N_5172);
or U5487 (N_5487,N_5333,N_5332);
nand U5488 (N_5488,N_5284,N_5386);
and U5489 (N_5489,N_5354,N_5330);
xor U5490 (N_5490,N_5231,N_5274);
nand U5491 (N_5491,N_5184,N_5108);
and U5492 (N_5492,N_5382,N_5148);
xor U5493 (N_5493,N_5185,N_5302);
nand U5494 (N_5494,N_5336,N_5359);
and U5495 (N_5495,N_5337,N_5127);
nor U5496 (N_5496,N_5230,N_5136);
and U5497 (N_5497,N_5367,N_5309);
nand U5498 (N_5498,N_5251,N_5300);
and U5499 (N_5499,N_5366,N_5241);
or U5500 (N_5500,N_5381,N_5259);
nand U5501 (N_5501,N_5225,N_5132);
or U5502 (N_5502,N_5249,N_5290);
nor U5503 (N_5503,N_5334,N_5376);
or U5504 (N_5504,N_5242,N_5177);
xnor U5505 (N_5505,N_5190,N_5392);
xnor U5506 (N_5506,N_5174,N_5111);
xor U5507 (N_5507,N_5267,N_5261);
nor U5508 (N_5508,N_5238,N_5206);
or U5509 (N_5509,N_5295,N_5383);
xnor U5510 (N_5510,N_5384,N_5244);
nand U5511 (N_5511,N_5181,N_5360);
and U5512 (N_5512,N_5207,N_5388);
nand U5513 (N_5513,N_5121,N_5257);
or U5514 (N_5514,N_5389,N_5260);
nand U5515 (N_5515,N_5315,N_5397);
and U5516 (N_5516,N_5171,N_5228);
xor U5517 (N_5517,N_5270,N_5353);
nor U5518 (N_5518,N_5236,N_5205);
nand U5519 (N_5519,N_5149,N_5167);
xor U5520 (N_5520,N_5297,N_5375);
nand U5521 (N_5521,N_5296,N_5141);
nor U5522 (N_5522,N_5145,N_5287);
or U5523 (N_5523,N_5311,N_5188);
nand U5524 (N_5524,N_5391,N_5232);
xnor U5525 (N_5525,N_5115,N_5126);
and U5526 (N_5526,N_5303,N_5168);
nor U5527 (N_5527,N_5372,N_5189);
xor U5528 (N_5528,N_5286,N_5264);
xnor U5529 (N_5529,N_5199,N_5265);
nand U5530 (N_5530,N_5131,N_5298);
or U5531 (N_5531,N_5138,N_5180);
xor U5532 (N_5532,N_5329,N_5379);
or U5533 (N_5533,N_5276,N_5301);
xor U5534 (N_5534,N_5152,N_5281);
or U5535 (N_5535,N_5266,N_5234);
or U5536 (N_5536,N_5125,N_5220);
nor U5537 (N_5537,N_5378,N_5202);
nor U5538 (N_5538,N_5158,N_5304);
or U5539 (N_5539,N_5253,N_5343);
nor U5540 (N_5540,N_5385,N_5245);
nor U5541 (N_5541,N_5342,N_5269);
nand U5542 (N_5542,N_5226,N_5356);
nand U5543 (N_5543,N_5157,N_5326);
and U5544 (N_5544,N_5341,N_5399);
or U5545 (N_5545,N_5100,N_5370);
xnor U5546 (N_5546,N_5237,N_5387);
xor U5547 (N_5547,N_5248,N_5374);
nor U5548 (N_5548,N_5151,N_5305);
xor U5549 (N_5549,N_5143,N_5198);
or U5550 (N_5550,N_5380,N_5297);
and U5551 (N_5551,N_5384,N_5150);
nor U5552 (N_5552,N_5267,N_5162);
xnor U5553 (N_5553,N_5102,N_5166);
xor U5554 (N_5554,N_5267,N_5300);
xor U5555 (N_5555,N_5149,N_5274);
nand U5556 (N_5556,N_5361,N_5207);
or U5557 (N_5557,N_5180,N_5380);
xnor U5558 (N_5558,N_5359,N_5205);
or U5559 (N_5559,N_5268,N_5313);
and U5560 (N_5560,N_5276,N_5287);
and U5561 (N_5561,N_5295,N_5350);
xnor U5562 (N_5562,N_5188,N_5379);
and U5563 (N_5563,N_5155,N_5225);
nor U5564 (N_5564,N_5158,N_5121);
nor U5565 (N_5565,N_5311,N_5220);
and U5566 (N_5566,N_5126,N_5124);
nand U5567 (N_5567,N_5182,N_5379);
nand U5568 (N_5568,N_5386,N_5287);
nor U5569 (N_5569,N_5137,N_5176);
nand U5570 (N_5570,N_5368,N_5130);
and U5571 (N_5571,N_5348,N_5375);
or U5572 (N_5572,N_5323,N_5380);
and U5573 (N_5573,N_5159,N_5265);
or U5574 (N_5574,N_5292,N_5256);
and U5575 (N_5575,N_5150,N_5265);
nor U5576 (N_5576,N_5144,N_5151);
or U5577 (N_5577,N_5211,N_5397);
nand U5578 (N_5578,N_5395,N_5335);
or U5579 (N_5579,N_5161,N_5347);
nor U5580 (N_5580,N_5240,N_5272);
nand U5581 (N_5581,N_5178,N_5211);
xor U5582 (N_5582,N_5222,N_5381);
and U5583 (N_5583,N_5305,N_5162);
or U5584 (N_5584,N_5102,N_5250);
nor U5585 (N_5585,N_5358,N_5204);
xor U5586 (N_5586,N_5132,N_5228);
xnor U5587 (N_5587,N_5278,N_5388);
and U5588 (N_5588,N_5296,N_5140);
xnor U5589 (N_5589,N_5283,N_5336);
and U5590 (N_5590,N_5300,N_5205);
and U5591 (N_5591,N_5212,N_5384);
nand U5592 (N_5592,N_5136,N_5280);
nand U5593 (N_5593,N_5163,N_5232);
and U5594 (N_5594,N_5229,N_5264);
xor U5595 (N_5595,N_5383,N_5233);
and U5596 (N_5596,N_5384,N_5364);
nand U5597 (N_5597,N_5192,N_5299);
and U5598 (N_5598,N_5140,N_5154);
nand U5599 (N_5599,N_5384,N_5339);
nand U5600 (N_5600,N_5227,N_5373);
nand U5601 (N_5601,N_5337,N_5215);
nor U5602 (N_5602,N_5289,N_5141);
and U5603 (N_5603,N_5270,N_5115);
nor U5604 (N_5604,N_5204,N_5316);
nor U5605 (N_5605,N_5268,N_5120);
nor U5606 (N_5606,N_5298,N_5155);
or U5607 (N_5607,N_5396,N_5340);
or U5608 (N_5608,N_5375,N_5121);
and U5609 (N_5609,N_5390,N_5201);
nor U5610 (N_5610,N_5282,N_5358);
nand U5611 (N_5611,N_5391,N_5177);
or U5612 (N_5612,N_5230,N_5384);
nor U5613 (N_5613,N_5363,N_5282);
nand U5614 (N_5614,N_5393,N_5136);
and U5615 (N_5615,N_5124,N_5341);
nand U5616 (N_5616,N_5276,N_5237);
xnor U5617 (N_5617,N_5110,N_5127);
and U5618 (N_5618,N_5281,N_5147);
xor U5619 (N_5619,N_5278,N_5144);
nand U5620 (N_5620,N_5248,N_5258);
or U5621 (N_5621,N_5305,N_5313);
or U5622 (N_5622,N_5373,N_5252);
nor U5623 (N_5623,N_5105,N_5229);
nand U5624 (N_5624,N_5302,N_5377);
and U5625 (N_5625,N_5203,N_5187);
nor U5626 (N_5626,N_5269,N_5396);
nand U5627 (N_5627,N_5393,N_5260);
nor U5628 (N_5628,N_5176,N_5275);
nand U5629 (N_5629,N_5240,N_5177);
xnor U5630 (N_5630,N_5366,N_5294);
and U5631 (N_5631,N_5300,N_5289);
or U5632 (N_5632,N_5271,N_5349);
or U5633 (N_5633,N_5204,N_5220);
and U5634 (N_5634,N_5192,N_5347);
nor U5635 (N_5635,N_5283,N_5324);
nand U5636 (N_5636,N_5395,N_5347);
or U5637 (N_5637,N_5251,N_5295);
nor U5638 (N_5638,N_5371,N_5217);
nor U5639 (N_5639,N_5395,N_5206);
xor U5640 (N_5640,N_5386,N_5148);
xor U5641 (N_5641,N_5119,N_5247);
and U5642 (N_5642,N_5339,N_5153);
and U5643 (N_5643,N_5198,N_5377);
and U5644 (N_5644,N_5183,N_5156);
nand U5645 (N_5645,N_5156,N_5220);
and U5646 (N_5646,N_5173,N_5313);
or U5647 (N_5647,N_5331,N_5103);
nand U5648 (N_5648,N_5332,N_5127);
xnor U5649 (N_5649,N_5117,N_5273);
and U5650 (N_5650,N_5381,N_5269);
nand U5651 (N_5651,N_5351,N_5296);
or U5652 (N_5652,N_5190,N_5166);
nor U5653 (N_5653,N_5221,N_5148);
or U5654 (N_5654,N_5357,N_5194);
xnor U5655 (N_5655,N_5224,N_5292);
xnor U5656 (N_5656,N_5115,N_5190);
or U5657 (N_5657,N_5106,N_5100);
or U5658 (N_5658,N_5295,N_5226);
nand U5659 (N_5659,N_5319,N_5152);
xnor U5660 (N_5660,N_5399,N_5237);
and U5661 (N_5661,N_5112,N_5226);
xor U5662 (N_5662,N_5380,N_5386);
nand U5663 (N_5663,N_5181,N_5159);
nor U5664 (N_5664,N_5174,N_5302);
xor U5665 (N_5665,N_5209,N_5313);
xor U5666 (N_5666,N_5308,N_5256);
nor U5667 (N_5667,N_5343,N_5259);
or U5668 (N_5668,N_5381,N_5341);
xor U5669 (N_5669,N_5149,N_5312);
nand U5670 (N_5670,N_5325,N_5351);
or U5671 (N_5671,N_5270,N_5224);
nand U5672 (N_5672,N_5258,N_5162);
and U5673 (N_5673,N_5201,N_5155);
and U5674 (N_5674,N_5319,N_5135);
nor U5675 (N_5675,N_5308,N_5266);
and U5676 (N_5676,N_5243,N_5397);
xnor U5677 (N_5677,N_5359,N_5122);
and U5678 (N_5678,N_5102,N_5188);
and U5679 (N_5679,N_5295,N_5327);
xor U5680 (N_5680,N_5151,N_5284);
and U5681 (N_5681,N_5385,N_5306);
or U5682 (N_5682,N_5241,N_5207);
nor U5683 (N_5683,N_5217,N_5386);
nand U5684 (N_5684,N_5289,N_5203);
xor U5685 (N_5685,N_5221,N_5169);
nand U5686 (N_5686,N_5198,N_5343);
and U5687 (N_5687,N_5395,N_5191);
and U5688 (N_5688,N_5187,N_5145);
and U5689 (N_5689,N_5261,N_5101);
xor U5690 (N_5690,N_5182,N_5322);
nor U5691 (N_5691,N_5187,N_5242);
nor U5692 (N_5692,N_5122,N_5345);
or U5693 (N_5693,N_5366,N_5206);
nor U5694 (N_5694,N_5198,N_5145);
xnor U5695 (N_5695,N_5241,N_5166);
nand U5696 (N_5696,N_5325,N_5237);
nand U5697 (N_5697,N_5383,N_5121);
xor U5698 (N_5698,N_5121,N_5287);
nor U5699 (N_5699,N_5376,N_5390);
nor U5700 (N_5700,N_5663,N_5661);
nor U5701 (N_5701,N_5496,N_5480);
nand U5702 (N_5702,N_5505,N_5434);
nor U5703 (N_5703,N_5407,N_5588);
xor U5704 (N_5704,N_5414,N_5648);
xnor U5705 (N_5705,N_5499,N_5699);
xor U5706 (N_5706,N_5637,N_5654);
nand U5707 (N_5707,N_5581,N_5600);
or U5708 (N_5708,N_5584,N_5506);
or U5709 (N_5709,N_5669,N_5463);
xor U5710 (N_5710,N_5538,N_5446);
or U5711 (N_5711,N_5482,N_5483);
and U5712 (N_5712,N_5668,N_5582);
or U5713 (N_5713,N_5556,N_5611);
or U5714 (N_5714,N_5417,N_5691);
xor U5715 (N_5715,N_5597,N_5469);
or U5716 (N_5716,N_5625,N_5612);
or U5717 (N_5717,N_5491,N_5686);
xor U5718 (N_5718,N_5546,N_5626);
xnor U5719 (N_5719,N_5695,N_5614);
nor U5720 (N_5720,N_5453,N_5440);
and U5721 (N_5721,N_5490,N_5497);
nor U5722 (N_5722,N_5411,N_5572);
xor U5723 (N_5723,N_5660,N_5529);
and U5724 (N_5724,N_5481,N_5460);
or U5725 (N_5725,N_5569,N_5461);
or U5726 (N_5726,N_5655,N_5579);
and U5727 (N_5727,N_5587,N_5647);
and U5728 (N_5728,N_5601,N_5590);
nor U5729 (N_5729,N_5642,N_5623);
nand U5730 (N_5730,N_5689,N_5478);
nand U5731 (N_5731,N_5641,N_5441);
nand U5732 (N_5732,N_5585,N_5489);
nand U5733 (N_5733,N_5462,N_5595);
xnor U5734 (N_5734,N_5653,N_5436);
nand U5735 (N_5735,N_5634,N_5456);
xor U5736 (N_5736,N_5630,N_5598);
nor U5737 (N_5737,N_5494,N_5594);
nand U5738 (N_5738,N_5692,N_5466);
nand U5739 (N_5739,N_5509,N_5474);
nor U5740 (N_5740,N_5658,N_5565);
nor U5741 (N_5741,N_5423,N_5685);
nand U5742 (N_5742,N_5656,N_5633);
xor U5743 (N_5743,N_5652,N_5425);
or U5744 (N_5744,N_5681,N_5560);
and U5745 (N_5745,N_5548,N_5559);
and U5746 (N_5746,N_5618,N_5694);
xnor U5747 (N_5747,N_5488,N_5540);
or U5748 (N_5748,N_5542,N_5528);
or U5749 (N_5749,N_5552,N_5455);
nor U5750 (N_5750,N_5541,N_5418);
and U5751 (N_5751,N_5532,N_5454);
xor U5752 (N_5752,N_5570,N_5687);
xnor U5753 (N_5753,N_5659,N_5433);
or U5754 (N_5754,N_5521,N_5646);
xnor U5755 (N_5755,N_5527,N_5606);
nand U5756 (N_5756,N_5602,N_5427);
nand U5757 (N_5757,N_5519,N_5696);
nand U5758 (N_5758,N_5467,N_5403);
nor U5759 (N_5759,N_5664,N_5406);
or U5760 (N_5760,N_5503,N_5635);
xor U5761 (N_5761,N_5688,N_5525);
or U5762 (N_5762,N_5617,N_5616);
and U5763 (N_5763,N_5530,N_5693);
xor U5764 (N_5764,N_5512,N_5543);
nor U5765 (N_5765,N_5421,N_5640);
nor U5766 (N_5766,N_5596,N_5645);
nand U5767 (N_5767,N_5471,N_5674);
or U5768 (N_5768,N_5487,N_5516);
xor U5769 (N_5769,N_5501,N_5452);
nor U5770 (N_5770,N_5666,N_5589);
nor U5771 (N_5771,N_5628,N_5680);
and U5772 (N_5772,N_5472,N_5558);
or U5773 (N_5773,N_5500,N_5415);
nand U5774 (N_5774,N_5574,N_5599);
nor U5775 (N_5775,N_5533,N_5408);
nor U5776 (N_5776,N_5522,N_5444);
nor U5777 (N_5777,N_5464,N_5493);
nor U5778 (N_5778,N_5429,N_5604);
and U5779 (N_5779,N_5537,N_5507);
and U5780 (N_5780,N_5622,N_5419);
xnor U5781 (N_5781,N_5672,N_5610);
or U5782 (N_5782,N_5449,N_5435);
or U5783 (N_5783,N_5431,N_5682);
nand U5784 (N_5784,N_5534,N_5555);
and U5785 (N_5785,N_5562,N_5510);
nand U5786 (N_5786,N_5524,N_5508);
xnor U5787 (N_5787,N_5586,N_5662);
or U5788 (N_5788,N_5549,N_5450);
xor U5789 (N_5789,N_5550,N_5677);
and U5790 (N_5790,N_5665,N_5420);
or U5791 (N_5791,N_5627,N_5475);
nand U5792 (N_5792,N_5451,N_5485);
xnor U5793 (N_5793,N_5644,N_5643);
or U5794 (N_5794,N_5670,N_5470);
xor U5795 (N_5795,N_5442,N_5486);
xnor U5796 (N_5796,N_5650,N_5424);
nor U5797 (N_5797,N_5445,N_5473);
or U5798 (N_5798,N_5520,N_5576);
and U5799 (N_5799,N_5636,N_5437);
and U5800 (N_5800,N_5575,N_5563);
or U5801 (N_5801,N_5613,N_5416);
and U5802 (N_5802,N_5631,N_5438);
and U5803 (N_5803,N_5426,N_5405);
xor U5804 (N_5804,N_5536,N_5608);
nand U5805 (N_5805,N_5539,N_5458);
nand U5806 (N_5806,N_5432,N_5573);
or U5807 (N_5807,N_5523,N_5553);
xor U5808 (N_5808,N_5675,N_5676);
nor U5809 (N_5809,N_5697,N_5544);
nand U5810 (N_5810,N_5412,N_5526);
xor U5811 (N_5811,N_5567,N_5413);
and U5812 (N_5812,N_5422,N_5443);
and U5813 (N_5813,N_5492,N_5684);
and U5814 (N_5814,N_5657,N_5678);
nor U5815 (N_5815,N_5621,N_5511);
xor U5816 (N_5816,N_5639,N_5402);
xor U5817 (N_5817,N_5607,N_5571);
or U5818 (N_5818,N_5401,N_5428);
xnor U5819 (N_5819,N_5578,N_5410);
nor U5820 (N_5820,N_5593,N_5409);
or U5821 (N_5821,N_5517,N_5498);
xor U5822 (N_5822,N_5459,N_5457);
and U5823 (N_5823,N_5698,N_5638);
nor U5824 (N_5824,N_5447,N_5583);
or U5825 (N_5825,N_5439,N_5404);
nor U5826 (N_5826,N_5564,N_5468);
nand U5827 (N_5827,N_5518,N_5603);
nor U5828 (N_5828,N_5577,N_5620);
or U5829 (N_5829,N_5624,N_5514);
nor U5830 (N_5830,N_5535,N_5591);
xor U5831 (N_5831,N_5476,N_5479);
and U5832 (N_5832,N_5554,N_5495);
nor U5833 (N_5833,N_5561,N_5651);
and U5834 (N_5834,N_5545,N_5683);
xor U5835 (N_5835,N_5580,N_5629);
nand U5836 (N_5836,N_5592,N_5515);
or U5837 (N_5837,N_5465,N_5679);
or U5838 (N_5838,N_5690,N_5484);
xor U5839 (N_5839,N_5667,N_5504);
nand U5840 (N_5840,N_5649,N_5632);
nor U5841 (N_5841,N_5400,N_5619);
xor U5842 (N_5842,N_5448,N_5547);
or U5843 (N_5843,N_5566,N_5531);
xnor U5844 (N_5844,N_5551,N_5430);
nand U5845 (N_5845,N_5502,N_5671);
or U5846 (N_5846,N_5557,N_5609);
xnor U5847 (N_5847,N_5568,N_5673);
or U5848 (N_5848,N_5615,N_5513);
or U5849 (N_5849,N_5605,N_5477);
nand U5850 (N_5850,N_5429,N_5443);
and U5851 (N_5851,N_5410,N_5669);
nand U5852 (N_5852,N_5490,N_5420);
nor U5853 (N_5853,N_5535,N_5629);
or U5854 (N_5854,N_5416,N_5519);
nor U5855 (N_5855,N_5475,N_5444);
or U5856 (N_5856,N_5665,N_5438);
and U5857 (N_5857,N_5637,N_5695);
xnor U5858 (N_5858,N_5501,N_5584);
xor U5859 (N_5859,N_5429,N_5650);
xor U5860 (N_5860,N_5429,N_5651);
and U5861 (N_5861,N_5693,N_5524);
or U5862 (N_5862,N_5585,N_5484);
nor U5863 (N_5863,N_5661,N_5456);
nor U5864 (N_5864,N_5580,N_5426);
nand U5865 (N_5865,N_5404,N_5465);
nand U5866 (N_5866,N_5488,N_5649);
and U5867 (N_5867,N_5612,N_5608);
nand U5868 (N_5868,N_5487,N_5531);
nand U5869 (N_5869,N_5640,N_5634);
and U5870 (N_5870,N_5488,N_5493);
xor U5871 (N_5871,N_5463,N_5454);
xnor U5872 (N_5872,N_5482,N_5667);
nor U5873 (N_5873,N_5459,N_5511);
nor U5874 (N_5874,N_5437,N_5581);
and U5875 (N_5875,N_5609,N_5406);
nand U5876 (N_5876,N_5643,N_5422);
xor U5877 (N_5877,N_5460,N_5465);
nand U5878 (N_5878,N_5518,N_5459);
nor U5879 (N_5879,N_5680,N_5581);
or U5880 (N_5880,N_5555,N_5448);
and U5881 (N_5881,N_5412,N_5615);
nor U5882 (N_5882,N_5483,N_5541);
nand U5883 (N_5883,N_5699,N_5578);
or U5884 (N_5884,N_5638,N_5539);
nand U5885 (N_5885,N_5660,N_5419);
nor U5886 (N_5886,N_5684,N_5601);
nand U5887 (N_5887,N_5562,N_5498);
nand U5888 (N_5888,N_5421,N_5502);
and U5889 (N_5889,N_5422,N_5509);
and U5890 (N_5890,N_5679,N_5618);
xnor U5891 (N_5891,N_5594,N_5485);
xor U5892 (N_5892,N_5615,N_5639);
or U5893 (N_5893,N_5589,N_5624);
nand U5894 (N_5894,N_5586,N_5465);
xor U5895 (N_5895,N_5537,N_5516);
xnor U5896 (N_5896,N_5502,N_5460);
nand U5897 (N_5897,N_5476,N_5680);
or U5898 (N_5898,N_5694,N_5489);
xnor U5899 (N_5899,N_5609,N_5529);
xor U5900 (N_5900,N_5599,N_5632);
or U5901 (N_5901,N_5508,N_5674);
and U5902 (N_5902,N_5691,N_5441);
and U5903 (N_5903,N_5560,N_5477);
and U5904 (N_5904,N_5655,N_5419);
or U5905 (N_5905,N_5697,N_5673);
or U5906 (N_5906,N_5603,N_5638);
and U5907 (N_5907,N_5654,N_5409);
xor U5908 (N_5908,N_5592,N_5417);
nand U5909 (N_5909,N_5438,N_5625);
nor U5910 (N_5910,N_5667,N_5625);
and U5911 (N_5911,N_5524,N_5641);
nor U5912 (N_5912,N_5596,N_5439);
nor U5913 (N_5913,N_5629,N_5421);
nand U5914 (N_5914,N_5682,N_5558);
or U5915 (N_5915,N_5403,N_5608);
xnor U5916 (N_5916,N_5649,N_5686);
nand U5917 (N_5917,N_5572,N_5431);
or U5918 (N_5918,N_5618,N_5552);
and U5919 (N_5919,N_5699,N_5648);
nand U5920 (N_5920,N_5510,N_5409);
and U5921 (N_5921,N_5638,N_5570);
xnor U5922 (N_5922,N_5460,N_5547);
or U5923 (N_5923,N_5645,N_5582);
nor U5924 (N_5924,N_5540,N_5414);
xnor U5925 (N_5925,N_5409,N_5612);
or U5926 (N_5926,N_5414,N_5632);
nand U5927 (N_5927,N_5433,N_5649);
xor U5928 (N_5928,N_5419,N_5556);
and U5929 (N_5929,N_5578,N_5599);
xnor U5930 (N_5930,N_5446,N_5654);
or U5931 (N_5931,N_5453,N_5468);
nand U5932 (N_5932,N_5498,N_5648);
nor U5933 (N_5933,N_5621,N_5557);
or U5934 (N_5934,N_5468,N_5542);
nor U5935 (N_5935,N_5585,N_5643);
or U5936 (N_5936,N_5484,N_5586);
xor U5937 (N_5937,N_5665,N_5609);
nand U5938 (N_5938,N_5586,N_5635);
or U5939 (N_5939,N_5633,N_5519);
or U5940 (N_5940,N_5545,N_5480);
xnor U5941 (N_5941,N_5487,N_5423);
nand U5942 (N_5942,N_5415,N_5433);
and U5943 (N_5943,N_5492,N_5488);
xnor U5944 (N_5944,N_5633,N_5439);
nor U5945 (N_5945,N_5444,N_5431);
nor U5946 (N_5946,N_5467,N_5509);
nand U5947 (N_5947,N_5500,N_5532);
or U5948 (N_5948,N_5539,N_5435);
xor U5949 (N_5949,N_5666,N_5453);
nor U5950 (N_5950,N_5425,N_5442);
xnor U5951 (N_5951,N_5415,N_5669);
and U5952 (N_5952,N_5463,N_5535);
xnor U5953 (N_5953,N_5687,N_5670);
or U5954 (N_5954,N_5454,N_5435);
xor U5955 (N_5955,N_5668,N_5573);
or U5956 (N_5956,N_5629,N_5664);
nor U5957 (N_5957,N_5656,N_5578);
and U5958 (N_5958,N_5606,N_5453);
nor U5959 (N_5959,N_5664,N_5433);
or U5960 (N_5960,N_5647,N_5554);
nor U5961 (N_5961,N_5427,N_5486);
xor U5962 (N_5962,N_5587,N_5600);
or U5963 (N_5963,N_5417,N_5513);
or U5964 (N_5964,N_5532,N_5540);
nand U5965 (N_5965,N_5556,N_5541);
nor U5966 (N_5966,N_5614,N_5631);
nand U5967 (N_5967,N_5593,N_5422);
nand U5968 (N_5968,N_5456,N_5566);
nand U5969 (N_5969,N_5571,N_5511);
nor U5970 (N_5970,N_5420,N_5593);
or U5971 (N_5971,N_5479,N_5585);
xnor U5972 (N_5972,N_5632,N_5543);
or U5973 (N_5973,N_5492,N_5474);
or U5974 (N_5974,N_5400,N_5571);
nand U5975 (N_5975,N_5679,N_5653);
nand U5976 (N_5976,N_5674,N_5689);
xnor U5977 (N_5977,N_5447,N_5489);
xnor U5978 (N_5978,N_5593,N_5461);
nand U5979 (N_5979,N_5554,N_5425);
or U5980 (N_5980,N_5577,N_5526);
or U5981 (N_5981,N_5528,N_5578);
or U5982 (N_5982,N_5618,N_5687);
xor U5983 (N_5983,N_5525,N_5448);
nand U5984 (N_5984,N_5420,N_5605);
xnor U5985 (N_5985,N_5468,N_5494);
nand U5986 (N_5986,N_5632,N_5475);
or U5987 (N_5987,N_5531,N_5546);
nand U5988 (N_5988,N_5684,N_5540);
nor U5989 (N_5989,N_5465,N_5570);
nand U5990 (N_5990,N_5507,N_5635);
nor U5991 (N_5991,N_5440,N_5461);
and U5992 (N_5992,N_5632,N_5535);
nor U5993 (N_5993,N_5663,N_5557);
and U5994 (N_5994,N_5654,N_5430);
and U5995 (N_5995,N_5663,N_5623);
nor U5996 (N_5996,N_5667,N_5600);
or U5997 (N_5997,N_5643,N_5400);
xnor U5998 (N_5998,N_5456,N_5556);
or U5999 (N_5999,N_5601,N_5566);
nand U6000 (N_6000,N_5931,N_5818);
or U6001 (N_6001,N_5802,N_5760);
nand U6002 (N_6002,N_5934,N_5959);
nor U6003 (N_6003,N_5814,N_5913);
and U6004 (N_6004,N_5797,N_5982);
or U6005 (N_6005,N_5891,N_5892);
xnor U6006 (N_6006,N_5904,N_5919);
and U6007 (N_6007,N_5878,N_5958);
and U6008 (N_6008,N_5908,N_5826);
xor U6009 (N_6009,N_5999,N_5733);
and U6010 (N_6010,N_5823,N_5924);
and U6011 (N_6011,N_5949,N_5994);
nand U6012 (N_6012,N_5922,N_5977);
or U6013 (N_6013,N_5819,N_5955);
xor U6014 (N_6014,N_5881,N_5722);
and U6015 (N_6015,N_5875,N_5824);
nor U6016 (N_6016,N_5727,N_5979);
or U6017 (N_6017,N_5796,N_5937);
or U6018 (N_6018,N_5846,N_5854);
or U6019 (N_6019,N_5858,N_5912);
or U6020 (N_6020,N_5728,N_5809);
nor U6021 (N_6021,N_5871,N_5963);
or U6022 (N_6022,N_5960,N_5843);
nor U6023 (N_6023,N_5750,N_5723);
nand U6024 (N_6024,N_5765,N_5896);
and U6025 (N_6025,N_5869,N_5948);
nand U6026 (N_6026,N_5753,N_5838);
and U6027 (N_6027,N_5942,N_5707);
and U6028 (N_6028,N_5724,N_5840);
xnor U6029 (N_6029,N_5860,N_5917);
nand U6030 (N_6030,N_5777,N_5983);
nor U6031 (N_6031,N_5830,N_5947);
and U6032 (N_6032,N_5730,N_5956);
nand U6033 (N_6033,N_5746,N_5738);
nor U6034 (N_6034,N_5754,N_5817);
nand U6035 (N_6035,N_5801,N_5714);
nand U6036 (N_6036,N_5886,N_5778);
nand U6037 (N_6037,N_5927,N_5907);
nand U6038 (N_6038,N_5720,N_5769);
or U6039 (N_6039,N_5758,N_5897);
xor U6040 (N_6040,N_5737,N_5872);
or U6041 (N_6041,N_5943,N_5713);
and U6042 (N_6042,N_5916,N_5807);
or U6043 (N_6043,N_5864,N_5879);
xnor U6044 (N_6044,N_5829,N_5990);
nor U6045 (N_6045,N_5828,N_5800);
xnor U6046 (N_6046,N_5899,N_5832);
xnor U6047 (N_6047,N_5716,N_5841);
xor U6048 (N_6048,N_5747,N_5873);
nor U6049 (N_6049,N_5839,N_5740);
nand U6050 (N_6050,N_5988,N_5836);
or U6051 (N_6051,N_5755,N_5941);
and U6052 (N_6052,N_5783,N_5835);
nand U6053 (N_6053,N_5966,N_5772);
nor U6054 (N_6054,N_5771,N_5751);
xnor U6055 (N_6055,N_5709,N_5885);
nor U6056 (N_6056,N_5876,N_5993);
xor U6057 (N_6057,N_5935,N_5757);
xor U6058 (N_6058,N_5770,N_5877);
or U6059 (N_6059,N_5790,N_5852);
or U6060 (N_6060,N_5779,N_5706);
and U6061 (N_6061,N_5773,N_5940);
xnor U6062 (N_6062,N_5861,N_5785);
or U6063 (N_6063,N_5782,N_5710);
and U6064 (N_6064,N_5853,N_5976);
nor U6065 (N_6065,N_5788,N_5822);
xor U6066 (N_6066,N_5890,N_5793);
or U6067 (N_6067,N_5857,N_5813);
nor U6068 (N_6068,N_5923,N_5974);
nand U6069 (N_6069,N_5887,N_5991);
or U6070 (N_6070,N_5969,N_5766);
or U6071 (N_6071,N_5911,N_5909);
and U6072 (N_6072,N_5957,N_5933);
and U6073 (N_6073,N_5902,N_5702);
or U6074 (N_6074,N_5711,N_5980);
xor U6075 (N_6075,N_5811,N_5978);
and U6076 (N_6076,N_5816,N_5821);
or U6077 (N_6077,N_5717,N_5996);
and U6078 (N_6078,N_5831,N_5851);
and U6079 (N_6079,N_5845,N_5950);
nand U6080 (N_6080,N_5764,N_5705);
nor U6081 (N_6081,N_5918,N_5930);
and U6082 (N_6082,N_5973,N_5898);
nand U6083 (N_6083,N_5774,N_5736);
nor U6084 (N_6084,N_5856,N_5944);
and U6085 (N_6085,N_5964,N_5834);
nor U6086 (N_6086,N_5812,N_5731);
or U6087 (N_6087,N_5929,N_5992);
or U6088 (N_6088,N_5847,N_5715);
nand U6089 (N_6089,N_5744,N_5926);
nand U6090 (N_6090,N_5905,N_5745);
and U6091 (N_6091,N_5789,N_5882);
nor U6092 (N_6092,N_5925,N_5849);
nand U6093 (N_6093,N_5863,N_5749);
xnor U6094 (N_6094,N_5921,N_5844);
nor U6095 (N_6095,N_5884,N_5954);
xnor U6096 (N_6096,N_5920,N_5915);
xnor U6097 (N_6097,N_5932,N_5748);
or U6098 (N_6098,N_5981,N_5708);
xor U6099 (N_6099,N_5704,N_5741);
nor U6100 (N_6100,N_5791,N_5971);
nand U6101 (N_6101,N_5725,N_5967);
or U6102 (N_6102,N_5756,N_5804);
and U6103 (N_6103,N_5910,N_5961);
nor U6104 (N_6104,N_5894,N_5968);
and U6105 (N_6105,N_5984,N_5742);
or U6106 (N_6106,N_5763,N_5700);
xnor U6107 (N_6107,N_5936,N_5953);
or U6108 (N_6108,N_5743,N_5712);
xor U6109 (N_6109,N_5972,N_5732);
or U6110 (N_6110,N_5719,N_5928);
xor U6111 (N_6111,N_5799,N_5952);
and U6112 (N_6112,N_5965,N_5867);
or U6113 (N_6113,N_5989,N_5951);
xor U6114 (N_6114,N_5850,N_5775);
and U6115 (N_6115,N_5975,N_5970);
and U6116 (N_6116,N_5833,N_5866);
or U6117 (N_6117,N_5718,N_5806);
or U6118 (N_6118,N_5842,N_5781);
or U6119 (N_6119,N_5998,N_5768);
and U6120 (N_6120,N_5985,N_5946);
or U6121 (N_6121,N_5729,N_5792);
xor U6122 (N_6122,N_5855,N_5862);
xnor U6123 (N_6123,N_5986,N_5987);
nand U6124 (N_6124,N_5808,N_5805);
nor U6125 (N_6125,N_5787,N_5895);
nor U6126 (N_6126,N_5889,N_5815);
xor U6127 (N_6127,N_5739,N_5767);
or U6128 (N_6128,N_5762,N_5734);
or U6129 (N_6129,N_5945,N_5752);
nor U6130 (N_6130,N_5914,N_5721);
nand U6131 (N_6131,N_5900,N_5893);
xor U6132 (N_6132,N_5865,N_5848);
or U6133 (N_6133,N_5803,N_5735);
and U6134 (N_6134,N_5780,N_5938);
or U6135 (N_6135,N_5995,N_5880);
or U6136 (N_6136,N_5776,N_5701);
nand U6137 (N_6137,N_5874,N_5939);
or U6138 (N_6138,N_5883,N_5726);
xor U6139 (N_6139,N_5859,N_5903);
nor U6140 (N_6140,N_5795,N_5962);
xnor U6141 (N_6141,N_5810,N_5825);
nor U6142 (N_6142,N_5786,N_5798);
nor U6143 (N_6143,N_5870,N_5906);
nor U6144 (N_6144,N_5827,N_5901);
xnor U6145 (N_6145,N_5784,N_5997);
and U6146 (N_6146,N_5761,N_5794);
and U6147 (N_6147,N_5820,N_5759);
nor U6148 (N_6148,N_5868,N_5837);
xnor U6149 (N_6149,N_5703,N_5888);
nor U6150 (N_6150,N_5850,N_5854);
nand U6151 (N_6151,N_5885,N_5950);
or U6152 (N_6152,N_5884,N_5811);
xnor U6153 (N_6153,N_5941,N_5810);
or U6154 (N_6154,N_5929,N_5738);
and U6155 (N_6155,N_5763,N_5789);
nand U6156 (N_6156,N_5771,N_5862);
nor U6157 (N_6157,N_5969,N_5990);
and U6158 (N_6158,N_5784,N_5798);
nand U6159 (N_6159,N_5800,N_5945);
nand U6160 (N_6160,N_5796,N_5832);
nor U6161 (N_6161,N_5814,N_5835);
nand U6162 (N_6162,N_5930,N_5917);
and U6163 (N_6163,N_5889,N_5741);
or U6164 (N_6164,N_5996,N_5882);
or U6165 (N_6165,N_5817,N_5988);
xnor U6166 (N_6166,N_5863,N_5753);
nor U6167 (N_6167,N_5733,N_5889);
nor U6168 (N_6168,N_5897,N_5718);
and U6169 (N_6169,N_5778,N_5898);
and U6170 (N_6170,N_5912,N_5948);
nand U6171 (N_6171,N_5800,N_5757);
nor U6172 (N_6172,N_5768,N_5762);
and U6173 (N_6173,N_5829,N_5801);
or U6174 (N_6174,N_5930,N_5947);
nand U6175 (N_6175,N_5773,N_5961);
nor U6176 (N_6176,N_5705,N_5817);
xor U6177 (N_6177,N_5744,N_5905);
nand U6178 (N_6178,N_5707,N_5884);
xor U6179 (N_6179,N_5957,N_5862);
or U6180 (N_6180,N_5903,N_5799);
nand U6181 (N_6181,N_5975,N_5797);
or U6182 (N_6182,N_5873,N_5733);
nand U6183 (N_6183,N_5973,N_5870);
and U6184 (N_6184,N_5860,N_5720);
or U6185 (N_6185,N_5827,N_5909);
nor U6186 (N_6186,N_5767,N_5761);
or U6187 (N_6187,N_5731,N_5866);
nor U6188 (N_6188,N_5811,N_5908);
and U6189 (N_6189,N_5937,N_5992);
and U6190 (N_6190,N_5888,N_5870);
nand U6191 (N_6191,N_5725,N_5972);
nor U6192 (N_6192,N_5796,N_5786);
nor U6193 (N_6193,N_5981,N_5821);
nor U6194 (N_6194,N_5849,N_5892);
nand U6195 (N_6195,N_5953,N_5781);
or U6196 (N_6196,N_5898,N_5922);
nand U6197 (N_6197,N_5979,N_5815);
or U6198 (N_6198,N_5887,N_5819);
and U6199 (N_6199,N_5834,N_5741);
nor U6200 (N_6200,N_5844,N_5996);
or U6201 (N_6201,N_5729,N_5773);
and U6202 (N_6202,N_5957,N_5730);
nor U6203 (N_6203,N_5758,N_5723);
or U6204 (N_6204,N_5954,N_5710);
and U6205 (N_6205,N_5780,N_5925);
and U6206 (N_6206,N_5791,N_5943);
nand U6207 (N_6207,N_5762,N_5952);
or U6208 (N_6208,N_5997,N_5780);
xor U6209 (N_6209,N_5978,N_5832);
nor U6210 (N_6210,N_5870,N_5875);
nand U6211 (N_6211,N_5850,N_5720);
and U6212 (N_6212,N_5932,N_5938);
nand U6213 (N_6213,N_5828,N_5722);
or U6214 (N_6214,N_5731,N_5950);
or U6215 (N_6215,N_5963,N_5714);
or U6216 (N_6216,N_5990,N_5938);
and U6217 (N_6217,N_5970,N_5883);
and U6218 (N_6218,N_5971,N_5913);
xnor U6219 (N_6219,N_5824,N_5990);
and U6220 (N_6220,N_5758,N_5839);
nand U6221 (N_6221,N_5775,N_5988);
or U6222 (N_6222,N_5897,N_5986);
xor U6223 (N_6223,N_5876,N_5921);
nand U6224 (N_6224,N_5803,N_5824);
nor U6225 (N_6225,N_5905,N_5892);
or U6226 (N_6226,N_5908,N_5794);
or U6227 (N_6227,N_5964,N_5898);
nand U6228 (N_6228,N_5783,N_5825);
nor U6229 (N_6229,N_5851,N_5791);
xnor U6230 (N_6230,N_5831,N_5850);
xnor U6231 (N_6231,N_5779,N_5940);
and U6232 (N_6232,N_5933,N_5716);
and U6233 (N_6233,N_5979,N_5820);
and U6234 (N_6234,N_5860,N_5876);
nand U6235 (N_6235,N_5775,N_5832);
nand U6236 (N_6236,N_5766,N_5973);
and U6237 (N_6237,N_5887,N_5794);
or U6238 (N_6238,N_5805,N_5884);
or U6239 (N_6239,N_5785,N_5923);
xor U6240 (N_6240,N_5769,N_5790);
xor U6241 (N_6241,N_5876,N_5928);
xnor U6242 (N_6242,N_5952,N_5918);
nand U6243 (N_6243,N_5860,N_5979);
xnor U6244 (N_6244,N_5964,N_5780);
xnor U6245 (N_6245,N_5820,N_5775);
or U6246 (N_6246,N_5943,N_5956);
nand U6247 (N_6247,N_5895,N_5842);
or U6248 (N_6248,N_5753,N_5709);
nand U6249 (N_6249,N_5836,N_5753);
and U6250 (N_6250,N_5869,N_5730);
nand U6251 (N_6251,N_5711,N_5775);
nand U6252 (N_6252,N_5994,N_5964);
nor U6253 (N_6253,N_5875,N_5780);
or U6254 (N_6254,N_5808,N_5897);
nand U6255 (N_6255,N_5769,N_5805);
nand U6256 (N_6256,N_5984,N_5923);
nand U6257 (N_6257,N_5971,N_5922);
nand U6258 (N_6258,N_5832,N_5867);
or U6259 (N_6259,N_5765,N_5700);
nor U6260 (N_6260,N_5769,N_5751);
and U6261 (N_6261,N_5951,N_5997);
and U6262 (N_6262,N_5756,N_5897);
nor U6263 (N_6263,N_5881,N_5798);
and U6264 (N_6264,N_5913,N_5828);
xor U6265 (N_6265,N_5863,N_5800);
xor U6266 (N_6266,N_5977,N_5885);
xnor U6267 (N_6267,N_5763,N_5999);
or U6268 (N_6268,N_5952,N_5706);
or U6269 (N_6269,N_5725,N_5973);
nand U6270 (N_6270,N_5999,N_5933);
or U6271 (N_6271,N_5942,N_5732);
nand U6272 (N_6272,N_5890,N_5756);
nand U6273 (N_6273,N_5885,N_5994);
nand U6274 (N_6274,N_5882,N_5978);
nor U6275 (N_6275,N_5815,N_5973);
or U6276 (N_6276,N_5942,N_5915);
nand U6277 (N_6277,N_5977,N_5786);
xnor U6278 (N_6278,N_5800,N_5929);
nand U6279 (N_6279,N_5724,N_5813);
nor U6280 (N_6280,N_5841,N_5712);
xnor U6281 (N_6281,N_5803,N_5994);
nor U6282 (N_6282,N_5947,N_5895);
and U6283 (N_6283,N_5970,N_5735);
nor U6284 (N_6284,N_5929,N_5912);
and U6285 (N_6285,N_5753,N_5825);
and U6286 (N_6286,N_5860,N_5948);
xor U6287 (N_6287,N_5896,N_5934);
xnor U6288 (N_6288,N_5910,N_5711);
or U6289 (N_6289,N_5778,N_5922);
and U6290 (N_6290,N_5854,N_5745);
nand U6291 (N_6291,N_5843,N_5894);
nor U6292 (N_6292,N_5768,N_5737);
or U6293 (N_6293,N_5706,N_5947);
xnor U6294 (N_6294,N_5703,N_5813);
and U6295 (N_6295,N_5911,N_5786);
xnor U6296 (N_6296,N_5985,N_5943);
and U6297 (N_6297,N_5740,N_5702);
and U6298 (N_6298,N_5914,N_5750);
or U6299 (N_6299,N_5981,N_5700);
and U6300 (N_6300,N_6038,N_6268);
or U6301 (N_6301,N_6061,N_6075);
nand U6302 (N_6302,N_6050,N_6086);
xor U6303 (N_6303,N_6287,N_6157);
nand U6304 (N_6304,N_6149,N_6035);
and U6305 (N_6305,N_6021,N_6181);
xor U6306 (N_6306,N_6285,N_6183);
xor U6307 (N_6307,N_6024,N_6293);
and U6308 (N_6308,N_6116,N_6148);
or U6309 (N_6309,N_6093,N_6191);
and U6310 (N_6310,N_6058,N_6256);
nor U6311 (N_6311,N_6074,N_6135);
xor U6312 (N_6312,N_6274,N_6254);
nor U6313 (N_6313,N_6132,N_6003);
nand U6314 (N_6314,N_6062,N_6138);
nand U6315 (N_6315,N_6053,N_6124);
or U6316 (N_6316,N_6097,N_6155);
and U6317 (N_6317,N_6039,N_6104);
nand U6318 (N_6318,N_6222,N_6223);
xnor U6319 (N_6319,N_6220,N_6156);
nor U6320 (N_6320,N_6275,N_6008);
nand U6321 (N_6321,N_6142,N_6173);
nand U6322 (N_6322,N_6091,N_6016);
xor U6323 (N_6323,N_6214,N_6203);
nor U6324 (N_6324,N_6296,N_6154);
xnor U6325 (N_6325,N_6001,N_6144);
nor U6326 (N_6326,N_6013,N_6204);
and U6327 (N_6327,N_6052,N_6202);
and U6328 (N_6328,N_6297,N_6047);
xnor U6329 (N_6329,N_6270,N_6169);
nor U6330 (N_6330,N_6034,N_6215);
and U6331 (N_6331,N_6007,N_6247);
xor U6332 (N_6332,N_6068,N_6098);
nor U6333 (N_6333,N_6289,N_6229);
nor U6334 (N_6334,N_6137,N_6162);
and U6335 (N_6335,N_6283,N_6070);
xor U6336 (N_6336,N_6272,N_6071);
nand U6337 (N_6337,N_6010,N_6037);
xor U6338 (N_6338,N_6252,N_6267);
nor U6339 (N_6339,N_6081,N_6226);
xnor U6340 (N_6340,N_6251,N_6193);
xor U6341 (N_6341,N_6205,N_6103);
and U6342 (N_6342,N_6244,N_6206);
xor U6343 (N_6343,N_6069,N_6029);
nor U6344 (N_6344,N_6151,N_6101);
or U6345 (N_6345,N_6082,N_6042);
nor U6346 (N_6346,N_6133,N_6192);
nand U6347 (N_6347,N_6266,N_6235);
nor U6348 (N_6348,N_6108,N_6243);
xnor U6349 (N_6349,N_6210,N_6140);
nor U6350 (N_6350,N_6022,N_6134);
xor U6351 (N_6351,N_6245,N_6117);
nor U6352 (N_6352,N_6129,N_6072);
or U6353 (N_6353,N_6253,N_6189);
xnor U6354 (N_6354,N_6041,N_6028);
xnor U6355 (N_6355,N_6088,N_6218);
or U6356 (N_6356,N_6127,N_6168);
xor U6357 (N_6357,N_6237,N_6176);
xor U6358 (N_6358,N_6002,N_6241);
and U6359 (N_6359,N_6248,N_6278);
and U6360 (N_6360,N_6049,N_6015);
and U6361 (N_6361,N_6113,N_6121);
and U6362 (N_6362,N_6294,N_6044);
or U6363 (N_6363,N_6064,N_6171);
nand U6364 (N_6364,N_6186,N_6126);
xor U6365 (N_6365,N_6230,N_6195);
or U6366 (N_6366,N_6115,N_6281);
xor U6367 (N_6367,N_6051,N_6128);
and U6368 (N_6368,N_6153,N_6045);
nor U6369 (N_6369,N_6290,N_6182);
nor U6370 (N_6370,N_6284,N_6054);
and U6371 (N_6371,N_6262,N_6299);
nand U6372 (N_6372,N_6141,N_6260);
nor U6373 (N_6373,N_6136,N_6221);
and U6374 (N_6374,N_6087,N_6099);
xor U6375 (N_6375,N_6282,N_6031);
or U6376 (N_6376,N_6250,N_6219);
xnor U6377 (N_6377,N_6213,N_6158);
nor U6378 (N_6378,N_6083,N_6159);
nor U6379 (N_6379,N_6032,N_6056);
xnor U6380 (N_6380,N_6179,N_6009);
nand U6381 (N_6381,N_6152,N_6277);
xnor U6382 (N_6382,N_6125,N_6123);
nor U6383 (N_6383,N_6232,N_6036);
nor U6384 (N_6384,N_6231,N_6177);
nor U6385 (N_6385,N_6018,N_6165);
and U6386 (N_6386,N_6295,N_6060);
or U6387 (N_6387,N_6067,N_6200);
or U6388 (N_6388,N_6109,N_6017);
or U6389 (N_6389,N_6106,N_6263);
and U6390 (N_6390,N_6030,N_6238);
xnor U6391 (N_6391,N_6092,N_6242);
nand U6392 (N_6392,N_6261,N_6163);
nor U6393 (N_6393,N_6265,N_6096);
nor U6394 (N_6394,N_6240,N_6094);
nor U6395 (N_6395,N_6014,N_6019);
nand U6396 (N_6396,N_6286,N_6199);
or U6397 (N_6397,N_6178,N_6227);
or U6398 (N_6398,N_6174,N_6066);
and U6399 (N_6399,N_6276,N_6194);
and U6400 (N_6400,N_6201,N_6105);
or U6401 (N_6401,N_6279,N_6209);
and U6402 (N_6402,N_6160,N_6122);
nor U6403 (N_6403,N_6043,N_6023);
nor U6404 (N_6404,N_6184,N_6234);
or U6405 (N_6405,N_6107,N_6216);
xnor U6406 (N_6406,N_6167,N_6118);
and U6407 (N_6407,N_6188,N_6273);
and U6408 (N_6408,N_6217,N_6080);
xnor U6409 (N_6409,N_6076,N_6059);
xnor U6410 (N_6410,N_6057,N_6264);
and U6411 (N_6411,N_6012,N_6233);
nor U6412 (N_6412,N_6288,N_6084);
and U6413 (N_6413,N_6026,N_6114);
or U6414 (N_6414,N_6175,N_6020);
or U6415 (N_6415,N_6090,N_6257);
nor U6416 (N_6416,N_6190,N_6258);
nand U6417 (N_6417,N_6033,N_6185);
nand U6418 (N_6418,N_6187,N_6004);
or U6419 (N_6419,N_6291,N_6078);
and U6420 (N_6420,N_6147,N_6046);
or U6421 (N_6421,N_6100,N_6280);
or U6422 (N_6422,N_6102,N_6063);
or U6423 (N_6423,N_6079,N_6211);
nor U6424 (N_6424,N_6271,N_6298);
nand U6425 (N_6425,N_6139,N_6172);
nand U6426 (N_6426,N_6198,N_6110);
nor U6427 (N_6427,N_6208,N_6228);
or U6428 (N_6428,N_6055,N_6249);
xnor U6429 (N_6429,N_6207,N_6000);
nand U6430 (N_6430,N_6089,N_6170);
and U6431 (N_6431,N_6027,N_6077);
and U6432 (N_6432,N_6150,N_6145);
nor U6433 (N_6433,N_6006,N_6025);
and U6434 (N_6434,N_6146,N_6292);
xor U6435 (N_6435,N_6259,N_6005);
or U6436 (N_6436,N_6225,N_6236);
or U6437 (N_6437,N_6112,N_6120);
xnor U6438 (N_6438,N_6166,N_6224);
nor U6439 (N_6439,N_6164,N_6197);
and U6440 (N_6440,N_6239,N_6119);
or U6441 (N_6441,N_6095,N_6073);
nand U6442 (N_6442,N_6143,N_6212);
or U6443 (N_6443,N_6085,N_6111);
nor U6444 (N_6444,N_6130,N_6131);
or U6445 (N_6445,N_6246,N_6255);
nand U6446 (N_6446,N_6161,N_6011);
nor U6447 (N_6447,N_6196,N_6180);
or U6448 (N_6448,N_6065,N_6048);
nor U6449 (N_6449,N_6040,N_6269);
nand U6450 (N_6450,N_6055,N_6035);
nor U6451 (N_6451,N_6114,N_6225);
xor U6452 (N_6452,N_6203,N_6028);
nor U6453 (N_6453,N_6211,N_6062);
xor U6454 (N_6454,N_6293,N_6135);
and U6455 (N_6455,N_6047,N_6052);
nand U6456 (N_6456,N_6298,N_6237);
and U6457 (N_6457,N_6167,N_6160);
or U6458 (N_6458,N_6058,N_6219);
or U6459 (N_6459,N_6204,N_6032);
nand U6460 (N_6460,N_6081,N_6032);
nand U6461 (N_6461,N_6228,N_6062);
xor U6462 (N_6462,N_6111,N_6266);
nand U6463 (N_6463,N_6045,N_6247);
nor U6464 (N_6464,N_6090,N_6028);
and U6465 (N_6465,N_6238,N_6268);
nand U6466 (N_6466,N_6242,N_6173);
or U6467 (N_6467,N_6035,N_6059);
or U6468 (N_6468,N_6127,N_6215);
nor U6469 (N_6469,N_6159,N_6243);
or U6470 (N_6470,N_6017,N_6296);
nand U6471 (N_6471,N_6106,N_6269);
and U6472 (N_6472,N_6017,N_6148);
and U6473 (N_6473,N_6111,N_6120);
nand U6474 (N_6474,N_6170,N_6071);
and U6475 (N_6475,N_6259,N_6134);
xnor U6476 (N_6476,N_6208,N_6160);
xnor U6477 (N_6477,N_6021,N_6078);
xor U6478 (N_6478,N_6064,N_6024);
and U6479 (N_6479,N_6185,N_6244);
xor U6480 (N_6480,N_6025,N_6009);
xor U6481 (N_6481,N_6152,N_6017);
xor U6482 (N_6482,N_6128,N_6168);
or U6483 (N_6483,N_6289,N_6157);
or U6484 (N_6484,N_6286,N_6026);
nand U6485 (N_6485,N_6128,N_6039);
xnor U6486 (N_6486,N_6280,N_6030);
nor U6487 (N_6487,N_6191,N_6282);
and U6488 (N_6488,N_6030,N_6108);
nor U6489 (N_6489,N_6292,N_6018);
and U6490 (N_6490,N_6203,N_6171);
nand U6491 (N_6491,N_6073,N_6040);
or U6492 (N_6492,N_6018,N_6219);
or U6493 (N_6493,N_6069,N_6297);
and U6494 (N_6494,N_6098,N_6263);
xor U6495 (N_6495,N_6229,N_6110);
xnor U6496 (N_6496,N_6001,N_6116);
nand U6497 (N_6497,N_6166,N_6004);
and U6498 (N_6498,N_6139,N_6237);
xor U6499 (N_6499,N_6205,N_6028);
and U6500 (N_6500,N_6058,N_6008);
or U6501 (N_6501,N_6045,N_6147);
xnor U6502 (N_6502,N_6100,N_6199);
xor U6503 (N_6503,N_6058,N_6112);
xor U6504 (N_6504,N_6141,N_6211);
nand U6505 (N_6505,N_6122,N_6043);
nor U6506 (N_6506,N_6216,N_6059);
nand U6507 (N_6507,N_6111,N_6170);
xnor U6508 (N_6508,N_6258,N_6092);
or U6509 (N_6509,N_6223,N_6276);
or U6510 (N_6510,N_6186,N_6057);
xor U6511 (N_6511,N_6079,N_6053);
nand U6512 (N_6512,N_6168,N_6268);
xnor U6513 (N_6513,N_6116,N_6204);
and U6514 (N_6514,N_6270,N_6005);
xnor U6515 (N_6515,N_6299,N_6291);
and U6516 (N_6516,N_6240,N_6117);
and U6517 (N_6517,N_6074,N_6077);
and U6518 (N_6518,N_6186,N_6103);
and U6519 (N_6519,N_6100,N_6037);
and U6520 (N_6520,N_6096,N_6072);
nor U6521 (N_6521,N_6035,N_6148);
nor U6522 (N_6522,N_6296,N_6094);
nand U6523 (N_6523,N_6105,N_6101);
or U6524 (N_6524,N_6227,N_6193);
or U6525 (N_6525,N_6036,N_6293);
nor U6526 (N_6526,N_6207,N_6155);
and U6527 (N_6527,N_6052,N_6088);
or U6528 (N_6528,N_6214,N_6001);
and U6529 (N_6529,N_6211,N_6264);
and U6530 (N_6530,N_6203,N_6240);
nand U6531 (N_6531,N_6144,N_6241);
nor U6532 (N_6532,N_6033,N_6148);
and U6533 (N_6533,N_6067,N_6170);
nor U6534 (N_6534,N_6152,N_6224);
nand U6535 (N_6535,N_6083,N_6133);
and U6536 (N_6536,N_6121,N_6163);
or U6537 (N_6537,N_6263,N_6094);
nand U6538 (N_6538,N_6244,N_6060);
nor U6539 (N_6539,N_6174,N_6043);
nor U6540 (N_6540,N_6053,N_6208);
nor U6541 (N_6541,N_6258,N_6024);
nand U6542 (N_6542,N_6217,N_6142);
and U6543 (N_6543,N_6070,N_6159);
and U6544 (N_6544,N_6155,N_6095);
or U6545 (N_6545,N_6202,N_6257);
and U6546 (N_6546,N_6090,N_6009);
and U6547 (N_6547,N_6012,N_6122);
nand U6548 (N_6548,N_6092,N_6137);
and U6549 (N_6549,N_6216,N_6139);
nor U6550 (N_6550,N_6292,N_6285);
nor U6551 (N_6551,N_6224,N_6031);
and U6552 (N_6552,N_6151,N_6212);
xnor U6553 (N_6553,N_6184,N_6132);
nor U6554 (N_6554,N_6132,N_6298);
or U6555 (N_6555,N_6121,N_6062);
nand U6556 (N_6556,N_6203,N_6123);
nor U6557 (N_6557,N_6200,N_6017);
or U6558 (N_6558,N_6161,N_6221);
xor U6559 (N_6559,N_6221,N_6241);
nand U6560 (N_6560,N_6029,N_6278);
nor U6561 (N_6561,N_6140,N_6221);
or U6562 (N_6562,N_6005,N_6107);
and U6563 (N_6563,N_6091,N_6104);
nor U6564 (N_6564,N_6084,N_6018);
nor U6565 (N_6565,N_6169,N_6242);
nor U6566 (N_6566,N_6241,N_6029);
or U6567 (N_6567,N_6111,N_6023);
nor U6568 (N_6568,N_6223,N_6287);
xor U6569 (N_6569,N_6269,N_6179);
or U6570 (N_6570,N_6234,N_6038);
xor U6571 (N_6571,N_6280,N_6194);
nor U6572 (N_6572,N_6240,N_6297);
xnor U6573 (N_6573,N_6153,N_6017);
or U6574 (N_6574,N_6019,N_6186);
or U6575 (N_6575,N_6232,N_6199);
nor U6576 (N_6576,N_6039,N_6232);
xor U6577 (N_6577,N_6196,N_6256);
nand U6578 (N_6578,N_6112,N_6117);
nor U6579 (N_6579,N_6205,N_6280);
xnor U6580 (N_6580,N_6201,N_6092);
xor U6581 (N_6581,N_6204,N_6298);
or U6582 (N_6582,N_6107,N_6070);
nor U6583 (N_6583,N_6112,N_6029);
nor U6584 (N_6584,N_6174,N_6007);
and U6585 (N_6585,N_6043,N_6028);
and U6586 (N_6586,N_6001,N_6052);
and U6587 (N_6587,N_6016,N_6027);
nand U6588 (N_6588,N_6120,N_6114);
and U6589 (N_6589,N_6237,N_6294);
and U6590 (N_6590,N_6258,N_6280);
nand U6591 (N_6591,N_6238,N_6274);
nor U6592 (N_6592,N_6299,N_6110);
nor U6593 (N_6593,N_6281,N_6187);
xnor U6594 (N_6594,N_6139,N_6014);
and U6595 (N_6595,N_6269,N_6049);
nor U6596 (N_6596,N_6219,N_6021);
or U6597 (N_6597,N_6168,N_6239);
xnor U6598 (N_6598,N_6232,N_6117);
nand U6599 (N_6599,N_6058,N_6115);
nand U6600 (N_6600,N_6301,N_6371);
xnor U6601 (N_6601,N_6439,N_6483);
or U6602 (N_6602,N_6537,N_6395);
nand U6603 (N_6603,N_6385,N_6319);
xnor U6604 (N_6604,N_6565,N_6560);
nand U6605 (N_6605,N_6528,N_6356);
nor U6606 (N_6606,N_6538,N_6544);
xnor U6607 (N_6607,N_6346,N_6318);
and U6608 (N_6608,N_6304,N_6479);
nor U6609 (N_6609,N_6530,N_6321);
or U6610 (N_6610,N_6591,N_6521);
and U6611 (N_6611,N_6495,N_6484);
nor U6612 (N_6612,N_6317,N_6442);
nor U6613 (N_6613,N_6396,N_6458);
and U6614 (N_6614,N_6429,N_6461);
xnor U6615 (N_6615,N_6574,N_6335);
xor U6616 (N_6616,N_6588,N_6545);
and U6617 (N_6617,N_6339,N_6333);
and U6618 (N_6618,N_6303,N_6407);
or U6619 (N_6619,N_6502,N_6421);
xnor U6620 (N_6620,N_6307,N_6403);
nor U6621 (N_6621,N_6523,N_6515);
xor U6622 (N_6622,N_6581,N_6388);
nor U6623 (N_6623,N_6448,N_6357);
nand U6624 (N_6624,N_6548,N_6526);
or U6625 (N_6625,N_6587,N_6363);
or U6626 (N_6626,N_6491,N_6367);
and U6627 (N_6627,N_6311,N_6422);
and U6628 (N_6628,N_6480,N_6563);
nor U6629 (N_6629,N_6453,N_6456);
nand U6630 (N_6630,N_6559,N_6500);
and U6631 (N_6631,N_6302,N_6350);
xnor U6632 (N_6632,N_6348,N_6419);
nand U6633 (N_6633,N_6323,N_6532);
xor U6634 (N_6634,N_6341,N_6380);
and U6635 (N_6635,N_6590,N_6330);
nor U6636 (N_6636,N_6576,N_6513);
and U6637 (N_6637,N_6472,N_6462);
or U6638 (N_6638,N_6522,N_6535);
nand U6639 (N_6639,N_6529,N_6313);
or U6640 (N_6640,N_6398,N_6354);
xnor U6641 (N_6641,N_6359,N_6441);
and U6642 (N_6642,N_6362,N_6597);
nor U6643 (N_6643,N_6399,N_6524);
nor U6644 (N_6644,N_6446,N_6437);
xnor U6645 (N_6645,N_6478,N_6579);
and U6646 (N_6646,N_6334,N_6489);
nand U6647 (N_6647,N_6556,N_6583);
and U6648 (N_6648,N_6497,N_6300);
xor U6649 (N_6649,N_6519,N_6487);
xor U6650 (N_6650,N_6410,N_6331);
nand U6651 (N_6651,N_6414,N_6488);
and U6652 (N_6652,N_6316,N_6332);
xor U6653 (N_6653,N_6444,N_6411);
and U6654 (N_6654,N_6546,N_6531);
xnor U6655 (N_6655,N_6562,N_6501);
nor U6656 (N_6656,N_6384,N_6520);
nand U6657 (N_6657,N_6571,N_6584);
xnor U6658 (N_6658,N_6372,N_6402);
nand U6659 (N_6659,N_6492,N_6505);
xnor U6660 (N_6660,N_6568,N_6394);
or U6661 (N_6661,N_6496,N_6432);
and U6662 (N_6662,N_6327,N_6434);
nand U6663 (N_6663,N_6409,N_6309);
nand U6664 (N_6664,N_6310,N_6425);
and U6665 (N_6665,N_6416,N_6338);
and U6666 (N_6666,N_6599,N_6504);
nor U6667 (N_6667,N_6578,N_6585);
or U6668 (N_6668,N_6557,N_6445);
xnor U6669 (N_6669,N_6352,N_6315);
and U6670 (N_6670,N_6469,N_6572);
nor U6671 (N_6671,N_6490,N_6379);
and U6672 (N_6672,N_6598,N_6375);
and U6673 (N_6673,N_6440,N_6549);
nand U6674 (N_6674,N_6471,N_6438);
nand U6675 (N_6675,N_6353,N_6383);
xor U6676 (N_6676,N_6358,N_6465);
or U6677 (N_6677,N_6401,N_6476);
or U6678 (N_6678,N_6326,N_6486);
nor U6679 (N_6679,N_6430,N_6593);
nand U6680 (N_6680,N_6506,N_6539);
nor U6681 (N_6681,N_6594,N_6470);
or U6682 (N_6682,N_6517,N_6328);
nor U6683 (N_6683,N_6423,N_6392);
or U6684 (N_6684,N_6569,N_6455);
or U6685 (N_6685,N_6525,N_6460);
or U6686 (N_6686,N_6424,N_6349);
and U6687 (N_6687,N_6305,N_6540);
nand U6688 (N_6688,N_6412,N_6516);
nand U6689 (N_6689,N_6381,N_6507);
nor U6690 (N_6690,N_6366,N_6413);
or U6691 (N_6691,N_6580,N_6449);
or U6692 (N_6692,N_6360,N_6485);
xor U6693 (N_6693,N_6509,N_6408);
nor U6694 (N_6694,N_6433,N_6527);
or U6695 (N_6695,N_6397,N_6466);
nor U6696 (N_6696,N_6499,N_6312);
or U6697 (N_6697,N_6417,N_6561);
xor U6698 (N_6698,N_6426,N_6365);
and U6699 (N_6699,N_6389,N_6386);
and U6700 (N_6700,N_6510,N_6351);
nand U6701 (N_6701,N_6306,N_6324);
xor U6702 (N_6702,N_6344,N_6477);
xor U6703 (N_6703,N_6481,N_6325);
xor U6704 (N_6704,N_6368,N_6406);
xnor U6705 (N_6705,N_6369,N_6420);
and U6706 (N_6706,N_6370,N_6558);
and U6707 (N_6707,N_6567,N_6582);
and U6708 (N_6708,N_6391,N_6550);
xnor U6709 (N_6709,N_6390,N_6382);
nand U6710 (N_6710,N_6427,N_6503);
xnor U6711 (N_6711,N_6512,N_6570);
or U6712 (N_6712,N_6314,N_6554);
nor U6713 (N_6713,N_6547,N_6536);
and U6714 (N_6714,N_6595,N_6575);
nor U6715 (N_6715,N_6459,N_6493);
or U6716 (N_6716,N_6364,N_6564);
xor U6717 (N_6717,N_6387,N_6457);
and U6718 (N_6718,N_6468,N_6343);
nor U6719 (N_6719,N_6577,N_6376);
and U6720 (N_6720,N_6447,N_6494);
nand U6721 (N_6721,N_6566,N_6552);
nor U6722 (N_6722,N_6443,N_6514);
xnor U6723 (N_6723,N_6336,N_6589);
xnor U6724 (N_6724,N_6415,N_6377);
and U6725 (N_6725,N_6308,N_6400);
nor U6726 (N_6726,N_6418,N_6405);
nor U6727 (N_6727,N_6428,N_6498);
xor U6728 (N_6728,N_6534,N_6596);
xor U6729 (N_6729,N_6543,N_6573);
and U6730 (N_6730,N_6435,N_6475);
and U6731 (N_6731,N_6518,N_6373);
and U6732 (N_6732,N_6320,N_6551);
nand U6733 (N_6733,N_6482,N_6340);
or U6734 (N_6734,N_6464,N_6322);
nand U6735 (N_6735,N_6586,N_6533);
or U6736 (N_6736,N_6508,N_6337);
or U6737 (N_6737,N_6378,N_6542);
nor U6738 (N_6738,N_6463,N_6555);
xnor U6739 (N_6739,N_6473,N_6467);
xor U6740 (N_6740,N_6553,N_6436);
nand U6741 (N_6741,N_6511,N_6454);
or U6742 (N_6742,N_6329,N_6374);
nand U6743 (N_6743,N_6450,N_6347);
nor U6744 (N_6744,N_6451,N_6393);
or U6745 (N_6745,N_6345,N_6452);
xnor U6746 (N_6746,N_6342,N_6404);
or U6747 (N_6747,N_6355,N_6431);
nand U6748 (N_6748,N_6541,N_6592);
and U6749 (N_6749,N_6361,N_6474);
nand U6750 (N_6750,N_6599,N_6388);
nand U6751 (N_6751,N_6409,N_6399);
nor U6752 (N_6752,N_6416,N_6304);
xor U6753 (N_6753,N_6521,N_6463);
or U6754 (N_6754,N_6499,N_6322);
or U6755 (N_6755,N_6431,N_6526);
nand U6756 (N_6756,N_6460,N_6335);
xnor U6757 (N_6757,N_6486,N_6523);
nand U6758 (N_6758,N_6333,N_6389);
or U6759 (N_6759,N_6404,N_6456);
or U6760 (N_6760,N_6354,N_6428);
nand U6761 (N_6761,N_6356,N_6339);
and U6762 (N_6762,N_6473,N_6392);
xor U6763 (N_6763,N_6401,N_6340);
nand U6764 (N_6764,N_6418,N_6573);
and U6765 (N_6765,N_6401,N_6362);
and U6766 (N_6766,N_6502,N_6524);
or U6767 (N_6767,N_6456,N_6468);
nand U6768 (N_6768,N_6442,N_6481);
xnor U6769 (N_6769,N_6378,N_6363);
nor U6770 (N_6770,N_6523,N_6436);
or U6771 (N_6771,N_6405,N_6598);
or U6772 (N_6772,N_6323,N_6539);
nor U6773 (N_6773,N_6444,N_6561);
and U6774 (N_6774,N_6568,N_6446);
or U6775 (N_6775,N_6574,N_6363);
nand U6776 (N_6776,N_6465,N_6545);
nor U6777 (N_6777,N_6429,N_6452);
xor U6778 (N_6778,N_6378,N_6490);
and U6779 (N_6779,N_6456,N_6563);
and U6780 (N_6780,N_6552,N_6527);
nand U6781 (N_6781,N_6374,N_6387);
or U6782 (N_6782,N_6562,N_6442);
or U6783 (N_6783,N_6481,N_6318);
nand U6784 (N_6784,N_6494,N_6574);
and U6785 (N_6785,N_6477,N_6339);
xor U6786 (N_6786,N_6545,N_6589);
or U6787 (N_6787,N_6307,N_6441);
xnor U6788 (N_6788,N_6389,N_6330);
nand U6789 (N_6789,N_6556,N_6408);
or U6790 (N_6790,N_6322,N_6487);
nand U6791 (N_6791,N_6492,N_6433);
nor U6792 (N_6792,N_6585,N_6403);
xnor U6793 (N_6793,N_6316,N_6447);
nor U6794 (N_6794,N_6353,N_6469);
nand U6795 (N_6795,N_6477,N_6402);
nor U6796 (N_6796,N_6339,N_6503);
or U6797 (N_6797,N_6363,N_6400);
nor U6798 (N_6798,N_6403,N_6535);
xnor U6799 (N_6799,N_6378,N_6518);
xnor U6800 (N_6800,N_6523,N_6346);
nor U6801 (N_6801,N_6470,N_6384);
nand U6802 (N_6802,N_6533,N_6354);
nor U6803 (N_6803,N_6562,N_6328);
or U6804 (N_6804,N_6390,N_6355);
nand U6805 (N_6805,N_6373,N_6548);
or U6806 (N_6806,N_6524,N_6508);
or U6807 (N_6807,N_6458,N_6342);
nor U6808 (N_6808,N_6407,N_6348);
nand U6809 (N_6809,N_6550,N_6372);
or U6810 (N_6810,N_6384,N_6370);
xor U6811 (N_6811,N_6347,N_6406);
or U6812 (N_6812,N_6475,N_6343);
nor U6813 (N_6813,N_6359,N_6577);
or U6814 (N_6814,N_6319,N_6415);
nand U6815 (N_6815,N_6354,N_6559);
and U6816 (N_6816,N_6452,N_6341);
and U6817 (N_6817,N_6406,N_6393);
and U6818 (N_6818,N_6310,N_6336);
nor U6819 (N_6819,N_6387,N_6303);
nor U6820 (N_6820,N_6394,N_6368);
nand U6821 (N_6821,N_6314,N_6327);
and U6822 (N_6822,N_6451,N_6436);
or U6823 (N_6823,N_6352,N_6418);
and U6824 (N_6824,N_6505,N_6354);
nand U6825 (N_6825,N_6372,N_6411);
or U6826 (N_6826,N_6527,N_6560);
or U6827 (N_6827,N_6463,N_6330);
nor U6828 (N_6828,N_6388,N_6520);
or U6829 (N_6829,N_6418,N_6474);
or U6830 (N_6830,N_6561,N_6443);
and U6831 (N_6831,N_6357,N_6595);
xor U6832 (N_6832,N_6301,N_6455);
or U6833 (N_6833,N_6599,N_6438);
xnor U6834 (N_6834,N_6552,N_6398);
nand U6835 (N_6835,N_6332,N_6371);
and U6836 (N_6836,N_6314,N_6300);
nor U6837 (N_6837,N_6578,N_6574);
or U6838 (N_6838,N_6420,N_6511);
nor U6839 (N_6839,N_6410,N_6599);
or U6840 (N_6840,N_6530,N_6509);
xnor U6841 (N_6841,N_6388,N_6457);
nor U6842 (N_6842,N_6562,N_6327);
xor U6843 (N_6843,N_6474,N_6525);
nor U6844 (N_6844,N_6537,N_6569);
or U6845 (N_6845,N_6446,N_6487);
nor U6846 (N_6846,N_6426,N_6548);
xor U6847 (N_6847,N_6339,N_6309);
nand U6848 (N_6848,N_6534,N_6431);
or U6849 (N_6849,N_6427,N_6383);
nand U6850 (N_6850,N_6344,N_6593);
xnor U6851 (N_6851,N_6582,N_6342);
xor U6852 (N_6852,N_6564,N_6475);
nand U6853 (N_6853,N_6351,N_6328);
and U6854 (N_6854,N_6572,N_6305);
nand U6855 (N_6855,N_6475,N_6400);
or U6856 (N_6856,N_6500,N_6399);
xnor U6857 (N_6857,N_6554,N_6479);
and U6858 (N_6858,N_6503,N_6488);
xor U6859 (N_6859,N_6547,N_6379);
or U6860 (N_6860,N_6530,N_6597);
xnor U6861 (N_6861,N_6587,N_6513);
or U6862 (N_6862,N_6475,N_6337);
nor U6863 (N_6863,N_6580,N_6394);
and U6864 (N_6864,N_6346,N_6588);
nand U6865 (N_6865,N_6355,N_6410);
nand U6866 (N_6866,N_6442,N_6359);
nand U6867 (N_6867,N_6314,N_6467);
and U6868 (N_6868,N_6421,N_6322);
nand U6869 (N_6869,N_6506,N_6553);
or U6870 (N_6870,N_6570,N_6390);
and U6871 (N_6871,N_6591,N_6373);
nor U6872 (N_6872,N_6353,N_6407);
or U6873 (N_6873,N_6462,N_6436);
nand U6874 (N_6874,N_6352,N_6452);
nand U6875 (N_6875,N_6517,N_6590);
nand U6876 (N_6876,N_6438,N_6425);
xnor U6877 (N_6877,N_6504,N_6412);
xor U6878 (N_6878,N_6490,N_6337);
xnor U6879 (N_6879,N_6385,N_6484);
xnor U6880 (N_6880,N_6556,N_6430);
nor U6881 (N_6881,N_6469,N_6316);
nor U6882 (N_6882,N_6469,N_6300);
nor U6883 (N_6883,N_6523,N_6511);
or U6884 (N_6884,N_6462,N_6318);
and U6885 (N_6885,N_6366,N_6494);
nand U6886 (N_6886,N_6599,N_6404);
nand U6887 (N_6887,N_6504,N_6472);
and U6888 (N_6888,N_6479,N_6548);
or U6889 (N_6889,N_6436,N_6403);
nor U6890 (N_6890,N_6382,N_6560);
or U6891 (N_6891,N_6499,N_6470);
xor U6892 (N_6892,N_6327,N_6302);
or U6893 (N_6893,N_6485,N_6568);
nor U6894 (N_6894,N_6388,N_6380);
xnor U6895 (N_6895,N_6454,N_6423);
nor U6896 (N_6896,N_6578,N_6407);
or U6897 (N_6897,N_6545,N_6514);
and U6898 (N_6898,N_6596,N_6334);
and U6899 (N_6899,N_6428,N_6311);
xnor U6900 (N_6900,N_6648,N_6609);
nor U6901 (N_6901,N_6890,N_6813);
nand U6902 (N_6902,N_6762,N_6725);
xor U6903 (N_6903,N_6872,N_6803);
or U6904 (N_6904,N_6863,N_6738);
xnor U6905 (N_6905,N_6669,N_6606);
or U6906 (N_6906,N_6732,N_6651);
xnor U6907 (N_6907,N_6770,N_6670);
or U6908 (N_6908,N_6826,N_6800);
nor U6909 (N_6909,N_6704,N_6897);
or U6910 (N_6910,N_6717,N_6878);
nand U6911 (N_6911,N_6786,N_6864);
nand U6912 (N_6912,N_6862,N_6846);
nor U6913 (N_6913,N_6691,N_6823);
nand U6914 (N_6914,N_6697,N_6811);
xor U6915 (N_6915,N_6640,N_6616);
nor U6916 (N_6916,N_6888,N_6707);
or U6917 (N_6917,N_6642,N_6849);
nand U6918 (N_6918,N_6714,N_6745);
nand U6919 (N_6919,N_6735,N_6664);
or U6920 (N_6920,N_6752,N_6782);
or U6921 (N_6921,N_6612,N_6604);
and U6922 (N_6922,N_6814,N_6620);
or U6923 (N_6923,N_6785,N_6624);
xor U6924 (N_6924,N_6812,N_6706);
and U6925 (N_6925,N_6600,N_6644);
and U6926 (N_6926,N_6774,N_6672);
nor U6927 (N_6927,N_6743,N_6737);
or U6928 (N_6928,N_6626,N_6840);
nand U6929 (N_6929,N_6764,N_6793);
xnor U6930 (N_6930,N_6754,N_6692);
xor U6931 (N_6931,N_6815,N_6772);
nand U6932 (N_6932,N_6755,N_6744);
nor U6933 (N_6933,N_6628,N_6850);
nor U6934 (N_6934,N_6729,N_6768);
nor U6935 (N_6935,N_6712,N_6666);
nand U6936 (N_6936,N_6833,N_6750);
or U6937 (N_6937,N_6667,N_6660);
nor U6938 (N_6938,N_6858,N_6638);
nand U6939 (N_6939,N_6733,N_6654);
xor U6940 (N_6940,N_6899,N_6771);
and U6941 (N_6941,N_6724,N_6865);
or U6942 (N_6942,N_6778,N_6731);
xor U6943 (N_6943,N_6810,N_6822);
or U6944 (N_6944,N_6649,N_6751);
xnor U6945 (N_6945,N_6859,N_6845);
and U6946 (N_6946,N_6690,N_6631);
and U6947 (N_6947,N_6795,N_6866);
and U6948 (N_6948,N_6877,N_6775);
and U6949 (N_6949,N_6898,N_6881);
nor U6950 (N_6950,N_6851,N_6821);
or U6951 (N_6951,N_6879,N_6788);
and U6952 (N_6952,N_6799,N_6883);
and U6953 (N_6953,N_6676,N_6875);
and U6954 (N_6954,N_6806,N_6791);
nor U6955 (N_6955,N_6838,N_6792);
xor U6956 (N_6956,N_6699,N_6721);
and U6957 (N_6957,N_6619,N_6686);
xor U6958 (N_6958,N_6645,N_6734);
and U6959 (N_6959,N_6759,N_6677);
nor U6960 (N_6960,N_6887,N_6643);
nand U6961 (N_6961,N_6684,N_6873);
xnor U6962 (N_6962,N_6694,N_6876);
nor U6963 (N_6963,N_6861,N_6632);
nor U6964 (N_6964,N_6831,N_6773);
nor U6965 (N_6965,N_6728,N_6659);
nand U6966 (N_6966,N_6709,N_6705);
or U6967 (N_6967,N_6746,N_6650);
xnor U6968 (N_6968,N_6767,N_6688);
nand U6969 (N_6969,N_6882,N_6629);
nand U6970 (N_6970,N_6622,N_6824);
xor U6971 (N_6971,N_6856,N_6653);
xnor U6972 (N_6972,N_6711,N_6718);
and U6973 (N_6973,N_6608,N_6753);
and U6974 (N_6974,N_6647,N_6675);
xnor U6975 (N_6975,N_6781,N_6830);
nor U6976 (N_6976,N_6844,N_6836);
xnor U6977 (N_6977,N_6683,N_6817);
nand U6978 (N_6978,N_6662,N_6860);
xnor U6979 (N_6979,N_6896,N_6842);
xnor U6980 (N_6980,N_6784,N_6723);
nand U6981 (N_6981,N_6868,N_6617);
xnor U6982 (N_6982,N_6852,N_6740);
nand U6983 (N_6983,N_6702,N_6713);
nand U6984 (N_6984,N_6671,N_6720);
or U6985 (N_6985,N_6889,N_6886);
nand U6986 (N_6986,N_6646,N_6804);
nand U6987 (N_6987,N_6805,N_6763);
and U6988 (N_6988,N_6656,N_6652);
and U6989 (N_6989,N_6736,N_6779);
nor U6990 (N_6990,N_6777,N_6818);
and U6991 (N_6991,N_6867,N_6603);
xnor U6992 (N_6992,N_6607,N_6801);
and U6993 (N_6993,N_6722,N_6621);
nand U6994 (N_6994,N_6829,N_6894);
or U6995 (N_6995,N_6657,N_6885);
xor U6996 (N_6996,N_6661,N_6708);
xor U6997 (N_6997,N_6655,N_6847);
or U6998 (N_6998,N_6613,N_6756);
and U6999 (N_6999,N_6841,N_6601);
and U7000 (N_7000,N_6627,N_6630);
or U7001 (N_7001,N_6780,N_6695);
and U7002 (N_7002,N_6816,N_6637);
and U7003 (N_7003,N_6741,N_6837);
or U7004 (N_7004,N_6835,N_6614);
or U7005 (N_7005,N_6820,N_6696);
and U7006 (N_7006,N_6854,N_6892);
and U7007 (N_7007,N_6698,N_6730);
nand U7008 (N_7008,N_6689,N_6633);
xor U7009 (N_7009,N_6749,N_6727);
or U7010 (N_7010,N_6674,N_6665);
xnor U7011 (N_7011,N_6819,N_6639);
or U7012 (N_7012,N_6700,N_6681);
nand U7013 (N_7013,N_6615,N_6832);
and U7014 (N_7014,N_6658,N_6769);
nand U7015 (N_7015,N_6807,N_6787);
or U7016 (N_7016,N_6869,N_6625);
nand U7017 (N_7017,N_6668,N_6760);
and U7018 (N_7018,N_6701,N_6739);
and U7019 (N_7019,N_6678,N_6874);
or U7020 (N_7020,N_6719,N_6687);
xor U7021 (N_7021,N_6680,N_6623);
nand U7022 (N_7022,N_6827,N_6747);
and U7023 (N_7023,N_6843,N_6891);
and U7024 (N_7024,N_6798,N_6857);
xnor U7025 (N_7025,N_6783,N_6839);
nor U7026 (N_7026,N_6825,N_6776);
and U7027 (N_7027,N_6828,N_6663);
and U7028 (N_7028,N_6802,N_6641);
nor U7029 (N_7029,N_6757,N_6685);
or U7030 (N_7030,N_6602,N_6790);
or U7031 (N_7031,N_6761,N_6618);
and U7032 (N_7032,N_6870,N_6742);
xnor U7033 (N_7033,N_6703,N_6635);
and U7034 (N_7034,N_6855,N_6853);
xor U7035 (N_7035,N_6834,N_6748);
xor U7036 (N_7036,N_6871,N_6679);
and U7037 (N_7037,N_6765,N_6895);
and U7038 (N_7038,N_6766,N_6693);
or U7039 (N_7039,N_6893,N_6796);
or U7040 (N_7040,N_6797,N_6884);
or U7041 (N_7041,N_6673,N_6880);
or U7042 (N_7042,N_6605,N_6758);
nor U7043 (N_7043,N_6848,N_6789);
nor U7044 (N_7044,N_6610,N_6794);
or U7045 (N_7045,N_6710,N_6808);
nand U7046 (N_7046,N_6726,N_6682);
nor U7047 (N_7047,N_6716,N_6634);
and U7048 (N_7048,N_6715,N_6611);
xor U7049 (N_7049,N_6809,N_6636);
or U7050 (N_7050,N_6646,N_6663);
or U7051 (N_7051,N_6626,N_6650);
and U7052 (N_7052,N_6768,N_6704);
and U7053 (N_7053,N_6671,N_6813);
and U7054 (N_7054,N_6842,N_6834);
nor U7055 (N_7055,N_6886,N_6627);
nor U7056 (N_7056,N_6751,N_6750);
and U7057 (N_7057,N_6773,N_6608);
or U7058 (N_7058,N_6832,N_6635);
xnor U7059 (N_7059,N_6882,N_6738);
xor U7060 (N_7060,N_6720,N_6630);
and U7061 (N_7061,N_6715,N_6722);
nand U7062 (N_7062,N_6760,N_6608);
nor U7063 (N_7063,N_6886,N_6780);
nor U7064 (N_7064,N_6789,N_6736);
xor U7065 (N_7065,N_6886,N_6661);
xnor U7066 (N_7066,N_6737,N_6738);
nand U7067 (N_7067,N_6685,N_6852);
and U7068 (N_7068,N_6604,N_6729);
nor U7069 (N_7069,N_6751,N_6618);
and U7070 (N_7070,N_6865,N_6893);
or U7071 (N_7071,N_6849,N_6877);
nor U7072 (N_7072,N_6852,N_6644);
or U7073 (N_7073,N_6603,N_6675);
nand U7074 (N_7074,N_6669,N_6758);
or U7075 (N_7075,N_6769,N_6713);
or U7076 (N_7076,N_6867,N_6793);
nor U7077 (N_7077,N_6733,N_6780);
nand U7078 (N_7078,N_6737,N_6615);
and U7079 (N_7079,N_6624,N_6682);
nor U7080 (N_7080,N_6715,N_6791);
or U7081 (N_7081,N_6842,N_6693);
or U7082 (N_7082,N_6804,N_6872);
nor U7083 (N_7083,N_6842,N_6607);
xor U7084 (N_7084,N_6795,N_6750);
and U7085 (N_7085,N_6874,N_6609);
nand U7086 (N_7086,N_6842,N_6637);
nor U7087 (N_7087,N_6893,N_6672);
or U7088 (N_7088,N_6678,N_6686);
xnor U7089 (N_7089,N_6893,N_6774);
and U7090 (N_7090,N_6792,N_6870);
xor U7091 (N_7091,N_6648,N_6823);
nand U7092 (N_7092,N_6763,N_6627);
nor U7093 (N_7093,N_6843,N_6768);
nand U7094 (N_7094,N_6803,N_6715);
and U7095 (N_7095,N_6859,N_6771);
xnor U7096 (N_7096,N_6880,N_6727);
xnor U7097 (N_7097,N_6789,N_6893);
or U7098 (N_7098,N_6863,N_6698);
nand U7099 (N_7099,N_6696,N_6803);
and U7100 (N_7100,N_6825,N_6791);
nor U7101 (N_7101,N_6898,N_6698);
or U7102 (N_7102,N_6729,N_6883);
nand U7103 (N_7103,N_6698,N_6834);
or U7104 (N_7104,N_6843,N_6836);
and U7105 (N_7105,N_6645,N_6757);
xnor U7106 (N_7106,N_6774,N_6694);
and U7107 (N_7107,N_6615,N_6841);
and U7108 (N_7108,N_6635,N_6718);
nand U7109 (N_7109,N_6858,N_6665);
or U7110 (N_7110,N_6897,N_6867);
and U7111 (N_7111,N_6886,N_6653);
and U7112 (N_7112,N_6822,N_6873);
and U7113 (N_7113,N_6861,N_6643);
or U7114 (N_7114,N_6669,N_6707);
nor U7115 (N_7115,N_6840,N_6718);
and U7116 (N_7116,N_6626,N_6852);
nand U7117 (N_7117,N_6674,N_6715);
nor U7118 (N_7118,N_6815,N_6825);
xnor U7119 (N_7119,N_6676,N_6695);
and U7120 (N_7120,N_6647,N_6634);
nor U7121 (N_7121,N_6841,N_6826);
xnor U7122 (N_7122,N_6857,N_6733);
nor U7123 (N_7123,N_6695,N_6603);
or U7124 (N_7124,N_6831,N_6843);
nor U7125 (N_7125,N_6736,N_6674);
or U7126 (N_7126,N_6742,N_6867);
nand U7127 (N_7127,N_6847,N_6750);
xnor U7128 (N_7128,N_6715,N_6760);
nand U7129 (N_7129,N_6869,N_6620);
nand U7130 (N_7130,N_6850,N_6722);
or U7131 (N_7131,N_6891,N_6862);
or U7132 (N_7132,N_6600,N_6655);
and U7133 (N_7133,N_6726,N_6812);
nand U7134 (N_7134,N_6771,N_6887);
nor U7135 (N_7135,N_6781,N_6648);
or U7136 (N_7136,N_6884,N_6791);
xnor U7137 (N_7137,N_6790,N_6647);
nor U7138 (N_7138,N_6692,N_6816);
or U7139 (N_7139,N_6754,N_6611);
nand U7140 (N_7140,N_6631,N_6620);
nand U7141 (N_7141,N_6752,N_6721);
or U7142 (N_7142,N_6686,N_6832);
xnor U7143 (N_7143,N_6628,N_6729);
nand U7144 (N_7144,N_6811,N_6656);
and U7145 (N_7145,N_6712,N_6810);
or U7146 (N_7146,N_6628,N_6859);
and U7147 (N_7147,N_6811,N_6669);
xnor U7148 (N_7148,N_6789,N_6747);
nor U7149 (N_7149,N_6688,N_6701);
and U7150 (N_7150,N_6789,N_6770);
nor U7151 (N_7151,N_6764,N_6713);
nand U7152 (N_7152,N_6727,N_6719);
and U7153 (N_7153,N_6707,N_6785);
nor U7154 (N_7154,N_6875,N_6735);
and U7155 (N_7155,N_6828,N_6820);
nand U7156 (N_7156,N_6837,N_6894);
nand U7157 (N_7157,N_6826,N_6687);
or U7158 (N_7158,N_6799,N_6694);
or U7159 (N_7159,N_6797,N_6615);
xnor U7160 (N_7160,N_6623,N_6683);
and U7161 (N_7161,N_6841,N_6605);
nor U7162 (N_7162,N_6677,N_6698);
nand U7163 (N_7163,N_6750,N_6660);
and U7164 (N_7164,N_6843,N_6842);
xnor U7165 (N_7165,N_6707,N_6741);
nor U7166 (N_7166,N_6858,N_6628);
and U7167 (N_7167,N_6648,N_6787);
xnor U7168 (N_7168,N_6689,N_6608);
and U7169 (N_7169,N_6713,N_6897);
nand U7170 (N_7170,N_6810,N_6619);
and U7171 (N_7171,N_6734,N_6794);
nand U7172 (N_7172,N_6793,N_6844);
xor U7173 (N_7173,N_6869,N_6775);
nand U7174 (N_7174,N_6783,N_6678);
or U7175 (N_7175,N_6752,N_6636);
xnor U7176 (N_7176,N_6633,N_6681);
nor U7177 (N_7177,N_6806,N_6605);
or U7178 (N_7178,N_6744,N_6827);
and U7179 (N_7179,N_6639,N_6695);
xor U7180 (N_7180,N_6818,N_6773);
nor U7181 (N_7181,N_6840,N_6831);
nor U7182 (N_7182,N_6643,N_6805);
xnor U7183 (N_7183,N_6669,N_6733);
or U7184 (N_7184,N_6622,N_6724);
and U7185 (N_7185,N_6737,N_6704);
nor U7186 (N_7186,N_6610,N_6654);
or U7187 (N_7187,N_6670,N_6708);
nand U7188 (N_7188,N_6640,N_6639);
and U7189 (N_7189,N_6814,N_6602);
nand U7190 (N_7190,N_6789,N_6850);
xor U7191 (N_7191,N_6743,N_6654);
nor U7192 (N_7192,N_6741,N_6854);
or U7193 (N_7193,N_6645,N_6792);
nand U7194 (N_7194,N_6768,N_6822);
nand U7195 (N_7195,N_6765,N_6888);
or U7196 (N_7196,N_6793,N_6868);
nor U7197 (N_7197,N_6866,N_6851);
or U7198 (N_7198,N_6847,N_6855);
xnor U7199 (N_7199,N_6739,N_6862);
nor U7200 (N_7200,N_6964,N_7139);
nand U7201 (N_7201,N_7102,N_6981);
nand U7202 (N_7202,N_6992,N_7010);
or U7203 (N_7203,N_7192,N_7170);
nand U7204 (N_7204,N_6998,N_7022);
nor U7205 (N_7205,N_6949,N_7001);
or U7206 (N_7206,N_6963,N_7061);
nand U7207 (N_7207,N_6936,N_6987);
xnor U7208 (N_7208,N_7028,N_7136);
xnor U7209 (N_7209,N_6991,N_7056);
or U7210 (N_7210,N_7162,N_7002);
and U7211 (N_7211,N_7097,N_6950);
nand U7212 (N_7212,N_6931,N_7089);
and U7213 (N_7213,N_7073,N_7103);
and U7214 (N_7214,N_6996,N_6916);
xor U7215 (N_7215,N_7081,N_7063);
xnor U7216 (N_7216,N_6958,N_6937);
nand U7217 (N_7217,N_6915,N_7155);
and U7218 (N_7218,N_7105,N_6925);
nor U7219 (N_7219,N_6944,N_7163);
nand U7220 (N_7220,N_7067,N_6960);
nor U7221 (N_7221,N_7033,N_7008);
nor U7222 (N_7222,N_7084,N_7101);
and U7223 (N_7223,N_7151,N_7126);
xnor U7224 (N_7224,N_6910,N_7172);
xnor U7225 (N_7225,N_6989,N_7032);
nand U7226 (N_7226,N_7177,N_6945);
xnor U7227 (N_7227,N_7121,N_7047);
and U7228 (N_7228,N_6968,N_7000);
or U7229 (N_7229,N_6900,N_6922);
xor U7230 (N_7230,N_7123,N_6933);
nor U7231 (N_7231,N_6965,N_6970);
nand U7232 (N_7232,N_7188,N_7074);
and U7233 (N_7233,N_7183,N_6903);
or U7234 (N_7234,N_6920,N_7058);
and U7235 (N_7235,N_7153,N_7026);
or U7236 (N_7236,N_6923,N_6914);
and U7237 (N_7237,N_7100,N_7112);
xor U7238 (N_7238,N_7087,N_7193);
nand U7239 (N_7239,N_6943,N_6974);
or U7240 (N_7240,N_7020,N_7159);
nand U7241 (N_7241,N_7118,N_7158);
or U7242 (N_7242,N_6940,N_7039);
or U7243 (N_7243,N_7117,N_7161);
and U7244 (N_7244,N_7044,N_6932);
or U7245 (N_7245,N_6985,N_6928);
and U7246 (N_7246,N_7122,N_6951);
or U7247 (N_7247,N_6942,N_7075);
or U7248 (N_7248,N_6962,N_7050);
nor U7249 (N_7249,N_7149,N_7066);
and U7250 (N_7250,N_6953,N_7070);
xor U7251 (N_7251,N_7168,N_7128);
nor U7252 (N_7252,N_7154,N_7140);
and U7253 (N_7253,N_7059,N_7182);
xor U7254 (N_7254,N_7072,N_7080);
nor U7255 (N_7255,N_7077,N_7052);
and U7256 (N_7256,N_7143,N_7009);
nand U7257 (N_7257,N_7131,N_6926);
or U7258 (N_7258,N_6902,N_6921);
nor U7259 (N_7259,N_6975,N_6979);
nor U7260 (N_7260,N_6911,N_7124);
xnor U7261 (N_7261,N_6918,N_7133);
xnor U7262 (N_7262,N_6907,N_7135);
and U7263 (N_7263,N_7173,N_6959);
nor U7264 (N_7264,N_7194,N_7069);
nand U7265 (N_7265,N_6939,N_7023);
nor U7266 (N_7266,N_7167,N_7197);
nor U7267 (N_7267,N_7152,N_6990);
or U7268 (N_7268,N_6924,N_7021);
xnor U7269 (N_7269,N_7109,N_7132);
or U7270 (N_7270,N_7005,N_6999);
nor U7271 (N_7271,N_7160,N_7006);
or U7272 (N_7272,N_7012,N_7079);
and U7273 (N_7273,N_7156,N_6956);
nor U7274 (N_7274,N_7038,N_7180);
xor U7275 (N_7275,N_7146,N_6934);
and U7276 (N_7276,N_7025,N_7013);
or U7277 (N_7277,N_7198,N_7065);
or U7278 (N_7278,N_7147,N_7106);
and U7279 (N_7279,N_7062,N_7191);
nand U7280 (N_7280,N_7018,N_6973);
xor U7281 (N_7281,N_7041,N_7196);
nor U7282 (N_7282,N_6955,N_7035);
xnor U7283 (N_7283,N_6901,N_7114);
and U7284 (N_7284,N_6982,N_7003);
and U7285 (N_7285,N_7043,N_7092);
xor U7286 (N_7286,N_7007,N_7071);
and U7287 (N_7287,N_6952,N_7099);
or U7288 (N_7288,N_7088,N_7108);
and U7289 (N_7289,N_6941,N_7157);
and U7290 (N_7290,N_6946,N_7019);
nand U7291 (N_7291,N_7185,N_7119);
xnor U7292 (N_7292,N_7016,N_6935);
and U7293 (N_7293,N_7051,N_6909);
nand U7294 (N_7294,N_6966,N_7094);
nor U7295 (N_7295,N_7085,N_7179);
or U7296 (N_7296,N_7060,N_6995);
nand U7297 (N_7297,N_7031,N_6905);
or U7298 (N_7298,N_7045,N_7148);
or U7299 (N_7299,N_7049,N_7053);
or U7300 (N_7300,N_7091,N_7137);
xnor U7301 (N_7301,N_7034,N_7030);
nand U7302 (N_7302,N_6938,N_7004);
xnor U7303 (N_7303,N_7096,N_7187);
xnor U7304 (N_7304,N_6961,N_7178);
and U7305 (N_7305,N_7166,N_7144);
nor U7306 (N_7306,N_7113,N_7027);
or U7307 (N_7307,N_6977,N_6927);
nand U7308 (N_7308,N_7090,N_6983);
nor U7309 (N_7309,N_6972,N_7104);
nor U7310 (N_7310,N_7098,N_7055);
and U7311 (N_7311,N_6986,N_6980);
nor U7312 (N_7312,N_7078,N_6997);
nand U7313 (N_7313,N_6976,N_7134);
or U7314 (N_7314,N_6913,N_7181);
or U7315 (N_7315,N_6917,N_7037);
nor U7316 (N_7316,N_7145,N_6904);
nand U7317 (N_7317,N_6930,N_7093);
nor U7318 (N_7318,N_7042,N_6948);
xnor U7319 (N_7319,N_7116,N_7169);
and U7320 (N_7320,N_7111,N_7199);
xor U7321 (N_7321,N_7130,N_6978);
or U7322 (N_7322,N_7171,N_7082);
xor U7323 (N_7323,N_7129,N_7048);
nand U7324 (N_7324,N_7138,N_7125);
xor U7325 (N_7325,N_7054,N_7017);
xor U7326 (N_7326,N_6912,N_7029);
nand U7327 (N_7327,N_7186,N_7046);
and U7328 (N_7328,N_7110,N_7036);
and U7329 (N_7329,N_7127,N_7184);
and U7330 (N_7330,N_6947,N_7064);
nand U7331 (N_7331,N_6954,N_7115);
nor U7332 (N_7332,N_7120,N_7076);
nor U7333 (N_7333,N_6994,N_6969);
and U7334 (N_7334,N_7107,N_6957);
or U7335 (N_7335,N_7150,N_6929);
nand U7336 (N_7336,N_7015,N_7095);
nor U7337 (N_7337,N_6906,N_6908);
nand U7338 (N_7338,N_7174,N_6967);
and U7339 (N_7339,N_6988,N_7040);
nor U7340 (N_7340,N_7057,N_7164);
nor U7341 (N_7341,N_7175,N_7141);
nor U7342 (N_7342,N_7176,N_6971);
or U7343 (N_7343,N_7086,N_7195);
xnor U7344 (N_7344,N_7083,N_7024);
and U7345 (N_7345,N_7014,N_7068);
nor U7346 (N_7346,N_7011,N_6993);
and U7347 (N_7347,N_7190,N_7142);
xor U7348 (N_7348,N_7165,N_6984);
or U7349 (N_7349,N_7189,N_6919);
and U7350 (N_7350,N_7080,N_7189);
and U7351 (N_7351,N_7014,N_7055);
nand U7352 (N_7352,N_7015,N_7102);
or U7353 (N_7353,N_7064,N_7124);
or U7354 (N_7354,N_6962,N_7106);
nor U7355 (N_7355,N_7125,N_7012);
xor U7356 (N_7356,N_6972,N_7050);
nor U7357 (N_7357,N_7029,N_6940);
nor U7358 (N_7358,N_6959,N_7060);
xnor U7359 (N_7359,N_7065,N_6958);
nor U7360 (N_7360,N_7079,N_7194);
or U7361 (N_7361,N_6904,N_7012);
or U7362 (N_7362,N_6971,N_7100);
nor U7363 (N_7363,N_6939,N_6985);
nand U7364 (N_7364,N_6930,N_6911);
xnor U7365 (N_7365,N_6967,N_7121);
nor U7366 (N_7366,N_7001,N_7125);
nand U7367 (N_7367,N_6918,N_7017);
or U7368 (N_7368,N_7144,N_6947);
and U7369 (N_7369,N_6952,N_6912);
xnor U7370 (N_7370,N_6930,N_6970);
nor U7371 (N_7371,N_7004,N_6985);
or U7372 (N_7372,N_7135,N_7159);
xor U7373 (N_7373,N_6946,N_6957);
nor U7374 (N_7374,N_7045,N_7195);
and U7375 (N_7375,N_7149,N_7025);
nand U7376 (N_7376,N_7184,N_7124);
and U7377 (N_7377,N_7194,N_7078);
or U7378 (N_7378,N_7049,N_6962);
nor U7379 (N_7379,N_7045,N_6900);
nor U7380 (N_7380,N_6991,N_7105);
or U7381 (N_7381,N_6981,N_6955);
and U7382 (N_7382,N_6905,N_7178);
nor U7383 (N_7383,N_7077,N_7135);
nor U7384 (N_7384,N_6979,N_6935);
and U7385 (N_7385,N_7064,N_7006);
nor U7386 (N_7386,N_6949,N_6947);
and U7387 (N_7387,N_6946,N_6928);
nand U7388 (N_7388,N_6914,N_7016);
xor U7389 (N_7389,N_6947,N_6942);
nand U7390 (N_7390,N_6943,N_6927);
or U7391 (N_7391,N_6935,N_7103);
and U7392 (N_7392,N_7008,N_6976);
or U7393 (N_7393,N_7179,N_6951);
nand U7394 (N_7394,N_7186,N_6904);
xnor U7395 (N_7395,N_6936,N_7118);
or U7396 (N_7396,N_7117,N_7192);
or U7397 (N_7397,N_7080,N_7155);
and U7398 (N_7398,N_7081,N_7085);
xnor U7399 (N_7399,N_6906,N_7014);
nand U7400 (N_7400,N_7094,N_6940);
nor U7401 (N_7401,N_6939,N_7006);
and U7402 (N_7402,N_7013,N_6958);
xor U7403 (N_7403,N_6923,N_7046);
or U7404 (N_7404,N_7105,N_6997);
xor U7405 (N_7405,N_7142,N_7162);
nand U7406 (N_7406,N_7122,N_6948);
xnor U7407 (N_7407,N_7106,N_6997);
nor U7408 (N_7408,N_6922,N_7174);
nor U7409 (N_7409,N_7176,N_7133);
and U7410 (N_7410,N_6938,N_7197);
xnor U7411 (N_7411,N_6935,N_6909);
or U7412 (N_7412,N_6995,N_6982);
and U7413 (N_7413,N_7149,N_7101);
nand U7414 (N_7414,N_6910,N_7030);
and U7415 (N_7415,N_7105,N_7153);
and U7416 (N_7416,N_6915,N_6914);
and U7417 (N_7417,N_6919,N_6984);
nor U7418 (N_7418,N_7064,N_7152);
and U7419 (N_7419,N_6987,N_7162);
nand U7420 (N_7420,N_6998,N_6988);
nand U7421 (N_7421,N_7162,N_7070);
or U7422 (N_7422,N_6916,N_7143);
or U7423 (N_7423,N_7163,N_7177);
or U7424 (N_7424,N_6905,N_7081);
or U7425 (N_7425,N_6994,N_7162);
xnor U7426 (N_7426,N_6996,N_7167);
nor U7427 (N_7427,N_6913,N_7088);
xor U7428 (N_7428,N_7013,N_7089);
nand U7429 (N_7429,N_6994,N_6944);
xor U7430 (N_7430,N_6907,N_7079);
nand U7431 (N_7431,N_6963,N_7185);
nor U7432 (N_7432,N_7062,N_7159);
or U7433 (N_7433,N_7126,N_6924);
nor U7434 (N_7434,N_7170,N_7155);
nor U7435 (N_7435,N_6973,N_6966);
nand U7436 (N_7436,N_6931,N_7111);
xor U7437 (N_7437,N_7140,N_6912);
nand U7438 (N_7438,N_6926,N_7027);
or U7439 (N_7439,N_7017,N_7050);
and U7440 (N_7440,N_7069,N_7132);
and U7441 (N_7441,N_6952,N_7171);
and U7442 (N_7442,N_7115,N_7170);
nand U7443 (N_7443,N_6945,N_7095);
nand U7444 (N_7444,N_6990,N_7009);
nor U7445 (N_7445,N_6995,N_7039);
xor U7446 (N_7446,N_7029,N_6980);
or U7447 (N_7447,N_7080,N_7150);
xor U7448 (N_7448,N_7022,N_7189);
or U7449 (N_7449,N_7180,N_7004);
nor U7450 (N_7450,N_7023,N_6905);
and U7451 (N_7451,N_7129,N_6955);
and U7452 (N_7452,N_6930,N_7189);
xnor U7453 (N_7453,N_7133,N_7006);
nor U7454 (N_7454,N_7145,N_7015);
or U7455 (N_7455,N_7123,N_7164);
nand U7456 (N_7456,N_6935,N_6904);
xor U7457 (N_7457,N_7121,N_7038);
nor U7458 (N_7458,N_7128,N_7133);
and U7459 (N_7459,N_6927,N_7038);
and U7460 (N_7460,N_6919,N_7009);
nand U7461 (N_7461,N_6940,N_6935);
nand U7462 (N_7462,N_7072,N_7107);
xor U7463 (N_7463,N_7198,N_7061);
xnor U7464 (N_7464,N_7063,N_7033);
nand U7465 (N_7465,N_7171,N_7106);
nand U7466 (N_7466,N_7174,N_7034);
nand U7467 (N_7467,N_7055,N_7126);
or U7468 (N_7468,N_6923,N_6909);
and U7469 (N_7469,N_6979,N_7127);
or U7470 (N_7470,N_7162,N_7059);
xor U7471 (N_7471,N_7175,N_6949);
nand U7472 (N_7472,N_6936,N_7091);
or U7473 (N_7473,N_7063,N_7135);
and U7474 (N_7474,N_7034,N_6933);
and U7475 (N_7475,N_6997,N_6954);
nand U7476 (N_7476,N_6955,N_7096);
or U7477 (N_7477,N_7087,N_7146);
xor U7478 (N_7478,N_7198,N_6973);
nand U7479 (N_7479,N_6939,N_6971);
xnor U7480 (N_7480,N_7053,N_7010);
xnor U7481 (N_7481,N_7077,N_7099);
nor U7482 (N_7482,N_6979,N_7050);
and U7483 (N_7483,N_7076,N_6947);
xor U7484 (N_7484,N_6929,N_6942);
and U7485 (N_7485,N_6904,N_7016);
and U7486 (N_7486,N_7123,N_6971);
and U7487 (N_7487,N_6966,N_7021);
nand U7488 (N_7488,N_6973,N_7005);
nor U7489 (N_7489,N_7132,N_6960);
nor U7490 (N_7490,N_6944,N_7148);
or U7491 (N_7491,N_7022,N_6926);
nor U7492 (N_7492,N_7195,N_7122);
and U7493 (N_7493,N_7007,N_7177);
or U7494 (N_7494,N_7100,N_6920);
nor U7495 (N_7495,N_7136,N_7146);
nor U7496 (N_7496,N_7100,N_6970);
nor U7497 (N_7497,N_7131,N_7166);
and U7498 (N_7498,N_7142,N_7046);
and U7499 (N_7499,N_6970,N_7043);
nand U7500 (N_7500,N_7474,N_7405);
or U7501 (N_7501,N_7400,N_7396);
or U7502 (N_7502,N_7330,N_7308);
nor U7503 (N_7503,N_7399,N_7200);
nand U7504 (N_7504,N_7226,N_7209);
nand U7505 (N_7505,N_7448,N_7472);
nand U7506 (N_7506,N_7411,N_7394);
xnor U7507 (N_7507,N_7408,N_7404);
nand U7508 (N_7508,N_7409,N_7468);
and U7509 (N_7509,N_7457,N_7208);
and U7510 (N_7510,N_7287,N_7325);
nor U7511 (N_7511,N_7428,N_7222);
nand U7512 (N_7512,N_7388,N_7353);
and U7513 (N_7513,N_7431,N_7333);
or U7514 (N_7514,N_7444,N_7237);
or U7515 (N_7515,N_7329,N_7268);
and U7516 (N_7516,N_7312,N_7340);
nor U7517 (N_7517,N_7410,N_7452);
nor U7518 (N_7518,N_7345,N_7294);
xor U7519 (N_7519,N_7305,N_7403);
nor U7520 (N_7520,N_7355,N_7424);
or U7521 (N_7521,N_7341,N_7414);
nand U7522 (N_7522,N_7401,N_7290);
xnor U7523 (N_7523,N_7358,N_7246);
or U7524 (N_7524,N_7331,N_7378);
nand U7525 (N_7525,N_7455,N_7495);
xnor U7526 (N_7526,N_7280,N_7429);
xor U7527 (N_7527,N_7234,N_7407);
or U7528 (N_7528,N_7447,N_7377);
nand U7529 (N_7529,N_7336,N_7462);
and U7530 (N_7530,N_7286,N_7393);
nand U7531 (N_7531,N_7368,N_7205);
nand U7532 (N_7532,N_7225,N_7202);
or U7533 (N_7533,N_7430,N_7276);
or U7534 (N_7534,N_7374,N_7427);
and U7535 (N_7535,N_7385,N_7423);
and U7536 (N_7536,N_7467,N_7316);
and U7537 (N_7537,N_7386,N_7485);
nand U7538 (N_7538,N_7315,N_7483);
xnor U7539 (N_7539,N_7247,N_7440);
and U7540 (N_7540,N_7220,N_7493);
or U7541 (N_7541,N_7362,N_7283);
or U7542 (N_7542,N_7470,N_7382);
xor U7543 (N_7543,N_7299,N_7488);
nor U7544 (N_7544,N_7391,N_7351);
nor U7545 (N_7545,N_7379,N_7487);
and U7546 (N_7546,N_7475,N_7446);
nor U7547 (N_7547,N_7346,N_7432);
and U7548 (N_7548,N_7207,N_7275);
and U7549 (N_7549,N_7381,N_7497);
and U7550 (N_7550,N_7288,N_7301);
nor U7551 (N_7551,N_7367,N_7491);
xnor U7552 (N_7552,N_7480,N_7257);
and U7553 (N_7553,N_7298,N_7376);
nor U7554 (N_7554,N_7266,N_7380);
nor U7555 (N_7555,N_7267,N_7383);
and U7556 (N_7556,N_7332,N_7252);
xor U7557 (N_7557,N_7434,N_7450);
or U7558 (N_7558,N_7461,N_7342);
nand U7559 (N_7559,N_7242,N_7221);
and U7560 (N_7560,N_7392,N_7296);
nand U7561 (N_7561,N_7343,N_7415);
or U7562 (N_7562,N_7489,N_7344);
and U7563 (N_7563,N_7473,N_7292);
nand U7564 (N_7564,N_7433,N_7321);
nor U7565 (N_7565,N_7369,N_7256);
or U7566 (N_7566,N_7241,N_7307);
nor U7567 (N_7567,N_7420,N_7232);
or U7568 (N_7568,N_7214,N_7387);
xor U7569 (N_7569,N_7212,N_7295);
nand U7570 (N_7570,N_7317,N_7261);
nand U7571 (N_7571,N_7435,N_7318);
xor U7572 (N_7572,N_7281,N_7459);
and U7573 (N_7573,N_7293,N_7204);
nor U7574 (N_7574,N_7398,N_7402);
xor U7575 (N_7575,N_7464,N_7313);
nor U7576 (N_7576,N_7322,N_7479);
nand U7577 (N_7577,N_7233,N_7311);
nand U7578 (N_7578,N_7370,N_7359);
or U7579 (N_7579,N_7463,N_7361);
nor U7580 (N_7580,N_7297,N_7412);
xnor U7581 (N_7581,N_7496,N_7278);
nand U7582 (N_7582,N_7328,N_7249);
xor U7583 (N_7583,N_7338,N_7436);
nand U7584 (N_7584,N_7319,N_7389);
nand U7585 (N_7585,N_7218,N_7310);
and U7586 (N_7586,N_7250,N_7289);
xnor U7587 (N_7587,N_7373,N_7445);
or U7588 (N_7588,N_7438,N_7265);
nand U7589 (N_7589,N_7255,N_7366);
and U7590 (N_7590,N_7360,N_7260);
or U7591 (N_7591,N_7456,N_7395);
nand U7592 (N_7592,N_7236,N_7270);
nand U7593 (N_7593,N_7215,N_7264);
nand U7594 (N_7594,N_7245,N_7478);
and U7595 (N_7595,N_7213,N_7284);
nor U7596 (N_7596,N_7384,N_7426);
nand U7597 (N_7597,N_7300,N_7486);
and U7598 (N_7598,N_7454,N_7248);
nand U7599 (N_7599,N_7258,N_7372);
or U7600 (N_7600,N_7498,N_7211);
or U7601 (N_7601,N_7302,N_7303);
nor U7602 (N_7602,N_7254,N_7269);
or U7603 (N_7603,N_7304,N_7458);
and U7604 (N_7604,N_7335,N_7244);
nand U7605 (N_7605,N_7352,N_7371);
xor U7606 (N_7606,N_7417,N_7324);
nand U7607 (N_7607,N_7285,N_7282);
nand U7608 (N_7608,N_7441,N_7219);
nor U7609 (N_7609,N_7263,N_7279);
and U7610 (N_7610,N_7419,N_7217);
or U7611 (N_7611,N_7397,N_7471);
xnor U7612 (N_7612,N_7469,N_7235);
xor U7613 (N_7613,N_7203,N_7350);
or U7614 (N_7614,N_7320,N_7449);
or U7615 (N_7615,N_7224,N_7425);
and U7616 (N_7616,N_7334,N_7476);
or U7617 (N_7617,N_7251,N_7243);
nor U7618 (N_7618,N_7206,N_7465);
or U7619 (N_7619,N_7439,N_7327);
xor U7620 (N_7620,N_7273,N_7437);
or U7621 (N_7621,N_7390,N_7201);
nand U7622 (N_7622,N_7323,N_7349);
and U7623 (N_7623,N_7337,N_7356);
xor U7624 (N_7624,N_7443,N_7363);
nor U7625 (N_7625,N_7365,N_7277);
nor U7626 (N_7626,N_7442,N_7348);
or U7627 (N_7627,N_7416,N_7421);
and U7628 (N_7628,N_7309,N_7259);
nand U7629 (N_7629,N_7484,N_7216);
or U7630 (N_7630,N_7210,N_7291);
or U7631 (N_7631,N_7262,N_7347);
xor U7632 (N_7632,N_7223,N_7364);
xor U7633 (N_7633,N_7326,N_7227);
nand U7634 (N_7634,N_7230,N_7481);
and U7635 (N_7635,N_7494,N_7240);
and U7636 (N_7636,N_7357,N_7499);
xnor U7637 (N_7637,N_7272,N_7460);
xor U7638 (N_7638,N_7375,N_7482);
nor U7639 (N_7639,N_7418,N_7406);
and U7640 (N_7640,N_7253,N_7238);
xnor U7641 (N_7641,N_7339,N_7231);
or U7642 (N_7642,N_7271,N_7306);
nor U7643 (N_7643,N_7477,N_7228);
or U7644 (N_7644,N_7453,N_7490);
nor U7645 (N_7645,N_7314,N_7466);
nor U7646 (N_7646,N_7422,N_7274);
nand U7647 (N_7647,N_7492,N_7229);
and U7648 (N_7648,N_7239,N_7354);
nor U7649 (N_7649,N_7413,N_7451);
and U7650 (N_7650,N_7332,N_7278);
or U7651 (N_7651,N_7300,N_7396);
nor U7652 (N_7652,N_7478,N_7232);
and U7653 (N_7653,N_7338,N_7363);
or U7654 (N_7654,N_7469,N_7285);
and U7655 (N_7655,N_7426,N_7217);
xor U7656 (N_7656,N_7347,N_7413);
xnor U7657 (N_7657,N_7314,N_7336);
or U7658 (N_7658,N_7424,N_7474);
and U7659 (N_7659,N_7219,N_7448);
nand U7660 (N_7660,N_7491,N_7354);
or U7661 (N_7661,N_7441,N_7210);
or U7662 (N_7662,N_7254,N_7375);
xnor U7663 (N_7663,N_7391,N_7499);
nand U7664 (N_7664,N_7444,N_7401);
and U7665 (N_7665,N_7404,N_7345);
nor U7666 (N_7666,N_7422,N_7264);
nand U7667 (N_7667,N_7441,N_7287);
xor U7668 (N_7668,N_7389,N_7368);
nor U7669 (N_7669,N_7278,N_7346);
and U7670 (N_7670,N_7343,N_7380);
xor U7671 (N_7671,N_7437,N_7297);
nand U7672 (N_7672,N_7362,N_7286);
nor U7673 (N_7673,N_7399,N_7260);
nor U7674 (N_7674,N_7266,N_7453);
xnor U7675 (N_7675,N_7294,N_7260);
nand U7676 (N_7676,N_7451,N_7320);
or U7677 (N_7677,N_7377,N_7309);
or U7678 (N_7678,N_7430,N_7286);
or U7679 (N_7679,N_7423,N_7221);
xor U7680 (N_7680,N_7203,N_7392);
nor U7681 (N_7681,N_7441,N_7381);
nor U7682 (N_7682,N_7388,N_7210);
nor U7683 (N_7683,N_7489,N_7246);
xnor U7684 (N_7684,N_7235,N_7343);
xor U7685 (N_7685,N_7262,N_7406);
xnor U7686 (N_7686,N_7485,N_7293);
and U7687 (N_7687,N_7294,N_7335);
nor U7688 (N_7688,N_7404,N_7409);
and U7689 (N_7689,N_7358,N_7234);
nor U7690 (N_7690,N_7459,N_7204);
or U7691 (N_7691,N_7219,N_7205);
or U7692 (N_7692,N_7289,N_7398);
nand U7693 (N_7693,N_7231,N_7289);
or U7694 (N_7694,N_7323,N_7269);
nand U7695 (N_7695,N_7240,N_7390);
nand U7696 (N_7696,N_7415,N_7447);
nand U7697 (N_7697,N_7381,N_7433);
xnor U7698 (N_7698,N_7220,N_7213);
nor U7699 (N_7699,N_7363,N_7313);
nand U7700 (N_7700,N_7357,N_7441);
xnor U7701 (N_7701,N_7434,N_7496);
xor U7702 (N_7702,N_7426,N_7447);
xnor U7703 (N_7703,N_7399,N_7470);
xor U7704 (N_7704,N_7370,N_7350);
xnor U7705 (N_7705,N_7493,N_7271);
nand U7706 (N_7706,N_7251,N_7397);
nand U7707 (N_7707,N_7278,N_7399);
or U7708 (N_7708,N_7269,N_7479);
or U7709 (N_7709,N_7401,N_7390);
xnor U7710 (N_7710,N_7243,N_7234);
and U7711 (N_7711,N_7222,N_7242);
nand U7712 (N_7712,N_7233,N_7348);
or U7713 (N_7713,N_7468,N_7320);
and U7714 (N_7714,N_7253,N_7397);
nand U7715 (N_7715,N_7375,N_7351);
and U7716 (N_7716,N_7211,N_7469);
xor U7717 (N_7717,N_7395,N_7417);
nor U7718 (N_7718,N_7365,N_7369);
or U7719 (N_7719,N_7432,N_7340);
nand U7720 (N_7720,N_7214,N_7363);
xor U7721 (N_7721,N_7383,N_7337);
xnor U7722 (N_7722,N_7204,N_7463);
nand U7723 (N_7723,N_7295,N_7323);
and U7724 (N_7724,N_7237,N_7303);
and U7725 (N_7725,N_7455,N_7477);
nor U7726 (N_7726,N_7484,N_7468);
nor U7727 (N_7727,N_7220,N_7379);
or U7728 (N_7728,N_7494,N_7326);
or U7729 (N_7729,N_7481,N_7270);
nor U7730 (N_7730,N_7303,N_7291);
nand U7731 (N_7731,N_7274,N_7259);
and U7732 (N_7732,N_7489,N_7238);
or U7733 (N_7733,N_7364,N_7486);
nand U7734 (N_7734,N_7456,N_7272);
nand U7735 (N_7735,N_7366,N_7432);
nand U7736 (N_7736,N_7417,N_7413);
and U7737 (N_7737,N_7319,N_7417);
or U7738 (N_7738,N_7290,N_7393);
nand U7739 (N_7739,N_7412,N_7346);
nor U7740 (N_7740,N_7220,N_7486);
nor U7741 (N_7741,N_7240,N_7473);
xnor U7742 (N_7742,N_7331,N_7286);
xor U7743 (N_7743,N_7270,N_7451);
xor U7744 (N_7744,N_7257,N_7324);
or U7745 (N_7745,N_7365,N_7371);
and U7746 (N_7746,N_7448,N_7355);
and U7747 (N_7747,N_7478,N_7292);
nor U7748 (N_7748,N_7260,N_7417);
nor U7749 (N_7749,N_7447,N_7459);
and U7750 (N_7750,N_7380,N_7459);
xnor U7751 (N_7751,N_7267,N_7217);
nor U7752 (N_7752,N_7213,N_7466);
or U7753 (N_7753,N_7245,N_7375);
or U7754 (N_7754,N_7209,N_7294);
xnor U7755 (N_7755,N_7206,N_7491);
nor U7756 (N_7756,N_7407,N_7466);
and U7757 (N_7757,N_7447,N_7233);
or U7758 (N_7758,N_7276,N_7494);
and U7759 (N_7759,N_7468,N_7332);
nor U7760 (N_7760,N_7234,N_7264);
or U7761 (N_7761,N_7304,N_7314);
nand U7762 (N_7762,N_7474,N_7229);
and U7763 (N_7763,N_7342,N_7401);
xnor U7764 (N_7764,N_7440,N_7462);
and U7765 (N_7765,N_7456,N_7209);
nor U7766 (N_7766,N_7486,N_7237);
xor U7767 (N_7767,N_7408,N_7346);
nand U7768 (N_7768,N_7361,N_7308);
or U7769 (N_7769,N_7272,N_7203);
nand U7770 (N_7770,N_7406,N_7287);
xnor U7771 (N_7771,N_7263,N_7345);
nand U7772 (N_7772,N_7238,N_7485);
and U7773 (N_7773,N_7302,N_7333);
nor U7774 (N_7774,N_7312,N_7457);
or U7775 (N_7775,N_7339,N_7254);
or U7776 (N_7776,N_7402,N_7216);
xor U7777 (N_7777,N_7412,N_7444);
nand U7778 (N_7778,N_7280,N_7391);
nand U7779 (N_7779,N_7288,N_7201);
nor U7780 (N_7780,N_7249,N_7222);
xnor U7781 (N_7781,N_7230,N_7409);
nand U7782 (N_7782,N_7383,N_7348);
or U7783 (N_7783,N_7489,N_7366);
or U7784 (N_7784,N_7263,N_7460);
nor U7785 (N_7785,N_7310,N_7377);
xor U7786 (N_7786,N_7379,N_7298);
and U7787 (N_7787,N_7281,N_7280);
or U7788 (N_7788,N_7406,N_7462);
nor U7789 (N_7789,N_7454,N_7263);
xnor U7790 (N_7790,N_7459,N_7375);
xor U7791 (N_7791,N_7230,N_7471);
and U7792 (N_7792,N_7281,N_7341);
nand U7793 (N_7793,N_7205,N_7331);
or U7794 (N_7794,N_7234,N_7203);
or U7795 (N_7795,N_7235,N_7251);
nor U7796 (N_7796,N_7254,N_7221);
and U7797 (N_7797,N_7296,N_7385);
nand U7798 (N_7798,N_7401,N_7298);
xor U7799 (N_7799,N_7380,N_7221);
nor U7800 (N_7800,N_7615,N_7639);
xor U7801 (N_7801,N_7627,N_7747);
and U7802 (N_7802,N_7735,N_7608);
xnor U7803 (N_7803,N_7515,N_7713);
or U7804 (N_7804,N_7611,N_7626);
or U7805 (N_7805,N_7507,N_7767);
or U7806 (N_7806,N_7592,N_7762);
nand U7807 (N_7807,N_7633,N_7622);
xor U7808 (N_7808,N_7560,N_7561);
or U7809 (N_7809,N_7524,N_7678);
and U7810 (N_7810,N_7728,N_7662);
and U7811 (N_7811,N_7787,N_7701);
nand U7812 (N_7812,N_7771,N_7697);
nand U7813 (N_7813,N_7518,N_7580);
or U7814 (N_7814,N_7573,N_7687);
and U7815 (N_7815,N_7621,N_7780);
nand U7816 (N_7816,N_7527,N_7690);
and U7817 (N_7817,N_7535,N_7723);
and U7818 (N_7818,N_7770,N_7731);
xnor U7819 (N_7819,N_7756,N_7794);
nor U7820 (N_7820,N_7636,N_7638);
and U7821 (N_7821,N_7676,N_7749);
or U7822 (N_7822,N_7606,N_7721);
and U7823 (N_7823,N_7763,N_7716);
nand U7824 (N_7824,N_7640,N_7620);
nor U7825 (N_7825,N_7565,N_7593);
xnor U7826 (N_7826,N_7665,N_7536);
xor U7827 (N_7827,N_7698,N_7790);
or U7828 (N_7828,N_7655,N_7543);
nor U7829 (N_7829,N_7774,N_7705);
or U7830 (N_7830,N_7623,N_7738);
nor U7831 (N_7831,N_7712,N_7526);
and U7832 (N_7832,N_7596,N_7793);
xnor U7833 (N_7833,N_7776,N_7558);
and U7834 (N_7834,N_7613,N_7521);
nor U7835 (N_7835,N_7643,N_7672);
and U7836 (N_7836,N_7778,N_7600);
and U7837 (N_7837,N_7538,N_7691);
and U7838 (N_7838,N_7694,N_7757);
or U7839 (N_7839,N_7579,N_7508);
and U7840 (N_7840,N_7556,N_7707);
nand U7841 (N_7841,N_7583,N_7619);
xor U7842 (N_7842,N_7797,N_7519);
nand U7843 (N_7843,N_7570,N_7542);
or U7844 (N_7844,N_7645,N_7750);
nand U7845 (N_7845,N_7704,N_7659);
nand U7846 (N_7846,N_7730,N_7562);
and U7847 (N_7847,N_7717,N_7520);
or U7848 (N_7848,N_7541,N_7796);
nor U7849 (N_7849,N_7513,N_7635);
and U7850 (N_7850,N_7737,N_7586);
xor U7851 (N_7851,N_7739,N_7604);
xnor U7852 (N_7852,N_7700,N_7599);
nor U7853 (N_7853,N_7710,N_7617);
or U7854 (N_7854,N_7528,N_7792);
or U7855 (N_7855,N_7540,N_7525);
or U7856 (N_7856,N_7715,N_7504);
or U7857 (N_7857,N_7624,N_7641);
xor U7858 (N_7858,N_7688,N_7696);
or U7859 (N_7859,N_7564,N_7501);
nor U7860 (N_7860,N_7637,N_7722);
and U7861 (N_7861,N_7695,N_7512);
xnor U7862 (N_7862,N_7625,N_7719);
and U7863 (N_7863,N_7663,N_7503);
nor U7864 (N_7864,N_7741,N_7648);
nand U7865 (N_7865,N_7725,N_7754);
and U7866 (N_7866,N_7755,N_7631);
xnor U7867 (N_7867,N_7582,N_7555);
or U7868 (N_7868,N_7514,N_7628);
or U7869 (N_7869,N_7609,N_7572);
xnor U7870 (N_7870,N_7791,N_7709);
nor U7871 (N_7871,N_7642,N_7670);
nor U7872 (N_7872,N_7759,N_7656);
and U7873 (N_7873,N_7733,N_7557);
nor U7874 (N_7874,N_7516,N_7782);
nand U7875 (N_7875,N_7603,N_7761);
nand U7876 (N_7876,N_7506,N_7587);
and U7877 (N_7877,N_7554,N_7783);
or U7878 (N_7878,N_7746,N_7509);
and U7879 (N_7879,N_7553,N_7764);
nor U7880 (N_7880,N_7772,N_7657);
xor U7881 (N_7881,N_7781,N_7567);
nor U7882 (N_7882,N_7758,N_7575);
nor U7883 (N_7883,N_7727,N_7714);
and U7884 (N_7884,N_7658,N_7597);
and U7885 (N_7885,N_7769,N_7534);
and U7886 (N_7886,N_7708,N_7692);
xnor U7887 (N_7887,N_7584,N_7748);
xor U7888 (N_7888,N_7724,N_7532);
nand U7889 (N_7889,N_7594,N_7616);
or U7890 (N_7890,N_7726,N_7667);
or U7891 (N_7891,N_7706,N_7753);
or U7892 (N_7892,N_7510,N_7589);
nor U7893 (N_7893,N_7779,N_7686);
or U7894 (N_7894,N_7588,N_7644);
or U7895 (N_7895,N_7568,N_7544);
and U7896 (N_7896,N_7559,N_7675);
nor U7897 (N_7897,N_7703,N_7547);
nand U7898 (N_7898,N_7654,N_7683);
or U7899 (N_7899,N_7546,N_7786);
or U7900 (N_7900,N_7777,N_7743);
xnor U7901 (N_7901,N_7751,N_7785);
and U7902 (N_7902,N_7653,N_7505);
and U7903 (N_7903,N_7685,N_7566);
or U7904 (N_7904,N_7732,N_7673);
nor U7905 (N_7905,N_7798,N_7614);
nand U7906 (N_7906,N_7539,N_7799);
xnor U7907 (N_7907,N_7548,N_7590);
xor U7908 (N_7908,N_7650,N_7552);
nand U7909 (N_7909,N_7775,N_7680);
and U7910 (N_7910,N_7684,N_7517);
nand U7911 (N_7911,N_7699,N_7634);
and U7912 (N_7912,N_7666,N_7742);
or U7913 (N_7913,N_7789,N_7549);
xor U7914 (N_7914,N_7577,N_7736);
or U7915 (N_7915,N_7618,N_7711);
or U7916 (N_7916,N_7569,N_7647);
nor U7917 (N_7917,N_7578,N_7661);
or U7918 (N_7918,N_7664,N_7605);
or U7919 (N_7919,N_7632,N_7682);
or U7920 (N_7920,N_7766,N_7740);
or U7921 (N_7921,N_7760,N_7537);
or U7922 (N_7922,N_7500,N_7550);
or U7923 (N_7923,N_7612,N_7660);
nor U7924 (N_7924,N_7563,N_7522);
and U7925 (N_7925,N_7551,N_7744);
nor U7926 (N_7926,N_7523,N_7649);
xor U7927 (N_7927,N_7545,N_7669);
nor U7928 (N_7928,N_7595,N_7574);
xnor U7929 (N_7929,N_7598,N_7630);
nor U7930 (N_7930,N_7530,N_7689);
xnor U7931 (N_7931,N_7502,N_7702);
or U7932 (N_7932,N_7677,N_7581);
xnor U7933 (N_7933,N_7652,N_7718);
nor U7934 (N_7934,N_7768,N_7765);
xor U7935 (N_7935,N_7720,N_7529);
xor U7936 (N_7936,N_7752,N_7674);
or U7937 (N_7937,N_7734,N_7629);
nor U7938 (N_7938,N_7671,N_7610);
or U7939 (N_7939,N_7602,N_7668);
nand U7940 (N_7940,N_7646,N_7601);
xor U7941 (N_7941,N_7591,N_7533);
xor U7942 (N_7942,N_7773,N_7511);
and U7943 (N_7943,N_7571,N_7531);
nor U7944 (N_7944,N_7788,N_7607);
and U7945 (N_7945,N_7681,N_7585);
xnor U7946 (N_7946,N_7795,N_7693);
and U7947 (N_7947,N_7576,N_7729);
xor U7948 (N_7948,N_7651,N_7745);
nand U7949 (N_7949,N_7679,N_7784);
xor U7950 (N_7950,N_7621,N_7660);
xor U7951 (N_7951,N_7626,N_7700);
and U7952 (N_7952,N_7618,N_7595);
and U7953 (N_7953,N_7599,N_7531);
and U7954 (N_7954,N_7651,N_7524);
or U7955 (N_7955,N_7778,N_7664);
and U7956 (N_7956,N_7762,N_7519);
nand U7957 (N_7957,N_7590,N_7612);
or U7958 (N_7958,N_7759,N_7701);
nor U7959 (N_7959,N_7642,N_7733);
and U7960 (N_7960,N_7560,N_7533);
xnor U7961 (N_7961,N_7632,N_7587);
xnor U7962 (N_7962,N_7632,N_7654);
or U7963 (N_7963,N_7527,N_7731);
xor U7964 (N_7964,N_7628,N_7672);
nor U7965 (N_7965,N_7739,N_7777);
nand U7966 (N_7966,N_7765,N_7713);
nor U7967 (N_7967,N_7628,N_7778);
nand U7968 (N_7968,N_7538,N_7522);
or U7969 (N_7969,N_7672,N_7644);
nand U7970 (N_7970,N_7774,N_7749);
xnor U7971 (N_7971,N_7770,N_7727);
nor U7972 (N_7972,N_7546,N_7781);
or U7973 (N_7973,N_7699,N_7711);
and U7974 (N_7974,N_7694,N_7678);
or U7975 (N_7975,N_7582,N_7651);
or U7976 (N_7976,N_7683,N_7731);
or U7977 (N_7977,N_7518,N_7582);
or U7978 (N_7978,N_7514,N_7606);
or U7979 (N_7979,N_7677,N_7557);
nor U7980 (N_7980,N_7672,N_7694);
nor U7981 (N_7981,N_7509,N_7553);
xnor U7982 (N_7982,N_7504,N_7695);
nand U7983 (N_7983,N_7714,N_7728);
nor U7984 (N_7984,N_7514,N_7799);
and U7985 (N_7985,N_7664,N_7723);
and U7986 (N_7986,N_7581,N_7551);
nand U7987 (N_7987,N_7650,N_7748);
and U7988 (N_7988,N_7556,N_7704);
or U7989 (N_7989,N_7713,N_7501);
nor U7990 (N_7990,N_7692,N_7726);
or U7991 (N_7991,N_7618,N_7672);
nand U7992 (N_7992,N_7524,N_7696);
nand U7993 (N_7993,N_7760,N_7685);
xor U7994 (N_7994,N_7538,N_7721);
nor U7995 (N_7995,N_7570,N_7576);
nor U7996 (N_7996,N_7644,N_7776);
or U7997 (N_7997,N_7654,N_7740);
nor U7998 (N_7998,N_7794,N_7560);
nand U7999 (N_7999,N_7667,N_7717);
nor U8000 (N_8000,N_7659,N_7626);
nor U8001 (N_8001,N_7504,N_7690);
xor U8002 (N_8002,N_7649,N_7505);
and U8003 (N_8003,N_7753,N_7746);
nand U8004 (N_8004,N_7670,N_7580);
xor U8005 (N_8005,N_7507,N_7526);
and U8006 (N_8006,N_7783,N_7711);
nor U8007 (N_8007,N_7703,N_7713);
nor U8008 (N_8008,N_7565,N_7736);
and U8009 (N_8009,N_7603,N_7758);
or U8010 (N_8010,N_7719,N_7676);
nor U8011 (N_8011,N_7674,N_7552);
and U8012 (N_8012,N_7701,N_7665);
nand U8013 (N_8013,N_7763,N_7512);
xnor U8014 (N_8014,N_7559,N_7782);
nor U8015 (N_8015,N_7552,N_7633);
xor U8016 (N_8016,N_7545,N_7732);
xor U8017 (N_8017,N_7758,N_7631);
or U8018 (N_8018,N_7553,N_7557);
nand U8019 (N_8019,N_7791,N_7741);
xnor U8020 (N_8020,N_7741,N_7793);
xnor U8021 (N_8021,N_7556,N_7601);
or U8022 (N_8022,N_7659,N_7644);
nor U8023 (N_8023,N_7597,N_7769);
nor U8024 (N_8024,N_7614,N_7554);
or U8025 (N_8025,N_7626,N_7548);
xor U8026 (N_8026,N_7611,N_7667);
xnor U8027 (N_8027,N_7694,N_7549);
or U8028 (N_8028,N_7655,N_7748);
or U8029 (N_8029,N_7742,N_7691);
xor U8030 (N_8030,N_7721,N_7577);
nor U8031 (N_8031,N_7713,N_7574);
nor U8032 (N_8032,N_7632,N_7663);
and U8033 (N_8033,N_7659,N_7645);
xnor U8034 (N_8034,N_7692,N_7694);
and U8035 (N_8035,N_7542,N_7697);
nand U8036 (N_8036,N_7799,N_7569);
and U8037 (N_8037,N_7584,N_7588);
xor U8038 (N_8038,N_7544,N_7507);
nor U8039 (N_8039,N_7784,N_7591);
nor U8040 (N_8040,N_7773,N_7792);
and U8041 (N_8041,N_7572,N_7698);
nor U8042 (N_8042,N_7500,N_7520);
nand U8043 (N_8043,N_7536,N_7541);
nand U8044 (N_8044,N_7607,N_7587);
xnor U8045 (N_8045,N_7688,N_7797);
and U8046 (N_8046,N_7543,N_7664);
and U8047 (N_8047,N_7613,N_7665);
xor U8048 (N_8048,N_7644,N_7679);
nand U8049 (N_8049,N_7726,N_7589);
and U8050 (N_8050,N_7634,N_7586);
xnor U8051 (N_8051,N_7512,N_7778);
and U8052 (N_8052,N_7755,N_7649);
xor U8053 (N_8053,N_7631,N_7645);
xor U8054 (N_8054,N_7575,N_7746);
xor U8055 (N_8055,N_7695,N_7658);
and U8056 (N_8056,N_7686,N_7604);
nor U8057 (N_8057,N_7718,N_7684);
nand U8058 (N_8058,N_7663,N_7643);
xnor U8059 (N_8059,N_7765,N_7676);
nand U8060 (N_8060,N_7670,N_7669);
nor U8061 (N_8061,N_7749,N_7572);
or U8062 (N_8062,N_7539,N_7506);
nand U8063 (N_8063,N_7643,N_7754);
nand U8064 (N_8064,N_7503,N_7771);
xnor U8065 (N_8065,N_7601,N_7606);
nand U8066 (N_8066,N_7798,N_7774);
nor U8067 (N_8067,N_7559,N_7672);
nand U8068 (N_8068,N_7615,N_7737);
xnor U8069 (N_8069,N_7669,N_7747);
or U8070 (N_8070,N_7667,N_7624);
and U8071 (N_8071,N_7572,N_7579);
nor U8072 (N_8072,N_7690,N_7507);
or U8073 (N_8073,N_7727,N_7678);
or U8074 (N_8074,N_7506,N_7659);
nor U8075 (N_8075,N_7586,N_7739);
or U8076 (N_8076,N_7511,N_7759);
xnor U8077 (N_8077,N_7524,N_7570);
nor U8078 (N_8078,N_7534,N_7553);
nor U8079 (N_8079,N_7658,N_7553);
nor U8080 (N_8080,N_7577,N_7724);
or U8081 (N_8081,N_7737,N_7690);
nand U8082 (N_8082,N_7539,N_7558);
or U8083 (N_8083,N_7719,N_7600);
nor U8084 (N_8084,N_7698,N_7750);
xor U8085 (N_8085,N_7663,N_7782);
or U8086 (N_8086,N_7526,N_7523);
xor U8087 (N_8087,N_7681,N_7623);
or U8088 (N_8088,N_7713,N_7577);
or U8089 (N_8089,N_7649,N_7662);
nand U8090 (N_8090,N_7570,N_7608);
or U8091 (N_8091,N_7562,N_7724);
or U8092 (N_8092,N_7768,N_7524);
or U8093 (N_8093,N_7762,N_7643);
nand U8094 (N_8094,N_7586,N_7544);
and U8095 (N_8095,N_7707,N_7690);
nor U8096 (N_8096,N_7508,N_7515);
xnor U8097 (N_8097,N_7526,N_7711);
nor U8098 (N_8098,N_7782,N_7685);
nand U8099 (N_8099,N_7719,N_7648);
nor U8100 (N_8100,N_8098,N_7958);
xnor U8101 (N_8101,N_8078,N_7932);
xnor U8102 (N_8102,N_7972,N_7855);
or U8103 (N_8103,N_7931,N_7956);
or U8104 (N_8104,N_8028,N_7815);
nand U8105 (N_8105,N_7869,N_7882);
or U8106 (N_8106,N_7953,N_7935);
or U8107 (N_8107,N_7888,N_8045);
xor U8108 (N_8108,N_7921,N_7933);
nand U8109 (N_8109,N_7996,N_8038);
nand U8110 (N_8110,N_7986,N_7893);
or U8111 (N_8111,N_7974,N_7963);
and U8112 (N_8112,N_7988,N_8096);
and U8113 (N_8113,N_8002,N_7802);
or U8114 (N_8114,N_8030,N_7993);
xor U8115 (N_8115,N_7891,N_7982);
and U8116 (N_8116,N_8073,N_7871);
nand U8117 (N_8117,N_7910,N_8026);
xnor U8118 (N_8118,N_8029,N_8095);
and U8119 (N_8119,N_8075,N_8094);
nand U8120 (N_8120,N_7889,N_8072);
nand U8121 (N_8121,N_7987,N_7989);
or U8122 (N_8122,N_8004,N_8008);
xnor U8123 (N_8123,N_8065,N_8074);
nor U8124 (N_8124,N_8016,N_7905);
or U8125 (N_8125,N_8060,N_7945);
nand U8126 (N_8126,N_7844,N_7890);
or U8127 (N_8127,N_8067,N_8093);
nor U8128 (N_8128,N_8090,N_7922);
nand U8129 (N_8129,N_7851,N_7809);
nand U8130 (N_8130,N_7915,N_8013);
or U8131 (N_8131,N_7954,N_7818);
nand U8132 (N_8132,N_7822,N_7824);
nor U8133 (N_8133,N_7941,N_7929);
and U8134 (N_8134,N_8037,N_7966);
nand U8135 (N_8135,N_7842,N_7816);
or U8136 (N_8136,N_7957,N_7858);
nor U8137 (N_8137,N_7947,N_8087);
xnor U8138 (N_8138,N_7876,N_7838);
and U8139 (N_8139,N_8027,N_7829);
nor U8140 (N_8140,N_7857,N_8050);
and U8141 (N_8141,N_7843,N_7961);
and U8142 (N_8142,N_8024,N_8070);
and U8143 (N_8143,N_7899,N_8019);
xor U8144 (N_8144,N_8066,N_8018);
xnor U8145 (N_8145,N_8035,N_7914);
nor U8146 (N_8146,N_7942,N_7997);
or U8147 (N_8147,N_7943,N_7845);
xnor U8148 (N_8148,N_7823,N_7885);
nor U8149 (N_8149,N_7859,N_7967);
nand U8150 (N_8150,N_7901,N_7813);
and U8151 (N_8151,N_7868,N_7965);
or U8152 (N_8152,N_8063,N_7902);
xnor U8153 (N_8153,N_7837,N_7970);
and U8154 (N_8154,N_8057,N_8000);
xor U8155 (N_8155,N_7917,N_8068);
and U8156 (N_8156,N_7831,N_8079);
or U8157 (N_8157,N_8025,N_7841);
or U8158 (N_8158,N_8056,N_8058);
nor U8159 (N_8159,N_7949,N_7919);
or U8160 (N_8160,N_7894,N_8033);
nor U8161 (N_8161,N_7826,N_7850);
nor U8162 (N_8162,N_7811,N_7976);
or U8163 (N_8163,N_7950,N_7923);
nand U8164 (N_8164,N_7960,N_8084);
nor U8165 (N_8165,N_7810,N_7969);
nor U8166 (N_8166,N_8005,N_7830);
nand U8167 (N_8167,N_7930,N_7825);
nand U8168 (N_8168,N_8046,N_7833);
xnor U8169 (N_8169,N_7918,N_7807);
xnor U8170 (N_8170,N_8040,N_7865);
nand U8171 (N_8171,N_7938,N_7820);
or U8172 (N_8172,N_8048,N_8007);
nand U8173 (N_8173,N_7827,N_8032);
and U8174 (N_8174,N_7806,N_8015);
xor U8175 (N_8175,N_8097,N_7874);
and U8176 (N_8176,N_7994,N_7946);
nand U8177 (N_8177,N_8061,N_7962);
or U8178 (N_8178,N_7854,N_7814);
and U8179 (N_8179,N_7911,N_8031);
nand U8180 (N_8180,N_7959,N_8051);
xor U8181 (N_8181,N_8092,N_8088);
nor U8182 (N_8182,N_7978,N_8089);
nand U8183 (N_8183,N_8017,N_7896);
or U8184 (N_8184,N_7800,N_8043);
or U8185 (N_8185,N_8064,N_8099);
nand U8186 (N_8186,N_7909,N_7999);
nor U8187 (N_8187,N_7846,N_8020);
nor U8188 (N_8188,N_7903,N_7980);
nand U8189 (N_8189,N_7895,N_7981);
nor U8190 (N_8190,N_8021,N_7975);
nand U8191 (N_8191,N_8085,N_7887);
and U8192 (N_8192,N_7808,N_7928);
or U8193 (N_8193,N_7883,N_7848);
and U8194 (N_8194,N_8059,N_7900);
or U8195 (N_8195,N_7944,N_7998);
nand U8196 (N_8196,N_7875,N_7812);
nor U8197 (N_8197,N_7924,N_8076);
and U8198 (N_8198,N_8052,N_7860);
nand U8199 (N_8199,N_7904,N_7867);
nand U8200 (N_8200,N_7934,N_8036);
nor U8201 (N_8201,N_7920,N_8022);
or U8202 (N_8202,N_7936,N_7955);
nor U8203 (N_8203,N_7864,N_7907);
or U8204 (N_8204,N_8091,N_8049);
nand U8205 (N_8205,N_7886,N_7853);
nand U8206 (N_8206,N_7995,N_7951);
xnor U8207 (N_8207,N_7912,N_7805);
or U8208 (N_8208,N_7897,N_8080);
xnor U8209 (N_8209,N_8055,N_7872);
or U8210 (N_8210,N_8083,N_7863);
nor U8211 (N_8211,N_8011,N_7964);
xnor U8212 (N_8212,N_7906,N_7916);
nor U8213 (N_8213,N_7925,N_7881);
xor U8214 (N_8214,N_7861,N_7801);
and U8215 (N_8215,N_7832,N_7852);
nand U8216 (N_8216,N_8010,N_7836);
and U8217 (N_8217,N_7984,N_8034);
nor U8218 (N_8218,N_8062,N_7939);
and U8219 (N_8219,N_7979,N_7856);
nand U8220 (N_8220,N_8014,N_7849);
or U8221 (N_8221,N_7977,N_7968);
or U8222 (N_8222,N_7880,N_7834);
xor U8223 (N_8223,N_7819,N_8039);
xor U8224 (N_8224,N_7908,N_7804);
and U8225 (N_8225,N_8053,N_7927);
or U8226 (N_8226,N_7847,N_8042);
and U8227 (N_8227,N_7991,N_7866);
or U8228 (N_8228,N_8071,N_8054);
xnor U8229 (N_8229,N_8082,N_8003);
nor U8230 (N_8230,N_8044,N_7948);
nand U8231 (N_8231,N_7990,N_8006);
nand U8232 (N_8232,N_7971,N_7879);
xor U8233 (N_8233,N_7870,N_7839);
or U8234 (N_8234,N_8077,N_7878);
and U8235 (N_8235,N_8012,N_8009);
nor U8236 (N_8236,N_7973,N_7892);
nand U8237 (N_8237,N_7877,N_8047);
or U8238 (N_8238,N_7828,N_7862);
and U8239 (N_8239,N_7940,N_7952);
xnor U8240 (N_8240,N_7926,N_8086);
and U8241 (N_8241,N_8069,N_7898);
xnor U8242 (N_8242,N_7835,N_8023);
xnor U8243 (N_8243,N_8041,N_7884);
or U8244 (N_8244,N_7803,N_8081);
nand U8245 (N_8245,N_7873,N_7821);
xor U8246 (N_8246,N_8001,N_7817);
and U8247 (N_8247,N_7992,N_7985);
nand U8248 (N_8248,N_7983,N_7840);
xnor U8249 (N_8249,N_7937,N_7913);
or U8250 (N_8250,N_7955,N_8020);
xnor U8251 (N_8251,N_7810,N_7906);
nand U8252 (N_8252,N_7890,N_8040);
and U8253 (N_8253,N_7977,N_7871);
nor U8254 (N_8254,N_7964,N_8002);
and U8255 (N_8255,N_8011,N_8074);
xnor U8256 (N_8256,N_7874,N_7853);
or U8257 (N_8257,N_7875,N_7831);
xnor U8258 (N_8258,N_8054,N_7822);
nand U8259 (N_8259,N_7837,N_7821);
nor U8260 (N_8260,N_7968,N_8098);
xnor U8261 (N_8261,N_8015,N_7882);
and U8262 (N_8262,N_8032,N_7969);
nor U8263 (N_8263,N_7826,N_7893);
and U8264 (N_8264,N_8043,N_8059);
xnor U8265 (N_8265,N_8011,N_8008);
and U8266 (N_8266,N_7967,N_7879);
or U8267 (N_8267,N_7856,N_7951);
xnor U8268 (N_8268,N_7843,N_7811);
xnor U8269 (N_8269,N_8088,N_8022);
or U8270 (N_8270,N_7825,N_7959);
and U8271 (N_8271,N_7975,N_7915);
and U8272 (N_8272,N_8039,N_7850);
nand U8273 (N_8273,N_7879,N_8059);
nor U8274 (N_8274,N_7812,N_7945);
or U8275 (N_8275,N_7954,N_7861);
xor U8276 (N_8276,N_7992,N_7916);
or U8277 (N_8277,N_7968,N_7883);
nor U8278 (N_8278,N_7871,N_7923);
nor U8279 (N_8279,N_8066,N_8050);
nor U8280 (N_8280,N_8019,N_8079);
nor U8281 (N_8281,N_7867,N_8011);
nand U8282 (N_8282,N_7971,N_7880);
xnor U8283 (N_8283,N_8079,N_7956);
nand U8284 (N_8284,N_8074,N_7802);
and U8285 (N_8285,N_8000,N_7999);
nor U8286 (N_8286,N_8087,N_7894);
xor U8287 (N_8287,N_7884,N_7819);
or U8288 (N_8288,N_7917,N_7983);
nor U8289 (N_8289,N_7835,N_7992);
or U8290 (N_8290,N_7958,N_7940);
and U8291 (N_8291,N_7811,N_8098);
nor U8292 (N_8292,N_7981,N_7823);
xor U8293 (N_8293,N_8047,N_7802);
or U8294 (N_8294,N_7828,N_7976);
xor U8295 (N_8295,N_7952,N_7823);
nor U8296 (N_8296,N_8024,N_7994);
or U8297 (N_8297,N_7889,N_8085);
or U8298 (N_8298,N_7881,N_7815);
nand U8299 (N_8299,N_7936,N_7886);
nor U8300 (N_8300,N_7856,N_7931);
nor U8301 (N_8301,N_8026,N_7858);
nor U8302 (N_8302,N_7988,N_7934);
or U8303 (N_8303,N_7856,N_7946);
and U8304 (N_8304,N_7957,N_8018);
xor U8305 (N_8305,N_7888,N_8015);
nor U8306 (N_8306,N_7808,N_7817);
xnor U8307 (N_8307,N_7872,N_7988);
and U8308 (N_8308,N_7949,N_8044);
nand U8309 (N_8309,N_7878,N_8093);
xor U8310 (N_8310,N_8062,N_7989);
nand U8311 (N_8311,N_7875,N_7901);
and U8312 (N_8312,N_7902,N_7848);
nor U8313 (N_8313,N_7844,N_7907);
or U8314 (N_8314,N_8077,N_7854);
nand U8315 (N_8315,N_7818,N_7909);
nand U8316 (N_8316,N_8078,N_7821);
nor U8317 (N_8317,N_8022,N_8014);
nor U8318 (N_8318,N_8053,N_8019);
or U8319 (N_8319,N_8092,N_7869);
nand U8320 (N_8320,N_8057,N_8095);
nand U8321 (N_8321,N_8021,N_8034);
nand U8322 (N_8322,N_8009,N_7877);
xnor U8323 (N_8323,N_7803,N_7816);
xnor U8324 (N_8324,N_7903,N_7899);
or U8325 (N_8325,N_7897,N_7832);
nand U8326 (N_8326,N_7829,N_7948);
and U8327 (N_8327,N_7964,N_7867);
xor U8328 (N_8328,N_8064,N_7815);
and U8329 (N_8329,N_7878,N_8041);
or U8330 (N_8330,N_8067,N_7952);
or U8331 (N_8331,N_7965,N_8040);
nand U8332 (N_8332,N_8074,N_7974);
nand U8333 (N_8333,N_7991,N_7879);
nor U8334 (N_8334,N_7825,N_7951);
nor U8335 (N_8335,N_7929,N_8064);
and U8336 (N_8336,N_8002,N_7806);
and U8337 (N_8337,N_8014,N_7962);
nor U8338 (N_8338,N_7892,N_7875);
and U8339 (N_8339,N_7937,N_7821);
or U8340 (N_8340,N_8010,N_7903);
nor U8341 (N_8341,N_7803,N_7842);
nor U8342 (N_8342,N_8049,N_8053);
and U8343 (N_8343,N_7950,N_8050);
xor U8344 (N_8344,N_7877,N_7980);
or U8345 (N_8345,N_8022,N_7860);
nand U8346 (N_8346,N_7985,N_8021);
or U8347 (N_8347,N_8055,N_7935);
and U8348 (N_8348,N_8075,N_8043);
and U8349 (N_8349,N_7924,N_8059);
and U8350 (N_8350,N_7837,N_7860);
and U8351 (N_8351,N_8081,N_7868);
and U8352 (N_8352,N_7951,N_7832);
nor U8353 (N_8353,N_7961,N_8008);
and U8354 (N_8354,N_7952,N_7943);
nor U8355 (N_8355,N_7839,N_8051);
nand U8356 (N_8356,N_8016,N_7901);
and U8357 (N_8357,N_8032,N_7918);
or U8358 (N_8358,N_7833,N_7850);
and U8359 (N_8359,N_7894,N_8026);
and U8360 (N_8360,N_8085,N_8025);
xor U8361 (N_8361,N_8049,N_7898);
and U8362 (N_8362,N_7822,N_7944);
xor U8363 (N_8363,N_7932,N_7951);
nor U8364 (N_8364,N_7970,N_8040);
nor U8365 (N_8365,N_7952,N_7862);
or U8366 (N_8366,N_7801,N_7931);
nor U8367 (N_8367,N_7849,N_8098);
nor U8368 (N_8368,N_7987,N_7882);
or U8369 (N_8369,N_7917,N_7966);
nor U8370 (N_8370,N_7922,N_7916);
or U8371 (N_8371,N_7974,N_8079);
nand U8372 (N_8372,N_7851,N_8005);
nor U8373 (N_8373,N_7977,N_7824);
and U8374 (N_8374,N_7926,N_7961);
and U8375 (N_8375,N_7841,N_7907);
nor U8376 (N_8376,N_8017,N_7869);
nand U8377 (N_8377,N_8011,N_8010);
nor U8378 (N_8378,N_7950,N_7962);
and U8379 (N_8379,N_8066,N_7873);
and U8380 (N_8380,N_8014,N_8054);
nor U8381 (N_8381,N_7986,N_8077);
or U8382 (N_8382,N_8086,N_7859);
or U8383 (N_8383,N_7863,N_7897);
and U8384 (N_8384,N_7936,N_8073);
or U8385 (N_8385,N_8091,N_7993);
or U8386 (N_8386,N_7863,N_8068);
or U8387 (N_8387,N_8005,N_7843);
and U8388 (N_8388,N_8042,N_7974);
nor U8389 (N_8389,N_8096,N_7835);
xor U8390 (N_8390,N_8009,N_8095);
or U8391 (N_8391,N_7841,N_7902);
xor U8392 (N_8392,N_7863,N_7941);
and U8393 (N_8393,N_8034,N_7824);
or U8394 (N_8394,N_8074,N_7844);
nand U8395 (N_8395,N_7843,N_7967);
and U8396 (N_8396,N_7895,N_7941);
nor U8397 (N_8397,N_7885,N_7934);
or U8398 (N_8398,N_7928,N_8044);
nand U8399 (N_8399,N_7960,N_8073);
nor U8400 (N_8400,N_8121,N_8300);
xor U8401 (N_8401,N_8151,N_8340);
xnor U8402 (N_8402,N_8264,N_8177);
or U8403 (N_8403,N_8172,N_8329);
and U8404 (N_8404,N_8262,N_8323);
nor U8405 (N_8405,N_8396,N_8245);
nand U8406 (N_8406,N_8307,N_8215);
xor U8407 (N_8407,N_8350,N_8252);
and U8408 (N_8408,N_8206,N_8283);
nor U8409 (N_8409,N_8312,N_8140);
and U8410 (N_8410,N_8389,N_8237);
and U8411 (N_8411,N_8311,N_8325);
nor U8412 (N_8412,N_8213,N_8296);
nor U8413 (N_8413,N_8136,N_8362);
or U8414 (N_8414,N_8379,N_8182);
or U8415 (N_8415,N_8327,N_8175);
or U8416 (N_8416,N_8265,N_8193);
xnor U8417 (N_8417,N_8103,N_8277);
or U8418 (N_8418,N_8272,N_8290);
and U8419 (N_8419,N_8124,N_8345);
and U8420 (N_8420,N_8288,N_8184);
nand U8421 (N_8421,N_8358,N_8348);
nor U8422 (N_8422,N_8114,N_8241);
nand U8423 (N_8423,N_8236,N_8118);
or U8424 (N_8424,N_8351,N_8143);
nand U8425 (N_8425,N_8149,N_8212);
and U8426 (N_8426,N_8301,N_8273);
and U8427 (N_8427,N_8353,N_8111);
and U8428 (N_8428,N_8235,N_8218);
nand U8429 (N_8429,N_8145,N_8195);
and U8430 (N_8430,N_8119,N_8382);
xnor U8431 (N_8431,N_8208,N_8308);
nor U8432 (N_8432,N_8170,N_8134);
and U8433 (N_8433,N_8132,N_8357);
nor U8434 (N_8434,N_8123,N_8216);
xnor U8435 (N_8435,N_8356,N_8392);
and U8436 (N_8436,N_8152,N_8336);
xnor U8437 (N_8437,N_8234,N_8228);
or U8438 (N_8438,N_8322,N_8319);
nand U8439 (N_8439,N_8219,N_8303);
xnor U8440 (N_8440,N_8183,N_8233);
nand U8441 (N_8441,N_8326,N_8238);
or U8442 (N_8442,N_8375,N_8243);
nor U8443 (N_8443,N_8203,N_8125);
nand U8444 (N_8444,N_8157,N_8279);
and U8445 (N_8445,N_8248,N_8302);
xnor U8446 (N_8446,N_8109,N_8332);
nor U8447 (N_8447,N_8287,N_8342);
nand U8448 (N_8448,N_8260,N_8102);
or U8449 (N_8449,N_8129,N_8160);
and U8450 (N_8450,N_8221,N_8158);
or U8451 (N_8451,N_8310,N_8131);
nand U8452 (N_8452,N_8168,N_8202);
xor U8453 (N_8453,N_8155,N_8197);
or U8454 (N_8454,N_8115,N_8179);
nand U8455 (N_8455,N_8343,N_8328);
or U8456 (N_8456,N_8341,N_8188);
and U8457 (N_8457,N_8280,N_8191);
and U8458 (N_8458,N_8333,N_8331);
nor U8459 (N_8459,N_8347,N_8286);
nor U8460 (N_8460,N_8104,N_8377);
nor U8461 (N_8461,N_8253,N_8196);
xor U8462 (N_8462,N_8167,N_8314);
nand U8463 (N_8463,N_8176,N_8293);
xnor U8464 (N_8464,N_8316,N_8222);
or U8465 (N_8465,N_8189,N_8205);
or U8466 (N_8466,N_8299,N_8144);
or U8467 (N_8467,N_8128,N_8164);
xnor U8468 (N_8468,N_8363,N_8291);
nand U8469 (N_8469,N_8261,N_8365);
nand U8470 (N_8470,N_8126,N_8180);
nand U8471 (N_8471,N_8366,N_8214);
nor U8472 (N_8472,N_8186,N_8395);
or U8473 (N_8473,N_8297,N_8313);
and U8474 (N_8474,N_8204,N_8394);
xor U8475 (N_8475,N_8122,N_8185);
or U8476 (N_8476,N_8330,N_8258);
xnor U8477 (N_8477,N_8199,N_8159);
nor U8478 (N_8478,N_8226,N_8100);
or U8479 (N_8479,N_8110,N_8268);
nor U8480 (N_8480,N_8225,N_8156);
and U8481 (N_8481,N_8106,N_8266);
nor U8482 (N_8482,N_8278,N_8148);
nor U8483 (N_8483,N_8230,N_8372);
nor U8484 (N_8484,N_8117,N_8255);
xor U8485 (N_8485,N_8380,N_8239);
nand U8486 (N_8486,N_8387,N_8281);
or U8487 (N_8487,N_8137,N_8178);
nand U8488 (N_8488,N_8232,N_8116);
xor U8489 (N_8489,N_8139,N_8173);
and U8490 (N_8490,N_8393,N_8108);
nand U8491 (N_8491,N_8378,N_8223);
or U8492 (N_8492,N_8309,N_8368);
and U8493 (N_8493,N_8163,N_8339);
xnor U8494 (N_8494,N_8304,N_8388);
nand U8495 (N_8495,N_8150,N_8289);
xnor U8496 (N_8496,N_8135,N_8130);
and U8497 (N_8497,N_8113,N_8370);
nor U8498 (N_8498,N_8320,N_8210);
nand U8499 (N_8499,N_8166,N_8259);
xor U8500 (N_8500,N_8101,N_8207);
nand U8501 (N_8501,N_8174,N_8105);
nand U8502 (N_8502,N_8318,N_8107);
xor U8503 (N_8503,N_8371,N_8364);
nand U8504 (N_8504,N_8201,N_8385);
or U8505 (N_8505,N_8346,N_8112);
or U8506 (N_8506,N_8256,N_8263);
xor U8507 (N_8507,N_8285,N_8269);
and U8508 (N_8508,N_8386,N_8317);
or U8509 (N_8509,N_8200,N_8190);
nor U8510 (N_8510,N_8249,N_8298);
and U8511 (N_8511,N_8391,N_8133);
nand U8512 (N_8512,N_8242,N_8246);
or U8513 (N_8513,N_8390,N_8220);
xor U8514 (N_8514,N_8374,N_8349);
or U8515 (N_8515,N_8352,N_8359);
or U8516 (N_8516,N_8276,N_8244);
nand U8517 (N_8517,N_8305,N_8142);
or U8518 (N_8518,N_8229,N_8231);
nand U8519 (N_8519,N_8384,N_8344);
or U8520 (N_8520,N_8120,N_8224);
nand U8521 (N_8521,N_8270,N_8169);
xnor U8522 (N_8522,N_8227,N_8355);
xnor U8523 (N_8523,N_8335,N_8217);
or U8524 (N_8524,N_8171,N_8162);
xor U8525 (N_8525,N_8373,N_8257);
or U8526 (N_8526,N_8251,N_8338);
xnor U8527 (N_8527,N_8282,N_8181);
xor U8528 (N_8528,N_8369,N_8141);
xnor U8529 (N_8529,N_8194,N_8306);
or U8530 (N_8530,N_8354,N_8240);
xnor U8531 (N_8531,N_8165,N_8376);
and U8532 (N_8532,N_8274,N_8337);
or U8533 (N_8533,N_8275,N_8284);
or U8534 (N_8534,N_8138,N_8250);
nand U8535 (N_8535,N_8334,N_8397);
nand U8536 (N_8536,N_8381,N_8292);
xnor U8537 (N_8537,N_8315,N_8399);
nor U8538 (N_8538,N_8127,N_8209);
and U8539 (N_8539,N_8146,N_8360);
or U8540 (N_8540,N_8211,N_8398);
xnor U8541 (N_8541,N_8383,N_8361);
nand U8542 (N_8542,N_8187,N_8294);
and U8543 (N_8543,N_8367,N_8271);
xor U8544 (N_8544,N_8247,N_8153);
or U8545 (N_8545,N_8154,N_8198);
or U8546 (N_8546,N_8192,N_8161);
xnor U8547 (N_8547,N_8267,N_8324);
xor U8548 (N_8548,N_8254,N_8295);
xnor U8549 (N_8549,N_8321,N_8147);
or U8550 (N_8550,N_8380,N_8210);
nand U8551 (N_8551,N_8293,N_8109);
and U8552 (N_8552,N_8357,N_8378);
nor U8553 (N_8553,N_8299,N_8217);
nand U8554 (N_8554,N_8384,N_8341);
or U8555 (N_8555,N_8239,N_8153);
nor U8556 (N_8556,N_8298,N_8384);
nand U8557 (N_8557,N_8136,N_8385);
xnor U8558 (N_8558,N_8314,N_8138);
nand U8559 (N_8559,N_8327,N_8311);
nand U8560 (N_8560,N_8118,N_8379);
nor U8561 (N_8561,N_8300,N_8299);
xnor U8562 (N_8562,N_8115,N_8364);
and U8563 (N_8563,N_8172,N_8227);
or U8564 (N_8564,N_8141,N_8105);
nor U8565 (N_8565,N_8165,N_8367);
xnor U8566 (N_8566,N_8375,N_8177);
and U8567 (N_8567,N_8315,N_8212);
xnor U8568 (N_8568,N_8240,N_8139);
or U8569 (N_8569,N_8108,N_8240);
nand U8570 (N_8570,N_8307,N_8369);
nor U8571 (N_8571,N_8137,N_8243);
nand U8572 (N_8572,N_8341,N_8250);
nand U8573 (N_8573,N_8180,N_8371);
and U8574 (N_8574,N_8315,N_8373);
xnor U8575 (N_8575,N_8174,N_8334);
xnor U8576 (N_8576,N_8335,N_8198);
xnor U8577 (N_8577,N_8123,N_8200);
or U8578 (N_8578,N_8128,N_8166);
xnor U8579 (N_8579,N_8340,N_8110);
nand U8580 (N_8580,N_8214,N_8156);
xor U8581 (N_8581,N_8370,N_8309);
and U8582 (N_8582,N_8352,N_8331);
xnor U8583 (N_8583,N_8382,N_8114);
nand U8584 (N_8584,N_8135,N_8163);
or U8585 (N_8585,N_8244,N_8326);
and U8586 (N_8586,N_8153,N_8388);
nand U8587 (N_8587,N_8183,N_8226);
or U8588 (N_8588,N_8377,N_8338);
nand U8589 (N_8589,N_8338,N_8237);
xnor U8590 (N_8590,N_8329,N_8271);
nor U8591 (N_8591,N_8261,N_8166);
or U8592 (N_8592,N_8382,N_8266);
and U8593 (N_8593,N_8195,N_8380);
nand U8594 (N_8594,N_8367,N_8377);
and U8595 (N_8595,N_8294,N_8188);
nand U8596 (N_8596,N_8201,N_8311);
and U8597 (N_8597,N_8111,N_8267);
xor U8598 (N_8598,N_8285,N_8327);
nand U8599 (N_8599,N_8391,N_8205);
nand U8600 (N_8600,N_8352,N_8138);
and U8601 (N_8601,N_8385,N_8127);
and U8602 (N_8602,N_8293,N_8313);
or U8603 (N_8603,N_8223,N_8193);
xor U8604 (N_8604,N_8280,N_8368);
xnor U8605 (N_8605,N_8378,N_8213);
and U8606 (N_8606,N_8109,N_8341);
and U8607 (N_8607,N_8229,N_8328);
nand U8608 (N_8608,N_8141,N_8261);
nor U8609 (N_8609,N_8172,N_8144);
nor U8610 (N_8610,N_8112,N_8282);
nand U8611 (N_8611,N_8272,N_8291);
and U8612 (N_8612,N_8269,N_8287);
and U8613 (N_8613,N_8360,N_8155);
and U8614 (N_8614,N_8257,N_8170);
nor U8615 (N_8615,N_8107,N_8140);
xnor U8616 (N_8616,N_8291,N_8237);
or U8617 (N_8617,N_8377,N_8393);
nor U8618 (N_8618,N_8336,N_8176);
nor U8619 (N_8619,N_8206,N_8253);
nand U8620 (N_8620,N_8127,N_8344);
or U8621 (N_8621,N_8342,N_8319);
and U8622 (N_8622,N_8189,N_8225);
and U8623 (N_8623,N_8252,N_8276);
or U8624 (N_8624,N_8308,N_8388);
nand U8625 (N_8625,N_8143,N_8180);
and U8626 (N_8626,N_8378,N_8292);
nand U8627 (N_8627,N_8356,N_8302);
or U8628 (N_8628,N_8288,N_8345);
xor U8629 (N_8629,N_8151,N_8264);
xor U8630 (N_8630,N_8345,N_8376);
or U8631 (N_8631,N_8221,N_8280);
nor U8632 (N_8632,N_8138,N_8310);
nand U8633 (N_8633,N_8308,N_8175);
nor U8634 (N_8634,N_8169,N_8218);
nor U8635 (N_8635,N_8273,N_8204);
xnor U8636 (N_8636,N_8324,N_8109);
nor U8637 (N_8637,N_8122,N_8299);
and U8638 (N_8638,N_8381,N_8256);
xnor U8639 (N_8639,N_8136,N_8252);
xnor U8640 (N_8640,N_8323,N_8276);
xnor U8641 (N_8641,N_8182,N_8376);
nor U8642 (N_8642,N_8108,N_8241);
nand U8643 (N_8643,N_8377,N_8335);
nand U8644 (N_8644,N_8261,N_8107);
xnor U8645 (N_8645,N_8303,N_8179);
nand U8646 (N_8646,N_8253,N_8227);
or U8647 (N_8647,N_8277,N_8172);
and U8648 (N_8648,N_8260,N_8151);
nand U8649 (N_8649,N_8149,N_8263);
or U8650 (N_8650,N_8237,N_8199);
xor U8651 (N_8651,N_8345,N_8340);
xnor U8652 (N_8652,N_8316,N_8202);
or U8653 (N_8653,N_8375,N_8104);
nor U8654 (N_8654,N_8346,N_8177);
or U8655 (N_8655,N_8256,N_8157);
nand U8656 (N_8656,N_8247,N_8182);
or U8657 (N_8657,N_8349,N_8394);
nand U8658 (N_8658,N_8330,N_8319);
and U8659 (N_8659,N_8176,N_8385);
xor U8660 (N_8660,N_8168,N_8254);
or U8661 (N_8661,N_8289,N_8271);
xnor U8662 (N_8662,N_8357,N_8245);
xor U8663 (N_8663,N_8325,N_8231);
or U8664 (N_8664,N_8181,N_8375);
and U8665 (N_8665,N_8158,N_8186);
xnor U8666 (N_8666,N_8194,N_8256);
nor U8667 (N_8667,N_8396,N_8295);
or U8668 (N_8668,N_8121,N_8103);
or U8669 (N_8669,N_8304,N_8383);
xnor U8670 (N_8670,N_8238,N_8169);
xnor U8671 (N_8671,N_8297,N_8243);
nor U8672 (N_8672,N_8313,N_8105);
nor U8673 (N_8673,N_8377,N_8178);
xor U8674 (N_8674,N_8249,N_8193);
nand U8675 (N_8675,N_8148,N_8339);
and U8676 (N_8676,N_8378,N_8317);
or U8677 (N_8677,N_8247,N_8127);
nor U8678 (N_8678,N_8268,N_8208);
xor U8679 (N_8679,N_8235,N_8371);
xnor U8680 (N_8680,N_8336,N_8214);
xor U8681 (N_8681,N_8175,N_8328);
nand U8682 (N_8682,N_8352,N_8291);
nor U8683 (N_8683,N_8316,N_8221);
xor U8684 (N_8684,N_8239,N_8150);
and U8685 (N_8685,N_8343,N_8245);
nor U8686 (N_8686,N_8103,N_8185);
or U8687 (N_8687,N_8129,N_8336);
and U8688 (N_8688,N_8314,N_8299);
or U8689 (N_8689,N_8261,N_8237);
and U8690 (N_8690,N_8145,N_8218);
or U8691 (N_8691,N_8311,N_8241);
and U8692 (N_8692,N_8192,N_8152);
xnor U8693 (N_8693,N_8329,N_8144);
xnor U8694 (N_8694,N_8387,N_8299);
and U8695 (N_8695,N_8286,N_8304);
or U8696 (N_8696,N_8235,N_8115);
or U8697 (N_8697,N_8112,N_8358);
nand U8698 (N_8698,N_8275,N_8348);
and U8699 (N_8699,N_8138,N_8129);
or U8700 (N_8700,N_8476,N_8606);
xor U8701 (N_8701,N_8561,N_8468);
nand U8702 (N_8702,N_8590,N_8671);
or U8703 (N_8703,N_8428,N_8513);
and U8704 (N_8704,N_8609,N_8638);
xnor U8705 (N_8705,N_8453,N_8510);
and U8706 (N_8706,N_8534,N_8615);
nor U8707 (N_8707,N_8568,N_8680);
nor U8708 (N_8708,N_8425,N_8450);
nand U8709 (N_8709,N_8578,N_8552);
or U8710 (N_8710,N_8665,N_8575);
or U8711 (N_8711,N_8417,N_8454);
nand U8712 (N_8712,N_8579,N_8576);
nand U8713 (N_8713,N_8586,N_8692);
nand U8714 (N_8714,N_8600,N_8555);
or U8715 (N_8715,N_8505,N_8622);
and U8716 (N_8716,N_8408,N_8518);
nor U8717 (N_8717,N_8444,N_8461);
xnor U8718 (N_8718,N_8628,N_8439);
nand U8719 (N_8719,N_8509,N_8677);
nand U8720 (N_8720,N_8598,N_8535);
nor U8721 (N_8721,N_8695,N_8456);
nand U8722 (N_8722,N_8673,N_8502);
or U8723 (N_8723,N_8459,N_8608);
or U8724 (N_8724,N_8511,N_8607);
nor U8725 (N_8725,N_8506,N_8487);
xor U8726 (N_8726,N_8637,N_8532);
nand U8727 (N_8727,N_8482,N_8524);
xnor U8728 (N_8728,N_8494,N_8619);
nand U8729 (N_8729,N_8406,N_8694);
nor U8730 (N_8730,N_8413,N_8441);
nor U8731 (N_8731,N_8641,N_8658);
nand U8732 (N_8732,N_8642,N_8650);
and U8733 (N_8733,N_8675,N_8593);
and U8734 (N_8734,N_8520,N_8530);
nand U8735 (N_8735,N_8596,N_8523);
and U8736 (N_8736,N_8447,N_8556);
or U8737 (N_8737,N_8499,N_8451);
nor U8738 (N_8738,N_8554,N_8624);
xnor U8739 (N_8739,N_8445,N_8491);
and U8740 (N_8740,N_8632,N_8653);
xnor U8741 (N_8741,N_8438,N_8660);
nor U8742 (N_8742,N_8630,N_8527);
xnor U8743 (N_8743,N_8640,N_8611);
and U8744 (N_8744,N_8681,N_8538);
nor U8745 (N_8745,N_8462,N_8631);
and U8746 (N_8746,N_8643,N_8669);
and U8747 (N_8747,N_8446,N_8626);
xnor U8748 (N_8748,N_8486,N_8644);
or U8749 (N_8749,N_8404,N_8411);
nand U8750 (N_8750,N_8551,N_8496);
nor U8751 (N_8751,N_8465,N_8560);
and U8752 (N_8752,N_8466,N_8563);
and U8753 (N_8753,N_8407,N_8566);
nor U8754 (N_8754,N_8687,N_8541);
or U8755 (N_8755,N_8443,N_8489);
and U8756 (N_8756,N_8549,N_8587);
nand U8757 (N_8757,N_8449,N_8431);
xnor U8758 (N_8758,N_8668,N_8503);
nor U8759 (N_8759,N_8580,N_8432);
nand U8760 (N_8760,N_8659,N_8592);
nor U8761 (N_8761,N_8636,N_8672);
or U8762 (N_8762,N_8436,N_8647);
or U8763 (N_8763,N_8562,N_8455);
and U8764 (N_8764,N_8661,N_8690);
nand U8765 (N_8765,N_8625,N_8648);
xor U8766 (N_8766,N_8564,N_8495);
nor U8767 (N_8767,N_8683,N_8540);
nor U8768 (N_8768,N_8612,N_8684);
nor U8769 (N_8769,N_8400,N_8514);
or U8770 (N_8770,N_8557,N_8480);
or U8771 (N_8771,N_8616,N_8458);
xor U8772 (N_8772,N_8492,N_8594);
or U8773 (N_8773,N_8548,N_8602);
or U8774 (N_8774,N_8691,N_8457);
nand U8775 (N_8775,N_8686,N_8610);
nor U8776 (N_8776,N_8674,N_8553);
nand U8777 (N_8777,N_8565,N_8663);
xor U8778 (N_8778,N_8547,N_8485);
and U8779 (N_8779,N_8473,N_8437);
nor U8780 (N_8780,N_8679,N_8639);
nor U8781 (N_8781,N_8655,N_8629);
xnor U8782 (N_8782,N_8605,N_8403);
and U8783 (N_8783,N_8414,N_8559);
xor U8784 (N_8784,N_8651,N_8662);
nand U8785 (N_8785,N_8401,N_8652);
nand U8786 (N_8786,N_8550,N_8490);
nor U8787 (N_8787,N_8529,N_8519);
nand U8788 (N_8788,N_8424,N_8604);
or U8789 (N_8789,N_8645,N_8500);
nor U8790 (N_8790,N_8498,N_8617);
or U8791 (N_8791,N_8682,N_8621);
and U8792 (N_8792,N_8464,N_8533);
and U8793 (N_8793,N_8526,N_8528);
and U8794 (N_8794,N_8430,N_8670);
nor U8795 (N_8795,N_8516,N_8531);
or U8796 (N_8796,N_8574,N_8649);
or U8797 (N_8797,N_8484,N_8440);
nor U8798 (N_8798,N_8603,N_8422);
xor U8799 (N_8799,N_8423,N_8688);
xnor U8800 (N_8800,N_8463,N_8442);
and U8801 (N_8801,N_8597,N_8483);
and U8802 (N_8802,N_8589,N_8601);
nand U8803 (N_8803,N_8536,N_8478);
and U8804 (N_8804,N_8623,N_8409);
xnor U8805 (N_8805,N_8699,N_8501);
nand U8806 (N_8806,N_8572,N_8525);
or U8807 (N_8807,N_8472,N_8543);
and U8808 (N_8808,N_8433,N_8588);
or U8809 (N_8809,N_8507,N_8577);
or U8810 (N_8810,N_8664,N_8689);
and U8811 (N_8811,N_8435,N_8676);
nand U8812 (N_8812,N_8479,N_8656);
xnor U8813 (N_8813,N_8635,N_8429);
or U8814 (N_8814,N_8678,N_8558);
nand U8815 (N_8815,N_8488,N_8416);
nor U8816 (N_8816,N_8595,N_8493);
nand U8817 (N_8817,N_8504,N_8481);
xor U8818 (N_8818,N_8497,N_8567);
nand U8819 (N_8819,N_8410,N_8581);
xor U8820 (N_8820,N_8508,N_8569);
nor U8821 (N_8821,N_8545,N_8522);
nand U8822 (N_8822,N_8646,N_8469);
or U8823 (N_8823,N_8415,N_8448);
nor U8824 (N_8824,N_8697,N_8539);
and U8825 (N_8825,N_8418,N_8427);
nor U8826 (N_8826,N_8618,N_8614);
and U8827 (N_8827,N_8421,N_8471);
and U8828 (N_8828,N_8667,N_8420);
nor U8829 (N_8829,N_8657,N_8515);
or U8830 (N_8830,N_8573,N_8419);
and U8831 (N_8831,N_8585,N_8537);
xor U8832 (N_8832,N_8627,N_8544);
xor U8833 (N_8833,N_8434,N_8460);
nand U8834 (N_8834,N_8467,N_8666);
xor U8835 (N_8835,N_8685,N_8542);
nand U8836 (N_8836,N_8583,N_8412);
and U8837 (N_8837,N_8452,N_8477);
nand U8838 (N_8838,N_8512,N_8654);
xor U8839 (N_8839,N_8426,N_8582);
xnor U8840 (N_8840,N_8521,N_8613);
nor U8841 (N_8841,N_8475,N_8474);
nand U8842 (N_8842,N_8620,N_8517);
xor U8843 (N_8843,N_8405,N_8570);
nor U8844 (N_8844,N_8571,N_8546);
or U8845 (N_8845,N_8591,N_8633);
or U8846 (N_8846,N_8599,N_8696);
or U8847 (N_8847,N_8584,N_8470);
xor U8848 (N_8848,N_8634,N_8693);
xnor U8849 (N_8849,N_8402,N_8698);
xnor U8850 (N_8850,N_8455,N_8668);
nor U8851 (N_8851,N_8460,N_8687);
and U8852 (N_8852,N_8620,N_8418);
nand U8853 (N_8853,N_8672,N_8563);
nand U8854 (N_8854,N_8602,N_8633);
and U8855 (N_8855,N_8557,N_8479);
or U8856 (N_8856,N_8432,N_8426);
or U8857 (N_8857,N_8646,N_8656);
xor U8858 (N_8858,N_8654,N_8474);
or U8859 (N_8859,N_8667,N_8424);
nor U8860 (N_8860,N_8665,N_8501);
and U8861 (N_8861,N_8468,N_8588);
nor U8862 (N_8862,N_8403,N_8469);
or U8863 (N_8863,N_8431,N_8630);
and U8864 (N_8864,N_8569,N_8491);
or U8865 (N_8865,N_8643,N_8689);
nand U8866 (N_8866,N_8445,N_8543);
nand U8867 (N_8867,N_8510,N_8692);
or U8868 (N_8868,N_8445,N_8681);
nand U8869 (N_8869,N_8659,N_8424);
and U8870 (N_8870,N_8560,N_8491);
or U8871 (N_8871,N_8599,N_8563);
nor U8872 (N_8872,N_8449,N_8475);
xor U8873 (N_8873,N_8668,N_8491);
or U8874 (N_8874,N_8521,N_8412);
nor U8875 (N_8875,N_8436,N_8619);
nor U8876 (N_8876,N_8477,N_8402);
nor U8877 (N_8877,N_8517,N_8456);
or U8878 (N_8878,N_8610,N_8588);
nor U8879 (N_8879,N_8417,N_8498);
and U8880 (N_8880,N_8484,N_8401);
and U8881 (N_8881,N_8660,N_8583);
xnor U8882 (N_8882,N_8498,N_8586);
or U8883 (N_8883,N_8559,N_8546);
and U8884 (N_8884,N_8413,N_8560);
nand U8885 (N_8885,N_8404,N_8609);
nor U8886 (N_8886,N_8535,N_8634);
and U8887 (N_8887,N_8464,N_8465);
nor U8888 (N_8888,N_8504,N_8581);
xnor U8889 (N_8889,N_8656,N_8604);
nand U8890 (N_8890,N_8503,N_8455);
or U8891 (N_8891,N_8543,N_8647);
nand U8892 (N_8892,N_8437,N_8563);
nor U8893 (N_8893,N_8626,N_8561);
or U8894 (N_8894,N_8609,N_8437);
nand U8895 (N_8895,N_8450,N_8557);
and U8896 (N_8896,N_8675,N_8418);
nand U8897 (N_8897,N_8520,N_8466);
nor U8898 (N_8898,N_8624,N_8466);
nor U8899 (N_8899,N_8474,N_8565);
nor U8900 (N_8900,N_8524,N_8694);
nor U8901 (N_8901,N_8679,N_8601);
or U8902 (N_8902,N_8407,N_8481);
nor U8903 (N_8903,N_8682,N_8649);
xor U8904 (N_8904,N_8583,N_8617);
and U8905 (N_8905,N_8511,N_8513);
xor U8906 (N_8906,N_8416,N_8644);
xnor U8907 (N_8907,N_8667,N_8684);
nand U8908 (N_8908,N_8572,N_8424);
nand U8909 (N_8909,N_8428,N_8470);
nor U8910 (N_8910,N_8548,N_8535);
or U8911 (N_8911,N_8422,N_8614);
xnor U8912 (N_8912,N_8506,N_8486);
nand U8913 (N_8913,N_8550,N_8499);
nor U8914 (N_8914,N_8435,N_8638);
nor U8915 (N_8915,N_8564,N_8488);
and U8916 (N_8916,N_8679,N_8429);
nand U8917 (N_8917,N_8535,N_8563);
nor U8918 (N_8918,N_8422,N_8639);
nand U8919 (N_8919,N_8670,N_8451);
or U8920 (N_8920,N_8622,N_8482);
or U8921 (N_8921,N_8526,N_8638);
xor U8922 (N_8922,N_8628,N_8642);
nand U8923 (N_8923,N_8412,N_8598);
and U8924 (N_8924,N_8435,N_8612);
or U8925 (N_8925,N_8482,N_8488);
xnor U8926 (N_8926,N_8401,N_8514);
nand U8927 (N_8927,N_8558,N_8416);
nand U8928 (N_8928,N_8671,N_8472);
nor U8929 (N_8929,N_8533,N_8549);
and U8930 (N_8930,N_8685,N_8503);
and U8931 (N_8931,N_8532,N_8404);
nor U8932 (N_8932,N_8443,N_8608);
nand U8933 (N_8933,N_8553,N_8471);
and U8934 (N_8934,N_8463,N_8620);
or U8935 (N_8935,N_8447,N_8545);
or U8936 (N_8936,N_8642,N_8472);
nand U8937 (N_8937,N_8514,N_8599);
or U8938 (N_8938,N_8656,N_8696);
or U8939 (N_8939,N_8510,N_8548);
xor U8940 (N_8940,N_8537,N_8682);
xor U8941 (N_8941,N_8519,N_8472);
and U8942 (N_8942,N_8611,N_8404);
or U8943 (N_8943,N_8546,N_8673);
and U8944 (N_8944,N_8527,N_8592);
nor U8945 (N_8945,N_8513,N_8624);
nand U8946 (N_8946,N_8690,N_8567);
and U8947 (N_8947,N_8428,N_8573);
and U8948 (N_8948,N_8444,N_8412);
nor U8949 (N_8949,N_8492,N_8419);
or U8950 (N_8950,N_8495,N_8599);
xnor U8951 (N_8951,N_8522,N_8686);
or U8952 (N_8952,N_8648,N_8453);
and U8953 (N_8953,N_8405,N_8425);
and U8954 (N_8954,N_8699,N_8585);
or U8955 (N_8955,N_8437,N_8501);
nor U8956 (N_8956,N_8449,N_8696);
xor U8957 (N_8957,N_8622,N_8547);
or U8958 (N_8958,N_8542,N_8526);
or U8959 (N_8959,N_8449,N_8447);
and U8960 (N_8960,N_8555,N_8448);
nand U8961 (N_8961,N_8650,N_8597);
nand U8962 (N_8962,N_8512,N_8552);
xnor U8963 (N_8963,N_8465,N_8574);
nand U8964 (N_8964,N_8551,N_8617);
nand U8965 (N_8965,N_8495,N_8540);
xnor U8966 (N_8966,N_8579,N_8656);
xor U8967 (N_8967,N_8432,N_8654);
nand U8968 (N_8968,N_8470,N_8402);
nand U8969 (N_8969,N_8563,N_8518);
nand U8970 (N_8970,N_8503,N_8551);
xor U8971 (N_8971,N_8439,N_8572);
or U8972 (N_8972,N_8513,N_8594);
nor U8973 (N_8973,N_8440,N_8600);
and U8974 (N_8974,N_8533,N_8445);
nand U8975 (N_8975,N_8425,N_8441);
xnor U8976 (N_8976,N_8402,N_8579);
or U8977 (N_8977,N_8403,N_8548);
nor U8978 (N_8978,N_8544,N_8591);
nor U8979 (N_8979,N_8498,N_8624);
or U8980 (N_8980,N_8656,N_8466);
xor U8981 (N_8981,N_8677,N_8410);
and U8982 (N_8982,N_8433,N_8537);
xor U8983 (N_8983,N_8640,N_8531);
nand U8984 (N_8984,N_8577,N_8575);
nor U8985 (N_8985,N_8671,N_8672);
and U8986 (N_8986,N_8653,N_8423);
or U8987 (N_8987,N_8587,N_8480);
and U8988 (N_8988,N_8644,N_8509);
or U8989 (N_8989,N_8464,N_8690);
nand U8990 (N_8990,N_8496,N_8680);
or U8991 (N_8991,N_8628,N_8577);
and U8992 (N_8992,N_8543,N_8571);
xnor U8993 (N_8993,N_8571,N_8455);
and U8994 (N_8994,N_8618,N_8481);
nor U8995 (N_8995,N_8651,N_8456);
xnor U8996 (N_8996,N_8550,N_8503);
nand U8997 (N_8997,N_8561,N_8693);
nor U8998 (N_8998,N_8695,N_8554);
or U8999 (N_8999,N_8567,N_8694);
xor U9000 (N_9000,N_8704,N_8726);
or U9001 (N_9001,N_8920,N_8885);
and U9002 (N_9002,N_8977,N_8746);
nor U9003 (N_9003,N_8931,N_8916);
and U9004 (N_9004,N_8995,N_8768);
xor U9005 (N_9005,N_8883,N_8976);
or U9006 (N_9006,N_8766,N_8993);
and U9007 (N_9007,N_8892,N_8829);
or U9008 (N_9008,N_8838,N_8730);
nand U9009 (N_9009,N_8859,N_8922);
xnor U9010 (N_9010,N_8813,N_8868);
nor U9011 (N_9011,N_8918,N_8964);
xor U9012 (N_9012,N_8744,N_8914);
or U9013 (N_9013,N_8850,N_8933);
nor U9014 (N_9014,N_8751,N_8783);
nor U9015 (N_9015,N_8937,N_8871);
and U9016 (N_9016,N_8737,N_8717);
or U9017 (N_9017,N_8724,N_8950);
xnor U9018 (N_9018,N_8946,N_8849);
nor U9019 (N_9019,N_8764,N_8841);
and U9020 (N_9020,N_8945,N_8845);
nor U9021 (N_9021,N_8742,N_8955);
and U9022 (N_9022,N_8784,N_8994);
xor U9023 (N_9023,N_8728,N_8992);
and U9024 (N_9024,N_8723,N_8959);
nand U9025 (N_9025,N_8798,N_8894);
nor U9026 (N_9026,N_8858,N_8747);
or U9027 (N_9027,N_8967,N_8758);
or U9028 (N_9028,N_8991,N_8881);
xnor U9029 (N_9029,N_8924,N_8949);
or U9030 (N_9030,N_8794,N_8939);
nor U9031 (N_9031,N_8759,N_8736);
or U9032 (N_9032,N_8823,N_8824);
xnor U9033 (N_9033,N_8806,N_8770);
and U9034 (N_9034,N_8917,N_8815);
nand U9035 (N_9035,N_8767,N_8782);
or U9036 (N_9036,N_8827,N_8769);
nor U9037 (N_9037,N_8734,N_8743);
xnor U9038 (N_9038,N_8873,N_8983);
nor U9039 (N_9039,N_8909,N_8864);
xnor U9040 (N_9040,N_8752,N_8989);
nor U9041 (N_9041,N_8904,N_8905);
nand U9042 (N_9042,N_8803,N_8943);
xor U9043 (N_9043,N_8971,N_8855);
or U9044 (N_9044,N_8880,N_8779);
xnor U9045 (N_9045,N_8848,N_8710);
nand U9046 (N_9046,N_8760,N_8851);
xnor U9047 (N_9047,N_8715,N_8739);
xnor U9048 (N_9048,N_8804,N_8825);
xor U9049 (N_9049,N_8707,N_8941);
or U9050 (N_9050,N_8853,N_8898);
xor U9051 (N_9051,N_8781,N_8966);
nor U9052 (N_9052,N_8954,N_8750);
nand U9053 (N_9053,N_8897,N_8833);
xnor U9054 (N_9054,N_8785,N_8812);
and U9055 (N_9055,N_8846,N_8874);
xnor U9056 (N_9056,N_8722,N_8990);
and U9057 (N_9057,N_8729,N_8840);
nand U9058 (N_9058,N_8862,N_8842);
and U9059 (N_9059,N_8800,N_8965);
xnor U9060 (N_9060,N_8786,N_8709);
xor U9061 (N_9061,N_8708,N_8795);
and U9062 (N_9062,N_8807,N_8997);
and U9063 (N_9063,N_8811,N_8884);
nor U9064 (N_9064,N_8765,N_8944);
nand U9065 (N_9065,N_8814,N_8738);
nor U9066 (N_9066,N_8876,N_8835);
nor U9067 (N_9067,N_8700,N_8857);
nor U9068 (N_9068,N_8951,N_8915);
or U9069 (N_9069,N_8836,N_8731);
xnor U9070 (N_9070,N_8908,N_8843);
nor U9071 (N_9071,N_8969,N_8972);
nand U9072 (N_9072,N_8961,N_8889);
and U9073 (N_9073,N_8773,N_8932);
or U9074 (N_9074,N_8928,N_8952);
or U9075 (N_9075,N_8839,N_8978);
or U9076 (N_9076,N_8973,N_8819);
nand U9077 (N_9077,N_8808,N_8870);
nand U9078 (N_9078,N_8847,N_8832);
nand U9079 (N_9079,N_8740,N_8778);
nor U9080 (N_9080,N_8895,N_8878);
nor U9081 (N_9081,N_8720,N_8763);
or U9082 (N_9082,N_8882,N_8791);
and U9083 (N_9083,N_8777,N_8822);
and U9084 (N_9084,N_8820,N_8877);
nor U9085 (N_9085,N_8856,N_8810);
nor U9086 (N_9086,N_8926,N_8867);
xnor U9087 (N_9087,N_8741,N_8711);
nor U9088 (N_9088,N_8831,N_8818);
or U9089 (N_9089,N_8716,N_8788);
and U9090 (N_9090,N_8893,N_8844);
or U9091 (N_9091,N_8996,N_8748);
nand U9092 (N_9092,N_8809,N_8887);
and U9093 (N_9093,N_8907,N_8956);
or U9094 (N_9094,N_8953,N_8930);
xnor U9095 (N_9095,N_8725,N_8960);
nor U9096 (N_9096,N_8934,N_8987);
xnor U9097 (N_9097,N_8910,N_8968);
and U9098 (N_9098,N_8714,N_8753);
nor U9099 (N_9099,N_8834,N_8912);
nand U9100 (N_9100,N_8828,N_8985);
nand U9101 (N_9101,N_8702,N_8963);
xor U9102 (N_9102,N_8911,N_8757);
nor U9103 (N_9103,N_8745,N_8797);
nor U9104 (N_9104,N_8982,N_8821);
xnor U9105 (N_9105,N_8923,N_8927);
and U9106 (N_9106,N_8888,N_8900);
xnor U9107 (N_9107,N_8817,N_8761);
or U9108 (N_9108,N_8942,N_8805);
nand U9109 (N_9109,N_8886,N_8792);
xor U9110 (N_9110,N_8999,N_8925);
nand U9111 (N_9111,N_8863,N_8756);
xnor U9112 (N_9112,N_8865,N_8875);
xnor U9113 (N_9113,N_8790,N_8718);
xnor U9114 (N_9114,N_8869,N_8854);
and U9115 (N_9115,N_8913,N_8860);
nor U9116 (N_9116,N_8891,N_8787);
xnor U9117 (N_9117,N_8776,N_8735);
or U9118 (N_9118,N_8935,N_8719);
or U9119 (N_9119,N_8852,N_8830);
nand U9120 (N_9120,N_8799,N_8879);
and U9121 (N_9121,N_8984,N_8774);
and U9122 (N_9122,N_8921,N_8929);
or U9123 (N_9123,N_8762,N_8902);
and U9124 (N_9124,N_8980,N_8772);
nor U9125 (N_9125,N_8936,N_8789);
nor U9126 (N_9126,N_8796,N_8919);
and U9127 (N_9127,N_8974,N_8962);
nor U9128 (N_9128,N_8801,N_8940);
or U9129 (N_9129,N_8749,N_8988);
nor U9130 (N_9130,N_8975,N_8947);
or U9131 (N_9131,N_8816,N_8701);
xnor U9132 (N_9132,N_8826,N_8938);
nand U9133 (N_9133,N_8780,N_8802);
nor U9134 (N_9134,N_8721,N_8866);
xnor U9135 (N_9135,N_8837,N_8901);
nand U9136 (N_9136,N_8906,N_8981);
nand U9137 (N_9137,N_8899,N_8998);
and U9138 (N_9138,N_8771,N_8713);
nand U9139 (N_9139,N_8705,N_8727);
and U9140 (N_9140,N_8754,N_8703);
nor U9141 (N_9141,N_8872,N_8732);
and U9142 (N_9142,N_8793,N_8896);
xnor U9143 (N_9143,N_8775,N_8903);
and U9144 (N_9144,N_8957,N_8890);
nand U9145 (N_9145,N_8986,N_8706);
xor U9146 (N_9146,N_8970,N_8979);
nor U9147 (N_9147,N_8712,N_8755);
and U9148 (N_9148,N_8958,N_8948);
and U9149 (N_9149,N_8733,N_8861);
nand U9150 (N_9150,N_8828,N_8873);
or U9151 (N_9151,N_8833,N_8969);
and U9152 (N_9152,N_8833,N_8944);
nor U9153 (N_9153,N_8970,N_8775);
nor U9154 (N_9154,N_8797,N_8997);
nor U9155 (N_9155,N_8791,N_8930);
xor U9156 (N_9156,N_8874,N_8908);
xor U9157 (N_9157,N_8975,N_8888);
or U9158 (N_9158,N_8778,N_8795);
or U9159 (N_9159,N_8775,N_8703);
or U9160 (N_9160,N_8848,N_8825);
nand U9161 (N_9161,N_8719,N_8750);
or U9162 (N_9162,N_8991,N_8949);
and U9163 (N_9163,N_8848,N_8918);
nand U9164 (N_9164,N_8891,N_8809);
xor U9165 (N_9165,N_8800,N_8803);
xor U9166 (N_9166,N_8874,N_8917);
or U9167 (N_9167,N_8886,N_8952);
or U9168 (N_9168,N_8890,N_8941);
xnor U9169 (N_9169,N_8964,N_8815);
xnor U9170 (N_9170,N_8933,N_8833);
nand U9171 (N_9171,N_8759,N_8815);
nor U9172 (N_9172,N_8951,N_8953);
nand U9173 (N_9173,N_8850,N_8982);
nor U9174 (N_9174,N_8961,N_8816);
and U9175 (N_9175,N_8792,N_8852);
xor U9176 (N_9176,N_8786,N_8730);
nor U9177 (N_9177,N_8878,N_8943);
and U9178 (N_9178,N_8749,N_8913);
nor U9179 (N_9179,N_8779,N_8776);
or U9180 (N_9180,N_8884,N_8967);
or U9181 (N_9181,N_8916,N_8853);
xor U9182 (N_9182,N_8808,N_8937);
nand U9183 (N_9183,N_8905,N_8911);
nand U9184 (N_9184,N_8947,N_8765);
nand U9185 (N_9185,N_8759,N_8976);
or U9186 (N_9186,N_8829,N_8768);
nand U9187 (N_9187,N_8975,N_8949);
or U9188 (N_9188,N_8874,N_8725);
nand U9189 (N_9189,N_8991,N_8785);
nand U9190 (N_9190,N_8997,N_8979);
nor U9191 (N_9191,N_8798,N_8837);
nand U9192 (N_9192,N_8768,N_8910);
or U9193 (N_9193,N_8964,N_8946);
xnor U9194 (N_9194,N_8759,N_8732);
or U9195 (N_9195,N_8971,N_8958);
xnor U9196 (N_9196,N_8700,N_8786);
nand U9197 (N_9197,N_8858,N_8806);
nand U9198 (N_9198,N_8871,N_8726);
xor U9199 (N_9199,N_8764,N_8757);
or U9200 (N_9200,N_8920,N_8918);
nand U9201 (N_9201,N_8704,N_8741);
or U9202 (N_9202,N_8829,N_8996);
xnor U9203 (N_9203,N_8878,N_8778);
or U9204 (N_9204,N_8850,N_8911);
or U9205 (N_9205,N_8888,N_8913);
and U9206 (N_9206,N_8758,N_8875);
nor U9207 (N_9207,N_8870,N_8716);
or U9208 (N_9208,N_8897,N_8987);
nor U9209 (N_9209,N_8999,N_8875);
nor U9210 (N_9210,N_8898,N_8919);
xor U9211 (N_9211,N_8814,N_8764);
xor U9212 (N_9212,N_8984,N_8857);
and U9213 (N_9213,N_8981,N_8874);
or U9214 (N_9214,N_8786,N_8986);
or U9215 (N_9215,N_8964,N_8973);
and U9216 (N_9216,N_8923,N_8852);
or U9217 (N_9217,N_8935,N_8793);
nand U9218 (N_9218,N_8931,N_8917);
nor U9219 (N_9219,N_8912,N_8726);
xor U9220 (N_9220,N_8872,N_8997);
xor U9221 (N_9221,N_8843,N_8784);
nor U9222 (N_9222,N_8852,N_8979);
xor U9223 (N_9223,N_8848,N_8851);
xnor U9224 (N_9224,N_8831,N_8819);
or U9225 (N_9225,N_8761,N_8990);
nor U9226 (N_9226,N_8826,N_8806);
and U9227 (N_9227,N_8815,N_8723);
or U9228 (N_9228,N_8810,N_8910);
xor U9229 (N_9229,N_8979,N_8985);
nand U9230 (N_9230,N_8986,N_8771);
nand U9231 (N_9231,N_8888,N_8934);
xnor U9232 (N_9232,N_8792,N_8982);
nand U9233 (N_9233,N_8725,N_8703);
nor U9234 (N_9234,N_8772,N_8792);
or U9235 (N_9235,N_8776,N_8901);
and U9236 (N_9236,N_8841,N_8944);
xor U9237 (N_9237,N_8823,N_8783);
and U9238 (N_9238,N_8785,N_8819);
and U9239 (N_9239,N_8827,N_8765);
or U9240 (N_9240,N_8801,N_8921);
and U9241 (N_9241,N_8912,N_8707);
nor U9242 (N_9242,N_8812,N_8987);
nor U9243 (N_9243,N_8791,N_8724);
or U9244 (N_9244,N_8952,N_8890);
and U9245 (N_9245,N_8835,N_8780);
and U9246 (N_9246,N_8932,N_8976);
nand U9247 (N_9247,N_8768,N_8748);
and U9248 (N_9248,N_8975,N_8833);
and U9249 (N_9249,N_8902,N_8928);
and U9250 (N_9250,N_8703,N_8850);
nand U9251 (N_9251,N_8952,N_8865);
and U9252 (N_9252,N_8727,N_8955);
xnor U9253 (N_9253,N_8814,N_8895);
nor U9254 (N_9254,N_8747,N_8766);
and U9255 (N_9255,N_8896,N_8754);
and U9256 (N_9256,N_8798,N_8709);
or U9257 (N_9257,N_8874,N_8760);
or U9258 (N_9258,N_8764,N_8880);
and U9259 (N_9259,N_8950,N_8949);
nand U9260 (N_9260,N_8711,N_8894);
nor U9261 (N_9261,N_8895,N_8730);
and U9262 (N_9262,N_8799,N_8779);
nor U9263 (N_9263,N_8855,N_8743);
or U9264 (N_9264,N_8824,N_8808);
xnor U9265 (N_9265,N_8822,N_8812);
xor U9266 (N_9266,N_8796,N_8845);
xnor U9267 (N_9267,N_8861,N_8814);
nor U9268 (N_9268,N_8770,N_8918);
or U9269 (N_9269,N_8969,N_8826);
and U9270 (N_9270,N_8853,N_8959);
nand U9271 (N_9271,N_8816,N_8805);
nor U9272 (N_9272,N_8784,N_8765);
nor U9273 (N_9273,N_8796,N_8920);
and U9274 (N_9274,N_8926,N_8732);
or U9275 (N_9275,N_8708,N_8789);
or U9276 (N_9276,N_8847,N_8868);
or U9277 (N_9277,N_8995,N_8749);
xor U9278 (N_9278,N_8943,N_8831);
nor U9279 (N_9279,N_8782,N_8995);
and U9280 (N_9280,N_8877,N_8866);
xor U9281 (N_9281,N_8823,N_8829);
xnor U9282 (N_9282,N_8917,N_8992);
nor U9283 (N_9283,N_8895,N_8804);
xnor U9284 (N_9284,N_8945,N_8771);
or U9285 (N_9285,N_8951,N_8896);
nor U9286 (N_9286,N_8738,N_8848);
and U9287 (N_9287,N_8880,N_8855);
xor U9288 (N_9288,N_8788,N_8964);
nor U9289 (N_9289,N_8972,N_8892);
or U9290 (N_9290,N_8815,N_8991);
xor U9291 (N_9291,N_8877,N_8879);
nand U9292 (N_9292,N_8705,N_8832);
xnor U9293 (N_9293,N_8761,N_8701);
or U9294 (N_9294,N_8778,N_8955);
nor U9295 (N_9295,N_8825,N_8849);
xor U9296 (N_9296,N_8817,N_8801);
nor U9297 (N_9297,N_8908,N_8830);
nand U9298 (N_9298,N_8844,N_8743);
nand U9299 (N_9299,N_8840,N_8812);
nor U9300 (N_9300,N_9039,N_9083);
xor U9301 (N_9301,N_9085,N_9075);
xor U9302 (N_9302,N_9263,N_9213);
nand U9303 (N_9303,N_9052,N_9105);
xnor U9304 (N_9304,N_9049,N_9141);
nand U9305 (N_9305,N_9020,N_9080);
xor U9306 (N_9306,N_9060,N_9242);
xnor U9307 (N_9307,N_9026,N_9233);
nor U9308 (N_9308,N_9250,N_9008);
nor U9309 (N_9309,N_9293,N_9179);
nand U9310 (N_9310,N_9191,N_9063);
nor U9311 (N_9311,N_9119,N_9042);
xor U9312 (N_9312,N_9210,N_9097);
or U9313 (N_9313,N_9082,N_9134);
and U9314 (N_9314,N_9151,N_9106);
and U9315 (N_9315,N_9099,N_9072);
nor U9316 (N_9316,N_9056,N_9013);
and U9317 (N_9317,N_9071,N_9285);
nor U9318 (N_9318,N_9275,N_9068);
or U9319 (N_9319,N_9247,N_9167);
nand U9320 (N_9320,N_9261,N_9208);
nand U9321 (N_9321,N_9093,N_9248);
nand U9322 (N_9322,N_9053,N_9079);
nor U9323 (N_9323,N_9066,N_9268);
nor U9324 (N_9324,N_9028,N_9288);
xnor U9325 (N_9325,N_9044,N_9209);
xnor U9326 (N_9326,N_9012,N_9264);
nor U9327 (N_9327,N_9102,N_9211);
nand U9328 (N_9328,N_9112,N_9243);
and U9329 (N_9329,N_9098,N_9017);
or U9330 (N_9330,N_9237,N_9043);
xnor U9331 (N_9331,N_9036,N_9192);
xor U9332 (N_9332,N_9190,N_9168);
nor U9333 (N_9333,N_9050,N_9158);
and U9334 (N_9334,N_9100,N_9219);
or U9335 (N_9335,N_9061,N_9260);
xnor U9336 (N_9336,N_9280,N_9070);
and U9337 (N_9337,N_9120,N_9113);
and U9338 (N_9338,N_9265,N_9088);
and U9339 (N_9339,N_9062,N_9027);
nand U9340 (N_9340,N_9007,N_9220);
and U9341 (N_9341,N_9198,N_9270);
nor U9342 (N_9342,N_9069,N_9018);
nor U9343 (N_9343,N_9235,N_9057);
and U9344 (N_9344,N_9162,N_9189);
nand U9345 (N_9345,N_9253,N_9148);
xnor U9346 (N_9346,N_9108,N_9298);
nand U9347 (N_9347,N_9153,N_9023);
xnor U9348 (N_9348,N_9299,N_9204);
nor U9349 (N_9349,N_9033,N_9232);
nor U9350 (N_9350,N_9031,N_9259);
nand U9351 (N_9351,N_9199,N_9107);
nor U9352 (N_9352,N_9122,N_9188);
and U9353 (N_9353,N_9239,N_9174);
or U9354 (N_9354,N_9257,N_9234);
nor U9355 (N_9355,N_9011,N_9177);
nor U9356 (N_9356,N_9032,N_9161);
nor U9357 (N_9357,N_9284,N_9121);
or U9358 (N_9358,N_9126,N_9067);
xor U9359 (N_9359,N_9181,N_9022);
nand U9360 (N_9360,N_9025,N_9021);
nor U9361 (N_9361,N_9214,N_9130);
xor U9362 (N_9362,N_9095,N_9240);
and U9363 (N_9363,N_9159,N_9218);
or U9364 (N_9364,N_9110,N_9173);
and U9365 (N_9365,N_9142,N_9271);
and U9366 (N_9366,N_9176,N_9054);
xor U9367 (N_9367,N_9004,N_9255);
nor U9368 (N_9368,N_9078,N_9183);
or U9369 (N_9369,N_9166,N_9172);
and U9370 (N_9370,N_9203,N_9048);
or U9371 (N_9371,N_9076,N_9178);
nor U9372 (N_9372,N_9096,N_9230);
nor U9373 (N_9373,N_9212,N_9258);
nand U9374 (N_9374,N_9103,N_9144);
and U9375 (N_9375,N_9207,N_9147);
nand U9376 (N_9376,N_9086,N_9267);
xnor U9377 (N_9377,N_9014,N_9087);
or U9378 (N_9378,N_9241,N_9046);
and U9379 (N_9379,N_9055,N_9051);
xnor U9380 (N_9380,N_9274,N_9139);
nor U9381 (N_9381,N_9037,N_9077);
and U9382 (N_9382,N_9155,N_9279);
nor U9383 (N_9383,N_9281,N_9143);
xor U9384 (N_9384,N_9278,N_9266);
and U9385 (N_9385,N_9038,N_9254);
nor U9386 (N_9386,N_9015,N_9195);
or U9387 (N_9387,N_9296,N_9276);
nand U9388 (N_9388,N_9133,N_9217);
nand U9389 (N_9389,N_9249,N_9005);
nand U9390 (N_9390,N_9149,N_9127);
nor U9391 (N_9391,N_9157,N_9059);
nor U9392 (N_9392,N_9231,N_9129);
xnor U9393 (N_9393,N_9140,N_9283);
or U9394 (N_9394,N_9150,N_9227);
nand U9395 (N_9395,N_9128,N_9091);
nand U9396 (N_9396,N_9045,N_9273);
or U9397 (N_9397,N_9244,N_9200);
xnor U9398 (N_9398,N_9202,N_9184);
xnor U9399 (N_9399,N_9109,N_9058);
or U9400 (N_9400,N_9000,N_9197);
xor U9401 (N_9401,N_9165,N_9295);
and U9402 (N_9402,N_9201,N_9035);
nor U9403 (N_9403,N_9009,N_9297);
xor U9404 (N_9404,N_9215,N_9132);
nor U9405 (N_9405,N_9294,N_9065);
and U9406 (N_9406,N_9131,N_9002);
nor U9407 (N_9407,N_9136,N_9003);
nand U9408 (N_9408,N_9081,N_9084);
nor U9409 (N_9409,N_9251,N_9252);
or U9410 (N_9410,N_9029,N_9224);
xor U9411 (N_9411,N_9282,N_9163);
nand U9412 (N_9412,N_9030,N_9170);
and U9413 (N_9413,N_9146,N_9040);
xor U9414 (N_9414,N_9118,N_9269);
xor U9415 (N_9415,N_9006,N_9262);
and U9416 (N_9416,N_9101,N_9291);
nor U9417 (N_9417,N_9135,N_9138);
xnor U9418 (N_9418,N_9245,N_9137);
or U9419 (N_9419,N_9104,N_9175);
nor U9420 (N_9420,N_9236,N_9186);
or U9421 (N_9421,N_9123,N_9205);
nand U9422 (N_9422,N_9222,N_9193);
or U9423 (N_9423,N_9238,N_9125);
and U9424 (N_9424,N_9216,N_9287);
nor U9425 (N_9425,N_9010,N_9115);
nand U9426 (N_9426,N_9114,N_9111);
nor U9427 (N_9427,N_9092,N_9272);
nor U9428 (N_9428,N_9117,N_9182);
or U9429 (N_9429,N_9073,N_9019);
xnor U9430 (N_9430,N_9206,N_9180);
or U9431 (N_9431,N_9164,N_9256);
or U9432 (N_9432,N_9124,N_9185);
or U9433 (N_9433,N_9221,N_9156);
and U9434 (N_9434,N_9286,N_9171);
nand U9435 (N_9435,N_9154,N_9228);
xor U9436 (N_9436,N_9090,N_9187);
xor U9437 (N_9437,N_9277,N_9116);
xor U9438 (N_9438,N_9041,N_9290);
and U9439 (N_9439,N_9016,N_9089);
or U9440 (N_9440,N_9292,N_9145);
or U9441 (N_9441,N_9064,N_9047);
and U9442 (N_9442,N_9160,N_9024);
nor U9443 (N_9443,N_9223,N_9152);
xor U9444 (N_9444,N_9289,N_9229);
xor U9445 (N_9445,N_9169,N_9226);
nor U9446 (N_9446,N_9246,N_9194);
and U9447 (N_9447,N_9196,N_9225);
or U9448 (N_9448,N_9094,N_9001);
and U9449 (N_9449,N_9074,N_9034);
and U9450 (N_9450,N_9238,N_9056);
nor U9451 (N_9451,N_9079,N_9145);
or U9452 (N_9452,N_9281,N_9239);
nand U9453 (N_9453,N_9191,N_9020);
xor U9454 (N_9454,N_9055,N_9226);
and U9455 (N_9455,N_9165,N_9161);
nor U9456 (N_9456,N_9152,N_9298);
xnor U9457 (N_9457,N_9123,N_9129);
nor U9458 (N_9458,N_9081,N_9064);
or U9459 (N_9459,N_9129,N_9065);
xor U9460 (N_9460,N_9135,N_9070);
xnor U9461 (N_9461,N_9090,N_9231);
nor U9462 (N_9462,N_9247,N_9110);
nand U9463 (N_9463,N_9257,N_9147);
xor U9464 (N_9464,N_9282,N_9047);
nand U9465 (N_9465,N_9238,N_9004);
and U9466 (N_9466,N_9035,N_9246);
xnor U9467 (N_9467,N_9187,N_9139);
or U9468 (N_9468,N_9264,N_9167);
nand U9469 (N_9469,N_9102,N_9210);
xnor U9470 (N_9470,N_9252,N_9034);
or U9471 (N_9471,N_9000,N_9149);
xor U9472 (N_9472,N_9112,N_9037);
or U9473 (N_9473,N_9030,N_9038);
xnor U9474 (N_9474,N_9003,N_9154);
nor U9475 (N_9475,N_9020,N_9128);
xor U9476 (N_9476,N_9287,N_9094);
or U9477 (N_9477,N_9053,N_9251);
and U9478 (N_9478,N_9247,N_9034);
or U9479 (N_9479,N_9160,N_9167);
and U9480 (N_9480,N_9176,N_9228);
xnor U9481 (N_9481,N_9058,N_9196);
and U9482 (N_9482,N_9143,N_9116);
or U9483 (N_9483,N_9014,N_9281);
nand U9484 (N_9484,N_9299,N_9061);
nor U9485 (N_9485,N_9032,N_9001);
xor U9486 (N_9486,N_9063,N_9165);
xnor U9487 (N_9487,N_9154,N_9041);
nor U9488 (N_9488,N_9154,N_9282);
and U9489 (N_9489,N_9089,N_9292);
nand U9490 (N_9490,N_9217,N_9201);
nand U9491 (N_9491,N_9134,N_9146);
nor U9492 (N_9492,N_9131,N_9296);
and U9493 (N_9493,N_9222,N_9026);
or U9494 (N_9494,N_9113,N_9008);
nand U9495 (N_9495,N_9043,N_9161);
nor U9496 (N_9496,N_9209,N_9139);
or U9497 (N_9497,N_9113,N_9149);
nand U9498 (N_9498,N_9155,N_9112);
xnor U9499 (N_9499,N_9248,N_9069);
nand U9500 (N_9500,N_9068,N_9255);
or U9501 (N_9501,N_9233,N_9194);
xor U9502 (N_9502,N_9233,N_9144);
or U9503 (N_9503,N_9096,N_9009);
nor U9504 (N_9504,N_9293,N_9153);
and U9505 (N_9505,N_9042,N_9043);
xnor U9506 (N_9506,N_9019,N_9216);
nand U9507 (N_9507,N_9237,N_9271);
and U9508 (N_9508,N_9018,N_9015);
or U9509 (N_9509,N_9252,N_9102);
nand U9510 (N_9510,N_9037,N_9121);
nand U9511 (N_9511,N_9071,N_9225);
xnor U9512 (N_9512,N_9250,N_9041);
xor U9513 (N_9513,N_9243,N_9201);
xor U9514 (N_9514,N_9072,N_9180);
and U9515 (N_9515,N_9228,N_9286);
nand U9516 (N_9516,N_9267,N_9089);
or U9517 (N_9517,N_9167,N_9078);
or U9518 (N_9518,N_9036,N_9246);
nor U9519 (N_9519,N_9113,N_9153);
xnor U9520 (N_9520,N_9078,N_9267);
and U9521 (N_9521,N_9208,N_9274);
or U9522 (N_9522,N_9104,N_9129);
nand U9523 (N_9523,N_9208,N_9285);
nor U9524 (N_9524,N_9207,N_9274);
nand U9525 (N_9525,N_9273,N_9065);
xnor U9526 (N_9526,N_9169,N_9275);
nand U9527 (N_9527,N_9005,N_9018);
nor U9528 (N_9528,N_9082,N_9034);
or U9529 (N_9529,N_9219,N_9240);
nand U9530 (N_9530,N_9084,N_9184);
and U9531 (N_9531,N_9221,N_9004);
xor U9532 (N_9532,N_9110,N_9234);
nor U9533 (N_9533,N_9210,N_9159);
and U9534 (N_9534,N_9258,N_9269);
nor U9535 (N_9535,N_9249,N_9199);
xor U9536 (N_9536,N_9073,N_9040);
xor U9537 (N_9537,N_9178,N_9292);
nand U9538 (N_9538,N_9068,N_9198);
or U9539 (N_9539,N_9120,N_9143);
nor U9540 (N_9540,N_9210,N_9008);
and U9541 (N_9541,N_9161,N_9162);
nand U9542 (N_9542,N_9056,N_9210);
or U9543 (N_9543,N_9106,N_9025);
nor U9544 (N_9544,N_9119,N_9025);
and U9545 (N_9545,N_9139,N_9184);
or U9546 (N_9546,N_9043,N_9190);
nor U9547 (N_9547,N_9049,N_9194);
and U9548 (N_9548,N_9237,N_9140);
or U9549 (N_9549,N_9105,N_9243);
and U9550 (N_9550,N_9241,N_9092);
nor U9551 (N_9551,N_9299,N_9070);
and U9552 (N_9552,N_9119,N_9233);
nor U9553 (N_9553,N_9012,N_9194);
nor U9554 (N_9554,N_9056,N_9135);
or U9555 (N_9555,N_9154,N_9121);
or U9556 (N_9556,N_9162,N_9035);
nor U9557 (N_9557,N_9025,N_9248);
xnor U9558 (N_9558,N_9275,N_9156);
xnor U9559 (N_9559,N_9236,N_9109);
or U9560 (N_9560,N_9209,N_9091);
or U9561 (N_9561,N_9204,N_9263);
xnor U9562 (N_9562,N_9242,N_9047);
xnor U9563 (N_9563,N_9145,N_9177);
nor U9564 (N_9564,N_9277,N_9234);
xor U9565 (N_9565,N_9109,N_9155);
and U9566 (N_9566,N_9204,N_9208);
nand U9567 (N_9567,N_9049,N_9040);
and U9568 (N_9568,N_9279,N_9078);
nand U9569 (N_9569,N_9291,N_9274);
xnor U9570 (N_9570,N_9044,N_9253);
nor U9571 (N_9571,N_9183,N_9081);
and U9572 (N_9572,N_9260,N_9159);
and U9573 (N_9573,N_9152,N_9241);
and U9574 (N_9574,N_9180,N_9286);
nor U9575 (N_9575,N_9033,N_9281);
or U9576 (N_9576,N_9205,N_9177);
nor U9577 (N_9577,N_9219,N_9173);
xnor U9578 (N_9578,N_9270,N_9036);
or U9579 (N_9579,N_9245,N_9125);
nand U9580 (N_9580,N_9144,N_9199);
and U9581 (N_9581,N_9017,N_9050);
nor U9582 (N_9582,N_9275,N_9257);
and U9583 (N_9583,N_9052,N_9099);
and U9584 (N_9584,N_9153,N_9039);
and U9585 (N_9585,N_9177,N_9296);
nand U9586 (N_9586,N_9153,N_9175);
nand U9587 (N_9587,N_9081,N_9012);
and U9588 (N_9588,N_9166,N_9278);
and U9589 (N_9589,N_9096,N_9228);
or U9590 (N_9590,N_9265,N_9272);
nor U9591 (N_9591,N_9038,N_9265);
and U9592 (N_9592,N_9294,N_9264);
xnor U9593 (N_9593,N_9034,N_9107);
nand U9594 (N_9594,N_9017,N_9254);
nor U9595 (N_9595,N_9087,N_9162);
nor U9596 (N_9596,N_9156,N_9033);
xor U9597 (N_9597,N_9187,N_9099);
xnor U9598 (N_9598,N_9059,N_9097);
xor U9599 (N_9599,N_9148,N_9110);
nand U9600 (N_9600,N_9316,N_9582);
or U9601 (N_9601,N_9575,N_9501);
xor U9602 (N_9602,N_9586,N_9389);
or U9603 (N_9603,N_9326,N_9318);
xor U9604 (N_9604,N_9359,N_9541);
and U9605 (N_9605,N_9415,N_9462);
xnor U9606 (N_9606,N_9366,N_9311);
or U9607 (N_9607,N_9447,N_9437);
xnor U9608 (N_9608,N_9578,N_9539);
or U9609 (N_9609,N_9442,N_9473);
and U9610 (N_9610,N_9587,N_9385);
or U9611 (N_9611,N_9428,N_9474);
nand U9612 (N_9612,N_9546,N_9333);
and U9613 (N_9613,N_9553,N_9485);
xor U9614 (N_9614,N_9490,N_9577);
or U9615 (N_9615,N_9497,N_9537);
and U9616 (N_9616,N_9379,N_9436);
nor U9617 (N_9617,N_9457,N_9482);
nand U9618 (N_9618,N_9346,N_9470);
xnor U9619 (N_9619,N_9516,N_9304);
or U9620 (N_9620,N_9592,N_9580);
xnor U9621 (N_9621,N_9365,N_9336);
nor U9622 (N_9622,N_9488,N_9305);
xnor U9623 (N_9623,N_9591,N_9418);
nor U9624 (N_9624,N_9469,N_9355);
and U9625 (N_9625,N_9569,N_9322);
nand U9626 (N_9626,N_9453,N_9441);
xor U9627 (N_9627,N_9324,N_9500);
and U9628 (N_9628,N_9398,N_9425);
or U9629 (N_9629,N_9378,N_9350);
xnor U9630 (N_9630,N_9420,N_9405);
and U9631 (N_9631,N_9545,N_9341);
nor U9632 (N_9632,N_9339,N_9487);
and U9633 (N_9633,N_9459,N_9535);
or U9634 (N_9634,N_9328,N_9446);
xor U9635 (N_9635,N_9448,N_9544);
or U9636 (N_9636,N_9563,N_9596);
nand U9637 (N_9637,N_9404,N_9383);
and U9638 (N_9638,N_9517,N_9536);
nor U9639 (N_9639,N_9595,N_9481);
and U9640 (N_9640,N_9460,N_9438);
or U9641 (N_9641,N_9330,N_9550);
xor U9642 (N_9642,N_9337,N_9367);
xor U9643 (N_9643,N_9495,N_9409);
xor U9644 (N_9644,N_9507,N_9354);
or U9645 (N_9645,N_9549,N_9467);
or U9646 (N_9646,N_9340,N_9509);
and U9647 (N_9647,N_9444,N_9407);
nand U9648 (N_9648,N_9526,N_9524);
nand U9649 (N_9649,N_9466,N_9494);
nand U9650 (N_9650,N_9363,N_9332);
xnor U9651 (N_9651,N_9308,N_9432);
nor U9652 (N_9652,N_9583,N_9471);
nand U9653 (N_9653,N_9522,N_9394);
nor U9654 (N_9654,N_9499,N_9373);
xnor U9655 (N_9655,N_9468,N_9313);
and U9656 (N_9656,N_9338,N_9434);
or U9657 (N_9657,N_9506,N_9342);
nand U9658 (N_9658,N_9542,N_9504);
nor U9659 (N_9659,N_9307,N_9371);
xnor U9660 (N_9660,N_9464,N_9588);
xor U9661 (N_9661,N_9375,N_9343);
nand U9662 (N_9662,N_9317,N_9449);
nand U9663 (N_9663,N_9310,N_9478);
xnor U9664 (N_9664,N_9579,N_9380);
and U9665 (N_9665,N_9568,N_9412);
or U9666 (N_9666,N_9493,N_9439);
nor U9667 (N_9667,N_9456,N_9557);
xnor U9668 (N_9668,N_9514,N_9452);
xor U9669 (N_9669,N_9559,N_9312);
or U9670 (N_9670,N_9486,N_9356);
or U9671 (N_9671,N_9556,N_9406);
nor U9672 (N_9672,N_9574,N_9554);
xor U9673 (N_9673,N_9388,N_9523);
nand U9674 (N_9674,N_9430,N_9567);
and U9675 (N_9675,N_9445,N_9463);
xor U9676 (N_9676,N_9594,N_9361);
or U9677 (N_9677,N_9528,N_9533);
and U9678 (N_9678,N_9325,N_9521);
or U9679 (N_9679,N_9331,N_9433);
nand U9680 (N_9680,N_9454,N_9593);
nand U9681 (N_9681,N_9547,N_9302);
xor U9682 (N_9682,N_9314,N_9525);
nand U9683 (N_9683,N_9570,N_9476);
or U9684 (N_9684,N_9477,N_9515);
and U9685 (N_9685,N_9530,N_9529);
and U9686 (N_9686,N_9369,N_9465);
or U9687 (N_9687,N_9450,N_9353);
xor U9688 (N_9688,N_9540,N_9562);
nand U9689 (N_9689,N_9303,N_9374);
xnor U9690 (N_9690,N_9344,N_9508);
and U9691 (N_9691,N_9370,N_9560);
xor U9692 (N_9692,N_9598,N_9599);
nor U9693 (N_9693,N_9391,N_9372);
nor U9694 (N_9694,N_9424,N_9315);
nor U9695 (N_9695,N_9548,N_9360);
nor U9696 (N_9696,N_9349,N_9413);
or U9697 (N_9697,N_9503,N_9309);
nand U9698 (N_9698,N_9345,N_9502);
nor U9699 (N_9699,N_9489,N_9455);
and U9700 (N_9700,N_9443,N_9520);
and U9701 (N_9701,N_9584,N_9561);
nor U9702 (N_9702,N_9572,N_9484);
nand U9703 (N_9703,N_9390,N_9351);
nand U9704 (N_9704,N_9410,N_9411);
and U9705 (N_9705,N_9401,N_9399);
xnor U9706 (N_9706,N_9451,N_9571);
and U9707 (N_9707,N_9396,N_9422);
and U9708 (N_9708,N_9368,N_9513);
xnor U9709 (N_9709,N_9321,N_9306);
nor U9710 (N_9710,N_9421,N_9479);
and U9711 (N_9711,N_9597,N_9402);
nand U9712 (N_9712,N_9397,N_9414);
and U9713 (N_9713,N_9565,N_9519);
xor U9714 (N_9714,N_9300,N_9395);
nor U9715 (N_9715,N_9498,N_9511);
or U9716 (N_9716,N_9382,N_9552);
nor U9717 (N_9717,N_9461,N_9393);
nand U9718 (N_9718,N_9564,N_9417);
or U9719 (N_9719,N_9387,N_9435);
and U9720 (N_9720,N_9329,N_9358);
xnor U9721 (N_9721,N_9510,N_9301);
nor U9722 (N_9722,N_9551,N_9423);
xor U9723 (N_9723,N_9532,N_9555);
nor U9724 (N_9724,N_9348,N_9419);
and U9725 (N_9725,N_9392,N_9429);
nand U9726 (N_9726,N_9431,N_9403);
xnor U9727 (N_9727,N_9319,N_9352);
xor U9728 (N_9728,N_9381,N_9362);
xor U9729 (N_9729,N_9483,N_9585);
xnor U9730 (N_9730,N_9573,N_9400);
and U9731 (N_9731,N_9491,N_9518);
or U9732 (N_9732,N_9386,N_9357);
xor U9733 (N_9733,N_9505,N_9377);
nand U9734 (N_9734,N_9492,N_9472);
and U9735 (N_9735,N_9534,N_9327);
nand U9736 (N_9736,N_9364,N_9334);
or U9737 (N_9737,N_9335,N_9527);
and U9738 (N_9738,N_9384,N_9440);
or U9739 (N_9739,N_9566,N_9376);
xor U9740 (N_9740,N_9427,N_9589);
xnor U9741 (N_9741,N_9581,N_9416);
or U9742 (N_9742,N_9558,N_9590);
nand U9743 (N_9743,N_9512,N_9531);
and U9744 (N_9744,N_9323,N_9475);
or U9745 (N_9745,N_9426,N_9347);
and U9746 (N_9746,N_9320,N_9496);
xor U9747 (N_9747,N_9458,N_9538);
xor U9748 (N_9748,N_9480,N_9543);
or U9749 (N_9749,N_9408,N_9576);
and U9750 (N_9750,N_9413,N_9381);
nor U9751 (N_9751,N_9585,N_9492);
nor U9752 (N_9752,N_9341,N_9551);
nand U9753 (N_9753,N_9394,N_9469);
and U9754 (N_9754,N_9544,N_9426);
and U9755 (N_9755,N_9343,N_9535);
or U9756 (N_9756,N_9348,N_9376);
xor U9757 (N_9757,N_9587,N_9416);
nor U9758 (N_9758,N_9567,N_9394);
nand U9759 (N_9759,N_9472,N_9324);
or U9760 (N_9760,N_9428,N_9480);
and U9761 (N_9761,N_9539,N_9562);
xnor U9762 (N_9762,N_9580,N_9371);
and U9763 (N_9763,N_9381,N_9531);
xor U9764 (N_9764,N_9358,N_9364);
xor U9765 (N_9765,N_9304,N_9554);
nand U9766 (N_9766,N_9458,N_9466);
nor U9767 (N_9767,N_9597,N_9466);
and U9768 (N_9768,N_9396,N_9574);
and U9769 (N_9769,N_9467,N_9503);
nor U9770 (N_9770,N_9319,N_9446);
nor U9771 (N_9771,N_9566,N_9574);
nand U9772 (N_9772,N_9327,N_9567);
or U9773 (N_9773,N_9512,N_9433);
nand U9774 (N_9774,N_9482,N_9401);
and U9775 (N_9775,N_9393,N_9488);
xnor U9776 (N_9776,N_9582,N_9417);
xnor U9777 (N_9777,N_9459,N_9429);
or U9778 (N_9778,N_9536,N_9487);
or U9779 (N_9779,N_9463,N_9365);
nand U9780 (N_9780,N_9409,N_9536);
nor U9781 (N_9781,N_9358,N_9494);
xor U9782 (N_9782,N_9335,N_9346);
nor U9783 (N_9783,N_9347,N_9461);
or U9784 (N_9784,N_9585,N_9524);
or U9785 (N_9785,N_9368,N_9592);
and U9786 (N_9786,N_9410,N_9525);
xnor U9787 (N_9787,N_9348,N_9527);
and U9788 (N_9788,N_9324,N_9304);
and U9789 (N_9789,N_9593,N_9415);
nor U9790 (N_9790,N_9552,N_9355);
nor U9791 (N_9791,N_9318,N_9307);
nand U9792 (N_9792,N_9520,N_9560);
and U9793 (N_9793,N_9546,N_9589);
and U9794 (N_9794,N_9482,N_9368);
and U9795 (N_9795,N_9439,N_9435);
and U9796 (N_9796,N_9451,N_9582);
or U9797 (N_9797,N_9308,N_9358);
xnor U9798 (N_9798,N_9470,N_9513);
xnor U9799 (N_9799,N_9480,N_9327);
nor U9800 (N_9800,N_9578,N_9503);
xor U9801 (N_9801,N_9340,N_9366);
and U9802 (N_9802,N_9370,N_9399);
or U9803 (N_9803,N_9520,N_9464);
xor U9804 (N_9804,N_9491,N_9326);
or U9805 (N_9805,N_9506,N_9451);
nor U9806 (N_9806,N_9478,N_9567);
xnor U9807 (N_9807,N_9363,N_9386);
nor U9808 (N_9808,N_9369,N_9431);
nand U9809 (N_9809,N_9372,N_9445);
nand U9810 (N_9810,N_9576,N_9481);
and U9811 (N_9811,N_9332,N_9360);
or U9812 (N_9812,N_9546,N_9424);
or U9813 (N_9813,N_9415,N_9404);
xor U9814 (N_9814,N_9517,N_9467);
and U9815 (N_9815,N_9491,N_9463);
and U9816 (N_9816,N_9506,N_9335);
nand U9817 (N_9817,N_9351,N_9447);
or U9818 (N_9818,N_9413,N_9481);
and U9819 (N_9819,N_9485,N_9454);
xor U9820 (N_9820,N_9313,N_9336);
and U9821 (N_9821,N_9457,N_9406);
and U9822 (N_9822,N_9458,N_9306);
nor U9823 (N_9823,N_9567,N_9492);
and U9824 (N_9824,N_9571,N_9598);
xor U9825 (N_9825,N_9567,N_9435);
nand U9826 (N_9826,N_9387,N_9517);
and U9827 (N_9827,N_9575,N_9428);
xor U9828 (N_9828,N_9581,N_9522);
nand U9829 (N_9829,N_9529,N_9433);
or U9830 (N_9830,N_9540,N_9394);
and U9831 (N_9831,N_9409,N_9458);
nor U9832 (N_9832,N_9504,N_9561);
nand U9833 (N_9833,N_9587,N_9490);
nand U9834 (N_9834,N_9413,N_9554);
and U9835 (N_9835,N_9424,N_9352);
nor U9836 (N_9836,N_9378,N_9560);
or U9837 (N_9837,N_9509,N_9316);
and U9838 (N_9838,N_9321,N_9303);
xor U9839 (N_9839,N_9406,N_9374);
or U9840 (N_9840,N_9318,N_9423);
xor U9841 (N_9841,N_9555,N_9353);
nand U9842 (N_9842,N_9403,N_9561);
or U9843 (N_9843,N_9587,N_9345);
or U9844 (N_9844,N_9585,N_9468);
or U9845 (N_9845,N_9553,N_9336);
nand U9846 (N_9846,N_9529,N_9514);
or U9847 (N_9847,N_9593,N_9558);
and U9848 (N_9848,N_9452,N_9376);
nand U9849 (N_9849,N_9339,N_9355);
xnor U9850 (N_9850,N_9576,N_9534);
nand U9851 (N_9851,N_9338,N_9436);
xnor U9852 (N_9852,N_9323,N_9433);
xnor U9853 (N_9853,N_9392,N_9330);
xor U9854 (N_9854,N_9437,N_9511);
nor U9855 (N_9855,N_9331,N_9316);
xnor U9856 (N_9856,N_9337,N_9511);
nor U9857 (N_9857,N_9480,N_9576);
or U9858 (N_9858,N_9501,N_9301);
or U9859 (N_9859,N_9535,N_9352);
nor U9860 (N_9860,N_9331,N_9363);
and U9861 (N_9861,N_9372,N_9351);
xor U9862 (N_9862,N_9374,N_9319);
and U9863 (N_9863,N_9377,N_9523);
nor U9864 (N_9864,N_9448,N_9482);
nor U9865 (N_9865,N_9371,N_9453);
nand U9866 (N_9866,N_9517,N_9568);
nor U9867 (N_9867,N_9586,N_9450);
nor U9868 (N_9868,N_9413,N_9304);
nor U9869 (N_9869,N_9515,N_9360);
nor U9870 (N_9870,N_9548,N_9581);
nor U9871 (N_9871,N_9364,N_9409);
and U9872 (N_9872,N_9500,N_9468);
or U9873 (N_9873,N_9572,N_9388);
xor U9874 (N_9874,N_9395,N_9339);
and U9875 (N_9875,N_9351,N_9585);
nand U9876 (N_9876,N_9510,N_9482);
nor U9877 (N_9877,N_9442,N_9332);
nand U9878 (N_9878,N_9560,N_9374);
xor U9879 (N_9879,N_9431,N_9566);
xor U9880 (N_9880,N_9567,N_9456);
and U9881 (N_9881,N_9569,N_9500);
and U9882 (N_9882,N_9322,N_9367);
nor U9883 (N_9883,N_9335,N_9320);
xnor U9884 (N_9884,N_9487,N_9314);
nand U9885 (N_9885,N_9417,N_9535);
and U9886 (N_9886,N_9471,N_9413);
xnor U9887 (N_9887,N_9525,N_9458);
or U9888 (N_9888,N_9549,N_9510);
and U9889 (N_9889,N_9468,N_9568);
or U9890 (N_9890,N_9406,N_9444);
nor U9891 (N_9891,N_9457,N_9460);
and U9892 (N_9892,N_9439,N_9593);
nor U9893 (N_9893,N_9507,N_9395);
nand U9894 (N_9894,N_9384,N_9396);
nand U9895 (N_9895,N_9335,N_9467);
nand U9896 (N_9896,N_9515,N_9341);
xor U9897 (N_9897,N_9339,N_9581);
nand U9898 (N_9898,N_9420,N_9426);
and U9899 (N_9899,N_9335,N_9321);
nor U9900 (N_9900,N_9630,N_9752);
nand U9901 (N_9901,N_9765,N_9891);
and U9902 (N_9902,N_9804,N_9818);
nor U9903 (N_9903,N_9869,N_9790);
xnor U9904 (N_9904,N_9874,N_9870);
xnor U9905 (N_9905,N_9830,N_9724);
nor U9906 (N_9906,N_9829,N_9863);
and U9907 (N_9907,N_9867,N_9602);
nand U9908 (N_9908,N_9730,N_9606);
nand U9909 (N_9909,N_9616,N_9875);
nor U9910 (N_9910,N_9739,N_9771);
or U9911 (N_9911,N_9899,N_9727);
nor U9912 (N_9912,N_9850,N_9607);
nand U9913 (N_9913,N_9643,N_9601);
or U9914 (N_9914,N_9784,N_9699);
and U9915 (N_9915,N_9849,N_9872);
xnor U9916 (N_9916,N_9675,N_9609);
nand U9917 (N_9917,N_9729,N_9682);
xnor U9918 (N_9918,N_9746,N_9839);
and U9919 (N_9919,N_9892,N_9707);
or U9920 (N_9920,N_9884,N_9705);
and U9921 (N_9921,N_9890,N_9761);
or U9922 (N_9922,N_9661,N_9670);
nand U9923 (N_9923,N_9858,N_9668);
xnor U9924 (N_9924,N_9774,N_9702);
xor U9925 (N_9925,N_9836,N_9728);
xor U9926 (N_9926,N_9660,N_9690);
nor U9927 (N_9927,N_9821,N_9676);
nor U9928 (N_9928,N_9600,N_9637);
nor U9929 (N_9929,N_9614,N_9855);
or U9930 (N_9930,N_9666,N_9859);
nor U9931 (N_9931,N_9671,N_9683);
xor U9932 (N_9932,N_9696,N_9664);
xor U9933 (N_9933,N_9827,N_9642);
or U9934 (N_9934,N_9810,N_9603);
or U9935 (N_9935,N_9805,N_9889);
or U9936 (N_9936,N_9613,N_9681);
nor U9937 (N_9937,N_9797,N_9716);
nand U9938 (N_9938,N_9706,N_9621);
and U9939 (N_9939,N_9896,N_9709);
or U9940 (N_9940,N_9733,N_9738);
nand U9941 (N_9941,N_9608,N_9799);
or U9942 (N_9942,N_9880,N_9641);
and U9943 (N_9943,N_9632,N_9680);
or U9944 (N_9944,N_9640,N_9841);
xor U9945 (N_9945,N_9747,N_9713);
xnor U9946 (N_9946,N_9831,N_9644);
and U9947 (N_9947,N_9897,N_9749);
nand U9948 (N_9948,N_9866,N_9835);
nor U9949 (N_9949,N_9865,N_9610);
and U9950 (N_9950,N_9758,N_9654);
or U9951 (N_9951,N_9624,N_9767);
nand U9952 (N_9952,N_9833,N_9878);
nand U9953 (N_9953,N_9822,N_9791);
xnor U9954 (N_9954,N_9781,N_9742);
nor U9955 (N_9955,N_9740,N_9698);
nor U9956 (N_9956,N_9677,N_9674);
and U9957 (N_9957,N_9751,N_9695);
and U9958 (N_9958,N_9652,N_9647);
xor U9959 (N_9959,N_9809,N_9672);
nor U9960 (N_9960,N_9843,N_9895);
nand U9961 (N_9961,N_9755,N_9667);
nor U9962 (N_9962,N_9851,N_9658);
or U9963 (N_9963,N_9622,N_9877);
xor U9964 (N_9964,N_9750,N_9745);
or U9965 (N_9965,N_9852,N_9636);
and U9966 (N_9966,N_9785,N_9620);
nor U9967 (N_9967,N_9689,N_9824);
xor U9968 (N_9968,N_9722,N_9625);
or U9969 (N_9969,N_9772,N_9832);
or U9970 (N_9970,N_9646,N_9619);
xor U9971 (N_9971,N_9812,N_9766);
xnor U9972 (N_9972,N_9684,N_9871);
nor U9973 (N_9973,N_9648,N_9720);
nand U9974 (N_9974,N_9725,N_9775);
and U9975 (N_9975,N_9834,N_9881);
nand U9976 (N_9976,N_9697,N_9762);
nor U9977 (N_9977,N_9825,N_9817);
or U9978 (N_9978,N_9717,N_9873);
nand U9979 (N_9979,N_9703,N_9757);
and U9980 (N_9980,N_9686,N_9811);
or U9981 (N_9981,N_9789,N_9687);
nand U9982 (N_9982,N_9898,N_9793);
and U9983 (N_9983,N_9788,N_9856);
xnor U9984 (N_9984,N_9826,N_9795);
or U9985 (N_9985,N_9768,N_9773);
and U9986 (N_9986,N_9885,N_9823);
nand U9987 (N_9987,N_9718,N_9876);
or U9988 (N_9988,N_9659,N_9688);
nand U9989 (N_9989,N_9678,N_9753);
and U9990 (N_9990,N_9715,N_9854);
and U9991 (N_9991,N_9803,N_9741);
nor U9992 (N_9992,N_9828,N_9612);
and U9993 (N_9993,N_9649,N_9615);
or U9994 (N_9994,N_9886,N_9769);
xnor U9995 (N_9995,N_9846,N_9759);
nand U9996 (N_9996,N_9853,N_9691);
xor U9997 (N_9997,N_9813,N_9737);
xnor U9998 (N_9998,N_9663,N_9662);
nand U9999 (N_9999,N_9845,N_9631);
and U10000 (N_10000,N_9888,N_9627);
nand U10001 (N_10001,N_9710,N_9657);
or U10002 (N_10002,N_9883,N_9712);
xnor U10003 (N_10003,N_9635,N_9633);
and U10004 (N_10004,N_9780,N_9879);
or U10005 (N_10005,N_9604,N_9744);
xnor U10006 (N_10006,N_9770,N_9882);
nand U10007 (N_10007,N_9779,N_9618);
and U10008 (N_10008,N_9794,N_9634);
and U10009 (N_10009,N_9650,N_9694);
xor U10010 (N_10010,N_9837,N_9669);
nor U10011 (N_10011,N_9665,N_9651);
nand U10012 (N_10012,N_9894,N_9864);
nand U10013 (N_10013,N_9814,N_9748);
and U10014 (N_10014,N_9655,N_9801);
and U10015 (N_10015,N_9816,N_9653);
xor U10016 (N_10016,N_9731,N_9798);
nand U10017 (N_10017,N_9819,N_9764);
nand U10018 (N_10018,N_9645,N_9685);
nor U10019 (N_10019,N_9778,N_9626);
or U10020 (N_10020,N_9763,N_9844);
xor U10021 (N_10021,N_9815,N_9796);
nand U10022 (N_10022,N_9629,N_9760);
nand U10023 (N_10023,N_9887,N_9692);
nor U10024 (N_10024,N_9714,N_9701);
nor U10025 (N_10025,N_9656,N_9617);
xnor U10026 (N_10026,N_9673,N_9776);
and U10027 (N_10027,N_9708,N_9806);
nand U10028 (N_10028,N_9719,N_9726);
xnor U10029 (N_10029,N_9623,N_9848);
nand U10030 (N_10030,N_9743,N_9787);
nor U10031 (N_10031,N_9860,N_9840);
nand U10032 (N_10032,N_9721,N_9807);
nand U10033 (N_10033,N_9704,N_9783);
nand U10034 (N_10034,N_9638,N_9736);
nor U10035 (N_10035,N_9857,N_9723);
xnor U10036 (N_10036,N_9732,N_9786);
nand U10037 (N_10037,N_9734,N_9802);
nor U10038 (N_10038,N_9842,N_9800);
and U10039 (N_10039,N_9782,N_9893);
and U10040 (N_10040,N_9868,N_9700);
nor U10041 (N_10041,N_9605,N_9754);
and U10042 (N_10042,N_9611,N_9693);
or U10043 (N_10043,N_9820,N_9792);
and U10044 (N_10044,N_9735,N_9861);
nor U10045 (N_10045,N_9628,N_9711);
nand U10046 (N_10046,N_9847,N_9756);
xor U10047 (N_10047,N_9838,N_9679);
or U10048 (N_10048,N_9777,N_9639);
and U10049 (N_10049,N_9862,N_9808);
xnor U10050 (N_10050,N_9779,N_9896);
and U10051 (N_10051,N_9777,N_9807);
and U10052 (N_10052,N_9796,N_9778);
nor U10053 (N_10053,N_9638,N_9748);
or U10054 (N_10054,N_9814,N_9669);
nand U10055 (N_10055,N_9850,N_9681);
or U10056 (N_10056,N_9742,N_9602);
and U10057 (N_10057,N_9726,N_9764);
and U10058 (N_10058,N_9634,N_9824);
nand U10059 (N_10059,N_9893,N_9625);
nor U10060 (N_10060,N_9824,N_9632);
nor U10061 (N_10061,N_9756,N_9867);
xor U10062 (N_10062,N_9838,N_9873);
or U10063 (N_10063,N_9824,N_9853);
xor U10064 (N_10064,N_9856,N_9796);
nor U10065 (N_10065,N_9893,N_9882);
nor U10066 (N_10066,N_9656,N_9785);
nor U10067 (N_10067,N_9668,N_9761);
xor U10068 (N_10068,N_9894,N_9861);
nor U10069 (N_10069,N_9812,N_9778);
nand U10070 (N_10070,N_9705,N_9701);
xor U10071 (N_10071,N_9641,N_9622);
xnor U10072 (N_10072,N_9678,N_9877);
or U10073 (N_10073,N_9835,N_9877);
and U10074 (N_10074,N_9623,N_9666);
xnor U10075 (N_10075,N_9648,N_9621);
nand U10076 (N_10076,N_9726,N_9656);
nor U10077 (N_10077,N_9871,N_9682);
xor U10078 (N_10078,N_9780,N_9633);
and U10079 (N_10079,N_9729,N_9718);
xnor U10080 (N_10080,N_9683,N_9612);
or U10081 (N_10081,N_9830,N_9670);
nand U10082 (N_10082,N_9731,N_9650);
or U10083 (N_10083,N_9848,N_9853);
or U10084 (N_10084,N_9654,N_9821);
nor U10085 (N_10085,N_9790,N_9708);
or U10086 (N_10086,N_9634,N_9815);
nor U10087 (N_10087,N_9699,N_9810);
nand U10088 (N_10088,N_9836,N_9871);
or U10089 (N_10089,N_9784,N_9771);
nor U10090 (N_10090,N_9842,N_9701);
and U10091 (N_10091,N_9762,N_9827);
nor U10092 (N_10092,N_9678,N_9819);
nor U10093 (N_10093,N_9745,N_9899);
and U10094 (N_10094,N_9703,N_9843);
nand U10095 (N_10095,N_9704,N_9601);
xnor U10096 (N_10096,N_9670,N_9668);
nand U10097 (N_10097,N_9808,N_9878);
nor U10098 (N_10098,N_9723,N_9837);
nand U10099 (N_10099,N_9888,N_9710);
xor U10100 (N_10100,N_9673,N_9662);
nand U10101 (N_10101,N_9818,N_9609);
xnor U10102 (N_10102,N_9663,N_9823);
nand U10103 (N_10103,N_9685,N_9609);
nand U10104 (N_10104,N_9647,N_9690);
xnor U10105 (N_10105,N_9649,N_9850);
nor U10106 (N_10106,N_9807,N_9655);
xor U10107 (N_10107,N_9657,N_9772);
xor U10108 (N_10108,N_9785,N_9844);
xor U10109 (N_10109,N_9680,N_9788);
or U10110 (N_10110,N_9835,N_9656);
and U10111 (N_10111,N_9653,N_9853);
nand U10112 (N_10112,N_9716,N_9675);
nor U10113 (N_10113,N_9683,N_9626);
xnor U10114 (N_10114,N_9606,N_9683);
xnor U10115 (N_10115,N_9676,N_9628);
nor U10116 (N_10116,N_9692,N_9774);
nand U10117 (N_10117,N_9733,N_9750);
xnor U10118 (N_10118,N_9860,N_9739);
or U10119 (N_10119,N_9849,N_9602);
nor U10120 (N_10120,N_9744,N_9685);
or U10121 (N_10121,N_9693,N_9667);
nand U10122 (N_10122,N_9660,N_9795);
and U10123 (N_10123,N_9698,N_9623);
nand U10124 (N_10124,N_9634,N_9662);
and U10125 (N_10125,N_9796,N_9635);
xnor U10126 (N_10126,N_9771,N_9661);
xor U10127 (N_10127,N_9770,N_9629);
or U10128 (N_10128,N_9680,N_9709);
xnor U10129 (N_10129,N_9883,N_9743);
and U10130 (N_10130,N_9634,N_9813);
nor U10131 (N_10131,N_9711,N_9804);
nand U10132 (N_10132,N_9716,N_9687);
or U10133 (N_10133,N_9778,N_9642);
and U10134 (N_10134,N_9608,N_9812);
nand U10135 (N_10135,N_9680,N_9742);
xor U10136 (N_10136,N_9701,N_9767);
xnor U10137 (N_10137,N_9638,N_9822);
xnor U10138 (N_10138,N_9682,N_9689);
nor U10139 (N_10139,N_9857,N_9664);
nand U10140 (N_10140,N_9845,N_9654);
nand U10141 (N_10141,N_9852,N_9804);
and U10142 (N_10142,N_9778,N_9838);
or U10143 (N_10143,N_9810,N_9705);
or U10144 (N_10144,N_9720,N_9654);
and U10145 (N_10145,N_9755,N_9615);
nor U10146 (N_10146,N_9811,N_9773);
or U10147 (N_10147,N_9789,N_9867);
nand U10148 (N_10148,N_9621,N_9732);
nand U10149 (N_10149,N_9851,N_9607);
nor U10150 (N_10150,N_9720,N_9839);
or U10151 (N_10151,N_9743,N_9794);
nor U10152 (N_10152,N_9699,N_9781);
or U10153 (N_10153,N_9774,N_9786);
or U10154 (N_10154,N_9668,N_9892);
nor U10155 (N_10155,N_9731,N_9862);
xor U10156 (N_10156,N_9761,N_9866);
nor U10157 (N_10157,N_9705,N_9717);
or U10158 (N_10158,N_9786,N_9663);
xor U10159 (N_10159,N_9846,N_9876);
nand U10160 (N_10160,N_9637,N_9737);
and U10161 (N_10161,N_9816,N_9661);
or U10162 (N_10162,N_9881,N_9615);
nand U10163 (N_10163,N_9742,N_9747);
or U10164 (N_10164,N_9868,N_9600);
or U10165 (N_10165,N_9869,N_9672);
and U10166 (N_10166,N_9751,N_9798);
and U10167 (N_10167,N_9752,N_9686);
and U10168 (N_10168,N_9765,N_9702);
or U10169 (N_10169,N_9703,N_9839);
nor U10170 (N_10170,N_9809,N_9859);
and U10171 (N_10171,N_9829,N_9824);
and U10172 (N_10172,N_9774,N_9882);
and U10173 (N_10173,N_9790,N_9652);
nor U10174 (N_10174,N_9637,N_9605);
nand U10175 (N_10175,N_9891,N_9786);
nor U10176 (N_10176,N_9758,N_9844);
nor U10177 (N_10177,N_9719,N_9802);
or U10178 (N_10178,N_9684,N_9836);
nand U10179 (N_10179,N_9780,N_9815);
xnor U10180 (N_10180,N_9794,N_9861);
or U10181 (N_10181,N_9799,N_9604);
xor U10182 (N_10182,N_9783,N_9790);
and U10183 (N_10183,N_9724,N_9655);
nand U10184 (N_10184,N_9820,N_9605);
or U10185 (N_10185,N_9789,N_9800);
nor U10186 (N_10186,N_9885,N_9600);
xnor U10187 (N_10187,N_9721,N_9882);
nand U10188 (N_10188,N_9892,N_9679);
or U10189 (N_10189,N_9732,N_9886);
xnor U10190 (N_10190,N_9871,N_9886);
or U10191 (N_10191,N_9797,N_9685);
xnor U10192 (N_10192,N_9802,N_9806);
or U10193 (N_10193,N_9839,N_9662);
and U10194 (N_10194,N_9647,N_9628);
or U10195 (N_10195,N_9676,N_9607);
or U10196 (N_10196,N_9663,N_9746);
or U10197 (N_10197,N_9612,N_9618);
nor U10198 (N_10198,N_9796,N_9805);
nor U10199 (N_10199,N_9880,N_9773);
nor U10200 (N_10200,N_10004,N_9998);
and U10201 (N_10201,N_9957,N_10187);
xor U10202 (N_10202,N_10092,N_10001);
or U10203 (N_10203,N_10182,N_9974);
nor U10204 (N_10204,N_10107,N_10086);
nor U10205 (N_10205,N_10079,N_10173);
nand U10206 (N_10206,N_10090,N_10109);
or U10207 (N_10207,N_10037,N_10171);
and U10208 (N_10208,N_10060,N_10024);
nand U10209 (N_10209,N_10198,N_10053);
or U10210 (N_10210,N_10080,N_10073);
nor U10211 (N_10211,N_10132,N_9990);
nor U10212 (N_10212,N_10137,N_10133);
nor U10213 (N_10213,N_9965,N_10180);
and U10214 (N_10214,N_10077,N_10027);
nor U10215 (N_10215,N_10046,N_10002);
or U10216 (N_10216,N_10050,N_9915);
or U10217 (N_10217,N_10070,N_9983);
nand U10218 (N_10218,N_9938,N_10156);
nand U10219 (N_10219,N_10081,N_10016);
nand U10220 (N_10220,N_10183,N_9981);
xnor U10221 (N_10221,N_10056,N_9958);
nand U10222 (N_10222,N_9970,N_9921);
nor U10223 (N_10223,N_10095,N_10121);
nand U10224 (N_10224,N_10075,N_10142);
nor U10225 (N_10225,N_10176,N_10150);
nand U10226 (N_10226,N_10148,N_10048);
xnor U10227 (N_10227,N_10055,N_9948);
nand U10228 (N_10228,N_10169,N_10188);
nand U10229 (N_10229,N_10094,N_10116);
or U10230 (N_10230,N_9950,N_9968);
and U10231 (N_10231,N_10194,N_9919);
nor U10232 (N_10232,N_9995,N_9929);
nor U10233 (N_10233,N_10172,N_10112);
nand U10234 (N_10234,N_10106,N_10102);
xnor U10235 (N_10235,N_9932,N_10043);
xor U10236 (N_10236,N_10145,N_10057);
nand U10237 (N_10237,N_9939,N_10098);
xor U10238 (N_10238,N_10199,N_10162);
or U10239 (N_10239,N_9914,N_10006);
xor U10240 (N_10240,N_10038,N_10120);
or U10241 (N_10241,N_10058,N_10104);
nor U10242 (N_10242,N_10147,N_10023);
nand U10243 (N_10243,N_10149,N_10039);
xor U10244 (N_10244,N_9991,N_10026);
nor U10245 (N_10245,N_9975,N_10178);
nand U10246 (N_10246,N_10101,N_10012);
nor U10247 (N_10247,N_10118,N_9993);
nor U10248 (N_10248,N_10139,N_9987);
xor U10249 (N_10249,N_9946,N_10193);
nand U10250 (N_10250,N_10088,N_9908);
or U10251 (N_10251,N_10007,N_9930);
nor U10252 (N_10252,N_10126,N_9935);
nand U10253 (N_10253,N_9927,N_9959);
xnor U10254 (N_10254,N_10168,N_10052);
and U10255 (N_10255,N_10017,N_10008);
nor U10256 (N_10256,N_10123,N_10034);
nor U10257 (N_10257,N_9985,N_9934);
or U10258 (N_10258,N_9996,N_10159);
nand U10259 (N_10259,N_10181,N_10136);
xor U10260 (N_10260,N_10059,N_9924);
and U10261 (N_10261,N_9951,N_9967);
xnor U10262 (N_10262,N_10113,N_10035);
or U10263 (N_10263,N_9902,N_9904);
nor U10264 (N_10264,N_10076,N_9909);
nor U10265 (N_10265,N_9907,N_9945);
xnor U10266 (N_10266,N_10018,N_10068);
xnor U10267 (N_10267,N_10146,N_10114);
or U10268 (N_10268,N_10042,N_10165);
and U10269 (N_10269,N_10031,N_10124);
or U10270 (N_10270,N_10011,N_9906);
or U10271 (N_10271,N_9933,N_9905);
or U10272 (N_10272,N_10019,N_10122);
xor U10273 (N_10273,N_10128,N_9940);
nand U10274 (N_10274,N_10108,N_9936);
or U10275 (N_10275,N_10161,N_10000);
and U10276 (N_10276,N_9964,N_10100);
and U10277 (N_10277,N_10190,N_10025);
xnor U10278 (N_10278,N_9997,N_10192);
nand U10279 (N_10279,N_10195,N_10189);
nand U10280 (N_10280,N_10044,N_9913);
and U10281 (N_10281,N_9989,N_10065);
or U10282 (N_10282,N_9963,N_9984);
nand U10283 (N_10283,N_10041,N_9973);
and U10284 (N_10284,N_10164,N_9971);
and U10285 (N_10285,N_10158,N_10045);
and U10286 (N_10286,N_10167,N_10117);
xnor U10287 (N_10287,N_9961,N_9947);
nand U10288 (N_10288,N_10028,N_9994);
nor U10289 (N_10289,N_9976,N_10141);
nor U10290 (N_10290,N_10096,N_9978);
and U10291 (N_10291,N_9900,N_10138);
xor U10292 (N_10292,N_9979,N_10066);
and U10293 (N_10293,N_10036,N_10071);
nand U10294 (N_10294,N_10040,N_10054);
and U10295 (N_10295,N_9926,N_10155);
or U10296 (N_10296,N_10089,N_10085);
xnor U10297 (N_10297,N_10022,N_9925);
xor U10298 (N_10298,N_10067,N_9986);
or U10299 (N_10299,N_10175,N_10051);
and U10300 (N_10300,N_10144,N_10115);
or U10301 (N_10301,N_10062,N_9918);
nor U10302 (N_10302,N_10072,N_10033);
nand U10303 (N_10303,N_9928,N_9910);
nand U10304 (N_10304,N_10134,N_10082);
nand U10305 (N_10305,N_10143,N_9955);
nand U10306 (N_10306,N_9988,N_10170);
nand U10307 (N_10307,N_10166,N_9916);
nor U10308 (N_10308,N_9942,N_10013);
and U10309 (N_10309,N_10103,N_10020);
nand U10310 (N_10310,N_10015,N_10069);
and U10311 (N_10311,N_9901,N_10030);
and U10312 (N_10312,N_10163,N_10135);
xnor U10313 (N_10313,N_9911,N_10152);
or U10314 (N_10314,N_10083,N_10021);
nor U10315 (N_10315,N_10047,N_9917);
or U10316 (N_10316,N_10177,N_10097);
nand U10317 (N_10317,N_10160,N_10009);
xnor U10318 (N_10318,N_9949,N_10078);
xnor U10319 (N_10319,N_10179,N_9944);
xor U10320 (N_10320,N_10196,N_9952);
xor U10321 (N_10321,N_10130,N_10110);
nand U10322 (N_10322,N_10131,N_9992);
nand U10323 (N_10323,N_10105,N_10061);
nand U10324 (N_10324,N_10111,N_10010);
or U10325 (N_10325,N_10084,N_9972);
nand U10326 (N_10326,N_10032,N_10197);
or U10327 (N_10327,N_10029,N_9980);
and U10328 (N_10328,N_9977,N_10151);
xor U10329 (N_10329,N_9969,N_10154);
nor U10330 (N_10330,N_10184,N_10125);
nor U10331 (N_10331,N_10087,N_10185);
and U10332 (N_10332,N_10191,N_9982);
and U10333 (N_10333,N_9943,N_10140);
nor U10334 (N_10334,N_10049,N_10174);
nand U10335 (N_10335,N_9941,N_10003);
nor U10336 (N_10336,N_9923,N_9920);
and U10337 (N_10337,N_10153,N_10186);
or U10338 (N_10338,N_10064,N_10129);
nor U10339 (N_10339,N_10074,N_9912);
xnor U10340 (N_10340,N_9966,N_10157);
or U10341 (N_10341,N_9960,N_9903);
nand U10342 (N_10342,N_10014,N_9937);
and U10343 (N_10343,N_9931,N_9954);
or U10344 (N_10344,N_9999,N_10091);
or U10345 (N_10345,N_9962,N_10099);
xor U10346 (N_10346,N_10127,N_9922);
and U10347 (N_10347,N_10063,N_10005);
nand U10348 (N_10348,N_9956,N_9953);
or U10349 (N_10349,N_10093,N_10119);
xnor U10350 (N_10350,N_10047,N_10119);
xor U10351 (N_10351,N_9909,N_10095);
nor U10352 (N_10352,N_10165,N_10060);
nor U10353 (N_10353,N_10015,N_10009);
nand U10354 (N_10354,N_9947,N_10044);
or U10355 (N_10355,N_10128,N_10033);
xnor U10356 (N_10356,N_9982,N_9910);
nand U10357 (N_10357,N_10199,N_9911);
xnor U10358 (N_10358,N_10089,N_10142);
xnor U10359 (N_10359,N_10080,N_9924);
and U10360 (N_10360,N_10127,N_10068);
nand U10361 (N_10361,N_9918,N_9915);
or U10362 (N_10362,N_10120,N_10133);
or U10363 (N_10363,N_9929,N_9924);
nand U10364 (N_10364,N_10131,N_10043);
nand U10365 (N_10365,N_10036,N_10146);
and U10366 (N_10366,N_10012,N_9954);
nor U10367 (N_10367,N_10172,N_10033);
nor U10368 (N_10368,N_10155,N_10020);
nor U10369 (N_10369,N_10176,N_10119);
nand U10370 (N_10370,N_10108,N_10062);
nand U10371 (N_10371,N_10055,N_9955);
xor U10372 (N_10372,N_10005,N_10170);
xnor U10373 (N_10373,N_9980,N_9926);
nand U10374 (N_10374,N_10187,N_10043);
or U10375 (N_10375,N_9900,N_9987);
or U10376 (N_10376,N_9997,N_9916);
xnor U10377 (N_10377,N_10091,N_9983);
nor U10378 (N_10378,N_10154,N_10084);
and U10379 (N_10379,N_10006,N_10091);
nand U10380 (N_10380,N_9926,N_9941);
xor U10381 (N_10381,N_10008,N_10136);
xor U10382 (N_10382,N_9943,N_10030);
nor U10383 (N_10383,N_10162,N_10128);
xor U10384 (N_10384,N_9914,N_10180);
xor U10385 (N_10385,N_9900,N_10150);
and U10386 (N_10386,N_10139,N_10028);
xor U10387 (N_10387,N_10090,N_9915);
and U10388 (N_10388,N_9952,N_9932);
and U10389 (N_10389,N_10070,N_10062);
or U10390 (N_10390,N_10133,N_10105);
xnor U10391 (N_10391,N_9985,N_10196);
nand U10392 (N_10392,N_10025,N_10143);
nor U10393 (N_10393,N_10158,N_10009);
nor U10394 (N_10394,N_10144,N_10079);
nor U10395 (N_10395,N_10061,N_10116);
xor U10396 (N_10396,N_10152,N_10018);
xnor U10397 (N_10397,N_10068,N_9968);
or U10398 (N_10398,N_10133,N_10130);
and U10399 (N_10399,N_10166,N_10140);
or U10400 (N_10400,N_9936,N_10010);
xnor U10401 (N_10401,N_10116,N_9965);
xor U10402 (N_10402,N_10050,N_9947);
nand U10403 (N_10403,N_10002,N_10013);
nor U10404 (N_10404,N_9926,N_10007);
or U10405 (N_10405,N_9920,N_9904);
nand U10406 (N_10406,N_9975,N_10040);
and U10407 (N_10407,N_10168,N_10158);
nand U10408 (N_10408,N_10039,N_10176);
nor U10409 (N_10409,N_10139,N_9923);
xor U10410 (N_10410,N_9983,N_10064);
and U10411 (N_10411,N_10189,N_10108);
nand U10412 (N_10412,N_10004,N_10186);
and U10413 (N_10413,N_9997,N_9917);
and U10414 (N_10414,N_9997,N_10184);
nor U10415 (N_10415,N_9960,N_10068);
nor U10416 (N_10416,N_9969,N_10123);
nor U10417 (N_10417,N_10090,N_10066);
nand U10418 (N_10418,N_10145,N_9912);
and U10419 (N_10419,N_10103,N_10183);
nand U10420 (N_10420,N_10057,N_9930);
or U10421 (N_10421,N_10034,N_10015);
and U10422 (N_10422,N_9968,N_10168);
nor U10423 (N_10423,N_10165,N_10044);
xor U10424 (N_10424,N_10081,N_10029);
and U10425 (N_10425,N_10184,N_10140);
xnor U10426 (N_10426,N_10039,N_10042);
and U10427 (N_10427,N_9923,N_9991);
or U10428 (N_10428,N_9913,N_10162);
and U10429 (N_10429,N_10189,N_9998);
or U10430 (N_10430,N_10026,N_10186);
nand U10431 (N_10431,N_10079,N_10049);
xor U10432 (N_10432,N_10142,N_10086);
xnor U10433 (N_10433,N_10025,N_10079);
xnor U10434 (N_10434,N_10077,N_9947);
or U10435 (N_10435,N_10149,N_9984);
xnor U10436 (N_10436,N_9943,N_10025);
nand U10437 (N_10437,N_9915,N_10121);
or U10438 (N_10438,N_10148,N_10035);
nand U10439 (N_10439,N_10142,N_10031);
nand U10440 (N_10440,N_10053,N_10083);
nor U10441 (N_10441,N_10143,N_10044);
and U10442 (N_10442,N_9929,N_10102);
and U10443 (N_10443,N_9946,N_9996);
and U10444 (N_10444,N_9999,N_9942);
and U10445 (N_10445,N_10042,N_10000);
nand U10446 (N_10446,N_9975,N_9918);
and U10447 (N_10447,N_10118,N_10177);
xor U10448 (N_10448,N_10039,N_10146);
and U10449 (N_10449,N_10157,N_9908);
and U10450 (N_10450,N_10025,N_10036);
xor U10451 (N_10451,N_10106,N_9977);
nand U10452 (N_10452,N_10092,N_10176);
nand U10453 (N_10453,N_10158,N_10004);
xor U10454 (N_10454,N_10059,N_9966);
or U10455 (N_10455,N_9922,N_10139);
nor U10456 (N_10456,N_10179,N_9935);
nand U10457 (N_10457,N_10046,N_10075);
and U10458 (N_10458,N_10045,N_10180);
and U10459 (N_10459,N_9918,N_10089);
and U10460 (N_10460,N_9900,N_9979);
and U10461 (N_10461,N_10149,N_9901);
or U10462 (N_10462,N_10009,N_10197);
or U10463 (N_10463,N_9940,N_10136);
and U10464 (N_10464,N_10031,N_10069);
nand U10465 (N_10465,N_10109,N_10026);
or U10466 (N_10466,N_10171,N_10056);
nand U10467 (N_10467,N_9980,N_10007);
and U10468 (N_10468,N_10198,N_10104);
and U10469 (N_10469,N_10084,N_10075);
nor U10470 (N_10470,N_10012,N_10029);
nand U10471 (N_10471,N_10122,N_9907);
xor U10472 (N_10472,N_9936,N_10149);
nor U10473 (N_10473,N_10061,N_10065);
or U10474 (N_10474,N_10147,N_9966);
and U10475 (N_10475,N_10155,N_10139);
nor U10476 (N_10476,N_9913,N_10001);
and U10477 (N_10477,N_9984,N_10002);
xor U10478 (N_10478,N_9988,N_9964);
or U10479 (N_10479,N_10154,N_9994);
nor U10480 (N_10480,N_10031,N_10106);
nand U10481 (N_10481,N_9991,N_9929);
nand U10482 (N_10482,N_9972,N_9978);
nor U10483 (N_10483,N_9948,N_10153);
nor U10484 (N_10484,N_9927,N_10012);
and U10485 (N_10485,N_9909,N_9912);
xor U10486 (N_10486,N_9913,N_10165);
and U10487 (N_10487,N_10143,N_10159);
nor U10488 (N_10488,N_9999,N_10004);
nand U10489 (N_10489,N_10199,N_10038);
xor U10490 (N_10490,N_9908,N_9946);
or U10491 (N_10491,N_10121,N_10077);
xnor U10492 (N_10492,N_10015,N_10178);
nand U10493 (N_10493,N_10112,N_10085);
and U10494 (N_10494,N_10071,N_10172);
and U10495 (N_10495,N_9945,N_9909);
or U10496 (N_10496,N_10193,N_10127);
and U10497 (N_10497,N_10107,N_10136);
xnor U10498 (N_10498,N_9925,N_9927);
nor U10499 (N_10499,N_9935,N_10082);
nand U10500 (N_10500,N_10303,N_10424);
or U10501 (N_10501,N_10436,N_10480);
and U10502 (N_10502,N_10333,N_10438);
nand U10503 (N_10503,N_10227,N_10340);
or U10504 (N_10504,N_10351,N_10223);
nor U10505 (N_10505,N_10263,N_10361);
nand U10506 (N_10506,N_10397,N_10426);
nor U10507 (N_10507,N_10413,N_10299);
nand U10508 (N_10508,N_10377,N_10238);
and U10509 (N_10509,N_10205,N_10217);
nor U10510 (N_10510,N_10250,N_10366);
and U10511 (N_10511,N_10326,N_10386);
nand U10512 (N_10512,N_10375,N_10401);
nor U10513 (N_10513,N_10433,N_10295);
nand U10514 (N_10514,N_10308,N_10497);
and U10515 (N_10515,N_10243,N_10364);
xor U10516 (N_10516,N_10395,N_10253);
nand U10517 (N_10517,N_10488,N_10210);
xor U10518 (N_10518,N_10249,N_10406);
xor U10519 (N_10519,N_10367,N_10486);
xor U10520 (N_10520,N_10272,N_10420);
and U10521 (N_10521,N_10264,N_10317);
and U10522 (N_10522,N_10437,N_10393);
nand U10523 (N_10523,N_10495,N_10476);
nand U10524 (N_10524,N_10347,N_10328);
and U10525 (N_10525,N_10311,N_10302);
or U10526 (N_10526,N_10468,N_10331);
nand U10527 (N_10527,N_10358,N_10493);
nand U10528 (N_10528,N_10465,N_10460);
and U10529 (N_10529,N_10434,N_10234);
nor U10530 (N_10530,N_10475,N_10415);
or U10531 (N_10531,N_10242,N_10284);
nor U10532 (N_10532,N_10481,N_10214);
nand U10533 (N_10533,N_10246,N_10298);
nand U10534 (N_10534,N_10384,N_10491);
nor U10535 (N_10535,N_10471,N_10289);
nor U10536 (N_10536,N_10320,N_10209);
nand U10537 (N_10537,N_10327,N_10484);
xor U10538 (N_10538,N_10266,N_10265);
or U10539 (N_10539,N_10279,N_10423);
and U10540 (N_10540,N_10292,N_10348);
xnor U10541 (N_10541,N_10408,N_10324);
and U10542 (N_10542,N_10342,N_10354);
or U10543 (N_10543,N_10306,N_10365);
and U10544 (N_10544,N_10483,N_10211);
or U10545 (N_10545,N_10430,N_10271);
nand U10546 (N_10546,N_10304,N_10280);
and U10547 (N_10547,N_10278,N_10204);
xor U10548 (N_10548,N_10498,N_10256);
xor U10549 (N_10549,N_10274,N_10441);
or U10550 (N_10550,N_10291,N_10203);
xor U10551 (N_10551,N_10370,N_10339);
nand U10552 (N_10552,N_10429,N_10477);
xnor U10553 (N_10553,N_10391,N_10411);
xor U10554 (N_10554,N_10276,N_10412);
or U10555 (N_10555,N_10363,N_10455);
or U10556 (N_10556,N_10494,N_10445);
and U10557 (N_10557,N_10452,N_10447);
nand U10558 (N_10558,N_10255,N_10432);
xor U10559 (N_10559,N_10442,N_10285);
nand U10560 (N_10560,N_10335,N_10334);
nor U10561 (N_10561,N_10296,N_10201);
nor U10562 (N_10562,N_10385,N_10294);
and U10563 (N_10563,N_10353,N_10282);
nand U10564 (N_10564,N_10257,N_10216);
and U10565 (N_10565,N_10245,N_10454);
and U10566 (N_10566,N_10208,N_10301);
nand U10567 (N_10567,N_10269,N_10372);
nand U10568 (N_10568,N_10376,N_10259);
nand U10569 (N_10569,N_10202,N_10275);
xnor U10570 (N_10570,N_10487,N_10207);
xor U10571 (N_10571,N_10337,N_10496);
or U10572 (N_10572,N_10458,N_10232);
nor U10573 (N_10573,N_10461,N_10261);
nand U10574 (N_10574,N_10312,N_10499);
and U10575 (N_10575,N_10383,N_10359);
xor U10576 (N_10576,N_10336,N_10389);
xor U10577 (N_10577,N_10319,N_10373);
nand U10578 (N_10578,N_10230,N_10360);
or U10579 (N_10579,N_10212,N_10262);
or U10580 (N_10580,N_10240,N_10407);
or U10581 (N_10581,N_10222,N_10310);
and U10582 (N_10582,N_10462,N_10231);
and U10583 (N_10583,N_10492,N_10220);
and U10584 (N_10584,N_10419,N_10396);
and U10585 (N_10585,N_10343,N_10346);
nand U10586 (N_10586,N_10405,N_10418);
nand U10587 (N_10587,N_10472,N_10307);
or U10588 (N_10588,N_10288,N_10239);
xor U10589 (N_10589,N_10247,N_10400);
xnor U10590 (N_10590,N_10435,N_10440);
and U10591 (N_10591,N_10425,N_10387);
nor U10592 (N_10592,N_10489,N_10305);
xnor U10593 (N_10593,N_10277,N_10382);
and U10594 (N_10594,N_10244,N_10235);
nor U10595 (N_10595,N_10381,N_10451);
nor U10596 (N_10596,N_10293,N_10226);
and U10597 (N_10597,N_10321,N_10218);
xor U10598 (N_10598,N_10273,N_10379);
nor U10599 (N_10599,N_10485,N_10478);
and U10600 (N_10600,N_10390,N_10267);
nor U10601 (N_10601,N_10341,N_10449);
xnor U10602 (N_10602,N_10374,N_10398);
nor U10603 (N_10603,N_10241,N_10332);
and U10604 (N_10604,N_10380,N_10228);
and U10605 (N_10605,N_10270,N_10268);
nand U10606 (N_10606,N_10251,N_10479);
or U10607 (N_10607,N_10446,N_10252);
and U10608 (N_10608,N_10428,N_10236);
xnor U10609 (N_10609,N_10421,N_10350);
nor U10610 (N_10610,N_10221,N_10469);
or U10611 (N_10611,N_10356,N_10219);
nor U10612 (N_10612,N_10330,N_10283);
xnor U10613 (N_10613,N_10399,N_10349);
and U10614 (N_10614,N_10431,N_10443);
nor U10615 (N_10615,N_10338,N_10416);
or U10616 (N_10616,N_10200,N_10345);
or U10617 (N_10617,N_10281,N_10388);
and U10618 (N_10618,N_10378,N_10286);
xor U10619 (N_10619,N_10409,N_10392);
nor U10620 (N_10620,N_10403,N_10402);
or U10621 (N_10621,N_10329,N_10344);
nor U10622 (N_10622,N_10422,N_10466);
nand U10623 (N_10623,N_10439,N_10224);
or U10624 (N_10624,N_10417,N_10323);
xnor U10625 (N_10625,N_10316,N_10362);
xnor U10626 (N_10626,N_10322,N_10233);
and U10627 (N_10627,N_10459,N_10450);
or U10628 (N_10628,N_10315,N_10325);
or U10629 (N_10629,N_10309,N_10394);
and U10630 (N_10630,N_10357,N_10404);
or U10631 (N_10631,N_10448,N_10248);
xnor U10632 (N_10632,N_10490,N_10287);
or U10633 (N_10633,N_10482,N_10225);
xnor U10634 (N_10634,N_10473,N_10213);
nand U10635 (N_10635,N_10474,N_10314);
nor U10636 (N_10636,N_10229,N_10410);
or U10637 (N_10637,N_10463,N_10352);
or U10638 (N_10638,N_10414,N_10444);
or U10639 (N_10639,N_10427,N_10456);
and U10640 (N_10640,N_10318,N_10300);
nor U10641 (N_10641,N_10297,N_10237);
or U10642 (N_10642,N_10371,N_10206);
nor U10643 (N_10643,N_10467,N_10260);
or U10644 (N_10644,N_10368,N_10464);
or U10645 (N_10645,N_10313,N_10453);
or U10646 (N_10646,N_10457,N_10290);
nor U10647 (N_10647,N_10470,N_10369);
xor U10648 (N_10648,N_10254,N_10215);
xnor U10649 (N_10649,N_10258,N_10355);
and U10650 (N_10650,N_10234,N_10396);
and U10651 (N_10651,N_10348,N_10373);
xor U10652 (N_10652,N_10201,N_10220);
or U10653 (N_10653,N_10360,N_10410);
xor U10654 (N_10654,N_10434,N_10408);
nand U10655 (N_10655,N_10274,N_10415);
or U10656 (N_10656,N_10414,N_10224);
or U10657 (N_10657,N_10317,N_10258);
nor U10658 (N_10658,N_10257,N_10375);
xnor U10659 (N_10659,N_10376,N_10454);
xnor U10660 (N_10660,N_10349,N_10393);
nor U10661 (N_10661,N_10208,N_10320);
nor U10662 (N_10662,N_10452,N_10256);
and U10663 (N_10663,N_10408,N_10497);
and U10664 (N_10664,N_10456,N_10477);
and U10665 (N_10665,N_10361,N_10261);
and U10666 (N_10666,N_10347,N_10287);
nand U10667 (N_10667,N_10397,N_10469);
xor U10668 (N_10668,N_10264,N_10484);
and U10669 (N_10669,N_10268,N_10280);
or U10670 (N_10670,N_10254,N_10373);
nand U10671 (N_10671,N_10224,N_10232);
nor U10672 (N_10672,N_10460,N_10276);
xnor U10673 (N_10673,N_10225,N_10322);
or U10674 (N_10674,N_10411,N_10474);
nor U10675 (N_10675,N_10478,N_10210);
nor U10676 (N_10676,N_10293,N_10437);
and U10677 (N_10677,N_10463,N_10495);
xnor U10678 (N_10678,N_10258,N_10487);
and U10679 (N_10679,N_10387,N_10353);
xor U10680 (N_10680,N_10208,N_10374);
and U10681 (N_10681,N_10291,N_10327);
xnor U10682 (N_10682,N_10329,N_10228);
xnor U10683 (N_10683,N_10339,N_10264);
xnor U10684 (N_10684,N_10301,N_10253);
xor U10685 (N_10685,N_10261,N_10322);
xor U10686 (N_10686,N_10373,N_10279);
nand U10687 (N_10687,N_10352,N_10435);
nor U10688 (N_10688,N_10200,N_10232);
nand U10689 (N_10689,N_10483,N_10280);
or U10690 (N_10690,N_10366,N_10388);
nor U10691 (N_10691,N_10229,N_10334);
or U10692 (N_10692,N_10401,N_10290);
nor U10693 (N_10693,N_10397,N_10320);
or U10694 (N_10694,N_10300,N_10490);
nor U10695 (N_10695,N_10364,N_10403);
or U10696 (N_10696,N_10358,N_10482);
nor U10697 (N_10697,N_10354,N_10420);
or U10698 (N_10698,N_10315,N_10200);
nor U10699 (N_10699,N_10491,N_10455);
or U10700 (N_10700,N_10233,N_10344);
xor U10701 (N_10701,N_10239,N_10447);
xnor U10702 (N_10702,N_10454,N_10203);
xor U10703 (N_10703,N_10442,N_10496);
nand U10704 (N_10704,N_10210,N_10377);
or U10705 (N_10705,N_10332,N_10296);
xor U10706 (N_10706,N_10246,N_10448);
nor U10707 (N_10707,N_10498,N_10476);
xor U10708 (N_10708,N_10345,N_10214);
nor U10709 (N_10709,N_10369,N_10326);
or U10710 (N_10710,N_10370,N_10245);
nor U10711 (N_10711,N_10391,N_10337);
or U10712 (N_10712,N_10431,N_10386);
nand U10713 (N_10713,N_10475,N_10279);
xnor U10714 (N_10714,N_10310,N_10350);
or U10715 (N_10715,N_10220,N_10277);
nor U10716 (N_10716,N_10238,N_10466);
or U10717 (N_10717,N_10228,N_10467);
nand U10718 (N_10718,N_10280,N_10284);
and U10719 (N_10719,N_10350,N_10497);
and U10720 (N_10720,N_10285,N_10228);
nand U10721 (N_10721,N_10427,N_10261);
nand U10722 (N_10722,N_10430,N_10466);
and U10723 (N_10723,N_10414,N_10303);
nand U10724 (N_10724,N_10337,N_10378);
or U10725 (N_10725,N_10209,N_10467);
nand U10726 (N_10726,N_10476,N_10367);
and U10727 (N_10727,N_10261,N_10370);
xnor U10728 (N_10728,N_10460,N_10352);
nor U10729 (N_10729,N_10245,N_10426);
nand U10730 (N_10730,N_10249,N_10234);
nand U10731 (N_10731,N_10304,N_10285);
or U10732 (N_10732,N_10349,N_10331);
nand U10733 (N_10733,N_10220,N_10325);
or U10734 (N_10734,N_10236,N_10355);
or U10735 (N_10735,N_10309,N_10427);
and U10736 (N_10736,N_10286,N_10477);
nand U10737 (N_10737,N_10225,N_10434);
nand U10738 (N_10738,N_10298,N_10398);
nor U10739 (N_10739,N_10385,N_10241);
or U10740 (N_10740,N_10448,N_10283);
xnor U10741 (N_10741,N_10335,N_10396);
and U10742 (N_10742,N_10489,N_10292);
nor U10743 (N_10743,N_10230,N_10248);
nand U10744 (N_10744,N_10467,N_10295);
nand U10745 (N_10745,N_10422,N_10401);
nand U10746 (N_10746,N_10327,N_10316);
nor U10747 (N_10747,N_10375,N_10403);
and U10748 (N_10748,N_10387,N_10465);
or U10749 (N_10749,N_10499,N_10390);
xnor U10750 (N_10750,N_10250,N_10206);
and U10751 (N_10751,N_10426,N_10438);
nand U10752 (N_10752,N_10210,N_10379);
xnor U10753 (N_10753,N_10382,N_10389);
nor U10754 (N_10754,N_10337,N_10463);
nand U10755 (N_10755,N_10357,N_10318);
xor U10756 (N_10756,N_10273,N_10272);
or U10757 (N_10757,N_10227,N_10264);
nor U10758 (N_10758,N_10351,N_10429);
xor U10759 (N_10759,N_10330,N_10484);
or U10760 (N_10760,N_10338,N_10481);
nand U10761 (N_10761,N_10345,N_10211);
xor U10762 (N_10762,N_10295,N_10257);
or U10763 (N_10763,N_10468,N_10435);
nor U10764 (N_10764,N_10499,N_10295);
or U10765 (N_10765,N_10253,N_10274);
and U10766 (N_10766,N_10497,N_10297);
nor U10767 (N_10767,N_10346,N_10331);
nor U10768 (N_10768,N_10301,N_10286);
xor U10769 (N_10769,N_10435,N_10464);
nor U10770 (N_10770,N_10456,N_10464);
nor U10771 (N_10771,N_10473,N_10406);
nand U10772 (N_10772,N_10291,N_10368);
or U10773 (N_10773,N_10416,N_10479);
nor U10774 (N_10774,N_10435,N_10279);
nand U10775 (N_10775,N_10406,N_10207);
xnor U10776 (N_10776,N_10356,N_10448);
xor U10777 (N_10777,N_10248,N_10262);
nor U10778 (N_10778,N_10216,N_10254);
nor U10779 (N_10779,N_10304,N_10467);
and U10780 (N_10780,N_10270,N_10234);
or U10781 (N_10781,N_10409,N_10256);
or U10782 (N_10782,N_10219,N_10229);
and U10783 (N_10783,N_10433,N_10291);
nor U10784 (N_10784,N_10305,N_10278);
and U10785 (N_10785,N_10477,N_10302);
or U10786 (N_10786,N_10489,N_10379);
xnor U10787 (N_10787,N_10389,N_10380);
and U10788 (N_10788,N_10499,N_10470);
or U10789 (N_10789,N_10261,N_10254);
nand U10790 (N_10790,N_10396,N_10394);
or U10791 (N_10791,N_10360,N_10222);
or U10792 (N_10792,N_10483,N_10399);
xnor U10793 (N_10793,N_10339,N_10348);
nand U10794 (N_10794,N_10301,N_10404);
nor U10795 (N_10795,N_10316,N_10307);
and U10796 (N_10796,N_10397,N_10355);
xnor U10797 (N_10797,N_10416,N_10265);
xor U10798 (N_10798,N_10232,N_10338);
or U10799 (N_10799,N_10258,N_10210);
or U10800 (N_10800,N_10601,N_10512);
nand U10801 (N_10801,N_10617,N_10578);
nand U10802 (N_10802,N_10638,N_10781);
nand U10803 (N_10803,N_10670,N_10634);
nor U10804 (N_10804,N_10725,N_10550);
nand U10805 (N_10805,N_10700,N_10795);
nor U10806 (N_10806,N_10783,N_10789);
xnor U10807 (N_10807,N_10716,N_10561);
nor U10808 (N_10808,N_10664,N_10787);
nand U10809 (N_10809,N_10508,N_10694);
nor U10810 (N_10810,N_10542,N_10671);
xnor U10811 (N_10811,N_10654,N_10657);
and U10812 (N_10812,N_10524,N_10636);
nor U10813 (N_10813,N_10730,N_10616);
nor U10814 (N_10814,N_10685,N_10751);
or U10815 (N_10815,N_10754,N_10621);
nor U10816 (N_10816,N_10585,N_10701);
or U10817 (N_10817,N_10529,N_10790);
xor U10818 (N_10818,N_10662,N_10572);
nand U10819 (N_10819,N_10780,N_10603);
nand U10820 (N_10820,N_10687,N_10568);
nor U10821 (N_10821,N_10506,N_10732);
nor U10822 (N_10822,N_10703,N_10676);
nor U10823 (N_10823,N_10784,N_10788);
nand U10824 (N_10824,N_10673,N_10643);
nand U10825 (N_10825,N_10760,N_10768);
and U10826 (N_10826,N_10628,N_10773);
nand U10827 (N_10827,N_10510,N_10635);
nor U10828 (N_10828,N_10766,N_10543);
or U10829 (N_10829,N_10520,N_10573);
nor U10830 (N_10830,N_10772,N_10624);
or U10831 (N_10831,N_10755,N_10713);
or U10832 (N_10832,N_10516,N_10569);
or U10833 (N_10833,N_10614,N_10746);
nor U10834 (N_10834,N_10762,N_10731);
and U10835 (N_10835,N_10600,N_10689);
xnor U10836 (N_10836,N_10799,N_10544);
xor U10837 (N_10837,N_10686,N_10672);
nor U10838 (N_10838,N_10593,N_10753);
and U10839 (N_10839,N_10525,N_10656);
and U10840 (N_10840,N_10574,N_10668);
nand U10841 (N_10841,N_10534,N_10774);
or U10842 (N_10842,N_10692,N_10717);
nand U10843 (N_10843,N_10591,N_10677);
and U10844 (N_10844,N_10737,N_10769);
or U10845 (N_10845,N_10604,N_10555);
xor U10846 (N_10846,N_10798,N_10632);
nand U10847 (N_10847,N_10528,N_10791);
xnor U10848 (N_10848,N_10583,N_10786);
and U10849 (N_10849,N_10704,N_10549);
xor U10850 (N_10850,N_10579,N_10666);
or U10851 (N_10851,N_10539,N_10580);
and U10852 (N_10852,N_10698,N_10563);
xor U10853 (N_10853,N_10536,N_10642);
xor U10854 (N_10854,N_10699,N_10681);
and U10855 (N_10855,N_10719,N_10546);
xnor U10856 (N_10856,N_10721,N_10782);
or U10857 (N_10857,N_10641,N_10586);
nor U10858 (N_10858,N_10674,N_10581);
or U10859 (N_10859,N_10532,N_10619);
nor U10860 (N_10860,N_10625,N_10533);
xor U10861 (N_10861,N_10639,N_10503);
xor U10862 (N_10862,N_10712,N_10658);
or U10863 (N_10863,N_10738,N_10776);
nor U10864 (N_10864,N_10566,N_10705);
and U10865 (N_10865,N_10763,N_10556);
and U10866 (N_10866,N_10767,N_10661);
nor U10867 (N_10867,N_10584,N_10599);
nor U10868 (N_10868,N_10627,N_10582);
and U10869 (N_10869,N_10640,N_10631);
or U10870 (N_10870,N_10551,N_10607);
or U10871 (N_10871,N_10511,N_10722);
and U10872 (N_10872,N_10613,N_10683);
nor U10873 (N_10873,N_10560,N_10757);
nor U10874 (N_10874,N_10761,N_10709);
nor U10875 (N_10875,N_10559,N_10541);
xor U10876 (N_10876,N_10736,N_10710);
nand U10877 (N_10877,N_10605,N_10502);
nor U10878 (N_10878,N_10562,N_10535);
nand U10879 (N_10879,N_10548,N_10606);
nor U10880 (N_10880,N_10720,N_10519);
nor U10881 (N_10881,N_10759,N_10655);
or U10882 (N_10882,N_10598,N_10558);
or U10883 (N_10883,N_10660,N_10618);
or U10884 (N_10884,N_10505,N_10623);
and U10885 (N_10885,N_10513,N_10734);
xnor U10886 (N_10886,N_10595,N_10779);
xnor U10887 (N_10887,N_10708,N_10567);
xor U10888 (N_10888,N_10575,N_10530);
or U10889 (N_10889,N_10626,N_10526);
and U10890 (N_10890,N_10696,N_10514);
xnor U10891 (N_10891,N_10500,N_10679);
nor U10892 (N_10892,N_10590,N_10596);
and U10893 (N_10893,N_10770,N_10777);
nor U10894 (N_10894,N_10684,N_10715);
xnor U10895 (N_10895,N_10758,N_10680);
xnor U10896 (N_10896,N_10577,N_10729);
nor U10897 (N_10897,N_10538,N_10748);
nand U10898 (N_10898,N_10501,N_10747);
and U10899 (N_10899,N_10678,N_10735);
and U10900 (N_10900,N_10650,N_10794);
nand U10901 (N_10901,N_10608,N_10706);
xnor U10902 (N_10902,N_10570,N_10764);
and U10903 (N_10903,N_10507,N_10714);
or U10904 (N_10904,N_10775,N_10665);
and U10905 (N_10905,N_10540,N_10765);
xnor U10906 (N_10906,N_10504,N_10521);
nor U10907 (N_10907,N_10518,N_10695);
or U10908 (N_10908,N_10545,N_10653);
or U10909 (N_10909,N_10647,N_10745);
xnor U10910 (N_10910,N_10644,N_10771);
and U10911 (N_10911,N_10744,N_10565);
or U10912 (N_10912,N_10523,N_10645);
xor U10913 (N_10913,N_10515,N_10597);
xnor U10914 (N_10914,N_10724,N_10630);
xor U10915 (N_10915,N_10742,N_10756);
xor U10916 (N_10916,N_10651,N_10537);
xor U10917 (N_10917,N_10554,N_10589);
nand U10918 (N_10918,N_10707,N_10609);
nand U10919 (N_10919,N_10741,N_10527);
xor U10920 (N_10920,N_10594,N_10667);
xnor U10921 (N_10921,N_10693,N_10612);
nor U10922 (N_10922,N_10509,N_10793);
nor U10923 (N_10923,N_10531,N_10792);
nor U10924 (N_10924,N_10785,N_10592);
nor U10925 (N_10925,N_10588,N_10669);
nor U10926 (N_10926,N_10675,N_10726);
or U10927 (N_10927,N_10522,N_10663);
xor U10928 (N_10928,N_10739,N_10571);
nand U10929 (N_10929,N_10576,N_10727);
nor U10930 (N_10930,N_10796,N_10652);
xor U10931 (N_10931,N_10564,N_10688);
xnor U10932 (N_10932,N_10691,N_10547);
or U10933 (N_10933,N_10723,N_10690);
and U10934 (N_10934,N_10749,N_10648);
nor U10935 (N_10935,N_10646,N_10610);
nor U10936 (N_10936,N_10517,N_10728);
or U10937 (N_10937,N_10697,N_10649);
xnor U10938 (N_10938,N_10620,N_10633);
xnor U10939 (N_10939,N_10629,N_10740);
or U10940 (N_10940,N_10553,N_10750);
xnor U10941 (N_10941,N_10797,N_10733);
nand U10942 (N_10942,N_10778,N_10743);
and U10943 (N_10943,N_10557,N_10682);
xnor U10944 (N_10944,N_10711,N_10552);
xnor U10945 (N_10945,N_10615,N_10637);
xor U10946 (N_10946,N_10622,N_10587);
or U10947 (N_10947,N_10602,N_10659);
and U10948 (N_10948,N_10752,N_10718);
xnor U10949 (N_10949,N_10611,N_10702);
nor U10950 (N_10950,N_10702,N_10537);
xor U10951 (N_10951,N_10709,N_10690);
or U10952 (N_10952,N_10717,N_10660);
or U10953 (N_10953,N_10754,N_10581);
nor U10954 (N_10954,N_10537,N_10631);
xnor U10955 (N_10955,N_10733,N_10738);
nand U10956 (N_10956,N_10606,N_10776);
and U10957 (N_10957,N_10593,N_10668);
or U10958 (N_10958,N_10777,N_10654);
xnor U10959 (N_10959,N_10625,N_10656);
or U10960 (N_10960,N_10739,N_10672);
xnor U10961 (N_10961,N_10687,N_10721);
or U10962 (N_10962,N_10685,N_10580);
nor U10963 (N_10963,N_10661,N_10630);
xnor U10964 (N_10964,N_10777,N_10577);
or U10965 (N_10965,N_10653,N_10541);
or U10966 (N_10966,N_10574,N_10638);
or U10967 (N_10967,N_10502,N_10790);
nor U10968 (N_10968,N_10568,N_10709);
or U10969 (N_10969,N_10561,N_10677);
or U10970 (N_10970,N_10633,N_10674);
and U10971 (N_10971,N_10772,N_10682);
and U10972 (N_10972,N_10730,N_10505);
nand U10973 (N_10973,N_10582,N_10737);
nand U10974 (N_10974,N_10664,N_10700);
nor U10975 (N_10975,N_10626,N_10620);
or U10976 (N_10976,N_10633,N_10658);
nor U10977 (N_10977,N_10690,N_10516);
and U10978 (N_10978,N_10799,N_10562);
or U10979 (N_10979,N_10552,N_10728);
nor U10980 (N_10980,N_10516,N_10715);
nand U10981 (N_10981,N_10728,N_10590);
nor U10982 (N_10982,N_10729,N_10512);
nor U10983 (N_10983,N_10717,N_10597);
nand U10984 (N_10984,N_10576,N_10507);
xnor U10985 (N_10985,N_10621,N_10515);
nand U10986 (N_10986,N_10766,N_10637);
xnor U10987 (N_10987,N_10555,N_10663);
and U10988 (N_10988,N_10613,N_10545);
nor U10989 (N_10989,N_10533,N_10676);
nand U10990 (N_10990,N_10559,N_10554);
nor U10991 (N_10991,N_10694,N_10594);
or U10992 (N_10992,N_10716,N_10772);
or U10993 (N_10993,N_10673,N_10584);
or U10994 (N_10994,N_10558,N_10573);
xor U10995 (N_10995,N_10763,N_10696);
nand U10996 (N_10996,N_10685,N_10764);
and U10997 (N_10997,N_10784,N_10765);
nand U10998 (N_10998,N_10778,N_10626);
xor U10999 (N_10999,N_10744,N_10595);
or U11000 (N_11000,N_10724,N_10552);
nand U11001 (N_11001,N_10799,N_10677);
xnor U11002 (N_11002,N_10743,N_10610);
xnor U11003 (N_11003,N_10770,N_10761);
nand U11004 (N_11004,N_10631,N_10673);
nand U11005 (N_11005,N_10687,N_10703);
nand U11006 (N_11006,N_10621,N_10774);
or U11007 (N_11007,N_10696,N_10624);
and U11008 (N_11008,N_10514,N_10706);
or U11009 (N_11009,N_10616,N_10555);
and U11010 (N_11010,N_10559,N_10715);
and U11011 (N_11011,N_10767,N_10656);
and U11012 (N_11012,N_10503,N_10622);
and U11013 (N_11013,N_10635,N_10568);
or U11014 (N_11014,N_10717,N_10764);
nor U11015 (N_11015,N_10687,N_10728);
nand U11016 (N_11016,N_10582,N_10566);
xor U11017 (N_11017,N_10772,N_10751);
and U11018 (N_11018,N_10778,N_10578);
nor U11019 (N_11019,N_10584,N_10651);
xor U11020 (N_11020,N_10647,N_10747);
xnor U11021 (N_11021,N_10729,N_10667);
xor U11022 (N_11022,N_10771,N_10788);
nand U11023 (N_11023,N_10650,N_10567);
nand U11024 (N_11024,N_10561,N_10549);
and U11025 (N_11025,N_10719,N_10532);
xor U11026 (N_11026,N_10580,N_10724);
nor U11027 (N_11027,N_10647,N_10553);
and U11028 (N_11028,N_10568,N_10534);
xnor U11029 (N_11029,N_10640,N_10612);
and U11030 (N_11030,N_10645,N_10504);
nand U11031 (N_11031,N_10536,N_10554);
or U11032 (N_11032,N_10702,N_10726);
nor U11033 (N_11033,N_10796,N_10560);
nor U11034 (N_11034,N_10578,N_10576);
or U11035 (N_11035,N_10595,N_10616);
nor U11036 (N_11036,N_10622,N_10525);
and U11037 (N_11037,N_10601,N_10552);
nand U11038 (N_11038,N_10740,N_10605);
xor U11039 (N_11039,N_10578,N_10732);
and U11040 (N_11040,N_10602,N_10761);
xor U11041 (N_11041,N_10503,N_10509);
nor U11042 (N_11042,N_10744,N_10773);
nor U11043 (N_11043,N_10773,N_10784);
nor U11044 (N_11044,N_10644,N_10743);
and U11045 (N_11045,N_10660,N_10666);
nor U11046 (N_11046,N_10580,N_10747);
and U11047 (N_11047,N_10528,N_10696);
nand U11048 (N_11048,N_10778,N_10560);
nand U11049 (N_11049,N_10531,N_10621);
xnor U11050 (N_11050,N_10722,N_10586);
xnor U11051 (N_11051,N_10628,N_10582);
or U11052 (N_11052,N_10595,N_10617);
nor U11053 (N_11053,N_10536,N_10572);
xor U11054 (N_11054,N_10591,N_10623);
nor U11055 (N_11055,N_10639,N_10686);
xor U11056 (N_11056,N_10634,N_10608);
or U11057 (N_11057,N_10734,N_10777);
nor U11058 (N_11058,N_10790,N_10739);
or U11059 (N_11059,N_10672,N_10653);
nor U11060 (N_11060,N_10732,N_10757);
and U11061 (N_11061,N_10541,N_10683);
and U11062 (N_11062,N_10604,N_10527);
and U11063 (N_11063,N_10697,N_10576);
nor U11064 (N_11064,N_10542,N_10714);
or U11065 (N_11065,N_10527,N_10730);
nor U11066 (N_11066,N_10794,N_10731);
and U11067 (N_11067,N_10557,N_10630);
and U11068 (N_11068,N_10709,N_10528);
nor U11069 (N_11069,N_10722,N_10555);
and U11070 (N_11070,N_10608,N_10541);
xnor U11071 (N_11071,N_10797,N_10562);
or U11072 (N_11072,N_10656,N_10711);
nor U11073 (N_11073,N_10507,N_10515);
nand U11074 (N_11074,N_10575,N_10686);
xor U11075 (N_11075,N_10709,N_10743);
xor U11076 (N_11076,N_10683,N_10655);
or U11077 (N_11077,N_10712,N_10651);
or U11078 (N_11078,N_10547,N_10701);
nand U11079 (N_11079,N_10599,N_10717);
nor U11080 (N_11080,N_10558,N_10632);
nand U11081 (N_11081,N_10644,N_10724);
and U11082 (N_11082,N_10583,N_10721);
xor U11083 (N_11083,N_10745,N_10760);
xor U11084 (N_11084,N_10762,N_10654);
nand U11085 (N_11085,N_10779,N_10695);
nand U11086 (N_11086,N_10560,N_10719);
nor U11087 (N_11087,N_10798,N_10731);
nand U11088 (N_11088,N_10510,N_10567);
nand U11089 (N_11089,N_10596,N_10562);
xnor U11090 (N_11090,N_10788,N_10603);
xor U11091 (N_11091,N_10523,N_10751);
and U11092 (N_11092,N_10720,N_10504);
nand U11093 (N_11093,N_10527,N_10556);
or U11094 (N_11094,N_10506,N_10659);
nor U11095 (N_11095,N_10578,N_10669);
nor U11096 (N_11096,N_10798,N_10655);
nand U11097 (N_11097,N_10533,N_10762);
or U11098 (N_11098,N_10531,N_10514);
xor U11099 (N_11099,N_10678,N_10616);
or U11100 (N_11100,N_10916,N_10981);
and U11101 (N_11101,N_10811,N_10861);
and U11102 (N_11102,N_11068,N_10915);
nand U11103 (N_11103,N_10883,N_11017);
and U11104 (N_11104,N_10887,N_11008);
xnor U11105 (N_11105,N_10991,N_10843);
nor U11106 (N_11106,N_10825,N_10923);
and U11107 (N_11107,N_10891,N_11084);
and U11108 (N_11108,N_10815,N_10902);
nor U11109 (N_11109,N_11056,N_10855);
nand U11110 (N_11110,N_10820,N_10876);
xor U11111 (N_11111,N_10961,N_10993);
or U11112 (N_11112,N_10997,N_10865);
nand U11113 (N_11113,N_10808,N_10879);
or U11114 (N_11114,N_10945,N_10839);
or U11115 (N_11115,N_10932,N_10833);
and U11116 (N_11116,N_10985,N_11064);
and U11117 (N_11117,N_10996,N_10901);
xnor U11118 (N_11118,N_11024,N_10920);
xor U11119 (N_11119,N_10957,N_10826);
nand U11120 (N_11120,N_10877,N_11065);
nor U11121 (N_11121,N_11041,N_11040);
nor U11122 (N_11122,N_10999,N_10832);
nor U11123 (N_11123,N_10908,N_10804);
or U11124 (N_11124,N_10805,N_10994);
nor U11125 (N_11125,N_10852,N_10869);
nor U11126 (N_11126,N_10892,N_10988);
xnor U11127 (N_11127,N_11057,N_10885);
xor U11128 (N_11128,N_10821,N_11009);
or U11129 (N_11129,N_11067,N_10922);
xor U11130 (N_11130,N_11020,N_10914);
nor U11131 (N_11131,N_11082,N_10943);
or U11132 (N_11132,N_10950,N_10859);
nand U11133 (N_11133,N_10851,N_10810);
nand U11134 (N_11134,N_10886,N_10871);
nand U11135 (N_11135,N_10936,N_10881);
xnor U11136 (N_11136,N_10980,N_11078);
xnor U11137 (N_11137,N_11058,N_10975);
nor U11138 (N_11138,N_10840,N_10873);
xnor U11139 (N_11139,N_11060,N_11001);
nand U11140 (N_11140,N_10953,N_10949);
nor U11141 (N_11141,N_11021,N_10866);
and U11142 (N_11142,N_10857,N_10965);
and U11143 (N_11143,N_11039,N_10894);
or U11144 (N_11144,N_10824,N_10806);
xnor U11145 (N_11145,N_10960,N_11051);
and U11146 (N_11146,N_10927,N_10946);
nand U11147 (N_11147,N_11032,N_10924);
xor U11148 (N_11148,N_10982,N_11034);
xor U11149 (N_11149,N_10983,N_10802);
nor U11150 (N_11150,N_10850,N_10942);
and U11151 (N_11151,N_10933,N_10974);
xnor U11152 (N_11152,N_11049,N_11069);
nand U11153 (N_11153,N_10801,N_11016);
nor U11154 (N_11154,N_10962,N_10870);
and U11155 (N_11155,N_10921,N_10926);
and U11156 (N_11156,N_10958,N_10992);
and U11157 (N_11157,N_11014,N_11003);
nand U11158 (N_11158,N_11022,N_10978);
and U11159 (N_11159,N_10903,N_11050);
nor U11160 (N_11160,N_10919,N_10998);
and U11161 (N_11161,N_11086,N_11000);
and U11162 (N_11162,N_10846,N_11096);
xnor U11163 (N_11163,N_10973,N_10912);
or U11164 (N_11164,N_11010,N_10911);
and U11165 (N_11165,N_10847,N_10835);
xnor U11166 (N_11166,N_11002,N_10809);
nor U11167 (N_11167,N_10858,N_10955);
nand U11168 (N_11168,N_11079,N_11018);
xnor U11169 (N_11169,N_10899,N_10929);
and U11170 (N_11170,N_11070,N_11011);
or U11171 (N_11171,N_10952,N_10812);
xor U11172 (N_11172,N_10979,N_11093);
and U11173 (N_11173,N_10934,N_10947);
nand U11174 (N_11174,N_11053,N_10963);
and U11175 (N_11175,N_10854,N_10937);
or U11176 (N_11176,N_10906,N_11026);
nand U11177 (N_11177,N_11019,N_11047);
nand U11178 (N_11178,N_10918,N_10853);
or U11179 (N_11179,N_10890,N_11013);
and U11180 (N_11180,N_10928,N_10990);
nand U11181 (N_11181,N_11087,N_10956);
nand U11182 (N_11182,N_10909,N_10941);
nand U11183 (N_11183,N_10989,N_10807);
and U11184 (N_11184,N_10818,N_11007);
and U11185 (N_11185,N_11029,N_10848);
xor U11186 (N_11186,N_11077,N_10837);
xor U11187 (N_11187,N_11035,N_10828);
nand U11188 (N_11188,N_11031,N_10842);
xor U11189 (N_11189,N_11094,N_10910);
or U11190 (N_11190,N_11015,N_10800);
xor U11191 (N_11191,N_10913,N_11042);
nand U11192 (N_11192,N_11052,N_10863);
nor U11193 (N_11193,N_11097,N_10875);
and U11194 (N_11194,N_11037,N_10813);
and U11195 (N_11195,N_10972,N_10856);
xor U11196 (N_11196,N_11089,N_10954);
xor U11197 (N_11197,N_11048,N_11038);
or U11198 (N_11198,N_10867,N_11095);
nand U11199 (N_11199,N_11005,N_11054);
or U11200 (N_11200,N_10904,N_10951);
xor U11201 (N_11201,N_11090,N_10938);
nand U11202 (N_11202,N_10905,N_10930);
and U11203 (N_11203,N_11045,N_11092);
xnor U11204 (N_11204,N_10829,N_11075);
and U11205 (N_11205,N_10836,N_10864);
or U11206 (N_11206,N_10872,N_10888);
nand U11207 (N_11207,N_10900,N_11081);
nor U11208 (N_11208,N_10984,N_10971);
nor U11209 (N_11209,N_11055,N_10862);
nor U11210 (N_11210,N_11046,N_11027);
and U11211 (N_11211,N_11063,N_10976);
nor U11212 (N_11212,N_10931,N_11099);
or U11213 (N_11213,N_10935,N_11083);
nand U11214 (N_11214,N_10898,N_10831);
xnor U11215 (N_11215,N_10917,N_10970);
or U11216 (N_11216,N_10860,N_10893);
nand U11217 (N_11217,N_10816,N_10884);
xor U11218 (N_11218,N_11036,N_10896);
or U11219 (N_11219,N_11028,N_11071);
nor U11220 (N_11220,N_11043,N_11030);
and U11221 (N_11221,N_11085,N_10830);
nand U11222 (N_11222,N_10967,N_10925);
or U11223 (N_11223,N_11076,N_11006);
nor U11224 (N_11224,N_10814,N_11012);
nand U11225 (N_11225,N_10838,N_10822);
xnor U11226 (N_11226,N_10880,N_10907);
nor U11227 (N_11227,N_10966,N_10895);
and U11228 (N_11228,N_10969,N_10986);
nor U11229 (N_11229,N_10968,N_11044);
and U11230 (N_11230,N_10897,N_10841);
nor U11231 (N_11231,N_11073,N_10987);
xor U11232 (N_11232,N_10889,N_11074);
xor U11233 (N_11233,N_10817,N_10803);
nand U11234 (N_11234,N_10849,N_11004);
nand U11235 (N_11235,N_11098,N_10874);
or U11236 (N_11236,N_10939,N_11033);
nor U11237 (N_11237,N_11072,N_11088);
xnor U11238 (N_11238,N_10940,N_11080);
nand U11239 (N_11239,N_10819,N_11061);
nand U11240 (N_11240,N_11059,N_10977);
nor U11241 (N_11241,N_11091,N_11023);
nand U11242 (N_11242,N_10959,N_10868);
xnor U11243 (N_11243,N_10944,N_10823);
nand U11244 (N_11244,N_10834,N_10878);
nor U11245 (N_11245,N_10845,N_10882);
nor U11246 (N_11246,N_10844,N_10995);
nor U11247 (N_11247,N_11025,N_10827);
or U11248 (N_11248,N_10948,N_10964);
or U11249 (N_11249,N_11062,N_11066);
nor U11250 (N_11250,N_11074,N_10929);
nor U11251 (N_11251,N_10815,N_11079);
and U11252 (N_11252,N_10897,N_10929);
xor U11253 (N_11253,N_10821,N_10974);
nand U11254 (N_11254,N_10927,N_10884);
nor U11255 (N_11255,N_10824,N_10825);
and U11256 (N_11256,N_11031,N_10919);
or U11257 (N_11257,N_10892,N_10938);
and U11258 (N_11258,N_11065,N_10961);
xor U11259 (N_11259,N_10994,N_11089);
and U11260 (N_11260,N_10871,N_10852);
or U11261 (N_11261,N_10899,N_11025);
xnor U11262 (N_11262,N_10816,N_10983);
nand U11263 (N_11263,N_10819,N_11055);
nor U11264 (N_11264,N_10954,N_10872);
or U11265 (N_11265,N_11035,N_11098);
and U11266 (N_11266,N_10991,N_11000);
nand U11267 (N_11267,N_11091,N_10978);
nand U11268 (N_11268,N_10898,N_11081);
nand U11269 (N_11269,N_10800,N_10993);
nor U11270 (N_11270,N_10838,N_10848);
nand U11271 (N_11271,N_11041,N_10869);
and U11272 (N_11272,N_11037,N_10896);
and U11273 (N_11273,N_11056,N_11070);
nor U11274 (N_11274,N_11072,N_10911);
or U11275 (N_11275,N_10800,N_11082);
and U11276 (N_11276,N_10900,N_11088);
nand U11277 (N_11277,N_10986,N_10833);
or U11278 (N_11278,N_10911,N_11007);
and U11279 (N_11279,N_10906,N_10806);
nor U11280 (N_11280,N_11093,N_11004);
or U11281 (N_11281,N_10934,N_11086);
xor U11282 (N_11282,N_10905,N_10876);
xnor U11283 (N_11283,N_10824,N_10907);
or U11284 (N_11284,N_10980,N_10888);
or U11285 (N_11285,N_11075,N_10974);
xor U11286 (N_11286,N_10869,N_10981);
nor U11287 (N_11287,N_10907,N_10834);
nor U11288 (N_11288,N_10899,N_10871);
nor U11289 (N_11289,N_11041,N_10913);
and U11290 (N_11290,N_11075,N_11076);
nor U11291 (N_11291,N_10846,N_11063);
nor U11292 (N_11292,N_10976,N_10982);
or U11293 (N_11293,N_10866,N_10918);
nand U11294 (N_11294,N_10832,N_11006);
nand U11295 (N_11295,N_10937,N_10835);
xor U11296 (N_11296,N_10853,N_10878);
and U11297 (N_11297,N_10826,N_10883);
and U11298 (N_11298,N_11072,N_10880);
nand U11299 (N_11299,N_11087,N_11035);
xor U11300 (N_11300,N_11066,N_10999);
and U11301 (N_11301,N_11013,N_10908);
and U11302 (N_11302,N_10931,N_10966);
xor U11303 (N_11303,N_10866,N_11030);
nand U11304 (N_11304,N_10908,N_11090);
nand U11305 (N_11305,N_10866,N_10919);
or U11306 (N_11306,N_10986,N_10967);
and U11307 (N_11307,N_11055,N_10844);
xnor U11308 (N_11308,N_11035,N_10915);
xor U11309 (N_11309,N_10899,N_10864);
and U11310 (N_11310,N_11007,N_10897);
or U11311 (N_11311,N_10853,N_10987);
xnor U11312 (N_11312,N_10967,N_10929);
xor U11313 (N_11313,N_10964,N_11069);
nor U11314 (N_11314,N_11026,N_10832);
nand U11315 (N_11315,N_11043,N_10874);
and U11316 (N_11316,N_10829,N_10882);
xor U11317 (N_11317,N_11078,N_10944);
nand U11318 (N_11318,N_11083,N_10863);
nor U11319 (N_11319,N_10951,N_11097);
xnor U11320 (N_11320,N_10968,N_10816);
or U11321 (N_11321,N_11026,N_10990);
xnor U11322 (N_11322,N_11066,N_11052);
or U11323 (N_11323,N_10826,N_10815);
or U11324 (N_11324,N_10885,N_10938);
and U11325 (N_11325,N_10852,N_10864);
nor U11326 (N_11326,N_10825,N_10888);
nor U11327 (N_11327,N_11056,N_10804);
and U11328 (N_11328,N_10856,N_10890);
nand U11329 (N_11329,N_10941,N_10976);
xnor U11330 (N_11330,N_10952,N_10894);
or U11331 (N_11331,N_10952,N_11075);
nor U11332 (N_11332,N_10902,N_10908);
and U11333 (N_11333,N_10952,N_10921);
and U11334 (N_11334,N_10936,N_10968);
nor U11335 (N_11335,N_11022,N_11097);
and U11336 (N_11336,N_11053,N_10909);
or U11337 (N_11337,N_10928,N_10997);
nor U11338 (N_11338,N_11031,N_10851);
and U11339 (N_11339,N_10835,N_11088);
or U11340 (N_11340,N_11079,N_10996);
xor U11341 (N_11341,N_11014,N_11051);
xnor U11342 (N_11342,N_10943,N_10900);
xnor U11343 (N_11343,N_10930,N_10827);
nand U11344 (N_11344,N_10904,N_10891);
xnor U11345 (N_11345,N_10904,N_11005);
nand U11346 (N_11346,N_10948,N_10835);
nand U11347 (N_11347,N_10983,N_10870);
or U11348 (N_11348,N_11046,N_10970);
or U11349 (N_11349,N_10950,N_11074);
nand U11350 (N_11350,N_10852,N_10982);
or U11351 (N_11351,N_10832,N_10926);
and U11352 (N_11352,N_11044,N_10800);
and U11353 (N_11353,N_11077,N_11033);
and U11354 (N_11354,N_11079,N_11031);
xnor U11355 (N_11355,N_10897,N_11060);
nor U11356 (N_11356,N_11043,N_11072);
nor U11357 (N_11357,N_11051,N_10993);
and U11358 (N_11358,N_11051,N_11052);
nand U11359 (N_11359,N_10994,N_11065);
nand U11360 (N_11360,N_10986,N_10895);
nand U11361 (N_11361,N_10884,N_10873);
or U11362 (N_11362,N_10853,N_10938);
nor U11363 (N_11363,N_10906,N_11098);
xnor U11364 (N_11364,N_11089,N_10984);
or U11365 (N_11365,N_10810,N_10992);
nand U11366 (N_11366,N_10862,N_10839);
nor U11367 (N_11367,N_10841,N_10807);
or U11368 (N_11368,N_11026,N_11054);
nand U11369 (N_11369,N_10869,N_10904);
xnor U11370 (N_11370,N_10814,N_10943);
nand U11371 (N_11371,N_10931,N_11011);
or U11372 (N_11372,N_11044,N_10975);
nor U11373 (N_11373,N_10840,N_11030);
nand U11374 (N_11374,N_10851,N_11018);
xnor U11375 (N_11375,N_11079,N_10941);
xnor U11376 (N_11376,N_10808,N_10913);
nor U11377 (N_11377,N_11028,N_10938);
and U11378 (N_11378,N_10996,N_10887);
or U11379 (N_11379,N_10967,N_11090);
or U11380 (N_11380,N_11042,N_11094);
nand U11381 (N_11381,N_10828,N_11056);
xnor U11382 (N_11382,N_10835,N_11094);
nor U11383 (N_11383,N_10950,N_10999);
nor U11384 (N_11384,N_11093,N_10948);
or U11385 (N_11385,N_11036,N_10960);
or U11386 (N_11386,N_10802,N_10822);
nor U11387 (N_11387,N_10800,N_10847);
xor U11388 (N_11388,N_10926,N_11092);
xor U11389 (N_11389,N_10908,N_10977);
nand U11390 (N_11390,N_10808,N_10996);
nand U11391 (N_11391,N_11060,N_11015);
xnor U11392 (N_11392,N_11043,N_11011);
and U11393 (N_11393,N_10890,N_10937);
xor U11394 (N_11394,N_10910,N_11034);
xor U11395 (N_11395,N_10924,N_11017);
and U11396 (N_11396,N_10801,N_11004);
xnor U11397 (N_11397,N_11019,N_10837);
and U11398 (N_11398,N_10925,N_10982);
or U11399 (N_11399,N_11040,N_10970);
and U11400 (N_11400,N_11225,N_11238);
nor U11401 (N_11401,N_11334,N_11189);
or U11402 (N_11402,N_11184,N_11342);
or U11403 (N_11403,N_11383,N_11289);
nand U11404 (N_11404,N_11192,N_11395);
or U11405 (N_11405,N_11309,N_11257);
nand U11406 (N_11406,N_11267,N_11252);
xnor U11407 (N_11407,N_11349,N_11165);
xnor U11408 (N_11408,N_11206,N_11320);
or U11409 (N_11409,N_11319,N_11374);
nor U11410 (N_11410,N_11261,N_11325);
nand U11411 (N_11411,N_11333,N_11392);
or U11412 (N_11412,N_11195,N_11211);
nor U11413 (N_11413,N_11306,N_11317);
nor U11414 (N_11414,N_11258,N_11324);
xor U11415 (N_11415,N_11230,N_11336);
nand U11416 (N_11416,N_11203,N_11265);
or U11417 (N_11417,N_11284,N_11399);
or U11418 (N_11418,N_11312,N_11108);
nor U11419 (N_11419,N_11326,N_11113);
xor U11420 (N_11420,N_11167,N_11356);
xnor U11421 (N_11421,N_11277,N_11185);
or U11422 (N_11422,N_11298,N_11367);
nand U11423 (N_11423,N_11218,N_11112);
nor U11424 (N_11424,N_11380,N_11368);
xor U11425 (N_11425,N_11246,N_11235);
xnor U11426 (N_11426,N_11316,N_11279);
or U11427 (N_11427,N_11194,N_11299);
nor U11428 (N_11428,N_11337,N_11118);
xor U11429 (N_11429,N_11353,N_11236);
and U11430 (N_11430,N_11359,N_11302);
and U11431 (N_11431,N_11205,N_11107);
nor U11432 (N_11432,N_11160,N_11172);
and U11433 (N_11433,N_11318,N_11210);
xnor U11434 (N_11434,N_11275,N_11243);
and U11435 (N_11435,N_11155,N_11385);
nand U11436 (N_11436,N_11181,N_11357);
or U11437 (N_11437,N_11276,N_11228);
xnor U11438 (N_11438,N_11291,N_11295);
nor U11439 (N_11439,N_11296,N_11119);
nor U11440 (N_11440,N_11348,N_11378);
and U11441 (N_11441,N_11137,N_11244);
nor U11442 (N_11442,N_11390,N_11332);
or U11443 (N_11443,N_11103,N_11240);
and U11444 (N_11444,N_11338,N_11127);
xnor U11445 (N_11445,N_11170,N_11335);
xor U11446 (N_11446,N_11153,N_11232);
nand U11447 (N_11447,N_11251,N_11161);
xnor U11448 (N_11448,N_11200,N_11239);
and U11449 (N_11449,N_11217,N_11190);
xor U11450 (N_11450,N_11158,N_11126);
nor U11451 (N_11451,N_11355,N_11162);
or U11452 (N_11452,N_11241,N_11343);
and U11453 (N_11453,N_11271,N_11171);
xnor U11454 (N_11454,N_11323,N_11339);
or U11455 (N_11455,N_11146,N_11109);
and U11456 (N_11456,N_11131,N_11231);
xor U11457 (N_11457,N_11386,N_11120);
nand U11458 (N_11458,N_11394,N_11233);
or U11459 (N_11459,N_11134,N_11204);
nand U11460 (N_11460,N_11197,N_11264);
and U11461 (N_11461,N_11382,N_11273);
nor U11462 (N_11462,N_11398,N_11187);
or U11463 (N_11463,N_11163,N_11110);
xnor U11464 (N_11464,N_11370,N_11292);
nor U11465 (N_11465,N_11169,N_11263);
nand U11466 (N_11466,N_11305,N_11361);
nand U11467 (N_11467,N_11144,N_11139);
nand U11468 (N_11468,N_11180,N_11226);
or U11469 (N_11469,N_11106,N_11345);
nand U11470 (N_11470,N_11154,N_11375);
nand U11471 (N_11471,N_11344,N_11173);
or U11472 (N_11472,N_11201,N_11346);
nand U11473 (N_11473,N_11330,N_11141);
xor U11474 (N_11474,N_11145,N_11100);
nor U11475 (N_11475,N_11117,N_11364);
or U11476 (N_11476,N_11388,N_11174);
or U11477 (N_11477,N_11340,N_11142);
xnor U11478 (N_11478,N_11290,N_11270);
and U11479 (N_11479,N_11331,N_11227);
and U11480 (N_11480,N_11269,N_11255);
and U11481 (N_11481,N_11242,N_11358);
nor U11482 (N_11482,N_11147,N_11188);
nor U11483 (N_11483,N_11186,N_11179);
or U11484 (N_11484,N_11389,N_11280);
or U11485 (N_11485,N_11259,N_11341);
nor U11486 (N_11486,N_11177,N_11114);
and U11487 (N_11487,N_11315,N_11278);
or U11488 (N_11488,N_11307,N_11363);
nand U11489 (N_11489,N_11151,N_11136);
nand U11490 (N_11490,N_11221,N_11369);
xor U11491 (N_11491,N_11249,N_11362);
xnor U11492 (N_11492,N_11322,N_11121);
nor U11493 (N_11493,N_11281,N_11152);
or U11494 (N_11494,N_11132,N_11351);
nor U11495 (N_11495,N_11216,N_11268);
xnor U11496 (N_11496,N_11256,N_11247);
or U11497 (N_11497,N_11198,N_11262);
nand U11498 (N_11498,N_11138,N_11166);
nand U11499 (N_11499,N_11266,N_11329);
xor U11500 (N_11500,N_11130,N_11377);
and U11501 (N_11501,N_11104,N_11274);
nand U11502 (N_11502,N_11254,N_11133);
nor U11503 (N_11503,N_11168,N_11202);
xnor U11504 (N_11504,N_11366,N_11253);
nor U11505 (N_11505,N_11245,N_11384);
or U11506 (N_11506,N_11379,N_11212);
or U11507 (N_11507,N_11229,N_11207);
nor U11508 (N_11508,N_11219,N_11283);
nor U11509 (N_11509,N_11123,N_11397);
or U11510 (N_11510,N_11156,N_11125);
xor U11511 (N_11511,N_11293,N_11237);
and U11512 (N_11512,N_11294,N_11101);
xnor U11513 (N_11513,N_11303,N_11148);
or U11514 (N_11514,N_11260,N_11373);
and U11515 (N_11515,N_11220,N_11304);
nand U11516 (N_11516,N_11314,N_11222);
nor U11517 (N_11517,N_11321,N_11327);
and U11518 (N_11518,N_11115,N_11149);
or U11519 (N_11519,N_11143,N_11376);
xor U11520 (N_11520,N_11272,N_11178);
and U11521 (N_11521,N_11193,N_11176);
nand U11522 (N_11522,N_11175,N_11301);
nand U11523 (N_11523,N_11287,N_11191);
and U11524 (N_11524,N_11164,N_11313);
nand U11525 (N_11525,N_11214,N_11116);
nand U11526 (N_11526,N_11354,N_11215);
nand U11527 (N_11527,N_11308,N_11310);
nand U11528 (N_11528,N_11105,N_11350);
nand U11529 (N_11529,N_11111,N_11286);
or U11530 (N_11530,N_11328,N_11372);
and U11531 (N_11531,N_11209,N_11157);
nor U11532 (N_11532,N_11223,N_11381);
xnor U11533 (N_11533,N_11213,N_11248);
or U11534 (N_11534,N_11288,N_11365);
or U11535 (N_11535,N_11159,N_11183);
xnor U11536 (N_11536,N_11297,N_11102);
nand U11537 (N_11537,N_11140,N_11393);
and U11538 (N_11538,N_11234,N_11124);
nand U11539 (N_11539,N_11396,N_11128);
nand U11540 (N_11540,N_11391,N_11150);
nand U11541 (N_11541,N_11300,N_11282);
and U11542 (N_11542,N_11122,N_11285);
nand U11543 (N_11543,N_11360,N_11208);
nand U11544 (N_11544,N_11129,N_11224);
xor U11545 (N_11545,N_11311,N_11352);
nand U11546 (N_11546,N_11199,N_11347);
or U11547 (N_11547,N_11387,N_11182);
nand U11548 (N_11548,N_11196,N_11250);
nand U11549 (N_11549,N_11135,N_11371);
or U11550 (N_11550,N_11267,N_11153);
nand U11551 (N_11551,N_11376,N_11133);
and U11552 (N_11552,N_11251,N_11387);
nor U11553 (N_11553,N_11283,N_11127);
nor U11554 (N_11554,N_11343,N_11350);
xor U11555 (N_11555,N_11362,N_11117);
nor U11556 (N_11556,N_11165,N_11396);
and U11557 (N_11557,N_11144,N_11362);
nor U11558 (N_11558,N_11267,N_11129);
xnor U11559 (N_11559,N_11377,N_11250);
or U11560 (N_11560,N_11173,N_11105);
xnor U11561 (N_11561,N_11356,N_11340);
and U11562 (N_11562,N_11222,N_11399);
xnor U11563 (N_11563,N_11202,N_11380);
and U11564 (N_11564,N_11108,N_11182);
nor U11565 (N_11565,N_11266,N_11257);
and U11566 (N_11566,N_11382,N_11397);
xnor U11567 (N_11567,N_11339,N_11137);
xor U11568 (N_11568,N_11283,N_11113);
or U11569 (N_11569,N_11294,N_11162);
nand U11570 (N_11570,N_11240,N_11223);
or U11571 (N_11571,N_11291,N_11261);
and U11572 (N_11572,N_11218,N_11227);
xnor U11573 (N_11573,N_11174,N_11371);
nor U11574 (N_11574,N_11150,N_11368);
nand U11575 (N_11575,N_11189,N_11293);
or U11576 (N_11576,N_11226,N_11138);
and U11577 (N_11577,N_11239,N_11107);
xor U11578 (N_11578,N_11261,N_11179);
and U11579 (N_11579,N_11141,N_11138);
nand U11580 (N_11580,N_11220,N_11335);
and U11581 (N_11581,N_11329,N_11319);
nor U11582 (N_11582,N_11138,N_11191);
nor U11583 (N_11583,N_11109,N_11293);
or U11584 (N_11584,N_11139,N_11312);
and U11585 (N_11585,N_11351,N_11246);
xnor U11586 (N_11586,N_11146,N_11357);
nor U11587 (N_11587,N_11256,N_11231);
nand U11588 (N_11588,N_11393,N_11186);
and U11589 (N_11589,N_11191,N_11367);
nand U11590 (N_11590,N_11274,N_11253);
xnor U11591 (N_11591,N_11391,N_11372);
nand U11592 (N_11592,N_11134,N_11211);
or U11593 (N_11593,N_11153,N_11370);
xor U11594 (N_11594,N_11254,N_11287);
and U11595 (N_11595,N_11351,N_11234);
xor U11596 (N_11596,N_11198,N_11235);
nor U11597 (N_11597,N_11352,N_11204);
xnor U11598 (N_11598,N_11234,N_11279);
or U11599 (N_11599,N_11356,N_11185);
nor U11600 (N_11600,N_11249,N_11261);
and U11601 (N_11601,N_11177,N_11319);
or U11602 (N_11602,N_11107,N_11336);
nor U11603 (N_11603,N_11113,N_11379);
and U11604 (N_11604,N_11180,N_11191);
and U11605 (N_11605,N_11193,N_11156);
nor U11606 (N_11606,N_11355,N_11267);
nor U11607 (N_11607,N_11279,N_11173);
or U11608 (N_11608,N_11370,N_11281);
nand U11609 (N_11609,N_11288,N_11202);
nand U11610 (N_11610,N_11195,N_11137);
nand U11611 (N_11611,N_11321,N_11350);
or U11612 (N_11612,N_11258,N_11193);
or U11613 (N_11613,N_11395,N_11156);
and U11614 (N_11614,N_11156,N_11207);
nand U11615 (N_11615,N_11352,N_11301);
and U11616 (N_11616,N_11294,N_11214);
nand U11617 (N_11617,N_11327,N_11244);
or U11618 (N_11618,N_11105,N_11301);
nor U11619 (N_11619,N_11155,N_11381);
xnor U11620 (N_11620,N_11133,N_11183);
nand U11621 (N_11621,N_11372,N_11253);
nor U11622 (N_11622,N_11146,N_11102);
and U11623 (N_11623,N_11285,N_11332);
nor U11624 (N_11624,N_11212,N_11273);
nand U11625 (N_11625,N_11201,N_11226);
and U11626 (N_11626,N_11317,N_11121);
xor U11627 (N_11627,N_11119,N_11242);
nand U11628 (N_11628,N_11225,N_11247);
or U11629 (N_11629,N_11380,N_11324);
nor U11630 (N_11630,N_11303,N_11171);
or U11631 (N_11631,N_11208,N_11329);
nor U11632 (N_11632,N_11313,N_11297);
xor U11633 (N_11633,N_11111,N_11246);
xor U11634 (N_11634,N_11162,N_11392);
and U11635 (N_11635,N_11222,N_11186);
and U11636 (N_11636,N_11132,N_11303);
and U11637 (N_11637,N_11257,N_11320);
and U11638 (N_11638,N_11201,N_11265);
or U11639 (N_11639,N_11258,N_11170);
xnor U11640 (N_11640,N_11276,N_11248);
or U11641 (N_11641,N_11135,N_11306);
or U11642 (N_11642,N_11277,N_11233);
nor U11643 (N_11643,N_11308,N_11387);
xor U11644 (N_11644,N_11172,N_11293);
and U11645 (N_11645,N_11362,N_11305);
or U11646 (N_11646,N_11247,N_11335);
nor U11647 (N_11647,N_11331,N_11170);
or U11648 (N_11648,N_11181,N_11370);
xor U11649 (N_11649,N_11191,N_11197);
nor U11650 (N_11650,N_11238,N_11261);
nor U11651 (N_11651,N_11100,N_11125);
xor U11652 (N_11652,N_11283,N_11171);
nor U11653 (N_11653,N_11265,N_11383);
or U11654 (N_11654,N_11326,N_11133);
nor U11655 (N_11655,N_11176,N_11341);
and U11656 (N_11656,N_11281,N_11347);
nor U11657 (N_11657,N_11216,N_11104);
xor U11658 (N_11658,N_11343,N_11246);
nor U11659 (N_11659,N_11399,N_11150);
nor U11660 (N_11660,N_11105,N_11340);
nor U11661 (N_11661,N_11103,N_11102);
or U11662 (N_11662,N_11386,N_11125);
and U11663 (N_11663,N_11392,N_11378);
nor U11664 (N_11664,N_11134,N_11295);
nor U11665 (N_11665,N_11114,N_11323);
or U11666 (N_11666,N_11163,N_11184);
xor U11667 (N_11667,N_11378,N_11324);
xor U11668 (N_11668,N_11329,N_11236);
xor U11669 (N_11669,N_11216,N_11107);
or U11670 (N_11670,N_11141,N_11373);
and U11671 (N_11671,N_11117,N_11342);
nand U11672 (N_11672,N_11172,N_11122);
nor U11673 (N_11673,N_11172,N_11269);
nand U11674 (N_11674,N_11197,N_11193);
and U11675 (N_11675,N_11109,N_11326);
xor U11676 (N_11676,N_11211,N_11150);
nor U11677 (N_11677,N_11188,N_11266);
and U11678 (N_11678,N_11350,N_11225);
nand U11679 (N_11679,N_11202,N_11307);
nor U11680 (N_11680,N_11272,N_11305);
xnor U11681 (N_11681,N_11167,N_11259);
nand U11682 (N_11682,N_11186,N_11302);
or U11683 (N_11683,N_11126,N_11105);
and U11684 (N_11684,N_11316,N_11312);
and U11685 (N_11685,N_11125,N_11204);
or U11686 (N_11686,N_11221,N_11240);
nand U11687 (N_11687,N_11348,N_11291);
or U11688 (N_11688,N_11144,N_11198);
and U11689 (N_11689,N_11386,N_11318);
nand U11690 (N_11690,N_11321,N_11167);
xnor U11691 (N_11691,N_11191,N_11396);
xnor U11692 (N_11692,N_11338,N_11373);
nor U11693 (N_11693,N_11215,N_11343);
nor U11694 (N_11694,N_11222,N_11304);
or U11695 (N_11695,N_11141,N_11263);
xnor U11696 (N_11696,N_11388,N_11253);
nor U11697 (N_11697,N_11150,N_11173);
xnor U11698 (N_11698,N_11354,N_11176);
nor U11699 (N_11699,N_11183,N_11111);
and U11700 (N_11700,N_11683,N_11626);
nor U11701 (N_11701,N_11587,N_11554);
nand U11702 (N_11702,N_11528,N_11437);
nand U11703 (N_11703,N_11568,N_11469);
or U11704 (N_11704,N_11531,N_11570);
and U11705 (N_11705,N_11603,N_11546);
and U11706 (N_11706,N_11592,N_11478);
nor U11707 (N_11707,N_11474,N_11460);
nor U11708 (N_11708,N_11645,N_11441);
nand U11709 (N_11709,N_11612,N_11566);
and U11710 (N_11710,N_11442,N_11553);
nand U11711 (N_11711,N_11640,N_11428);
xor U11712 (N_11712,N_11614,N_11471);
nand U11713 (N_11713,N_11473,N_11615);
nand U11714 (N_11714,N_11682,N_11608);
or U11715 (N_11715,N_11430,N_11506);
or U11716 (N_11716,N_11485,N_11527);
and U11717 (N_11717,N_11650,N_11618);
xnor U11718 (N_11718,N_11464,N_11691);
xnor U11719 (N_11719,N_11627,N_11405);
nor U11720 (N_11720,N_11569,N_11468);
and U11721 (N_11721,N_11481,N_11556);
and U11722 (N_11722,N_11449,N_11545);
nand U11723 (N_11723,N_11492,N_11551);
nand U11724 (N_11724,N_11681,N_11687);
or U11725 (N_11725,N_11567,N_11661);
and U11726 (N_11726,N_11417,N_11654);
and U11727 (N_11727,N_11605,N_11600);
xor U11728 (N_11728,N_11511,N_11439);
xor U11729 (N_11729,N_11524,N_11581);
nand U11730 (N_11730,N_11659,N_11542);
or U11731 (N_11731,N_11558,N_11678);
or U11732 (N_11732,N_11697,N_11443);
or U11733 (N_11733,N_11622,N_11418);
xnor U11734 (N_11734,N_11550,N_11504);
nand U11735 (N_11735,N_11571,N_11540);
xnor U11736 (N_11736,N_11619,N_11457);
xor U11737 (N_11737,N_11631,N_11672);
xor U11738 (N_11738,N_11412,N_11467);
or U11739 (N_11739,N_11580,N_11692);
or U11740 (N_11740,N_11561,N_11557);
xnor U11741 (N_11741,N_11611,N_11657);
and U11742 (N_11742,N_11610,N_11634);
and U11743 (N_11743,N_11680,N_11564);
xor U11744 (N_11744,N_11695,N_11547);
and U11745 (N_11745,N_11572,N_11498);
or U11746 (N_11746,N_11676,N_11693);
or U11747 (N_11747,N_11447,N_11532);
and U11748 (N_11748,N_11646,N_11422);
and U11749 (N_11749,N_11671,N_11414);
and U11750 (N_11750,N_11409,N_11625);
nor U11751 (N_11751,N_11477,N_11491);
or U11752 (N_11752,N_11549,N_11628);
and U11753 (N_11753,N_11451,N_11589);
xnor U11754 (N_11754,N_11617,N_11529);
nand U11755 (N_11755,N_11520,N_11413);
and U11756 (N_11756,N_11643,N_11655);
or U11757 (N_11757,N_11544,N_11501);
nand U11758 (N_11758,N_11679,N_11548);
xor U11759 (N_11759,N_11578,N_11456);
xor U11760 (N_11760,N_11674,N_11694);
nand U11761 (N_11761,N_11484,N_11486);
or U11762 (N_11762,N_11688,N_11462);
nor U11763 (N_11763,N_11642,N_11653);
and U11764 (N_11764,N_11593,N_11660);
nor U11765 (N_11765,N_11475,N_11648);
or U11766 (N_11766,N_11601,N_11510);
and U11767 (N_11767,N_11662,N_11526);
nor U11768 (N_11768,N_11472,N_11508);
nor U11769 (N_11769,N_11584,N_11543);
and U11770 (N_11770,N_11480,N_11665);
nand U11771 (N_11771,N_11401,N_11555);
nand U11772 (N_11772,N_11696,N_11470);
nand U11773 (N_11773,N_11502,N_11639);
xor U11774 (N_11774,N_11582,N_11533);
or U11775 (N_11775,N_11579,N_11416);
nand U11776 (N_11776,N_11522,N_11434);
xor U11777 (N_11777,N_11512,N_11466);
xor U11778 (N_11778,N_11597,N_11652);
and U11779 (N_11779,N_11596,N_11499);
xor U11780 (N_11780,N_11559,N_11591);
xnor U11781 (N_11781,N_11667,N_11541);
nor U11782 (N_11782,N_11440,N_11433);
and U11783 (N_11783,N_11641,N_11429);
nand U11784 (N_11784,N_11586,N_11656);
xor U11785 (N_11785,N_11535,N_11431);
and U11786 (N_11786,N_11613,N_11560);
and U11787 (N_11787,N_11454,N_11609);
nand U11788 (N_11788,N_11415,N_11523);
or U11789 (N_11789,N_11624,N_11452);
nor U11790 (N_11790,N_11500,N_11463);
nand U11791 (N_11791,N_11583,N_11668);
nor U11792 (N_11792,N_11632,N_11699);
nor U11793 (N_11793,N_11664,N_11515);
and U11794 (N_11794,N_11517,N_11419);
and U11795 (N_11795,N_11493,N_11516);
nor U11796 (N_11796,N_11444,N_11505);
nor U11797 (N_11797,N_11436,N_11448);
nand U11798 (N_11798,N_11513,N_11420);
xnor U11799 (N_11799,N_11423,N_11651);
or U11800 (N_11800,N_11530,N_11489);
xnor U11801 (N_11801,N_11590,N_11573);
or U11802 (N_11802,N_11621,N_11686);
xor U11803 (N_11803,N_11574,N_11604);
and U11804 (N_11804,N_11446,N_11607);
nand U11805 (N_11805,N_11488,N_11636);
nand U11806 (N_11806,N_11459,N_11509);
nand U11807 (N_11807,N_11514,N_11616);
xor U11808 (N_11808,N_11689,N_11534);
nor U11809 (N_11809,N_11407,N_11518);
and U11810 (N_11810,N_11690,N_11404);
nor U11811 (N_11811,N_11461,N_11482);
and U11812 (N_11812,N_11487,N_11411);
xnor U11813 (N_11813,N_11503,N_11666);
nand U11814 (N_11814,N_11408,N_11403);
and U11815 (N_11815,N_11406,N_11400);
nand U11816 (N_11816,N_11453,N_11519);
or U11817 (N_11817,N_11644,N_11649);
nand U11818 (N_11818,N_11675,N_11563);
xor U11819 (N_11819,N_11450,N_11495);
nor U11820 (N_11820,N_11565,N_11496);
nor U11821 (N_11821,N_11562,N_11435);
nor U11822 (N_11822,N_11685,N_11635);
or U11823 (N_11823,N_11426,N_11476);
nor U11824 (N_11824,N_11637,N_11536);
xnor U11825 (N_11825,N_11494,N_11673);
xnor U11826 (N_11826,N_11669,N_11537);
xor U11827 (N_11827,N_11677,N_11585);
and U11828 (N_11828,N_11698,N_11658);
nor U11829 (N_11829,N_11602,N_11521);
xor U11830 (N_11830,N_11445,N_11647);
nor U11831 (N_11831,N_11630,N_11629);
and U11832 (N_11832,N_11424,N_11432);
or U11833 (N_11833,N_11490,N_11575);
xnor U11834 (N_11834,N_11497,N_11479);
or U11835 (N_11835,N_11620,N_11670);
nand U11836 (N_11836,N_11507,N_11421);
nor U11837 (N_11837,N_11595,N_11663);
or U11838 (N_11838,N_11483,N_11402);
and U11839 (N_11839,N_11633,N_11538);
nand U11840 (N_11840,N_11599,N_11465);
nand U11841 (N_11841,N_11425,N_11598);
nand U11842 (N_11842,N_11410,N_11623);
or U11843 (N_11843,N_11684,N_11606);
nor U11844 (N_11844,N_11525,N_11594);
nand U11845 (N_11845,N_11539,N_11458);
xor U11846 (N_11846,N_11438,N_11552);
or U11847 (N_11847,N_11576,N_11638);
xnor U11848 (N_11848,N_11455,N_11577);
xor U11849 (N_11849,N_11427,N_11588);
or U11850 (N_11850,N_11590,N_11471);
nand U11851 (N_11851,N_11638,N_11675);
nand U11852 (N_11852,N_11625,N_11684);
or U11853 (N_11853,N_11602,N_11636);
xnor U11854 (N_11854,N_11610,N_11674);
nand U11855 (N_11855,N_11559,N_11589);
nor U11856 (N_11856,N_11521,N_11508);
nand U11857 (N_11857,N_11536,N_11646);
nor U11858 (N_11858,N_11444,N_11464);
nand U11859 (N_11859,N_11638,N_11429);
xnor U11860 (N_11860,N_11627,N_11451);
and U11861 (N_11861,N_11447,N_11594);
nand U11862 (N_11862,N_11605,N_11472);
xnor U11863 (N_11863,N_11513,N_11694);
or U11864 (N_11864,N_11577,N_11524);
xor U11865 (N_11865,N_11622,N_11696);
xor U11866 (N_11866,N_11510,N_11421);
nor U11867 (N_11867,N_11694,N_11554);
and U11868 (N_11868,N_11681,N_11666);
nor U11869 (N_11869,N_11495,N_11400);
or U11870 (N_11870,N_11458,N_11519);
xor U11871 (N_11871,N_11642,N_11511);
xnor U11872 (N_11872,N_11673,N_11567);
or U11873 (N_11873,N_11603,N_11454);
nor U11874 (N_11874,N_11468,N_11541);
and U11875 (N_11875,N_11624,N_11462);
nand U11876 (N_11876,N_11623,N_11698);
or U11877 (N_11877,N_11513,N_11548);
nor U11878 (N_11878,N_11402,N_11677);
xor U11879 (N_11879,N_11497,N_11543);
nand U11880 (N_11880,N_11653,N_11485);
or U11881 (N_11881,N_11623,N_11423);
or U11882 (N_11882,N_11678,N_11610);
and U11883 (N_11883,N_11516,N_11447);
nor U11884 (N_11884,N_11618,N_11668);
xnor U11885 (N_11885,N_11601,N_11516);
nand U11886 (N_11886,N_11683,N_11491);
nor U11887 (N_11887,N_11440,N_11676);
nand U11888 (N_11888,N_11503,N_11542);
nand U11889 (N_11889,N_11642,N_11523);
nand U11890 (N_11890,N_11434,N_11587);
or U11891 (N_11891,N_11408,N_11469);
and U11892 (N_11892,N_11515,N_11608);
xnor U11893 (N_11893,N_11505,N_11598);
or U11894 (N_11894,N_11436,N_11437);
or U11895 (N_11895,N_11474,N_11415);
and U11896 (N_11896,N_11660,N_11418);
xor U11897 (N_11897,N_11544,N_11526);
and U11898 (N_11898,N_11614,N_11466);
and U11899 (N_11899,N_11534,N_11611);
nor U11900 (N_11900,N_11433,N_11450);
nand U11901 (N_11901,N_11686,N_11648);
nor U11902 (N_11902,N_11463,N_11672);
nor U11903 (N_11903,N_11488,N_11456);
xnor U11904 (N_11904,N_11625,N_11558);
xnor U11905 (N_11905,N_11665,N_11690);
or U11906 (N_11906,N_11587,N_11614);
xnor U11907 (N_11907,N_11610,N_11565);
or U11908 (N_11908,N_11657,N_11583);
nor U11909 (N_11909,N_11563,N_11456);
and U11910 (N_11910,N_11451,N_11674);
xor U11911 (N_11911,N_11519,N_11466);
nand U11912 (N_11912,N_11591,N_11688);
or U11913 (N_11913,N_11509,N_11472);
nand U11914 (N_11914,N_11400,N_11421);
or U11915 (N_11915,N_11416,N_11632);
and U11916 (N_11916,N_11590,N_11604);
or U11917 (N_11917,N_11639,N_11657);
xnor U11918 (N_11918,N_11582,N_11664);
nand U11919 (N_11919,N_11515,N_11502);
nand U11920 (N_11920,N_11625,N_11445);
nor U11921 (N_11921,N_11683,N_11663);
nor U11922 (N_11922,N_11458,N_11513);
or U11923 (N_11923,N_11542,N_11689);
and U11924 (N_11924,N_11432,N_11670);
nor U11925 (N_11925,N_11633,N_11445);
xor U11926 (N_11926,N_11507,N_11686);
nand U11927 (N_11927,N_11455,N_11554);
xor U11928 (N_11928,N_11688,N_11427);
or U11929 (N_11929,N_11458,N_11588);
xnor U11930 (N_11930,N_11521,N_11647);
nand U11931 (N_11931,N_11510,N_11650);
xnor U11932 (N_11932,N_11557,N_11621);
and U11933 (N_11933,N_11515,N_11600);
nor U11934 (N_11934,N_11529,N_11480);
and U11935 (N_11935,N_11522,N_11505);
nand U11936 (N_11936,N_11549,N_11637);
xnor U11937 (N_11937,N_11495,N_11631);
nand U11938 (N_11938,N_11462,N_11588);
or U11939 (N_11939,N_11586,N_11693);
xnor U11940 (N_11940,N_11451,N_11592);
xor U11941 (N_11941,N_11449,N_11573);
or U11942 (N_11942,N_11452,N_11641);
nand U11943 (N_11943,N_11497,N_11699);
xor U11944 (N_11944,N_11611,N_11415);
or U11945 (N_11945,N_11640,N_11471);
or U11946 (N_11946,N_11661,N_11483);
or U11947 (N_11947,N_11604,N_11513);
nand U11948 (N_11948,N_11429,N_11555);
or U11949 (N_11949,N_11522,N_11591);
xor U11950 (N_11950,N_11536,N_11690);
and U11951 (N_11951,N_11430,N_11608);
nor U11952 (N_11952,N_11431,N_11657);
and U11953 (N_11953,N_11664,N_11696);
and U11954 (N_11954,N_11653,N_11567);
and U11955 (N_11955,N_11425,N_11675);
xor U11956 (N_11956,N_11672,N_11517);
and U11957 (N_11957,N_11645,N_11638);
nor U11958 (N_11958,N_11666,N_11591);
or U11959 (N_11959,N_11500,N_11444);
nor U11960 (N_11960,N_11519,N_11408);
or U11961 (N_11961,N_11604,N_11584);
or U11962 (N_11962,N_11690,N_11597);
and U11963 (N_11963,N_11551,N_11572);
xor U11964 (N_11964,N_11639,N_11440);
and U11965 (N_11965,N_11443,N_11505);
and U11966 (N_11966,N_11555,N_11570);
xnor U11967 (N_11967,N_11524,N_11429);
nor U11968 (N_11968,N_11684,N_11550);
nor U11969 (N_11969,N_11537,N_11547);
nor U11970 (N_11970,N_11553,N_11584);
xor U11971 (N_11971,N_11531,N_11557);
xnor U11972 (N_11972,N_11408,N_11419);
or U11973 (N_11973,N_11644,N_11596);
and U11974 (N_11974,N_11694,N_11529);
and U11975 (N_11975,N_11582,N_11587);
nand U11976 (N_11976,N_11683,N_11604);
and U11977 (N_11977,N_11557,N_11448);
and U11978 (N_11978,N_11679,N_11480);
and U11979 (N_11979,N_11649,N_11445);
and U11980 (N_11980,N_11595,N_11486);
or U11981 (N_11981,N_11636,N_11600);
nand U11982 (N_11982,N_11612,N_11425);
or U11983 (N_11983,N_11602,N_11480);
and U11984 (N_11984,N_11688,N_11546);
xor U11985 (N_11985,N_11547,N_11400);
nor U11986 (N_11986,N_11401,N_11672);
or U11987 (N_11987,N_11471,N_11684);
xor U11988 (N_11988,N_11663,N_11499);
nand U11989 (N_11989,N_11443,N_11661);
and U11990 (N_11990,N_11661,N_11647);
xnor U11991 (N_11991,N_11570,N_11536);
nand U11992 (N_11992,N_11410,N_11520);
nor U11993 (N_11993,N_11493,N_11468);
nand U11994 (N_11994,N_11580,N_11697);
nor U11995 (N_11995,N_11692,N_11575);
and U11996 (N_11996,N_11454,N_11467);
or U11997 (N_11997,N_11647,N_11585);
nor U11998 (N_11998,N_11653,N_11526);
nor U11999 (N_11999,N_11695,N_11556);
nor U12000 (N_12000,N_11898,N_11887);
xor U12001 (N_12001,N_11897,N_11750);
nand U12002 (N_12002,N_11822,N_11793);
and U12003 (N_12003,N_11998,N_11716);
and U12004 (N_12004,N_11771,N_11896);
xnor U12005 (N_12005,N_11916,N_11746);
and U12006 (N_12006,N_11962,N_11761);
nand U12007 (N_12007,N_11739,N_11745);
and U12008 (N_12008,N_11828,N_11755);
nor U12009 (N_12009,N_11711,N_11843);
and U12010 (N_12010,N_11769,N_11809);
xnor U12011 (N_12011,N_11965,N_11768);
xor U12012 (N_12012,N_11732,N_11800);
nand U12013 (N_12013,N_11770,N_11879);
nand U12014 (N_12014,N_11859,N_11777);
nor U12015 (N_12015,N_11984,N_11886);
xor U12016 (N_12016,N_11774,N_11786);
xor U12017 (N_12017,N_11707,N_11999);
xor U12018 (N_12018,N_11747,N_11900);
nor U12019 (N_12019,N_11811,N_11954);
nand U12020 (N_12020,N_11977,N_11776);
and U12021 (N_12021,N_11851,N_11881);
nor U12022 (N_12022,N_11903,N_11705);
or U12023 (N_12023,N_11955,N_11704);
nand U12024 (N_12024,N_11748,N_11890);
nand U12025 (N_12025,N_11812,N_11784);
and U12026 (N_12026,N_11922,N_11734);
or U12027 (N_12027,N_11972,N_11714);
nor U12028 (N_12028,N_11789,N_11971);
nor U12029 (N_12029,N_11844,N_11960);
nor U12030 (N_12030,N_11966,N_11724);
nand U12031 (N_12031,N_11835,N_11940);
nand U12032 (N_12032,N_11762,N_11941);
xnor U12033 (N_12033,N_11866,N_11969);
and U12034 (N_12034,N_11939,N_11968);
nand U12035 (N_12035,N_11782,N_11970);
xnor U12036 (N_12036,N_11953,N_11820);
nor U12037 (N_12037,N_11723,N_11833);
xor U12038 (N_12038,N_11823,N_11801);
or U12039 (N_12039,N_11810,N_11956);
and U12040 (N_12040,N_11904,N_11985);
xor U12041 (N_12041,N_11925,N_11760);
nor U12042 (N_12042,N_11710,N_11997);
nor U12043 (N_12043,N_11738,N_11882);
and U12044 (N_12044,N_11753,N_11974);
and U12045 (N_12045,N_11749,N_11908);
nor U12046 (N_12046,N_11807,N_11781);
and U12047 (N_12047,N_11778,N_11743);
or U12048 (N_12048,N_11964,N_11715);
nor U12049 (N_12049,N_11744,N_11740);
nand U12050 (N_12050,N_11899,N_11867);
nor U12051 (N_12051,N_11799,N_11934);
and U12052 (N_12052,N_11913,N_11936);
nand U12053 (N_12053,N_11856,N_11952);
nand U12054 (N_12054,N_11795,N_11728);
xor U12055 (N_12055,N_11868,N_11901);
or U12056 (N_12056,N_11788,N_11979);
or U12057 (N_12057,N_11730,N_11860);
nand U12058 (N_12058,N_11864,N_11923);
nor U12059 (N_12059,N_11836,N_11871);
nand U12060 (N_12060,N_11764,N_11891);
nand U12061 (N_12061,N_11862,N_11992);
nand U12062 (N_12062,N_11990,N_11712);
and U12063 (N_12063,N_11910,N_11931);
or U12064 (N_12064,N_11830,N_11794);
nand U12065 (N_12065,N_11973,N_11987);
nand U12066 (N_12066,N_11829,N_11976);
xor U12067 (N_12067,N_11855,N_11736);
and U12068 (N_12068,N_11785,N_11709);
or U12069 (N_12069,N_11909,N_11727);
nor U12070 (N_12070,N_11889,N_11995);
xor U12071 (N_12071,N_11991,N_11927);
and U12072 (N_12072,N_11919,N_11779);
xnor U12073 (N_12073,N_11702,N_11834);
xnor U12074 (N_12074,N_11842,N_11735);
and U12075 (N_12075,N_11967,N_11854);
xor U12076 (N_12076,N_11983,N_11751);
nor U12077 (N_12077,N_11752,N_11975);
and U12078 (N_12078,N_11847,N_11877);
nand U12079 (N_12079,N_11825,N_11959);
or U12080 (N_12080,N_11827,N_11920);
nor U12081 (N_12081,N_11905,N_11872);
and U12082 (N_12082,N_11846,N_11733);
xor U12083 (N_12083,N_11742,N_11837);
nand U12084 (N_12084,N_11957,N_11758);
nor U12085 (N_12085,N_11848,N_11773);
or U12086 (N_12086,N_11763,N_11792);
nand U12087 (N_12087,N_11857,N_11849);
nor U12088 (N_12088,N_11943,N_11850);
and U12089 (N_12089,N_11708,N_11845);
nand U12090 (N_12090,N_11918,N_11721);
xnor U12091 (N_12091,N_11982,N_11933);
nor U12092 (N_12092,N_11852,N_11924);
and U12093 (N_12093,N_11902,N_11767);
or U12094 (N_12094,N_11884,N_11719);
and U12095 (N_12095,N_11892,N_11858);
nor U12096 (N_12096,N_11808,N_11963);
xnor U12097 (N_12097,N_11726,N_11949);
nor U12098 (N_12098,N_11951,N_11706);
nor U12099 (N_12099,N_11865,N_11831);
nor U12100 (N_12100,N_11894,N_11791);
nand U12101 (N_12101,N_11988,N_11765);
nand U12102 (N_12102,N_11814,N_11821);
and U12103 (N_12103,N_11838,N_11701);
or U12104 (N_12104,N_11895,N_11945);
or U12105 (N_12105,N_11840,N_11928);
and U12106 (N_12106,N_11797,N_11861);
nor U12107 (N_12107,N_11802,N_11935);
nor U12108 (N_12108,N_11880,N_11790);
and U12109 (N_12109,N_11841,N_11722);
nor U12110 (N_12110,N_11921,N_11937);
nor U12111 (N_12111,N_11870,N_11805);
xor U12112 (N_12112,N_11873,N_11832);
or U12113 (N_12113,N_11826,N_11875);
xor U12114 (N_12114,N_11725,N_11766);
nor U12115 (N_12115,N_11819,N_11942);
and U12116 (N_12116,N_11796,N_11981);
and U12117 (N_12117,N_11803,N_11729);
or U12118 (N_12118,N_11772,N_11944);
xnor U12119 (N_12119,N_11888,N_11938);
nor U12120 (N_12120,N_11914,N_11932);
xnor U12121 (N_12121,N_11915,N_11713);
nand U12122 (N_12122,N_11783,N_11839);
nor U12123 (N_12123,N_11961,N_11718);
and U12124 (N_12124,N_11893,N_11885);
nor U12125 (N_12125,N_11780,N_11816);
and U12126 (N_12126,N_11703,N_11817);
xnor U12127 (N_12127,N_11720,N_11929);
xnor U12128 (N_12128,N_11756,N_11930);
xnor U12129 (N_12129,N_11989,N_11950);
nor U12130 (N_12130,N_11717,N_11759);
nor U12131 (N_12131,N_11804,N_11993);
xnor U12132 (N_12132,N_11986,N_11876);
or U12133 (N_12133,N_11947,N_11757);
or U12134 (N_12134,N_11948,N_11878);
and U12135 (N_12135,N_11853,N_11911);
xor U12136 (N_12136,N_11754,N_11863);
or U12137 (N_12137,N_11737,N_11806);
or U12138 (N_12138,N_11741,N_11996);
xor U12139 (N_12139,N_11912,N_11700);
xor U12140 (N_12140,N_11926,N_11883);
xnor U12141 (N_12141,N_11798,N_11907);
nand U12142 (N_12142,N_11818,N_11731);
and U12143 (N_12143,N_11787,N_11824);
or U12144 (N_12144,N_11917,N_11813);
xor U12145 (N_12145,N_11978,N_11980);
nor U12146 (N_12146,N_11874,N_11958);
and U12147 (N_12147,N_11906,N_11775);
xnor U12148 (N_12148,N_11994,N_11815);
nand U12149 (N_12149,N_11869,N_11946);
nand U12150 (N_12150,N_11895,N_11833);
nand U12151 (N_12151,N_11886,N_11916);
xor U12152 (N_12152,N_11720,N_11976);
nand U12153 (N_12153,N_11965,N_11789);
nor U12154 (N_12154,N_11883,N_11846);
or U12155 (N_12155,N_11770,N_11973);
nor U12156 (N_12156,N_11958,N_11833);
xnor U12157 (N_12157,N_11879,N_11864);
or U12158 (N_12158,N_11894,N_11958);
nor U12159 (N_12159,N_11781,N_11880);
nand U12160 (N_12160,N_11773,N_11763);
nor U12161 (N_12161,N_11954,N_11745);
nor U12162 (N_12162,N_11893,N_11733);
and U12163 (N_12163,N_11902,N_11985);
nand U12164 (N_12164,N_11702,N_11844);
nor U12165 (N_12165,N_11754,N_11971);
nor U12166 (N_12166,N_11978,N_11883);
xor U12167 (N_12167,N_11796,N_11868);
nor U12168 (N_12168,N_11788,N_11838);
and U12169 (N_12169,N_11837,N_11789);
nand U12170 (N_12170,N_11939,N_11875);
xnor U12171 (N_12171,N_11863,N_11946);
and U12172 (N_12172,N_11829,N_11711);
or U12173 (N_12173,N_11721,N_11868);
or U12174 (N_12174,N_11704,N_11813);
and U12175 (N_12175,N_11765,N_11713);
or U12176 (N_12176,N_11763,N_11844);
nand U12177 (N_12177,N_11814,N_11986);
or U12178 (N_12178,N_11818,N_11980);
and U12179 (N_12179,N_11742,N_11956);
and U12180 (N_12180,N_11970,N_11956);
and U12181 (N_12181,N_11875,N_11845);
nor U12182 (N_12182,N_11927,N_11996);
nand U12183 (N_12183,N_11881,N_11858);
nor U12184 (N_12184,N_11954,N_11785);
nor U12185 (N_12185,N_11904,N_11810);
or U12186 (N_12186,N_11838,N_11743);
nand U12187 (N_12187,N_11760,N_11849);
and U12188 (N_12188,N_11727,N_11759);
xnor U12189 (N_12189,N_11997,N_11876);
and U12190 (N_12190,N_11788,N_11781);
nor U12191 (N_12191,N_11747,N_11833);
or U12192 (N_12192,N_11941,N_11958);
or U12193 (N_12193,N_11758,N_11941);
and U12194 (N_12194,N_11970,N_11964);
and U12195 (N_12195,N_11862,N_11969);
nand U12196 (N_12196,N_11736,N_11763);
nand U12197 (N_12197,N_11748,N_11941);
nand U12198 (N_12198,N_11721,N_11786);
and U12199 (N_12199,N_11973,N_11729);
or U12200 (N_12200,N_11907,N_11725);
nor U12201 (N_12201,N_11859,N_11876);
or U12202 (N_12202,N_11800,N_11749);
nor U12203 (N_12203,N_11895,N_11943);
nand U12204 (N_12204,N_11809,N_11937);
nand U12205 (N_12205,N_11974,N_11852);
nand U12206 (N_12206,N_11938,N_11790);
and U12207 (N_12207,N_11779,N_11795);
nor U12208 (N_12208,N_11994,N_11891);
xor U12209 (N_12209,N_11822,N_11892);
nor U12210 (N_12210,N_11957,N_11750);
nand U12211 (N_12211,N_11756,N_11810);
and U12212 (N_12212,N_11931,N_11748);
xnor U12213 (N_12213,N_11804,N_11755);
and U12214 (N_12214,N_11761,N_11801);
or U12215 (N_12215,N_11932,N_11827);
nand U12216 (N_12216,N_11981,N_11760);
or U12217 (N_12217,N_11958,N_11922);
nor U12218 (N_12218,N_11756,N_11993);
and U12219 (N_12219,N_11981,N_11952);
and U12220 (N_12220,N_11907,N_11930);
xnor U12221 (N_12221,N_11912,N_11882);
and U12222 (N_12222,N_11861,N_11770);
and U12223 (N_12223,N_11851,N_11709);
and U12224 (N_12224,N_11886,N_11746);
xnor U12225 (N_12225,N_11781,N_11802);
nor U12226 (N_12226,N_11830,N_11776);
nor U12227 (N_12227,N_11994,N_11936);
nand U12228 (N_12228,N_11964,N_11800);
xor U12229 (N_12229,N_11716,N_11809);
nand U12230 (N_12230,N_11787,N_11721);
nand U12231 (N_12231,N_11858,N_11755);
nand U12232 (N_12232,N_11783,N_11768);
nor U12233 (N_12233,N_11751,N_11956);
nand U12234 (N_12234,N_11742,N_11781);
and U12235 (N_12235,N_11839,N_11708);
nand U12236 (N_12236,N_11888,N_11709);
and U12237 (N_12237,N_11806,N_11902);
nand U12238 (N_12238,N_11857,N_11723);
and U12239 (N_12239,N_11768,N_11715);
nand U12240 (N_12240,N_11721,N_11906);
and U12241 (N_12241,N_11883,N_11726);
xor U12242 (N_12242,N_11900,N_11730);
xor U12243 (N_12243,N_11737,N_11908);
nor U12244 (N_12244,N_11967,N_11800);
or U12245 (N_12245,N_11785,N_11783);
or U12246 (N_12246,N_11799,N_11706);
xnor U12247 (N_12247,N_11747,N_11731);
nor U12248 (N_12248,N_11727,N_11769);
nand U12249 (N_12249,N_11934,N_11928);
and U12250 (N_12250,N_11889,N_11734);
xor U12251 (N_12251,N_11886,N_11995);
nand U12252 (N_12252,N_11976,N_11822);
nor U12253 (N_12253,N_11959,N_11702);
xnor U12254 (N_12254,N_11844,N_11807);
nand U12255 (N_12255,N_11825,N_11874);
nand U12256 (N_12256,N_11952,N_11914);
nand U12257 (N_12257,N_11710,N_11800);
xor U12258 (N_12258,N_11882,N_11724);
and U12259 (N_12259,N_11892,N_11931);
and U12260 (N_12260,N_11939,N_11805);
nor U12261 (N_12261,N_11827,N_11971);
or U12262 (N_12262,N_11861,N_11847);
xnor U12263 (N_12263,N_11779,N_11882);
or U12264 (N_12264,N_11998,N_11786);
nor U12265 (N_12265,N_11797,N_11940);
and U12266 (N_12266,N_11903,N_11807);
or U12267 (N_12267,N_11882,N_11838);
xor U12268 (N_12268,N_11984,N_11710);
nor U12269 (N_12269,N_11727,N_11839);
nor U12270 (N_12270,N_11856,N_11872);
nor U12271 (N_12271,N_11777,N_11984);
xor U12272 (N_12272,N_11847,N_11810);
nand U12273 (N_12273,N_11818,N_11931);
and U12274 (N_12274,N_11729,N_11870);
nand U12275 (N_12275,N_11860,N_11888);
nand U12276 (N_12276,N_11949,N_11976);
and U12277 (N_12277,N_11776,N_11846);
or U12278 (N_12278,N_11935,N_11867);
and U12279 (N_12279,N_11772,N_11797);
nor U12280 (N_12280,N_11994,N_11742);
xnor U12281 (N_12281,N_11900,N_11781);
xor U12282 (N_12282,N_11751,N_11790);
nand U12283 (N_12283,N_11981,N_11806);
and U12284 (N_12284,N_11770,N_11743);
and U12285 (N_12285,N_11908,N_11848);
and U12286 (N_12286,N_11933,N_11752);
or U12287 (N_12287,N_11993,N_11712);
nor U12288 (N_12288,N_11744,N_11882);
nor U12289 (N_12289,N_11912,N_11727);
or U12290 (N_12290,N_11832,N_11818);
and U12291 (N_12291,N_11911,N_11982);
xnor U12292 (N_12292,N_11735,N_11806);
xnor U12293 (N_12293,N_11853,N_11796);
or U12294 (N_12294,N_11877,N_11849);
nand U12295 (N_12295,N_11940,N_11763);
nor U12296 (N_12296,N_11912,N_11714);
nor U12297 (N_12297,N_11834,N_11932);
nor U12298 (N_12298,N_11750,N_11852);
nand U12299 (N_12299,N_11733,N_11997);
nor U12300 (N_12300,N_12299,N_12081);
and U12301 (N_12301,N_12236,N_12246);
and U12302 (N_12302,N_12148,N_12279);
nor U12303 (N_12303,N_12225,N_12056);
nor U12304 (N_12304,N_12182,N_12166);
xor U12305 (N_12305,N_12152,N_12180);
and U12306 (N_12306,N_12256,N_12178);
nor U12307 (N_12307,N_12289,N_12202);
or U12308 (N_12308,N_12006,N_12031);
xor U12309 (N_12309,N_12083,N_12224);
or U12310 (N_12310,N_12276,N_12046);
nand U12311 (N_12311,N_12297,N_12282);
nor U12312 (N_12312,N_12157,N_12238);
xor U12313 (N_12313,N_12112,N_12141);
and U12314 (N_12314,N_12292,N_12001);
nor U12315 (N_12315,N_12003,N_12160);
xnor U12316 (N_12316,N_12219,N_12241);
or U12317 (N_12317,N_12154,N_12260);
nand U12318 (N_12318,N_12275,N_12145);
xnor U12319 (N_12319,N_12211,N_12125);
or U12320 (N_12320,N_12071,N_12229);
and U12321 (N_12321,N_12095,N_12084);
and U12322 (N_12322,N_12207,N_12209);
nor U12323 (N_12323,N_12203,N_12281);
nor U12324 (N_12324,N_12082,N_12103);
and U12325 (N_12325,N_12264,N_12023);
xnor U12326 (N_12326,N_12263,N_12106);
xnor U12327 (N_12327,N_12052,N_12069);
nand U12328 (N_12328,N_12242,N_12042);
and U12329 (N_12329,N_12284,N_12220);
or U12330 (N_12330,N_12265,N_12005);
nand U12331 (N_12331,N_12129,N_12198);
nor U12332 (N_12332,N_12155,N_12065);
or U12333 (N_12333,N_12000,N_12175);
and U12334 (N_12334,N_12146,N_12015);
nand U12335 (N_12335,N_12033,N_12269);
or U12336 (N_12336,N_12171,N_12009);
or U12337 (N_12337,N_12113,N_12210);
nor U12338 (N_12338,N_12019,N_12123);
nand U12339 (N_12339,N_12294,N_12067);
nand U12340 (N_12340,N_12161,N_12205);
and U12341 (N_12341,N_12101,N_12173);
nand U12342 (N_12342,N_12085,N_12286);
nand U12343 (N_12343,N_12233,N_12190);
and U12344 (N_12344,N_12298,N_12092);
xor U12345 (N_12345,N_12114,N_12057);
and U12346 (N_12346,N_12017,N_12119);
nor U12347 (N_12347,N_12077,N_12251);
xor U12348 (N_12348,N_12290,N_12247);
nor U12349 (N_12349,N_12087,N_12226);
nor U12350 (N_12350,N_12061,N_12127);
nand U12351 (N_12351,N_12147,N_12158);
xor U12352 (N_12352,N_12194,N_12250);
nand U12353 (N_12353,N_12159,N_12266);
and U12354 (N_12354,N_12107,N_12140);
xnor U12355 (N_12355,N_12218,N_12075);
xnor U12356 (N_12356,N_12039,N_12153);
or U12357 (N_12357,N_12104,N_12167);
nor U12358 (N_12358,N_12184,N_12115);
nor U12359 (N_12359,N_12164,N_12174);
or U12360 (N_12360,N_12035,N_12197);
nor U12361 (N_12361,N_12016,N_12192);
nor U12362 (N_12362,N_12130,N_12183);
xnor U12363 (N_12363,N_12122,N_12285);
nand U12364 (N_12364,N_12041,N_12079);
or U12365 (N_12365,N_12037,N_12252);
xnor U12366 (N_12366,N_12062,N_12026);
or U12367 (N_12367,N_12287,N_12199);
xor U12368 (N_12368,N_12195,N_12168);
nor U12369 (N_12369,N_12230,N_12124);
or U12370 (N_12370,N_12191,N_12268);
or U12371 (N_12371,N_12172,N_12138);
nand U12372 (N_12372,N_12050,N_12267);
nor U12373 (N_12373,N_12208,N_12237);
nor U12374 (N_12374,N_12010,N_12278);
xor U12375 (N_12375,N_12165,N_12272);
nor U12376 (N_12376,N_12111,N_12188);
nor U12377 (N_12377,N_12086,N_12169);
or U12378 (N_12378,N_12110,N_12170);
nor U12379 (N_12379,N_12098,N_12249);
xnor U12380 (N_12380,N_12021,N_12228);
nand U12381 (N_12381,N_12002,N_12270);
and U12382 (N_12382,N_12248,N_12259);
or U12383 (N_12383,N_12150,N_12080);
or U12384 (N_12384,N_12055,N_12096);
nand U12385 (N_12385,N_12043,N_12206);
nand U12386 (N_12386,N_12060,N_12213);
and U12387 (N_12387,N_12244,N_12227);
xor U12388 (N_12388,N_12036,N_12288);
nor U12389 (N_12389,N_12291,N_12089);
nand U12390 (N_12390,N_12070,N_12094);
or U12391 (N_12391,N_12013,N_12216);
nand U12392 (N_12392,N_12121,N_12176);
and U12393 (N_12393,N_12120,N_12038);
nand U12394 (N_12394,N_12131,N_12133);
or U12395 (N_12395,N_12186,N_12018);
xnor U12396 (N_12396,N_12102,N_12118);
and U12397 (N_12397,N_12091,N_12044);
or U12398 (N_12398,N_12200,N_12142);
and U12399 (N_12399,N_12024,N_12296);
or U12400 (N_12400,N_12163,N_12239);
nand U12401 (N_12401,N_12240,N_12262);
nand U12402 (N_12402,N_12217,N_12047);
or U12403 (N_12403,N_12004,N_12105);
or U12404 (N_12404,N_12135,N_12221);
nor U12405 (N_12405,N_12196,N_12073);
nand U12406 (N_12406,N_12068,N_12204);
nand U12407 (N_12407,N_12030,N_12254);
nor U12408 (N_12408,N_12177,N_12283);
nand U12409 (N_12409,N_12231,N_12078);
or U12410 (N_12410,N_12189,N_12020);
nor U12411 (N_12411,N_12066,N_12201);
xnor U12412 (N_12412,N_12134,N_12007);
or U12413 (N_12413,N_12257,N_12076);
nand U12414 (N_12414,N_12149,N_12090);
nor U12415 (N_12415,N_12045,N_12097);
nor U12416 (N_12416,N_12048,N_12014);
nand U12417 (N_12417,N_12222,N_12215);
xnor U12418 (N_12418,N_12063,N_12100);
or U12419 (N_12419,N_12144,N_12008);
nand U12420 (N_12420,N_12059,N_12088);
nor U12421 (N_12421,N_12032,N_12093);
nand U12422 (N_12422,N_12185,N_12109);
or U12423 (N_12423,N_12234,N_12099);
and U12424 (N_12424,N_12253,N_12028);
xnor U12425 (N_12425,N_12049,N_12223);
xor U12426 (N_12426,N_12271,N_12235);
or U12427 (N_12427,N_12162,N_12293);
and U12428 (N_12428,N_12151,N_12040);
xnor U12429 (N_12429,N_12132,N_12280);
nand U12430 (N_12430,N_12295,N_12212);
and U12431 (N_12431,N_12128,N_12179);
and U12432 (N_12432,N_12214,N_12072);
nor U12433 (N_12433,N_12058,N_12232);
and U12434 (N_12434,N_12181,N_12274);
nand U12435 (N_12435,N_12139,N_12277);
xnor U12436 (N_12436,N_12273,N_12156);
nor U12437 (N_12437,N_12143,N_12029);
and U12438 (N_12438,N_12193,N_12137);
nor U12439 (N_12439,N_12074,N_12136);
xor U12440 (N_12440,N_12012,N_12245);
nand U12441 (N_12441,N_12255,N_12027);
or U12442 (N_12442,N_12025,N_12258);
or U12443 (N_12443,N_12054,N_12108);
xnor U12444 (N_12444,N_12243,N_12053);
and U12445 (N_12445,N_12117,N_12011);
or U12446 (N_12446,N_12051,N_12022);
and U12447 (N_12447,N_12034,N_12126);
and U12448 (N_12448,N_12261,N_12116);
nand U12449 (N_12449,N_12064,N_12187);
or U12450 (N_12450,N_12077,N_12237);
or U12451 (N_12451,N_12201,N_12245);
nor U12452 (N_12452,N_12267,N_12060);
and U12453 (N_12453,N_12132,N_12279);
xor U12454 (N_12454,N_12102,N_12235);
and U12455 (N_12455,N_12219,N_12108);
and U12456 (N_12456,N_12162,N_12069);
and U12457 (N_12457,N_12129,N_12210);
xnor U12458 (N_12458,N_12172,N_12102);
nor U12459 (N_12459,N_12263,N_12295);
xnor U12460 (N_12460,N_12041,N_12223);
nor U12461 (N_12461,N_12115,N_12286);
nor U12462 (N_12462,N_12225,N_12162);
nor U12463 (N_12463,N_12208,N_12138);
nand U12464 (N_12464,N_12062,N_12157);
xnor U12465 (N_12465,N_12078,N_12142);
or U12466 (N_12466,N_12069,N_12032);
and U12467 (N_12467,N_12230,N_12266);
and U12468 (N_12468,N_12259,N_12081);
xor U12469 (N_12469,N_12018,N_12264);
nand U12470 (N_12470,N_12203,N_12137);
nand U12471 (N_12471,N_12050,N_12091);
or U12472 (N_12472,N_12298,N_12255);
nand U12473 (N_12473,N_12063,N_12228);
or U12474 (N_12474,N_12284,N_12213);
nor U12475 (N_12475,N_12030,N_12057);
xnor U12476 (N_12476,N_12102,N_12031);
xor U12477 (N_12477,N_12236,N_12273);
or U12478 (N_12478,N_12066,N_12039);
xor U12479 (N_12479,N_12055,N_12270);
xor U12480 (N_12480,N_12276,N_12170);
and U12481 (N_12481,N_12056,N_12257);
nand U12482 (N_12482,N_12133,N_12262);
or U12483 (N_12483,N_12132,N_12135);
xnor U12484 (N_12484,N_12176,N_12080);
xnor U12485 (N_12485,N_12274,N_12075);
nand U12486 (N_12486,N_12017,N_12100);
nand U12487 (N_12487,N_12229,N_12233);
xnor U12488 (N_12488,N_12146,N_12280);
nand U12489 (N_12489,N_12197,N_12254);
nor U12490 (N_12490,N_12137,N_12204);
and U12491 (N_12491,N_12013,N_12263);
and U12492 (N_12492,N_12122,N_12171);
nor U12493 (N_12493,N_12157,N_12264);
and U12494 (N_12494,N_12014,N_12203);
and U12495 (N_12495,N_12189,N_12143);
and U12496 (N_12496,N_12128,N_12111);
nand U12497 (N_12497,N_12051,N_12238);
or U12498 (N_12498,N_12173,N_12066);
nand U12499 (N_12499,N_12200,N_12075);
nand U12500 (N_12500,N_12284,N_12021);
and U12501 (N_12501,N_12006,N_12190);
nand U12502 (N_12502,N_12027,N_12196);
or U12503 (N_12503,N_12209,N_12148);
xor U12504 (N_12504,N_12034,N_12099);
nor U12505 (N_12505,N_12204,N_12142);
nand U12506 (N_12506,N_12227,N_12110);
nor U12507 (N_12507,N_12031,N_12215);
or U12508 (N_12508,N_12077,N_12185);
xnor U12509 (N_12509,N_12173,N_12220);
nor U12510 (N_12510,N_12299,N_12120);
or U12511 (N_12511,N_12224,N_12060);
or U12512 (N_12512,N_12051,N_12218);
nand U12513 (N_12513,N_12001,N_12117);
nor U12514 (N_12514,N_12079,N_12075);
nor U12515 (N_12515,N_12020,N_12051);
xor U12516 (N_12516,N_12195,N_12154);
nor U12517 (N_12517,N_12249,N_12085);
or U12518 (N_12518,N_12271,N_12173);
nand U12519 (N_12519,N_12171,N_12124);
or U12520 (N_12520,N_12241,N_12195);
and U12521 (N_12521,N_12040,N_12173);
xnor U12522 (N_12522,N_12162,N_12027);
nand U12523 (N_12523,N_12280,N_12183);
or U12524 (N_12524,N_12146,N_12155);
or U12525 (N_12525,N_12183,N_12040);
and U12526 (N_12526,N_12136,N_12113);
and U12527 (N_12527,N_12205,N_12044);
nor U12528 (N_12528,N_12292,N_12067);
nor U12529 (N_12529,N_12287,N_12208);
nor U12530 (N_12530,N_12106,N_12187);
and U12531 (N_12531,N_12115,N_12134);
xor U12532 (N_12532,N_12193,N_12148);
and U12533 (N_12533,N_12067,N_12268);
nand U12534 (N_12534,N_12041,N_12199);
or U12535 (N_12535,N_12144,N_12248);
xnor U12536 (N_12536,N_12204,N_12260);
xor U12537 (N_12537,N_12269,N_12144);
nor U12538 (N_12538,N_12270,N_12236);
and U12539 (N_12539,N_12218,N_12029);
and U12540 (N_12540,N_12035,N_12052);
nand U12541 (N_12541,N_12055,N_12219);
nand U12542 (N_12542,N_12221,N_12018);
nand U12543 (N_12543,N_12131,N_12125);
xor U12544 (N_12544,N_12264,N_12139);
or U12545 (N_12545,N_12144,N_12089);
xnor U12546 (N_12546,N_12140,N_12089);
nand U12547 (N_12547,N_12278,N_12252);
xor U12548 (N_12548,N_12015,N_12218);
xor U12549 (N_12549,N_12040,N_12188);
and U12550 (N_12550,N_12028,N_12058);
nand U12551 (N_12551,N_12170,N_12098);
xnor U12552 (N_12552,N_12264,N_12138);
xnor U12553 (N_12553,N_12213,N_12002);
nor U12554 (N_12554,N_12148,N_12050);
and U12555 (N_12555,N_12072,N_12121);
or U12556 (N_12556,N_12035,N_12103);
nand U12557 (N_12557,N_12008,N_12113);
or U12558 (N_12558,N_12290,N_12194);
and U12559 (N_12559,N_12148,N_12132);
nor U12560 (N_12560,N_12087,N_12090);
nor U12561 (N_12561,N_12075,N_12231);
nor U12562 (N_12562,N_12244,N_12180);
nand U12563 (N_12563,N_12153,N_12104);
or U12564 (N_12564,N_12199,N_12172);
nor U12565 (N_12565,N_12089,N_12166);
or U12566 (N_12566,N_12164,N_12251);
xnor U12567 (N_12567,N_12046,N_12206);
and U12568 (N_12568,N_12172,N_12001);
or U12569 (N_12569,N_12158,N_12247);
xor U12570 (N_12570,N_12093,N_12242);
or U12571 (N_12571,N_12247,N_12280);
or U12572 (N_12572,N_12227,N_12273);
nor U12573 (N_12573,N_12265,N_12006);
or U12574 (N_12574,N_12162,N_12093);
xnor U12575 (N_12575,N_12175,N_12016);
and U12576 (N_12576,N_12049,N_12221);
xor U12577 (N_12577,N_12123,N_12146);
and U12578 (N_12578,N_12271,N_12132);
or U12579 (N_12579,N_12208,N_12133);
and U12580 (N_12580,N_12098,N_12077);
xor U12581 (N_12581,N_12286,N_12262);
nand U12582 (N_12582,N_12223,N_12244);
nand U12583 (N_12583,N_12098,N_12100);
or U12584 (N_12584,N_12057,N_12094);
xor U12585 (N_12585,N_12089,N_12102);
or U12586 (N_12586,N_12297,N_12288);
nand U12587 (N_12587,N_12213,N_12169);
nor U12588 (N_12588,N_12228,N_12208);
nor U12589 (N_12589,N_12192,N_12280);
or U12590 (N_12590,N_12065,N_12156);
or U12591 (N_12591,N_12199,N_12006);
xor U12592 (N_12592,N_12068,N_12148);
xor U12593 (N_12593,N_12169,N_12296);
and U12594 (N_12594,N_12072,N_12021);
nor U12595 (N_12595,N_12026,N_12215);
xor U12596 (N_12596,N_12053,N_12264);
or U12597 (N_12597,N_12013,N_12073);
nand U12598 (N_12598,N_12214,N_12252);
nand U12599 (N_12599,N_12009,N_12155);
nand U12600 (N_12600,N_12469,N_12549);
nor U12601 (N_12601,N_12455,N_12539);
nand U12602 (N_12602,N_12378,N_12457);
nor U12603 (N_12603,N_12490,N_12321);
nand U12604 (N_12604,N_12374,N_12421);
nor U12605 (N_12605,N_12325,N_12550);
xor U12606 (N_12606,N_12481,N_12564);
nand U12607 (N_12607,N_12470,N_12500);
nand U12608 (N_12608,N_12369,N_12530);
nor U12609 (N_12609,N_12551,N_12487);
and U12610 (N_12610,N_12473,N_12462);
xor U12611 (N_12611,N_12301,N_12568);
or U12612 (N_12612,N_12522,N_12498);
nand U12613 (N_12613,N_12366,N_12465);
or U12614 (N_12614,N_12414,N_12367);
nand U12615 (N_12615,N_12331,N_12453);
or U12616 (N_12616,N_12518,N_12589);
and U12617 (N_12617,N_12525,N_12488);
and U12618 (N_12618,N_12476,N_12506);
or U12619 (N_12619,N_12483,N_12359);
nand U12620 (N_12620,N_12489,N_12409);
nor U12621 (N_12621,N_12395,N_12358);
or U12622 (N_12622,N_12365,N_12531);
or U12623 (N_12623,N_12460,N_12461);
and U12624 (N_12624,N_12332,N_12338);
nand U12625 (N_12625,N_12327,N_12557);
and U12626 (N_12626,N_12424,N_12349);
xnor U12627 (N_12627,N_12334,N_12306);
nand U12628 (N_12628,N_12388,N_12527);
nand U12629 (N_12629,N_12423,N_12554);
nand U12630 (N_12630,N_12422,N_12428);
nor U12631 (N_12631,N_12593,N_12510);
nor U12632 (N_12632,N_12415,N_12363);
nor U12633 (N_12633,N_12380,N_12302);
nand U12634 (N_12634,N_12391,N_12492);
nor U12635 (N_12635,N_12537,N_12429);
nand U12636 (N_12636,N_12390,N_12376);
nor U12637 (N_12637,N_12373,N_12377);
nand U12638 (N_12638,N_12398,N_12571);
nand U12639 (N_12639,N_12532,N_12324);
nand U12640 (N_12640,N_12310,N_12574);
nor U12641 (N_12641,N_12472,N_12326);
nand U12642 (N_12642,N_12548,N_12355);
nand U12643 (N_12643,N_12406,N_12381);
or U12644 (N_12644,N_12573,N_12452);
nor U12645 (N_12645,N_12520,N_12512);
nor U12646 (N_12646,N_12405,N_12475);
and U12647 (N_12647,N_12439,N_12426);
nor U12648 (N_12648,N_12567,N_12482);
nand U12649 (N_12649,N_12508,N_12352);
and U12650 (N_12650,N_12474,N_12596);
xor U12651 (N_12651,N_12347,N_12552);
or U12652 (N_12652,N_12300,N_12434);
and U12653 (N_12653,N_12392,N_12467);
or U12654 (N_12654,N_12346,N_12497);
nand U12655 (N_12655,N_12372,N_12404);
nand U12656 (N_12656,N_12587,N_12572);
xnor U12657 (N_12657,N_12303,N_12307);
and U12658 (N_12658,N_12560,N_12534);
nand U12659 (N_12659,N_12353,N_12544);
nor U12660 (N_12660,N_12496,N_12480);
nor U12661 (N_12661,N_12595,N_12399);
or U12662 (N_12662,N_12581,N_12454);
or U12663 (N_12663,N_12533,N_12451);
xor U12664 (N_12664,N_12582,N_12420);
nor U12665 (N_12665,N_12316,N_12342);
and U12666 (N_12666,N_12456,N_12394);
xor U12667 (N_12667,N_12591,N_12408);
or U12668 (N_12668,N_12495,N_12562);
or U12669 (N_12669,N_12333,N_12553);
nand U12670 (N_12670,N_12511,N_12584);
xor U12671 (N_12671,N_12598,N_12412);
or U12672 (N_12672,N_12410,N_12578);
nand U12673 (N_12673,N_12370,N_12493);
nand U12674 (N_12674,N_12443,N_12330);
nor U12675 (N_12675,N_12559,N_12445);
nand U12676 (N_12676,N_12590,N_12328);
and U12677 (N_12677,N_12484,N_12385);
and U12678 (N_12678,N_12384,N_12393);
or U12679 (N_12679,N_12477,N_12516);
nand U12680 (N_12680,N_12466,N_12354);
nor U12681 (N_12681,N_12547,N_12304);
or U12682 (N_12682,N_12343,N_12463);
nor U12683 (N_12683,N_12526,N_12416);
xor U12684 (N_12684,N_12442,N_12535);
and U12685 (N_12685,N_12345,N_12397);
and U12686 (N_12686,N_12313,N_12323);
or U12687 (N_12687,N_12433,N_12305);
or U12688 (N_12688,N_12446,N_12309);
nand U12689 (N_12689,N_12543,N_12320);
or U12690 (N_12690,N_12371,N_12335);
xnor U12691 (N_12691,N_12386,N_12538);
and U12692 (N_12692,N_12440,N_12444);
or U12693 (N_12693,N_12382,N_12501);
nor U12694 (N_12694,N_12458,N_12566);
and U12695 (N_12695,N_12337,N_12364);
or U12696 (N_12696,N_12515,N_12485);
xnor U12697 (N_12697,N_12509,N_12569);
and U12698 (N_12698,N_12514,N_12565);
nor U12699 (N_12699,N_12494,N_12402);
and U12700 (N_12700,N_12479,N_12317);
nor U12701 (N_12701,N_12401,N_12585);
or U12702 (N_12702,N_12502,N_12417);
xnor U12703 (N_12703,N_12425,N_12503);
or U12704 (N_12704,N_12468,N_12464);
xor U12705 (N_12705,N_12312,N_12576);
nor U12706 (N_12706,N_12396,N_12579);
nand U12707 (N_12707,N_12308,N_12351);
and U12708 (N_12708,N_12383,N_12542);
xor U12709 (N_12709,N_12361,N_12450);
xnor U12710 (N_12710,N_12400,N_12314);
xor U12711 (N_12711,N_12430,N_12447);
nand U12712 (N_12712,N_12441,N_12389);
nand U12713 (N_12713,N_12563,N_12419);
xor U12714 (N_12714,N_12505,N_12586);
nor U12715 (N_12715,N_12592,N_12471);
nand U12716 (N_12716,N_12523,N_12362);
nor U12717 (N_12717,N_12491,N_12427);
nor U12718 (N_12718,N_12322,N_12379);
and U12719 (N_12719,N_12575,N_12448);
nand U12720 (N_12720,N_12555,N_12418);
nor U12721 (N_12721,N_12545,N_12329);
nand U12722 (N_12722,N_12340,N_12436);
xnor U12723 (N_12723,N_12594,N_12403);
xnor U12724 (N_12724,N_12577,N_12407);
nand U12725 (N_12725,N_12597,N_12517);
nor U12726 (N_12726,N_12524,N_12315);
nor U12727 (N_12727,N_12375,N_12319);
and U12728 (N_12728,N_12311,N_12536);
and U12729 (N_12729,N_12519,N_12387);
nand U12730 (N_12730,N_12504,N_12438);
nor U12731 (N_12731,N_12529,N_12558);
nor U12732 (N_12732,N_12318,N_12437);
or U12733 (N_12733,N_12507,N_12528);
or U12734 (N_12734,N_12348,N_12368);
xnor U12735 (N_12735,N_12341,N_12336);
and U12736 (N_12736,N_12459,N_12432);
and U12737 (N_12737,N_12513,N_12540);
and U12738 (N_12738,N_12478,N_12486);
nand U12739 (N_12739,N_12541,N_12546);
and U12740 (N_12740,N_12431,N_12521);
nor U12741 (N_12741,N_12360,N_12561);
xor U12742 (N_12742,N_12588,N_12350);
nand U12743 (N_12743,N_12583,N_12339);
xor U12744 (N_12744,N_12357,N_12356);
or U12745 (N_12745,N_12499,N_12411);
nand U12746 (N_12746,N_12599,N_12413);
nor U12747 (N_12747,N_12570,N_12580);
or U12748 (N_12748,N_12449,N_12344);
and U12749 (N_12749,N_12556,N_12435);
or U12750 (N_12750,N_12580,N_12451);
and U12751 (N_12751,N_12428,N_12415);
or U12752 (N_12752,N_12395,N_12345);
or U12753 (N_12753,N_12492,N_12576);
nor U12754 (N_12754,N_12565,N_12359);
or U12755 (N_12755,N_12583,N_12384);
or U12756 (N_12756,N_12449,N_12508);
xor U12757 (N_12757,N_12400,N_12338);
and U12758 (N_12758,N_12396,N_12470);
nor U12759 (N_12759,N_12326,N_12371);
nand U12760 (N_12760,N_12410,N_12363);
or U12761 (N_12761,N_12382,N_12340);
nand U12762 (N_12762,N_12331,N_12343);
or U12763 (N_12763,N_12429,N_12457);
xnor U12764 (N_12764,N_12592,N_12386);
and U12765 (N_12765,N_12543,N_12304);
nor U12766 (N_12766,N_12585,N_12533);
or U12767 (N_12767,N_12576,N_12466);
nor U12768 (N_12768,N_12440,N_12325);
or U12769 (N_12769,N_12516,N_12523);
xnor U12770 (N_12770,N_12527,N_12370);
xnor U12771 (N_12771,N_12521,N_12574);
and U12772 (N_12772,N_12569,N_12555);
nand U12773 (N_12773,N_12434,N_12488);
and U12774 (N_12774,N_12355,N_12494);
and U12775 (N_12775,N_12414,N_12433);
nor U12776 (N_12776,N_12596,N_12324);
nand U12777 (N_12777,N_12512,N_12530);
and U12778 (N_12778,N_12309,N_12367);
nor U12779 (N_12779,N_12316,N_12305);
or U12780 (N_12780,N_12437,N_12319);
nand U12781 (N_12781,N_12394,N_12303);
and U12782 (N_12782,N_12366,N_12317);
and U12783 (N_12783,N_12454,N_12584);
nor U12784 (N_12784,N_12325,N_12532);
and U12785 (N_12785,N_12543,N_12410);
nand U12786 (N_12786,N_12320,N_12519);
and U12787 (N_12787,N_12399,N_12497);
nor U12788 (N_12788,N_12383,N_12535);
and U12789 (N_12789,N_12593,N_12499);
and U12790 (N_12790,N_12357,N_12530);
nand U12791 (N_12791,N_12446,N_12490);
nor U12792 (N_12792,N_12571,N_12552);
nand U12793 (N_12793,N_12319,N_12540);
nor U12794 (N_12794,N_12457,N_12520);
xnor U12795 (N_12795,N_12390,N_12550);
xor U12796 (N_12796,N_12315,N_12591);
and U12797 (N_12797,N_12461,N_12455);
or U12798 (N_12798,N_12416,N_12567);
nor U12799 (N_12799,N_12571,N_12418);
and U12800 (N_12800,N_12363,N_12331);
nand U12801 (N_12801,N_12398,N_12465);
xnor U12802 (N_12802,N_12328,N_12355);
xnor U12803 (N_12803,N_12306,N_12521);
xnor U12804 (N_12804,N_12429,N_12337);
nand U12805 (N_12805,N_12357,N_12591);
nor U12806 (N_12806,N_12587,N_12332);
or U12807 (N_12807,N_12353,N_12425);
xnor U12808 (N_12808,N_12544,N_12515);
or U12809 (N_12809,N_12312,N_12543);
nand U12810 (N_12810,N_12369,N_12490);
or U12811 (N_12811,N_12473,N_12478);
and U12812 (N_12812,N_12388,N_12507);
nor U12813 (N_12813,N_12595,N_12315);
nor U12814 (N_12814,N_12374,N_12446);
nor U12815 (N_12815,N_12540,N_12464);
or U12816 (N_12816,N_12312,N_12421);
nor U12817 (N_12817,N_12479,N_12553);
and U12818 (N_12818,N_12366,N_12329);
xor U12819 (N_12819,N_12578,N_12460);
xnor U12820 (N_12820,N_12501,N_12321);
and U12821 (N_12821,N_12353,N_12438);
xnor U12822 (N_12822,N_12593,N_12451);
or U12823 (N_12823,N_12580,N_12351);
nor U12824 (N_12824,N_12549,N_12514);
and U12825 (N_12825,N_12349,N_12568);
or U12826 (N_12826,N_12405,N_12387);
xor U12827 (N_12827,N_12353,N_12595);
and U12828 (N_12828,N_12487,N_12519);
xnor U12829 (N_12829,N_12304,N_12408);
nor U12830 (N_12830,N_12358,N_12570);
nor U12831 (N_12831,N_12454,N_12532);
nand U12832 (N_12832,N_12360,N_12475);
nand U12833 (N_12833,N_12499,N_12304);
or U12834 (N_12834,N_12323,N_12332);
or U12835 (N_12835,N_12351,N_12379);
xnor U12836 (N_12836,N_12351,N_12585);
nand U12837 (N_12837,N_12351,N_12599);
and U12838 (N_12838,N_12416,N_12399);
and U12839 (N_12839,N_12322,N_12303);
xor U12840 (N_12840,N_12432,N_12430);
or U12841 (N_12841,N_12482,N_12446);
nor U12842 (N_12842,N_12513,N_12307);
and U12843 (N_12843,N_12398,N_12336);
nand U12844 (N_12844,N_12547,N_12444);
xnor U12845 (N_12845,N_12558,N_12538);
or U12846 (N_12846,N_12362,N_12486);
and U12847 (N_12847,N_12314,N_12507);
and U12848 (N_12848,N_12473,N_12569);
nand U12849 (N_12849,N_12404,N_12306);
nor U12850 (N_12850,N_12578,N_12588);
nor U12851 (N_12851,N_12535,N_12560);
xnor U12852 (N_12852,N_12381,N_12503);
xnor U12853 (N_12853,N_12332,N_12403);
and U12854 (N_12854,N_12506,N_12309);
xor U12855 (N_12855,N_12425,N_12431);
xnor U12856 (N_12856,N_12382,N_12418);
nor U12857 (N_12857,N_12410,N_12537);
nor U12858 (N_12858,N_12585,N_12417);
xnor U12859 (N_12859,N_12377,N_12439);
nand U12860 (N_12860,N_12383,N_12332);
or U12861 (N_12861,N_12573,N_12495);
nor U12862 (N_12862,N_12417,N_12338);
and U12863 (N_12863,N_12557,N_12319);
xor U12864 (N_12864,N_12474,N_12467);
nand U12865 (N_12865,N_12476,N_12459);
and U12866 (N_12866,N_12346,N_12303);
xor U12867 (N_12867,N_12558,N_12579);
xor U12868 (N_12868,N_12372,N_12473);
xnor U12869 (N_12869,N_12477,N_12550);
and U12870 (N_12870,N_12553,N_12444);
nand U12871 (N_12871,N_12419,N_12541);
xor U12872 (N_12872,N_12554,N_12523);
or U12873 (N_12873,N_12453,N_12462);
nor U12874 (N_12874,N_12387,N_12528);
nand U12875 (N_12875,N_12573,N_12346);
and U12876 (N_12876,N_12340,N_12431);
or U12877 (N_12877,N_12554,N_12364);
or U12878 (N_12878,N_12363,N_12349);
and U12879 (N_12879,N_12439,N_12531);
and U12880 (N_12880,N_12429,N_12495);
and U12881 (N_12881,N_12578,N_12481);
nor U12882 (N_12882,N_12473,N_12476);
and U12883 (N_12883,N_12579,N_12438);
or U12884 (N_12884,N_12355,N_12514);
xnor U12885 (N_12885,N_12317,N_12463);
or U12886 (N_12886,N_12520,N_12540);
nand U12887 (N_12887,N_12482,N_12301);
xnor U12888 (N_12888,N_12564,N_12540);
or U12889 (N_12889,N_12571,N_12337);
nand U12890 (N_12890,N_12383,N_12489);
and U12891 (N_12891,N_12320,N_12524);
nand U12892 (N_12892,N_12542,N_12529);
and U12893 (N_12893,N_12421,N_12368);
xor U12894 (N_12894,N_12472,N_12533);
xnor U12895 (N_12895,N_12358,N_12446);
nor U12896 (N_12896,N_12474,N_12415);
nor U12897 (N_12897,N_12344,N_12593);
or U12898 (N_12898,N_12522,N_12385);
and U12899 (N_12899,N_12507,N_12316);
xor U12900 (N_12900,N_12707,N_12631);
and U12901 (N_12901,N_12628,N_12764);
nand U12902 (N_12902,N_12886,N_12660);
xnor U12903 (N_12903,N_12852,N_12626);
or U12904 (N_12904,N_12804,N_12808);
and U12905 (N_12905,N_12622,N_12891);
and U12906 (N_12906,N_12895,N_12614);
nor U12907 (N_12907,N_12795,N_12755);
nor U12908 (N_12908,N_12676,N_12818);
nor U12909 (N_12909,N_12640,N_12790);
or U12910 (N_12910,N_12899,N_12772);
nor U12911 (N_12911,N_12604,N_12682);
or U12912 (N_12912,N_12815,N_12603);
xnor U12913 (N_12913,N_12620,N_12726);
nor U12914 (N_12914,N_12840,N_12885);
nand U12915 (N_12915,N_12865,N_12783);
nor U12916 (N_12916,N_12692,N_12624);
nor U12917 (N_12917,N_12735,N_12610);
xor U12918 (N_12918,N_12758,N_12711);
xor U12919 (N_12919,N_12847,N_12834);
nor U12920 (N_12920,N_12837,N_12722);
nand U12921 (N_12921,N_12831,N_12841);
nor U12922 (N_12922,N_12715,N_12752);
and U12923 (N_12923,N_12657,N_12663);
nor U12924 (N_12924,N_12756,N_12741);
nand U12925 (N_12925,N_12748,N_12613);
xor U12926 (N_12926,N_12661,N_12606);
xor U12927 (N_12927,N_12653,N_12777);
xor U12928 (N_12928,N_12646,N_12892);
nand U12929 (N_12929,N_12883,N_12778);
nand U12930 (N_12930,N_12800,N_12762);
nor U12931 (N_12931,N_12718,N_12680);
xnor U12932 (N_12932,N_12861,N_12890);
and U12933 (N_12933,N_12801,N_12671);
or U12934 (N_12934,N_12856,N_12759);
xor U12935 (N_12935,N_12706,N_12673);
or U12936 (N_12936,N_12807,N_12652);
nand U12937 (N_12937,N_12791,N_12686);
and U12938 (N_12938,N_12674,N_12814);
and U12939 (N_12939,N_12827,N_12785);
and U12940 (N_12940,N_12730,N_12789);
or U12941 (N_12941,N_12787,N_12727);
nor U12942 (N_12942,N_12630,N_12609);
nor U12943 (N_12943,N_12839,N_12881);
nand U12944 (N_12944,N_12702,N_12893);
xnor U12945 (N_12945,N_12643,N_12737);
xor U12946 (N_12946,N_12659,N_12802);
nand U12947 (N_12947,N_12869,N_12824);
or U12948 (N_12948,N_12894,N_12687);
nand U12949 (N_12949,N_12879,N_12838);
and U12950 (N_12950,N_12749,N_12782);
and U12951 (N_12951,N_12848,N_12829);
xnor U12952 (N_12952,N_12612,N_12708);
nor U12953 (N_12953,N_12705,N_12780);
and U12954 (N_12954,N_12880,N_12751);
and U12955 (N_12955,N_12898,N_12683);
xnor U12956 (N_12956,N_12863,N_12639);
and U12957 (N_12957,N_12832,N_12700);
and U12958 (N_12958,N_12719,N_12849);
or U12959 (N_12959,N_12689,N_12621);
nor U12960 (N_12960,N_12773,N_12792);
nand U12961 (N_12961,N_12647,N_12862);
or U12962 (N_12962,N_12623,N_12677);
or U12963 (N_12963,N_12732,N_12658);
nor U12964 (N_12964,N_12878,N_12638);
nand U12965 (N_12965,N_12618,N_12828);
or U12966 (N_12966,N_12889,N_12876);
nand U12967 (N_12967,N_12798,N_12654);
nor U12968 (N_12968,N_12636,N_12884);
xnor U12969 (N_12969,N_12794,N_12655);
and U12970 (N_12970,N_12611,N_12854);
xor U12971 (N_12971,N_12864,N_12701);
or U12972 (N_12972,N_12750,N_12836);
and U12973 (N_12973,N_12691,N_12743);
nand U12974 (N_12974,N_12601,N_12786);
or U12975 (N_12975,N_12738,N_12816);
and U12976 (N_12976,N_12681,N_12775);
and U12977 (N_12977,N_12767,N_12627);
and U12978 (N_12978,N_12810,N_12757);
or U12979 (N_12979,N_12799,N_12615);
and U12980 (N_12980,N_12742,N_12670);
or U12981 (N_12981,N_12820,N_12779);
and U12982 (N_12982,N_12608,N_12728);
or U12983 (N_12983,N_12872,N_12843);
xor U12984 (N_12984,N_12760,N_12733);
nor U12985 (N_12985,N_12853,N_12695);
or U12986 (N_12986,N_12684,N_12678);
or U12987 (N_12987,N_12712,N_12888);
nand U12988 (N_12988,N_12859,N_12747);
or U12989 (N_12989,N_12835,N_12897);
nand U12990 (N_12990,N_12641,N_12716);
nand U12991 (N_12991,N_12868,N_12887);
xnor U12992 (N_12992,N_12871,N_12817);
and U12993 (N_12993,N_12664,N_12704);
or U12994 (N_12994,N_12870,N_12720);
xor U12995 (N_12995,N_12635,N_12809);
nor U12996 (N_12996,N_12826,N_12784);
nand U12997 (N_12997,N_12731,N_12693);
xor U12998 (N_12998,N_12896,N_12629);
nand U12999 (N_12999,N_12637,N_12830);
nand U13000 (N_13000,N_12698,N_12617);
nand U13001 (N_13001,N_12768,N_12644);
and U13002 (N_13002,N_12648,N_12668);
nor U13003 (N_13003,N_12746,N_12781);
nand U13004 (N_13004,N_12665,N_12669);
nand U13005 (N_13005,N_12844,N_12600);
xor U13006 (N_13006,N_12855,N_12806);
and U13007 (N_13007,N_12619,N_12717);
nor U13008 (N_13008,N_12822,N_12607);
and U13009 (N_13009,N_12703,N_12873);
xor U13010 (N_13010,N_12770,N_12845);
nand U13011 (N_13011,N_12874,N_12788);
nor U13012 (N_13012,N_12723,N_12709);
xnor U13013 (N_13013,N_12833,N_12763);
nand U13014 (N_13014,N_12725,N_12714);
nand U13015 (N_13015,N_12846,N_12666);
nand U13016 (N_13016,N_12649,N_12651);
nand U13017 (N_13017,N_12688,N_12805);
nor U13018 (N_13018,N_12690,N_12823);
nand U13019 (N_13019,N_12821,N_12744);
nand U13020 (N_13020,N_12813,N_12616);
xor U13021 (N_13021,N_12721,N_12662);
or U13022 (N_13022,N_12858,N_12685);
nand U13023 (N_13023,N_12882,N_12875);
nand U13024 (N_13024,N_12645,N_12739);
and U13025 (N_13025,N_12797,N_12656);
nor U13026 (N_13026,N_12851,N_12860);
and U13027 (N_13027,N_12753,N_12867);
nor U13028 (N_13028,N_12632,N_12602);
nand U13029 (N_13029,N_12771,N_12825);
nand U13030 (N_13030,N_12605,N_12774);
or U13031 (N_13031,N_12672,N_12625);
xnor U13032 (N_13032,N_12745,N_12811);
nor U13033 (N_13033,N_12812,N_12857);
nor U13034 (N_13034,N_12633,N_12766);
and U13035 (N_13035,N_12769,N_12729);
nor U13036 (N_13036,N_12713,N_12761);
nor U13037 (N_13037,N_12877,N_12710);
xnor U13038 (N_13038,N_12765,N_12850);
and U13039 (N_13039,N_12694,N_12740);
nor U13040 (N_13040,N_12803,N_12724);
and U13041 (N_13041,N_12699,N_12842);
nor U13042 (N_13042,N_12634,N_12696);
and U13043 (N_13043,N_12734,N_12697);
or U13044 (N_13044,N_12819,N_12642);
or U13045 (N_13045,N_12675,N_12667);
nor U13046 (N_13046,N_12776,N_12866);
nor U13047 (N_13047,N_12754,N_12796);
xor U13048 (N_13048,N_12793,N_12650);
and U13049 (N_13049,N_12679,N_12736);
or U13050 (N_13050,N_12871,N_12619);
nor U13051 (N_13051,N_12728,N_12627);
and U13052 (N_13052,N_12854,N_12619);
and U13053 (N_13053,N_12690,N_12636);
xor U13054 (N_13054,N_12609,N_12724);
nand U13055 (N_13055,N_12849,N_12679);
nand U13056 (N_13056,N_12856,N_12802);
nor U13057 (N_13057,N_12867,N_12787);
xor U13058 (N_13058,N_12791,N_12777);
or U13059 (N_13059,N_12633,N_12677);
and U13060 (N_13060,N_12738,N_12656);
or U13061 (N_13061,N_12880,N_12853);
nor U13062 (N_13062,N_12862,N_12878);
or U13063 (N_13063,N_12621,N_12615);
nand U13064 (N_13064,N_12756,N_12681);
and U13065 (N_13065,N_12844,N_12629);
or U13066 (N_13066,N_12811,N_12722);
or U13067 (N_13067,N_12637,N_12880);
nor U13068 (N_13068,N_12669,N_12867);
or U13069 (N_13069,N_12655,N_12656);
or U13070 (N_13070,N_12703,N_12807);
nand U13071 (N_13071,N_12775,N_12776);
nor U13072 (N_13072,N_12676,N_12733);
nor U13073 (N_13073,N_12813,N_12666);
nor U13074 (N_13074,N_12794,N_12723);
xnor U13075 (N_13075,N_12638,N_12736);
and U13076 (N_13076,N_12627,N_12825);
and U13077 (N_13077,N_12682,N_12635);
xor U13078 (N_13078,N_12789,N_12817);
xnor U13079 (N_13079,N_12740,N_12878);
nand U13080 (N_13080,N_12765,N_12712);
or U13081 (N_13081,N_12897,N_12630);
xnor U13082 (N_13082,N_12659,N_12830);
nand U13083 (N_13083,N_12677,N_12896);
nor U13084 (N_13084,N_12647,N_12693);
or U13085 (N_13085,N_12871,N_12621);
nand U13086 (N_13086,N_12891,N_12627);
xnor U13087 (N_13087,N_12683,N_12778);
nand U13088 (N_13088,N_12848,N_12662);
and U13089 (N_13089,N_12867,N_12875);
xnor U13090 (N_13090,N_12877,N_12799);
nor U13091 (N_13091,N_12603,N_12742);
nor U13092 (N_13092,N_12629,N_12741);
nor U13093 (N_13093,N_12881,N_12890);
xor U13094 (N_13094,N_12751,N_12808);
nand U13095 (N_13095,N_12801,N_12822);
and U13096 (N_13096,N_12736,N_12772);
and U13097 (N_13097,N_12772,N_12882);
nand U13098 (N_13098,N_12828,N_12851);
and U13099 (N_13099,N_12877,N_12683);
nand U13100 (N_13100,N_12663,N_12612);
nor U13101 (N_13101,N_12750,N_12603);
xor U13102 (N_13102,N_12799,N_12821);
xor U13103 (N_13103,N_12795,N_12736);
or U13104 (N_13104,N_12624,N_12651);
and U13105 (N_13105,N_12765,N_12793);
xnor U13106 (N_13106,N_12847,N_12626);
xor U13107 (N_13107,N_12765,N_12835);
nor U13108 (N_13108,N_12699,N_12828);
nor U13109 (N_13109,N_12600,N_12706);
or U13110 (N_13110,N_12767,N_12625);
or U13111 (N_13111,N_12710,N_12752);
or U13112 (N_13112,N_12707,N_12838);
nor U13113 (N_13113,N_12878,N_12886);
nor U13114 (N_13114,N_12712,N_12754);
xor U13115 (N_13115,N_12714,N_12739);
nor U13116 (N_13116,N_12684,N_12732);
xnor U13117 (N_13117,N_12701,N_12609);
nor U13118 (N_13118,N_12624,N_12824);
nand U13119 (N_13119,N_12646,N_12722);
xnor U13120 (N_13120,N_12738,N_12871);
xor U13121 (N_13121,N_12717,N_12792);
xor U13122 (N_13122,N_12680,N_12880);
nor U13123 (N_13123,N_12811,N_12794);
and U13124 (N_13124,N_12605,N_12852);
nor U13125 (N_13125,N_12734,N_12833);
nor U13126 (N_13126,N_12773,N_12879);
xnor U13127 (N_13127,N_12655,N_12601);
or U13128 (N_13128,N_12832,N_12636);
xnor U13129 (N_13129,N_12623,N_12819);
or U13130 (N_13130,N_12620,N_12769);
xor U13131 (N_13131,N_12640,N_12888);
xnor U13132 (N_13132,N_12632,N_12803);
xnor U13133 (N_13133,N_12668,N_12878);
or U13134 (N_13134,N_12694,N_12665);
xor U13135 (N_13135,N_12825,N_12648);
and U13136 (N_13136,N_12696,N_12757);
nor U13137 (N_13137,N_12792,N_12779);
and U13138 (N_13138,N_12864,N_12806);
or U13139 (N_13139,N_12610,N_12813);
or U13140 (N_13140,N_12843,N_12712);
and U13141 (N_13141,N_12870,N_12782);
nand U13142 (N_13142,N_12803,N_12870);
nand U13143 (N_13143,N_12885,N_12787);
xnor U13144 (N_13144,N_12654,N_12645);
xor U13145 (N_13145,N_12851,N_12730);
nor U13146 (N_13146,N_12686,N_12644);
and U13147 (N_13147,N_12858,N_12662);
xnor U13148 (N_13148,N_12778,N_12679);
nand U13149 (N_13149,N_12861,N_12664);
nor U13150 (N_13150,N_12775,N_12772);
or U13151 (N_13151,N_12759,N_12662);
nor U13152 (N_13152,N_12755,N_12729);
or U13153 (N_13153,N_12684,N_12751);
nand U13154 (N_13154,N_12673,N_12884);
nand U13155 (N_13155,N_12639,N_12651);
or U13156 (N_13156,N_12894,N_12699);
nand U13157 (N_13157,N_12802,N_12656);
xor U13158 (N_13158,N_12797,N_12821);
nand U13159 (N_13159,N_12611,N_12813);
nand U13160 (N_13160,N_12682,N_12693);
nor U13161 (N_13161,N_12733,N_12648);
xnor U13162 (N_13162,N_12709,N_12863);
or U13163 (N_13163,N_12642,N_12705);
xnor U13164 (N_13164,N_12707,N_12649);
xor U13165 (N_13165,N_12888,N_12730);
and U13166 (N_13166,N_12663,N_12815);
nor U13167 (N_13167,N_12779,N_12629);
xnor U13168 (N_13168,N_12791,N_12622);
or U13169 (N_13169,N_12794,N_12848);
or U13170 (N_13170,N_12856,N_12610);
xnor U13171 (N_13171,N_12649,N_12710);
nor U13172 (N_13172,N_12621,N_12821);
xor U13173 (N_13173,N_12611,N_12651);
or U13174 (N_13174,N_12785,N_12820);
or U13175 (N_13175,N_12839,N_12844);
xnor U13176 (N_13176,N_12893,N_12750);
nand U13177 (N_13177,N_12689,N_12718);
xnor U13178 (N_13178,N_12868,N_12731);
xnor U13179 (N_13179,N_12795,N_12698);
xnor U13180 (N_13180,N_12887,N_12734);
xor U13181 (N_13181,N_12863,N_12833);
or U13182 (N_13182,N_12718,N_12628);
nor U13183 (N_13183,N_12629,N_12859);
nand U13184 (N_13184,N_12878,N_12864);
nand U13185 (N_13185,N_12604,N_12673);
xnor U13186 (N_13186,N_12766,N_12621);
or U13187 (N_13187,N_12790,N_12683);
nor U13188 (N_13188,N_12726,N_12729);
nor U13189 (N_13189,N_12636,N_12817);
nand U13190 (N_13190,N_12651,N_12723);
xor U13191 (N_13191,N_12856,N_12734);
or U13192 (N_13192,N_12869,N_12750);
nor U13193 (N_13193,N_12818,N_12836);
xnor U13194 (N_13194,N_12639,N_12797);
nor U13195 (N_13195,N_12767,N_12817);
or U13196 (N_13196,N_12837,N_12616);
or U13197 (N_13197,N_12760,N_12794);
or U13198 (N_13198,N_12659,N_12871);
nor U13199 (N_13199,N_12847,N_12686);
xnor U13200 (N_13200,N_13181,N_13035);
or U13201 (N_13201,N_13177,N_13024);
nor U13202 (N_13202,N_13139,N_13016);
or U13203 (N_13203,N_13040,N_13014);
nor U13204 (N_13204,N_13055,N_13013);
nor U13205 (N_13205,N_13087,N_13146);
nor U13206 (N_13206,N_13086,N_12993);
and U13207 (N_13207,N_12979,N_12932);
nand U13208 (N_13208,N_12971,N_13007);
or U13209 (N_13209,N_13187,N_12915);
xnor U13210 (N_13210,N_12918,N_13053);
or U13211 (N_13211,N_13073,N_13160);
and U13212 (N_13212,N_12942,N_13039);
and U13213 (N_13213,N_12927,N_13030);
xor U13214 (N_13214,N_13197,N_13151);
and U13215 (N_13215,N_12934,N_12998);
nand U13216 (N_13216,N_13095,N_13071);
or U13217 (N_13217,N_13033,N_12951);
or U13218 (N_13218,N_12945,N_12995);
xor U13219 (N_13219,N_12969,N_12909);
nor U13220 (N_13220,N_13064,N_13079);
and U13221 (N_13221,N_13198,N_13162);
nand U13222 (N_13222,N_12923,N_12962);
nor U13223 (N_13223,N_13001,N_13005);
nor U13224 (N_13224,N_13124,N_13043);
or U13225 (N_13225,N_12968,N_13034);
and U13226 (N_13226,N_13131,N_13165);
and U13227 (N_13227,N_13117,N_13057);
xor U13228 (N_13228,N_13076,N_13004);
nand U13229 (N_13229,N_13061,N_13130);
or U13230 (N_13230,N_12977,N_13152);
and U13231 (N_13231,N_13107,N_13120);
nand U13232 (N_13232,N_13183,N_12978);
xor U13233 (N_13233,N_13171,N_13099);
and U13234 (N_13234,N_13068,N_13052);
nand U13235 (N_13235,N_12950,N_12939);
nand U13236 (N_13236,N_13191,N_13047);
nand U13237 (N_13237,N_12988,N_13142);
nor U13238 (N_13238,N_13137,N_12958);
xor U13239 (N_13239,N_13159,N_13116);
nand U13240 (N_13240,N_13140,N_13077);
nor U13241 (N_13241,N_13048,N_13075);
xnor U13242 (N_13242,N_12999,N_13050);
and U13243 (N_13243,N_13002,N_13155);
or U13244 (N_13244,N_13037,N_13065);
nand U13245 (N_13245,N_12965,N_13062);
nand U13246 (N_13246,N_13009,N_13018);
xor U13247 (N_13247,N_13031,N_13106);
xnor U13248 (N_13248,N_12912,N_12952);
xnor U13249 (N_13249,N_12926,N_13179);
nand U13250 (N_13250,N_12928,N_13006);
or U13251 (N_13251,N_13168,N_12982);
or U13252 (N_13252,N_13122,N_12957);
or U13253 (N_13253,N_12960,N_13022);
or U13254 (N_13254,N_13025,N_13083);
nand U13255 (N_13255,N_13127,N_12986);
nand U13256 (N_13256,N_13172,N_13104);
nor U13257 (N_13257,N_13167,N_13113);
xnor U13258 (N_13258,N_13185,N_12910);
nand U13259 (N_13259,N_12984,N_12976);
xnor U13260 (N_13260,N_13153,N_13145);
nor U13261 (N_13261,N_12930,N_12916);
or U13262 (N_13262,N_13056,N_12966);
nor U13263 (N_13263,N_13119,N_13192);
and U13264 (N_13264,N_13150,N_13103);
nor U13265 (N_13265,N_12944,N_12992);
nand U13266 (N_13266,N_13045,N_12963);
nor U13267 (N_13267,N_13149,N_13134);
nand U13268 (N_13268,N_13060,N_13147);
nor U13269 (N_13269,N_13015,N_13078);
xor U13270 (N_13270,N_13136,N_13123);
nor U13271 (N_13271,N_13058,N_13108);
or U13272 (N_13272,N_13036,N_12972);
nand U13273 (N_13273,N_13190,N_12900);
or U13274 (N_13274,N_13161,N_13020);
nor U13275 (N_13275,N_12975,N_12996);
nor U13276 (N_13276,N_12991,N_12953);
nor U13277 (N_13277,N_13012,N_12905);
nand U13278 (N_13278,N_13118,N_13148);
nand U13279 (N_13279,N_12941,N_13041);
or U13280 (N_13280,N_13070,N_12907);
nand U13281 (N_13281,N_13189,N_12921);
nor U13282 (N_13282,N_13038,N_13084);
xnor U13283 (N_13283,N_13135,N_13098);
xnor U13284 (N_13284,N_13169,N_13000);
nand U13285 (N_13285,N_12908,N_13097);
nand U13286 (N_13286,N_13184,N_13042);
nand U13287 (N_13287,N_12987,N_13112);
or U13288 (N_13288,N_12917,N_12985);
nor U13289 (N_13289,N_13173,N_13125);
nor U13290 (N_13290,N_13069,N_12906);
nor U13291 (N_13291,N_12901,N_13046);
or U13292 (N_13292,N_12911,N_12955);
nand U13293 (N_13293,N_13128,N_13132);
nor U13294 (N_13294,N_12981,N_13074);
or U13295 (N_13295,N_12937,N_13182);
xnor U13296 (N_13296,N_13094,N_12938);
nand U13297 (N_13297,N_12936,N_12925);
nand U13298 (N_13298,N_13011,N_13089);
nand U13299 (N_13299,N_12959,N_13017);
nand U13300 (N_13300,N_12980,N_13054);
and U13301 (N_13301,N_13010,N_13032);
nand U13302 (N_13302,N_13141,N_13059);
and U13303 (N_13303,N_13195,N_13114);
nand U13304 (N_13304,N_13003,N_13144);
and U13305 (N_13305,N_12913,N_13157);
nand U13306 (N_13306,N_13090,N_13143);
xnor U13307 (N_13307,N_13170,N_13029);
xor U13308 (N_13308,N_13110,N_13067);
nor U13309 (N_13309,N_13111,N_13180);
and U13310 (N_13310,N_13164,N_12947);
nor U13311 (N_13311,N_13027,N_13166);
or U13312 (N_13312,N_13028,N_13008);
xor U13313 (N_13313,N_13115,N_12940);
nor U13314 (N_13314,N_13093,N_13019);
nor U13315 (N_13315,N_13080,N_12997);
or U13316 (N_13316,N_12954,N_13105);
nor U13317 (N_13317,N_13178,N_13063);
nand U13318 (N_13318,N_13156,N_13081);
or U13319 (N_13319,N_13158,N_13129);
nand U13320 (N_13320,N_12989,N_13051);
nand U13321 (N_13321,N_13023,N_13121);
nand U13322 (N_13322,N_13138,N_12920);
xnor U13323 (N_13323,N_12956,N_13026);
and U13324 (N_13324,N_13193,N_12902);
or U13325 (N_13325,N_12943,N_12961);
xor U13326 (N_13326,N_13186,N_13092);
nor U13327 (N_13327,N_13088,N_13072);
nor U13328 (N_13328,N_12929,N_13102);
nand U13329 (N_13329,N_13100,N_13196);
nand U13330 (N_13330,N_13085,N_12919);
nand U13331 (N_13331,N_13154,N_12946);
nor U13332 (N_13332,N_13163,N_13101);
nor U13333 (N_13333,N_12973,N_13188);
xor U13334 (N_13334,N_12994,N_13082);
or U13335 (N_13335,N_12967,N_12935);
and U13336 (N_13336,N_12983,N_13096);
or U13337 (N_13337,N_12949,N_12974);
and U13338 (N_13338,N_12964,N_13109);
or U13339 (N_13339,N_12931,N_12948);
or U13340 (N_13340,N_12922,N_13049);
or U13341 (N_13341,N_12903,N_13199);
nor U13342 (N_13342,N_13176,N_13133);
and U13343 (N_13343,N_13194,N_13021);
and U13344 (N_13344,N_12970,N_13091);
nor U13345 (N_13345,N_12914,N_13044);
nor U13346 (N_13346,N_13175,N_12933);
or U13347 (N_13347,N_12924,N_12990);
xnor U13348 (N_13348,N_13126,N_13066);
nor U13349 (N_13349,N_13174,N_12904);
and U13350 (N_13350,N_13160,N_13169);
xor U13351 (N_13351,N_12953,N_13172);
nor U13352 (N_13352,N_13083,N_13156);
nand U13353 (N_13353,N_12995,N_13167);
nor U13354 (N_13354,N_13114,N_12950);
or U13355 (N_13355,N_12941,N_13003);
or U13356 (N_13356,N_13158,N_12956);
nor U13357 (N_13357,N_13071,N_13190);
and U13358 (N_13358,N_13187,N_12941);
or U13359 (N_13359,N_13026,N_13138);
xor U13360 (N_13360,N_13035,N_12909);
nor U13361 (N_13361,N_12979,N_12978);
xor U13362 (N_13362,N_13017,N_13196);
nand U13363 (N_13363,N_12984,N_13173);
nand U13364 (N_13364,N_12954,N_13066);
or U13365 (N_13365,N_13005,N_13034);
nor U13366 (N_13366,N_13182,N_13053);
xnor U13367 (N_13367,N_13130,N_12920);
or U13368 (N_13368,N_13098,N_13053);
and U13369 (N_13369,N_13137,N_13101);
xor U13370 (N_13370,N_13001,N_13045);
and U13371 (N_13371,N_13082,N_13058);
nand U13372 (N_13372,N_13090,N_13058);
nand U13373 (N_13373,N_13109,N_13006);
nand U13374 (N_13374,N_13118,N_13003);
or U13375 (N_13375,N_12938,N_13124);
nand U13376 (N_13376,N_12998,N_12997);
and U13377 (N_13377,N_13112,N_13085);
or U13378 (N_13378,N_13032,N_13013);
nand U13379 (N_13379,N_13060,N_12929);
or U13380 (N_13380,N_13044,N_13039);
xor U13381 (N_13381,N_13125,N_12953);
xnor U13382 (N_13382,N_13145,N_12975);
or U13383 (N_13383,N_13057,N_12937);
xor U13384 (N_13384,N_12931,N_12940);
or U13385 (N_13385,N_13147,N_13167);
nor U13386 (N_13386,N_13042,N_12902);
xnor U13387 (N_13387,N_13107,N_13159);
nand U13388 (N_13388,N_12971,N_13075);
nand U13389 (N_13389,N_13168,N_13078);
xnor U13390 (N_13390,N_13047,N_12906);
nor U13391 (N_13391,N_12994,N_13058);
nor U13392 (N_13392,N_13006,N_13082);
or U13393 (N_13393,N_12989,N_13056);
nand U13394 (N_13394,N_13017,N_12929);
and U13395 (N_13395,N_13051,N_12929);
or U13396 (N_13396,N_13153,N_12965);
nor U13397 (N_13397,N_13056,N_12940);
nor U13398 (N_13398,N_12924,N_13138);
or U13399 (N_13399,N_12977,N_12945);
nor U13400 (N_13400,N_13006,N_13146);
xnor U13401 (N_13401,N_12950,N_13053);
nand U13402 (N_13402,N_13173,N_13101);
xor U13403 (N_13403,N_12992,N_13038);
and U13404 (N_13404,N_13117,N_12919);
xor U13405 (N_13405,N_12988,N_12992);
nand U13406 (N_13406,N_13012,N_13105);
nand U13407 (N_13407,N_13111,N_13198);
nor U13408 (N_13408,N_13158,N_13066);
and U13409 (N_13409,N_13009,N_13032);
or U13410 (N_13410,N_13170,N_13026);
xor U13411 (N_13411,N_13023,N_13177);
and U13412 (N_13412,N_13089,N_13130);
and U13413 (N_13413,N_13018,N_13174);
nand U13414 (N_13414,N_12980,N_13052);
and U13415 (N_13415,N_13124,N_13084);
nor U13416 (N_13416,N_13114,N_12985);
nor U13417 (N_13417,N_12952,N_12949);
nand U13418 (N_13418,N_12900,N_13130);
or U13419 (N_13419,N_12959,N_13060);
nor U13420 (N_13420,N_13110,N_12912);
nand U13421 (N_13421,N_13006,N_13115);
or U13422 (N_13422,N_13098,N_13178);
or U13423 (N_13423,N_12997,N_13061);
and U13424 (N_13424,N_12982,N_13133);
or U13425 (N_13425,N_13013,N_13064);
nand U13426 (N_13426,N_13017,N_13105);
nor U13427 (N_13427,N_13055,N_13163);
nor U13428 (N_13428,N_13175,N_12956);
and U13429 (N_13429,N_13083,N_13054);
nand U13430 (N_13430,N_13101,N_13148);
or U13431 (N_13431,N_13019,N_13097);
xor U13432 (N_13432,N_12940,N_12915);
and U13433 (N_13433,N_13188,N_13160);
or U13434 (N_13434,N_12910,N_13127);
nand U13435 (N_13435,N_13003,N_12927);
nand U13436 (N_13436,N_12930,N_12912);
and U13437 (N_13437,N_13023,N_13008);
xor U13438 (N_13438,N_13106,N_13119);
nor U13439 (N_13439,N_13142,N_13067);
nor U13440 (N_13440,N_13163,N_13133);
nor U13441 (N_13441,N_13140,N_13180);
or U13442 (N_13442,N_12910,N_13116);
and U13443 (N_13443,N_13016,N_12935);
nand U13444 (N_13444,N_12995,N_13079);
xor U13445 (N_13445,N_13192,N_12947);
xnor U13446 (N_13446,N_13191,N_13196);
xor U13447 (N_13447,N_12975,N_13167);
or U13448 (N_13448,N_13088,N_13103);
nand U13449 (N_13449,N_13112,N_13126);
or U13450 (N_13450,N_13190,N_12971);
or U13451 (N_13451,N_13057,N_13142);
or U13452 (N_13452,N_12924,N_12963);
or U13453 (N_13453,N_13175,N_12903);
or U13454 (N_13454,N_13059,N_12987);
or U13455 (N_13455,N_13175,N_13131);
and U13456 (N_13456,N_13124,N_13082);
xor U13457 (N_13457,N_13190,N_13077);
and U13458 (N_13458,N_12938,N_13102);
and U13459 (N_13459,N_13110,N_12986);
nand U13460 (N_13460,N_13053,N_13171);
or U13461 (N_13461,N_13165,N_13054);
and U13462 (N_13462,N_13050,N_12962);
nand U13463 (N_13463,N_13039,N_13178);
nand U13464 (N_13464,N_12958,N_13015);
nor U13465 (N_13465,N_13163,N_12912);
nor U13466 (N_13466,N_13108,N_13003);
nand U13467 (N_13467,N_13197,N_13147);
or U13468 (N_13468,N_13168,N_13147);
or U13469 (N_13469,N_12983,N_13045);
and U13470 (N_13470,N_13163,N_13075);
and U13471 (N_13471,N_13130,N_13164);
or U13472 (N_13472,N_13173,N_13053);
xnor U13473 (N_13473,N_13000,N_12905);
or U13474 (N_13474,N_13131,N_12999);
or U13475 (N_13475,N_13133,N_13178);
or U13476 (N_13476,N_12925,N_13182);
nor U13477 (N_13477,N_13165,N_13020);
and U13478 (N_13478,N_13039,N_12901);
xnor U13479 (N_13479,N_12925,N_13106);
nor U13480 (N_13480,N_12969,N_13105);
xor U13481 (N_13481,N_12917,N_12979);
or U13482 (N_13482,N_13170,N_13095);
xnor U13483 (N_13483,N_12901,N_12950);
xor U13484 (N_13484,N_13111,N_13079);
nor U13485 (N_13485,N_12914,N_12959);
nor U13486 (N_13486,N_12904,N_12921);
or U13487 (N_13487,N_12930,N_12913);
or U13488 (N_13488,N_12951,N_13079);
or U13489 (N_13489,N_13165,N_13137);
nand U13490 (N_13490,N_13136,N_13149);
xor U13491 (N_13491,N_13161,N_13090);
and U13492 (N_13492,N_13012,N_12982);
and U13493 (N_13493,N_13091,N_12916);
or U13494 (N_13494,N_12977,N_12912);
or U13495 (N_13495,N_13069,N_13042);
and U13496 (N_13496,N_13029,N_13106);
nor U13497 (N_13497,N_13133,N_12952);
or U13498 (N_13498,N_12998,N_12925);
nor U13499 (N_13499,N_12963,N_12942);
nand U13500 (N_13500,N_13365,N_13479);
and U13501 (N_13501,N_13347,N_13370);
or U13502 (N_13502,N_13230,N_13249);
nand U13503 (N_13503,N_13383,N_13407);
xor U13504 (N_13504,N_13462,N_13257);
nand U13505 (N_13505,N_13281,N_13367);
xnor U13506 (N_13506,N_13314,N_13375);
or U13507 (N_13507,N_13282,N_13286);
and U13508 (N_13508,N_13266,N_13213);
or U13509 (N_13509,N_13467,N_13497);
or U13510 (N_13510,N_13487,N_13481);
xnor U13511 (N_13511,N_13373,N_13469);
or U13512 (N_13512,N_13260,N_13341);
and U13513 (N_13513,N_13325,N_13237);
nor U13514 (N_13514,N_13490,N_13466);
or U13515 (N_13515,N_13381,N_13312);
xnor U13516 (N_13516,N_13356,N_13328);
nand U13517 (N_13517,N_13430,N_13436);
nand U13518 (N_13518,N_13464,N_13399);
nor U13519 (N_13519,N_13372,N_13216);
or U13520 (N_13520,N_13321,N_13387);
nor U13521 (N_13521,N_13425,N_13359);
and U13522 (N_13522,N_13262,N_13404);
nor U13523 (N_13523,N_13461,N_13374);
xor U13524 (N_13524,N_13258,N_13444);
or U13525 (N_13525,N_13343,N_13491);
and U13526 (N_13526,N_13248,N_13412);
nand U13527 (N_13527,N_13360,N_13364);
nor U13528 (N_13528,N_13468,N_13437);
and U13529 (N_13529,N_13303,N_13219);
nand U13530 (N_13530,N_13203,N_13322);
nand U13531 (N_13531,N_13274,N_13483);
or U13532 (N_13532,N_13405,N_13366);
or U13533 (N_13533,N_13254,N_13484);
nand U13534 (N_13534,N_13352,N_13304);
nor U13535 (N_13535,N_13496,N_13295);
nor U13536 (N_13536,N_13250,N_13401);
and U13537 (N_13537,N_13231,N_13358);
and U13538 (N_13538,N_13238,N_13276);
nand U13539 (N_13539,N_13457,N_13267);
nor U13540 (N_13540,N_13362,N_13220);
nand U13541 (N_13541,N_13392,N_13334);
nor U13542 (N_13542,N_13287,N_13298);
xnor U13543 (N_13543,N_13278,N_13434);
and U13544 (N_13544,N_13465,N_13205);
nand U13545 (N_13545,N_13446,N_13299);
or U13546 (N_13546,N_13209,N_13236);
nand U13547 (N_13547,N_13391,N_13415);
or U13548 (N_13548,N_13335,N_13337);
or U13549 (N_13549,N_13460,N_13445);
nor U13550 (N_13550,N_13413,N_13470);
nor U13551 (N_13551,N_13453,N_13488);
and U13552 (N_13552,N_13290,N_13400);
or U13553 (N_13553,N_13357,N_13439);
nand U13554 (N_13554,N_13403,N_13330);
xnor U13555 (N_13555,N_13476,N_13417);
nand U13556 (N_13556,N_13492,N_13349);
nor U13557 (N_13557,N_13218,N_13423);
nor U13558 (N_13558,N_13285,N_13376);
and U13559 (N_13559,N_13275,N_13448);
nor U13560 (N_13560,N_13431,N_13390);
or U13561 (N_13561,N_13240,N_13316);
xnor U13562 (N_13562,N_13211,N_13306);
and U13563 (N_13563,N_13416,N_13477);
and U13564 (N_13564,N_13206,N_13244);
nor U13565 (N_13565,N_13293,N_13478);
or U13566 (N_13566,N_13271,N_13429);
or U13567 (N_13567,N_13200,N_13264);
or U13568 (N_13568,N_13212,N_13410);
xor U13569 (N_13569,N_13292,N_13251);
nand U13570 (N_13570,N_13255,N_13493);
and U13571 (N_13571,N_13296,N_13452);
or U13572 (N_13572,N_13253,N_13263);
xor U13573 (N_13573,N_13380,N_13397);
and U13574 (N_13574,N_13311,N_13319);
xor U13575 (N_13575,N_13318,N_13329);
or U13576 (N_13576,N_13388,N_13498);
xor U13577 (N_13577,N_13459,N_13424);
and U13578 (N_13578,N_13259,N_13421);
nor U13579 (N_13579,N_13208,N_13449);
nor U13580 (N_13580,N_13382,N_13447);
and U13581 (N_13581,N_13340,N_13471);
xnor U13582 (N_13582,N_13280,N_13458);
nand U13583 (N_13583,N_13393,N_13351);
nor U13584 (N_13584,N_13350,N_13420);
xnor U13585 (N_13585,N_13432,N_13378);
nand U13586 (N_13586,N_13409,N_13346);
xor U13587 (N_13587,N_13385,N_13228);
and U13588 (N_13588,N_13438,N_13289);
xor U13589 (N_13589,N_13338,N_13411);
xor U13590 (N_13590,N_13336,N_13402);
or U13591 (N_13591,N_13226,N_13494);
nor U13592 (N_13592,N_13398,N_13339);
and U13593 (N_13593,N_13474,N_13361);
nand U13594 (N_13594,N_13422,N_13368);
nand U13595 (N_13595,N_13215,N_13480);
nand U13596 (N_13596,N_13224,N_13241);
nor U13597 (N_13597,N_13463,N_13389);
xor U13598 (N_13598,N_13307,N_13252);
or U13599 (N_13599,N_13419,N_13247);
xnor U13600 (N_13600,N_13235,N_13377);
nand U13601 (N_13601,N_13222,N_13210);
nor U13602 (N_13602,N_13291,N_13427);
or U13603 (N_13603,N_13369,N_13473);
and U13604 (N_13604,N_13332,N_13265);
and U13605 (N_13605,N_13426,N_13270);
xnor U13606 (N_13606,N_13261,N_13256);
and U13607 (N_13607,N_13406,N_13418);
nor U13608 (N_13608,N_13333,N_13441);
or U13609 (N_13609,N_13394,N_13284);
nand U13610 (N_13610,N_13269,N_13204);
nand U13611 (N_13611,N_13433,N_13344);
xnor U13612 (N_13612,N_13313,N_13489);
nor U13613 (N_13613,N_13279,N_13408);
xnor U13614 (N_13614,N_13345,N_13227);
nand U13615 (N_13615,N_13342,N_13239);
nor U13616 (N_13616,N_13371,N_13456);
xor U13617 (N_13617,N_13246,N_13232);
and U13618 (N_13618,N_13245,N_13443);
xnor U13619 (N_13619,N_13207,N_13475);
or U13620 (N_13620,N_13315,N_13268);
xor U13621 (N_13621,N_13233,N_13428);
or U13622 (N_13622,N_13472,N_13482);
nor U13623 (N_13623,N_13363,N_13217);
or U13624 (N_13624,N_13242,N_13234);
nand U13625 (N_13625,N_13451,N_13308);
nand U13626 (N_13626,N_13310,N_13272);
and U13627 (N_13627,N_13486,N_13288);
nor U13628 (N_13628,N_13450,N_13495);
and U13629 (N_13629,N_13317,N_13300);
and U13630 (N_13630,N_13348,N_13379);
xnor U13631 (N_13631,N_13323,N_13354);
and U13632 (N_13632,N_13320,N_13386);
and U13633 (N_13633,N_13243,N_13225);
and U13634 (N_13634,N_13499,N_13353);
nand U13635 (N_13635,N_13454,N_13384);
nor U13636 (N_13636,N_13294,N_13201);
and U13637 (N_13637,N_13355,N_13309);
nand U13638 (N_13638,N_13277,N_13485);
and U13639 (N_13639,N_13326,N_13331);
nand U13640 (N_13640,N_13221,N_13414);
xnor U13641 (N_13641,N_13301,N_13229);
nor U13642 (N_13642,N_13305,N_13440);
and U13643 (N_13643,N_13202,N_13302);
nand U13644 (N_13644,N_13223,N_13297);
or U13645 (N_13645,N_13442,N_13435);
xnor U13646 (N_13646,N_13327,N_13273);
and U13647 (N_13647,N_13324,N_13395);
xor U13648 (N_13648,N_13283,N_13396);
and U13649 (N_13649,N_13214,N_13455);
nand U13650 (N_13650,N_13330,N_13271);
nand U13651 (N_13651,N_13492,N_13456);
nor U13652 (N_13652,N_13343,N_13424);
nor U13653 (N_13653,N_13494,N_13216);
nor U13654 (N_13654,N_13440,N_13247);
nand U13655 (N_13655,N_13397,N_13499);
xnor U13656 (N_13656,N_13281,N_13303);
nor U13657 (N_13657,N_13408,N_13313);
and U13658 (N_13658,N_13353,N_13360);
and U13659 (N_13659,N_13224,N_13286);
nand U13660 (N_13660,N_13238,N_13318);
xor U13661 (N_13661,N_13417,N_13434);
xor U13662 (N_13662,N_13333,N_13443);
nor U13663 (N_13663,N_13386,N_13436);
nor U13664 (N_13664,N_13420,N_13243);
and U13665 (N_13665,N_13360,N_13323);
or U13666 (N_13666,N_13408,N_13333);
nor U13667 (N_13667,N_13268,N_13307);
nor U13668 (N_13668,N_13318,N_13493);
xor U13669 (N_13669,N_13276,N_13243);
and U13670 (N_13670,N_13251,N_13372);
and U13671 (N_13671,N_13323,N_13453);
xnor U13672 (N_13672,N_13278,N_13424);
or U13673 (N_13673,N_13337,N_13373);
nand U13674 (N_13674,N_13365,N_13280);
and U13675 (N_13675,N_13463,N_13337);
nand U13676 (N_13676,N_13200,N_13330);
or U13677 (N_13677,N_13213,N_13409);
or U13678 (N_13678,N_13471,N_13256);
xnor U13679 (N_13679,N_13218,N_13417);
and U13680 (N_13680,N_13416,N_13443);
xnor U13681 (N_13681,N_13462,N_13387);
nand U13682 (N_13682,N_13204,N_13412);
or U13683 (N_13683,N_13245,N_13241);
or U13684 (N_13684,N_13436,N_13489);
xor U13685 (N_13685,N_13349,N_13386);
or U13686 (N_13686,N_13229,N_13388);
and U13687 (N_13687,N_13200,N_13238);
and U13688 (N_13688,N_13389,N_13455);
xnor U13689 (N_13689,N_13407,N_13491);
nand U13690 (N_13690,N_13322,N_13275);
nand U13691 (N_13691,N_13368,N_13218);
and U13692 (N_13692,N_13436,N_13423);
xor U13693 (N_13693,N_13435,N_13357);
nand U13694 (N_13694,N_13391,N_13478);
nor U13695 (N_13695,N_13450,N_13397);
or U13696 (N_13696,N_13258,N_13222);
nand U13697 (N_13697,N_13220,N_13371);
and U13698 (N_13698,N_13420,N_13300);
nand U13699 (N_13699,N_13450,N_13373);
nor U13700 (N_13700,N_13309,N_13246);
nor U13701 (N_13701,N_13221,N_13446);
or U13702 (N_13702,N_13364,N_13215);
and U13703 (N_13703,N_13440,N_13430);
xnor U13704 (N_13704,N_13339,N_13340);
nand U13705 (N_13705,N_13425,N_13378);
or U13706 (N_13706,N_13238,N_13270);
nor U13707 (N_13707,N_13231,N_13416);
nand U13708 (N_13708,N_13227,N_13215);
xor U13709 (N_13709,N_13290,N_13480);
nor U13710 (N_13710,N_13427,N_13208);
nand U13711 (N_13711,N_13230,N_13324);
nand U13712 (N_13712,N_13490,N_13437);
nor U13713 (N_13713,N_13465,N_13393);
xor U13714 (N_13714,N_13282,N_13354);
nand U13715 (N_13715,N_13237,N_13490);
xnor U13716 (N_13716,N_13403,N_13459);
nand U13717 (N_13717,N_13237,N_13387);
and U13718 (N_13718,N_13331,N_13493);
xnor U13719 (N_13719,N_13444,N_13371);
xnor U13720 (N_13720,N_13488,N_13342);
and U13721 (N_13721,N_13437,N_13445);
and U13722 (N_13722,N_13463,N_13298);
nor U13723 (N_13723,N_13448,N_13238);
nand U13724 (N_13724,N_13406,N_13246);
or U13725 (N_13725,N_13224,N_13444);
and U13726 (N_13726,N_13313,N_13442);
nor U13727 (N_13727,N_13493,N_13428);
nor U13728 (N_13728,N_13263,N_13456);
nor U13729 (N_13729,N_13434,N_13357);
or U13730 (N_13730,N_13476,N_13449);
and U13731 (N_13731,N_13209,N_13353);
nor U13732 (N_13732,N_13280,N_13463);
and U13733 (N_13733,N_13344,N_13251);
xnor U13734 (N_13734,N_13299,N_13458);
and U13735 (N_13735,N_13225,N_13251);
or U13736 (N_13736,N_13490,N_13213);
or U13737 (N_13737,N_13449,N_13420);
nor U13738 (N_13738,N_13283,N_13334);
xor U13739 (N_13739,N_13413,N_13332);
xor U13740 (N_13740,N_13347,N_13274);
nor U13741 (N_13741,N_13325,N_13376);
and U13742 (N_13742,N_13488,N_13451);
nand U13743 (N_13743,N_13418,N_13273);
or U13744 (N_13744,N_13387,N_13322);
nor U13745 (N_13745,N_13376,N_13372);
and U13746 (N_13746,N_13441,N_13498);
xor U13747 (N_13747,N_13404,N_13206);
xor U13748 (N_13748,N_13286,N_13222);
and U13749 (N_13749,N_13222,N_13372);
xnor U13750 (N_13750,N_13355,N_13496);
or U13751 (N_13751,N_13210,N_13325);
nand U13752 (N_13752,N_13324,N_13449);
and U13753 (N_13753,N_13338,N_13256);
nor U13754 (N_13754,N_13284,N_13397);
nand U13755 (N_13755,N_13238,N_13409);
nor U13756 (N_13756,N_13438,N_13320);
and U13757 (N_13757,N_13326,N_13382);
and U13758 (N_13758,N_13432,N_13260);
xor U13759 (N_13759,N_13293,N_13232);
nor U13760 (N_13760,N_13246,N_13311);
nor U13761 (N_13761,N_13498,N_13233);
or U13762 (N_13762,N_13317,N_13439);
xnor U13763 (N_13763,N_13389,N_13381);
and U13764 (N_13764,N_13293,N_13408);
and U13765 (N_13765,N_13368,N_13426);
nand U13766 (N_13766,N_13452,N_13453);
and U13767 (N_13767,N_13402,N_13284);
nor U13768 (N_13768,N_13490,N_13468);
xnor U13769 (N_13769,N_13484,N_13226);
and U13770 (N_13770,N_13269,N_13220);
or U13771 (N_13771,N_13313,N_13346);
or U13772 (N_13772,N_13379,N_13318);
nor U13773 (N_13773,N_13214,N_13341);
or U13774 (N_13774,N_13203,N_13384);
nand U13775 (N_13775,N_13234,N_13452);
and U13776 (N_13776,N_13417,N_13346);
and U13777 (N_13777,N_13233,N_13397);
nor U13778 (N_13778,N_13384,N_13429);
or U13779 (N_13779,N_13440,N_13465);
and U13780 (N_13780,N_13321,N_13392);
xor U13781 (N_13781,N_13219,N_13252);
or U13782 (N_13782,N_13496,N_13473);
and U13783 (N_13783,N_13295,N_13327);
nor U13784 (N_13784,N_13485,N_13439);
or U13785 (N_13785,N_13241,N_13418);
and U13786 (N_13786,N_13380,N_13366);
nand U13787 (N_13787,N_13409,N_13381);
nor U13788 (N_13788,N_13358,N_13494);
xnor U13789 (N_13789,N_13488,N_13261);
nor U13790 (N_13790,N_13314,N_13403);
or U13791 (N_13791,N_13413,N_13221);
nand U13792 (N_13792,N_13369,N_13277);
xnor U13793 (N_13793,N_13485,N_13233);
and U13794 (N_13794,N_13370,N_13360);
and U13795 (N_13795,N_13304,N_13378);
nand U13796 (N_13796,N_13433,N_13342);
nand U13797 (N_13797,N_13286,N_13362);
nand U13798 (N_13798,N_13226,N_13202);
nor U13799 (N_13799,N_13210,N_13360);
or U13800 (N_13800,N_13710,N_13509);
xnor U13801 (N_13801,N_13538,N_13570);
or U13802 (N_13802,N_13604,N_13504);
xnor U13803 (N_13803,N_13699,N_13720);
xor U13804 (N_13804,N_13781,N_13630);
xor U13805 (N_13805,N_13760,N_13778);
or U13806 (N_13806,N_13680,N_13740);
nand U13807 (N_13807,N_13662,N_13571);
and U13808 (N_13808,N_13721,N_13732);
nor U13809 (N_13809,N_13637,N_13785);
and U13810 (N_13810,N_13739,N_13549);
xnor U13811 (N_13811,N_13718,N_13764);
nor U13812 (N_13812,N_13582,N_13546);
and U13813 (N_13813,N_13735,N_13500);
nor U13814 (N_13814,N_13779,N_13529);
nor U13815 (N_13815,N_13793,N_13695);
nor U13816 (N_13816,N_13745,N_13759);
xnor U13817 (N_13817,N_13667,N_13705);
nand U13818 (N_13818,N_13591,N_13693);
nor U13819 (N_13819,N_13614,N_13645);
xnor U13820 (N_13820,N_13598,N_13643);
nor U13821 (N_13821,N_13661,N_13775);
nand U13822 (N_13822,N_13550,N_13737);
xor U13823 (N_13823,N_13545,N_13722);
xor U13824 (N_13824,N_13756,N_13505);
nand U13825 (N_13825,N_13729,N_13703);
nand U13826 (N_13826,N_13715,N_13569);
and U13827 (N_13827,N_13748,N_13543);
nor U13828 (N_13828,N_13586,N_13743);
nor U13829 (N_13829,N_13572,N_13724);
xnor U13830 (N_13830,N_13664,N_13553);
nor U13831 (N_13831,N_13607,N_13601);
xor U13832 (N_13832,N_13554,N_13762);
xnor U13833 (N_13833,N_13669,N_13501);
or U13834 (N_13834,N_13653,N_13565);
and U13835 (N_13835,N_13518,N_13594);
or U13836 (N_13836,N_13711,N_13640);
or U13837 (N_13837,N_13683,N_13573);
nand U13838 (N_13838,N_13770,N_13516);
nor U13839 (N_13839,N_13686,N_13736);
xor U13840 (N_13840,N_13668,N_13583);
nand U13841 (N_13841,N_13780,N_13615);
and U13842 (N_13842,N_13691,N_13741);
or U13843 (N_13843,N_13787,N_13557);
nor U13844 (N_13844,N_13663,N_13773);
xnor U13845 (N_13845,N_13655,N_13709);
xor U13846 (N_13846,N_13541,N_13520);
nand U13847 (N_13847,N_13690,N_13707);
nor U13848 (N_13848,N_13580,N_13584);
nand U13849 (N_13849,N_13629,N_13552);
xor U13850 (N_13850,N_13613,N_13752);
and U13851 (N_13851,N_13647,N_13673);
xor U13852 (N_13852,N_13763,N_13542);
and U13853 (N_13853,N_13652,N_13589);
xnor U13854 (N_13854,N_13659,N_13547);
nor U13855 (N_13855,N_13731,N_13527);
xnor U13856 (N_13856,N_13517,N_13755);
nor U13857 (N_13857,N_13566,N_13757);
nor U13858 (N_13858,N_13784,N_13749);
nand U13859 (N_13859,N_13798,N_13679);
and U13860 (N_13860,N_13726,N_13638);
or U13861 (N_13861,N_13765,N_13531);
and U13862 (N_13862,N_13644,N_13609);
nor U13863 (N_13863,N_13634,N_13666);
and U13864 (N_13864,N_13617,N_13587);
xnor U13865 (N_13865,N_13767,N_13612);
xnor U13866 (N_13866,N_13562,N_13648);
nand U13867 (N_13867,N_13533,N_13623);
nor U13868 (N_13868,N_13551,N_13649);
nand U13869 (N_13869,N_13610,N_13631);
nor U13870 (N_13870,N_13717,N_13523);
xor U13871 (N_13871,N_13766,N_13596);
xnor U13872 (N_13872,N_13588,N_13506);
nor U13873 (N_13873,N_13620,N_13665);
nor U13874 (N_13874,N_13747,N_13513);
nor U13875 (N_13875,N_13642,N_13611);
nand U13876 (N_13876,N_13579,N_13753);
or U13877 (N_13877,N_13646,N_13657);
and U13878 (N_13878,N_13561,N_13744);
and U13879 (N_13879,N_13592,N_13660);
or U13880 (N_13880,N_13700,N_13532);
nor U13881 (N_13881,N_13602,N_13540);
xnor U13882 (N_13882,N_13618,N_13639);
nor U13883 (N_13883,N_13577,N_13563);
nor U13884 (N_13884,N_13719,N_13564);
xnor U13885 (N_13885,N_13761,N_13599);
nand U13886 (N_13886,N_13578,N_13742);
and U13887 (N_13887,N_13537,N_13692);
nor U13888 (N_13888,N_13674,N_13783);
nor U13889 (N_13889,N_13799,N_13702);
xnor U13890 (N_13890,N_13585,N_13654);
or U13891 (N_13891,N_13603,N_13530);
xnor U13892 (N_13892,N_13725,N_13600);
and U13893 (N_13893,N_13704,N_13696);
xor U13894 (N_13894,N_13574,N_13526);
or U13895 (N_13895,N_13560,N_13777);
nand U13896 (N_13896,N_13670,N_13535);
and U13897 (N_13897,N_13728,N_13524);
nor U13898 (N_13898,N_13624,N_13685);
and U13899 (N_13899,N_13675,N_13567);
xnor U13900 (N_13900,N_13519,N_13672);
nand U13901 (N_13901,N_13619,N_13684);
nand U13902 (N_13902,N_13708,N_13575);
and U13903 (N_13903,N_13627,N_13790);
or U13904 (N_13904,N_13727,N_13713);
or U13905 (N_13905,N_13650,N_13701);
nor U13906 (N_13906,N_13622,N_13733);
nand U13907 (N_13907,N_13568,N_13606);
xor U13908 (N_13908,N_13681,N_13789);
xor U13909 (N_13909,N_13712,N_13698);
nand U13910 (N_13910,N_13633,N_13608);
nor U13911 (N_13911,N_13694,N_13593);
and U13912 (N_13912,N_13628,N_13514);
xnor U13913 (N_13913,N_13671,N_13641);
nand U13914 (N_13914,N_13734,N_13677);
xnor U13915 (N_13915,N_13636,N_13794);
or U13916 (N_13916,N_13597,N_13786);
nand U13917 (N_13917,N_13510,N_13750);
nand U13918 (N_13918,N_13706,N_13626);
nand U13919 (N_13919,N_13697,N_13658);
xnor U13920 (N_13920,N_13512,N_13621);
and U13921 (N_13921,N_13723,N_13656);
or U13922 (N_13922,N_13792,N_13576);
nor U13923 (N_13923,N_13515,N_13714);
and U13924 (N_13924,N_13605,N_13536);
nand U13925 (N_13925,N_13595,N_13544);
or U13926 (N_13926,N_13556,N_13508);
nand U13927 (N_13927,N_13751,N_13503);
nand U13928 (N_13928,N_13581,N_13511);
or U13929 (N_13929,N_13635,N_13791);
or U13930 (N_13930,N_13689,N_13769);
and U13931 (N_13931,N_13539,N_13738);
nand U13932 (N_13932,N_13625,N_13555);
and U13933 (N_13933,N_13796,N_13687);
or U13934 (N_13934,N_13797,N_13774);
and U13935 (N_13935,N_13772,N_13754);
xnor U13936 (N_13936,N_13507,N_13782);
or U13937 (N_13937,N_13558,N_13758);
nor U13938 (N_13938,N_13632,N_13525);
and U13939 (N_13939,N_13730,N_13590);
and U13940 (N_13940,N_13651,N_13688);
xor U13941 (N_13941,N_13616,N_13771);
or U13942 (N_13942,N_13528,N_13502);
nor U13943 (N_13943,N_13768,N_13716);
xor U13944 (N_13944,N_13682,N_13678);
nand U13945 (N_13945,N_13521,N_13559);
and U13946 (N_13946,N_13795,N_13548);
nand U13947 (N_13947,N_13676,N_13522);
or U13948 (N_13948,N_13776,N_13746);
xnor U13949 (N_13949,N_13534,N_13788);
nand U13950 (N_13950,N_13595,N_13662);
nor U13951 (N_13951,N_13553,N_13653);
nor U13952 (N_13952,N_13532,N_13581);
xnor U13953 (N_13953,N_13763,N_13658);
nor U13954 (N_13954,N_13617,N_13561);
xor U13955 (N_13955,N_13549,N_13652);
nand U13956 (N_13956,N_13672,N_13733);
nand U13957 (N_13957,N_13649,N_13735);
and U13958 (N_13958,N_13569,N_13743);
xnor U13959 (N_13959,N_13569,N_13633);
or U13960 (N_13960,N_13532,N_13683);
and U13961 (N_13961,N_13552,N_13722);
xor U13962 (N_13962,N_13588,N_13529);
xnor U13963 (N_13963,N_13538,N_13502);
or U13964 (N_13964,N_13782,N_13562);
xor U13965 (N_13965,N_13506,N_13778);
and U13966 (N_13966,N_13604,N_13721);
or U13967 (N_13967,N_13740,N_13705);
and U13968 (N_13968,N_13665,N_13748);
nor U13969 (N_13969,N_13724,N_13609);
xor U13970 (N_13970,N_13542,N_13696);
and U13971 (N_13971,N_13579,N_13543);
and U13972 (N_13972,N_13792,N_13525);
nand U13973 (N_13973,N_13755,N_13609);
nor U13974 (N_13974,N_13582,N_13763);
xor U13975 (N_13975,N_13694,N_13769);
nor U13976 (N_13976,N_13682,N_13654);
and U13977 (N_13977,N_13621,N_13543);
or U13978 (N_13978,N_13545,N_13748);
or U13979 (N_13979,N_13793,N_13626);
xor U13980 (N_13980,N_13792,N_13647);
and U13981 (N_13981,N_13541,N_13756);
xor U13982 (N_13982,N_13694,N_13588);
and U13983 (N_13983,N_13661,N_13630);
and U13984 (N_13984,N_13515,N_13739);
nor U13985 (N_13985,N_13796,N_13747);
nor U13986 (N_13986,N_13667,N_13563);
and U13987 (N_13987,N_13554,N_13776);
nand U13988 (N_13988,N_13669,N_13722);
or U13989 (N_13989,N_13686,N_13700);
nand U13990 (N_13990,N_13788,N_13555);
or U13991 (N_13991,N_13594,N_13577);
or U13992 (N_13992,N_13780,N_13682);
nand U13993 (N_13993,N_13532,N_13747);
and U13994 (N_13994,N_13604,N_13740);
nor U13995 (N_13995,N_13624,N_13711);
and U13996 (N_13996,N_13702,N_13719);
nand U13997 (N_13997,N_13756,N_13754);
or U13998 (N_13998,N_13781,N_13651);
xor U13999 (N_13999,N_13717,N_13654);
or U14000 (N_14000,N_13694,N_13669);
nand U14001 (N_14001,N_13787,N_13737);
or U14002 (N_14002,N_13543,N_13565);
or U14003 (N_14003,N_13722,N_13623);
or U14004 (N_14004,N_13506,N_13752);
nor U14005 (N_14005,N_13789,N_13593);
and U14006 (N_14006,N_13767,N_13555);
and U14007 (N_14007,N_13786,N_13530);
nand U14008 (N_14008,N_13759,N_13558);
xor U14009 (N_14009,N_13589,N_13762);
nand U14010 (N_14010,N_13795,N_13699);
xor U14011 (N_14011,N_13618,N_13583);
and U14012 (N_14012,N_13601,N_13662);
and U14013 (N_14013,N_13681,N_13553);
nor U14014 (N_14014,N_13682,N_13694);
nand U14015 (N_14015,N_13709,N_13584);
nand U14016 (N_14016,N_13696,N_13720);
or U14017 (N_14017,N_13766,N_13632);
and U14018 (N_14018,N_13554,N_13620);
and U14019 (N_14019,N_13678,N_13652);
or U14020 (N_14020,N_13571,N_13683);
and U14021 (N_14021,N_13571,N_13695);
nand U14022 (N_14022,N_13753,N_13723);
nand U14023 (N_14023,N_13566,N_13777);
nor U14024 (N_14024,N_13692,N_13688);
and U14025 (N_14025,N_13777,N_13708);
nor U14026 (N_14026,N_13518,N_13584);
or U14027 (N_14027,N_13584,N_13724);
or U14028 (N_14028,N_13738,N_13631);
and U14029 (N_14029,N_13576,N_13509);
nand U14030 (N_14030,N_13584,N_13692);
and U14031 (N_14031,N_13795,N_13651);
and U14032 (N_14032,N_13597,N_13538);
or U14033 (N_14033,N_13626,N_13514);
and U14034 (N_14034,N_13794,N_13726);
nor U14035 (N_14035,N_13729,N_13536);
nand U14036 (N_14036,N_13737,N_13742);
nor U14037 (N_14037,N_13720,N_13655);
or U14038 (N_14038,N_13507,N_13624);
or U14039 (N_14039,N_13742,N_13696);
or U14040 (N_14040,N_13529,N_13664);
and U14041 (N_14041,N_13719,N_13683);
and U14042 (N_14042,N_13630,N_13534);
nor U14043 (N_14043,N_13529,N_13600);
xor U14044 (N_14044,N_13727,N_13678);
nor U14045 (N_14045,N_13751,N_13558);
or U14046 (N_14046,N_13545,N_13701);
or U14047 (N_14047,N_13726,N_13655);
nor U14048 (N_14048,N_13695,N_13524);
nand U14049 (N_14049,N_13750,N_13543);
nand U14050 (N_14050,N_13787,N_13728);
nand U14051 (N_14051,N_13733,N_13706);
xnor U14052 (N_14052,N_13515,N_13598);
nand U14053 (N_14053,N_13665,N_13608);
nand U14054 (N_14054,N_13763,N_13717);
or U14055 (N_14055,N_13590,N_13634);
nor U14056 (N_14056,N_13506,N_13696);
nor U14057 (N_14057,N_13529,N_13531);
nor U14058 (N_14058,N_13594,N_13774);
or U14059 (N_14059,N_13748,N_13639);
xor U14060 (N_14060,N_13612,N_13790);
nand U14061 (N_14061,N_13572,N_13697);
and U14062 (N_14062,N_13722,N_13768);
and U14063 (N_14063,N_13510,N_13574);
nand U14064 (N_14064,N_13694,N_13585);
xnor U14065 (N_14065,N_13666,N_13721);
xor U14066 (N_14066,N_13628,N_13703);
and U14067 (N_14067,N_13657,N_13585);
nor U14068 (N_14068,N_13643,N_13613);
xnor U14069 (N_14069,N_13564,N_13519);
and U14070 (N_14070,N_13650,N_13545);
xnor U14071 (N_14071,N_13796,N_13739);
and U14072 (N_14072,N_13648,N_13723);
or U14073 (N_14073,N_13526,N_13630);
nand U14074 (N_14074,N_13509,N_13716);
or U14075 (N_14075,N_13640,N_13550);
or U14076 (N_14076,N_13782,N_13522);
nand U14077 (N_14077,N_13513,N_13653);
xnor U14078 (N_14078,N_13685,N_13757);
or U14079 (N_14079,N_13698,N_13590);
and U14080 (N_14080,N_13695,N_13747);
and U14081 (N_14081,N_13560,N_13749);
nor U14082 (N_14082,N_13619,N_13763);
and U14083 (N_14083,N_13563,N_13598);
xor U14084 (N_14084,N_13546,N_13547);
and U14085 (N_14085,N_13728,N_13781);
and U14086 (N_14086,N_13540,N_13603);
or U14087 (N_14087,N_13562,N_13760);
nor U14088 (N_14088,N_13710,N_13619);
and U14089 (N_14089,N_13709,N_13556);
and U14090 (N_14090,N_13787,N_13629);
and U14091 (N_14091,N_13789,N_13588);
and U14092 (N_14092,N_13791,N_13546);
nand U14093 (N_14093,N_13681,N_13755);
or U14094 (N_14094,N_13735,N_13637);
xor U14095 (N_14095,N_13646,N_13631);
xnor U14096 (N_14096,N_13526,N_13668);
nand U14097 (N_14097,N_13723,N_13775);
and U14098 (N_14098,N_13630,N_13606);
nor U14099 (N_14099,N_13726,N_13700);
or U14100 (N_14100,N_14084,N_13865);
nand U14101 (N_14101,N_13812,N_13876);
nand U14102 (N_14102,N_13951,N_13878);
nand U14103 (N_14103,N_13938,N_13954);
xnor U14104 (N_14104,N_13918,N_13926);
or U14105 (N_14105,N_13939,N_14044);
and U14106 (N_14106,N_13905,N_13891);
xnor U14107 (N_14107,N_13853,N_14083);
nand U14108 (N_14108,N_13934,N_13815);
or U14109 (N_14109,N_14033,N_14047);
or U14110 (N_14110,N_13826,N_13854);
nor U14111 (N_14111,N_13965,N_13829);
nor U14112 (N_14112,N_13869,N_13916);
and U14113 (N_14113,N_13925,N_13836);
or U14114 (N_14114,N_14071,N_14017);
nor U14115 (N_14115,N_13800,N_13949);
xnor U14116 (N_14116,N_14079,N_14015);
nor U14117 (N_14117,N_14048,N_13927);
xnor U14118 (N_14118,N_13945,N_13802);
nor U14119 (N_14119,N_13845,N_13960);
xor U14120 (N_14120,N_14096,N_14072);
or U14121 (N_14121,N_13811,N_14050);
nand U14122 (N_14122,N_14009,N_14073);
nand U14123 (N_14123,N_13838,N_13913);
nor U14124 (N_14124,N_13848,N_14081);
nand U14125 (N_14125,N_14002,N_13807);
and U14126 (N_14126,N_13994,N_13941);
xor U14127 (N_14127,N_14077,N_13944);
nand U14128 (N_14128,N_13874,N_13929);
or U14129 (N_14129,N_14075,N_13942);
xnor U14130 (N_14130,N_13962,N_14091);
and U14131 (N_14131,N_13990,N_14024);
and U14132 (N_14132,N_13983,N_14093);
nand U14133 (N_14133,N_13915,N_14087);
nor U14134 (N_14134,N_14094,N_13861);
nand U14135 (N_14135,N_14032,N_14012);
and U14136 (N_14136,N_13898,N_14008);
nand U14137 (N_14137,N_13816,N_13920);
or U14138 (N_14138,N_14051,N_13988);
and U14139 (N_14139,N_14035,N_14039);
nor U14140 (N_14140,N_13970,N_14003);
and U14141 (N_14141,N_13893,N_13818);
nand U14142 (N_14142,N_13937,N_13914);
xnor U14143 (N_14143,N_14082,N_13888);
xnor U14144 (N_14144,N_13866,N_14059);
or U14145 (N_14145,N_13834,N_13864);
xor U14146 (N_14146,N_13922,N_13863);
nor U14147 (N_14147,N_13832,N_13950);
and U14148 (N_14148,N_13843,N_13917);
and U14149 (N_14149,N_13872,N_13986);
and U14150 (N_14150,N_13856,N_13857);
xor U14151 (N_14151,N_14043,N_14013);
nand U14152 (N_14152,N_14038,N_13956);
nand U14153 (N_14153,N_14052,N_13825);
xnor U14154 (N_14154,N_13882,N_13852);
or U14155 (N_14155,N_13946,N_13849);
or U14156 (N_14156,N_14026,N_13979);
or U14157 (N_14157,N_14067,N_13961);
and U14158 (N_14158,N_14016,N_13881);
nand U14159 (N_14159,N_13907,N_13821);
nor U14160 (N_14160,N_14099,N_13880);
and U14161 (N_14161,N_13996,N_14063);
or U14162 (N_14162,N_14007,N_13931);
or U14163 (N_14163,N_13844,N_13971);
nor U14164 (N_14164,N_13984,N_13987);
nand U14165 (N_14165,N_13885,N_14042);
or U14166 (N_14166,N_14053,N_14064);
and U14167 (N_14167,N_13982,N_13896);
and U14168 (N_14168,N_13894,N_13813);
or U14169 (N_14169,N_13980,N_14005);
nand U14170 (N_14170,N_14022,N_13933);
xor U14171 (N_14171,N_13912,N_14010);
nor U14172 (N_14172,N_13850,N_14001);
or U14173 (N_14173,N_13859,N_13909);
nor U14174 (N_14174,N_13824,N_14074);
and U14175 (N_14175,N_13883,N_13958);
xor U14176 (N_14176,N_13835,N_14061);
nand U14177 (N_14177,N_13801,N_13921);
nand U14178 (N_14178,N_14021,N_13977);
nand U14179 (N_14179,N_13999,N_13957);
or U14180 (N_14180,N_13884,N_14097);
and U14181 (N_14181,N_14068,N_13955);
xor U14182 (N_14182,N_13964,N_13842);
nand U14183 (N_14183,N_13991,N_14019);
and U14184 (N_14184,N_13935,N_13998);
or U14185 (N_14185,N_13901,N_13879);
nor U14186 (N_14186,N_13810,N_13972);
nand U14187 (N_14187,N_13841,N_13870);
nor U14188 (N_14188,N_14089,N_13817);
nand U14189 (N_14189,N_14027,N_13992);
and U14190 (N_14190,N_13887,N_14098);
nand U14191 (N_14191,N_13868,N_13966);
nor U14192 (N_14192,N_13851,N_13846);
nand U14193 (N_14193,N_13959,N_13831);
nor U14194 (N_14194,N_14041,N_13919);
and U14195 (N_14195,N_13936,N_14090);
and U14196 (N_14196,N_13828,N_14037);
nor U14197 (N_14197,N_13837,N_13860);
nand U14198 (N_14198,N_14095,N_13908);
or U14199 (N_14199,N_14028,N_14085);
or U14200 (N_14200,N_13814,N_14049);
or U14201 (N_14201,N_13932,N_14046);
nand U14202 (N_14202,N_13871,N_13975);
nand U14203 (N_14203,N_13974,N_14036);
nor U14204 (N_14204,N_13827,N_13895);
nor U14205 (N_14205,N_13809,N_13886);
and U14206 (N_14206,N_13862,N_14030);
nor U14207 (N_14207,N_13899,N_14076);
xor U14208 (N_14208,N_13858,N_14000);
nand U14209 (N_14209,N_14078,N_13847);
nor U14210 (N_14210,N_13985,N_13875);
and U14211 (N_14211,N_13855,N_13822);
or U14212 (N_14212,N_14018,N_13808);
or U14213 (N_14213,N_14070,N_14060);
nor U14214 (N_14214,N_13804,N_13963);
xor U14215 (N_14215,N_13805,N_13892);
nor U14216 (N_14216,N_13904,N_13897);
xnor U14217 (N_14217,N_14031,N_14055);
and U14218 (N_14218,N_14020,N_14066);
nand U14219 (N_14219,N_13900,N_14092);
nor U14220 (N_14220,N_14069,N_13997);
or U14221 (N_14221,N_13973,N_13943);
nor U14222 (N_14222,N_14034,N_13952);
and U14223 (N_14223,N_14057,N_13978);
nor U14224 (N_14224,N_14065,N_13989);
nand U14225 (N_14225,N_14088,N_14086);
nor U14226 (N_14226,N_14056,N_13911);
xnor U14227 (N_14227,N_13906,N_13993);
and U14228 (N_14228,N_14023,N_14029);
and U14229 (N_14229,N_14054,N_13819);
nor U14230 (N_14230,N_13830,N_14025);
or U14231 (N_14231,N_14004,N_13981);
nand U14232 (N_14232,N_13976,N_14045);
nor U14233 (N_14233,N_13820,N_13833);
or U14234 (N_14234,N_13947,N_13968);
nand U14235 (N_14235,N_13803,N_13930);
and U14236 (N_14236,N_13967,N_14080);
and U14237 (N_14237,N_13902,N_13840);
nand U14238 (N_14238,N_13877,N_13839);
nor U14239 (N_14239,N_14062,N_13940);
nand U14240 (N_14240,N_13873,N_13953);
xor U14241 (N_14241,N_14040,N_14006);
and U14242 (N_14242,N_14014,N_14058);
or U14243 (N_14243,N_13923,N_13889);
xnor U14244 (N_14244,N_13928,N_13903);
nand U14245 (N_14245,N_13890,N_13823);
nor U14246 (N_14246,N_13948,N_13806);
nor U14247 (N_14247,N_14011,N_13969);
or U14248 (N_14248,N_13995,N_13924);
and U14249 (N_14249,N_13867,N_13910);
or U14250 (N_14250,N_13806,N_13868);
and U14251 (N_14251,N_14081,N_14048);
or U14252 (N_14252,N_14086,N_13865);
nor U14253 (N_14253,N_14009,N_14090);
and U14254 (N_14254,N_14029,N_13830);
xor U14255 (N_14255,N_14006,N_13970);
xor U14256 (N_14256,N_14096,N_13988);
nor U14257 (N_14257,N_13903,N_14001);
nor U14258 (N_14258,N_14059,N_14064);
or U14259 (N_14259,N_14069,N_13900);
nor U14260 (N_14260,N_14063,N_13920);
xor U14261 (N_14261,N_13991,N_14042);
or U14262 (N_14262,N_13913,N_14072);
nand U14263 (N_14263,N_14094,N_14002);
nor U14264 (N_14264,N_13802,N_13901);
nand U14265 (N_14265,N_13996,N_13826);
and U14266 (N_14266,N_14067,N_13908);
or U14267 (N_14267,N_13917,N_13841);
nand U14268 (N_14268,N_14093,N_14080);
or U14269 (N_14269,N_13853,N_13916);
nor U14270 (N_14270,N_14027,N_13938);
or U14271 (N_14271,N_13960,N_13957);
nand U14272 (N_14272,N_13836,N_13946);
xnor U14273 (N_14273,N_13938,N_13945);
or U14274 (N_14274,N_13910,N_14033);
xnor U14275 (N_14275,N_13809,N_13894);
or U14276 (N_14276,N_13815,N_14019);
xor U14277 (N_14277,N_13948,N_14033);
nor U14278 (N_14278,N_13972,N_13960);
nor U14279 (N_14279,N_13897,N_13929);
and U14280 (N_14280,N_13960,N_13953);
and U14281 (N_14281,N_13906,N_14030);
nor U14282 (N_14282,N_13979,N_14047);
and U14283 (N_14283,N_13865,N_13845);
nor U14284 (N_14284,N_13861,N_13989);
nor U14285 (N_14285,N_13948,N_14071);
nand U14286 (N_14286,N_14075,N_14061);
and U14287 (N_14287,N_14059,N_13816);
nand U14288 (N_14288,N_14026,N_13978);
and U14289 (N_14289,N_13976,N_13902);
nand U14290 (N_14290,N_13868,N_14029);
xor U14291 (N_14291,N_13839,N_13927);
nor U14292 (N_14292,N_14040,N_13972);
xor U14293 (N_14293,N_13937,N_13813);
and U14294 (N_14294,N_13872,N_13988);
nand U14295 (N_14295,N_13860,N_14028);
nor U14296 (N_14296,N_14020,N_14029);
xor U14297 (N_14297,N_14000,N_13811);
xnor U14298 (N_14298,N_13887,N_14069);
xnor U14299 (N_14299,N_14010,N_13954);
xor U14300 (N_14300,N_14059,N_13900);
or U14301 (N_14301,N_13957,N_13843);
or U14302 (N_14302,N_13843,N_13809);
and U14303 (N_14303,N_13853,N_13964);
nor U14304 (N_14304,N_13984,N_13868);
and U14305 (N_14305,N_13801,N_13907);
or U14306 (N_14306,N_14041,N_14044);
nand U14307 (N_14307,N_13837,N_13955);
nor U14308 (N_14308,N_13991,N_13869);
and U14309 (N_14309,N_13905,N_14049);
nand U14310 (N_14310,N_14071,N_14080);
nand U14311 (N_14311,N_13902,N_14046);
nor U14312 (N_14312,N_13865,N_13837);
nand U14313 (N_14313,N_14069,N_13880);
or U14314 (N_14314,N_14000,N_14033);
nor U14315 (N_14315,N_13885,N_13996);
or U14316 (N_14316,N_13914,N_14012);
or U14317 (N_14317,N_13838,N_13918);
nand U14318 (N_14318,N_14096,N_13960);
nand U14319 (N_14319,N_13862,N_13960);
or U14320 (N_14320,N_13806,N_13929);
or U14321 (N_14321,N_13971,N_14003);
or U14322 (N_14322,N_13845,N_13806);
xor U14323 (N_14323,N_14010,N_13884);
nor U14324 (N_14324,N_13867,N_13911);
xor U14325 (N_14325,N_14035,N_13885);
nand U14326 (N_14326,N_13970,N_13982);
or U14327 (N_14327,N_13800,N_14035);
nand U14328 (N_14328,N_14046,N_14047);
or U14329 (N_14329,N_13842,N_14067);
nor U14330 (N_14330,N_14074,N_14021);
or U14331 (N_14331,N_14034,N_14053);
nor U14332 (N_14332,N_13928,N_14009);
nor U14333 (N_14333,N_13989,N_14071);
nor U14334 (N_14334,N_13853,N_13846);
nand U14335 (N_14335,N_14064,N_14081);
xnor U14336 (N_14336,N_13966,N_13844);
nand U14337 (N_14337,N_14019,N_14027);
xnor U14338 (N_14338,N_13975,N_14095);
nor U14339 (N_14339,N_13911,N_13939);
nor U14340 (N_14340,N_14011,N_13960);
nor U14341 (N_14341,N_13981,N_14008);
or U14342 (N_14342,N_13967,N_13819);
xor U14343 (N_14343,N_14072,N_13972);
or U14344 (N_14344,N_13984,N_13916);
and U14345 (N_14345,N_13940,N_14037);
nand U14346 (N_14346,N_13837,N_13866);
or U14347 (N_14347,N_13815,N_13845);
nand U14348 (N_14348,N_13929,N_13817);
nand U14349 (N_14349,N_13859,N_14096);
or U14350 (N_14350,N_13896,N_13988);
nand U14351 (N_14351,N_13937,N_13845);
xor U14352 (N_14352,N_14075,N_14060);
or U14353 (N_14353,N_14085,N_14087);
and U14354 (N_14354,N_13836,N_13851);
xnor U14355 (N_14355,N_14025,N_13918);
nand U14356 (N_14356,N_14070,N_13932);
and U14357 (N_14357,N_13997,N_13912);
nor U14358 (N_14358,N_13991,N_13963);
nor U14359 (N_14359,N_13824,N_14001);
and U14360 (N_14360,N_14085,N_14012);
xor U14361 (N_14361,N_14066,N_13927);
and U14362 (N_14362,N_13868,N_14091);
nand U14363 (N_14363,N_13907,N_13895);
or U14364 (N_14364,N_14067,N_14086);
and U14365 (N_14365,N_13801,N_13915);
xor U14366 (N_14366,N_13991,N_14064);
nor U14367 (N_14367,N_13851,N_13901);
or U14368 (N_14368,N_13867,N_13856);
nor U14369 (N_14369,N_13933,N_13894);
nor U14370 (N_14370,N_13875,N_14036);
xnor U14371 (N_14371,N_14077,N_14026);
nand U14372 (N_14372,N_14026,N_13867);
nand U14373 (N_14373,N_13833,N_14044);
or U14374 (N_14374,N_13935,N_13982);
nor U14375 (N_14375,N_14036,N_13956);
xor U14376 (N_14376,N_14041,N_13890);
nor U14377 (N_14377,N_13930,N_13988);
and U14378 (N_14378,N_14043,N_13830);
xnor U14379 (N_14379,N_14019,N_13871);
or U14380 (N_14380,N_14035,N_14037);
nor U14381 (N_14381,N_13967,N_13848);
xor U14382 (N_14382,N_13890,N_14038);
or U14383 (N_14383,N_13985,N_13842);
and U14384 (N_14384,N_13850,N_13904);
and U14385 (N_14385,N_13935,N_14094);
xor U14386 (N_14386,N_14020,N_13881);
nor U14387 (N_14387,N_13909,N_13820);
and U14388 (N_14388,N_13803,N_14009);
nand U14389 (N_14389,N_13844,N_14097);
nand U14390 (N_14390,N_14015,N_14045);
nor U14391 (N_14391,N_14042,N_14007);
and U14392 (N_14392,N_13986,N_13870);
and U14393 (N_14393,N_14053,N_13955);
nand U14394 (N_14394,N_13970,N_14087);
and U14395 (N_14395,N_13941,N_13983);
and U14396 (N_14396,N_13940,N_13913);
nand U14397 (N_14397,N_13957,N_14080);
xnor U14398 (N_14398,N_14042,N_13970);
xor U14399 (N_14399,N_14091,N_13974);
or U14400 (N_14400,N_14119,N_14126);
or U14401 (N_14401,N_14230,N_14392);
nor U14402 (N_14402,N_14130,N_14102);
nand U14403 (N_14403,N_14363,N_14173);
or U14404 (N_14404,N_14393,N_14237);
nand U14405 (N_14405,N_14103,N_14251);
nor U14406 (N_14406,N_14279,N_14360);
nor U14407 (N_14407,N_14244,N_14311);
or U14408 (N_14408,N_14328,N_14137);
xnor U14409 (N_14409,N_14180,N_14161);
and U14410 (N_14410,N_14341,N_14302);
or U14411 (N_14411,N_14377,N_14201);
nand U14412 (N_14412,N_14179,N_14389);
nor U14413 (N_14413,N_14358,N_14202);
and U14414 (N_14414,N_14379,N_14219);
xnor U14415 (N_14415,N_14218,N_14252);
nand U14416 (N_14416,N_14142,N_14200);
nor U14417 (N_14417,N_14212,N_14347);
and U14418 (N_14418,N_14308,N_14197);
and U14419 (N_14419,N_14366,N_14185);
nand U14420 (N_14420,N_14123,N_14293);
and U14421 (N_14421,N_14198,N_14143);
nor U14422 (N_14422,N_14221,N_14214);
nand U14423 (N_14423,N_14213,N_14345);
xnor U14424 (N_14424,N_14163,N_14110);
or U14425 (N_14425,N_14340,N_14235);
or U14426 (N_14426,N_14171,N_14304);
or U14427 (N_14427,N_14263,N_14106);
nand U14428 (N_14428,N_14270,N_14354);
xor U14429 (N_14429,N_14210,N_14275);
nor U14430 (N_14430,N_14280,N_14339);
nor U14431 (N_14431,N_14116,N_14211);
or U14432 (N_14432,N_14240,N_14146);
nand U14433 (N_14433,N_14124,N_14284);
and U14434 (N_14434,N_14167,N_14134);
nor U14435 (N_14435,N_14316,N_14307);
nor U14436 (N_14436,N_14314,N_14289);
nand U14437 (N_14437,N_14325,N_14374);
and U14438 (N_14438,N_14370,N_14188);
and U14439 (N_14439,N_14256,N_14331);
or U14440 (N_14440,N_14350,N_14365);
xor U14441 (N_14441,N_14343,N_14248);
xnor U14442 (N_14442,N_14391,N_14385);
xnor U14443 (N_14443,N_14208,N_14382);
and U14444 (N_14444,N_14395,N_14177);
nand U14445 (N_14445,N_14136,N_14108);
nor U14446 (N_14446,N_14181,N_14111);
or U14447 (N_14447,N_14264,N_14132);
and U14448 (N_14448,N_14128,N_14267);
and U14449 (N_14449,N_14149,N_14351);
nor U14450 (N_14450,N_14274,N_14150);
nor U14451 (N_14451,N_14151,N_14156);
nand U14452 (N_14452,N_14259,N_14310);
nor U14453 (N_14453,N_14176,N_14381);
or U14454 (N_14454,N_14352,N_14165);
and U14455 (N_14455,N_14329,N_14399);
nor U14456 (N_14456,N_14193,N_14216);
and U14457 (N_14457,N_14288,N_14120);
or U14458 (N_14458,N_14135,N_14258);
and U14459 (N_14459,N_14182,N_14320);
xnor U14460 (N_14460,N_14349,N_14376);
and U14461 (N_14461,N_14355,N_14159);
xor U14462 (N_14462,N_14315,N_14305);
and U14463 (N_14463,N_14361,N_14330);
xor U14464 (N_14464,N_14217,N_14204);
nor U14465 (N_14465,N_14138,N_14291);
nand U14466 (N_14466,N_14246,N_14286);
or U14467 (N_14467,N_14317,N_14322);
and U14468 (N_14468,N_14139,N_14394);
nand U14469 (N_14469,N_14282,N_14100);
or U14470 (N_14470,N_14371,N_14226);
or U14471 (N_14471,N_14309,N_14236);
nor U14472 (N_14472,N_14312,N_14190);
xnor U14473 (N_14473,N_14373,N_14342);
or U14474 (N_14474,N_14206,N_14195);
nor U14475 (N_14475,N_14144,N_14323);
nand U14476 (N_14476,N_14262,N_14294);
nor U14477 (N_14477,N_14148,N_14306);
and U14478 (N_14478,N_14301,N_14249);
nand U14479 (N_14479,N_14234,N_14155);
and U14480 (N_14480,N_14166,N_14112);
or U14481 (N_14481,N_14285,N_14114);
nor U14482 (N_14482,N_14245,N_14129);
or U14483 (N_14483,N_14327,N_14368);
nand U14484 (N_14484,N_14162,N_14318);
nand U14485 (N_14485,N_14276,N_14222);
xnor U14486 (N_14486,N_14261,N_14141);
nor U14487 (N_14487,N_14319,N_14337);
xor U14488 (N_14488,N_14260,N_14292);
nor U14489 (N_14489,N_14272,N_14125);
nor U14490 (N_14490,N_14115,N_14196);
and U14491 (N_14491,N_14191,N_14187);
and U14492 (N_14492,N_14220,N_14287);
and U14493 (N_14493,N_14170,N_14160);
xnor U14494 (N_14494,N_14344,N_14283);
xnor U14495 (N_14495,N_14117,N_14239);
nor U14496 (N_14496,N_14192,N_14133);
xor U14497 (N_14497,N_14326,N_14247);
and U14498 (N_14498,N_14168,N_14298);
or U14499 (N_14499,N_14215,N_14300);
and U14500 (N_14500,N_14357,N_14253);
and U14501 (N_14501,N_14223,N_14225);
nor U14502 (N_14502,N_14209,N_14254);
or U14503 (N_14503,N_14348,N_14296);
nand U14504 (N_14504,N_14388,N_14233);
nand U14505 (N_14505,N_14383,N_14333);
xor U14506 (N_14506,N_14127,N_14378);
or U14507 (N_14507,N_14397,N_14290);
and U14508 (N_14508,N_14153,N_14295);
xnor U14509 (N_14509,N_14122,N_14207);
and U14510 (N_14510,N_14158,N_14268);
or U14511 (N_14511,N_14242,N_14396);
and U14512 (N_14512,N_14109,N_14375);
or U14513 (N_14513,N_14121,N_14189);
nor U14514 (N_14514,N_14224,N_14324);
xnor U14515 (N_14515,N_14147,N_14297);
and U14516 (N_14516,N_14265,N_14243);
xnor U14517 (N_14517,N_14369,N_14232);
xnor U14518 (N_14518,N_14199,N_14157);
nor U14519 (N_14519,N_14269,N_14338);
and U14520 (N_14520,N_14299,N_14172);
or U14521 (N_14521,N_14184,N_14107);
or U14522 (N_14522,N_14281,N_14131);
and U14523 (N_14523,N_14390,N_14205);
nor U14524 (N_14524,N_14178,N_14321);
or U14525 (N_14525,N_14227,N_14277);
and U14526 (N_14526,N_14332,N_14346);
and U14527 (N_14527,N_14387,N_14113);
xor U14528 (N_14528,N_14105,N_14255);
nand U14529 (N_14529,N_14257,N_14271);
nand U14530 (N_14530,N_14145,N_14356);
and U14531 (N_14531,N_14336,N_14359);
nand U14532 (N_14532,N_14384,N_14194);
and U14533 (N_14533,N_14398,N_14203);
or U14534 (N_14534,N_14101,N_14353);
nor U14535 (N_14535,N_14278,N_14380);
xnor U14536 (N_14536,N_14241,N_14362);
xnor U14537 (N_14537,N_14386,N_14372);
nor U14538 (N_14538,N_14169,N_14152);
nand U14539 (N_14539,N_14273,N_14266);
xnor U14540 (N_14540,N_14183,N_14303);
nor U14541 (N_14541,N_14174,N_14238);
xor U14542 (N_14542,N_14118,N_14250);
nand U14543 (N_14543,N_14186,N_14175);
or U14544 (N_14544,N_14335,N_14313);
and U14545 (N_14545,N_14334,N_14104);
and U14546 (N_14546,N_14154,N_14228);
nor U14547 (N_14547,N_14229,N_14164);
and U14548 (N_14548,N_14364,N_14367);
or U14549 (N_14549,N_14231,N_14140);
or U14550 (N_14550,N_14182,N_14352);
nor U14551 (N_14551,N_14248,N_14186);
and U14552 (N_14552,N_14146,N_14248);
or U14553 (N_14553,N_14167,N_14197);
nand U14554 (N_14554,N_14284,N_14188);
nand U14555 (N_14555,N_14366,N_14309);
and U14556 (N_14556,N_14344,N_14186);
or U14557 (N_14557,N_14233,N_14289);
or U14558 (N_14558,N_14230,N_14364);
xor U14559 (N_14559,N_14140,N_14389);
and U14560 (N_14560,N_14217,N_14261);
nor U14561 (N_14561,N_14157,N_14164);
and U14562 (N_14562,N_14279,N_14110);
xnor U14563 (N_14563,N_14281,N_14200);
nand U14564 (N_14564,N_14257,N_14290);
or U14565 (N_14565,N_14188,N_14116);
nor U14566 (N_14566,N_14284,N_14357);
nor U14567 (N_14567,N_14226,N_14389);
or U14568 (N_14568,N_14327,N_14107);
nand U14569 (N_14569,N_14299,N_14129);
and U14570 (N_14570,N_14326,N_14394);
nor U14571 (N_14571,N_14163,N_14214);
or U14572 (N_14572,N_14152,N_14386);
nor U14573 (N_14573,N_14396,N_14339);
and U14574 (N_14574,N_14107,N_14230);
nand U14575 (N_14575,N_14161,N_14384);
and U14576 (N_14576,N_14389,N_14257);
nand U14577 (N_14577,N_14194,N_14217);
xor U14578 (N_14578,N_14378,N_14166);
nand U14579 (N_14579,N_14209,N_14380);
nor U14580 (N_14580,N_14383,N_14163);
and U14581 (N_14581,N_14196,N_14258);
xnor U14582 (N_14582,N_14355,N_14354);
xnor U14583 (N_14583,N_14143,N_14385);
nor U14584 (N_14584,N_14277,N_14329);
nor U14585 (N_14585,N_14280,N_14209);
xor U14586 (N_14586,N_14170,N_14153);
nand U14587 (N_14587,N_14201,N_14138);
nor U14588 (N_14588,N_14171,N_14246);
and U14589 (N_14589,N_14252,N_14363);
or U14590 (N_14590,N_14167,N_14195);
xnor U14591 (N_14591,N_14158,N_14336);
or U14592 (N_14592,N_14317,N_14187);
and U14593 (N_14593,N_14137,N_14359);
or U14594 (N_14594,N_14304,N_14337);
nand U14595 (N_14595,N_14271,N_14280);
or U14596 (N_14596,N_14114,N_14203);
or U14597 (N_14597,N_14123,N_14121);
and U14598 (N_14598,N_14199,N_14368);
nor U14599 (N_14599,N_14374,N_14169);
xnor U14600 (N_14600,N_14145,N_14315);
and U14601 (N_14601,N_14238,N_14260);
and U14602 (N_14602,N_14141,N_14119);
nand U14603 (N_14603,N_14153,N_14346);
nor U14604 (N_14604,N_14386,N_14388);
xnor U14605 (N_14605,N_14162,N_14331);
or U14606 (N_14606,N_14311,N_14135);
nor U14607 (N_14607,N_14168,N_14244);
nand U14608 (N_14608,N_14342,N_14326);
xnor U14609 (N_14609,N_14223,N_14193);
and U14610 (N_14610,N_14103,N_14265);
and U14611 (N_14611,N_14113,N_14105);
xnor U14612 (N_14612,N_14173,N_14380);
nand U14613 (N_14613,N_14344,N_14321);
and U14614 (N_14614,N_14382,N_14249);
nand U14615 (N_14615,N_14228,N_14233);
nor U14616 (N_14616,N_14334,N_14210);
and U14617 (N_14617,N_14220,N_14347);
or U14618 (N_14618,N_14302,N_14330);
nor U14619 (N_14619,N_14113,N_14396);
nand U14620 (N_14620,N_14217,N_14312);
nand U14621 (N_14621,N_14269,N_14296);
nand U14622 (N_14622,N_14111,N_14296);
nor U14623 (N_14623,N_14374,N_14354);
or U14624 (N_14624,N_14330,N_14124);
nor U14625 (N_14625,N_14124,N_14145);
and U14626 (N_14626,N_14223,N_14262);
and U14627 (N_14627,N_14135,N_14215);
xnor U14628 (N_14628,N_14357,N_14217);
and U14629 (N_14629,N_14254,N_14338);
xor U14630 (N_14630,N_14222,N_14186);
xor U14631 (N_14631,N_14222,N_14315);
xor U14632 (N_14632,N_14295,N_14279);
nor U14633 (N_14633,N_14348,N_14234);
nand U14634 (N_14634,N_14116,N_14353);
nand U14635 (N_14635,N_14182,N_14124);
nand U14636 (N_14636,N_14172,N_14170);
nor U14637 (N_14637,N_14239,N_14288);
xnor U14638 (N_14638,N_14380,N_14326);
nor U14639 (N_14639,N_14170,N_14168);
xnor U14640 (N_14640,N_14220,N_14329);
nor U14641 (N_14641,N_14278,N_14357);
nand U14642 (N_14642,N_14278,N_14245);
and U14643 (N_14643,N_14399,N_14210);
and U14644 (N_14644,N_14295,N_14123);
nor U14645 (N_14645,N_14297,N_14237);
or U14646 (N_14646,N_14387,N_14321);
nor U14647 (N_14647,N_14334,N_14276);
xnor U14648 (N_14648,N_14197,N_14399);
and U14649 (N_14649,N_14334,N_14118);
nor U14650 (N_14650,N_14348,N_14122);
and U14651 (N_14651,N_14273,N_14363);
or U14652 (N_14652,N_14265,N_14280);
nor U14653 (N_14653,N_14260,N_14290);
nor U14654 (N_14654,N_14376,N_14365);
and U14655 (N_14655,N_14280,N_14110);
xor U14656 (N_14656,N_14194,N_14112);
nor U14657 (N_14657,N_14260,N_14226);
xnor U14658 (N_14658,N_14331,N_14302);
and U14659 (N_14659,N_14166,N_14158);
nand U14660 (N_14660,N_14102,N_14337);
and U14661 (N_14661,N_14221,N_14171);
nand U14662 (N_14662,N_14194,N_14387);
nand U14663 (N_14663,N_14244,N_14351);
nand U14664 (N_14664,N_14211,N_14347);
nand U14665 (N_14665,N_14340,N_14227);
or U14666 (N_14666,N_14225,N_14239);
xnor U14667 (N_14667,N_14299,N_14261);
xnor U14668 (N_14668,N_14152,N_14285);
xor U14669 (N_14669,N_14277,N_14345);
and U14670 (N_14670,N_14245,N_14166);
nor U14671 (N_14671,N_14239,N_14217);
and U14672 (N_14672,N_14355,N_14306);
nor U14673 (N_14673,N_14344,N_14177);
and U14674 (N_14674,N_14364,N_14237);
and U14675 (N_14675,N_14189,N_14390);
nand U14676 (N_14676,N_14122,N_14109);
and U14677 (N_14677,N_14378,N_14379);
nand U14678 (N_14678,N_14117,N_14340);
nor U14679 (N_14679,N_14279,N_14354);
and U14680 (N_14680,N_14156,N_14208);
xor U14681 (N_14681,N_14388,N_14325);
xnor U14682 (N_14682,N_14263,N_14350);
xnor U14683 (N_14683,N_14329,N_14170);
or U14684 (N_14684,N_14201,N_14224);
or U14685 (N_14685,N_14341,N_14296);
or U14686 (N_14686,N_14274,N_14391);
and U14687 (N_14687,N_14243,N_14289);
nor U14688 (N_14688,N_14282,N_14281);
nor U14689 (N_14689,N_14362,N_14158);
and U14690 (N_14690,N_14299,N_14240);
xnor U14691 (N_14691,N_14102,N_14114);
and U14692 (N_14692,N_14338,N_14355);
nor U14693 (N_14693,N_14238,N_14300);
and U14694 (N_14694,N_14322,N_14167);
nor U14695 (N_14695,N_14177,N_14285);
or U14696 (N_14696,N_14126,N_14312);
xor U14697 (N_14697,N_14322,N_14115);
nor U14698 (N_14698,N_14318,N_14320);
and U14699 (N_14699,N_14343,N_14245);
nor U14700 (N_14700,N_14493,N_14656);
nor U14701 (N_14701,N_14515,N_14440);
nor U14702 (N_14702,N_14499,N_14542);
or U14703 (N_14703,N_14682,N_14590);
or U14704 (N_14704,N_14678,N_14520);
xor U14705 (N_14705,N_14665,N_14626);
and U14706 (N_14706,N_14482,N_14405);
or U14707 (N_14707,N_14488,N_14662);
and U14708 (N_14708,N_14413,N_14483);
nand U14709 (N_14709,N_14593,N_14492);
nor U14710 (N_14710,N_14543,N_14504);
nand U14711 (N_14711,N_14580,N_14638);
nand U14712 (N_14712,N_14489,N_14695);
nand U14713 (N_14713,N_14636,N_14581);
xor U14714 (N_14714,N_14446,N_14574);
nor U14715 (N_14715,N_14655,N_14664);
or U14716 (N_14716,N_14685,N_14417);
nand U14717 (N_14717,N_14582,N_14452);
xor U14718 (N_14718,N_14619,N_14475);
nand U14719 (N_14719,N_14432,N_14651);
nor U14720 (N_14720,N_14552,N_14553);
nand U14721 (N_14721,N_14647,N_14532);
or U14722 (N_14722,N_14420,N_14676);
nand U14723 (N_14723,N_14568,N_14539);
xor U14724 (N_14724,N_14439,N_14622);
nand U14725 (N_14725,N_14434,N_14663);
nor U14726 (N_14726,N_14579,N_14567);
nand U14727 (N_14727,N_14607,N_14572);
and U14728 (N_14728,N_14536,N_14545);
nor U14729 (N_14729,N_14465,N_14627);
or U14730 (N_14730,N_14550,N_14598);
nand U14731 (N_14731,N_14654,N_14642);
nor U14732 (N_14732,N_14497,N_14674);
and U14733 (N_14733,N_14584,N_14407);
nand U14734 (N_14734,N_14672,N_14697);
nand U14735 (N_14735,N_14606,N_14524);
nor U14736 (N_14736,N_14670,N_14435);
nand U14737 (N_14737,N_14408,N_14612);
nor U14738 (N_14738,N_14681,N_14591);
xnor U14739 (N_14739,N_14538,N_14621);
nand U14740 (N_14740,N_14464,N_14560);
nand U14741 (N_14741,N_14510,N_14433);
nor U14742 (N_14742,N_14570,N_14437);
or U14743 (N_14743,N_14523,N_14611);
nand U14744 (N_14744,N_14625,N_14595);
and U14745 (N_14745,N_14461,N_14491);
or U14746 (N_14746,N_14617,N_14644);
nor U14747 (N_14747,N_14605,N_14427);
and U14748 (N_14748,N_14571,N_14506);
xnor U14749 (N_14749,N_14573,N_14691);
nor U14750 (N_14750,N_14529,N_14406);
xnor U14751 (N_14751,N_14615,N_14438);
and U14752 (N_14752,N_14501,N_14460);
nand U14753 (N_14753,N_14618,N_14423);
xnor U14754 (N_14754,N_14409,N_14528);
nor U14755 (N_14755,N_14657,N_14425);
nor U14756 (N_14756,N_14609,N_14457);
and U14757 (N_14757,N_14601,N_14634);
and U14758 (N_14758,N_14480,N_14496);
nand U14759 (N_14759,N_14455,N_14470);
nor U14760 (N_14760,N_14462,N_14479);
or U14761 (N_14761,N_14402,N_14505);
xnor U14762 (N_14762,N_14551,N_14445);
xnor U14763 (N_14763,N_14535,N_14577);
and U14764 (N_14764,N_14679,N_14694);
xnor U14765 (N_14765,N_14426,N_14419);
and U14766 (N_14766,N_14667,N_14646);
nand U14767 (N_14767,N_14661,N_14521);
nor U14768 (N_14768,N_14507,N_14444);
xnor U14769 (N_14769,N_14671,N_14564);
nor U14770 (N_14770,N_14546,N_14549);
xor U14771 (N_14771,N_14513,N_14699);
xnor U14772 (N_14772,N_14487,N_14451);
xor U14773 (N_14773,N_14599,N_14533);
nand U14774 (N_14774,N_14473,N_14589);
nor U14775 (N_14775,N_14540,N_14525);
nor U14776 (N_14776,N_14404,N_14698);
nand U14777 (N_14777,N_14410,N_14453);
nor U14778 (N_14778,N_14516,N_14411);
nor U14779 (N_14779,N_14639,N_14641);
or U14780 (N_14780,N_14680,N_14458);
and U14781 (N_14781,N_14512,N_14422);
or U14782 (N_14782,N_14643,N_14631);
nand U14783 (N_14783,N_14576,N_14696);
nor U14784 (N_14784,N_14517,N_14594);
nand U14785 (N_14785,N_14463,N_14485);
or U14786 (N_14786,N_14401,N_14624);
or U14787 (N_14787,N_14562,N_14459);
xor U14788 (N_14788,N_14467,N_14565);
and U14789 (N_14789,N_14415,N_14561);
nor U14790 (N_14790,N_14469,N_14414);
nor U14791 (N_14791,N_14548,N_14478);
nor U14792 (N_14792,N_14660,N_14400);
and U14793 (N_14793,N_14658,N_14403);
nor U14794 (N_14794,N_14466,N_14428);
and U14795 (N_14795,N_14687,N_14632);
nor U14796 (N_14796,N_14556,N_14602);
and U14797 (N_14797,N_14441,N_14472);
and U14798 (N_14798,N_14494,N_14669);
and U14799 (N_14799,N_14587,N_14531);
nand U14800 (N_14800,N_14650,N_14637);
nor U14801 (N_14801,N_14675,N_14603);
xnor U14802 (N_14802,N_14692,N_14673);
xor U14803 (N_14803,N_14508,N_14511);
xor U14804 (N_14804,N_14514,N_14436);
xor U14805 (N_14805,N_14592,N_14683);
nor U14806 (N_14806,N_14690,N_14623);
nand U14807 (N_14807,N_14559,N_14454);
nor U14808 (N_14808,N_14490,N_14486);
or U14809 (N_14809,N_14530,N_14557);
xnor U14810 (N_14810,N_14421,N_14563);
or U14811 (N_14811,N_14575,N_14484);
or U14812 (N_14812,N_14544,N_14443);
nand U14813 (N_14813,N_14430,N_14537);
or U14814 (N_14814,N_14554,N_14447);
xnor U14815 (N_14815,N_14471,N_14500);
or U14816 (N_14816,N_14630,N_14610);
xor U14817 (N_14817,N_14498,N_14527);
or U14818 (N_14818,N_14468,N_14600);
and U14819 (N_14819,N_14693,N_14547);
or U14820 (N_14820,N_14450,N_14534);
or U14821 (N_14821,N_14648,N_14653);
or U14822 (N_14822,N_14649,N_14519);
and U14823 (N_14823,N_14566,N_14456);
nand U14824 (N_14824,N_14583,N_14596);
nand U14825 (N_14825,N_14613,N_14666);
nor U14826 (N_14826,N_14502,N_14588);
nor U14827 (N_14827,N_14616,N_14555);
nand U14828 (N_14828,N_14604,N_14614);
or U14829 (N_14829,N_14569,N_14448);
nand U14830 (N_14830,N_14476,N_14503);
xnor U14831 (N_14831,N_14659,N_14431);
nor U14832 (N_14832,N_14597,N_14418);
xnor U14833 (N_14833,N_14684,N_14558);
nor U14834 (N_14834,N_14449,N_14629);
xor U14835 (N_14835,N_14586,N_14424);
and U14836 (N_14836,N_14578,N_14645);
and U14837 (N_14837,N_14509,N_14635);
nor U14838 (N_14838,N_14677,N_14686);
nor U14839 (N_14839,N_14474,N_14526);
xnor U14840 (N_14840,N_14688,N_14412);
xnor U14841 (N_14841,N_14416,N_14495);
nand U14842 (N_14842,N_14628,N_14652);
or U14843 (N_14843,N_14689,N_14633);
xor U14844 (N_14844,N_14640,N_14541);
nand U14845 (N_14845,N_14429,N_14585);
and U14846 (N_14846,N_14620,N_14518);
xor U14847 (N_14847,N_14481,N_14442);
nand U14848 (N_14848,N_14608,N_14477);
nor U14849 (N_14849,N_14668,N_14522);
and U14850 (N_14850,N_14466,N_14447);
and U14851 (N_14851,N_14420,N_14604);
and U14852 (N_14852,N_14636,N_14579);
nor U14853 (N_14853,N_14440,N_14529);
nor U14854 (N_14854,N_14484,N_14496);
nand U14855 (N_14855,N_14562,N_14456);
nand U14856 (N_14856,N_14498,N_14592);
nand U14857 (N_14857,N_14443,N_14520);
nor U14858 (N_14858,N_14530,N_14566);
and U14859 (N_14859,N_14651,N_14504);
nor U14860 (N_14860,N_14511,N_14458);
or U14861 (N_14861,N_14596,N_14503);
nand U14862 (N_14862,N_14547,N_14562);
nand U14863 (N_14863,N_14492,N_14673);
nand U14864 (N_14864,N_14478,N_14490);
or U14865 (N_14865,N_14416,N_14574);
nor U14866 (N_14866,N_14594,N_14595);
or U14867 (N_14867,N_14683,N_14628);
nor U14868 (N_14868,N_14404,N_14584);
and U14869 (N_14869,N_14495,N_14431);
or U14870 (N_14870,N_14681,N_14464);
or U14871 (N_14871,N_14422,N_14598);
and U14872 (N_14872,N_14661,N_14530);
nand U14873 (N_14873,N_14420,N_14606);
nor U14874 (N_14874,N_14413,N_14500);
and U14875 (N_14875,N_14557,N_14523);
and U14876 (N_14876,N_14674,N_14699);
nor U14877 (N_14877,N_14506,N_14575);
or U14878 (N_14878,N_14535,N_14536);
or U14879 (N_14879,N_14496,N_14477);
nor U14880 (N_14880,N_14408,N_14690);
and U14881 (N_14881,N_14483,N_14488);
nor U14882 (N_14882,N_14686,N_14599);
and U14883 (N_14883,N_14510,N_14423);
nor U14884 (N_14884,N_14484,N_14528);
xor U14885 (N_14885,N_14548,N_14685);
and U14886 (N_14886,N_14418,N_14401);
nor U14887 (N_14887,N_14528,N_14582);
xnor U14888 (N_14888,N_14443,N_14602);
and U14889 (N_14889,N_14584,N_14499);
or U14890 (N_14890,N_14461,N_14547);
nand U14891 (N_14891,N_14442,N_14474);
or U14892 (N_14892,N_14417,N_14454);
nand U14893 (N_14893,N_14692,N_14604);
or U14894 (N_14894,N_14666,N_14578);
nor U14895 (N_14895,N_14541,N_14469);
nand U14896 (N_14896,N_14622,N_14450);
or U14897 (N_14897,N_14577,N_14589);
nand U14898 (N_14898,N_14608,N_14438);
or U14899 (N_14899,N_14431,N_14494);
nand U14900 (N_14900,N_14433,N_14425);
xnor U14901 (N_14901,N_14469,N_14584);
and U14902 (N_14902,N_14509,N_14513);
and U14903 (N_14903,N_14467,N_14602);
and U14904 (N_14904,N_14566,N_14691);
nor U14905 (N_14905,N_14450,N_14547);
xnor U14906 (N_14906,N_14596,N_14686);
xnor U14907 (N_14907,N_14615,N_14467);
and U14908 (N_14908,N_14432,N_14578);
and U14909 (N_14909,N_14404,N_14690);
xor U14910 (N_14910,N_14620,N_14493);
and U14911 (N_14911,N_14524,N_14472);
xnor U14912 (N_14912,N_14598,N_14520);
or U14913 (N_14913,N_14603,N_14617);
xnor U14914 (N_14914,N_14462,N_14644);
nand U14915 (N_14915,N_14447,N_14450);
nand U14916 (N_14916,N_14523,N_14468);
xnor U14917 (N_14917,N_14552,N_14457);
nand U14918 (N_14918,N_14600,N_14637);
or U14919 (N_14919,N_14616,N_14688);
nand U14920 (N_14920,N_14618,N_14586);
xor U14921 (N_14921,N_14645,N_14640);
xor U14922 (N_14922,N_14612,N_14534);
nand U14923 (N_14923,N_14637,N_14403);
nor U14924 (N_14924,N_14546,N_14417);
nand U14925 (N_14925,N_14427,N_14406);
nand U14926 (N_14926,N_14568,N_14525);
or U14927 (N_14927,N_14661,N_14600);
or U14928 (N_14928,N_14573,N_14518);
xnor U14929 (N_14929,N_14490,N_14577);
or U14930 (N_14930,N_14538,N_14463);
or U14931 (N_14931,N_14607,N_14410);
or U14932 (N_14932,N_14433,N_14646);
xnor U14933 (N_14933,N_14511,N_14673);
or U14934 (N_14934,N_14622,N_14614);
or U14935 (N_14935,N_14619,N_14686);
nor U14936 (N_14936,N_14538,N_14520);
xnor U14937 (N_14937,N_14484,N_14511);
nand U14938 (N_14938,N_14443,N_14627);
nor U14939 (N_14939,N_14459,N_14675);
or U14940 (N_14940,N_14573,N_14675);
xor U14941 (N_14941,N_14548,N_14675);
and U14942 (N_14942,N_14672,N_14510);
and U14943 (N_14943,N_14412,N_14583);
xor U14944 (N_14944,N_14461,N_14448);
nand U14945 (N_14945,N_14630,N_14501);
or U14946 (N_14946,N_14565,N_14630);
xor U14947 (N_14947,N_14531,N_14551);
xor U14948 (N_14948,N_14479,N_14641);
or U14949 (N_14949,N_14678,N_14580);
and U14950 (N_14950,N_14597,N_14679);
or U14951 (N_14951,N_14686,N_14461);
nor U14952 (N_14952,N_14567,N_14513);
or U14953 (N_14953,N_14687,N_14456);
nor U14954 (N_14954,N_14681,N_14615);
xnor U14955 (N_14955,N_14433,N_14610);
or U14956 (N_14956,N_14625,N_14513);
or U14957 (N_14957,N_14433,N_14682);
nor U14958 (N_14958,N_14454,N_14520);
nand U14959 (N_14959,N_14446,N_14556);
nand U14960 (N_14960,N_14455,N_14663);
nor U14961 (N_14961,N_14529,N_14474);
xor U14962 (N_14962,N_14677,N_14641);
or U14963 (N_14963,N_14476,N_14573);
or U14964 (N_14964,N_14645,N_14444);
or U14965 (N_14965,N_14475,N_14465);
nand U14966 (N_14966,N_14543,N_14616);
and U14967 (N_14967,N_14427,N_14580);
and U14968 (N_14968,N_14634,N_14486);
nand U14969 (N_14969,N_14467,N_14646);
nand U14970 (N_14970,N_14467,N_14563);
nand U14971 (N_14971,N_14403,N_14537);
or U14972 (N_14972,N_14482,N_14659);
xnor U14973 (N_14973,N_14593,N_14519);
xnor U14974 (N_14974,N_14635,N_14673);
nor U14975 (N_14975,N_14418,N_14698);
nand U14976 (N_14976,N_14690,N_14403);
nand U14977 (N_14977,N_14630,N_14596);
xor U14978 (N_14978,N_14664,N_14619);
nand U14979 (N_14979,N_14635,N_14614);
or U14980 (N_14980,N_14437,N_14506);
and U14981 (N_14981,N_14655,N_14609);
nor U14982 (N_14982,N_14667,N_14423);
or U14983 (N_14983,N_14546,N_14598);
or U14984 (N_14984,N_14670,N_14498);
nand U14985 (N_14985,N_14612,N_14609);
xor U14986 (N_14986,N_14575,N_14592);
and U14987 (N_14987,N_14628,N_14426);
nand U14988 (N_14988,N_14635,N_14452);
or U14989 (N_14989,N_14698,N_14508);
nor U14990 (N_14990,N_14626,N_14507);
or U14991 (N_14991,N_14693,N_14430);
xnor U14992 (N_14992,N_14408,N_14559);
nor U14993 (N_14993,N_14585,N_14671);
nand U14994 (N_14994,N_14518,N_14679);
nor U14995 (N_14995,N_14538,N_14548);
and U14996 (N_14996,N_14438,N_14431);
and U14997 (N_14997,N_14640,N_14417);
xnor U14998 (N_14998,N_14479,N_14476);
nand U14999 (N_14999,N_14624,N_14531);
xnor U15000 (N_15000,N_14895,N_14930);
nand U15001 (N_15001,N_14734,N_14738);
xor U15002 (N_15002,N_14727,N_14902);
nor U15003 (N_15003,N_14759,N_14985);
and U15004 (N_15004,N_14980,N_14712);
xor U15005 (N_15005,N_14748,N_14894);
or U15006 (N_15006,N_14812,N_14720);
nand U15007 (N_15007,N_14883,N_14929);
xnor U15008 (N_15008,N_14804,N_14999);
nand U15009 (N_15009,N_14992,N_14993);
nor U15010 (N_15010,N_14885,N_14799);
nor U15011 (N_15011,N_14805,N_14852);
nor U15012 (N_15012,N_14763,N_14907);
or U15013 (N_15013,N_14719,N_14713);
and U15014 (N_15014,N_14771,N_14953);
nand U15015 (N_15015,N_14906,N_14728);
xnor U15016 (N_15016,N_14781,N_14753);
nor U15017 (N_15017,N_14939,N_14811);
and U15018 (N_15018,N_14867,N_14908);
xnor U15019 (N_15019,N_14888,N_14705);
nand U15020 (N_15020,N_14944,N_14875);
and U15021 (N_15021,N_14795,N_14722);
nand U15022 (N_15022,N_14864,N_14785);
nand U15023 (N_15023,N_14898,N_14987);
or U15024 (N_15024,N_14945,N_14779);
or U15025 (N_15025,N_14965,N_14765);
nor U15026 (N_15026,N_14813,N_14994);
nand U15027 (N_15027,N_14958,N_14851);
or U15028 (N_15028,N_14830,N_14900);
nand U15029 (N_15029,N_14941,N_14866);
nand U15030 (N_15030,N_14797,N_14701);
and U15031 (N_15031,N_14772,N_14706);
nor U15032 (N_15032,N_14882,N_14726);
nor U15033 (N_15033,N_14767,N_14715);
and U15034 (N_15034,N_14787,N_14912);
or U15035 (N_15035,N_14909,N_14744);
or U15036 (N_15036,N_14931,N_14959);
nor U15037 (N_15037,N_14950,N_14951);
xor U15038 (N_15038,N_14755,N_14732);
and U15039 (N_15039,N_14904,N_14818);
nand U15040 (N_15040,N_14923,N_14741);
or U15041 (N_15041,N_14717,N_14998);
nand U15042 (N_15042,N_14833,N_14820);
xor U15043 (N_15043,N_14822,N_14920);
nand U15044 (N_15044,N_14889,N_14873);
or U15045 (N_15045,N_14915,N_14709);
and U15046 (N_15046,N_14780,N_14981);
xor U15047 (N_15047,N_14777,N_14943);
or U15048 (N_15048,N_14775,N_14828);
nor U15049 (N_15049,N_14844,N_14846);
and U15050 (N_15050,N_14737,N_14725);
nand U15051 (N_15051,N_14986,N_14816);
nand U15052 (N_15052,N_14896,N_14925);
xnor U15053 (N_15053,N_14903,N_14761);
xor U15054 (N_15054,N_14967,N_14760);
nand U15055 (N_15055,N_14764,N_14714);
xor U15056 (N_15056,N_14802,N_14946);
xor U15057 (N_15057,N_14983,N_14917);
and U15058 (N_15058,N_14750,N_14740);
nor U15059 (N_15059,N_14836,N_14932);
xnor U15060 (N_15060,N_14808,N_14838);
xor U15061 (N_15061,N_14868,N_14803);
nand U15062 (N_15062,N_14918,N_14971);
nand U15063 (N_15063,N_14842,N_14794);
nor U15064 (N_15064,N_14910,N_14921);
xor U15065 (N_15065,N_14707,N_14960);
and U15066 (N_15066,N_14934,N_14845);
xor U15067 (N_15067,N_14938,N_14859);
nor U15068 (N_15068,N_14916,N_14927);
nand U15069 (N_15069,N_14913,N_14823);
nand U15070 (N_15070,N_14881,N_14721);
and U15071 (N_15071,N_14758,N_14982);
xor U15072 (N_15072,N_14817,N_14747);
nand U15073 (N_15073,N_14814,N_14847);
nor U15074 (N_15074,N_14968,N_14834);
nor U15075 (N_15075,N_14793,N_14751);
or U15076 (N_15076,N_14890,N_14984);
and U15077 (N_15077,N_14807,N_14757);
xor U15078 (N_15078,N_14857,N_14988);
nand U15079 (N_15079,N_14774,N_14743);
xor U15080 (N_15080,N_14877,N_14790);
and U15081 (N_15081,N_14933,N_14990);
and U15082 (N_15082,N_14825,N_14824);
or U15083 (N_15083,N_14978,N_14879);
xnor U15084 (N_15084,N_14850,N_14952);
and U15085 (N_15085,N_14831,N_14724);
nand U15086 (N_15086,N_14855,N_14869);
or U15087 (N_15087,N_14871,N_14948);
xor U15088 (N_15088,N_14703,N_14940);
or U15089 (N_15089,N_14700,N_14880);
or U15090 (N_15090,N_14853,N_14969);
nand U15091 (N_15091,N_14957,N_14922);
or U15092 (N_15092,N_14815,N_14949);
and U15093 (N_15093,N_14892,N_14975);
xnor U15094 (N_15094,N_14800,N_14928);
xor U15095 (N_15095,N_14937,N_14964);
and U15096 (N_15096,N_14977,N_14783);
xnor U15097 (N_15097,N_14966,N_14862);
xnor U15098 (N_15098,N_14954,N_14711);
or U15099 (N_15099,N_14766,N_14970);
and U15100 (N_15100,N_14963,N_14792);
nor U15101 (N_15101,N_14796,N_14899);
or U15102 (N_15102,N_14806,N_14749);
or U15103 (N_15103,N_14778,N_14729);
or U15104 (N_15104,N_14878,N_14789);
and U15105 (N_15105,N_14897,N_14996);
or U15106 (N_15106,N_14798,N_14935);
nand U15107 (N_15107,N_14710,N_14974);
or U15108 (N_15108,N_14704,N_14865);
nor U15109 (N_15109,N_14874,N_14947);
xor U15110 (N_15110,N_14924,N_14776);
xor U15111 (N_15111,N_14962,N_14768);
nand U15112 (N_15112,N_14791,N_14835);
and U15113 (N_15113,N_14936,N_14870);
nor U15114 (N_15114,N_14861,N_14809);
xor U15115 (N_15115,N_14723,N_14773);
nand U15116 (N_15116,N_14718,N_14827);
or U15117 (N_15117,N_14801,N_14976);
nand U15118 (N_15118,N_14891,N_14942);
nor U15119 (N_15119,N_14955,N_14730);
and U15120 (N_15120,N_14810,N_14754);
or U15121 (N_15121,N_14858,N_14872);
nor U15122 (N_15122,N_14839,N_14731);
xnor U15123 (N_15123,N_14769,N_14821);
and U15124 (N_15124,N_14854,N_14848);
xor U15125 (N_15125,N_14826,N_14884);
and U15126 (N_15126,N_14919,N_14746);
and U15127 (N_15127,N_14926,N_14905);
and U15128 (N_15128,N_14849,N_14893);
nor U15129 (N_15129,N_14876,N_14736);
nor U15130 (N_15130,N_14840,N_14784);
xnor U15131 (N_15131,N_14860,N_14735);
xor U15132 (N_15132,N_14762,N_14973);
and U15133 (N_15133,N_14989,N_14739);
xor U15134 (N_15134,N_14911,N_14956);
xor U15135 (N_15135,N_14886,N_14887);
xnor U15136 (N_15136,N_14788,N_14832);
nor U15137 (N_15137,N_14752,N_14961);
and U15138 (N_15138,N_14708,N_14856);
nor U15139 (N_15139,N_14901,N_14702);
nor U15140 (N_15140,N_14829,N_14716);
nor U15141 (N_15141,N_14979,N_14995);
or U15142 (N_15142,N_14863,N_14782);
nor U15143 (N_15143,N_14837,N_14742);
nor U15144 (N_15144,N_14991,N_14914);
or U15145 (N_15145,N_14745,N_14972);
and U15146 (N_15146,N_14841,N_14770);
or U15147 (N_15147,N_14819,N_14733);
and U15148 (N_15148,N_14786,N_14997);
or U15149 (N_15149,N_14756,N_14843);
nor U15150 (N_15150,N_14992,N_14960);
and U15151 (N_15151,N_14901,N_14928);
nor U15152 (N_15152,N_14954,N_14701);
xnor U15153 (N_15153,N_14780,N_14928);
or U15154 (N_15154,N_14986,N_14757);
nand U15155 (N_15155,N_14827,N_14830);
or U15156 (N_15156,N_14911,N_14779);
nand U15157 (N_15157,N_14934,N_14765);
xnor U15158 (N_15158,N_14915,N_14876);
nand U15159 (N_15159,N_14798,N_14896);
and U15160 (N_15160,N_14914,N_14903);
or U15161 (N_15161,N_14796,N_14971);
nor U15162 (N_15162,N_14966,N_14777);
and U15163 (N_15163,N_14903,N_14973);
nor U15164 (N_15164,N_14896,N_14759);
xor U15165 (N_15165,N_14827,N_14885);
or U15166 (N_15166,N_14821,N_14897);
xor U15167 (N_15167,N_14960,N_14702);
xor U15168 (N_15168,N_14991,N_14971);
nor U15169 (N_15169,N_14791,N_14755);
nor U15170 (N_15170,N_14840,N_14788);
or U15171 (N_15171,N_14943,N_14787);
and U15172 (N_15172,N_14846,N_14943);
and U15173 (N_15173,N_14863,N_14866);
nor U15174 (N_15174,N_14816,N_14988);
nand U15175 (N_15175,N_14961,N_14824);
or U15176 (N_15176,N_14985,N_14719);
nand U15177 (N_15177,N_14712,N_14839);
nand U15178 (N_15178,N_14705,N_14784);
xnor U15179 (N_15179,N_14882,N_14919);
and U15180 (N_15180,N_14759,N_14823);
xor U15181 (N_15181,N_14758,N_14907);
or U15182 (N_15182,N_14877,N_14981);
and U15183 (N_15183,N_14734,N_14931);
nor U15184 (N_15184,N_14889,N_14874);
or U15185 (N_15185,N_14829,N_14943);
nand U15186 (N_15186,N_14773,N_14984);
or U15187 (N_15187,N_14781,N_14866);
xor U15188 (N_15188,N_14837,N_14834);
nor U15189 (N_15189,N_14719,N_14914);
and U15190 (N_15190,N_14738,N_14890);
nand U15191 (N_15191,N_14823,N_14857);
and U15192 (N_15192,N_14959,N_14772);
and U15193 (N_15193,N_14788,N_14756);
nand U15194 (N_15194,N_14911,N_14933);
or U15195 (N_15195,N_14860,N_14932);
nor U15196 (N_15196,N_14723,N_14906);
xnor U15197 (N_15197,N_14894,N_14810);
or U15198 (N_15198,N_14883,N_14926);
nor U15199 (N_15199,N_14782,N_14734);
nor U15200 (N_15200,N_14973,N_14879);
and U15201 (N_15201,N_14733,N_14990);
or U15202 (N_15202,N_14817,N_14800);
xnor U15203 (N_15203,N_14870,N_14779);
nand U15204 (N_15204,N_14937,N_14898);
or U15205 (N_15205,N_14943,N_14788);
nand U15206 (N_15206,N_14946,N_14836);
nor U15207 (N_15207,N_14873,N_14711);
xor U15208 (N_15208,N_14998,N_14758);
nand U15209 (N_15209,N_14815,N_14792);
and U15210 (N_15210,N_14830,N_14933);
nor U15211 (N_15211,N_14935,N_14768);
nor U15212 (N_15212,N_14852,N_14762);
nand U15213 (N_15213,N_14729,N_14992);
nand U15214 (N_15214,N_14989,N_14718);
or U15215 (N_15215,N_14814,N_14918);
or U15216 (N_15216,N_14949,N_14922);
nor U15217 (N_15217,N_14731,N_14748);
nand U15218 (N_15218,N_14987,N_14801);
nand U15219 (N_15219,N_14870,N_14988);
xor U15220 (N_15220,N_14729,N_14919);
nand U15221 (N_15221,N_14954,N_14881);
xor U15222 (N_15222,N_14825,N_14812);
or U15223 (N_15223,N_14968,N_14966);
or U15224 (N_15224,N_14785,N_14722);
nor U15225 (N_15225,N_14798,N_14773);
or U15226 (N_15226,N_14933,N_14895);
or U15227 (N_15227,N_14920,N_14975);
nand U15228 (N_15228,N_14829,N_14887);
nor U15229 (N_15229,N_14996,N_14708);
xor U15230 (N_15230,N_14755,N_14921);
xnor U15231 (N_15231,N_14872,N_14964);
xnor U15232 (N_15232,N_14916,N_14757);
nand U15233 (N_15233,N_14774,N_14839);
nand U15234 (N_15234,N_14837,N_14991);
nor U15235 (N_15235,N_14857,N_14999);
xnor U15236 (N_15236,N_14771,N_14763);
nor U15237 (N_15237,N_14981,N_14746);
and U15238 (N_15238,N_14884,N_14793);
nor U15239 (N_15239,N_14842,N_14792);
and U15240 (N_15240,N_14797,N_14879);
or U15241 (N_15241,N_14907,N_14813);
nand U15242 (N_15242,N_14992,N_14782);
xnor U15243 (N_15243,N_14837,N_14935);
nor U15244 (N_15244,N_14712,N_14858);
nand U15245 (N_15245,N_14844,N_14960);
xnor U15246 (N_15246,N_14798,N_14811);
and U15247 (N_15247,N_14838,N_14875);
nand U15248 (N_15248,N_14860,N_14924);
nor U15249 (N_15249,N_14780,N_14921);
nand U15250 (N_15250,N_14903,N_14797);
nor U15251 (N_15251,N_14978,N_14997);
nor U15252 (N_15252,N_14745,N_14866);
nand U15253 (N_15253,N_14710,N_14866);
xor U15254 (N_15254,N_14715,N_14839);
xnor U15255 (N_15255,N_14862,N_14749);
xor U15256 (N_15256,N_14875,N_14957);
nor U15257 (N_15257,N_14853,N_14799);
nand U15258 (N_15258,N_14979,N_14906);
nand U15259 (N_15259,N_14755,N_14768);
nor U15260 (N_15260,N_14950,N_14938);
or U15261 (N_15261,N_14896,N_14841);
nand U15262 (N_15262,N_14822,N_14850);
nor U15263 (N_15263,N_14936,N_14739);
nand U15264 (N_15264,N_14922,N_14804);
or U15265 (N_15265,N_14985,N_14714);
nor U15266 (N_15266,N_14928,N_14741);
and U15267 (N_15267,N_14743,N_14978);
and U15268 (N_15268,N_14910,N_14834);
xor U15269 (N_15269,N_14747,N_14860);
and U15270 (N_15270,N_14923,N_14906);
nor U15271 (N_15271,N_14793,N_14713);
nand U15272 (N_15272,N_14732,N_14983);
and U15273 (N_15273,N_14731,N_14824);
or U15274 (N_15274,N_14980,N_14800);
and U15275 (N_15275,N_14755,N_14751);
nand U15276 (N_15276,N_14983,N_14820);
nand U15277 (N_15277,N_14874,N_14701);
nor U15278 (N_15278,N_14731,N_14983);
or U15279 (N_15279,N_14733,N_14915);
nor U15280 (N_15280,N_14909,N_14892);
nor U15281 (N_15281,N_14984,N_14994);
xor U15282 (N_15282,N_14803,N_14981);
nor U15283 (N_15283,N_14833,N_14947);
and U15284 (N_15284,N_14771,N_14870);
xor U15285 (N_15285,N_14716,N_14941);
nand U15286 (N_15286,N_14731,N_14710);
and U15287 (N_15287,N_14979,N_14884);
and U15288 (N_15288,N_14796,N_14725);
and U15289 (N_15289,N_14783,N_14806);
nor U15290 (N_15290,N_14748,N_14977);
nand U15291 (N_15291,N_14793,N_14879);
or U15292 (N_15292,N_14766,N_14816);
nor U15293 (N_15293,N_14818,N_14700);
nor U15294 (N_15294,N_14856,N_14847);
nand U15295 (N_15295,N_14844,N_14835);
xor U15296 (N_15296,N_14757,N_14987);
and U15297 (N_15297,N_14882,N_14997);
or U15298 (N_15298,N_14796,N_14888);
xnor U15299 (N_15299,N_14951,N_14880);
and U15300 (N_15300,N_15242,N_15151);
nor U15301 (N_15301,N_15077,N_15032);
nand U15302 (N_15302,N_15196,N_15218);
xnor U15303 (N_15303,N_15094,N_15237);
or U15304 (N_15304,N_15098,N_15116);
nand U15305 (N_15305,N_15229,N_15035);
xor U15306 (N_15306,N_15187,N_15292);
or U15307 (N_15307,N_15043,N_15093);
and U15308 (N_15308,N_15288,N_15066);
and U15309 (N_15309,N_15248,N_15265);
xor U15310 (N_15310,N_15123,N_15080);
nand U15311 (N_15311,N_15230,N_15029);
and U15312 (N_15312,N_15165,N_15294);
and U15313 (N_15313,N_15212,N_15289);
xnor U15314 (N_15314,N_15100,N_15130);
or U15315 (N_15315,N_15023,N_15156);
nor U15316 (N_15316,N_15221,N_15086);
nor U15317 (N_15317,N_15026,N_15287);
nand U15318 (N_15318,N_15008,N_15259);
nor U15319 (N_15319,N_15233,N_15075);
nor U15320 (N_15320,N_15183,N_15190);
and U15321 (N_15321,N_15181,N_15079);
and U15322 (N_15322,N_15296,N_15074);
nand U15323 (N_15323,N_15214,N_15009);
and U15324 (N_15324,N_15042,N_15127);
xnor U15325 (N_15325,N_15092,N_15231);
and U15326 (N_15326,N_15217,N_15089);
xor U15327 (N_15327,N_15076,N_15063);
or U15328 (N_15328,N_15238,N_15108);
or U15329 (N_15329,N_15247,N_15112);
nand U15330 (N_15330,N_15203,N_15131);
xnor U15331 (N_15331,N_15251,N_15166);
nand U15332 (N_15332,N_15284,N_15021);
nor U15333 (N_15333,N_15149,N_15096);
and U15334 (N_15334,N_15117,N_15260);
or U15335 (N_15335,N_15264,N_15227);
nand U15336 (N_15336,N_15107,N_15038);
xor U15337 (N_15337,N_15213,N_15083);
or U15338 (N_15338,N_15073,N_15139);
nand U15339 (N_15339,N_15215,N_15241);
xnor U15340 (N_15340,N_15223,N_15144);
nand U15341 (N_15341,N_15102,N_15004);
nand U15342 (N_15342,N_15087,N_15252);
or U15343 (N_15343,N_15201,N_15095);
xnor U15344 (N_15344,N_15244,N_15148);
xor U15345 (N_15345,N_15271,N_15268);
nand U15346 (N_15346,N_15031,N_15145);
nor U15347 (N_15347,N_15298,N_15054);
and U15348 (N_15348,N_15068,N_15153);
xnor U15349 (N_15349,N_15273,N_15200);
or U15350 (N_15350,N_15034,N_15245);
or U15351 (N_15351,N_15055,N_15278);
and U15352 (N_15352,N_15113,N_15006);
and U15353 (N_15353,N_15143,N_15180);
xor U15354 (N_15354,N_15125,N_15224);
or U15355 (N_15355,N_15277,N_15137);
and U15356 (N_15356,N_15118,N_15085);
and U15357 (N_15357,N_15140,N_15184);
xor U15358 (N_15358,N_15136,N_15071);
and U15359 (N_15359,N_15266,N_15062);
xnor U15360 (N_15360,N_15164,N_15236);
nand U15361 (N_15361,N_15082,N_15047);
xor U15362 (N_15362,N_15276,N_15222);
nand U15363 (N_15363,N_15010,N_15036);
or U15364 (N_15364,N_15186,N_15104);
or U15365 (N_15365,N_15120,N_15141);
nor U15366 (N_15366,N_15163,N_15013);
nor U15367 (N_15367,N_15262,N_15020);
nor U15368 (N_15368,N_15007,N_15030);
or U15369 (N_15369,N_15056,N_15174);
nor U15370 (N_15370,N_15158,N_15282);
nand U15371 (N_15371,N_15015,N_15161);
or U15372 (N_15372,N_15293,N_15255);
nor U15373 (N_15373,N_15177,N_15129);
and U15374 (N_15374,N_15270,N_15099);
xor U15375 (N_15375,N_15016,N_15059);
nor U15376 (N_15376,N_15065,N_15115);
nand U15377 (N_15377,N_15199,N_15235);
and U15378 (N_15378,N_15189,N_15297);
nand U15379 (N_15379,N_15061,N_15272);
and U15380 (N_15380,N_15128,N_15005);
nor U15381 (N_15381,N_15103,N_15012);
xnor U15382 (N_15382,N_15001,N_15246);
nor U15383 (N_15383,N_15147,N_15053);
nor U15384 (N_15384,N_15135,N_15159);
xor U15385 (N_15385,N_15220,N_15088);
nor U15386 (N_15386,N_15188,N_15160);
xor U15387 (N_15387,N_15206,N_15041);
nor U15388 (N_15388,N_15173,N_15003);
nor U15389 (N_15389,N_15044,N_15150);
nor U15390 (N_15390,N_15046,N_15033);
xnor U15391 (N_15391,N_15138,N_15170);
or U15392 (N_15392,N_15225,N_15195);
xor U15393 (N_15393,N_15208,N_15169);
nand U15394 (N_15394,N_15011,N_15258);
nand U15395 (N_15395,N_15263,N_15072);
nor U15396 (N_15396,N_15198,N_15014);
xnor U15397 (N_15397,N_15280,N_15228);
nand U15398 (N_15398,N_15191,N_15142);
xnor U15399 (N_15399,N_15179,N_15097);
or U15400 (N_15400,N_15018,N_15279);
or U15401 (N_15401,N_15205,N_15050);
and U15402 (N_15402,N_15240,N_15257);
or U15403 (N_15403,N_15267,N_15070);
nand U15404 (N_15404,N_15204,N_15154);
nand U15405 (N_15405,N_15106,N_15261);
or U15406 (N_15406,N_15175,N_15226);
xor U15407 (N_15407,N_15167,N_15022);
nand U15408 (N_15408,N_15048,N_15197);
nand U15409 (N_15409,N_15162,N_15024);
or U15410 (N_15410,N_15124,N_15114);
nor U15411 (N_15411,N_15134,N_15152);
xor U15412 (N_15412,N_15239,N_15019);
and U15413 (N_15413,N_15194,N_15045);
xnor U15414 (N_15414,N_15101,N_15078);
xor U15415 (N_15415,N_15254,N_15052);
or U15416 (N_15416,N_15040,N_15269);
xor U15417 (N_15417,N_15295,N_15049);
xor U15418 (N_15418,N_15234,N_15126);
nor U15419 (N_15419,N_15090,N_15105);
or U15420 (N_15420,N_15219,N_15111);
nor U15421 (N_15421,N_15275,N_15146);
and U15422 (N_15422,N_15067,N_15202);
nand U15423 (N_15423,N_15171,N_15028);
and U15424 (N_15424,N_15286,N_15025);
and U15425 (N_15425,N_15249,N_15176);
nand U15426 (N_15426,N_15243,N_15002);
nor U15427 (N_15427,N_15256,N_15274);
nand U15428 (N_15428,N_15069,N_15133);
and U15429 (N_15429,N_15157,N_15172);
xor U15430 (N_15430,N_15121,N_15091);
nand U15431 (N_15431,N_15178,N_15017);
and U15432 (N_15432,N_15182,N_15207);
nor U15433 (N_15433,N_15253,N_15060);
and U15434 (N_15434,N_15281,N_15193);
or U15435 (N_15435,N_15210,N_15283);
nand U15436 (N_15436,N_15192,N_15211);
nand U15437 (N_15437,N_15291,N_15037);
or U15438 (N_15438,N_15185,N_15081);
nor U15439 (N_15439,N_15122,N_15232);
nor U15440 (N_15440,N_15084,N_15039);
nand U15441 (N_15441,N_15285,N_15119);
nand U15442 (N_15442,N_15110,N_15299);
and U15443 (N_15443,N_15155,N_15250);
nand U15444 (N_15444,N_15109,N_15051);
nor U15445 (N_15445,N_15209,N_15168);
or U15446 (N_15446,N_15064,N_15216);
nand U15447 (N_15447,N_15027,N_15000);
xor U15448 (N_15448,N_15290,N_15058);
nor U15449 (N_15449,N_15057,N_15132);
and U15450 (N_15450,N_15165,N_15146);
or U15451 (N_15451,N_15263,N_15122);
nand U15452 (N_15452,N_15238,N_15065);
xor U15453 (N_15453,N_15174,N_15237);
nor U15454 (N_15454,N_15091,N_15278);
and U15455 (N_15455,N_15281,N_15288);
nor U15456 (N_15456,N_15192,N_15257);
nand U15457 (N_15457,N_15105,N_15162);
nor U15458 (N_15458,N_15296,N_15121);
xor U15459 (N_15459,N_15258,N_15124);
and U15460 (N_15460,N_15007,N_15264);
and U15461 (N_15461,N_15200,N_15140);
and U15462 (N_15462,N_15147,N_15145);
or U15463 (N_15463,N_15152,N_15191);
nand U15464 (N_15464,N_15111,N_15043);
xnor U15465 (N_15465,N_15059,N_15121);
nor U15466 (N_15466,N_15228,N_15174);
xor U15467 (N_15467,N_15253,N_15223);
nor U15468 (N_15468,N_15130,N_15121);
and U15469 (N_15469,N_15172,N_15233);
nor U15470 (N_15470,N_15255,N_15290);
or U15471 (N_15471,N_15033,N_15198);
nor U15472 (N_15472,N_15220,N_15141);
xor U15473 (N_15473,N_15267,N_15298);
and U15474 (N_15474,N_15243,N_15028);
and U15475 (N_15475,N_15234,N_15227);
nand U15476 (N_15476,N_15128,N_15160);
or U15477 (N_15477,N_15147,N_15005);
nor U15478 (N_15478,N_15284,N_15134);
xnor U15479 (N_15479,N_15280,N_15132);
or U15480 (N_15480,N_15270,N_15178);
xor U15481 (N_15481,N_15041,N_15192);
or U15482 (N_15482,N_15044,N_15057);
nor U15483 (N_15483,N_15249,N_15136);
nand U15484 (N_15484,N_15234,N_15112);
xnor U15485 (N_15485,N_15177,N_15172);
nand U15486 (N_15486,N_15258,N_15007);
and U15487 (N_15487,N_15294,N_15048);
or U15488 (N_15488,N_15129,N_15148);
xor U15489 (N_15489,N_15212,N_15046);
nor U15490 (N_15490,N_15185,N_15211);
xnor U15491 (N_15491,N_15159,N_15254);
nor U15492 (N_15492,N_15278,N_15010);
nand U15493 (N_15493,N_15009,N_15100);
nor U15494 (N_15494,N_15143,N_15144);
nor U15495 (N_15495,N_15139,N_15120);
nor U15496 (N_15496,N_15134,N_15097);
and U15497 (N_15497,N_15251,N_15151);
xnor U15498 (N_15498,N_15103,N_15059);
and U15499 (N_15499,N_15018,N_15196);
and U15500 (N_15500,N_15247,N_15270);
nand U15501 (N_15501,N_15221,N_15277);
nor U15502 (N_15502,N_15133,N_15094);
and U15503 (N_15503,N_15238,N_15073);
xor U15504 (N_15504,N_15042,N_15072);
and U15505 (N_15505,N_15011,N_15080);
or U15506 (N_15506,N_15009,N_15124);
nor U15507 (N_15507,N_15239,N_15203);
and U15508 (N_15508,N_15230,N_15191);
nand U15509 (N_15509,N_15263,N_15227);
nand U15510 (N_15510,N_15056,N_15239);
nand U15511 (N_15511,N_15243,N_15123);
or U15512 (N_15512,N_15052,N_15190);
or U15513 (N_15513,N_15249,N_15100);
xor U15514 (N_15514,N_15030,N_15228);
or U15515 (N_15515,N_15257,N_15176);
xor U15516 (N_15516,N_15054,N_15261);
xnor U15517 (N_15517,N_15166,N_15201);
xor U15518 (N_15518,N_15104,N_15257);
nand U15519 (N_15519,N_15128,N_15076);
nand U15520 (N_15520,N_15130,N_15249);
and U15521 (N_15521,N_15215,N_15109);
and U15522 (N_15522,N_15034,N_15244);
nand U15523 (N_15523,N_15240,N_15239);
xnor U15524 (N_15524,N_15212,N_15008);
xor U15525 (N_15525,N_15114,N_15188);
and U15526 (N_15526,N_15032,N_15024);
nand U15527 (N_15527,N_15127,N_15209);
or U15528 (N_15528,N_15238,N_15188);
nand U15529 (N_15529,N_15111,N_15197);
or U15530 (N_15530,N_15116,N_15071);
nand U15531 (N_15531,N_15296,N_15010);
and U15532 (N_15532,N_15038,N_15291);
and U15533 (N_15533,N_15298,N_15161);
nand U15534 (N_15534,N_15064,N_15072);
and U15535 (N_15535,N_15135,N_15228);
xnor U15536 (N_15536,N_15261,N_15253);
or U15537 (N_15537,N_15057,N_15275);
nand U15538 (N_15538,N_15018,N_15174);
nor U15539 (N_15539,N_15203,N_15133);
nand U15540 (N_15540,N_15129,N_15244);
xnor U15541 (N_15541,N_15278,N_15049);
or U15542 (N_15542,N_15120,N_15054);
xor U15543 (N_15543,N_15021,N_15283);
xor U15544 (N_15544,N_15203,N_15155);
and U15545 (N_15545,N_15036,N_15235);
nor U15546 (N_15546,N_15299,N_15170);
or U15547 (N_15547,N_15249,N_15038);
nor U15548 (N_15548,N_15089,N_15047);
and U15549 (N_15549,N_15024,N_15183);
and U15550 (N_15550,N_15229,N_15081);
nand U15551 (N_15551,N_15066,N_15071);
and U15552 (N_15552,N_15000,N_15181);
nand U15553 (N_15553,N_15130,N_15219);
nor U15554 (N_15554,N_15032,N_15017);
xnor U15555 (N_15555,N_15002,N_15069);
xor U15556 (N_15556,N_15156,N_15258);
or U15557 (N_15557,N_15090,N_15109);
nor U15558 (N_15558,N_15166,N_15264);
nor U15559 (N_15559,N_15173,N_15004);
xor U15560 (N_15560,N_15145,N_15183);
and U15561 (N_15561,N_15244,N_15156);
or U15562 (N_15562,N_15261,N_15193);
xnor U15563 (N_15563,N_15111,N_15243);
nand U15564 (N_15564,N_15065,N_15205);
xnor U15565 (N_15565,N_15217,N_15265);
nor U15566 (N_15566,N_15160,N_15045);
xor U15567 (N_15567,N_15134,N_15110);
xnor U15568 (N_15568,N_15122,N_15030);
nor U15569 (N_15569,N_15048,N_15239);
or U15570 (N_15570,N_15157,N_15202);
nor U15571 (N_15571,N_15121,N_15105);
nand U15572 (N_15572,N_15048,N_15012);
or U15573 (N_15573,N_15083,N_15071);
xor U15574 (N_15574,N_15068,N_15094);
xnor U15575 (N_15575,N_15188,N_15075);
nand U15576 (N_15576,N_15284,N_15190);
nor U15577 (N_15577,N_15223,N_15035);
xor U15578 (N_15578,N_15284,N_15017);
xor U15579 (N_15579,N_15197,N_15010);
xor U15580 (N_15580,N_15248,N_15122);
xor U15581 (N_15581,N_15203,N_15186);
nand U15582 (N_15582,N_15144,N_15212);
and U15583 (N_15583,N_15083,N_15107);
nand U15584 (N_15584,N_15016,N_15268);
and U15585 (N_15585,N_15165,N_15288);
and U15586 (N_15586,N_15173,N_15165);
nand U15587 (N_15587,N_15083,N_15030);
nor U15588 (N_15588,N_15043,N_15071);
xor U15589 (N_15589,N_15023,N_15022);
and U15590 (N_15590,N_15284,N_15025);
nor U15591 (N_15591,N_15251,N_15229);
or U15592 (N_15592,N_15246,N_15195);
xnor U15593 (N_15593,N_15020,N_15230);
xnor U15594 (N_15594,N_15009,N_15199);
and U15595 (N_15595,N_15051,N_15010);
or U15596 (N_15596,N_15050,N_15222);
xnor U15597 (N_15597,N_15140,N_15173);
xnor U15598 (N_15598,N_15081,N_15055);
xnor U15599 (N_15599,N_15039,N_15171);
nand U15600 (N_15600,N_15552,N_15377);
nor U15601 (N_15601,N_15494,N_15595);
or U15602 (N_15602,N_15329,N_15499);
and U15603 (N_15603,N_15566,N_15526);
nor U15604 (N_15604,N_15445,N_15375);
or U15605 (N_15605,N_15484,N_15575);
nand U15606 (N_15606,N_15585,N_15343);
xnor U15607 (N_15607,N_15503,N_15596);
and U15608 (N_15608,N_15332,N_15455);
or U15609 (N_15609,N_15515,N_15330);
nor U15610 (N_15610,N_15392,N_15589);
and U15611 (N_15611,N_15504,N_15486);
and U15612 (N_15612,N_15367,N_15374);
nor U15613 (N_15613,N_15417,N_15338);
or U15614 (N_15614,N_15557,N_15317);
and U15615 (N_15615,N_15598,N_15413);
or U15616 (N_15616,N_15453,N_15387);
nor U15617 (N_15617,N_15364,N_15522);
nor U15618 (N_15618,N_15542,N_15406);
nor U15619 (N_15619,N_15373,N_15433);
xor U15620 (N_15620,N_15449,N_15501);
nand U15621 (N_15621,N_15578,N_15422);
nand U15622 (N_15622,N_15335,N_15593);
nand U15623 (N_15623,N_15415,N_15544);
nand U15624 (N_15624,N_15310,N_15462);
or U15625 (N_15625,N_15381,N_15410);
nor U15626 (N_15626,N_15480,N_15309);
or U15627 (N_15627,N_15320,N_15394);
nand U15628 (N_15628,N_15372,N_15446);
nor U15629 (N_15629,N_15371,N_15326);
or U15630 (N_15630,N_15519,N_15531);
or U15631 (N_15631,N_15431,N_15590);
nand U15632 (N_15632,N_15349,N_15420);
and U15633 (N_15633,N_15354,N_15489);
and U15634 (N_15634,N_15506,N_15458);
xnor U15635 (N_15635,N_15380,N_15540);
or U15636 (N_15636,N_15481,N_15399);
xnor U15637 (N_15637,N_15398,N_15450);
and U15638 (N_15638,N_15305,N_15586);
xor U15639 (N_15639,N_15581,N_15565);
or U15640 (N_15640,N_15512,N_15571);
xnor U15641 (N_15641,N_15348,N_15313);
and U15642 (N_15642,N_15302,N_15334);
or U15643 (N_15643,N_15390,N_15591);
nor U15644 (N_15644,N_15548,N_15533);
or U15645 (N_15645,N_15437,N_15535);
or U15646 (N_15646,N_15430,N_15572);
nor U15647 (N_15647,N_15474,N_15439);
nor U15648 (N_15648,N_15477,N_15322);
nor U15649 (N_15649,N_15307,N_15304);
nor U15650 (N_15650,N_15541,N_15525);
and U15651 (N_15651,N_15385,N_15358);
and U15652 (N_15652,N_15550,N_15356);
nand U15653 (N_15653,N_15391,N_15587);
or U15654 (N_15654,N_15321,N_15493);
or U15655 (N_15655,N_15341,N_15397);
and U15656 (N_15656,N_15551,N_15303);
nor U15657 (N_15657,N_15404,N_15538);
nor U15658 (N_15658,N_15312,N_15537);
and U15659 (N_15659,N_15470,N_15363);
nand U15660 (N_15660,N_15547,N_15523);
and U15661 (N_15661,N_15574,N_15558);
xnor U15662 (N_15662,N_15436,N_15520);
or U15663 (N_15663,N_15543,N_15554);
or U15664 (N_15664,N_15418,N_15340);
nor U15665 (N_15665,N_15314,N_15528);
nor U15666 (N_15666,N_15301,N_15393);
and U15667 (N_15667,N_15524,N_15403);
nand U15668 (N_15668,N_15564,N_15510);
nand U15669 (N_15669,N_15383,N_15389);
and U15670 (N_15670,N_15475,N_15459);
nor U15671 (N_15671,N_15511,N_15376);
and U15672 (N_15672,N_15419,N_15402);
nor U15673 (N_15673,N_15467,N_15315);
nand U15674 (N_15674,N_15434,N_15382);
or U15675 (N_15675,N_15577,N_15432);
nor U15676 (N_15676,N_15479,N_15333);
and U15677 (N_15677,N_15388,N_15411);
nand U15678 (N_15678,N_15563,N_15583);
nand U15679 (N_15679,N_15345,N_15507);
nand U15680 (N_15680,N_15549,N_15318);
nand U15681 (N_15681,N_15441,N_15461);
xor U15682 (N_15682,N_15408,N_15412);
or U15683 (N_15683,N_15560,N_15357);
xnor U15684 (N_15684,N_15319,N_15440);
or U15685 (N_15685,N_15324,N_15546);
nand U15686 (N_15686,N_15460,N_15407);
nor U15687 (N_15687,N_15556,N_15352);
or U15688 (N_15688,N_15346,N_15469);
xor U15689 (N_15689,N_15514,N_15342);
or U15690 (N_15690,N_15495,N_15360);
nand U15691 (N_15691,N_15478,N_15456);
xnor U15692 (N_15692,N_15534,N_15444);
xor U15693 (N_15693,N_15328,N_15428);
xnor U15694 (N_15694,N_15457,N_15414);
and U15695 (N_15695,N_15353,N_15502);
nor U15696 (N_15696,N_15508,N_15421);
nor U15697 (N_15697,N_15435,N_15569);
or U15698 (N_15698,N_15487,N_15366);
xnor U15699 (N_15699,N_15573,N_15347);
xor U15700 (N_15700,N_15579,N_15466);
nor U15701 (N_15701,N_15311,N_15369);
xor U15702 (N_15702,N_15454,N_15529);
or U15703 (N_15703,N_15567,N_15500);
nor U15704 (N_15704,N_15424,N_15536);
or U15705 (N_15705,N_15361,N_15427);
or U15706 (N_15706,N_15447,N_15359);
or U15707 (N_15707,N_15452,N_15473);
xor U15708 (N_15708,N_15463,N_15468);
nand U15709 (N_15709,N_15350,N_15530);
nand U15710 (N_15710,N_15497,N_15423);
and U15711 (N_15711,N_15513,N_15539);
and U15712 (N_15712,N_15599,N_15576);
and U15713 (N_15713,N_15553,N_15465);
xnor U15714 (N_15714,N_15490,N_15488);
or U15715 (N_15715,N_15555,N_15442);
nor U15716 (N_15716,N_15327,N_15344);
xor U15717 (N_15717,N_15464,N_15300);
nor U15718 (N_15718,N_15409,N_15509);
nand U15719 (N_15719,N_15443,N_15379);
or U15720 (N_15720,N_15308,N_15498);
and U15721 (N_15721,N_15492,N_15491);
nor U15722 (N_15722,N_15570,N_15448);
and U15723 (N_15723,N_15438,N_15316);
and U15724 (N_15724,N_15568,N_15368);
or U15725 (N_15725,N_15325,N_15580);
nand U15726 (N_15726,N_15323,N_15588);
nor U15727 (N_15727,N_15562,N_15396);
or U15728 (N_15728,N_15485,N_15416);
nand U15729 (N_15729,N_15386,N_15592);
and U15730 (N_15730,N_15401,N_15496);
xor U15731 (N_15731,N_15306,N_15331);
and U15732 (N_15732,N_15532,N_15594);
xnor U15733 (N_15733,N_15395,N_15521);
xor U15734 (N_15734,N_15483,N_15355);
nor U15735 (N_15735,N_15370,N_15582);
nor U15736 (N_15736,N_15425,N_15545);
nand U15737 (N_15737,N_15559,N_15365);
or U15738 (N_15738,N_15384,N_15339);
nor U15739 (N_15739,N_15561,N_15472);
nand U15740 (N_15740,N_15471,N_15378);
and U15741 (N_15741,N_15505,N_15518);
nor U15742 (N_15742,N_15400,N_15405);
xor U15743 (N_15743,N_15584,N_15476);
xor U15744 (N_15744,N_15362,N_15426);
or U15745 (N_15745,N_15351,N_15429);
nand U15746 (N_15746,N_15336,N_15337);
nand U15747 (N_15747,N_15451,N_15516);
nor U15748 (N_15748,N_15527,N_15517);
nand U15749 (N_15749,N_15482,N_15597);
xnor U15750 (N_15750,N_15584,N_15595);
xnor U15751 (N_15751,N_15406,N_15301);
or U15752 (N_15752,N_15354,N_15596);
nor U15753 (N_15753,N_15465,N_15424);
or U15754 (N_15754,N_15442,N_15494);
xnor U15755 (N_15755,N_15327,N_15320);
xor U15756 (N_15756,N_15395,N_15390);
or U15757 (N_15757,N_15365,N_15326);
nor U15758 (N_15758,N_15493,N_15506);
nand U15759 (N_15759,N_15402,N_15325);
nand U15760 (N_15760,N_15529,N_15330);
nor U15761 (N_15761,N_15526,N_15524);
nor U15762 (N_15762,N_15564,N_15483);
and U15763 (N_15763,N_15443,N_15344);
nor U15764 (N_15764,N_15428,N_15534);
nand U15765 (N_15765,N_15593,N_15329);
and U15766 (N_15766,N_15449,N_15511);
xor U15767 (N_15767,N_15594,N_15510);
and U15768 (N_15768,N_15323,N_15395);
nand U15769 (N_15769,N_15485,N_15469);
nor U15770 (N_15770,N_15596,N_15534);
and U15771 (N_15771,N_15311,N_15319);
and U15772 (N_15772,N_15415,N_15512);
or U15773 (N_15773,N_15599,N_15432);
nand U15774 (N_15774,N_15344,N_15418);
nor U15775 (N_15775,N_15386,N_15537);
and U15776 (N_15776,N_15345,N_15492);
xor U15777 (N_15777,N_15572,N_15598);
and U15778 (N_15778,N_15539,N_15429);
xor U15779 (N_15779,N_15418,N_15408);
and U15780 (N_15780,N_15511,N_15422);
nor U15781 (N_15781,N_15443,N_15519);
or U15782 (N_15782,N_15306,N_15506);
or U15783 (N_15783,N_15325,N_15544);
xnor U15784 (N_15784,N_15445,N_15366);
or U15785 (N_15785,N_15314,N_15372);
or U15786 (N_15786,N_15493,N_15338);
nor U15787 (N_15787,N_15390,N_15569);
nor U15788 (N_15788,N_15588,N_15457);
xnor U15789 (N_15789,N_15360,N_15446);
xnor U15790 (N_15790,N_15302,N_15470);
nor U15791 (N_15791,N_15322,N_15329);
xor U15792 (N_15792,N_15486,N_15576);
nand U15793 (N_15793,N_15508,N_15367);
nor U15794 (N_15794,N_15575,N_15538);
xnor U15795 (N_15795,N_15594,N_15414);
or U15796 (N_15796,N_15565,N_15587);
nor U15797 (N_15797,N_15318,N_15380);
and U15798 (N_15798,N_15430,N_15564);
nor U15799 (N_15799,N_15524,N_15541);
nor U15800 (N_15800,N_15369,N_15500);
nor U15801 (N_15801,N_15304,N_15552);
nand U15802 (N_15802,N_15449,N_15517);
and U15803 (N_15803,N_15346,N_15489);
nor U15804 (N_15804,N_15580,N_15381);
nor U15805 (N_15805,N_15458,N_15592);
and U15806 (N_15806,N_15574,N_15548);
nand U15807 (N_15807,N_15428,N_15446);
nand U15808 (N_15808,N_15441,N_15393);
and U15809 (N_15809,N_15479,N_15304);
nand U15810 (N_15810,N_15360,N_15565);
nor U15811 (N_15811,N_15313,N_15531);
nand U15812 (N_15812,N_15556,N_15517);
and U15813 (N_15813,N_15501,N_15573);
or U15814 (N_15814,N_15321,N_15359);
and U15815 (N_15815,N_15387,N_15536);
xnor U15816 (N_15816,N_15393,N_15448);
nor U15817 (N_15817,N_15397,N_15418);
xnor U15818 (N_15818,N_15533,N_15350);
xor U15819 (N_15819,N_15320,N_15443);
nor U15820 (N_15820,N_15505,N_15362);
xnor U15821 (N_15821,N_15493,N_15578);
and U15822 (N_15822,N_15487,N_15419);
xnor U15823 (N_15823,N_15366,N_15544);
or U15824 (N_15824,N_15415,N_15572);
xnor U15825 (N_15825,N_15552,N_15471);
nor U15826 (N_15826,N_15423,N_15478);
and U15827 (N_15827,N_15507,N_15464);
and U15828 (N_15828,N_15343,N_15379);
xor U15829 (N_15829,N_15425,N_15416);
and U15830 (N_15830,N_15570,N_15493);
or U15831 (N_15831,N_15421,N_15482);
and U15832 (N_15832,N_15465,N_15447);
nor U15833 (N_15833,N_15315,N_15414);
xnor U15834 (N_15834,N_15426,N_15480);
and U15835 (N_15835,N_15509,N_15594);
xor U15836 (N_15836,N_15584,N_15524);
nand U15837 (N_15837,N_15347,N_15427);
and U15838 (N_15838,N_15544,N_15403);
nor U15839 (N_15839,N_15515,N_15382);
xnor U15840 (N_15840,N_15370,N_15563);
xor U15841 (N_15841,N_15454,N_15371);
nor U15842 (N_15842,N_15358,N_15419);
or U15843 (N_15843,N_15476,N_15312);
and U15844 (N_15844,N_15462,N_15440);
and U15845 (N_15845,N_15439,N_15543);
nor U15846 (N_15846,N_15407,N_15484);
nor U15847 (N_15847,N_15469,N_15517);
or U15848 (N_15848,N_15561,N_15332);
and U15849 (N_15849,N_15548,N_15425);
and U15850 (N_15850,N_15507,N_15367);
or U15851 (N_15851,N_15586,N_15573);
nor U15852 (N_15852,N_15387,N_15443);
and U15853 (N_15853,N_15444,N_15384);
nand U15854 (N_15854,N_15520,N_15525);
and U15855 (N_15855,N_15399,N_15452);
xor U15856 (N_15856,N_15475,N_15569);
nand U15857 (N_15857,N_15356,N_15386);
and U15858 (N_15858,N_15356,N_15486);
or U15859 (N_15859,N_15450,N_15561);
nand U15860 (N_15860,N_15582,N_15560);
and U15861 (N_15861,N_15530,N_15574);
or U15862 (N_15862,N_15512,N_15555);
nand U15863 (N_15863,N_15478,N_15532);
nand U15864 (N_15864,N_15396,N_15518);
nor U15865 (N_15865,N_15356,N_15361);
or U15866 (N_15866,N_15371,N_15568);
xnor U15867 (N_15867,N_15458,N_15568);
nand U15868 (N_15868,N_15589,N_15407);
nor U15869 (N_15869,N_15569,N_15316);
nor U15870 (N_15870,N_15511,N_15508);
xor U15871 (N_15871,N_15365,N_15376);
nand U15872 (N_15872,N_15487,N_15496);
or U15873 (N_15873,N_15358,N_15309);
nor U15874 (N_15874,N_15346,N_15402);
and U15875 (N_15875,N_15581,N_15499);
nand U15876 (N_15876,N_15355,N_15548);
nor U15877 (N_15877,N_15381,N_15367);
or U15878 (N_15878,N_15410,N_15352);
xor U15879 (N_15879,N_15494,N_15538);
nor U15880 (N_15880,N_15522,N_15437);
nand U15881 (N_15881,N_15508,N_15527);
or U15882 (N_15882,N_15516,N_15529);
or U15883 (N_15883,N_15507,N_15373);
nand U15884 (N_15884,N_15401,N_15529);
nand U15885 (N_15885,N_15541,N_15343);
or U15886 (N_15886,N_15484,N_15340);
or U15887 (N_15887,N_15569,N_15430);
nand U15888 (N_15888,N_15540,N_15458);
or U15889 (N_15889,N_15521,N_15448);
xor U15890 (N_15890,N_15350,N_15357);
nand U15891 (N_15891,N_15457,N_15577);
nand U15892 (N_15892,N_15492,N_15523);
nor U15893 (N_15893,N_15564,N_15357);
and U15894 (N_15894,N_15598,N_15370);
nand U15895 (N_15895,N_15408,N_15574);
and U15896 (N_15896,N_15597,N_15332);
or U15897 (N_15897,N_15592,N_15379);
nor U15898 (N_15898,N_15336,N_15394);
nor U15899 (N_15899,N_15397,N_15588);
and U15900 (N_15900,N_15659,N_15889);
or U15901 (N_15901,N_15821,N_15779);
nor U15902 (N_15902,N_15605,N_15726);
nor U15903 (N_15903,N_15819,N_15891);
xor U15904 (N_15904,N_15653,N_15663);
xnor U15905 (N_15905,N_15666,N_15787);
nand U15906 (N_15906,N_15766,N_15632);
xor U15907 (N_15907,N_15865,N_15637);
nor U15908 (N_15908,N_15780,N_15796);
or U15909 (N_15909,N_15795,N_15675);
nor U15910 (N_15910,N_15898,N_15767);
and U15911 (N_15911,N_15716,N_15644);
or U15912 (N_15912,N_15661,N_15822);
xnor U15913 (N_15913,N_15629,N_15722);
xnor U15914 (N_15914,N_15652,N_15873);
and U15915 (N_15915,N_15718,N_15888);
xnor U15916 (N_15916,N_15702,N_15601);
nand U15917 (N_15917,N_15698,N_15850);
xnor U15918 (N_15918,N_15757,N_15733);
nand U15919 (N_15919,N_15893,N_15816);
and U15920 (N_15920,N_15823,N_15635);
nor U15921 (N_15921,N_15639,N_15754);
nor U15922 (N_15922,N_15619,N_15790);
xnor U15923 (N_15923,N_15805,N_15769);
or U15924 (N_15924,N_15687,N_15633);
or U15925 (N_15925,N_15781,N_15614);
xnor U15926 (N_15926,N_15774,N_15752);
or U15927 (N_15927,N_15641,N_15843);
nor U15928 (N_15928,N_15717,N_15876);
nand U15929 (N_15929,N_15669,N_15667);
xnor U15930 (N_15930,N_15673,N_15874);
xor U15931 (N_15931,N_15699,N_15734);
nor U15932 (N_15932,N_15640,N_15615);
and U15933 (N_15933,N_15768,N_15728);
xnor U15934 (N_15934,N_15806,N_15600);
and U15935 (N_15935,N_15680,N_15657);
nor U15936 (N_15936,N_15642,N_15836);
or U15937 (N_15937,N_15712,N_15606);
nand U15938 (N_15938,N_15760,N_15880);
nand U15939 (N_15939,N_15678,N_15753);
nor U15940 (N_15940,N_15801,N_15820);
nand U15941 (N_15941,N_15704,N_15895);
nand U15942 (N_15942,N_15782,N_15869);
xor U15943 (N_15943,N_15624,N_15812);
and U15944 (N_15944,N_15773,N_15839);
xnor U15945 (N_15945,N_15671,N_15685);
xor U15946 (N_15946,N_15825,N_15723);
nor U15947 (N_15947,N_15844,N_15747);
and U15948 (N_15948,N_15651,N_15677);
xnor U15949 (N_15949,N_15740,N_15604);
and U15950 (N_15950,N_15607,N_15786);
nand U15951 (N_15951,N_15725,N_15701);
and U15952 (N_15952,N_15849,N_15761);
xnor U15953 (N_15953,N_15799,N_15835);
and U15954 (N_15954,N_15602,N_15785);
nor U15955 (N_15955,N_15616,N_15867);
xor U15956 (N_15956,N_15832,N_15711);
nor U15957 (N_15957,N_15634,N_15729);
nand U15958 (N_15958,N_15755,N_15750);
and U15959 (N_15959,N_15764,N_15638);
and U15960 (N_15960,N_15828,N_15643);
or U15961 (N_15961,N_15883,N_15811);
or U15962 (N_15962,N_15877,N_15897);
and U15963 (N_15963,N_15676,N_15636);
or U15964 (N_15964,N_15628,N_15697);
nor U15965 (N_15965,N_15868,N_15703);
or U15966 (N_15966,N_15772,N_15756);
and U15967 (N_15967,N_15804,N_15608);
xnor U15968 (N_15968,N_15744,N_15784);
xor U15969 (N_15969,N_15890,N_15815);
or U15970 (N_15970,N_15885,N_15826);
xnor U15971 (N_15971,N_15739,N_15656);
xnor U15972 (N_15972,N_15700,N_15803);
nor U15973 (N_15973,N_15771,N_15846);
and U15974 (N_15974,N_15864,N_15748);
nor U15975 (N_15975,N_15834,N_15794);
nand U15976 (N_15976,N_15856,N_15899);
nand U15977 (N_15977,N_15645,N_15824);
and U15978 (N_15978,N_15791,N_15848);
or U15979 (N_15979,N_15847,N_15681);
xnor U15980 (N_15980,N_15737,N_15797);
xnor U15981 (N_15981,N_15866,N_15730);
and U15982 (N_15982,N_15751,N_15684);
xnor U15983 (N_15983,N_15618,N_15724);
nand U15984 (N_15984,N_15691,N_15875);
xnor U15985 (N_15985,N_15713,N_15617);
nor U15986 (N_15986,N_15679,N_15829);
or U15987 (N_15987,N_15738,N_15626);
and U15988 (N_15988,N_15732,N_15743);
or U15989 (N_15989,N_15705,N_15646);
xor U15990 (N_15990,N_15777,N_15841);
or U15991 (N_15991,N_15665,N_15833);
nand U15992 (N_15992,N_15783,N_15709);
nand U15993 (N_15993,N_15620,N_15655);
and U15994 (N_15994,N_15852,N_15845);
or U15995 (N_15995,N_15670,N_15683);
or U15996 (N_15996,N_15778,N_15623);
nand U15997 (N_15997,N_15647,N_15792);
nand U15998 (N_15998,N_15610,N_15818);
xnor U15999 (N_15999,N_15837,N_15692);
or U16000 (N_16000,N_15627,N_15870);
and U16001 (N_16001,N_15674,N_15727);
nor U16002 (N_16002,N_15622,N_15660);
nor U16003 (N_16003,N_15814,N_15706);
nand U16004 (N_16004,N_15860,N_15735);
or U16005 (N_16005,N_15789,N_15721);
nor U16006 (N_16006,N_15882,N_15649);
nand U16007 (N_16007,N_15621,N_15872);
xnor U16008 (N_16008,N_15631,N_15763);
or U16009 (N_16009,N_15731,N_15765);
or U16010 (N_16010,N_15887,N_15817);
nand U16011 (N_16011,N_15793,N_15892);
nand U16012 (N_16012,N_15648,N_15693);
or U16013 (N_16013,N_15625,N_15658);
nand U16014 (N_16014,N_15664,N_15749);
nand U16015 (N_16015,N_15894,N_15813);
or U16016 (N_16016,N_15830,N_15742);
and U16017 (N_16017,N_15831,N_15863);
nor U16018 (N_16018,N_15827,N_15776);
and U16019 (N_16019,N_15886,N_15720);
xnor U16020 (N_16020,N_15871,N_15858);
and U16021 (N_16021,N_15854,N_15842);
nand U16022 (N_16022,N_15609,N_15710);
or U16023 (N_16023,N_15688,N_15603);
nand U16024 (N_16024,N_15798,N_15878);
nand U16025 (N_16025,N_15775,N_15695);
nor U16026 (N_16026,N_15650,N_15809);
or U16027 (N_16027,N_15715,N_15682);
xor U16028 (N_16028,N_15851,N_15861);
xnor U16029 (N_16029,N_15714,N_15690);
xnor U16030 (N_16030,N_15630,N_15745);
xor U16031 (N_16031,N_15719,N_15800);
nand U16032 (N_16032,N_15613,N_15654);
nand U16033 (N_16033,N_15853,N_15694);
or U16034 (N_16034,N_15840,N_15881);
xor U16035 (N_16035,N_15807,N_15808);
nand U16036 (N_16036,N_15884,N_15759);
nand U16037 (N_16037,N_15862,N_15736);
xor U16038 (N_16038,N_15859,N_15857);
xnor U16039 (N_16039,N_15788,N_15896);
and U16040 (N_16040,N_15612,N_15672);
or U16041 (N_16041,N_15762,N_15696);
or U16042 (N_16042,N_15708,N_15686);
or U16043 (N_16043,N_15662,N_15707);
nand U16044 (N_16044,N_15879,N_15668);
or U16045 (N_16045,N_15741,N_15802);
and U16046 (N_16046,N_15689,N_15758);
nand U16047 (N_16047,N_15838,N_15810);
nand U16048 (N_16048,N_15855,N_15746);
xor U16049 (N_16049,N_15611,N_15770);
or U16050 (N_16050,N_15701,N_15851);
or U16051 (N_16051,N_15763,N_15792);
nand U16052 (N_16052,N_15613,N_15741);
xnor U16053 (N_16053,N_15641,N_15635);
nand U16054 (N_16054,N_15657,N_15787);
or U16055 (N_16055,N_15729,N_15703);
nand U16056 (N_16056,N_15788,N_15897);
or U16057 (N_16057,N_15618,N_15875);
nor U16058 (N_16058,N_15658,N_15887);
xor U16059 (N_16059,N_15876,N_15767);
xnor U16060 (N_16060,N_15829,N_15659);
nand U16061 (N_16061,N_15601,N_15677);
nand U16062 (N_16062,N_15741,N_15824);
and U16063 (N_16063,N_15718,N_15602);
nor U16064 (N_16064,N_15755,N_15765);
nand U16065 (N_16065,N_15810,N_15870);
nor U16066 (N_16066,N_15756,N_15622);
xnor U16067 (N_16067,N_15892,N_15834);
and U16068 (N_16068,N_15655,N_15652);
or U16069 (N_16069,N_15857,N_15708);
nor U16070 (N_16070,N_15721,N_15623);
nand U16071 (N_16071,N_15690,N_15623);
or U16072 (N_16072,N_15899,N_15794);
and U16073 (N_16073,N_15783,N_15879);
nor U16074 (N_16074,N_15886,N_15669);
or U16075 (N_16075,N_15797,N_15866);
nand U16076 (N_16076,N_15816,N_15680);
xor U16077 (N_16077,N_15800,N_15686);
xnor U16078 (N_16078,N_15688,N_15635);
nand U16079 (N_16079,N_15658,N_15791);
nand U16080 (N_16080,N_15870,N_15858);
and U16081 (N_16081,N_15649,N_15863);
and U16082 (N_16082,N_15740,N_15856);
or U16083 (N_16083,N_15673,N_15798);
nor U16084 (N_16084,N_15616,N_15720);
xnor U16085 (N_16085,N_15656,N_15881);
or U16086 (N_16086,N_15675,N_15783);
nand U16087 (N_16087,N_15830,N_15715);
nor U16088 (N_16088,N_15779,N_15643);
and U16089 (N_16089,N_15750,N_15872);
nor U16090 (N_16090,N_15632,N_15826);
nor U16091 (N_16091,N_15629,N_15809);
and U16092 (N_16092,N_15776,N_15645);
and U16093 (N_16093,N_15738,N_15769);
nor U16094 (N_16094,N_15666,N_15601);
or U16095 (N_16095,N_15654,N_15684);
xor U16096 (N_16096,N_15660,N_15895);
and U16097 (N_16097,N_15823,N_15818);
nor U16098 (N_16098,N_15863,N_15833);
or U16099 (N_16099,N_15873,N_15624);
nand U16100 (N_16100,N_15698,N_15685);
and U16101 (N_16101,N_15805,N_15739);
nor U16102 (N_16102,N_15864,N_15899);
or U16103 (N_16103,N_15668,N_15801);
nor U16104 (N_16104,N_15603,N_15658);
nor U16105 (N_16105,N_15653,N_15706);
or U16106 (N_16106,N_15740,N_15799);
and U16107 (N_16107,N_15888,N_15656);
and U16108 (N_16108,N_15856,N_15687);
nor U16109 (N_16109,N_15782,N_15634);
nor U16110 (N_16110,N_15813,N_15653);
or U16111 (N_16111,N_15896,N_15745);
or U16112 (N_16112,N_15826,N_15763);
nand U16113 (N_16113,N_15833,N_15757);
xor U16114 (N_16114,N_15897,N_15711);
or U16115 (N_16115,N_15870,N_15741);
nand U16116 (N_16116,N_15735,N_15776);
or U16117 (N_16117,N_15846,N_15861);
nand U16118 (N_16118,N_15643,N_15649);
xor U16119 (N_16119,N_15848,N_15842);
nand U16120 (N_16120,N_15808,N_15716);
or U16121 (N_16121,N_15729,N_15792);
and U16122 (N_16122,N_15800,N_15650);
xor U16123 (N_16123,N_15733,N_15715);
or U16124 (N_16124,N_15723,N_15636);
nor U16125 (N_16125,N_15793,N_15715);
and U16126 (N_16126,N_15728,N_15719);
nor U16127 (N_16127,N_15708,N_15638);
xnor U16128 (N_16128,N_15742,N_15778);
xnor U16129 (N_16129,N_15690,N_15668);
xnor U16130 (N_16130,N_15743,N_15600);
and U16131 (N_16131,N_15702,N_15799);
nor U16132 (N_16132,N_15760,N_15774);
and U16133 (N_16133,N_15796,N_15636);
nor U16134 (N_16134,N_15771,N_15697);
and U16135 (N_16135,N_15650,N_15840);
nand U16136 (N_16136,N_15610,N_15688);
nand U16137 (N_16137,N_15819,N_15763);
nor U16138 (N_16138,N_15759,N_15658);
nor U16139 (N_16139,N_15722,N_15658);
and U16140 (N_16140,N_15620,N_15695);
nand U16141 (N_16141,N_15696,N_15826);
and U16142 (N_16142,N_15841,N_15876);
or U16143 (N_16143,N_15699,N_15680);
nand U16144 (N_16144,N_15834,N_15803);
or U16145 (N_16145,N_15718,N_15740);
nand U16146 (N_16146,N_15826,N_15794);
and U16147 (N_16147,N_15862,N_15654);
and U16148 (N_16148,N_15782,N_15874);
or U16149 (N_16149,N_15863,N_15758);
nand U16150 (N_16150,N_15771,N_15852);
xor U16151 (N_16151,N_15673,N_15639);
nor U16152 (N_16152,N_15893,N_15628);
xnor U16153 (N_16153,N_15672,N_15640);
and U16154 (N_16154,N_15703,N_15735);
nor U16155 (N_16155,N_15613,N_15769);
nor U16156 (N_16156,N_15812,N_15742);
nand U16157 (N_16157,N_15896,N_15690);
xor U16158 (N_16158,N_15858,N_15837);
and U16159 (N_16159,N_15751,N_15841);
nand U16160 (N_16160,N_15838,N_15788);
xnor U16161 (N_16161,N_15881,N_15677);
nor U16162 (N_16162,N_15663,N_15640);
nand U16163 (N_16163,N_15830,N_15647);
or U16164 (N_16164,N_15871,N_15893);
nand U16165 (N_16165,N_15887,N_15782);
nand U16166 (N_16166,N_15823,N_15749);
or U16167 (N_16167,N_15870,N_15679);
or U16168 (N_16168,N_15658,N_15783);
xnor U16169 (N_16169,N_15730,N_15790);
nor U16170 (N_16170,N_15831,N_15601);
nor U16171 (N_16171,N_15709,N_15683);
and U16172 (N_16172,N_15601,N_15867);
nand U16173 (N_16173,N_15796,N_15611);
nand U16174 (N_16174,N_15618,N_15899);
and U16175 (N_16175,N_15713,N_15765);
xnor U16176 (N_16176,N_15673,N_15751);
xnor U16177 (N_16177,N_15866,N_15763);
nand U16178 (N_16178,N_15762,N_15718);
and U16179 (N_16179,N_15839,N_15722);
xnor U16180 (N_16180,N_15859,N_15825);
nor U16181 (N_16181,N_15829,N_15862);
nor U16182 (N_16182,N_15877,N_15696);
or U16183 (N_16183,N_15751,N_15715);
xor U16184 (N_16184,N_15741,N_15850);
and U16185 (N_16185,N_15729,N_15775);
or U16186 (N_16186,N_15602,N_15704);
or U16187 (N_16187,N_15723,N_15834);
nor U16188 (N_16188,N_15689,N_15628);
nand U16189 (N_16189,N_15670,N_15873);
or U16190 (N_16190,N_15835,N_15786);
nand U16191 (N_16191,N_15652,N_15807);
xnor U16192 (N_16192,N_15786,N_15667);
nor U16193 (N_16193,N_15708,N_15622);
nor U16194 (N_16194,N_15621,N_15653);
xor U16195 (N_16195,N_15720,N_15774);
nor U16196 (N_16196,N_15749,N_15776);
nor U16197 (N_16197,N_15821,N_15669);
xnor U16198 (N_16198,N_15759,N_15838);
nand U16199 (N_16199,N_15839,N_15677);
and U16200 (N_16200,N_15963,N_16180);
and U16201 (N_16201,N_15904,N_16048);
or U16202 (N_16202,N_15931,N_16013);
nor U16203 (N_16203,N_16062,N_16082);
nor U16204 (N_16204,N_16040,N_15993);
or U16205 (N_16205,N_16070,N_15906);
xor U16206 (N_16206,N_16164,N_15916);
nand U16207 (N_16207,N_15961,N_15985);
or U16208 (N_16208,N_16058,N_15950);
nand U16209 (N_16209,N_16068,N_16030);
xnor U16210 (N_16210,N_15965,N_15964);
nor U16211 (N_16211,N_15972,N_16081);
nor U16212 (N_16212,N_15986,N_16021);
and U16213 (N_16213,N_15974,N_16135);
and U16214 (N_16214,N_16092,N_15923);
nand U16215 (N_16215,N_15928,N_16090);
nand U16216 (N_16216,N_15940,N_15919);
nand U16217 (N_16217,N_16019,N_16067);
or U16218 (N_16218,N_16143,N_16093);
nor U16219 (N_16219,N_16183,N_15934);
nor U16220 (N_16220,N_16002,N_16140);
or U16221 (N_16221,N_15996,N_15920);
nand U16222 (N_16222,N_15922,N_16077);
nand U16223 (N_16223,N_16116,N_16184);
nand U16224 (N_16224,N_16034,N_16165);
nand U16225 (N_16225,N_15951,N_15936);
or U16226 (N_16226,N_16195,N_16099);
or U16227 (N_16227,N_16174,N_16188);
or U16228 (N_16228,N_16009,N_16051);
xnor U16229 (N_16229,N_16000,N_15977);
xnor U16230 (N_16230,N_16071,N_16098);
xnor U16231 (N_16231,N_16138,N_16127);
xnor U16232 (N_16232,N_15967,N_16031);
xor U16233 (N_16233,N_16193,N_16029);
and U16234 (N_16234,N_15988,N_16028);
or U16235 (N_16235,N_15924,N_16055);
nor U16236 (N_16236,N_16069,N_16007);
and U16237 (N_16237,N_16157,N_15911);
nand U16238 (N_16238,N_15959,N_15960);
xnor U16239 (N_16239,N_16131,N_16154);
or U16240 (N_16240,N_16094,N_15909);
xor U16241 (N_16241,N_16146,N_16148);
nand U16242 (N_16242,N_16163,N_16089);
xnor U16243 (N_16243,N_16198,N_16141);
and U16244 (N_16244,N_16169,N_16044);
or U16245 (N_16245,N_16107,N_16024);
or U16246 (N_16246,N_16168,N_16086);
nor U16247 (N_16247,N_16022,N_16177);
nor U16248 (N_16248,N_16102,N_16113);
nor U16249 (N_16249,N_16061,N_15918);
nand U16250 (N_16250,N_16197,N_16073);
or U16251 (N_16251,N_16014,N_15927);
or U16252 (N_16252,N_15937,N_15952);
or U16253 (N_16253,N_16003,N_16057);
or U16254 (N_16254,N_16144,N_16050);
nand U16255 (N_16255,N_16039,N_16110);
nor U16256 (N_16256,N_16015,N_16156);
xor U16257 (N_16257,N_15999,N_16145);
and U16258 (N_16258,N_15968,N_16192);
or U16259 (N_16259,N_16152,N_15938);
or U16260 (N_16260,N_15966,N_15998);
nor U16261 (N_16261,N_16104,N_15948);
nand U16262 (N_16262,N_15981,N_16016);
and U16263 (N_16263,N_16196,N_16052);
or U16264 (N_16264,N_16046,N_16078);
or U16265 (N_16265,N_16121,N_16134);
or U16266 (N_16266,N_15935,N_16109);
and U16267 (N_16267,N_16056,N_16179);
xor U16268 (N_16268,N_16065,N_16012);
nand U16269 (N_16269,N_15942,N_15910);
or U16270 (N_16270,N_15921,N_16185);
nor U16271 (N_16271,N_15903,N_15997);
nand U16272 (N_16272,N_15958,N_16175);
nand U16273 (N_16273,N_16149,N_15932);
and U16274 (N_16274,N_16153,N_16128);
nand U16275 (N_16275,N_15929,N_16137);
and U16276 (N_16276,N_15914,N_16059);
and U16277 (N_16277,N_16041,N_15901);
xor U16278 (N_16278,N_15979,N_16032);
nor U16279 (N_16279,N_16150,N_15900);
and U16280 (N_16280,N_16043,N_15944);
nand U16281 (N_16281,N_16033,N_15905);
or U16282 (N_16282,N_15915,N_16049);
and U16283 (N_16283,N_16063,N_15945);
nor U16284 (N_16284,N_16124,N_16114);
nor U16285 (N_16285,N_16182,N_16194);
or U16286 (N_16286,N_15926,N_16117);
xor U16287 (N_16287,N_15943,N_16160);
xor U16288 (N_16288,N_15939,N_16047);
xor U16289 (N_16289,N_16125,N_16027);
nor U16290 (N_16290,N_16088,N_16167);
nor U16291 (N_16291,N_16187,N_15949);
xor U16292 (N_16292,N_16023,N_16074);
nor U16293 (N_16293,N_15976,N_16008);
or U16294 (N_16294,N_16147,N_16142);
nand U16295 (N_16295,N_16136,N_16045);
xor U16296 (N_16296,N_16101,N_15941);
nor U16297 (N_16297,N_16079,N_16005);
xnor U16298 (N_16298,N_16018,N_16026);
nor U16299 (N_16299,N_16006,N_16126);
or U16300 (N_16300,N_15995,N_16112);
nor U16301 (N_16301,N_15956,N_16190);
and U16302 (N_16302,N_15947,N_16158);
nand U16303 (N_16303,N_15990,N_16053);
nor U16304 (N_16304,N_15933,N_16181);
and U16305 (N_16305,N_16035,N_16097);
or U16306 (N_16306,N_15930,N_16155);
xnor U16307 (N_16307,N_16087,N_15970);
nand U16308 (N_16308,N_16020,N_15912);
xor U16309 (N_16309,N_15992,N_16001);
xnor U16310 (N_16310,N_16106,N_16115);
and U16311 (N_16311,N_16199,N_16083);
xor U16312 (N_16312,N_16004,N_15954);
xnor U16313 (N_16313,N_16178,N_16130);
or U16314 (N_16314,N_16017,N_16189);
or U16315 (N_16315,N_16066,N_16054);
nor U16316 (N_16316,N_16132,N_16038);
or U16317 (N_16317,N_16119,N_16037);
or U16318 (N_16318,N_15980,N_16176);
or U16319 (N_16319,N_16191,N_16036);
and U16320 (N_16320,N_16010,N_16111);
nand U16321 (N_16321,N_16133,N_15987);
nand U16322 (N_16322,N_15983,N_16085);
or U16323 (N_16323,N_16129,N_15957);
xnor U16324 (N_16324,N_16096,N_16105);
nand U16325 (N_16325,N_15908,N_16151);
or U16326 (N_16326,N_16173,N_16060);
nor U16327 (N_16327,N_16171,N_15913);
and U16328 (N_16328,N_15953,N_16072);
nor U16329 (N_16329,N_16166,N_16042);
nand U16330 (N_16330,N_16011,N_15982);
nor U16331 (N_16331,N_15902,N_16076);
xnor U16332 (N_16332,N_15925,N_16025);
and U16333 (N_16333,N_15969,N_16186);
nor U16334 (N_16334,N_15946,N_16084);
nor U16335 (N_16335,N_16120,N_16161);
nor U16336 (N_16336,N_15978,N_15994);
nor U16337 (N_16337,N_16122,N_15991);
and U16338 (N_16338,N_16091,N_16064);
nor U16339 (N_16339,N_16162,N_15917);
nand U16340 (N_16340,N_15984,N_16139);
or U16341 (N_16341,N_15907,N_15971);
or U16342 (N_16342,N_16080,N_15989);
or U16343 (N_16343,N_16103,N_15975);
and U16344 (N_16344,N_16095,N_15962);
and U16345 (N_16345,N_16170,N_16108);
nor U16346 (N_16346,N_15955,N_16159);
xor U16347 (N_16347,N_16172,N_16123);
nor U16348 (N_16348,N_16075,N_15973);
or U16349 (N_16349,N_16118,N_16100);
nand U16350 (N_16350,N_15907,N_16193);
or U16351 (N_16351,N_15998,N_16025);
or U16352 (N_16352,N_15986,N_16146);
nand U16353 (N_16353,N_16199,N_16116);
or U16354 (N_16354,N_15912,N_16171);
and U16355 (N_16355,N_15963,N_16102);
nand U16356 (N_16356,N_16174,N_16076);
xnor U16357 (N_16357,N_16038,N_16082);
xnor U16358 (N_16358,N_16036,N_16108);
xnor U16359 (N_16359,N_15970,N_16096);
nand U16360 (N_16360,N_16149,N_15960);
and U16361 (N_16361,N_15912,N_15979);
and U16362 (N_16362,N_16038,N_15923);
and U16363 (N_16363,N_16087,N_16114);
xnor U16364 (N_16364,N_16000,N_16102);
xor U16365 (N_16365,N_16006,N_16196);
or U16366 (N_16366,N_15990,N_15908);
and U16367 (N_16367,N_16125,N_15940);
or U16368 (N_16368,N_16120,N_16128);
nand U16369 (N_16369,N_16130,N_16022);
or U16370 (N_16370,N_15928,N_16157);
nand U16371 (N_16371,N_16079,N_15947);
nor U16372 (N_16372,N_15930,N_16149);
or U16373 (N_16373,N_16151,N_16074);
and U16374 (N_16374,N_16108,N_15912);
nand U16375 (N_16375,N_16066,N_15939);
nand U16376 (N_16376,N_16065,N_15950);
nor U16377 (N_16377,N_16133,N_16124);
or U16378 (N_16378,N_16095,N_15935);
nor U16379 (N_16379,N_15931,N_16104);
or U16380 (N_16380,N_15960,N_16105);
or U16381 (N_16381,N_16074,N_16125);
xor U16382 (N_16382,N_16162,N_16184);
nand U16383 (N_16383,N_16012,N_16024);
nor U16384 (N_16384,N_15952,N_15939);
xor U16385 (N_16385,N_16058,N_15905);
xnor U16386 (N_16386,N_16143,N_15998);
or U16387 (N_16387,N_16148,N_16170);
xnor U16388 (N_16388,N_16131,N_16091);
nor U16389 (N_16389,N_15918,N_16152);
nand U16390 (N_16390,N_16001,N_16019);
nor U16391 (N_16391,N_16132,N_16131);
nor U16392 (N_16392,N_15902,N_15958);
and U16393 (N_16393,N_15970,N_16101);
and U16394 (N_16394,N_16012,N_16194);
nand U16395 (N_16395,N_16089,N_15992);
xnor U16396 (N_16396,N_16029,N_15941);
xor U16397 (N_16397,N_16012,N_16040);
xnor U16398 (N_16398,N_15951,N_15937);
nand U16399 (N_16399,N_16128,N_16064);
nand U16400 (N_16400,N_16057,N_16156);
or U16401 (N_16401,N_15940,N_16042);
and U16402 (N_16402,N_16099,N_16007);
xor U16403 (N_16403,N_15929,N_16195);
or U16404 (N_16404,N_16152,N_16077);
or U16405 (N_16405,N_15962,N_15938);
xnor U16406 (N_16406,N_16108,N_15935);
nand U16407 (N_16407,N_16180,N_16062);
nor U16408 (N_16408,N_15914,N_16021);
nor U16409 (N_16409,N_16068,N_15956);
nand U16410 (N_16410,N_16137,N_16057);
nor U16411 (N_16411,N_15983,N_16052);
nor U16412 (N_16412,N_15982,N_15977);
and U16413 (N_16413,N_16144,N_16169);
nand U16414 (N_16414,N_16042,N_15982);
xor U16415 (N_16415,N_16105,N_15950);
xor U16416 (N_16416,N_16089,N_16173);
nand U16417 (N_16417,N_16184,N_16159);
xnor U16418 (N_16418,N_16061,N_15959);
nand U16419 (N_16419,N_16177,N_15953);
and U16420 (N_16420,N_16040,N_16015);
and U16421 (N_16421,N_16010,N_16004);
and U16422 (N_16422,N_16064,N_16152);
nand U16423 (N_16423,N_16190,N_16053);
and U16424 (N_16424,N_16185,N_15968);
and U16425 (N_16425,N_15917,N_15998);
nand U16426 (N_16426,N_15941,N_15928);
xnor U16427 (N_16427,N_16176,N_16006);
nor U16428 (N_16428,N_16031,N_16110);
nor U16429 (N_16429,N_16145,N_15974);
and U16430 (N_16430,N_16135,N_15988);
xor U16431 (N_16431,N_15936,N_16153);
and U16432 (N_16432,N_16009,N_16124);
nor U16433 (N_16433,N_16061,N_16173);
nand U16434 (N_16434,N_15981,N_16119);
and U16435 (N_16435,N_16181,N_16074);
or U16436 (N_16436,N_15924,N_16028);
nor U16437 (N_16437,N_16088,N_16115);
nand U16438 (N_16438,N_15946,N_16012);
and U16439 (N_16439,N_16105,N_16133);
and U16440 (N_16440,N_15943,N_16116);
nand U16441 (N_16441,N_16010,N_16052);
or U16442 (N_16442,N_16016,N_16040);
or U16443 (N_16443,N_15966,N_16013);
nor U16444 (N_16444,N_16112,N_16150);
and U16445 (N_16445,N_16090,N_15923);
nand U16446 (N_16446,N_15983,N_16082);
xnor U16447 (N_16447,N_16115,N_15945);
or U16448 (N_16448,N_15967,N_16066);
and U16449 (N_16449,N_15944,N_16164);
xor U16450 (N_16450,N_16179,N_15976);
nand U16451 (N_16451,N_15949,N_15937);
or U16452 (N_16452,N_16118,N_16132);
nand U16453 (N_16453,N_16130,N_16054);
nor U16454 (N_16454,N_16153,N_16164);
and U16455 (N_16455,N_15954,N_16116);
nand U16456 (N_16456,N_15980,N_16131);
nand U16457 (N_16457,N_16036,N_16092);
xnor U16458 (N_16458,N_15959,N_16158);
nand U16459 (N_16459,N_16152,N_15926);
and U16460 (N_16460,N_15965,N_16115);
and U16461 (N_16461,N_15971,N_15967);
or U16462 (N_16462,N_16131,N_15959);
nand U16463 (N_16463,N_16088,N_16170);
xor U16464 (N_16464,N_16197,N_16035);
xor U16465 (N_16465,N_16123,N_16002);
nand U16466 (N_16466,N_16027,N_15911);
nor U16467 (N_16467,N_16095,N_16103);
and U16468 (N_16468,N_16067,N_16123);
and U16469 (N_16469,N_15960,N_15953);
and U16470 (N_16470,N_16029,N_16187);
nor U16471 (N_16471,N_15901,N_16175);
xor U16472 (N_16472,N_15949,N_15992);
xnor U16473 (N_16473,N_16070,N_16147);
xor U16474 (N_16474,N_16038,N_16069);
xnor U16475 (N_16475,N_15943,N_15919);
nand U16476 (N_16476,N_16092,N_16131);
nor U16477 (N_16477,N_15981,N_15961);
or U16478 (N_16478,N_16060,N_16180);
nor U16479 (N_16479,N_16140,N_16113);
and U16480 (N_16480,N_15980,N_15913);
or U16481 (N_16481,N_16143,N_15977);
nand U16482 (N_16482,N_16059,N_16132);
nor U16483 (N_16483,N_16051,N_16028);
and U16484 (N_16484,N_15957,N_16102);
or U16485 (N_16485,N_15979,N_15945);
xor U16486 (N_16486,N_15934,N_15920);
nor U16487 (N_16487,N_16062,N_16024);
nand U16488 (N_16488,N_16130,N_16080);
nand U16489 (N_16489,N_16096,N_16178);
nor U16490 (N_16490,N_16057,N_15951);
or U16491 (N_16491,N_15965,N_15980);
nand U16492 (N_16492,N_15938,N_16129);
or U16493 (N_16493,N_16101,N_15978);
and U16494 (N_16494,N_16099,N_16179);
and U16495 (N_16495,N_15989,N_15970);
nor U16496 (N_16496,N_15952,N_15973);
nor U16497 (N_16497,N_16171,N_16051);
nor U16498 (N_16498,N_16148,N_16118);
xor U16499 (N_16499,N_16151,N_15959);
xor U16500 (N_16500,N_16209,N_16395);
nor U16501 (N_16501,N_16378,N_16431);
xor U16502 (N_16502,N_16414,N_16430);
and U16503 (N_16503,N_16381,N_16478);
nand U16504 (N_16504,N_16264,N_16481);
nor U16505 (N_16505,N_16295,N_16296);
xor U16506 (N_16506,N_16224,N_16260);
nor U16507 (N_16507,N_16306,N_16238);
or U16508 (N_16508,N_16272,N_16343);
nand U16509 (N_16509,N_16396,N_16281);
or U16510 (N_16510,N_16356,N_16248);
and U16511 (N_16511,N_16461,N_16347);
or U16512 (N_16512,N_16266,N_16398);
and U16513 (N_16513,N_16445,N_16307);
and U16514 (N_16514,N_16473,N_16474);
and U16515 (N_16515,N_16397,N_16417);
or U16516 (N_16516,N_16375,N_16348);
nor U16517 (N_16517,N_16488,N_16441);
nor U16518 (N_16518,N_16489,N_16285);
xnor U16519 (N_16519,N_16210,N_16391);
and U16520 (N_16520,N_16207,N_16354);
and U16521 (N_16521,N_16280,N_16440);
nor U16522 (N_16522,N_16475,N_16349);
nor U16523 (N_16523,N_16448,N_16233);
nor U16524 (N_16524,N_16476,N_16384);
xnor U16525 (N_16525,N_16402,N_16371);
xnor U16526 (N_16526,N_16342,N_16230);
xnor U16527 (N_16527,N_16428,N_16340);
or U16528 (N_16528,N_16362,N_16442);
nor U16529 (N_16529,N_16450,N_16420);
and U16530 (N_16530,N_16232,N_16373);
nand U16531 (N_16531,N_16487,N_16482);
and U16532 (N_16532,N_16419,N_16495);
or U16533 (N_16533,N_16304,N_16490);
and U16534 (N_16534,N_16245,N_16225);
nand U16535 (N_16535,N_16261,N_16374);
or U16536 (N_16536,N_16492,N_16409);
and U16537 (N_16537,N_16303,N_16425);
nand U16538 (N_16538,N_16453,N_16426);
nand U16539 (N_16539,N_16421,N_16333);
and U16540 (N_16540,N_16467,N_16389);
or U16541 (N_16541,N_16439,N_16462);
or U16542 (N_16542,N_16383,N_16336);
and U16543 (N_16543,N_16360,N_16289);
xnor U16544 (N_16544,N_16221,N_16290);
and U16545 (N_16545,N_16202,N_16454);
or U16546 (N_16546,N_16324,N_16410);
or U16547 (N_16547,N_16294,N_16205);
or U16548 (N_16548,N_16213,N_16345);
and U16549 (N_16549,N_16480,N_16404);
xnor U16550 (N_16550,N_16255,N_16339);
or U16551 (N_16551,N_16317,N_16386);
and U16552 (N_16552,N_16271,N_16466);
or U16553 (N_16553,N_16321,N_16382);
or U16554 (N_16554,N_16403,N_16226);
or U16555 (N_16555,N_16385,N_16468);
nor U16556 (N_16556,N_16412,N_16313);
nand U16557 (N_16557,N_16352,N_16499);
nor U16558 (N_16558,N_16228,N_16203);
or U16559 (N_16559,N_16325,N_16400);
or U16560 (N_16560,N_16262,N_16493);
or U16561 (N_16561,N_16483,N_16310);
xnor U16562 (N_16562,N_16265,N_16498);
and U16563 (N_16563,N_16355,N_16223);
xnor U16564 (N_16564,N_16364,N_16334);
xnor U16565 (N_16565,N_16405,N_16460);
nand U16566 (N_16566,N_16332,N_16211);
and U16567 (N_16567,N_16366,N_16456);
and U16568 (N_16568,N_16387,N_16444);
and U16569 (N_16569,N_16267,N_16240);
xor U16570 (N_16570,N_16367,N_16299);
nor U16571 (N_16571,N_16350,N_16413);
or U16572 (N_16572,N_16415,N_16286);
xnor U16573 (N_16573,N_16287,N_16312);
and U16574 (N_16574,N_16243,N_16305);
and U16575 (N_16575,N_16315,N_16335);
xor U16576 (N_16576,N_16455,N_16250);
nor U16577 (N_16577,N_16311,N_16215);
nor U16578 (N_16578,N_16427,N_16254);
xnor U16579 (N_16579,N_16263,N_16330);
and U16580 (N_16580,N_16446,N_16268);
nand U16581 (N_16581,N_16491,N_16463);
nor U16582 (N_16582,N_16256,N_16407);
or U16583 (N_16583,N_16392,N_16201);
or U16584 (N_16584,N_16437,N_16472);
and U16585 (N_16585,N_16244,N_16322);
nand U16586 (N_16586,N_16316,N_16459);
xor U16587 (N_16587,N_16283,N_16406);
xor U16588 (N_16588,N_16249,N_16436);
and U16589 (N_16589,N_16270,N_16423);
or U16590 (N_16590,N_16331,N_16432);
nand U16591 (N_16591,N_16220,N_16300);
and U16592 (N_16592,N_16429,N_16219);
and U16593 (N_16593,N_16358,N_16273);
or U16594 (N_16594,N_16229,N_16451);
nand U16595 (N_16595,N_16284,N_16408);
nand U16596 (N_16596,N_16206,N_16253);
nor U16597 (N_16597,N_16320,N_16323);
nand U16598 (N_16598,N_16216,N_16231);
xor U16599 (N_16599,N_16298,N_16443);
and U16600 (N_16600,N_16302,N_16435);
or U16601 (N_16601,N_16314,N_16394);
nand U16602 (N_16602,N_16239,N_16319);
nor U16603 (N_16603,N_16236,N_16496);
nand U16604 (N_16604,N_16247,N_16365);
nand U16605 (N_16605,N_16372,N_16297);
or U16606 (N_16606,N_16237,N_16208);
xnor U16607 (N_16607,N_16361,N_16337);
nand U16608 (N_16608,N_16388,N_16329);
or U16609 (N_16609,N_16449,N_16357);
or U16610 (N_16610,N_16494,N_16416);
xnor U16611 (N_16611,N_16309,N_16470);
nor U16612 (N_16612,N_16368,N_16212);
or U16613 (N_16613,N_16327,N_16269);
and U16614 (N_16614,N_16486,N_16291);
xnor U16615 (N_16615,N_16204,N_16379);
or U16616 (N_16616,N_16464,N_16438);
nand U16617 (N_16617,N_16293,N_16344);
xnor U16618 (N_16618,N_16222,N_16452);
nand U16619 (N_16619,N_16258,N_16257);
or U16620 (N_16620,N_16369,N_16252);
and U16621 (N_16621,N_16422,N_16217);
and U16622 (N_16622,N_16471,N_16235);
nor U16623 (N_16623,N_16308,N_16376);
nand U16624 (N_16624,N_16484,N_16301);
and U16625 (N_16625,N_16282,N_16259);
or U16626 (N_16626,N_16363,N_16278);
and U16627 (N_16627,N_16465,N_16214);
xnor U16628 (N_16628,N_16401,N_16377);
nand U16629 (N_16629,N_16288,N_16424);
and U16630 (N_16630,N_16393,N_16251);
nand U16631 (N_16631,N_16218,N_16276);
nor U16632 (N_16632,N_16275,N_16457);
and U16633 (N_16633,N_16485,N_16200);
nand U16634 (N_16634,N_16328,N_16338);
or U16635 (N_16635,N_16434,N_16234);
or U16636 (N_16636,N_16353,N_16326);
nand U16637 (N_16637,N_16241,N_16370);
xor U16638 (N_16638,N_16341,N_16246);
nand U16639 (N_16639,N_16447,N_16242);
xor U16640 (N_16640,N_16418,N_16477);
xor U16641 (N_16641,N_16274,N_16351);
nor U16642 (N_16642,N_16380,N_16346);
and U16643 (N_16643,N_16497,N_16411);
xnor U16644 (N_16644,N_16359,N_16479);
xor U16645 (N_16645,N_16279,N_16399);
and U16646 (N_16646,N_16227,N_16318);
or U16647 (N_16647,N_16292,N_16469);
xnor U16648 (N_16648,N_16390,N_16277);
or U16649 (N_16649,N_16433,N_16458);
or U16650 (N_16650,N_16386,N_16451);
or U16651 (N_16651,N_16475,N_16275);
and U16652 (N_16652,N_16412,N_16217);
and U16653 (N_16653,N_16250,N_16333);
xnor U16654 (N_16654,N_16336,N_16211);
and U16655 (N_16655,N_16256,N_16471);
nand U16656 (N_16656,N_16460,N_16328);
xor U16657 (N_16657,N_16230,N_16265);
xnor U16658 (N_16658,N_16430,N_16315);
and U16659 (N_16659,N_16351,N_16327);
and U16660 (N_16660,N_16234,N_16222);
and U16661 (N_16661,N_16458,N_16209);
and U16662 (N_16662,N_16408,N_16438);
xnor U16663 (N_16663,N_16216,N_16488);
and U16664 (N_16664,N_16398,N_16239);
or U16665 (N_16665,N_16245,N_16323);
nor U16666 (N_16666,N_16395,N_16444);
nand U16667 (N_16667,N_16217,N_16288);
nand U16668 (N_16668,N_16349,N_16414);
xor U16669 (N_16669,N_16421,N_16331);
nor U16670 (N_16670,N_16285,N_16303);
xnor U16671 (N_16671,N_16396,N_16373);
nand U16672 (N_16672,N_16263,N_16358);
nor U16673 (N_16673,N_16363,N_16379);
nand U16674 (N_16674,N_16326,N_16209);
and U16675 (N_16675,N_16225,N_16288);
xnor U16676 (N_16676,N_16273,N_16326);
or U16677 (N_16677,N_16228,N_16222);
and U16678 (N_16678,N_16331,N_16334);
nand U16679 (N_16679,N_16398,N_16489);
xnor U16680 (N_16680,N_16470,N_16422);
xor U16681 (N_16681,N_16363,N_16366);
and U16682 (N_16682,N_16226,N_16313);
xnor U16683 (N_16683,N_16283,N_16290);
and U16684 (N_16684,N_16466,N_16308);
and U16685 (N_16685,N_16233,N_16397);
and U16686 (N_16686,N_16486,N_16273);
nor U16687 (N_16687,N_16331,N_16441);
and U16688 (N_16688,N_16426,N_16347);
nand U16689 (N_16689,N_16367,N_16289);
and U16690 (N_16690,N_16427,N_16355);
nand U16691 (N_16691,N_16237,N_16357);
xor U16692 (N_16692,N_16290,N_16350);
xnor U16693 (N_16693,N_16432,N_16208);
or U16694 (N_16694,N_16231,N_16256);
nor U16695 (N_16695,N_16427,N_16231);
or U16696 (N_16696,N_16223,N_16401);
or U16697 (N_16697,N_16205,N_16478);
or U16698 (N_16698,N_16470,N_16243);
and U16699 (N_16699,N_16314,N_16494);
nand U16700 (N_16700,N_16214,N_16434);
and U16701 (N_16701,N_16439,N_16492);
nand U16702 (N_16702,N_16443,N_16263);
and U16703 (N_16703,N_16458,N_16297);
or U16704 (N_16704,N_16264,N_16338);
xor U16705 (N_16705,N_16321,N_16285);
xnor U16706 (N_16706,N_16407,N_16238);
or U16707 (N_16707,N_16395,N_16305);
and U16708 (N_16708,N_16442,N_16443);
or U16709 (N_16709,N_16459,N_16490);
or U16710 (N_16710,N_16213,N_16434);
xor U16711 (N_16711,N_16247,N_16384);
and U16712 (N_16712,N_16437,N_16346);
and U16713 (N_16713,N_16475,N_16251);
nand U16714 (N_16714,N_16363,N_16362);
xnor U16715 (N_16715,N_16387,N_16364);
and U16716 (N_16716,N_16489,N_16327);
xor U16717 (N_16717,N_16390,N_16250);
and U16718 (N_16718,N_16378,N_16321);
xor U16719 (N_16719,N_16277,N_16262);
nand U16720 (N_16720,N_16401,N_16265);
xnor U16721 (N_16721,N_16395,N_16336);
and U16722 (N_16722,N_16378,N_16390);
nand U16723 (N_16723,N_16488,N_16386);
xnor U16724 (N_16724,N_16315,N_16255);
xor U16725 (N_16725,N_16212,N_16308);
or U16726 (N_16726,N_16288,N_16406);
nor U16727 (N_16727,N_16318,N_16365);
and U16728 (N_16728,N_16268,N_16356);
nand U16729 (N_16729,N_16309,N_16488);
xnor U16730 (N_16730,N_16455,N_16232);
nor U16731 (N_16731,N_16299,N_16262);
and U16732 (N_16732,N_16309,N_16466);
nand U16733 (N_16733,N_16353,N_16336);
or U16734 (N_16734,N_16307,N_16327);
and U16735 (N_16735,N_16350,N_16384);
nor U16736 (N_16736,N_16413,N_16408);
or U16737 (N_16737,N_16405,N_16427);
and U16738 (N_16738,N_16321,N_16412);
and U16739 (N_16739,N_16499,N_16403);
nor U16740 (N_16740,N_16322,N_16342);
nor U16741 (N_16741,N_16431,N_16292);
nand U16742 (N_16742,N_16238,N_16427);
and U16743 (N_16743,N_16494,N_16428);
nand U16744 (N_16744,N_16334,N_16360);
nand U16745 (N_16745,N_16222,N_16218);
or U16746 (N_16746,N_16284,N_16371);
xor U16747 (N_16747,N_16451,N_16417);
and U16748 (N_16748,N_16418,N_16347);
nand U16749 (N_16749,N_16364,N_16369);
nor U16750 (N_16750,N_16431,N_16238);
xor U16751 (N_16751,N_16460,N_16448);
or U16752 (N_16752,N_16310,N_16202);
xor U16753 (N_16753,N_16476,N_16386);
and U16754 (N_16754,N_16273,N_16388);
or U16755 (N_16755,N_16238,N_16384);
nor U16756 (N_16756,N_16325,N_16364);
nor U16757 (N_16757,N_16249,N_16321);
and U16758 (N_16758,N_16305,N_16211);
or U16759 (N_16759,N_16430,N_16244);
and U16760 (N_16760,N_16293,N_16361);
nor U16761 (N_16761,N_16260,N_16342);
and U16762 (N_16762,N_16487,N_16204);
nor U16763 (N_16763,N_16453,N_16384);
or U16764 (N_16764,N_16415,N_16211);
nand U16765 (N_16765,N_16281,N_16335);
xor U16766 (N_16766,N_16334,N_16337);
or U16767 (N_16767,N_16482,N_16228);
or U16768 (N_16768,N_16405,N_16458);
xor U16769 (N_16769,N_16305,N_16365);
or U16770 (N_16770,N_16295,N_16476);
nor U16771 (N_16771,N_16286,N_16261);
nand U16772 (N_16772,N_16213,N_16245);
and U16773 (N_16773,N_16248,N_16330);
or U16774 (N_16774,N_16229,N_16260);
and U16775 (N_16775,N_16322,N_16283);
nand U16776 (N_16776,N_16381,N_16453);
xor U16777 (N_16777,N_16350,N_16414);
xnor U16778 (N_16778,N_16328,N_16388);
and U16779 (N_16779,N_16450,N_16226);
and U16780 (N_16780,N_16206,N_16333);
and U16781 (N_16781,N_16458,N_16290);
and U16782 (N_16782,N_16481,N_16210);
or U16783 (N_16783,N_16283,N_16255);
nand U16784 (N_16784,N_16325,N_16482);
nand U16785 (N_16785,N_16361,N_16436);
xnor U16786 (N_16786,N_16300,N_16226);
or U16787 (N_16787,N_16324,N_16444);
and U16788 (N_16788,N_16317,N_16303);
xnor U16789 (N_16789,N_16264,N_16316);
nand U16790 (N_16790,N_16224,N_16496);
or U16791 (N_16791,N_16293,N_16357);
and U16792 (N_16792,N_16264,N_16324);
or U16793 (N_16793,N_16447,N_16203);
xor U16794 (N_16794,N_16386,N_16494);
nand U16795 (N_16795,N_16226,N_16302);
nand U16796 (N_16796,N_16236,N_16230);
or U16797 (N_16797,N_16473,N_16412);
and U16798 (N_16798,N_16386,N_16431);
nand U16799 (N_16799,N_16283,N_16461);
nand U16800 (N_16800,N_16511,N_16577);
nor U16801 (N_16801,N_16738,N_16692);
or U16802 (N_16802,N_16745,N_16565);
or U16803 (N_16803,N_16530,N_16652);
or U16804 (N_16804,N_16515,N_16784);
and U16805 (N_16805,N_16676,N_16750);
nand U16806 (N_16806,N_16659,N_16520);
nand U16807 (N_16807,N_16727,N_16535);
or U16808 (N_16808,N_16672,N_16605);
or U16809 (N_16809,N_16749,N_16572);
and U16810 (N_16810,N_16697,N_16613);
nand U16811 (N_16811,N_16512,N_16654);
or U16812 (N_16812,N_16788,N_16688);
nor U16813 (N_16813,N_16773,N_16606);
nor U16814 (N_16814,N_16502,N_16768);
nand U16815 (N_16815,N_16614,N_16592);
or U16816 (N_16816,N_16508,N_16513);
nor U16817 (N_16817,N_16782,N_16668);
nor U16818 (N_16818,N_16709,N_16564);
xor U16819 (N_16819,N_16763,N_16776);
xnor U16820 (N_16820,N_16761,N_16716);
nor U16821 (N_16821,N_16537,N_16648);
nor U16822 (N_16822,N_16787,N_16724);
nor U16823 (N_16823,N_16552,N_16667);
or U16824 (N_16824,N_16578,N_16562);
nor U16825 (N_16825,N_16705,N_16673);
xor U16826 (N_16826,N_16755,N_16781);
nor U16827 (N_16827,N_16793,N_16785);
nand U16828 (N_16828,N_16585,N_16597);
or U16829 (N_16829,N_16608,N_16767);
or U16830 (N_16830,N_16504,N_16573);
nand U16831 (N_16831,N_16700,N_16607);
or U16832 (N_16832,N_16567,N_16798);
nand U16833 (N_16833,N_16647,N_16725);
nand U16834 (N_16834,N_16551,N_16757);
nor U16835 (N_16835,N_16505,N_16501);
xnor U16836 (N_16836,N_16538,N_16542);
nor U16837 (N_16837,N_16590,N_16526);
xnor U16838 (N_16838,N_16758,N_16766);
nor U16839 (N_16839,N_16547,N_16517);
and U16840 (N_16840,N_16625,N_16529);
and U16841 (N_16841,N_16594,N_16645);
and U16842 (N_16842,N_16778,N_16588);
nand U16843 (N_16843,N_16717,N_16674);
or U16844 (N_16844,N_16695,N_16579);
nor U16845 (N_16845,N_16683,N_16701);
or U16846 (N_16846,N_16704,N_16698);
nor U16847 (N_16847,N_16633,N_16617);
xor U16848 (N_16848,N_16616,N_16739);
or U16849 (N_16849,N_16710,N_16558);
nand U16850 (N_16850,N_16561,N_16733);
xor U16851 (N_16851,N_16591,N_16675);
or U16852 (N_16852,N_16678,N_16549);
nand U16853 (N_16853,N_16621,N_16651);
and U16854 (N_16854,N_16533,N_16560);
xor U16855 (N_16855,N_16630,N_16677);
nor U16856 (N_16856,N_16660,N_16563);
nor U16857 (N_16857,N_16665,N_16792);
nand U16858 (N_16858,N_16619,N_16743);
xor U16859 (N_16859,N_16797,N_16687);
nor U16860 (N_16860,N_16521,N_16627);
xor U16861 (N_16861,N_16794,N_16569);
and U16862 (N_16862,N_16663,N_16615);
and U16863 (N_16863,N_16507,N_16694);
nor U16864 (N_16864,N_16711,N_16707);
or U16865 (N_16865,N_16731,N_16671);
nand U16866 (N_16866,N_16669,N_16602);
nand U16867 (N_16867,N_16748,N_16680);
nand U16868 (N_16868,N_16586,N_16769);
and U16869 (N_16869,N_16516,N_16601);
and U16870 (N_16870,N_16644,N_16679);
xnor U16871 (N_16871,N_16759,N_16772);
xnor U16872 (N_16872,N_16756,N_16500);
nor U16873 (N_16873,N_16544,N_16771);
and U16874 (N_16874,N_16628,N_16664);
or U16875 (N_16875,N_16640,N_16568);
and U16876 (N_16876,N_16791,N_16662);
xor U16877 (N_16877,N_16634,N_16531);
nand U16878 (N_16878,N_16523,N_16624);
xor U16879 (N_16879,N_16650,N_16553);
nand U16880 (N_16880,N_16612,N_16661);
xor U16881 (N_16881,N_16545,N_16596);
and U16882 (N_16882,N_16539,N_16574);
nor U16883 (N_16883,N_16638,N_16693);
xnor U16884 (N_16884,N_16783,N_16556);
nor U16885 (N_16885,N_16670,N_16587);
and U16886 (N_16886,N_16681,N_16635);
or U16887 (N_16887,N_16584,N_16656);
nor U16888 (N_16888,N_16580,N_16599);
and U16889 (N_16889,N_16744,N_16554);
and U16890 (N_16890,N_16751,N_16543);
nand U16891 (N_16891,N_16754,N_16631);
nor U16892 (N_16892,N_16746,N_16598);
or U16893 (N_16893,N_16593,N_16719);
nor U16894 (N_16894,N_16742,N_16546);
and U16895 (N_16895,N_16715,N_16777);
and U16896 (N_16896,N_16548,N_16510);
nor U16897 (N_16897,N_16703,N_16774);
nor U16898 (N_16898,N_16706,N_16509);
and U16899 (N_16899,N_16740,N_16583);
nor U16900 (N_16900,N_16770,N_16790);
xnor U16901 (N_16901,N_16714,N_16646);
or U16902 (N_16902,N_16559,N_16557);
or U16903 (N_16903,N_16532,N_16789);
xnor U16904 (N_16904,N_16604,N_16666);
xor U16905 (N_16905,N_16519,N_16637);
or U16906 (N_16906,N_16582,N_16775);
xnor U16907 (N_16907,N_16726,N_16595);
xor U16908 (N_16908,N_16689,N_16796);
xor U16909 (N_16909,N_16575,N_16686);
xnor U16910 (N_16910,N_16799,N_16641);
or U16911 (N_16911,N_16795,N_16609);
nor U16912 (N_16912,N_16603,N_16723);
nor U16913 (N_16913,N_16642,N_16722);
xor U16914 (N_16914,N_16540,N_16684);
nor U16915 (N_16915,N_16581,N_16699);
and U16916 (N_16916,N_16657,N_16721);
xor U16917 (N_16917,N_16620,N_16736);
or U16918 (N_16918,N_16622,N_16729);
and U16919 (N_16919,N_16753,N_16525);
or U16920 (N_16920,N_16655,N_16752);
or U16921 (N_16921,N_16524,N_16555);
nor U16922 (N_16922,N_16780,N_16610);
nand U16923 (N_16923,N_16629,N_16747);
and U16924 (N_16924,N_16718,N_16534);
and U16925 (N_16925,N_16636,N_16536);
or U16926 (N_16926,N_16626,N_16632);
xnor U16927 (N_16927,N_16611,N_16762);
xnor U16928 (N_16928,N_16765,N_16734);
or U16929 (N_16929,N_16720,N_16639);
or U16930 (N_16930,N_16702,N_16541);
nand U16931 (N_16931,N_16786,N_16589);
and U16932 (N_16932,N_16735,N_16732);
nand U16933 (N_16933,N_16760,N_16708);
xnor U16934 (N_16934,N_16730,N_16623);
xnor U16935 (N_16935,N_16653,N_16779);
or U16936 (N_16936,N_16737,N_16685);
and U16937 (N_16937,N_16571,N_16600);
nor U16938 (N_16938,N_16712,N_16682);
or U16939 (N_16939,N_16570,N_16649);
and U16940 (N_16940,N_16696,N_16713);
nor U16941 (N_16941,N_16764,N_16691);
nor U16942 (N_16942,N_16576,N_16728);
and U16943 (N_16943,N_16550,N_16658);
or U16944 (N_16944,N_16503,N_16522);
and U16945 (N_16945,N_16506,N_16690);
nand U16946 (N_16946,N_16528,N_16741);
or U16947 (N_16947,N_16527,N_16518);
nor U16948 (N_16948,N_16618,N_16643);
xor U16949 (N_16949,N_16514,N_16566);
xor U16950 (N_16950,N_16706,N_16563);
nor U16951 (N_16951,N_16782,N_16698);
xnor U16952 (N_16952,N_16758,N_16616);
or U16953 (N_16953,N_16661,N_16702);
or U16954 (N_16954,N_16677,N_16548);
and U16955 (N_16955,N_16611,N_16770);
and U16956 (N_16956,N_16794,N_16653);
nor U16957 (N_16957,N_16671,N_16516);
nor U16958 (N_16958,N_16725,N_16534);
xnor U16959 (N_16959,N_16664,N_16610);
or U16960 (N_16960,N_16715,N_16563);
nor U16961 (N_16961,N_16596,N_16795);
or U16962 (N_16962,N_16717,N_16516);
or U16963 (N_16963,N_16786,N_16590);
nor U16964 (N_16964,N_16543,N_16544);
nor U16965 (N_16965,N_16679,N_16783);
and U16966 (N_16966,N_16505,N_16509);
and U16967 (N_16967,N_16610,N_16734);
nor U16968 (N_16968,N_16600,N_16590);
nand U16969 (N_16969,N_16665,N_16662);
or U16970 (N_16970,N_16789,N_16620);
xnor U16971 (N_16971,N_16647,N_16542);
nand U16972 (N_16972,N_16769,N_16500);
xnor U16973 (N_16973,N_16733,N_16786);
xnor U16974 (N_16974,N_16545,N_16507);
or U16975 (N_16975,N_16735,N_16587);
and U16976 (N_16976,N_16561,N_16521);
or U16977 (N_16977,N_16665,N_16778);
or U16978 (N_16978,N_16520,N_16691);
nand U16979 (N_16979,N_16644,N_16704);
nor U16980 (N_16980,N_16556,N_16752);
or U16981 (N_16981,N_16732,N_16595);
xor U16982 (N_16982,N_16533,N_16708);
and U16983 (N_16983,N_16601,N_16662);
or U16984 (N_16984,N_16523,N_16630);
and U16985 (N_16985,N_16604,N_16520);
xnor U16986 (N_16986,N_16689,N_16570);
and U16987 (N_16987,N_16510,N_16505);
nor U16988 (N_16988,N_16541,N_16768);
xnor U16989 (N_16989,N_16750,N_16682);
nor U16990 (N_16990,N_16500,N_16623);
or U16991 (N_16991,N_16523,N_16568);
xnor U16992 (N_16992,N_16763,N_16770);
nor U16993 (N_16993,N_16530,N_16674);
nand U16994 (N_16994,N_16533,N_16597);
and U16995 (N_16995,N_16509,N_16751);
xor U16996 (N_16996,N_16642,N_16541);
nor U16997 (N_16997,N_16545,N_16745);
nor U16998 (N_16998,N_16596,N_16792);
xor U16999 (N_16999,N_16692,N_16752);
xor U17000 (N_17000,N_16707,N_16601);
or U17001 (N_17001,N_16630,N_16543);
nor U17002 (N_17002,N_16513,N_16751);
xor U17003 (N_17003,N_16602,N_16736);
and U17004 (N_17004,N_16572,N_16637);
and U17005 (N_17005,N_16649,N_16729);
xnor U17006 (N_17006,N_16520,N_16574);
xnor U17007 (N_17007,N_16720,N_16666);
and U17008 (N_17008,N_16715,N_16615);
nand U17009 (N_17009,N_16556,N_16659);
or U17010 (N_17010,N_16732,N_16593);
xor U17011 (N_17011,N_16700,N_16511);
or U17012 (N_17012,N_16506,N_16663);
xor U17013 (N_17013,N_16677,N_16770);
nand U17014 (N_17014,N_16536,N_16671);
nor U17015 (N_17015,N_16600,N_16734);
or U17016 (N_17016,N_16708,N_16699);
nand U17017 (N_17017,N_16701,N_16601);
xnor U17018 (N_17018,N_16742,N_16632);
nand U17019 (N_17019,N_16512,N_16521);
or U17020 (N_17020,N_16536,N_16777);
xnor U17021 (N_17021,N_16744,N_16682);
or U17022 (N_17022,N_16548,N_16633);
and U17023 (N_17023,N_16720,N_16616);
or U17024 (N_17024,N_16656,N_16655);
nand U17025 (N_17025,N_16716,N_16644);
and U17026 (N_17026,N_16731,N_16606);
nor U17027 (N_17027,N_16687,N_16695);
nand U17028 (N_17028,N_16664,N_16668);
and U17029 (N_17029,N_16532,N_16666);
nor U17030 (N_17030,N_16561,N_16639);
xor U17031 (N_17031,N_16662,N_16653);
and U17032 (N_17032,N_16633,N_16628);
nor U17033 (N_17033,N_16704,N_16747);
nor U17034 (N_17034,N_16623,N_16727);
xnor U17035 (N_17035,N_16535,N_16754);
or U17036 (N_17036,N_16755,N_16521);
and U17037 (N_17037,N_16521,N_16799);
nor U17038 (N_17038,N_16797,N_16618);
nand U17039 (N_17039,N_16595,N_16707);
or U17040 (N_17040,N_16504,N_16613);
nand U17041 (N_17041,N_16594,N_16775);
nor U17042 (N_17042,N_16528,N_16765);
or U17043 (N_17043,N_16718,N_16688);
and U17044 (N_17044,N_16756,N_16654);
nor U17045 (N_17045,N_16758,N_16514);
nor U17046 (N_17046,N_16586,N_16587);
or U17047 (N_17047,N_16729,N_16786);
nor U17048 (N_17048,N_16623,N_16699);
and U17049 (N_17049,N_16681,N_16732);
nand U17050 (N_17050,N_16639,N_16723);
and U17051 (N_17051,N_16640,N_16540);
xnor U17052 (N_17052,N_16643,N_16763);
and U17053 (N_17053,N_16660,N_16557);
and U17054 (N_17054,N_16694,N_16718);
or U17055 (N_17055,N_16525,N_16684);
nand U17056 (N_17056,N_16607,N_16621);
nand U17057 (N_17057,N_16570,N_16665);
nand U17058 (N_17058,N_16529,N_16512);
xor U17059 (N_17059,N_16727,N_16648);
or U17060 (N_17060,N_16778,N_16706);
nor U17061 (N_17061,N_16551,N_16786);
and U17062 (N_17062,N_16625,N_16570);
nor U17063 (N_17063,N_16704,N_16553);
or U17064 (N_17064,N_16511,N_16763);
nor U17065 (N_17065,N_16698,N_16785);
nor U17066 (N_17066,N_16687,N_16795);
nand U17067 (N_17067,N_16696,N_16503);
and U17068 (N_17068,N_16555,N_16578);
xor U17069 (N_17069,N_16722,N_16720);
nand U17070 (N_17070,N_16720,N_16575);
nor U17071 (N_17071,N_16799,N_16582);
nor U17072 (N_17072,N_16510,N_16735);
or U17073 (N_17073,N_16522,N_16733);
or U17074 (N_17074,N_16582,N_16796);
xor U17075 (N_17075,N_16547,N_16783);
nand U17076 (N_17076,N_16511,N_16792);
nand U17077 (N_17077,N_16769,N_16570);
or U17078 (N_17078,N_16695,N_16670);
nor U17079 (N_17079,N_16612,N_16698);
or U17080 (N_17080,N_16767,N_16662);
nand U17081 (N_17081,N_16782,N_16780);
and U17082 (N_17082,N_16525,N_16787);
nor U17083 (N_17083,N_16552,N_16651);
xnor U17084 (N_17084,N_16583,N_16527);
or U17085 (N_17085,N_16516,N_16697);
nor U17086 (N_17086,N_16765,N_16551);
xor U17087 (N_17087,N_16568,N_16540);
nor U17088 (N_17088,N_16569,N_16699);
or U17089 (N_17089,N_16799,N_16612);
and U17090 (N_17090,N_16788,N_16663);
or U17091 (N_17091,N_16638,N_16523);
nand U17092 (N_17092,N_16791,N_16735);
xnor U17093 (N_17093,N_16662,N_16711);
nand U17094 (N_17094,N_16542,N_16526);
nand U17095 (N_17095,N_16663,N_16524);
or U17096 (N_17096,N_16590,N_16537);
and U17097 (N_17097,N_16549,N_16700);
and U17098 (N_17098,N_16746,N_16711);
or U17099 (N_17099,N_16695,N_16692);
nand U17100 (N_17100,N_17031,N_16859);
nor U17101 (N_17101,N_16914,N_16985);
and U17102 (N_17102,N_16830,N_17019);
or U17103 (N_17103,N_17012,N_16996);
nor U17104 (N_17104,N_17003,N_17066);
nand U17105 (N_17105,N_17037,N_16942);
and U17106 (N_17106,N_16896,N_16915);
or U17107 (N_17107,N_16906,N_16894);
nor U17108 (N_17108,N_16892,N_16988);
nor U17109 (N_17109,N_17047,N_16964);
nor U17110 (N_17110,N_17073,N_16806);
xor U17111 (N_17111,N_16845,N_17077);
xor U17112 (N_17112,N_16812,N_17079);
xnor U17113 (N_17113,N_16975,N_16981);
nor U17114 (N_17114,N_16930,N_17083);
and U17115 (N_17115,N_17011,N_17049);
xor U17116 (N_17116,N_16840,N_16917);
or U17117 (N_17117,N_16874,N_16961);
and U17118 (N_17118,N_16873,N_17075);
nor U17119 (N_17119,N_17028,N_17080);
and U17120 (N_17120,N_16986,N_16870);
xnor U17121 (N_17121,N_16867,N_17045);
nand U17122 (N_17122,N_16932,N_16811);
and U17123 (N_17123,N_16955,N_17093);
nor U17124 (N_17124,N_16935,N_16834);
nor U17125 (N_17125,N_16853,N_17084);
nand U17126 (N_17126,N_17023,N_17053);
xor U17127 (N_17127,N_17004,N_17040);
or U17128 (N_17128,N_16803,N_17070);
xor U17129 (N_17129,N_16848,N_16990);
and U17130 (N_17130,N_17048,N_17016);
and U17131 (N_17131,N_16900,N_16881);
and U17132 (N_17132,N_16882,N_17069);
or U17133 (N_17133,N_16814,N_16861);
or U17134 (N_17134,N_16851,N_17082);
nand U17135 (N_17135,N_16864,N_17025);
or U17136 (N_17136,N_16916,N_16852);
nor U17137 (N_17137,N_16951,N_16836);
nor U17138 (N_17138,N_16862,N_16888);
nand U17139 (N_17139,N_16837,N_16832);
nand U17140 (N_17140,N_16855,N_16994);
or U17141 (N_17141,N_16946,N_16993);
xor U17142 (N_17142,N_17074,N_17052);
nand U17143 (N_17143,N_17026,N_16967);
and U17144 (N_17144,N_17068,N_17007);
nand U17145 (N_17145,N_16885,N_16801);
xnor U17146 (N_17146,N_16823,N_16866);
or U17147 (N_17147,N_17076,N_16802);
nand U17148 (N_17148,N_17089,N_16982);
nand U17149 (N_17149,N_17097,N_16819);
xor U17150 (N_17150,N_17081,N_16965);
or U17151 (N_17151,N_16856,N_16849);
or U17152 (N_17152,N_16841,N_16911);
nand U17153 (N_17153,N_16880,N_16983);
xnor U17154 (N_17154,N_16850,N_17056);
xnor U17155 (N_17155,N_16843,N_16865);
or U17156 (N_17156,N_17098,N_17071);
nand U17157 (N_17157,N_17027,N_16931);
nand U17158 (N_17158,N_16828,N_17014);
nor U17159 (N_17159,N_16947,N_17043);
nor U17160 (N_17160,N_17085,N_16991);
and U17161 (N_17161,N_16977,N_16875);
xnor U17162 (N_17162,N_16846,N_17030);
nand U17163 (N_17163,N_16813,N_16963);
nand U17164 (N_17164,N_16927,N_16992);
and U17165 (N_17165,N_16928,N_16948);
and U17166 (N_17166,N_16902,N_17021);
and U17167 (N_17167,N_16956,N_17042);
xor U17168 (N_17168,N_16926,N_17013);
or U17169 (N_17169,N_17091,N_17096);
xor U17170 (N_17170,N_16970,N_17024);
or U17171 (N_17171,N_17065,N_16937);
nor U17172 (N_17172,N_16943,N_16829);
and U17173 (N_17173,N_17002,N_16922);
and U17174 (N_17174,N_16824,N_17061);
nand U17175 (N_17175,N_16895,N_16839);
and U17176 (N_17176,N_16899,N_16872);
or U17177 (N_17177,N_17064,N_17046);
and U17178 (N_17178,N_16998,N_16997);
or U17179 (N_17179,N_16921,N_16938);
nor U17180 (N_17180,N_17005,N_17029);
and U17181 (N_17181,N_16987,N_16960);
nand U17182 (N_17182,N_16976,N_16858);
nand U17183 (N_17183,N_17055,N_16807);
nor U17184 (N_17184,N_16929,N_16810);
nor U17185 (N_17185,N_16959,N_16816);
nor U17186 (N_17186,N_16889,N_17009);
or U17187 (N_17187,N_16905,N_16989);
and U17188 (N_17188,N_16854,N_16950);
or U17189 (N_17189,N_16941,N_16919);
nand U17190 (N_17190,N_16907,N_16958);
and U17191 (N_17191,N_16876,N_16969);
and U17192 (N_17192,N_17041,N_17051);
xor U17193 (N_17193,N_16953,N_17057);
or U17194 (N_17194,N_16968,N_16999);
or U17195 (N_17195,N_16912,N_17088);
nor U17196 (N_17196,N_16940,N_16936);
xnor U17197 (N_17197,N_16826,N_17078);
and U17198 (N_17198,N_16893,N_16908);
or U17199 (N_17199,N_16974,N_16877);
nand U17200 (N_17200,N_17059,N_16890);
and U17201 (N_17201,N_16980,N_16800);
nand U17202 (N_17202,N_16820,N_16972);
xnor U17203 (N_17203,N_16857,N_17035);
or U17204 (N_17204,N_16903,N_16886);
and U17205 (N_17205,N_16863,N_16897);
and U17206 (N_17206,N_17054,N_16847);
and U17207 (N_17207,N_16827,N_17060);
nor U17208 (N_17208,N_17018,N_17010);
xnor U17209 (N_17209,N_17039,N_16978);
nor U17210 (N_17210,N_16825,N_16944);
xor U17211 (N_17211,N_16818,N_16934);
xor U17212 (N_17212,N_16805,N_17092);
or U17213 (N_17213,N_16957,N_16817);
nor U17214 (N_17214,N_17015,N_16984);
xor U17215 (N_17215,N_16920,N_16891);
nor U17216 (N_17216,N_17032,N_17062);
and U17217 (N_17217,N_17020,N_16831);
and U17218 (N_17218,N_16879,N_17094);
nor U17219 (N_17219,N_16869,N_17044);
xor U17220 (N_17220,N_16945,N_16871);
or U17221 (N_17221,N_16933,N_17036);
and U17222 (N_17222,N_17000,N_16939);
nor U17223 (N_17223,N_16822,N_16838);
nor U17224 (N_17224,N_16904,N_16924);
and U17225 (N_17225,N_16883,N_16809);
or U17226 (N_17226,N_16925,N_16878);
xnor U17227 (N_17227,N_16966,N_17086);
nor U17228 (N_17228,N_16954,N_16884);
or U17229 (N_17229,N_16949,N_17022);
or U17230 (N_17230,N_16901,N_16844);
nand U17231 (N_17231,N_17067,N_17099);
nand U17232 (N_17232,N_16910,N_16898);
xor U17233 (N_17233,N_17050,N_16808);
and U17234 (N_17234,N_16913,N_16979);
nor U17235 (N_17235,N_17087,N_16835);
or U17236 (N_17236,N_16887,N_17095);
and U17237 (N_17237,N_16833,N_16842);
or U17238 (N_17238,N_17063,N_16918);
nor U17239 (N_17239,N_17072,N_16868);
xor U17240 (N_17240,N_16952,N_17090);
nand U17241 (N_17241,N_16804,N_17034);
and U17242 (N_17242,N_16923,N_16971);
nand U17243 (N_17243,N_16815,N_16860);
and U17244 (N_17244,N_16909,N_16973);
nand U17245 (N_17245,N_17006,N_17017);
and U17246 (N_17246,N_17058,N_17033);
xnor U17247 (N_17247,N_17001,N_17038);
xnor U17248 (N_17248,N_16821,N_16962);
and U17249 (N_17249,N_16995,N_17008);
nand U17250 (N_17250,N_16814,N_16956);
or U17251 (N_17251,N_17087,N_16954);
or U17252 (N_17252,N_17021,N_16810);
nand U17253 (N_17253,N_17083,N_17010);
and U17254 (N_17254,N_17092,N_17036);
and U17255 (N_17255,N_16860,N_17007);
or U17256 (N_17256,N_16910,N_16831);
xnor U17257 (N_17257,N_16803,N_17014);
xor U17258 (N_17258,N_17062,N_17050);
and U17259 (N_17259,N_16975,N_16854);
xnor U17260 (N_17260,N_17073,N_16895);
nor U17261 (N_17261,N_17012,N_16982);
nand U17262 (N_17262,N_16890,N_16965);
xor U17263 (N_17263,N_16973,N_16914);
and U17264 (N_17264,N_16837,N_17017);
and U17265 (N_17265,N_16897,N_16806);
xnor U17266 (N_17266,N_16844,N_17005);
and U17267 (N_17267,N_16953,N_16938);
xnor U17268 (N_17268,N_16911,N_16862);
xor U17269 (N_17269,N_16955,N_16903);
nor U17270 (N_17270,N_16924,N_16910);
or U17271 (N_17271,N_16970,N_16930);
xor U17272 (N_17272,N_16830,N_16871);
or U17273 (N_17273,N_17040,N_17027);
xor U17274 (N_17274,N_16807,N_16939);
and U17275 (N_17275,N_16936,N_16856);
or U17276 (N_17276,N_17074,N_16887);
xor U17277 (N_17277,N_17059,N_17000);
xnor U17278 (N_17278,N_16927,N_16930);
and U17279 (N_17279,N_16999,N_17051);
and U17280 (N_17280,N_16955,N_16950);
and U17281 (N_17281,N_16949,N_16908);
xor U17282 (N_17282,N_17018,N_17086);
xnor U17283 (N_17283,N_17027,N_16907);
xnor U17284 (N_17284,N_17085,N_17003);
nor U17285 (N_17285,N_16831,N_16997);
and U17286 (N_17286,N_17069,N_16948);
and U17287 (N_17287,N_17029,N_17036);
nand U17288 (N_17288,N_16927,N_16943);
and U17289 (N_17289,N_17056,N_16880);
and U17290 (N_17290,N_16817,N_16866);
or U17291 (N_17291,N_16906,N_16800);
or U17292 (N_17292,N_16948,N_16988);
nor U17293 (N_17293,N_16816,N_16971);
xnor U17294 (N_17294,N_16806,N_17008);
or U17295 (N_17295,N_16886,N_17060);
nand U17296 (N_17296,N_17002,N_16814);
and U17297 (N_17297,N_16945,N_16878);
or U17298 (N_17298,N_16970,N_17037);
xnor U17299 (N_17299,N_16922,N_17057);
nor U17300 (N_17300,N_16921,N_16912);
or U17301 (N_17301,N_16867,N_16856);
nor U17302 (N_17302,N_16967,N_16960);
or U17303 (N_17303,N_16921,N_16843);
xor U17304 (N_17304,N_17077,N_16827);
xnor U17305 (N_17305,N_17058,N_16889);
xnor U17306 (N_17306,N_17036,N_16869);
or U17307 (N_17307,N_17053,N_16968);
nand U17308 (N_17308,N_17079,N_16967);
and U17309 (N_17309,N_17035,N_16966);
or U17310 (N_17310,N_16898,N_16970);
nand U17311 (N_17311,N_17082,N_17052);
xnor U17312 (N_17312,N_16959,N_17088);
or U17313 (N_17313,N_16936,N_16875);
and U17314 (N_17314,N_16950,N_16876);
or U17315 (N_17315,N_17069,N_16905);
xor U17316 (N_17316,N_16908,N_16841);
xnor U17317 (N_17317,N_16849,N_17036);
nor U17318 (N_17318,N_16973,N_16891);
and U17319 (N_17319,N_16841,N_16943);
or U17320 (N_17320,N_17039,N_17069);
or U17321 (N_17321,N_17073,N_17037);
and U17322 (N_17322,N_17062,N_16969);
nand U17323 (N_17323,N_16886,N_17047);
nor U17324 (N_17324,N_17027,N_16839);
or U17325 (N_17325,N_16966,N_16969);
xor U17326 (N_17326,N_16956,N_16985);
nor U17327 (N_17327,N_16843,N_16928);
xor U17328 (N_17328,N_16969,N_16936);
nor U17329 (N_17329,N_16854,N_16907);
and U17330 (N_17330,N_17054,N_17052);
or U17331 (N_17331,N_17091,N_16819);
or U17332 (N_17332,N_16849,N_16985);
nand U17333 (N_17333,N_17095,N_17070);
nand U17334 (N_17334,N_16868,N_16887);
xor U17335 (N_17335,N_16824,N_17067);
nor U17336 (N_17336,N_16802,N_16842);
or U17337 (N_17337,N_16970,N_16960);
nand U17338 (N_17338,N_17092,N_17006);
xnor U17339 (N_17339,N_16898,N_17077);
nor U17340 (N_17340,N_16965,N_16906);
nor U17341 (N_17341,N_17081,N_16843);
xnor U17342 (N_17342,N_16970,N_16815);
nand U17343 (N_17343,N_16948,N_17060);
nor U17344 (N_17344,N_16881,N_16854);
and U17345 (N_17345,N_16920,N_16937);
xor U17346 (N_17346,N_17037,N_16832);
nor U17347 (N_17347,N_16924,N_16931);
or U17348 (N_17348,N_16921,N_17062);
nor U17349 (N_17349,N_17078,N_16820);
nor U17350 (N_17350,N_16931,N_16826);
xnor U17351 (N_17351,N_17065,N_16997);
nor U17352 (N_17352,N_16889,N_16920);
nand U17353 (N_17353,N_16994,N_16813);
and U17354 (N_17354,N_16864,N_16818);
or U17355 (N_17355,N_16840,N_17071);
nor U17356 (N_17356,N_16887,N_16856);
and U17357 (N_17357,N_16886,N_16990);
xnor U17358 (N_17358,N_16908,N_16948);
xnor U17359 (N_17359,N_16870,N_16910);
nand U17360 (N_17360,N_17086,N_16834);
nor U17361 (N_17361,N_16896,N_17006);
or U17362 (N_17362,N_16931,N_16881);
nand U17363 (N_17363,N_16873,N_16938);
nor U17364 (N_17364,N_16874,N_16887);
nor U17365 (N_17365,N_17083,N_16926);
nand U17366 (N_17366,N_16999,N_16830);
and U17367 (N_17367,N_16966,N_16922);
or U17368 (N_17368,N_16867,N_16843);
xnor U17369 (N_17369,N_16808,N_16846);
nor U17370 (N_17370,N_16805,N_16984);
or U17371 (N_17371,N_16926,N_16904);
nor U17372 (N_17372,N_16817,N_16803);
nand U17373 (N_17373,N_16942,N_17010);
and U17374 (N_17374,N_17054,N_17024);
or U17375 (N_17375,N_16905,N_16894);
and U17376 (N_17376,N_16902,N_16988);
nor U17377 (N_17377,N_17097,N_17043);
or U17378 (N_17378,N_16823,N_16816);
nor U17379 (N_17379,N_17057,N_17065);
nor U17380 (N_17380,N_17038,N_17035);
and U17381 (N_17381,N_16849,N_16976);
xor U17382 (N_17382,N_16932,N_17022);
and U17383 (N_17383,N_16813,N_17019);
or U17384 (N_17384,N_17021,N_16838);
and U17385 (N_17385,N_16848,N_16827);
nand U17386 (N_17386,N_17067,N_16914);
nand U17387 (N_17387,N_16958,N_17042);
or U17388 (N_17388,N_16848,N_16907);
nand U17389 (N_17389,N_16903,N_16824);
xnor U17390 (N_17390,N_17007,N_17051);
or U17391 (N_17391,N_16894,N_16854);
nand U17392 (N_17392,N_17049,N_17074);
xnor U17393 (N_17393,N_17098,N_16803);
or U17394 (N_17394,N_16820,N_17049);
and U17395 (N_17395,N_17083,N_16848);
nand U17396 (N_17396,N_16864,N_17034);
nor U17397 (N_17397,N_16808,N_16950);
xnor U17398 (N_17398,N_16909,N_16836);
or U17399 (N_17399,N_17095,N_17049);
xnor U17400 (N_17400,N_17153,N_17205);
xor U17401 (N_17401,N_17211,N_17257);
nor U17402 (N_17402,N_17285,N_17200);
xor U17403 (N_17403,N_17304,N_17324);
and U17404 (N_17404,N_17279,N_17364);
and U17405 (N_17405,N_17176,N_17297);
or U17406 (N_17406,N_17278,N_17122);
and U17407 (N_17407,N_17160,N_17224);
or U17408 (N_17408,N_17262,N_17273);
nor U17409 (N_17409,N_17238,N_17107);
xnor U17410 (N_17410,N_17235,N_17294);
or U17411 (N_17411,N_17121,N_17203);
xor U17412 (N_17412,N_17112,N_17335);
and U17413 (N_17413,N_17250,N_17221);
nand U17414 (N_17414,N_17269,N_17266);
nor U17415 (N_17415,N_17334,N_17223);
nor U17416 (N_17416,N_17371,N_17254);
or U17417 (N_17417,N_17138,N_17328);
nor U17418 (N_17418,N_17299,N_17191);
nand U17419 (N_17419,N_17377,N_17378);
or U17420 (N_17420,N_17208,N_17363);
or U17421 (N_17421,N_17291,N_17379);
nand U17422 (N_17422,N_17118,N_17368);
nand U17423 (N_17423,N_17249,N_17157);
nor U17424 (N_17424,N_17240,N_17226);
and U17425 (N_17425,N_17197,N_17142);
nor U17426 (N_17426,N_17355,N_17316);
or U17427 (N_17427,N_17358,N_17166);
or U17428 (N_17428,N_17325,N_17244);
or U17429 (N_17429,N_17380,N_17275);
nand U17430 (N_17430,N_17111,N_17163);
or U17431 (N_17431,N_17286,N_17232);
or U17432 (N_17432,N_17337,N_17156);
xnor U17433 (N_17433,N_17330,N_17336);
nor U17434 (N_17434,N_17346,N_17247);
and U17435 (N_17435,N_17161,N_17222);
nand U17436 (N_17436,N_17341,N_17149);
nand U17437 (N_17437,N_17241,N_17272);
xor U17438 (N_17438,N_17227,N_17154);
nand U17439 (N_17439,N_17356,N_17395);
nand U17440 (N_17440,N_17229,N_17323);
nor U17441 (N_17441,N_17217,N_17125);
nor U17442 (N_17442,N_17196,N_17102);
or U17443 (N_17443,N_17347,N_17296);
and U17444 (N_17444,N_17135,N_17362);
xnor U17445 (N_17445,N_17137,N_17220);
and U17446 (N_17446,N_17155,N_17381);
and U17447 (N_17447,N_17116,N_17327);
and U17448 (N_17448,N_17390,N_17169);
and U17449 (N_17449,N_17367,N_17357);
nand U17450 (N_17450,N_17225,N_17302);
and U17451 (N_17451,N_17300,N_17369);
nor U17452 (N_17452,N_17314,N_17234);
and U17453 (N_17453,N_17150,N_17298);
xnor U17454 (N_17454,N_17237,N_17168);
and U17455 (N_17455,N_17216,N_17382);
and U17456 (N_17456,N_17104,N_17180);
and U17457 (N_17457,N_17398,N_17255);
xor U17458 (N_17458,N_17287,N_17148);
nand U17459 (N_17459,N_17373,N_17342);
or U17460 (N_17460,N_17389,N_17282);
nand U17461 (N_17461,N_17361,N_17393);
and U17462 (N_17462,N_17386,N_17397);
nand U17463 (N_17463,N_17271,N_17119);
and U17464 (N_17464,N_17280,N_17186);
and U17465 (N_17465,N_17248,N_17376);
or U17466 (N_17466,N_17326,N_17396);
or U17467 (N_17467,N_17320,N_17394);
and U17468 (N_17468,N_17352,N_17242);
or U17469 (N_17469,N_17338,N_17312);
nand U17470 (N_17470,N_17190,N_17214);
nor U17471 (N_17471,N_17259,N_17231);
nand U17472 (N_17472,N_17195,N_17295);
and U17473 (N_17473,N_17129,N_17167);
or U17474 (N_17474,N_17201,N_17359);
nand U17475 (N_17475,N_17170,N_17130);
nand U17476 (N_17476,N_17184,N_17159);
or U17477 (N_17477,N_17311,N_17263);
and U17478 (N_17478,N_17332,N_17132);
nand U17479 (N_17479,N_17268,N_17264);
nor U17480 (N_17480,N_17383,N_17276);
xnor U17481 (N_17481,N_17145,N_17188);
or U17482 (N_17482,N_17318,N_17139);
nor U17483 (N_17483,N_17215,N_17164);
xnor U17484 (N_17484,N_17349,N_17251);
nand U17485 (N_17485,N_17113,N_17308);
or U17486 (N_17486,N_17109,N_17124);
nor U17487 (N_17487,N_17131,N_17319);
nand U17488 (N_17488,N_17245,N_17385);
and U17489 (N_17489,N_17366,N_17175);
xnor U17490 (N_17490,N_17140,N_17270);
and U17491 (N_17491,N_17100,N_17290);
and U17492 (N_17492,N_17136,N_17277);
nor U17493 (N_17493,N_17350,N_17147);
xnor U17494 (N_17494,N_17115,N_17199);
and U17495 (N_17495,N_17182,N_17152);
nor U17496 (N_17496,N_17339,N_17303);
nor U17497 (N_17497,N_17370,N_17246);
xnor U17498 (N_17498,N_17236,N_17392);
nor U17499 (N_17499,N_17210,N_17194);
nor U17500 (N_17500,N_17114,N_17239);
or U17501 (N_17501,N_17123,N_17120);
nand U17502 (N_17502,N_17261,N_17253);
nand U17503 (N_17503,N_17348,N_17134);
or U17504 (N_17504,N_17384,N_17256);
nand U17505 (N_17505,N_17126,N_17228);
nor U17506 (N_17506,N_17258,N_17172);
or U17507 (N_17507,N_17305,N_17174);
or U17508 (N_17508,N_17365,N_17333);
or U17509 (N_17509,N_17307,N_17179);
nor U17510 (N_17510,N_17207,N_17162);
or U17511 (N_17511,N_17322,N_17212);
xor U17512 (N_17512,N_17372,N_17313);
nor U17513 (N_17513,N_17354,N_17151);
nand U17514 (N_17514,N_17105,N_17213);
xnor U17515 (N_17515,N_17306,N_17388);
nand U17516 (N_17516,N_17292,N_17181);
nand U17517 (N_17517,N_17351,N_17144);
xnor U17518 (N_17518,N_17283,N_17202);
xor U17519 (N_17519,N_17143,N_17281);
or U17520 (N_17520,N_17301,N_17391);
nor U17521 (N_17521,N_17165,N_17274);
or U17522 (N_17522,N_17128,N_17204);
xor U17523 (N_17523,N_17193,N_17108);
nor U17524 (N_17524,N_17141,N_17178);
nand U17525 (N_17525,N_17189,N_17192);
nor U17526 (N_17526,N_17206,N_17230);
nor U17527 (N_17527,N_17387,N_17233);
or U17528 (N_17528,N_17185,N_17127);
xor U17529 (N_17529,N_17284,N_17173);
nor U17530 (N_17530,N_17293,N_17315);
nand U17531 (N_17531,N_17260,N_17177);
xnor U17532 (N_17532,N_17374,N_17219);
or U17533 (N_17533,N_17198,N_17331);
nand U17534 (N_17534,N_17343,N_17310);
or U17535 (N_17535,N_17218,N_17353);
nand U17536 (N_17536,N_17243,N_17103);
nor U17537 (N_17537,N_17133,N_17183);
nor U17538 (N_17538,N_17110,N_17288);
and U17539 (N_17539,N_17158,N_17340);
nor U17540 (N_17540,N_17345,N_17309);
and U17541 (N_17541,N_17399,N_17375);
nand U17542 (N_17542,N_17329,N_17317);
nor U17543 (N_17543,N_17106,N_17252);
and U17544 (N_17544,N_17267,N_17146);
and U17545 (N_17545,N_17321,N_17344);
nor U17546 (N_17546,N_17209,N_17101);
nand U17547 (N_17547,N_17360,N_17171);
and U17548 (N_17548,N_17117,N_17265);
nor U17549 (N_17549,N_17289,N_17187);
nor U17550 (N_17550,N_17203,N_17308);
and U17551 (N_17551,N_17282,N_17281);
xnor U17552 (N_17552,N_17216,N_17159);
and U17553 (N_17553,N_17227,N_17252);
xnor U17554 (N_17554,N_17109,N_17296);
xnor U17555 (N_17555,N_17122,N_17267);
nor U17556 (N_17556,N_17136,N_17275);
xnor U17557 (N_17557,N_17305,N_17244);
nor U17558 (N_17558,N_17230,N_17338);
nand U17559 (N_17559,N_17388,N_17284);
and U17560 (N_17560,N_17139,N_17390);
or U17561 (N_17561,N_17306,N_17173);
and U17562 (N_17562,N_17175,N_17363);
xnor U17563 (N_17563,N_17366,N_17290);
nor U17564 (N_17564,N_17255,N_17330);
and U17565 (N_17565,N_17324,N_17201);
xor U17566 (N_17566,N_17175,N_17389);
nand U17567 (N_17567,N_17394,N_17135);
xor U17568 (N_17568,N_17217,N_17233);
xor U17569 (N_17569,N_17253,N_17159);
or U17570 (N_17570,N_17343,N_17135);
or U17571 (N_17571,N_17233,N_17306);
nand U17572 (N_17572,N_17165,N_17375);
or U17573 (N_17573,N_17373,N_17272);
and U17574 (N_17574,N_17183,N_17347);
xnor U17575 (N_17575,N_17303,N_17360);
nand U17576 (N_17576,N_17105,N_17232);
nand U17577 (N_17577,N_17294,N_17258);
and U17578 (N_17578,N_17359,N_17200);
or U17579 (N_17579,N_17219,N_17322);
xor U17580 (N_17580,N_17185,N_17115);
nand U17581 (N_17581,N_17221,N_17373);
or U17582 (N_17582,N_17244,N_17153);
or U17583 (N_17583,N_17337,N_17100);
or U17584 (N_17584,N_17149,N_17223);
and U17585 (N_17585,N_17252,N_17303);
and U17586 (N_17586,N_17296,N_17395);
nor U17587 (N_17587,N_17268,N_17350);
and U17588 (N_17588,N_17179,N_17100);
or U17589 (N_17589,N_17189,N_17160);
nand U17590 (N_17590,N_17120,N_17369);
and U17591 (N_17591,N_17115,N_17264);
xor U17592 (N_17592,N_17214,N_17290);
or U17593 (N_17593,N_17398,N_17392);
nand U17594 (N_17594,N_17224,N_17301);
nand U17595 (N_17595,N_17375,N_17179);
xor U17596 (N_17596,N_17308,N_17146);
and U17597 (N_17597,N_17166,N_17219);
nor U17598 (N_17598,N_17219,N_17109);
nand U17599 (N_17599,N_17308,N_17147);
xnor U17600 (N_17600,N_17167,N_17254);
or U17601 (N_17601,N_17291,N_17337);
nand U17602 (N_17602,N_17233,N_17345);
or U17603 (N_17603,N_17394,N_17163);
and U17604 (N_17604,N_17278,N_17121);
xnor U17605 (N_17605,N_17316,N_17244);
nand U17606 (N_17606,N_17343,N_17318);
and U17607 (N_17607,N_17335,N_17347);
xor U17608 (N_17608,N_17299,N_17204);
nand U17609 (N_17609,N_17185,N_17309);
or U17610 (N_17610,N_17146,N_17175);
xor U17611 (N_17611,N_17355,N_17338);
xor U17612 (N_17612,N_17169,N_17276);
nand U17613 (N_17613,N_17326,N_17209);
xnor U17614 (N_17614,N_17158,N_17384);
nor U17615 (N_17615,N_17312,N_17246);
nand U17616 (N_17616,N_17296,N_17224);
and U17617 (N_17617,N_17266,N_17158);
xnor U17618 (N_17618,N_17144,N_17305);
nor U17619 (N_17619,N_17172,N_17130);
xnor U17620 (N_17620,N_17112,N_17150);
nor U17621 (N_17621,N_17139,N_17161);
nor U17622 (N_17622,N_17378,N_17394);
nand U17623 (N_17623,N_17140,N_17230);
xnor U17624 (N_17624,N_17390,N_17168);
and U17625 (N_17625,N_17332,N_17277);
nor U17626 (N_17626,N_17381,N_17130);
xnor U17627 (N_17627,N_17256,N_17171);
or U17628 (N_17628,N_17221,N_17343);
or U17629 (N_17629,N_17128,N_17308);
xor U17630 (N_17630,N_17157,N_17128);
nand U17631 (N_17631,N_17141,N_17382);
or U17632 (N_17632,N_17150,N_17139);
and U17633 (N_17633,N_17290,N_17331);
nand U17634 (N_17634,N_17159,N_17324);
xor U17635 (N_17635,N_17236,N_17170);
xnor U17636 (N_17636,N_17394,N_17386);
nand U17637 (N_17637,N_17332,N_17237);
nand U17638 (N_17638,N_17239,N_17308);
xnor U17639 (N_17639,N_17181,N_17336);
nand U17640 (N_17640,N_17246,N_17282);
xnor U17641 (N_17641,N_17353,N_17220);
and U17642 (N_17642,N_17127,N_17243);
xnor U17643 (N_17643,N_17236,N_17293);
or U17644 (N_17644,N_17341,N_17108);
and U17645 (N_17645,N_17264,N_17395);
and U17646 (N_17646,N_17201,N_17345);
nor U17647 (N_17647,N_17149,N_17297);
or U17648 (N_17648,N_17219,N_17317);
nor U17649 (N_17649,N_17265,N_17274);
or U17650 (N_17650,N_17240,N_17344);
nand U17651 (N_17651,N_17260,N_17118);
or U17652 (N_17652,N_17228,N_17149);
nand U17653 (N_17653,N_17319,N_17294);
xnor U17654 (N_17654,N_17129,N_17338);
and U17655 (N_17655,N_17126,N_17357);
nand U17656 (N_17656,N_17369,N_17334);
nor U17657 (N_17657,N_17261,N_17299);
nor U17658 (N_17658,N_17318,N_17314);
xor U17659 (N_17659,N_17217,N_17357);
nand U17660 (N_17660,N_17284,N_17168);
or U17661 (N_17661,N_17307,N_17158);
xor U17662 (N_17662,N_17137,N_17353);
nor U17663 (N_17663,N_17398,N_17254);
nand U17664 (N_17664,N_17320,N_17298);
nand U17665 (N_17665,N_17393,N_17396);
or U17666 (N_17666,N_17305,N_17374);
xnor U17667 (N_17667,N_17371,N_17216);
or U17668 (N_17668,N_17383,N_17181);
xor U17669 (N_17669,N_17379,N_17108);
or U17670 (N_17670,N_17187,N_17179);
nor U17671 (N_17671,N_17148,N_17290);
nor U17672 (N_17672,N_17230,N_17377);
nor U17673 (N_17673,N_17117,N_17287);
xor U17674 (N_17674,N_17392,N_17300);
nand U17675 (N_17675,N_17259,N_17209);
nand U17676 (N_17676,N_17114,N_17392);
and U17677 (N_17677,N_17126,N_17223);
nand U17678 (N_17678,N_17162,N_17113);
and U17679 (N_17679,N_17322,N_17280);
and U17680 (N_17680,N_17222,N_17361);
nand U17681 (N_17681,N_17317,N_17397);
xor U17682 (N_17682,N_17361,N_17278);
or U17683 (N_17683,N_17185,N_17172);
nor U17684 (N_17684,N_17139,N_17239);
xor U17685 (N_17685,N_17285,N_17120);
nand U17686 (N_17686,N_17269,N_17288);
and U17687 (N_17687,N_17363,N_17340);
nor U17688 (N_17688,N_17221,N_17386);
nand U17689 (N_17689,N_17264,N_17342);
nand U17690 (N_17690,N_17203,N_17360);
and U17691 (N_17691,N_17338,N_17175);
and U17692 (N_17692,N_17397,N_17290);
or U17693 (N_17693,N_17285,N_17111);
and U17694 (N_17694,N_17111,N_17293);
and U17695 (N_17695,N_17300,N_17306);
nor U17696 (N_17696,N_17337,N_17211);
xnor U17697 (N_17697,N_17106,N_17184);
nand U17698 (N_17698,N_17162,N_17164);
nand U17699 (N_17699,N_17339,N_17102);
nor U17700 (N_17700,N_17410,N_17478);
nor U17701 (N_17701,N_17682,N_17536);
nand U17702 (N_17702,N_17474,N_17551);
and U17703 (N_17703,N_17577,N_17592);
and U17704 (N_17704,N_17658,N_17548);
or U17705 (N_17705,N_17683,N_17659);
nand U17706 (N_17706,N_17624,N_17453);
and U17707 (N_17707,N_17586,N_17441);
or U17708 (N_17708,N_17581,N_17429);
or U17709 (N_17709,N_17483,N_17442);
nand U17710 (N_17710,N_17665,N_17531);
and U17711 (N_17711,N_17402,N_17675);
nand U17712 (N_17712,N_17469,N_17457);
nand U17713 (N_17713,N_17666,N_17496);
or U17714 (N_17714,N_17595,N_17468);
nand U17715 (N_17715,N_17549,N_17564);
nand U17716 (N_17716,N_17590,N_17699);
xor U17717 (N_17717,N_17561,N_17427);
xnor U17718 (N_17718,N_17506,N_17677);
nor U17719 (N_17719,N_17504,N_17602);
and U17720 (N_17720,N_17588,N_17597);
nand U17721 (N_17721,N_17641,N_17634);
or U17722 (N_17722,N_17511,N_17430);
nand U17723 (N_17723,N_17609,N_17480);
or U17724 (N_17724,N_17567,N_17539);
nand U17725 (N_17725,N_17637,N_17559);
or U17726 (N_17726,N_17670,N_17458);
or U17727 (N_17727,N_17556,N_17565);
xnor U17728 (N_17728,N_17685,N_17403);
nor U17729 (N_17729,N_17555,N_17582);
or U17730 (N_17730,N_17495,N_17423);
nor U17731 (N_17731,N_17507,N_17547);
xnor U17732 (N_17732,N_17412,N_17618);
or U17733 (N_17733,N_17678,N_17640);
or U17734 (N_17734,N_17541,N_17428);
and U17735 (N_17735,N_17572,N_17575);
or U17736 (N_17736,N_17638,N_17432);
and U17737 (N_17737,N_17407,N_17434);
and U17738 (N_17738,N_17585,N_17414);
nand U17739 (N_17739,N_17463,N_17594);
xnor U17740 (N_17740,N_17426,N_17542);
and U17741 (N_17741,N_17464,N_17569);
nand U17742 (N_17742,N_17574,N_17604);
or U17743 (N_17743,N_17409,N_17697);
xor U17744 (N_17744,N_17573,N_17443);
xnor U17745 (N_17745,N_17523,N_17627);
nand U17746 (N_17746,N_17466,N_17562);
and U17747 (N_17747,N_17571,N_17681);
or U17748 (N_17748,N_17625,N_17450);
nand U17749 (N_17749,N_17516,N_17525);
or U17750 (N_17750,N_17690,N_17519);
nor U17751 (N_17751,N_17522,N_17467);
and U17752 (N_17752,N_17417,N_17653);
nand U17753 (N_17753,N_17596,N_17687);
and U17754 (N_17754,N_17517,N_17411);
nand U17755 (N_17755,N_17643,N_17494);
and U17756 (N_17756,N_17521,N_17461);
and U17757 (N_17757,N_17626,N_17557);
nand U17758 (N_17758,N_17419,N_17405);
xor U17759 (N_17759,N_17485,N_17465);
xor U17760 (N_17760,N_17598,N_17647);
nor U17761 (N_17761,N_17663,N_17433);
nand U17762 (N_17762,N_17477,N_17578);
or U17763 (N_17763,N_17619,N_17648);
xnor U17764 (N_17764,N_17470,N_17669);
or U17765 (N_17765,N_17520,N_17591);
xnor U17766 (N_17766,N_17688,N_17664);
xor U17767 (N_17767,N_17420,N_17438);
or U17768 (N_17768,N_17694,N_17608);
nor U17769 (N_17769,N_17656,N_17473);
and U17770 (N_17770,N_17605,N_17462);
xnor U17771 (N_17771,N_17679,N_17482);
nand U17772 (N_17772,N_17632,N_17689);
or U17773 (N_17773,N_17460,N_17532);
nand U17774 (N_17774,N_17513,N_17489);
or U17775 (N_17775,N_17554,N_17538);
and U17776 (N_17776,N_17501,N_17580);
nor U17777 (N_17777,N_17472,N_17503);
nor U17778 (N_17778,N_17667,N_17543);
nor U17779 (N_17779,N_17589,N_17654);
nor U17780 (N_17780,N_17673,N_17639);
and U17781 (N_17781,N_17599,N_17437);
or U17782 (N_17782,N_17451,N_17490);
nor U17783 (N_17783,N_17454,N_17487);
nor U17784 (N_17784,N_17509,N_17445);
nor U17785 (N_17785,N_17644,N_17421);
or U17786 (N_17786,N_17449,N_17695);
and U17787 (N_17787,N_17610,N_17518);
nor U17788 (N_17788,N_17439,N_17440);
or U17789 (N_17789,N_17413,N_17540);
or U17790 (N_17790,N_17416,N_17533);
or U17791 (N_17791,N_17649,N_17435);
xnor U17792 (N_17792,N_17651,N_17661);
or U17793 (N_17793,N_17424,N_17422);
or U17794 (N_17794,N_17479,N_17500);
xor U17795 (N_17795,N_17606,N_17534);
or U17796 (N_17796,N_17415,N_17530);
xnor U17797 (N_17797,N_17512,N_17635);
nor U17798 (N_17798,N_17493,N_17404);
nand U17799 (N_17799,N_17447,N_17436);
xor U17800 (N_17800,N_17459,N_17444);
or U17801 (N_17801,N_17537,N_17524);
nor U17802 (N_17802,N_17455,N_17502);
and U17803 (N_17803,N_17498,N_17552);
and U17804 (N_17804,N_17613,N_17611);
xor U17805 (N_17805,N_17508,N_17452);
or U17806 (N_17806,N_17566,N_17629);
xor U17807 (N_17807,N_17545,N_17528);
or U17808 (N_17808,N_17499,N_17584);
nor U17809 (N_17809,N_17676,N_17620);
xnor U17810 (N_17810,N_17671,N_17680);
xnor U17811 (N_17811,N_17628,N_17527);
xnor U17812 (N_17812,N_17481,N_17550);
xor U17813 (N_17813,N_17630,N_17431);
nor U17814 (N_17814,N_17486,N_17579);
xor U17815 (N_17815,N_17510,N_17617);
nand U17816 (N_17816,N_17633,N_17615);
nand U17817 (N_17817,N_17446,N_17497);
and U17818 (N_17818,N_17686,N_17563);
xor U17819 (N_17819,N_17526,N_17607);
nand U17820 (N_17820,N_17660,N_17698);
nand U17821 (N_17821,N_17612,N_17515);
nand U17822 (N_17822,N_17576,N_17621);
or U17823 (N_17823,N_17691,N_17645);
xor U17824 (N_17824,N_17408,N_17505);
and U17825 (N_17825,N_17616,N_17560);
xor U17826 (N_17826,N_17668,N_17488);
nor U17827 (N_17827,N_17492,N_17587);
and U17828 (N_17828,N_17568,N_17406);
and U17829 (N_17829,N_17514,N_17583);
nand U17830 (N_17830,N_17593,N_17544);
nand U17831 (N_17831,N_17692,N_17642);
nor U17832 (N_17832,N_17603,N_17696);
xor U17833 (N_17833,N_17622,N_17646);
or U17834 (N_17834,N_17623,N_17674);
xnor U17835 (N_17835,N_17491,N_17614);
xor U17836 (N_17836,N_17401,N_17425);
and U17837 (N_17837,N_17600,N_17529);
nand U17838 (N_17838,N_17662,N_17570);
nor U17839 (N_17839,N_17456,N_17553);
xor U17840 (N_17840,N_17655,N_17672);
nand U17841 (N_17841,N_17652,N_17558);
or U17842 (N_17842,N_17601,N_17475);
nor U17843 (N_17843,N_17657,N_17684);
nor U17844 (N_17844,N_17400,N_17448);
xnor U17845 (N_17845,N_17418,N_17636);
or U17846 (N_17846,N_17476,N_17650);
nand U17847 (N_17847,N_17546,N_17535);
nor U17848 (N_17848,N_17631,N_17471);
nand U17849 (N_17849,N_17484,N_17693);
or U17850 (N_17850,N_17606,N_17653);
xor U17851 (N_17851,N_17404,N_17433);
xor U17852 (N_17852,N_17565,N_17445);
or U17853 (N_17853,N_17680,N_17456);
or U17854 (N_17854,N_17503,N_17611);
nand U17855 (N_17855,N_17430,N_17515);
xnor U17856 (N_17856,N_17695,N_17490);
nand U17857 (N_17857,N_17645,N_17669);
and U17858 (N_17858,N_17417,N_17594);
nand U17859 (N_17859,N_17572,N_17616);
or U17860 (N_17860,N_17487,N_17402);
nor U17861 (N_17861,N_17688,N_17413);
xnor U17862 (N_17862,N_17525,N_17551);
or U17863 (N_17863,N_17488,N_17623);
and U17864 (N_17864,N_17562,N_17407);
or U17865 (N_17865,N_17624,N_17572);
and U17866 (N_17866,N_17418,N_17632);
and U17867 (N_17867,N_17433,N_17638);
nand U17868 (N_17868,N_17520,N_17463);
or U17869 (N_17869,N_17497,N_17585);
nor U17870 (N_17870,N_17435,N_17547);
or U17871 (N_17871,N_17465,N_17608);
and U17872 (N_17872,N_17659,N_17484);
xnor U17873 (N_17873,N_17446,N_17543);
nor U17874 (N_17874,N_17598,N_17682);
xnor U17875 (N_17875,N_17497,N_17556);
nor U17876 (N_17876,N_17644,N_17419);
and U17877 (N_17877,N_17667,N_17586);
or U17878 (N_17878,N_17659,N_17590);
xnor U17879 (N_17879,N_17558,N_17542);
xor U17880 (N_17880,N_17441,N_17578);
or U17881 (N_17881,N_17596,N_17410);
nand U17882 (N_17882,N_17682,N_17448);
xor U17883 (N_17883,N_17516,N_17434);
xnor U17884 (N_17884,N_17456,N_17449);
xnor U17885 (N_17885,N_17584,N_17411);
xnor U17886 (N_17886,N_17492,N_17595);
xor U17887 (N_17887,N_17507,N_17676);
or U17888 (N_17888,N_17593,N_17572);
or U17889 (N_17889,N_17670,N_17418);
nand U17890 (N_17890,N_17472,N_17479);
nor U17891 (N_17891,N_17417,N_17483);
and U17892 (N_17892,N_17668,N_17621);
xnor U17893 (N_17893,N_17693,N_17564);
xnor U17894 (N_17894,N_17630,N_17452);
or U17895 (N_17895,N_17652,N_17613);
nor U17896 (N_17896,N_17651,N_17576);
nand U17897 (N_17897,N_17491,N_17461);
nor U17898 (N_17898,N_17543,N_17535);
nor U17899 (N_17899,N_17613,N_17424);
nand U17900 (N_17900,N_17433,N_17443);
nand U17901 (N_17901,N_17620,N_17458);
and U17902 (N_17902,N_17411,N_17595);
and U17903 (N_17903,N_17529,N_17495);
and U17904 (N_17904,N_17504,N_17559);
xor U17905 (N_17905,N_17442,N_17510);
nor U17906 (N_17906,N_17551,N_17568);
and U17907 (N_17907,N_17596,N_17487);
and U17908 (N_17908,N_17670,N_17543);
or U17909 (N_17909,N_17524,N_17441);
nor U17910 (N_17910,N_17536,N_17577);
nor U17911 (N_17911,N_17493,N_17616);
or U17912 (N_17912,N_17686,N_17628);
nand U17913 (N_17913,N_17552,N_17466);
or U17914 (N_17914,N_17435,N_17607);
or U17915 (N_17915,N_17676,N_17455);
or U17916 (N_17916,N_17519,N_17605);
xor U17917 (N_17917,N_17615,N_17428);
or U17918 (N_17918,N_17620,N_17434);
or U17919 (N_17919,N_17532,N_17413);
nand U17920 (N_17920,N_17479,N_17562);
and U17921 (N_17921,N_17597,N_17602);
and U17922 (N_17922,N_17646,N_17659);
xor U17923 (N_17923,N_17698,N_17560);
and U17924 (N_17924,N_17493,N_17537);
nand U17925 (N_17925,N_17401,N_17413);
and U17926 (N_17926,N_17480,N_17479);
and U17927 (N_17927,N_17480,N_17486);
or U17928 (N_17928,N_17603,N_17571);
xor U17929 (N_17929,N_17643,N_17527);
nand U17930 (N_17930,N_17448,N_17540);
and U17931 (N_17931,N_17565,N_17620);
and U17932 (N_17932,N_17646,N_17469);
and U17933 (N_17933,N_17613,N_17594);
xor U17934 (N_17934,N_17694,N_17563);
nor U17935 (N_17935,N_17431,N_17569);
nand U17936 (N_17936,N_17605,N_17407);
or U17937 (N_17937,N_17616,N_17591);
or U17938 (N_17938,N_17553,N_17612);
and U17939 (N_17939,N_17601,N_17407);
nand U17940 (N_17940,N_17479,N_17694);
or U17941 (N_17941,N_17647,N_17612);
xnor U17942 (N_17942,N_17597,N_17528);
and U17943 (N_17943,N_17611,N_17429);
xor U17944 (N_17944,N_17687,N_17627);
nand U17945 (N_17945,N_17621,N_17633);
and U17946 (N_17946,N_17548,N_17639);
and U17947 (N_17947,N_17431,N_17612);
nor U17948 (N_17948,N_17569,N_17435);
or U17949 (N_17949,N_17697,N_17423);
xnor U17950 (N_17950,N_17469,N_17586);
xnor U17951 (N_17951,N_17548,N_17690);
nor U17952 (N_17952,N_17605,N_17448);
and U17953 (N_17953,N_17402,N_17427);
xnor U17954 (N_17954,N_17652,N_17480);
xnor U17955 (N_17955,N_17517,N_17610);
nor U17956 (N_17956,N_17582,N_17445);
nand U17957 (N_17957,N_17699,N_17440);
or U17958 (N_17958,N_17418,N_17675);
nor U17959 (N_17959,N_17630,N_17529);
or U17960 (N_17960,N_17409,N_17515);
xor U17961 (N_17961,N_17558,N_17623);
or U17962 (N_17962,N_17526,N_17529);
and U17963 (N_17963,N_17588,N_17670);
and U17964 (N_17964,N_17581,N_17426);
nor U17965 (N_17965,N_17444,N_17464);
or U17966 (N_17966,N_17526,N_17691);
xor U17967 (N_17967,N_17520,N_17505);
xor U17968 (N_17968,N_17421,N_17645);
nor U17969 (N_17969,N_17530,N_17413);
and U17970 (N_17970,N_17534,N_17501);
nor U17971 (N_17971,N_17572,N_17534);
and U17972 (N_17972,N_17539,N_17596);
nand U17973 (N_17973,N_17629,N_17407);
or U17974 (N_17974,N_17503,N_17603);
xor U17975 (N_17975,N_17551,N_17554);
xnor U17976 (N_17976,N_17539,N_17432);
nand U17977 (N_17977,N_17462,N_17428);
or U17978 (N_17978,N_17646,N_17540);
nor U17979 (N_17979,N_17422,N_17431);
nand U17980 (N_17980,N_17642,N_17411);
xnor U17981 (N_17981,N_17649,N_17487);
nand U17982 (N_17982,N_17450,N_17445);
and U17983 (N_17983,N_17595,N_17420);
xnor U17984 (N_17984,N_17504,N_17615);
nand U17985 (N_17985,N_17662,N_17676);
or U17986 (N_17986,N_17565,N_17558);
and U17987 (N_17987,N_17491,N_17604);
or U17988 (N_17988,N_17593,N_17634);
nand U17989 (N_17989,N_17465,N_17538);
and U17990 (N_17990,N_17436,N_17545);
and U17991 (N_17991,N_17451,N_17482);
or U17992 (N_17992,N_17546,N_17693);
nand U17993 (N_17993,N_17444,N_17522);
or U17994 (N_17994,N_17656,N_17548);
and U17995 (N_17995,N_17691,N_17648);
nor U17996 (N_17996,N_17463,N_17402);
nor U17997 (N_17997,N_17690,N_17567);
nand U17998 (N_17998,N_17625,N_17655);
nor U17999 (N_17999,N_17652,N_17509);
and U18000 (N_18000,N_17954,N_17744);
xor U18001 (N_18001,N_17988,N_17930);
and U18002 (N_18002,N_17980,N_17967);
nor U18003 (N_18003,N_17764,N_17853);
nand U18004 (N_18004,N_17736,N_17915);
xnor U18005 (N_18005,N_17724,N_17788);
and U18006 (N_18006,N_17892,N_17798);
or U18007 (N_18007,N_17821,N_17904);
nor U18008 (N_18008,N_17709,N_17971);
xnor U18009 (N_18009,N_17845,N_17813);
and U18010 (N_18010,N_17885,N_17778);
and U18011 (N_18011,N_17718,N_17893);
nor U18012 (N_18012,N_17909,N_17983);
and U18013 (N_18013,N_17940,N_17874);
nor U18014 (N_18014,N_17923,N_17876);
nand U18015 (N_18015,N_17721,N_17762);
nor U18016 (N_18016,N_17975,N_17819);
xor U18017 (N_18017,N_17816,N_17838);
nand U18018 (N_18018,N_17911,N_17942);
or U18019 (N_18019,N_17842,N_17922);
nand U18020 (N_18020,N_17831,N_17896);
xor U18021 (N_18021,N_17886,N_17841);
and U18022 (N_18022,N_17800,N_17960);
nand U18023 (N_18023,N_17818,N_17792);
and U18024 (N_18024,N_17747,N_17977);
and U18025 (N_18025,N_17864,N_17972);
and U18026 (N_18026,N_17847,N_17903);
or U18027 (N_18027,N_17997,N_17740);
or U18028 (N_18028,N_17839,N_17772);
nor U18029 (N_18029,N_17700,N_17925);
and U18030 (N_18030,N_17739,N_17873);
xnor U18031 (N_18031,N_17716,N_17731);
xnor U18032 (N_18032,N_17982,N_17941);
or U18033 (N_18033,N_17926,N_17797);
and U18034 (N_18034,N_17801,N_17761);
or U18035 (N_18035,N_17745,N_17871);
nor U18036 (N_18036,N_17882,N_17757);
xor U18037 (N_18037,N_17832,N_17751);
xnor U18038 (N_18038,N_17949,N_17962);
nor U18039 (N_18039,N_17730,N_17998);
nor U18040 (N_18040,N_17992,N_17888);
nor U18041 (N_18041,N_17770,N_17902);
and U18042 (N_18042,N_17914,N_17900);
xnor U18043 (N_18043,N_17704,N_17765);
nand U18044 (N_18044,N_17701,N_17866);
nor U18045 (N_18045,N_17848,N_17991);
or U18046 (N_18046,N_17970,N_17867);
and U18047 (N_18047,N_17766,N_17937);
xor U18048 (N_18048,N_17944,N_17771);
and U18049 (N_18049,N_17933,N_17833);
nor U18050 (N_18050,N_17861,N_17965);
and U18051 (N_18051,N_17990,N_17763);
xor U18052 (N_18052,N_17830,N_17768);
nor U18053 (N_18053,N_17702,N_17817);
or U18054 (N_18054,N_17750,N_17907);
xnor U18055 (N_18055,N_17826,N_17946);
nand U18056 (N_18056,N_17795,N_17979);
nor U18057 (N_18057,N_17823,N_17985);
and U18058 (N_18058,N_17755,N_17934);
and U18059 (N_18059,N_17780,N_17722);
or U18060 (N_18060,N_17756,N_17857);
or U18061 (N_18061,N_17956,N_17735);
nor U18062 (N_18062,N_17727,N_17791);
or U18063 (N_18063,N_17726,N_17929);
and U18064 (N_18064,N_17938,N_17805);
nor U18065 (N_18065,N_17889,N_17835);
xor U18066 (N_18066,N_17849,N_17917);
and U18067 (N_18067,N_17981,N_17734);
or U18068 (N_18068,N_17928,N_17943);
and U18069 (N_18069,N_17905,N_17748);
or U18070 (N_18070,N_17738,N_17746);
xor U18071 (N_18071,N_17884,N_17963);
nand U18072 (N_18072,N_17913,N_17872);
or U18073 (N_18073,N_17959,N_17955);
nor U18074 (N_18074,N_17712,N_17879);
or U18075 (N_18075,N_17786,N_17968);
and U18076 (N_18076,N_17978,N_17749);
nand U18077 (N_18077,N_17790,N_17808);
and U18078 (N_18078,N_17912,N_17927);
nand U18079 (N_18079,N_17875,N_17843);
xor U18080 (N_18080,N_17758,N_17899);
xnor U18081 (N_18081,N_17860,N_17769);
and U18082 (N_18082,N_17901,N_17741);
or U18083 (N_18083,N_17767,N_17793);
nand U18084 (N_18084,N_17785,N_17865);
or U18085 (N_18085,N_17759,N_17862);
nor U18086 (N_18086,N_17891,N_17775);
and U18087 (N_18087,N_17812,N_17969);
or U18088 (N_18088,N_17811,N_17733);
or U18089 (N_18089,N_17868,N_17999);
nor U18090 (N_18090,N_17952,N_17883);
nor U18091 (N_18091,N_17707,N_17732);
xnor U18092 (N_18092,N_17713,N_17994);
nand U18093 (N_18093,N_17824,N_17920);
and U18094 (N_18094,N_17710,N_17881);
nor U18095 (N_18095,N_17945,N_17863);
xor U18096 (N_18096,N_17895,N_17728);
nand U18097 (N_18097,N_17825,N_17807);
nor U18098 (N_18098,N_17752,N_17851);
and U18099 (N_18099,N_17737,N_17995);
xnor U18100 (N_18100,N_17957,N_17951);
or U18101 (N_18101,N_17987,N_17958);
or U18102 (N_18102,N_17779,N_17815);
nand U18103 (N_18103,N_17802,N_17859);
and U18104 (N_18104,N_17711,N_17754);
nor U18105 (N_18105,N_17715,N_17924);
or U18106 (N_18106,N_17809,N_17753);
nor U18107 (N_18107,N_17878,N_17950);
xor U18108 (N_18108,N_17774,N_17717);
xnor U18109 (N_18109,N_17939,N_17989);
or U18110 (N_18110,N_17858,N_17789);
and U18111 (N_18111,N_17720,N_17725);
or U18112 (N_18112,N_17856,N_17953);
or U18113 (N_18113,N_17996,N_17799);
nor U18114 (N_18114,N_17708,N_17837);
nor U18115 (N_18115,N_17852,N_17840);
nand U18116 (N_18116,N_17935,N_17908);
and U18117 (N_18117,N_17828,N_17964);
and U18118 (N_18118,N_17887,N_17973);
xnor U18119 (N_18119,N_17760,N_17846);
and U18120 (N_18120,N_17966,N_17993);
xnor U18121 (N_18121,N_17729,N_17827);
and U18122 (N_18122,N_17820,N_17931);
nor U18123 (N_18123,N_17803,N_17703);
nor U18124 (N_18124,N_17869,N_17880);
or U18125 (N_18125,N_17850,N_17877);
nor U18126 (N_18126,N_17836,N_17706);
nand U18127 (N_18127,N_17870,N_17804);
or U18128 (N_18128,N_17714,N_17919);
nand U18129 (N_18129,N_17787,N_17782);
or U18130 (N_18130,N_17719,N_17784);
and U18131 (N_18131,N_17844,N_17948);
and U18132 (N_18132,N_17898,N_17705);
xor U18133 (N_18133,N_17810,N_17777);
nor U18134 (N_18134,N_17806,N_17796);
nand U18135 (N_18135,N_17961,N_17986);
nor U18136 (N_18136,N_17932,N_17814);
xor U18137 (N_18137,N_17916,N_17743);
or U18138 (N_18138,N_17910,N_17822);
nor U18139 (N_18139,N_17794,N_17776);
and U18140 (N_18140,N_17773,N_17783);
xor U18141 (N_18141,N_17947,N_17834);
nor U18142 (N_18142,N_17781,N_17829);
and U18143 (N_18143,N_17974,N_17854);
and U18144 (N_18144,N_17890,N_17921);
or U18145 (N_18145,N_17936,N_17897);
xnor U18146 (N_18146,N_17906,N_17984);
or U18147 (N_18147,N_17894,N_17976);
and U18148 (N_18148,N_17855,N_17918);
xnor U18149 (N_18149,N_17723,N_17742);
nand U18150 (N_18150,N_17987,N_17800);
or U18151 (N_18151,N_17786,N_17976);
and U18152 (N_18152,N_17754,N_17742);
and U18153 (N_18153,N_17718,N_17758);
or U18154 (N_18154,N_17760,N_17821);
nand U18155 (N_18155,N_17725,N_17860);
and U18156 (N_18156,N_17790,N_17972);
nand U18157 (N_18157,N_17888,N_17785);
nand U18158 (N_18158,N_17900,N_17789);
xor U18159 (N_18159,N_17991,N_17835);
nor U18160 (N_18160,N_17864,N_17881);
xnor U18161 (N_18161,N_17892,N_17880);
nor U18162 (N_18162,N_17940,N_17839);
or U18163 (N_18163,N_17760,N_17726);
nor U18164 (N_18164,N_17918,N_17994);
or U18165 (N_18165,N_17955,N_17757);
nand U18166 (N_18166,N_17999,N_17754);
or U18167 (N_18167,N_17918,N_17993);
or U18168 (N_18168,N_17772,N_17985);
nand U18169 (N_18169,N_17845,N_17911);
and U18170 (N_18170,N_17841,N_17866);
nand U18171 (N_18171,N_17809,N_17796);
xor U18172 (N_18172,N_17868,N_17889);
and U18173 (N_18173,N_17701,N_17734);
nand U18174 (N_18174,N_17717,N_17809);
nor U18175 (N_18175,N_17926,N_17823);
xnor U18176 (N_18176,N_17742,N_17982);
xor U18177 (N_18177,N_17788,N_17725);
xnor U18178 (N_18178,N_17914,N_17893);
nand U18179 (N_18179,N_17994,N_17851);
nand U18180 (N_18180,N_17977,N_17991);
xor U18181 (N_18181,N_17915,N_17832);
nor U18182 (N_18182,N_17857,N_17946);
xnor U18183 (N_18183,N_17748,N_17775);
and U18184 (N_18184,N_17736,N_17871);
nand U18185 (N_18185,N_17798,N_17976);
or U18186 (N_18186,N_17838,N_17817);
or U18187 (N_18187,N_17926,N_17922);
xnor U18188 (N_18188,N_17884,N_17715);
xor U18189 (N_18189,N_17889,N_17706);
nor U18190 (N_18190,N_17943,N_17896);
xor U18191 (N_18191,N_17916,N_17875);
or U18192 (N_18192,N_17888,N_17750);
nand U18193 (N_18193,N_17997,N_17822);
nor U18194 (N_18194,N_17845,N_17973);
nand U18195 (N_18195,N_17861,N_17785);
nor U18196 (N_18196,N_17808,N_17975);
nor U18197 (N_18197,N_17999,N_17912);
nand U18198 (N_18198,N_17947,N_17919);
nand U18199 (N_18199,N_17964,N_17922);
nand U18200 (N_18200,N_17843,N_17878);
and U18201 (N_18201,N_17993,N_17719);
nor U18202 (N_18202,N_17860,N_17772);
nand U18203 (N_18203,N_17770,N_17731);
nor U18204 (N_18204,N_17920,N_17827);
nor U18205 (N_18205,N_17844,N_17759);
or U18206 (N_18206,N_17929,N_17715);
or U18207 (N_18207,N_17944,N_17806);
and U18208 (N_18208,N_17817,N_17729);
xor U18209 (N_18209,N_17834,N_17733);
xnor U18210 (N_18210,N_17764,N_17746);
nand U18211 (N_18211,N_17771,N_17873);
nand U18212 (N_18212,N_17813,N_17833);
nor U18213 (N_18213,N_17959,N_17976);
and U18214 (N_18214,N_17999,N_17979);
nor U18215 (N_18215,N_17715,N_17887);
nand U18216 (N_18216,N_17763,N_17719);
xnor U18217 (N_18217,N_17968,N_17710);
nor U18218 (N_18218,N_17899,N_17794);
or U18219 (N_18219,N_17724,N_17931);
xnor U18220 (N_18220,N_17876,N_17727);
and U18221 (N_18221,N_17865,N_17863);
nand U18222 (N_18222,N_17856,N_17816);
xnor U18223 (N_18223,N_17741,N_17797);
nor U18224 (N_18224,N_17809,N_17815);
nor U18225 (N_18225,N_17794,N_17868);
xnor U18226 (N_18226,N_17950,N_17866);
xor U18227 (N_18227,N_17741,N_17859);
xor U18228 (N_18228,N_17701,N_17727);
xor U18229 (N_18229,N_17795,N_17836);
and U18230 (N_18230,N_17910,N_17950);
nor U18231 (N_18231,N_17933,N_17774);
or U18232 (N_18232,N_17892,N_17884);
or U18233 (N_18233,N_17703,N_17841);
or U18234 (N_18234,N_17960,N_17953);
nand U18235 (N_18235,N_17821,N_17994);
and U18236 (N_18236,N_17721,N_17789);
nor U18237 (N_18237,N_17793,N_17907);
nor U18238 (N_18238,N_17922,N_17823);
and U18239 (N_18239,N_17826,N_17908);
xnor U18240 (N_18240,N_17857,N_17789);
xor U18241 (N_18241,N_17875,N_17861);
nand U18242 (N_18242,N_17843,N_17773);
and U18243 (N_18243,N_17850,N_17732);
xor U18244 (N_18244,N_17791,N_17955);
and U18245 (N_18245,N_17786,N_17901);
or U18246 (N_18246,N_17823,N_17708);
and U18247 (N_18247,N_17915,N_17968);
nor U18248 (N_18248,N_17809,N_17928);
xnor U18249 (N_18249,N_17791,N_17822);
nand U18250 (N_18250,N_17837,N_17744);
xor U18251 (N_18251,N_17952,N_17899);
or U18252 (N_18252,N_17913,N_17799);
or U18253 (N_18253,N_17741,N_17928);
nor U18254 (N_18254,N_17740,N_17862);
or U18255 (N_18255,N_17905,N_17844);
xnor U18256 (N_18256,N_17869,N_17953);
nor U18257 (N_18257,N_17887,N_17895);
xor U18258 (N_18258,N_17799,N_17855);
nor U18259 (N_18259,N_17910,N_17732);
and U18260 (N_18260,N_17798,N_17830);
and U18261 (N_18261,N_17924,N_17897);
nand U18262 (N_18262,N_17720,N_17997);
and U18263 (N_18263,N_17936,N_17723);
and U18264 (N_18264,N_17912,N_17717);
nand U18265 (N_18265,N_17921,N_17768);
and U18266 (N_18266,N_17706,N_17926);
xnor U18267 (N_18267,N_17985,N_17757);
xnor U18268 (N_18268,N_17814,N_17820);
xnor U18269 (N_18269,N_17733,N_17758);
xor U18270 (N_18270,N_17773,N_17818);
xnor U18271 (N_18271,N_17834,N_17860);
or U18272 (N_18272,N_17948,N_17994);
and U18273 (N_18273,N_17866,N_17859);
nor U18274 (N_18274,N_17790,N_17943);
xor U18275 (N_18275,N_17892,N_17757);
xnor U18276 (N_18276,N_17863,N_17720);
xnor U18277 (N_18277,N_17872,N_17898);
nand U18278 (N_18278,N_17865,N_17883);
xnor U18279 (N_18279,N_17825,N_17937);
xor U18280 (N_18280,N_17842,N_17882);
or U18281 (N_18281,N_17861,N_17956);
and U18282 (N_18282,N_17817,N_17893);
nor U18283 (N_18283,N_17845,N_17883);
nand U18284 (N_18284,N_17747,N_17796);
or U18285 (N_18285,N_17861,N_17711);
or U18286 (N_18286,N_17882,N_17774);
and U18287 (N_18287,N_17863,N_17705);
xnor U18288 (N_18288,N_17929,N_17807);
or U18289 (N_18289,N_17717,N_17910);
nand U18290 (N_18290,N_17849,N_17738);
nand U18291 (N_18291,N_17724,N_17900);
and U18292 (N_18292,N_17879,N_17709);
or U18293 (N_18293,N_17968,N_17872);
and U18294 (N_18294,N_17977,N_17864);
and U18295 (N_18295,N_17808,N_17987);
nand U18296 (N_18296,N_17828,N_17852);
xnor U18297 (N_18297,N_17987,N_17957);
nand U18298 (N_18298,N_17981,N_17899);
or U18299 (N_18299,N_17887,N_17886);
and U18300 (N_18300,N_18063,N_18119);
and U18301 (N_18301,N_18281,N_18116);
xnor U18302 (N_18302,N_18088,N_18004);
or U18303 (N_18303,N_18047,N_18020);
nor U18304 (N_18304,N_18008,N_18220);
nor U18305 (N_18305,N_18169,N_18288);
nand U18306 (N_18306,N_18283,N_18298);
nor U18307 (N_18307,N_18135,N_18182);
xor U18308 (N_18308,N_18018,N_18037);
nand U18309 (N_18309,N_18231,N_18087);
and U18310 (N_18310,N_18214,N_18236);
or U18311 (N_18311,N_18096,N_18078);
or U18312 (N_18312,N_18093,N_18221);
nand U18313 (N_18313,N_18043,N_18068);
nand U18314 (N_18314,N_18145,N_18065);
and U18315 (N_18315,N_18164,N_18014);
xor U18316 (N_18316,N_18045,N_18155);
xor U18317 (N_18317,N_18051,N_18227);
and U18318 (N_18318,N_18044,N_18115);
nor U18319 (N_18319,N_18266,N_18090);
and U18320 (N_18320,N_18242,N_18059);
or U18321 (N_18321,N_18041,N_18027);
and U18322 (N_18322,N_18292,N_18091);
xnor U18323 (N_18323,N_18147,N_18042);
and U18324 (N_18324,N_18171,N_18212);
and U18325 (N_18325,N_18295,N_18028);
or U18326 (N_18326,N_18279,N_18204);
nand U18327 (N_18327,N_18112,N_18253);
or U18328 (N_18328,N_18262,N_18163);
or U18329 (N_18329,N_18180,N_18278);
xor U18330 (N_18330,N_18206,N_18124);
xor U18331 (N_18331,N_18229,N_18086);
nor U18332 (N_18332,N_18024,N_18218);
or U18333 (N_18333,N_18170,N_18114);
xnor U18334 (N_18334,N_18156,N_18141);
xnor U18335 (N_18335,N_18244,N_18261);
or U18336 (N_18336,N_18176,N_18174);
nor U18337 (N_18337,N_18021,N_18131);
and U18338 (N_18338,N_18210,N_18082);
and U18339 (N_18339,N_18293,N_18032);
xnor U18340 (N_18340,N_18194,N_18161);
and U18341 (N_18341,N_18255,N_18064);
or U18342 (N_18342,N_18069,N_18039);
and U18343 (N_18343,N_18187,N_18175);
and U18344 (N_18344,N_18201,N_18077);
xor U18345 (N_18345,N_18256,N_18005);
and U18346 (N_18346,N_18151,N_18002);
or U18347 (N_18347,N_18084,N_18081);
nand U18348 (N_18348,N_18061,N_18294);
nand U18349 (N_18349,N_18166,N_18085);
nand U18350 (N_18350,N_18132,N_18183);
nor U18351 (N_18351,N_18052,N_18209);
nor U18352 (N_18352,N_18033,N_18035);
nand U18353 (N_18353,N_18122,N_18172);
and U18354 (N_18354,N_18271,N_18006);
nand U18355 (N_18355,N_18127,N_18101);
or U18356 (N_18356,N_18029,N_18267);
nand U18357 (N_18357,N_18009,N_18275);
nand U18358 (N_18358,N_18226,N_18110);
xor U18359 (N_18359,N_18297,N_18259);
and U18360 (N_18360,N_18058,N_18282);
and U18361 (N_18361,N_18010,N_18067);
nor U18362 (N_18362,N_18017,N_18277);
and U18363 (N_18363,N_18079,N_18103);
nor U18364 (N_18364,N_18142,N_18143);
and U18365 (N_18365,N_18177,N_18076);
nor U18366 (N_18366,N_18191,N_18286);
nand U18367 (N_18367,N_18239,N_18159);
nand U18368 (N_18368,N_18246,N_18289);
nor U18369 (N_18369,N_18097,N_18276);
and U18370 (N_18370,N_18238,N_18034);
nand U18371 (N_18371,N_18038,N_18225);
nand U18372 (N_18372,N_18268,N_18046);
nand U18373 (N_18373,N_18228,N_18092);
nand U18374 (N_18374,N_18146,N_18126);
and U18375 (N_18375,N_18150,N_18152);
xor U18376 (N_18376,N_18190,N_18031);
nor U18377 (N_18377,N_18060,N_18181);
xor U18378 (N_18378,N_18269,N_18094);
nor U18379 (N_18379,N_18025,N_18036);
nor U18380 (N_18380,N_18184,N_18208);
or U18381 (N_18381,N_18066,N_18193);
nand U18382 (N_18382,N_18128,N_18049);
or U18383 (N_18383,N_18108,N_18178);
nor U18384 (N_18384,N_18284,N_18160);
nor U18385 (N_18385,N_18230,N_18167);
nor U18386 (N_18386,N_18280,N_18215);
and U18387 (N_18387,N_18012,N_18245);
nor U18388 (N_18388,N_18200,N_18264);
xnor U18389 (N_18389,N_18232,N_18107);
xnor U18390 (N_18390,N_18192,N_18057);
or U18391 (N_18391,N_18137,N_18140);
xnor U18392 (N_18392,N_18007,N_18083);
nand U18393 (N_18393,N_18123,N_18205);
nand U18394 (N_18394,N_18254,N_18075);
and U18395 (N_18395,N_18040,N_18179);
nor U18396 (N_18396,N_18168,N_18100);
nand U18397 (N_18397,N_18157,N_18257);
or U18398 (N_18398,N_18117,N_18023);
nand U18399 (N_18399,N_18197,N_18098);
nand U18400 (N_18400,N_18270,N_18149);
or U18401 (N_18401,N_18089,N_18048);
xnor U18402 (N_18402,N_18263,N_18173);
xnor U18403 (N_18403,N_18153,N_18016);
and U18404 (N_18404,N_18062,N_18055);
nor U18405 (N_18405,N_18189,N_18105);
nand U18406 (N_18406,N_18213,N_18195);
nor U18407 (N_18407,N_18241,N_18291);
and U18408 (N_18408,N_18134,N_18000);
nand U18409 (N_18409,N_18162,N_18222);
or U18410 (N_18410,N_18273,N_18249);
xnor U18411 (N_18411,N_18138,N_18247);
and U18412 (N_18412,N_18265,N_18074);
or U18413 (N_18413,N_18290,N_18274);
or U18414 (N_18414,N_18054,N_18251);
nand U18415 (N_18415,N_18158,N_18237);
nand U18416 (N_18416,N_18233,N_18113);
and U18417 (N_18417,N_18019,N_18154);
nor U18418 (N_18418,N_18186,N_18073);
and U18419 (N_18419,N_18219,N_18070);
or U18420 (N_18420,N_18248,N_18296);
or U18421 (N_18421,N_18080,N_18203);
nor U18422 (N_18422,N_18258,N_18260);
xnor U18423 (N_18423,N_18129,N_18243);
nand U18424 (N_18424,N_18050,N_18216);
xnor U18425 (N_18425,N_18196,N_18102);
nand U18426 (N_18426,N_18234,N_18011);
xnor U18427 (N_18427,N_18139,N_18056);
and U18428 (N_18428,N_18022,N_18003);
or U18429 (N_18429,N_18240,N_18285);
or U18430 (N_18430,N_18198,N_18133);
xor U18431 (N_18431,N_18111,N_18272);
xnor U18432 (N_18432,N_18207,N_18099);
and U18433 (N_18433,N_18252,N_18223);
nand U18434 (N_18434,N_18071,N_18121);
nand U18435 (N_18435,N_18120,N_18202);
nor U18436 (N_18436,N_18118,N_18217);
or U18437 (N_18437,N_18165,N_18235);
nor U18438 (N_18438,N_18125,N_18130);
nand U18439 (N_18439,N_18026,N_18013);
and U18440 (N_18440,N_18144,N_18072);
and U18441 (N_18441,N_18104,N_18106);
and U18442 (N_18442,N_18199,N_18015);
nor U18443 (N_18443,N_18224,N_18053);
or U18444 (N_18444,N_18109,N_18250);
or U18445 (N_18445,N_18188,N_18001);
or U18446 (N_18446,N_18299,N_18287);
nand U18447 (N_18447,N_18185,N_18030);
and U18448 (N_18448,N_18136,N_18095);
nand U18449 (N_18449,N_18148,N_18211);
nand U18450 (N_18450,N_18107,N_18187);
nor U18451 (N_18451,N_18287,N_18190);
nor U18452 (N_18452,N_18139,N_18112);
xor U18453 (N_18453,N_18296,N_18297);
or U18454 (N_18454,N_18254,N_18051);
nand U18455 (N_18455,N_18279,N_18070);
nand U18456 (N_18456,N_18090,N_18105);
nand U18457 (N_18457,N_18004,N_18107);
or U18458 (N_18458,N_18209,N_18249);
xor U18459 (N_18459,N_18230,N_18262);
xnor U18460 (N_18460,N_18257,N_18172);
xor U18461 (N_18461,N_18134,N_18069);
xor U18462 (N_18462,N_18095,N_18144);
xnor U18463 (N_18463,N_18029,N_18100);
and U18464 (N_18464,N_18126,N_18280);
or U18465 (N_18465,N_18038,N_18201);
nand U18466 (N_18466,N_18284,N_18013);
and U18467 (N_18467,N_18008,N_18038);
and U18468 (N_18468,N_18255,N_18017);
nand U18469 (N_18469,N_18048,N_18176);
nand U18470 (N_18470,N_18179,N_18256);
nand U18471 (N_18471,N_18225,N_18033);
nor U18472 (N_18472,N_18094,N_18104);
nor U18473 (N_18473,N_18097,N_18271);
nor U18474 (N_18474,N_18283,N_18184);
nor U18475 (N_18475,N_18064,N_18118);
or U18476 (N_18476,N_18031,N_18053);
nand U18477 (N_18477,N_18257,N_18208);
nand U18478 (N_18478,N_18239,N_18170);
nand U18479 (N_18479,N_18192,N_18260);
or U18480 (N_18480,N_18235,N_18033);
nand U18481 (N_18481,N_18108,N_18075);
nand U18482 (N_18482,N_18120,N_18165);
xor U18483 (N_18483,N_18258,N_18183);
xnor U18484 (N_18484,N_18167,N_18140);
and U18485 (N_18485,N_18215,N_18175);
xor U18486 (N_18486,N_18013,N_18227);
xnor U18487 (N_18487,N_18275,N_18238);
and U18488 (N_18488,N_18050,N_18266);
xor U18489 (N_18489,N_18299,N_18178);
xnor U18490 (N_18490,N_18051,N_18144);
and U18491 (N_18491,N_18053,N_18243);
nor U18492 (N_18492,N_18042,N_18205);
nor U18493 (N_18493,N_18275,N_18072);
nor U18494 (N_18494,N_18177,N_18102);
or U18495 (N_18495,N_18059,N_18198);
or U18496 (N_18496,N_18114,N_18184);
xor U18497 (N_18497,N_18115,N_18239);
or U18498 (N_18498,N_18151,N_18113);
or U18499 (N_18499,N_18052,N_18176);
nor U18500 (N_18500,N_18043,N_18096);
nor U18501 (N_18501,N_18265,N_18053);
nand U18502 (N_18502,N_18050,N_18273);
xor U18503 (N_18503,N_18116,N_18064);
nand U18504 (N_18504,N_18105,N_18260);
and U18505 (N_18505,N_18175,N_18221);
xnor U18506 (N_18506,N_18292,N_18259);
and U18507 (N_18507,N_18031,N_18104);
xnor U18508 (N_18508,N_18017,N_18231);
and U18509 (N_18509,N_18100,N_18265);
nor U18510 (N_18510,N_18250,N_18204);
and U18511 (N_18511,N_18016,N_18178);
nor U18512 (N_18512,N_18210,N_18061);
nand U18513 (N_18513,N_18138,N_18018);
nand U18514 (N_18514,N_18173,N_18132);
and U18515 (N_18515,N_18272,N_18064);
nand U18516 (N_18516,N_18269,N_18096);
xor U18517 (N_18517,N_18138,N_18244);
nor U18518 (N_18518,N_18201,N_18193);
or U18519 (N_18519,N_18099,N_18021);
xor U18520 (N_18520,N_18173,N_18117);
or U18521 (N_18521,N_18265,N_18021);
nand U18522 (N_18522,N_18268,N_18194);
or U18523 (N_18523,N_18189,N_18214);
or U18524 (N_18524,N_18220,N_18231);
xnor U18525 (N_18525,N_18209,N_18014);
nor U18526 (N_18526,N_18012,N_18171);
xor U18527 (N_18527,N_18207,N_18164);
xnor U18528 (N_18528,N_18253,N_18166);
nor U18529 (N_18529,N_18290,N_18037);
and U18530 (N_18530,N_18133,N_18203);
nor U18531 (N_18531,N_18162,N_18086);
xor U18532 (N_18532,N_18118,N_18199);
or U18533 (N_18533,N_18286,N_18009);
nor U18534 (N_18534,N_18051,N_18055);
xnor U18535 (N_18535,N_18290,N_18264);
and U18536 (N_18536,N_18271,N_18030);
xnor U18537 (N_18537,N_18130,N_18189);
nand U18538 (N_18538,N_18083,N_18233);
nand U18539 (N_18539,N_18031,N_18230);
nand U18540 (N_18540,N_18094,N_18274);
nand U18541 (N_18541,N_18192,N_18029);
nor U18542 (N_18542,N_18165,N_18119);
or U18543 (N_18543,N_18284,N_18188);
or U18544 (N_18544,N_18147,N_18139);
xor U18545 (N_18545,N_18133,N_18185);
nor U18546 (N_18546,N_18045,N_18255);
xnor U18547 (N_18547,N_18246,N_18269);
and U18548 (N_18548,N_18239,N_18099);
xnor U18549 (N_18549,N_18293,N_18250);
nor U18550 (N_18550,N_18032,N_18079);
xnor U18551 (N_18551,N_18062,N_18061);
xor U18552 (N_18552,N_18156,N_18008);
or U18553 (N_18553,N_18212,N_18252);
and U18554 (N_18554,N_18200,N_18128);
nand U18555 (N_18555,N_18013,N_18110);
nand U18556 (N_18556,N_18034,N_18289);
nor U18557 (N_18557,N_18003,N_18188);
xor U18558 (N_18558,N_18182,N_18160);
and U18559 (N_18559,N_18276,N_18020);
or U18560 (N_18560,N_18100,N_18077);
and U18561 (N_18561,N_18241,N_18124);
and U18562 (N_18562,N_18087,N_18234);
and U18563 (N_18563,N_18252,N_18288);
xor U18564 (N_18564,N_18119,N_18289);
and U18565 (N_18565,N_18202,N_18096);
or U18566 (N_18566,N_18119,N_18161);
xnor U18567 (N_18567,N_18059,N_18192);
or U18568 (N_18568,N_18045,N_18108);
nand U18569 (N_18569,N_18194,N_18059);
nand U18570 (N_18570,N_18078,N_18159);
nand U18571 (N_18571,N_18216,N_18155);
xor U18572 (N_18572,N_18069,N_18008);
nor U18573 (N_18573,N_18180,N_18027);
nor U18574 (N_18574,N_18248,N_18201);
xnor U18575 (N_18575,N_18082,N_18057);
or U18576 (N_18576,N_18160,N_18066);
and U18577 (N_18577,N_18049,N_18198);
or U18578 (N_18578,N_18069,N_18138);
or U18579 (N_18579,N_18198,N_18122);
nor U18580 (N_18580,N_18189,N_18050);
nand U18581 (N_18581,N_18109,N_18228);
and U18582 (N_18582,N_18228,N_18086);
nor U18583 (N_18583,N_18220,N_18109);
or U18584 (N_18584,N_18115,N_18205);
nor U18585 (N_18585,N_18140,N_18285);
and U18586 (N_18586,N_18035,N_18109);
or U18587 (N_18587,N_18020,N_18154);
nor U18588 (N_18588,N_18214,N_18139);
xor U18589 (N_18589,N_18012,N_18244);
xnor U18590 (N_18590,N_18292,N_18061);
nor U18591 (N_18591,N_18115,N_18149);
nor U18592 (N_18592,N_18186,N_18202);
and U18593 (N_18593,N_18208,N_18135);
nor U18594 (N_18594,N_18134,N_18171);
or U18595 (N_18595,N_18023,N_18179);
nand U18596 (N_18596,N_18150,N_18036);
nor U18597 (N_18597,N_18051,N_18259);
or U18598 (N_18598,N_18104,N_18243);
or U18599 (N_18599,N_18073,N_18001);
xor U18600 (N_18600,N_18316,N_18363);
or U18601 (N_18601,N_18460,N_18349);
and U18602 (N_18602,N_18525,N_18335);
nand U18603 (N_18603,N_18502,N_18497);
and U18604 (N_18604,N_18463,N_18441);
and U18605 (N_18605,N_18402,N_18478);
and U18606 (N_18606,N_18531,N_18545);
and U18607 (N_18607,N_18474,N_18374);
xor U18608 (N_18608,N_18354,N_18410);
xor U18609 (N_18609,N_18304,N_18309);
or U18610 (N_18610,N_18429,N_18358);
or U18611 (N_18611,N_18489,N_18526);
and U18612 (N_18612,N_18448,N_18428);
nor U18613 (N_18613,N_18574,N_18510);
nor U18614 (N_18614,N_18317,N_18416);
xnor U18615 (N_18615,N_18324,N_18303);
xnor U18616 (N_18616,N_18355,N_18342);
nand U18617 (N_18617,N_18369,N_18508);
and U18618 (N_18618,N_18313,N_18401);
nand U18619 (N_18619,N_18341,N_18507);
or U18620 (N_18620,N_18479,N_18403);
and U18621 (N_18621,N_18443,N_18315);
xnor U18622 (N_18622,N_18435,N_18327);
xor U18623 (N_18623,N_18565,N_18585);
nor U18624 (N_18624,N_18394,N_18576);
nor U18625 (N_18625,N_18559,N_18372);
and U18626 (N_18626,N_18509,N_18396);
nor U18627 (N_18627,N_18453,N_18382);
xnor U18628 (N_18628,N_18464,N_18530);
and U18629 (N_18629,N_18557,N_18541);
or U18630 (N_18630,N_18325,N_18424);
or U18631 (N_18631,N_18500,N_18570);
nor U18632 (N_18632,N_18482,N_18521);
nor U18633 (N_18633,N_18554,N_18381);
and U18634 (N_18634,N_18484,N_18498);
and U18635 (N_18635,N_18340,N_18377);
xnor U18636 (N_18636,N_18469,N_18449);
nand U18637 (N_18637,N_18346,N_18456);
and U18638 (N_18638,N_18450,N_18535);
nor U18639 (N_18639,N_18522,N_18433);
xor U18640 (N_18640,N_18584,N_18561);
nand U18641 (N_18641,N_18505,N_18552);
or U18642 (N_18642,N_18577,N_18551);
nand U18643 (N_18643,N_18527,N_18490);
nand U18644 (N_18644,N_18445,N_18312);
nand U18645 (N_18645,N_18417,N_18593);
nand U18646 (N_18646,N_18571,N_18459);
or U18647 (N_18647,N_18398,N_18553);
nand U18648 (N_18648,N_18431,N_18564);
or U18649 (N_18649,N_18386,N_18582);
nor U18650 (N_18650,N_18408,N_18462);
nor U18651 (N_18651,N_18421,N_18543);
or U18652 (N_18652,N_18523,N_18353);
nor U18653 (N_18653,N_18483,N_18359);
nand U18654 (N_18654,N_18400,N_18356);
xor U18655 (N_18655,N_18512,N_18332);
nand U18656 (N_18656,N_18536,N_18370);
xor U18657 (N_18657,N_18437,N_18520);
xnor U18658 (N_18658,N_18360,N_18348);
and U18659 (N_18659,N_18589,N_18391);
xnor U18660 (N_18660,N_18384,N_18580);
nand U18661 (N_18661,N_18393,N_18302);
and U18662 (N_18662,N_18555,N_18420);
nand U18663 (N_18663,N_18390,N_18501);
xor U18664 (N_18664,N_18307,N_18426);
and U18665 (N_18665,N_18319,N_18539);
and U18666 (N_18666,N_18488,N_18477);
nor U18667 (N_18667,N_18432,N_18563);
xor U18668 (N_18668,N_18533,N_18328);
or U18669 (N_18669,N_18331,N_18573);
nor U18670 (N_18670,N_18515,N_18493);
xor U18671 (N_18671,N_18430,N_18326);
and U18672 (N_18672,N_18440,N_18308);
nand U18673 (N_18673,N_18367,N_18486);
nor U18674 (N_18674,N_18376,N_18419);
and U18675 (N_18675,N_18562,N_18590);
xnor U18676 (N_18676,N_18494,N_18472);
nand U18677 (N_18677,N_18444,N_18364);
and U18678 (N_18678,N_18513,N_18537);
xor U18679 (N_18679,N_18528,N_18351);
or U18680 (N_18680,N_18339,N_18503);
xnor U18681 (N_18681,N_18454,N_18300);
nand U18682 (N_18682,N_18572,N_18379);
xor U18683 (N_18683,N_18540,N_18506);
nand U18684 (N_18684,N_18361,N_18547);
nor U18685 (N_18685,N_18495,N_18422);
nand U18686 (N_18686,N_18487,N_18392);
nor U18687 (N_18687,N_18597,N_18524);
or U18688 (N_18688,N_18399,N_18405);
nand U18689 (N_18689,N_18514,N_18314);
or U18690 (N_18690,N_18511,N_18544);
nor U18691 (N_18691,N_18362,N_18404);
xor U18692 (N_18692,N_18365,N_18587);
or U18693 (N_18693,N_18414,N_18334);
nor U18694 (N_18694,N_18436,N_18338);
xnor U18695 (N_18695,N_18442,N_18387);
nor U18696 (N_18696,N_18476,N_18546);
nand U18697 (N_18697,N_18594,N_18438);
and U18698 (N_18698,N_18468,N_18407);
xor U18699 (N_18699,N_18383,N_18470);
nor U18700 (N_18700,N_18485,N_18592);
nand U18701 (N_18701,N_18465,N_18491);
nand U18702 (N_18702,N_18447,N_18366);
and U18703 (N_18703,N_18534,N_18323);
xnor U18704 (N_18704,N_18578,N_18595);
xor U18705 (N_18705,N_18583,N_18415);
nand U18706 (N_18706,N_18467,N_18343);
nand U18707 (N_18707,N_18305,N_18591);
nor U18708 (N_18708,N_18344,N_18517);
xor U18709 (N_18709,N_18368,N_18588);
nand U18710 (N_18710,N_18519,N_18397);
or U18711 (N_18711,N_18466,N_18518);
and U18712 (N_18712,N_18598,N_18538);
nor U18713 (N_18713,N_18439,N_18542);
nand U18714 (N_18714,N_18318,N_18579);
and U18715 (N_18715,N_18333,N_18492);
nor U18716 (N_18716,N_18347,N_18395);
xnor U18717 (N_18717,N_18352,N_18499);
or U18718 (N_18718,N_18389,N_18306);
or U18719 (N_18719,N_18350,N_18418);
nand U18720 (N_18720,N_18457,N_18311);
or U18721 (N_18721,N_18452,N_18567);
nand U18722 (N_18722,N_18423,N_18337);
nand U18723 (N_18723,N_18461,N_18473);
xor U18724 (N_18724,N_18458,N_18480);
nand U18725 (N_18725,N_18301,N_18427);
or U18726 (N_18726,N_18569,N_18549);
nand U18727 (N_18727,N_18336,N_18586);
and U18728 (N_18728,N_18529,N_18596);
nand U18729 (N_18729,N_18550,N_18373);
nand U18730 (N_18730,N_18504,N_18475);
nand U18731 (N_18731,N_18471,N_18446);
nor U18732 (N_18732,N_18575,N_18556);
xor U18733 (N_18733,N_18345,N_18320);
nand U18734 (N_18734,N_18357,N_18378);
or U18735 (N_18735,N_18380,N_18560);
and U18736 (N_18736,N_18371,N_18329);
and U18737 (N_18737,N_18581,N_18322);
and U18738 (N_18738,N_18409,N_18310);
nor U18739 (N_18739,N_18411,N_18532);
xnor U18740 (N_18740,N_18330,N_18568);
and U18741 (N_18741,N_18375,N_18434);
nand U18742 (N_18742,N_18455,N_18406);
nand U18743 (N_18743,N_18516,N_18388);
nor U18744 (N_18744,N_18451,N_18496);
or U18745 (N_18745,N_18566,N_18599);
xor U18746 (N_18746,N_18412,N_18413);
and U18747 (N_18747,N_18425,N_18481);
or U18748 (N_18748,N_18385,N_18321);
and U18749 (N_18749,N_18548,N_18558);
nand U18750 (N_18750,N_18331,N_18481);
nor U18751 (N_18751,N_18328,N_18561);
nor U18752 (N_18752,N_18343,N_18395);
or U18753 (N_18753,N_18361,N_18331);
nand U18754 (N_18754,N_18511,N_18318);
or U18755 (N_18755,N_18529,N_18515);
xnor U18756 (N_18756,N_18523,N_18515);
or U18757 (N_18757,N_18441,N_18328);
nand U18758 (N_18758,N_18364,N_18356);
nor U18759 (N_18759,N_18490,N_18498);
nand U18760 (N_18760,N_18539,N_18588);
nor U18761 (N_18761,N_18302,N_18575);
and U18762 (N_18762,N_18320,N_18539);
or U18763 (N_18763,N_18588,N_18314);
nand U18764 (N_18764,N_18505,N_18431);
or U18765 (N_18765,N_18342,N_18480);
or U18766 (N_18766,N_18382,N_18362);
or U18767 (N_18767,N_18546,N_18470);
nand U18768 (N_18768,N_18392,N_18404);
or U18769 (N_18769,N_18476,N_18524);
or U18770 (N_18770,N_18335,N_18592);
nand U18771 (N_18771,N_18551,N_18492);
nand U18772 (N_18772,N_18590,N_18302);
xor U18773 (N_18773,N_18584,N_18386);
or U18774 (N_18774,N_18437,N_18518);
xor U18775 (N_18775,N_18345,N_18382);
and U18776 (N_18776,N_18395,N_18459);
xor U18777 (N_18777,N_18483,N_18487);
and U18778 (N_18778,N_18492,N_18401);
or U18779 (N_18779,N_18301,N_18546);
xnor U18780 (N_18780,N_18309,N_18333);
nand U18781 (N_18781,N_18314,N_18321);
nand U18782 (N_18782,N_18421,N_18532);
and U18783 (N_18783,N_18312,N_18431);
nand U18784 (N_18784,N_18453,N_18468);
nand U18785 (N_18785,N_18503,N_18561);
or U18786 (N_18786,N_18416,N_18387);
and U18787 (N_18787,N_18338,N_18316);
xor U18788 (N_18788,N_18454,N_18339);
and U18789 (N_18789,N_18581,N_18477);
xnor U18790 (N_18790,N_18555,N_18373);
nor U18791 (N_18791,N_18363,N_18460);
and U18792 (N_18792,N_18369,N_18407);
nand U18793 (N_18793,N_18450,N_18492);
nor U18794 (N_18794,N_18451,N_18574);
nor U18795 (N_18795,N_18309,N_18564);
xnor U18796 (N_18796,N_18300,N_18479);
nor U18797 (N_18797,N_18497,N_18397);
or U18798 (N_18798,N_18484,N_18517);
xor U18799 (N_18799,N_18346,N_18589);
or U18800 (N_18800,N_18591,N_18465);
or U18801 (N_18801,N_18523,N_18559);
nand U18802 (N_18802,N_18555,N_18406);
or U18803 (N_18803,N_18586,N_18315);
and U18804 (N_18804,N_18599,N_18314);
xor U18805 (N_18805,N_18332,N_18579);
xor U18806 (N_18806,N_18466,N_18485);
nand U18807 (N_18807,N_18435,N_18321);
nand U18808 (N_18808,N_18594,N_18598);
or U18809 (N_18809,N_18437,N_18423);
nor U18810 (N_18810,N_18327,N_18561);
xor U18811 (N_18811,N_18382,N_18366);
nand U18812 (N_18812,N_18465,N_18438);
and U18813 (N_18813,N_18370,N_18544);
and U18814 (N_18814,N_18506,N_18315);
xor U18815 (N_18815,N_18404,N_18397);
nand U18816 (N_18816,N_18305,N_18568);
or U18817 (N_18817,N_18439,N_18349);
or U18818 (N_18818,N_18498,N_18527);
xnor U18819 (N_18819,N_18424,N_18449);
nor U18820 (N_18820,N_18590,N_18452);
nor U18821 (N_18821,N_18463,N_18519);
or U18822 (N_18822,N_18354,N_18359);
or U18823 (N_18823,N_18457,N_18550);
and U18824 (N_18824,N_18524,N_18495);
or U18825 (N_18825,N_18434,N_18437);
or U18826 (N_18826,N_18420,N_18497);
nor U18827 (N_18827,N_18331,N_18492);
xor U18828 (N_18828,N_18528,N_18349);
or U18829 (N_18829,N_18507,N_18327);
or U18830 (N_18830,N_18403,N_18591);
xor U18831 (N_18831,N_18512,N_18340);
and U18832 (N_18832,N_18428,N_18372);
or U18833 (N_18833,N_18539,N_18337);
nand U18834 (N_18834,N_18595,N_18367);
or U18835 (N_18835,N_18591,N_18396);
xnor U18836 (N_18836,N_18479,N_18310);
nor U18837 (N_18837,N_18493,N_18301);
and U18838 (N_18838,N_18472,N_18522);
xor U18839 (N_18839,N_18385,N_18531);
xnor U18840 (N_18840,N_18477,N_18563);
nand U18841 (N_18841,N_18403,N_18400);
or U18842 (N_18842,N_18399,N_18504);
nor U18843 (N_18843,N_18408,N_18407);
and U18844 (N_18844,N_18571,N_18565);
xor U18845 (N_18845,N_18393,N_18459);
nor U18846 (N_18846,N_18544,N_18517);
nand U18847 (N_18847,N_18595,N_18546);
or U18848 (N_18848,N_18408,N_18581);
and U18849 (N_18849,N_18577,N_18531);
xor U18850 (N_18850,N_18432,N_18324);
nor U18851 (N_18851,N_18326,N_18559);
nor U18852 (N_18852,N_18547,N_18392);
nor U18853 (N_18853,N_18581,N_18454);
and U18854 (N_18854,N_18352,N_18342);
xnor U18855 (N_18855,N_18570,N_18483);
nand U18856 (N_18856,N_18371,N_18550);
nand U18857 (N_18857,N_18471,N_18559);
nor U18858 (N_18858,N_18398,N_18509);
nor U18859 (N_18859,N_18531,N_18521);
xnor U18860 (N_18860,N_18382,N_18494);
xor U18861 (N_18861,N_18386,N_18534);
and U18862 (N_18862,N_18372,N_18581);
xor U18863 (N_18863,N_18478,N_18506);
nand U18864 (N_18864,N_18563,N_18384);
and U18865 (N_18865,N_18463,N_18507);
or U18866 (N_18866,N_18596,N_18477);
or U18867 (N_18867,N_18565,N_18550);
xnor U18868 (N_18868,N_18321,N_18374);
xnor U18869 (N_18869,N_18397,N_18310);
nand U18870 (N_18870,N_18338,N_18405);
xor U18871 (N_18871,N_18560,N_18378);
nand U18872 (N_18872,N_18590,N_18381);
xnor U18873 (N_18873,N_18363,N_18573);
xnor U18874 (N_18874,N_18383,N_18392);
xor U18875 (N_18875,N_18575,N_18485);
xor U18876 (N_18876,N_18340,N_18396);
nor U18877 (N_18877,N_18336,N_18350);
and U18878 (N_18878,N_18476,N_18594);
xnor U18879 (N_18879,N_18399,N_18433);
or U18880 (N_18880,N_18338,N_18336);
or U18881 (N_18881,N_18544,N_18447);
xor U18882 (N_18882,N_18393,N_18525);
and U18883 (N_18883,N_18426,N_18436);
xnor U18884 (N_18884,N_18559,N_18528);
xnor U18885 (N_18885,N_18411,N_18443);
nand U18886 (N_18886,N_18447,N_18474);
xnor U18887 (N_18887,N_18463,N_18555);
nor U18888 (N_18888,N_18390,N_18325);
or U18889 (N_18889,N_18457,N_18325);
xnor U18890 (N_18890,N_18469,N_18381);
xor U18891 (N_18891,N_18429,N_18378);
xor U18892 (N_18892,N_18500,N_18558);
nand U18893 (N_18893,N_18540,N_18503);
xnor U18894 (N_18894,N_18588,N_18556);
and U18895 (N_18895,N_18591,N_18341);
nand U18896 (N_18896,N_18362,N_18457);
nor U18897 (N_18897,N_18452,N_18384);
or U18898 (N_18898,N_18454,N_18584);
xor U18899 (N_18899,N_18486,N_18415);
nor U18900 (N_18900,N_18678,N_18724);
nor U18901 (N_18901,N_18867,N_18838);
and U18902 (N_18902,N_18852,N_18812);
xor U18903 (N_18903,N_18839,N_18674);
or U18904 (N_18904,N_18794,N_18792);
or U18905 (N_18905,N_18788,N_18833);
nand U18906 (N_18906,N_18733,N_18649);
xnor U18907 (N_18907,N_18816,N_18662);
or U18908 (N_18908,N_18778,N_18661);
xor U18909 (N_18909,N_18784,N_18898);
and U18910 (N_18910,N_18738,N_18845);
or U18911 (N_18911,N_18817,N_18781);
xnor U18912 (N_18912,N_18896,N_18858);
and U18913 (N_18913,N_18883,N_18766);
nor U18914 (N_18914,N_18870,N_18657);
or U18915 (N_18915,N_18654,N_18653);
and U18916 (N_18916,N_18720,N_18861);
or U18917 (N_18917,N_18765,N_18634);
xor U18918 (N_18918,N_18630,N_18848);
or U18919 (N_18919,N_18892,N_18669);
nor U18920 (N_18920,N_18756,N_18632);
and U18921 (N_18921,N_18628,N_18686);
and U18922 (N_18922,N_18789,N_18715);
nor U18923 (N_18923,N_18783,N_18796);
nand U18924 (N_18924,N_18739,N_18605);
or U18925 (N_18925,N_18727,N_18790);
nand U18926 (N_18926,N_18735,N_18732);
and U18927 (N_18927,N_18606,N_18680);
xnor U18928 (N_18928,N_18889,N_18797);
or U18929 (N_18929,N_18785,N_18691);
nand U18930 (N_18930,N_18682,N_18846);
or U18931 (N_18931,N_18828,N_18791);
and U18932 (N_18932,N_18805,N_18762);
nor U18933 (N_18933,N_18659,N_18814);
or U18934 (N_18934,N_18882,N_18786);
and U18935 (N_18935,N_18642,N_18713);
nor U18936 (N_18936,N_18847,N_18744);
xnor U18937 (N_18937,N_18664,N_18800);
and U18938 (N_18938,N_18779,N_18831);
xor U18939 (N_18939,N_18868,N_18866);
or U18940 (N_18940,N_18830,N_18651);
and U18941 (N_18941,N_18853,N_18834);
and U18942 (N_18942,N_18712,N_18714);
or U18943 (N_18943,N_18660,N_18667);
or U18944 (N_18944,N_18887,N_18886);
or U18945 (N_18945,N_18769,N_18849);
xor U18946 (N_18946,N_18822,N_18730);
nor U18947 (N_18947,N_18695,N_18871);
nand U18948 (N_18948,N_18708,N_18857);
or U18949 (N_18949,N_18802,N_18641);
or U18950 (N_18950,N_18767,N_18742);
nand U18951 (N_18951,N_18676,N_18747);
nand U18952 (N_18952,N_18795,N_18803);
nor U18953 (N_18953,N_18754,N_18683);
or U18954 (N_18954,N_18780,N_18723);
nor U18955 (N_18955,N_18675,N_18635);
and U18956 (N_18956,N_18692,N_18821);
or U18957 (N_18957,N_18804,N_18772);
xor U18958 (N_18958,N_18865,N_18703);
xor U18959 (N_18959,N_18627,N_18824);
or U18960 (N_18960,N_18897,N_18699);
nor U18961 (N_18961,N_18652,N_18602);
and U18962 (N_18962,N_18891,N_18787);
xnor U18963 (N_18963,N_18726,N_18716);
and U18964 (N_18964,N_18601,N_18737);
or U18965 (N_18965,N_18644,N_18646);
nand U18966 (N_18966,N_18827,N_18707);
and U18967 (N_18967,N_18689,N_18687);
and U18968 (N_18968,N_18618,N_18837);
and U18969 (N_18969,N_18776,N_18679);
and U18970 (N_18970,N_18874,N_18709);
and U18971 (N_18971,N_18823,N_18734);
xor U18972 (N_18972,N_18607,N_18629);
or U18973 (N_18973,N_18684,N_18835);
or U18974 (N_18974,N_18806,N_18869);
nand U18975 (N_18975,N_18647,N_18843);
or U18976 (N_18976,N_18700,N_18899);
nor U18977 (N_18977,N_18878,N_18620);
or U18978 (N_18978,N_18836,N_18637);
xnor U18979 (N_18979,N_18609,N_18807);
nor U18980 (N_18980,N_18768,N_18877);
or U18981 (N_18981,N_18777,N_18633);
nor U18982 (N_18982,N_18740,N_18706);
and U18983 (N_18983,N_18728,N_18701);
xnor U18984 (N_18984,N_18622,N_18650);
and U18985 (N_18985,N_18656,N_18719);
xnor U18986 (N_18986,N_18743,N_18697);
or U18987 (N_18987,N_18617,N_18759);
or U18988 (N_18988,N_18610,N_18619);
nor U18989 (N_18989,N_18764,N_18844);
nor U18990 (N_18990,N_18614,N_18893);
and U18991 (N_18991,N_18808,N_18810);
nand U18992 (N_18992,N_18862,N_18611);
and U18993 (N_18993,N_18752,N_18748);
nand U18994 (N_18994,N_18639,N_18623);
or U18995 (N_18995,N_18826,N_18864);
and U18996 (N_18996,N_18895,N_18872);
or U18997 (N_18997,N_18655,N_18717);
nand U18998 (N_18998,N_18645,N_18888);
nand U18999 (N_18999,N_18718,N_18763);
nand U19000 (N_19000,N_18801,N_18859);
nor U19001 (N_19001,N_18850,N_18774);
nand U19002 (N_19002,N_18666,N_18636);
xnor U19003 (N_19003,N_18819,N_18825);
xor U19004 (N_19004,N_18782,N_18860);
xnor U19005 (N_19005,N_18670,N_18600);
nor U19006 (N_19006,N_18832,N_18885);
nand U19007 (N_19007,N_18829,N_18710);
nand U19008 (N_19008,N_18875,N_18881);
or U19009 (N_19009,N_18625,N_18751);
nand U19010 (N_19010,N_18705,N_18753);
xnor U19011 (N_19011,N_18879,N_18818);
or U19012 (N_19012,N_18638,N_18880);
and U19013 (N_19013,N_18729,N_18755);
and U19014 (N_19014,N_18722,N_18603);
nand U19015 (N_19015,N_18626,N_18631);
xnor U19016 (N_19016,N_18698,N_18770);
nand U19017 (N_19017,N_18604,N_18672);
xnor U19018 (N_19018,N_18761,N_18624);
nor U19019 (N_19019,N_18813,N_18685);
nand U19020 (N_19020,N_18890,N_18725);
or U19021 (N_19021,N_18757,N_18809);
nor U19022 (N_19022,N_18773,N_18736);
nand U19023 (N_19023,N_18894,N_18663);
nor U19024 (N_19024,N_18693,N_18677);
and U19025 (N_19025,N_18702,N_18690);
xnor U19026 (N_19026,N_18608,N_18615);
nand U19027 (N_19027,N_18671,N_18640);
xnor U19028 (N_19028,N_18820,N_18643);
nand U19029 (N_19029,N_18884,N_18731);
nor U19030 (N_19030,N_18793,N_18842);
nand U19031 (N_19031,N_18811,N_18851);
xor U19032 (N_19032,N_18749,N_18621);
xnor U19033 (N_19033,N_18721,N_18771);
or U19034 (N_19034,N_18758,N_18694);
and U19035 (N_19035,N_18798,N_18745);
or U19036 (N_19036,N_18799,N_18746);
or U19037 (N_19037,N_18863,N_18854);
nand U19038 (N_19038,N_18760,N_18815);
or U19039 (N_19039,N_18750,N_18775);
and U19040 (N_19040,N_18704,N_18696);
xnor U19041 (N_19041,N_18741,N_18711);
and U19042 (N_19042,N_18668,N_18841);
and U19043 (N_19043,N_18688,N_18665);
xnor U19044 (N_19044,N_18681,N_18613);
xnor U19045 (N_19045,N_18876,N_18840);
nor U19046 (N_19046,N_18616,N_18658);
nand U19047 (N_19047,N_18648,N_18612);
nor U19048 (N_19048,N_18855,N_18856);
and U19049 (N_19049,N_18873,N_18673);
nand U19050 (N_19050,N_18773,N_18667);
nand U19051 (N_19051,N_18730,N_18794);
nor U19052 (N_19052,N_18874,N_18879);
and U19053 (N_19053,N_18654,N_18726);
nand U19054 (N_19054,N_18634,N_18810);
and U19055 (N_19055,N_18683,N_18821);
nor U19056 (N_19056,N_18850,N_18727);
or U19057 (N_19057,N_18763,N_18670);
nand U19058 (N_19058,N_18759,N_18758);
nor U19059 (N_19059,N_18892,N_18779);
or U19060 (N_19060,N_18805,N_18838);
nand U19061 (N_19061,N_18757,N_18818);
nand U19062 (N_19062,N_18740,N_18853);
or U19063 (N_19063,N_18894,N_18776);
or U19064 (N_19064,N_18733,N_18830);
and U19065 (N_19065,N_18859,N_18811);
and U19066 (N_19066,N_18746,N_18602);
nor U19067 (N_19067,N_18795,N_18767);
nor U19068 (N_19068,N_18790,N_18869);
xnor U19069 (N_19069,N_18685,N_18846);
and U19070 (N_19070,N_18842,N_18877);
and U19071 (N_19071,N_18703,N_18646);
or U19072 (N_19072,N_18732,N_18605);
nand U19073 (N_19073,N_18770,N_18690);
nand U19074 (N_19074,N_18853,N_18616);
nand U19075 (N_19075,N_18722,N_18840);
and U19076 (N_19076,N_18737,N_18651);
or U19077 (N_19077,N_18886,N_18749);
nand U19078 (N_19078,N_18891,N_18880);
nand U19079 (N_19079,N_18765,N_18660);
and U19080 (N_19080,N_18744,N_18821);
or U19081 (N_19081,N_18652,N_18841);
nor U19082 (N_19082,N_18788,N_18727);
nor U19083 (N_19083,N_18836,N_18806);
or U19084 (N_19084,N_18757,N_18863);
and U19085 (N_19085,N_18675,N_18773);
nand U19086 (N_19086,N_18797,N_18839);
and U19087 (N_19087,N_18784,N_18831);
nand U19088 (N_19088,N_18836,N_18659);
nand U19089 (N_19089,N_18615,N_18879);
nor U19090 (N_19090,N_18607,N_18706);
nand U19091 (N_19091,N_18887,N_18605);
or U19092 (N_19092,N_18674,N_18616);
nor U19093 (N_19093,N_18837,N_18643);
and U19094 (N_19094,N_18833,N_18720);
nand U19095 (N_19095,N_18601,N_18603);
or U19096 (N_19096,N_18720,N_18893);
nand U19097 (N_19097,N_18766,N_18615);
and U19098 (N_19098,N_18617,N_18895);
nand U19099 (N_19099,N_18681,N_18648);
or U19100 (N_19100,N_18845,N_18691);
and U19101 (N_19101,N_18694,N_18719);
nor U19102 (N_19102,N_18802,N_18678);
nor U19103 (N_19103,N_18702,N_18663);
nor U19104 (N_19104,N_18616,N_18785);
or U19105 (N_19105,N_18613,N_18639);
or U19106 (N_19106,N_18650,N_18831);
and U19107 (N_19107,N_18617,N_18801);
or U19108 (N_19108,N_18854,N_18828);
nor U19109 (N_19109,N_18688,N_18779);
or U19110 (N_19110,N_18612,N_18762);
nand U19111 (N_19111,N_18611,N_18828);
xor U19112 (N_19112,N_18862,N_18787);
or U19113 (N_19113,N_18843,N_18796);
or U19114 (N_19114,N_18759,N_18839);
or U19115 (N_19115,N_18632,N_18611);
nor U19116 (N_19116,N_18637,N_18862);
xnor U19117 (N_19117,N_18621,N_18894);
xor U19118 (N_19118,N_18772,N_18767);
xor U19119 (N_19119,N_18637,N_18627);
nor U19120 (N_19120,N_18698,N_18785);
nor U19121 (N_19121,N_18680,N_18724);
or U19122 (N_19122,N_18616,N_18626);
nor U19123 (N_19123,N_18731,N_18721);
nor U19124 (N_19124,N_18631,N_18806);
or U19125 (N_19125,N_18753,N_18678);
nand U19126 (N_19126,N_18757,N_18647);
nand U19127 (N_19127,N_18614,N_18627);
and U19128 (N_19128,N_18837,N_18689);
and U19129 (N_19129,N_18825,N_18802);
and U19130 (N_19130,N_18702,N_18736);
or U19131 (N_19131,N_18720,N_18892);
nand U19132 (N_19132,N_18638,N_18871);
xor U19133 (N_19133,N_18637,N_18640);
xor U19134 (N_19134,N_18896,N_18849);
or U19135 (N_19135,N_18747,N_18855);
and U19136 (N_19136,N_18724,N_18715);
nor U19137 (N_19137,N_18883,N_18807);
xor U19138 (N_19138,N_18608,N_18604);
nor U19139 (N_19139,N_18840,N_18609);
nand U19140 (N_19140,N_18836,N_18634);
or U19141 (N_19141,N_18770,N_18749);
or U19142 (N_19142,N_18899,N_18618);
nand U19143 (N_19143,N_18633,N_18844);
or U19144 (N_19144,N_18850,N_18690);
xnor U19145 (N_19145,N_18698,N_18875);
xor U19146 (N_19146,N_18702,N_18885);
nor U19147 (N_19147,N_18831,N_18620);
or U19148 (N_19148,N_18788,N_18784);
and U19149 (N_19149,N_18705,N_18765);
nor U19150 (N_19150,N_18875,N_18729);
nor U19151 (N_19151,N_18799,N_18650);
nor U19152 (N_19152,N_18697,N_18764);
xor U19153 (N_19153,N_18820,N_18649);
nand U19154 (N_19154,N_18806,N_18720);
and U19155 (N_19155,N_18748,N_18713);
or U19156 (N_19156,N_18760,N_18717);
nor U19157 (N_19157,N_18891,N_18615);
nand U19158 (N_19158,N_18800,N_18881);
or U19159 (N_19159,N_18668,N_18813);
nor U19160 (N_19160,N_18633,N_18634);
nand U19161 (N_19161,N_18858,N_18742);
xnor U19162 (N_19162,N_18731,N_18655);
nor U19163 (N_19163,N_18696,N_18814);
and U19164 (N_19164,N_18681,N_18852);
nand U19165 (N_19165,N_18774,N_18867);
and U19166 (N_19166,N_18801,N_18635);
xor U19167 (N_19167,N_18786,N_18691);
or U19168 (N_19168,N_18886,N_18629);
xor U19169 (N_19169,N_18602,N_18645);
nand U19170 (N_19170,N_18728,N_18757);
nor U19171 (N_19171,N_18763,N_18745);
nor U19172 (N_19172,N_18702,N_18617);
nor U19173 (N_19173,N_18826,N_18806);
nor U19174 (N_19174,N_18643,N_18845);
and U19175 (N_19175,N_18733,N_18795);
nor U19176 (N_19176,N_18690,N_18667);
or U19177 (N_19177,N_18706,N_18846);
xnor U19178 (N_19178,N_18693,N_18718);
and U19179 (N_19179,N_18678,N_18609);
nor U19180 (N_19180,N_18822,N_18706);
nor U19181 (N_19181,N_18692,N_18881);
and U19182 (N_19182,N_18847,N_18849);
nor U19183 (N_19183,N_18835,N_18848);
nor U19184 (N_19184,N_18874,N_18824);
nor U19185 (N_19185,N_18819,N_18749);
or U19186 (N_19186,N_18706,N_18785);
xnor U19187 (N_19187,N_18612,N_18735);
xor U19188 (N_19188,N_18802,N_18807);
xnor U19189 (N_19189,N_18643,N_18685);
nand U19190 (N_19190,N_18695,N_18800);
nand U19191 (N_19191,N_18667,N_18772);
nand U19192 (N_19192,N_18897,N_18645);
nor U19193 (N_19193,N_18696,N_18748);
xnor U19194 (N_19194,N_18682,N_18819);
nor U19195 (N_19195,N_18830,N_18711);
nand U19196 (N_19196,N_18822,N_18679);
or U19197 (N_19197,N_18728,N_18655);
xor U19198 (N_19198,N_18790,N_18697);
or U19199 (N_19199,N_18736,N_18857);
and U19200 (N_19200,N_19088,N_19086);
nand U19201 (N_19201,N_18948,N_18934);
nor U19202 (N_19202,N_18972,N_18973);
and U19203 (N_19203,N_19112,N_19055);
xnor U19204 (N_19204,N_19113,N_19105);
nor U19205 (N_19205,N_18927,N_18946);
nor U19206 (N_19206,N_19017,N_19035);
and U19207 (N_19207,N_18904,N_18908);
xnor U19208 (N_19208,N_19102,N_19019);
xor U19209 (N_19209,N_19126,N_18903);
nor U19210 (N_19210,N_18937,N_19183);
xor U19211 (N_19211,N_19106,N_18906);
and U19212 (N_19212,N_18967,N_18993);
and U19213 (N_19213,N_19178,N_18975);
and U19214 (N_19214,N_19038,N_18901);
or U19215 (N_19215,N_19002,N_19018);
nand U19216 (N_19216,N_19152,N_18965);
or U19217 (N_19217,N_19172,N_19093);
nand U19218 (N_19218,N_18925,N_19137);
xnor U19219 (N_19219,N_19171,N_18947);
nor U19220 (N_19220,N_19039,N_19095);
nand U19221 (N_19221,N_19162,N_19164);
nor U19222 (N_19222,N_19087,N_19057);
and U19223 (N_19223,N_19129,N_18938);
nand U19224 (N_19224,N_19060,N_18952);
nand U19225 (N_19225,N_18987,N_19121);
or U19226 (N_19226,N_18998,N_18914);
nand U19227 (N_19227,N_19101,N_19096);
xor U19228 (N_19228,N_18910,N_18961);
nand U19229 (N_19229,N_19177,N_18942);
or U19230 (N_19230,N_19168,N_19193);
nand U19231 (N_19231,N_19157,N_19160);
nor U19232 (N_19232,N_19056,N_19027);
xnor U19233 (N_19233,N_19196,N_19182);
nand U19234 (N_19234,N_19098,N_19179);
nor U19235 (N_19235,N_19170,N_18939);
nor U19236 (N_19236,N_19081,N_19030);
nand U19237 (N_19237,N_19007,N_19051);
xor U19238 (N_19238,N_18926,N_18979);
xnor U19239 (N_19239,N_19180,N_19189);
or U19240 (N_19240,N_18913,N_19117);
xnor U19241 (N_19241,N_18922,N_18940);
nor U19242 (N_19242,N_19050,N_18988);
nor U19243 (N_19243,N_19003,N_19071);
nand U19244 (N_19244,N_19059,N_19166);
nand U19245 (N_19245,N_18983,N_19009);
nand U19246 (N_19246,N_19042,N_19010);
nor U19247 (N_19247,N_19135,N_19076);
and U19248 (N_19248,N_19174,N_19120);
or U19249 (N_19249,N_19012,N_19001);
or U19250 (N_19250,N_18981,N_18918);
nor U19251 (N_19251,N_19107,N_19130);
and U19252 (N_19252,N_18955,N_19029);
nor U19253 (N_19253,N_19058,N_19141);
nand U19254 (N_19254,N_19147,N_19192);
or U19255 (N_19255,N_19125,N_19099);
or U19256 (N_19256,N_18936,N_19104);
or U19257 (N_19257,N_19014,N_18909);
or U19258 (N_19258,N_19085,N_19070);
nand U19259 (N_19259,N_19115,N_19063);
nand U19260 (N_19260,N_19084,N_19143);
xnor U19261 (N_19261,N_18985,N_18977);
nand U19262 (N_19262,N_19127,N_19199);
nand U19263 (N_19263,N_19025,N_18976);
or U19264 (N_19264,N_19068,N_19080);
nor U19265 (N_19265,N_19048,N_19054);
and U19266 (N_19266,N_18917,N_19142);
and U19267 (N_19267,N_19184,N_18902);
and U19268 (N_19268,N_18916,N_19067);
and U19269 (N_19269,N_18912,N_18905);
nand U19270 (N_19270,N_18989,N_19026);
xnor U19271 (N_19271,N_18941,N_19065);
nor U19272 (N_19272,N_19069,N_19116);
nand U19273 (N_19273,N_19198,N_19092);
and U19274 (N_19274,N_19140,N_19124);
xnor U19275 (N_19275,N_19109,N_19153);
and U19276 (N_19276,N_18968,N_19008);
nand U19277 (N_19277,N_18944,N_19165);
nor U19278 (N_19278,N_19016,N_19138);
and U19279 (N_19279,N_19064,N_18969);
nor U19280 (N_19280,N_18931,N_19190);
and U19281 (N_19281,N_18954,N_19074);
nand U19282 (N_19282,N_19072,N_19191);
and U19283 (N_19283,N_18970,N_19062);
and U19284 (N_19284,N_18929,N_19024);
nand U19285 (N_19285,N_18984,N_19132);
nor U19286 (N_19286,N_18924,N_19197);
xnor U19287 (N_19287,N_19046,N_19036);
nor U19288 (N_19288,N_18978,N_19006);
nand U19289 (N_19289,N_18900,N_19015);
nand U19290 (N_19290,N_19149,N_19134);
or U19291 (N_19291,N_18957,N_19128);
nor U19292 (N_19292,N_19167,N_19195);
xor U19293 (N_19293,N_18960,N_19021);
and U19294 (N_19294,N_18921,N_19169);
and U19295 (N_19295,N_19052,N_19108);
nand U19296 (N_19296,N_19151,N_18992);
and U19297 (N_19297,N_19122,N_19011);
nor U19298 (N_19298,N_18966,N_19161);
nand U19299 (N_19299,N_19049,N_18991);
nor U19300 (N_19300,N_19022,N_19020);
or U19301 (N_19301,N_18953,N_18920);
and U19302 (N_19302,N_18951,N_19158);
and U19303 (N_19303,N_19145,N_19186);
nand U19304 (N_19304,N_19139,N_18945);
and U19305 (N_19305,N_19045,N_18911);
nand U19306 (N_19306,N_19110,N_18950);
xor U19307 (N_19307,N_19041,N_19004);
and U19308 (N_19308,N_18932,N_19023);
nor U19309 (N_19309,N_19073,N_19078);
xnor U19310 (N_19310,N_18962,N_19123);
xnor U19311 (N_19311,N_19148,N_19032);
xor U19312 (N_19312,N_19188,N_19097);
or U19313 (N_19313,N_19103,N_19118);
or U19314 (N_19314,N_19159,N_19176);
xor U19315 (N_19315,N_19082,N_19083);
nor U19316 (N_19316,N_19044,N_19146);
nand U19317 (N_19317,N_19131,N_18915);
nand U19318 (N_19318,N_19136,N_19005);
or U19319 (N_19319,N_18919,N_19034);
nor U19320 (N_19320,N_19079,N_18996);
and U19321 (N_19321,N_18980,N_19077);
and U19322 (N_19322,N_18935,N_18907);
and U19323 (N_19323,N_18933,N_18923);
nand U19324 (N_19324,N_19163,N_19040);
nand U19325 (N_19325,N_19111,N_18964);
nor U19326 (N_19326,N_19119,N_19053);
and U19327 (N_19327,N_19091,N_19144);
nand U19328 (N_19328,N_19075,N_19181);
xnor U19329 (N_19329,N_19033,N_19175);
nor U19330 (N_19330,N_19013,N_18958);
nor U19331 (N_19331,N_18959,N_19185);
or U19332 (N_19332,N_19155,N_19089);
nor U19333 (N_19333,N_18994,N_18997);
and U19334 (N_19334,N_18928,N_19133);
nand U19335 (N_19335,N_19114,N_19194);
nor U19336 (N_19336,N_18963,N_19150);
or U19337 (N_19337,N_19090,N_18995);
and U19338 (N_19338,N_19043,N_18986);
and U19339 (N_19339,N_18949,N_18943);
nor U19340 (N_19340,N_19047,N_19031);
xnor U19341 (N_19341,N_18971,N_19173);
nand U19342 (N_19342,N_19100,N_19187);
and U19343 (N_19343,N_19037,N_19061);
nor U19344 (N_19344,N_18974,N_18982);
nand U19345 (N_19345,N_18990,N_19156);
and U19346 (N_19346,N_19028,N_18930);
nand U19347 (N_19347,N_19066,N_18999);
and U19348 (N_19348,N_19094,N_19154);
xor U19349 (N_19349,N_19000,N_18956);
or U19350 (N_19350,N_19045,N_19042);
nor U19351 (N_19351,N_19023,N_18916);
or U19352 (N_19352,N_19082,N_19120);
and U19353 (N_19353,N_18959,N_18923);
and U19354 (N_19354,N_19190,N_18924);
xnor U19355 (N_19355,N_18958,N_19120);
xnor U19356 (N_19356,N_19056,N_19009);
or U19357 (N_19357,N_19060,N_18962);
nor U19358 (N_19358,N_19078,N_19085);
xor U19359 (N_19359,N_19125,N_19145);
xnor U19360 (N_19360,N_19103,N_18995);
nand U19361 (N_19361,N_19079,N_19160);
nor U19362 (N_19362,N_19018,N_18972);
nor U19363 (N_19363,N_19085,N_19089);
or U19364 (N_19364,N_19052,N_19100);
and U19365 (N_19365,N_19061,N_19189);
or U19366 (N_19366,N_19085,N_19054);
nor U19367 (N_19367,N_19047,N_18944);
xor U19368 (N_19368,N_19159,N_18952);
and U19369 (N_19369,N_18952,N_19040);
nand U19370 (N_19370,N_18990,N_18984);
nand U19371 (N_19371,N_18972,N_19154);
or U19372 (N_19372,N_19108,N_18990);
xor U19373 (N_19373,N_19025,N_19153);
xor U19374 (N_19374,N_18957,N_19069);
or U19375 (N_19375,N_18933,N_19088);
and U19376 (N_19376,N_19002,N_18976);
nor U19377 (N_19377,N_19076,N_18947);
nand U19378 (N_19378,N_19067,N_19188);
and U19379 (N_19379,N_18931,N_18932);
or U19380 (N_19380,N_19134,N_19100);
nor U19381 (N_19381,N_19091,N_18950);
or U19382 (N_19382,N_18928,N_19005);
and U19383 (N_19383,N_19018,N_19146);
nor U19384 (N_19384,N_19071,N_19177);
and U19385 (N_19385,N_18910,N_19160);
nand U19386 (N_19386,N_18969,N_19046);
nor U19387 (N_19387,N_19025,N_18961);
nor U19388 (N_19388,N_18972,N_18989);
or U19389 (N_19389,N_18953,N_18963);
or U19390 (N_19390,N_18955,N_19159);
nor U19391 (N_19391,N_18983,N_19115);
xor U19392 (N_19392,N_18914,N_19063);
xnor U19393 (N_19393,N_18947,N_19050);
and U19394 (N_19394,N_19024,N_19193);
nor U19395 (N_19395,N_19136,N_19054);
xor U19396 (N_19396,N_18953,N_18947);
xnor U19397 (N_19397,N_19063,N_19107);
and U19398 (N_19398,N_19070,N_19056);
and U19399 (N_19399,N_19020,N_19149);
xor U19400 (N_19400,N_19156,N_18937);
nand U19401 (N_19401,N_18972,N_18988);
xor U19402 (N_19402,N_19133,N_19016);
or U19403 (N_19403,N_19124,N_19127);
or U19404 (N_19404,N_19063,N_18928);
nor U19405 (N_19405,N_18962,N_18983);
or U19406 (N_19406,N_19021,N_18917);
xnor U19407 (N_19407,N_18966,N_19148);
xnor U19408 (N_19408,N_19100,N_19137);
nor U19409 (N_19409,N_19116,N_19097);
and U19410 (N_19410,N_18938,N_19157);
or U19411 (N_19411,N_19132,N_19003);
and U19412 (N_19412,N_19007,N_18957);
and U19413 (N_19413,N_19176,N_19023);
or U19414 (N_19414,N_18906,N_18966);
nand U19415 (N_19415,N_18961,N_19038);
and U19416 (N_19416,N_18910,N_19056);
nand U19417 (N_19417,N_18954,N_19131);
or U19418 (N_19418,N_19083,N_19053);
nand U19419 (N_19419,N_19025,N_19084);
and U19420 (N_19420,N_18986,N_18980);
xor U19421 (N_19421,N_19080,N_19071);
nor U19422 (N_19422,N_19174,N_19029);
and U19423 (N_19423,N_19048,N_18933);
xnor U19424 (N_19424,N_19111,N_19054);
and U19425 (N_19425,N_19067,N_19084);
xnor U19426 (N_19426,N_19024,N_19004);
and U19427 (N_19427,N_19019,N_19097);
or U19428 (N_19428,N_19094,N_19052);
xnor U19429 (N_19429,N_18979,N_18960);
xnor U19430 (N_19430,N_18957,N_18905);
or U19431 (N_19431,N_18977,N_19015);
nand U19432 (N_19432,N_19020,N_19099);
or U19433 (N_19433,N_19135,N_18992);
xnor U19434 (N_19434,N_19042,N_19118);
nand U19435 (N_19435,N_18949,N_19065);
nand U19436 (N_19436,N_19003,N_19018);
and U19437 (N_19437,N_18922,N_19134);
xor U19438 (N_19438,N_19059,N_19002);
nor U19439 (N_19439,N_19039,N_18984);
nand U19440 (N_19440,N_19129,N_19010);
nor U19441 (N_19441,N_19059,N_19019);
xnor U19442 (N_19442,N_18931,N_19157);
nand U19443 (N_19443,N_19003,N_19145);
or U19444 (N_19444,N_19071,N_19199);
xnor U19445 (N_19445,N_18929,N_18964);
nor U19446 (N_19446,N_18970,N_19148);
nand U19447 (N_19447,N_18984,N_19090);
nor U19448 (N_19448,N_19192,N_18941);
xor U19449 (N_19449,N_19077,N_18953);
nand U19450 (N_19450,N_19136,N_18903);
nand U19451 (N_19451,N_19115,N_19073);
or U19452 (N_19452,N_19183,N_19016);
xnor U19453 (N_19453,N_19049,N_18963);
nor U19454 (N_19454,N_19121,N_19047);
nor U19455 (N_19455,N_18952,N_18992);
or U19456 (N_19456,N_19020,N_18945);
nor U19457 (N_19457,N_18970,N_19100);
nor U19458 (N_19458,N_19037,N_19041);
or U19459 (N_19459,N_18989,N_19148);
and U19460 (N_19460,N_19073,N_19131);
or U19461 (N_19461,N_19029,N_19034);
or U19462 (N_19462,N_18947,N_19194);
xnor U19463 (N_19463,N_19132,N_18910);
nor U19464 (N_19464,N_18923,N_19063);
nor U19465 (N_19465,N_19044,N_19196);
nor U19466 (N_19466,N_18936,N_19002);
and U19467 (N_19467,N_19007,N_18984);
and U19468 (N_19468,N_19029,N_19181);
xnor U19469 (N_19469,N_19021,N_19040);
nor U19470 (N_19470,N_18988,N_19175);
and U19471 (N_19471,N_18918,N_18901);
nand U19472 (N_19472,N_18984,N_19197);
xor U19473 (N_19473,N_19001,N_19033);
or U19474 (N_19474,N_19025,N_19049);
and U19475 (N_19475,N_19177,N_19135);
nor U19476 (N_19476,N_19058,N_18901);
xnor U19477 (N_19477,N_19075,N_18956);
and U19478 (N_19478,N_19014,N_19041);
nor U19479 (N_19479,N_18942,N_19042);
nand U19480 (N_19480,N_18901,N_19193);
nor U19481 (N_19481,N_19172,N_19098);
nor U19482 (N_19482,N_19071,N_18983);
or U19483 (N_19483,N_18926,N_19039);
or U19484 (N_19484,N_18921,N_19136);
xnor U19485 (N_19485,N_19177,N_19167);
and U19486 (N_19486,N_19167,N_18934);
and U19487 (N_19487,N_19105,N_18915);
nand U19488 (N_19488,N_18921,N_18927);
nor U19489 (N_19489,N_19063,N_18980);
nor U19490 (N_19490,N_19061,N_18912);
nand U19491 (N_19491,N_19134,N_19076);
nand U19492 (N_19492,N_19158,N_19112);
nand U19493 (N_19493,N_19160,N_19048);
and U19494 (N_19494,N_19090,N_19146);
or U19495 (N_19495,N_18972,N_18920);
xnor U19496 (N_19496,N_19111,N_18928);
nand U19497 (N_19497,N_18975,N_19017);
and U19498 (N_19498,N_19124,N_19031);
nand U19499 (N_19499,N_19134,N_19019);
nor U19500 (N_19500,N_19381,N_19429);
nor U19501 (N_19501,N_19318,N_19263);
and U19502 (N_19502,N_19360,N_19350);
xor U19503 (N_19503,N_19416,N_19316);
or U19504 (N_19504,N_19465,N_19309);
nand U19505 (N_19505,N_19365,N_19414);
or U19506 (N_19506,N_19262,N_19255);
xnor U19507 (N_19507,N_19479,N_19388);
and U19508 (N_19508,N_19389,N_19302);
and U19509 (N_19509,N_19272,N_19346);
nor U19510 (N_19510,N_19203,N_19433);
xor U19511 (N_19511,N_19271,N_19415);
or U19512 (N_19512,N_19292,N_19289);
nor U19513 (N_19513,N_19205,N_19482);
nand U19514 (N_19514,N_19361,N_19435);
and U19515 (N_19515,N_19495,N_19339);
nand U19516 (N_19516,N_19457,N_19370);
and U19517 (N_19517,N_19234,N_19215);
nand U19518 (N_19518,N_19296,N_19440);
nor U19519 (N_19519,N_19409,N_19397);
or U19520 (N_19520,N_19474,N_19281);
and U19521 (N_19521,N_19209,N_19400);
nand U19522 (N_19522,N_19250,N_19471);
or U19523 (N_19523,N_19320,N_19453);
xnor U19524 (N_19524,N_19357,N_19264);
or U19525 (N_19525,N_19385,N_19458);
or U19526 (N_19526,N_19244,N_19488);
xor U19527 (N_19527,N_19448,N_19493);
xor U19528 (N_19528,N_19232,N_19403);
nor U19529 (N_19529,N_19386,N_19268);
and U19530 (N_19530,N_19283,N_19480);
and U19531 (N_19531,N_19329,N_19475);
or U19532 (N_19532,N_19221,N_19413);
and U19533 (N_19533,N_19254,N_19379);
xnor U19534 (N_19534,N_19301,N_19242);
nand U19535 (N_19535,N_19477,N_19432);
or U19536 (N_19536,N_19390,N_19355);
nor U19537 (N_19537,N_19472,N_19417);
xnor U19538 (N_19538,N_19335,N_19330);
xnor U19539 (N_19539,N_19406,N_19280);
and U19540 (N_19540,N_19491,N_19277);
or U19541 (N_19541,N_19362,N_19208);
and U19542 (N_19542,N_19229,N_19438);
nor U19543 (N_19543,N_19384,N_19241);
and U19544 (N_19544,N_19430,N_19497);
and U19545 (N_19545,N_19315,N_19455);
xor U19546 (N_19546,N_19256,N_19291);
nor U19547 (N_19547,N_19233,N_19434);
nand U19548 (N_19548,N_19359,N_19286);
nand U19549 (N_19549,N_19237,N_19352);
nand U19550 (N_19550,N_19240,N_19211);
xor U19551 (N_19551,N_19421,N_19344);
and U19552 (N_19552,N_19285,N_19260);
and U19553 (N_19553,N_19239,N_19425);
nand U19554 (N_19554,N_19424,N_19396);
and U19555 (N_19555,N_19478,N_19319);
and U19556 (N_19556,N_19227,N_19364);
nand U19557 (N_19557,N_19265,N_19368);
xor U19558 (N_19558,N_19243,N_19444);
and U19559 (N_19559,N_19249,N_19328);
xnor U19560 (N_19560,N_19276,N_19422);
nand U19561 (N_19561,N_19468,N_19235);
and U19562 (N_19562,N_19418,N_19445);
nand U19563 (N_19563,N_19443,N_19294);
nor U19564 (N_19564,N_19214,N_19251);
nor U19565 (N_19565,N_19420,N_19216);
nor U19566 (N_19566,N_19306,N_19220);
xnor U19567 (N_19567,N_19340,N_19342);
and U19568 (N_19568,N_19231,N_19466);
nor U19569 (N_19569,N_19224,N_19467);
nor U19570 (N_19570,N_19275,N_19353);
xnor U19571 (N_19571,N_19206,N_19253);
and U19572 (N_19572,N_19481,N_19399);
nand U19573 (N_19573,N_19333,N_19373);
or U19574 (N_19574,N_19372,N_19257);
or U19575 (N_19575,N_19469,N_19354);
xnor U19576 (N_19576,N_19382,N_19236);
nand U19577 (N_19577,N_19431,N_19470);
nor U19578 (N_19578,N_19489,N_19423);
nor U19579 (N_19579,N_19369,N_19295);
and U19580 (N_19580,N_19419,N_19392);
nor U19581 (N_19581,N_19483,N_19278);
nand U19582 (N_19582,N_19336,N_19314);
or U19583 (N_19583,N_19473,N_19298);
nand U19584 (N_19584,N_19338,N_19383);
xor U19585 (N_19585,N_19312,N_19323);
xor U19586 (N_19586,N_19274,N_19437);
xnor U19587 (N_19587,N_19258,N_19486);
xor U19588 (N_19588,N_19394,N_19219);
or U19589 (N_19589,N_19487,N_19492);
xor U19590 (N_19590,N_19310,N_19499);
and U19591 (N_19591,N_19322,N_19485);
nor U19592 (N_19592,N_19299,N_19332);
and U19593 (N_19593,N_19349,N_19405);
xor U19594 (N_19594,N_19267,N_19452);
nand U19595 (N_19595,N_19305,N_19225);
nor U19596 (N_19596,N_19436,N_19459);
or U19597 (N_19597,N_19439,N_19463);
xnor U19598 (N_19598,N_19202,N_19270);
nor U19599 (N_19599,N_19311,N_19218);
or U19600 (N_19600,N_19376,N_19427);
nor U19601 (N_19601,N_19345,N_19371);
nand U19602 (N_19602,N_19200,N_19284);
nand U19603 (N_19603,N_19282,N_19226);
nor U19604 (N_19604,N_19327,N_19246);
nor U19605 (N_19605,N_19248,N_19451);
xor U19606 (N_19606,N_19410,N_19393);
xor U19607 (N_19607,N_19207,N_19351);
and U19608 (N_19608,N_19341,N_19450);
and U19609 (N_19609,N_19498,N_19378);
xor U19610 (N_19610,N_19331,N_19449);
nand U19611 (N_19611,N_19404,N_19279);
or U19612 (N_19612,N_19261,N_19496);
and U19613 (N_19613,N_19293,N_19343);
nor U19614 (N_19614,N_19337,N_19307);
or U19615 (N_19615,N_19401,N_19366);
and U19616 (N_19616,N_19407,N_19456);
and U19617 (N_19617,N_19358,N_19308);
and U19618 (N_19618,N_19212,N_19304);
nor U19619 (N_19619,N_19408,N_19266);
nor U19620 (N_19620,N_19462,N_19347);
or U19621 (N_19621,N_19387,N_19297);
or U19622 (N_19622,N_19367,N_19484);
and U19623 (N_19623,N_19288,N_19490);
nor U19624 (N_19624,N_19428,N_19228);
xor U19625 (N_19625,N_19441,N_19210);
nand U19626 (N_19626,N_19252,N_19245);
nand U19627 (N_19627,N_19321,N_19461);
or U19628 (N_19628,N_19238,N_19412);
xnor U19629 (N_19629,N_19377,N_19334);
xnor U19630 (N_19630,N_19374,N_19380);
nor U19631 (N_19631,N_19375,N_19201);
xnor U19632 (N_19632,N_19287,N_19395);
or U19633 (N_19633,N_19290,N_19300);
nor U19634 (N_19634,N_19223,N_19303);
or U19635 (N_19635,N_19325,N_19213);
nand U19636 (N_19636,N_19247,N_19204);
nor U19637 (N_19637,N_19356,N_19464);
xnor U19638 (N_19638,N_19269,N_19398);
or U19639 (N_19639,N_19494,N_19317);
xor U19640 (N_19640,N_19446,N_19426);
and U19641 (N_19641,N_19313,N_19391);
or U19642 (N_19642,N_19454,N_19411);
nor U19643 (N_19643,N_19442,N_19222);
nor U19644 (N_19644,N_19324,N_19447);
and U19645 (N_19645,N_19348,N_19363);
or U19646 (N_19646,N_19273,N_19460);
or U19647 (N_19647,N_19230,N_19326);
xor U19648 (N_19648,N_19259,N_19476);
or U19649 (N_19649,N_19402,N_19217);
or U19650 (N_19650,N_19292,N_19252);
xor U19651 (N_19651,N_19216,N_19361);
and U19652 (N_19652,N_19200,N_19313);
xor U19653 (N_19653,N_19279,N_19278);
or U19654 (N_19654,N_19325,N_19279);
nand U19655 (N_19655,N_19221,N_19262);
and U19656 (N_19656,N_19232,N_19442);
xnor U19657 (N_19657,N_19292,N_19378);
and U19658 (N_19658,N_19393,N_19313);
nor U19659 (N_19659,N_19467,N_19325);
or U19660 (N_19660,N_19417,N_19210);
nand U19661 (N_19661,N_19489,N_19471);
and U19662 (N_19662,N_19356,N_19300);
nand U19663 (N_19663,N_19397,N_19471);
nor U19664 (N_19664,N_19287,N_19475);
nor U19665 (N_19665,N_19449,N_19446);
xor U19666 (N_19666,N_19312,N_19342);
or U19667 (N_19667,N_19233,N_19354);
or U19668 (N_19668,N_19219,N_19202);
nor U19669 (N_19669,N_19397,N_19312);
or U19670 (N_19670,N_19230,N_19435);
and U19671 (N_19671,N_19303,N_19269);
or U19672 (N_19672,N_19212,N_19253);
nor U19673 (N_19673,N_19276,N_19264);
or U19674 (N_19674,N_19355,N_19219);
and U19675 (N_19675,N_19373,N_19478);
and U19676 (N_19676,N_19365,N_19331);
and U19677 (N_19677,N_19404,N_19480);
and U19678 (N_19678,N_19252,N_19213);
and U19679 (N_19679,N_19277,N_19441);
xnor U19680 (N_19680,N_19351,N_19411);
nand U19681 (N_19681,N_19353,N_19489);
or U19682 (N_19682,N_19350,N_19443);
nand U19683 (N_19683,N_19264,N_19456);
xor U19684 (N_19684,N_19454,N_19346);
and U19685 (N_19685,N_19337,N_19247);
nand U19686 (N_19686,N_19288,N_19357);
nand U19687 (N_19687,N_19312,N_19203);
xor U19688 (N_19688,N_19262,N_19404);
and U19689 (N_19689,N_19223,N_19204);
or U19690 (N_19690,N_19312,N_19346);
xor U19691 (N_19691,N_19338,N_19418);
xor U19692 (N_19692,N_19274,N_19463);
xnor U19693 (N_19693,N_19317,N_19475);
xor U19694 (N_19694,N_19333,N_19270);
nand U19695 (N_19695,N_19491,N_19418);
xor U19696 (N_19696,N_19393,N_19273);
xnor U19697 (N_19697,N_19441,N_19208);
and U19698 (N_19698,N_19289,N_19347);
or U19699 (N_19699,N_19206,N_19205);
xor U19700 (N_19700,N_19420,N_19445);
nand U19701 (N_19701,N_19384,N_19206);
and U19702 (N_19702,N_19311,N_19343);
nor U19703 (N_19703,N_19330,N_19388);
or U19704 (N_19704,N_19270,N_19381);
nor U19705 (N_19705,N_19299,N_19315);
nand U19706 (N_19706,N_19483,N_19393);
nand U19707 (N_19707,N_19365,N_19446);
or U19708 (N_19708,N_19277,N_19263);
and U19709 (N_19709,N_19491,N_19487);
xor U19710 (N_19710,N_19274,N_19296);
nor U19711 (N_19711,N_19406,N_19206);
nor U19712 (N_19712,N_19368,N_19365);
nand U19713 (N_19713,N_19459,N_19375);
nor U19714 (N_19714,N_19302,N_19401);
and U19715 (N_19715,N_19472,N_19388);
xnor U19716 (N_19716,N_19284,N_19325);
nand U19717 (N_19717,N_19268,N_19282);
nor U19718 (N_19718,N_19310,N_19279);
nor U19719 (N_19719,N_19493,N_19236);
nand U19720 (N_19720,N_19357,N_19483);
or U19721 (N_19721,N_19256,N_19456);
xor U19722 (N_19722,N_19250,N_19418);
or U19723 (N_19723,N_19411,N_19303);
nor U19724 (N_19724,N_19459,N_19201);
or U19725 (N_19725,N_19211,N_19450);
xor U19726 (N_19726,N_19480,N_19352);
or U19727 (N_19727,N_19257,N_19339);
xnor U19728 (N_19728,N_19265,N_19466);
nor U19729 (N_19729,N_19434,N_19449);
nand U19730 (N_19730,N_19471,N_19231);
nand U19731 (N_19731,N_19333,N_19495);
nor U19732 (N_19732,N_19290,N_19404);
or U19733 (N_19733,N_19219,N_19450);
or U19734 (N_19734,N_19346,N_19247);
nand U19735 (N_19735,N_19246,N_19326);
or U19736 (N_19736,N_19331,N_19479);
nand U19737 (N_19737,N_19418,N_19214);
nor U19738 (N_19738,N_19264,N_19326);
xnor U19739 (N_19739,N_19309,N_19422);
xor U19740 (N_19740,N_19262,N_19312);
and U19741 (N_19741,N_19351,N_19339);
xnor U19742 (N_19742,N_19490,N_19456);
xnor U19743 (N_19743,N_19206,N_19473);
or U19744 (N_19744,N_19330,N_19368);
and U19745 (N_19745,N_19436,N_19294);
and U19746 (N_19746,N_19437,N_19289);
or U19747 (N_19747,N_19457,N_19467);
or U19748 (N_19748,N_19330,N_19354);
nor U19749 (N_19749,N_19224,N_19216);
xnor U19750 (N_19750,N_19296,N_19276);
or U19751 (N_19751,N_19289,N_19471);
xnor U19752 (N_19752,N_19219,N_19314);
xor U19753 (N_19753,N_19466,N_19346);
nor U19754 (N_19754,N_19225,N_19397);
nor U19755 (N_19755,N_19266,N_19440);
and U19756 (N_19756,N_19256,N_19367);
xor U19757 (N_19757,N_19341,N_19332);
xnor U19758 (N_19758,N_19335,N_19465);
or U19759 (N_19759,N_19497,N_19288);
xor U19760 (N_19760,N_19487,N_19204);
nand U19761 (N_19761,N_19334,N_19475);
or U19762 (N_19762,N_19446,N_19430);
or U19763 (N_19763,N_19339,N_19231);
nand U19764 (N_19764,N_19435,N_19298);
nand U19765 (N_19765,N_19472,N_19230);
nor U19766 (N_19766,N_19385,N_19215);
xor U19767 (N_19767,N_19283,N_19395);
xnor U19768 (N_19768,N_19336,N_19445);
and U19769 (N_19769,N_19324,N_19273);
nor U19770 (N_19770,N_19403,N_19395);
or U19771 (N_19771,N_19257,N_19209);
and U19772 (N_19772,N_19246,N_19243);
nand U19773 (N_19773,N_19315,N_19476);
or U19774 (N_19774,N_19367,N_19232);
and U19775 (N_19775,N_19305,N_19268);
or U19776 (N_19776,N_19410,N_19314);
xnor U19777 (N_19777,N_19348,N_19435);
xor U19778 (N_19778,N_19436,N_19359);
or U19779 (N_19779,N_19466,N_19497);
and U19780 (N_19780,N_19308,N_19391);
nor U19781 (N_19781,N_19214,N_19322);
xnor U19782 (N_19782,N_19260,N_19344);
xnor U19783 (N_19783,N_19239,N_19327);
xnor U19784 (N_19784,N_19294,N_19371);
nor U19785 (N_19785,N_19236,N_19329);
nand U19786 (N_19786,N_19208,N_19303);
and U19787 (N_19787,N_19211,N_19497);
or U19788 (N_19788,N_19239,N_19417);
or U19789 (N_19789,N_19249,N_19462);
nor U19790 (N_19790,N_19357,N_19254);
and U19791 (N_19791,N_19327,N_19275);
nand U19792 (N_19792,N_19303,N_19205);
xor U19793 (N_19793,N_19486,N_19440);
and U19794 (N_19794,N_19408,N_19290);
nor U19795 (N_19795,N_19375,N_19480);
or U19796 (N_19796,N_19205,N_19436);
nand U19797 (N_19797,N_19400,N_19229);
xor U19798 (N_19798,N_19210,N_19205);
nor U19799 (N_19799,N_19214,N_19372);
nand U19800 (N_19800,N_19558,N_19726);
xor U19801 (N_19801,N_19730,N_19565);
xnor U19802 (N_19802,N_19764,N_19788);
xor U19803 (N_19803,N_19670,N_19671);
and U19804 (N_19804,N_19537,N_19566);
or U19805 (N_19805,N_19744,N_19756);
and U19806 (N_19806,N_19599,N_19592);
nor U19807 (N_19807,N_19614,N_19704);
nor U19808 (N_19808,N_19669,N_19607);
nor U19809 (N_19809,N_19560,N_19602);
xnor U19810 (N_19810,N_19604,N_19725);
nor U19811 (N_19811,N_19683,N_19742);
nand U19812 (N_19812,N_19572,N_19612);
nand U19813 (N_19813,N_19555,N_19674);
or U19814 (N_19814,N_19628,N_19751);
or U19815 (N_19815,N_19775,N_19644);
nor U19816 (N_19816,N_19777,N_19780);
and U19817 (N_19817,N_19773,N_19701);
or U19818 (N_19818,N_19650,N_19584);
xnor U19819 (N_19819,N_19506,N_19544);
and U19820 (N_19820,N_19507,N_19731);
and U19821 (N_19821,N_19649,N_19750);
nand U19822 (N_19822,N_19527,N_19790);
nand U19823 (N_19823,N_19700,N_19522);
nor U19824 (N_19824,N_19706,N_19711);
nor U19825 (N_19825,N_19760,N_19797);
nor U19826 (N_19826,N_19747,N_19697);
or U19827 (N_19827,N_19647,N_19517);
and U19828 (N_19828,N_19651,N_19564);
or U19829 (N_19829,N_19745,N_19574);
or U19830 (N_19830,N_19720,N_19518);
xnor U19831 (N_19831,N_19677,N_19682);
nand U19832 (N_19832,N_19695,N_19765);
and U19833 (N_19833,N_19668,N_19769);
xor U19834 (N_19834,N_19571,N_19637);
or U19835 (N_19835,N_19660,N_19792);
nand U19836 (N_19836,N_19579,N_19728);
and U19837 (N_19837,N_19559,N_19707);
nor U19838 (N_19838,N_19646,N_19641);
or U19839 (N_19839,N_19575,N_19676);
xor U19840 (N_19840,N_19580,N_19761);
nand U19841 (N_19841,N_19759,N_19534);
or U19842 (N_19842,N_19684,N_19620);
nand U19843 (N_19843,N_19638,N_19783);
xnor U19844 (N_19844,N_19784,N_19598);
and U19845 (N_19845,N_19548,N_19772);
xnor U19846 (N_19846,N_19787,N_19521);
xnor U19847 (N_19847,N_19531,N_19547);
xor U19848 (N_19848,N_19734,N_19736);
nand U19849 (N_19849,N_19729,N_19689);
or U19850 (N_19850,N_19500,N_19746);
and U19851 (N_19851,N_19743,N_19524);
nand U19852 (N_19852,N_19662,N_19755);
xor U19853 (N_19853,N_19569,N_19648);
nand U19854 (N_19854,N_19545,N_19699);
xnor U19855 (N_19855,N_19675,N_19610);
and U19856 (N_19856,N_19779,N_19563);
nor U19857 (N_19857,N_19738,N_19654);
nand U19858 (N_19858,N_19735,N_19741);
nand U19859 (N_19859,N_19640,N_19538);
or U19860 (N_19860,N_19724,N_19549);
or U19861 (N_19861,N_19526,N_19514);
nand U19862 (N_19862,N_19757,N_19794);
and U19863 (N_19863,N_19578,N_19611);
and U19864 (N_19864,N_19619,N_19634);
and U19865 (N_19865,N_19515,N_19632);
nand U19866 (N_19866,N_19661,N_19719);
nor U19867 (N_19867,N_19615,N_19656);
nor U19868 (N_19868,N_19696,N_19723);
nand U19869 (N_19869,N_19550,N_19593);
nand U19870 (N_19870,N_19588,N_19519);
or U19871 (N_19871,N_19766,N_19561);
xor U19872 (N_19872,N_19739,N_19582);
and U19873 (N_19873,N_19771,N_19733);
nor U19874 (N_19874,N_19636,N_19600);
or U19875 (N_19875,N_19710,N_19606);
and U19876 (N_19876,N_19781,N_19631);
nand U19877 (N_19877,N_19655,N_19520);
nand U19878 (N_19878,N_19786,N_19796);
nor U19879 (N_19879,N_19658,N_19504);
xnor U19880 (N_19880,N_19552,N_19703);
and U19881 (N_19881,N_19645,N_19732);
nand U19882 (N_19882,N_19618,N_19768);
and U19883 (N_19883,N_19798,N_19546);
and U19884 (N_19884,N_19530,N_19663);
or U19885 (N_19885,N_19613,N_19740);
nor U19886 (N_19886,N_19659,N_19597);
xor U19887 (N_19887,N_19554,N_19627);
nand U19888 (N_19888,N_19688,N_19562);
or U19889 (N_19889,N_19687,N_19528);
nor U19890 (N_19890,N_19727,N_19587);
and U19891 (N_19891,N_19667,N_19541);
or U19892 (N_19892,N_19774,N_19573);
nand U19893 (N_19893,N_19502,N_19539);
and U19894 (N_19894,N_19625,N_19789);
nand U19895 (N_19895,N_19754,N_19693);
xnor U19896 (N_19896,N_19595,N_19623);
nand U19897 (N_19897,N_19763,N_19679);
nand U19898 (N_19898,N_19624,N_19510);
nor U19899 (N_19899,N_19712,N_19568);
or U19900 (N_19900,N_19605,N_19666);
and U19901 (N_19901,N_19785,N_19553);
nor U19902 (N_19902,N_19664,N_19694);
or U19903 (N_19903,N_19749,N_19673);
and U19904 (N_19904,N_19702,N_19608);
nand U19905 (N_19905,N_19770,N_19533);
nand U19906 (N_19906,N_19799,N_19525);
nand U19907 (N_19907,N_19715,N_19503);
or U19908 (N_19908,N_19680,N_19714);
xnor U19909 (N_19909,N_19616,N_19629);
nand U19910 (N_19910,N_19653,N_19685);
or U19911 (N_19911,N_19508,N_19591);
nand U19912 (N_19912,N_19551,N_19639);
or U19913 (N_19913,N_19718,N_19795);
nand U19914 (N_19914,N_19652,N_19642);
xnor U19915 (N_19915,N_19776,N_19512);
xor U19916 (N_19916,N_19705,N_19630);
or U19917 (N_19917,N_19557,N_19617);
or U19918 (N_19918,N_19535,N_19635);
nor U19919 (N_19919,N_19511,N_19713);
nand U19920 (N_19920,N_19692,N_19516);
xnor U19921 (N_19921,N_19657,N_19621);
xor U19922 (N_19922,N_19708,N_19716);
and U19923 (N_19923,N_19532,N_19603);
and U19924 (N_19924,N_19633,N_19509);
and U19925 (N_19925,N_19542,N_19583);
xor U19926 (N_19926,N_19793,N_19622);
xor U19927 (N_19927,N_19540,N_19594);
or U19928 (N_19928,N_19556,N_19536);
xor U19929 (N_19929,N_19513,N_19505);
nand U19930 (N_19930,N_19678,N_19681);
xnor U19931 (N_19931,N_19665,N_19529);
and U19932 (N_19932,N_19782,N_19601);
xnor U19933 (N_19933,N_19778,N_19581);
nand U19934 (N_19934,N_19643,N_19672);
nor U19935 (N_19935,N_19758,N_19698);
or U19936 (N_19936,N_19709,N_19543);
or U19937 (N_19937,N_19791,N_19686);
and U19938 (N_19938,N_19596,N_19609);
or U19939 (N_19939,N_19570,N_19753);
and U19940 (N_19940,N_19589,N_19585);
nand U19941 (N_19941,N_19762,N_19767);
and U19942 (N_19942,N_19717,N_19691);
and U19943 (N_19943,N_19523,N_19690);
nor U19944 (N_19944,N_19748,N_19752);
nand U19945 (N_19945,N_19722,N_19626);
nand U19946 (N_19946,N_19737,N_19576);
or U19947 (N_19947,N_19586,N_19721);
and U19948 (N_19948,N_19567,N_19577);
and U19949 (N_19949,N_19590,N_19501);
and U19950 (N_19950,N_19731,N_19610);
nand U19951 (N_19951,N_19579,N_19706);
or U19952 (N_19952,N_19651,N_19626);
nand U19953 (N_19953,N_19769,N_19624);
xnor U19954 (N_19954,N_19738,N_19627);
xnor U19955 (N_19955,N_19534,N_19785);
or U19956 (N_19956,N_19688,N_19706);
xnor U19957 (N_19957,N_19634,N_19675);
and U19958 (N_19958,N_19796,N_19547);
xor U19959 (N_19959,N_19620,N_19743);
xnor U19960 (N_19960,N_19563,N_19530);
xor U19961 (N_19961,N_19640,N_19611);
xnor U19962 (N_19962,N_19772,N_19774);
or U19963 (N_19963,N_19534,N_19529);
nand U19964 (N_19964,N_19655,N_19792);
or U19965 (N_19965,N_19695,N_19546);
or U19966 (N_19966,N_19531,N_19751);
and U19967 (N_19967,N_19566,N_19525);
nor U19968 (N_19968,N_19627,N_19513);
and U19969 (N_19969,N_19757,N_19508);
xor U19970 (N_19970,N_19727,N_19626);
or U19971 (N_19971,N_19721,N_19732);
xnor U19972 (N_19972,N_19706,N_19695);
or U19973 (N_19973,N_19753,N_19789);
xor U19974 (N_19974,N_19742,N_19522);
or U19975 (N_19975,N_19727,N_19741);
and U19976 (N_19976,N_19730,N_19593);
or U19977 (N_19977,N_19758,N_19600);
or U19978 (N_19978,N_19718,N_19672);
nor U19979 (N_19979,N_19555,N_19551);
xor U19980 (N_19980,N_19695,N_19794);
nor U19981 (N_19981,N_19530,N_19733);
nand U19982 (N_19982,N_19618,N_19657);
and U19983 (N_19983,N_19677,N_19690);
nor U19984 (N_19984,N_19799,N_19573);
or U19985 (N_19985,N_19547,N_19506);
or U19986 (N_19986,N_19506,N_19765);
and U19987 (N_19987,N_19614,N_19560);
and U19988 (N_19988,N_19522,N_19643);
xor U19989 (N_19989,N_19585,N_19508);
and U19990 (N_19990,N_19718,N_19604);
nand U19991 (N_19991,N_19595,N_19752);
nand U19992 (N_19992,N_19741,N_19797);
or U19993 (N_19993,N_19510,N_19793);
nor U19994 (N_19994,N_19781,N_19771);
nand U19995 (N_19995,N_19639,N_19589);
and U19996 (N_19996,N_19583,N_19540);
and U19997 (N_19997,N_19773,N_19697);
or U19998 (N_19998,N_19727,N_19561);
nor U19999 (N_19999,N_19617,N_19770);
nand U20000 (N_20000,N_19663,N_19565);
or U20001 (N_20001,N_19608,N_19606);
xnor U20002 (N_20002,N_19706,N_19558);
nand U20003 (N_20003,N_19679,N_19712);
and U20004 (N_20004,N_19797,N_19704);
nor U20005 (N_20005,N_19502,N_19553);
nand U20006 (N_20006,N_19512,N_19575);
nor U20007 (N_20007,N_19615,N_19616);
and U20008 (N_20008,N_19618,N_19785);
nand U20009 (N_20009,N_19763,N_19783);
xnor U20010 (N_20010,N_19681,N_19512);
xor U20011 (N_20011,N_19692,N_19574);
and U20012 (N_20012,N_19610,N_19556);
or U20013 (N_20013,N_19743,N_19717);
xor U20014 (N_20014,N_19700,N_19723);
or U20015 (N_20015,N_19699,N_19600);
nand U20016 (N_20016,N_19714,N_19534);
xor U20017 (N_20017,N_19692,N_19747);
xor U20018 (N_20018,N_19665,N_19584);
xor U20019 (N_20019,N_19609,N_19681);
xor U20020 (N_20020,N_19622,N_19794);
nor U20021 (N_20021,N_19629,N_19518);
or U20022 (N_20022,N_19694,N_19750);
nand U20023 (N_20023,N_19732,N_19770);
nor U20024 (N_20024,N_19766,N_19786);
or U20025 (N_20025,N_19738,N_19735);
xor U20026 (N_20026,N_19567,N_19543);
nand U20027 (N_20027,N_19597,N_19546);
xor U20028 (N_20028,N_19597,N_19570);
nor U20029 (N_20029,N_19501,N_19601);
xor U20030 (N_20030,N_19690,N_19682);
xor U20031 (N_20031,N_19606,N_19744);
nand U20032 (N_20032,N_19646,N_19552);
xor U20033 (N_20033,N_19617,N_19763);
and U20034 (N_20034,N_19733,N_19716);
and U20035 (N_20035,N_19581,N_19501);
or U20036 (N_20036,N_19720,N_19511);
or U20037 (N_20037,N_19607,N_19711);
xor U20038 (N_20038,N_19690,N_19708);
or U20039 (N_20039,N_19623,N_19679);
xnor U20040 (N_20040,N_19598,N_19707);
nor U20041 (N_20041,N_19635,N_19555);
or U20042 (N_20042,N_19547,N_19569);
or U20043 (N_20043,N_19758,N_19689);
and U20044 (N_20044,N_19748,N_19781);
xor U20045 (N_20045,N_19784,N_19768);
nor U20046 (N_20046,N_19728,N_19595);
xor U20047 (N_20047,N_19715,N_19780);
or U20048 (N_20048,N_19576,N_19774);
xor U20049 (N_20049,N_19694,N_19692);
and U20050 (N_20050,N_19684,N_19744);
and U20051 (N_20051,N_19568,N_19644);
xor U20052 (N_20052,N_19790,N_19682);
and U20053 (N_20053,N_19661,N_19767);
xor U20054 (N_20054,N_19644,N_19681);
and U20055 (N_20055,N_19793,N_19555);
nor U20056 (N_20056,N_19667,N_19591);
and U20057 (N_20057,N_19563,N_19708);
nand U20058 (N_20058,N_19666,N_19796);
or U20059 (N_20059,N_19775,N_19539);
xor U20060 (N_20060,N_19504,N_19537);
and U20061 (N_20061,N_19545,N_19720);
or U20062 (N_20062,N_19580,N_19757);
nand U20063 (N_20063,N_19630,N_19598);
nor U20064 (N_20064,N_19755,N_19690);
nor U20065 (N_20065,N_19678,N_19557);
nand U20066 (N_20066,N_19712,N_19678);
nand U20067 (N_20067,N_19775,N_19677);
or U20068 (N_20068,N_19620,N_19788);
and U20069 (N_20069,N_19518,N_19561);
or U20070 (N_20070,N_19631,N_19573);
nand U20071 (N_20071,N_19631,N_19768);
and U20072 (N_20072,N_19584,N_19601);
or U20073 (N_20073,N_19523,N_19547);
and U20074 (N_20074,N_19727,N_19510);
or U20075 (N_20075,N_19566,N_19757);
or U20076 (N_20076,N_19655,N_19608);
nand U20077 (N_20077,N_19771,N_19743);
and U20078 (N_20078,N_19762,N_19580);
or U20079 (N_20079,N_19623,N_19516);
or U20080 (N_20080,N_19662,N_19611);
or U20081 (N_20081,N_19635,N_19717);
and U20082 (N_20082,N_19530,N_19610);
nor U20083 (N_20083,N_19657,N_19717);
nor U20084 (N_20084,N_19627,N_19707);
nor U20085 (N_20085,N_19579,N_19738);
xnor U20086 (N_20086,N_19778,N_19682);
nand U20087 (N_20087,N_19798,N_19566);
nand U20088 (N_20088,N_19521,N_19694);
nor U20089 (N_20089,N_19616,N_19685);
xnor U20090 (N_20090,N_19753,N_19761);
or U20091 (N_20091,N_19694,N_19568);
or U20092 (N_20092,N_19518,N_19558);
and U20093 (N_20093,N_19598,N_19572);
nor U20094 (N_20094,N_19541,N_19789);
or U20095 (N_20095,N_19617,N_19538);
and U20096 (N_20096,N_19616,N_19753);
nand U20097 (N_20097,N_19603,N_19663);
and U20098 (N_20098,N_19574,N_19761);
and U20099 (N_20099,N_19568,N_19725);
and U20100 (N_20100,N_19820,N_20093);
nor U20101 (N_20101,N_20049,N_19813);
and U20102 (N_20102,N_19832,N_20053);
nand U20103 (N_20103,N_19874,N_20003);
or U20104 (N_20104,N_19964,N_19912);
xor U20105 (N_20105,N_19816,N_20031);
xor U20106 (N_20106,N_19908,N_19935);
and U20107 (N_20107,N_19992,N_20009);
and U20108 (N_20108,N_19986,N_19914);
and U20109 (N_20109,N_19839,N_19865);
nor U20110 (N_20110,N_19965,N_19825);
or U20111 (N_20111,N_20072,N_19971);
nor U20112 (N_20112,N_20043,N_19940);
xor U20113 (N_20113,N_19847,N_19920);
xnor U20114 (N_20114,N_19999,N_19862);
nor U20115 (N_20115,N_19909,N_19899);
or U20116 (N_20116,N_19973,N_20007);
xor U20117 (N_20117,N_19824,N_20061);
nor U20118 (N_20118,N_19948,N_20099);
xnor U20119 (N_20119,N_19900,N_19919);
or U20120 (N_20120,N_19924,N_19843);
and U20121 (N_20121,N_19864,N_19962);
nand U20122 (N_20122,N_19903,N_20075);
and U20123 (N_20123,N_19810,N_20037);
nand U20124 (N_20124,N_19979,N_20096);
xor U20125 (N_20125,N_19907,N_19978);
nor U20126 (N_20126,N_19995,N_19845);
and U20127 (N_20127,N_19927,N_20006);
or U20128 (N_20128,N_19980,N_20088);
nand U20129 (N_20129,N_20079,N_19819);
and U20130 (N_20130,N_19858,N_19829);
and U20131 (N_20131,N_20056,N_19991);
nor U20132 (N_20132,N_19837,N_19906);
xor U20133 (N_20133,N_19806,N_19939);
xnor U20134 (N_20134,N_20091,N_19867);
or U20135 (N_20135,N_19803,N_19976);
nor U20136 (N_20136,N_19898,N_19852);
or U20137 (N_20137,N_19996,N_19882);
and U20138 (N_20138,N_20055,N_19823);
nor U20139 (N_20139,N_19990,N_19884);
xor U20140 (N_20140,N_19835,N_19818);
and U20141 (N_20141,N_20012,N_20021);
nand U20142 (N_20142,N_19970,N_19896);
nor U20143 (N_20143,N_20022,N_19915);
xor U20144 (N_20144,N_20074,N_19840);
nand U20145 (N_20145,N_20014,N_19945);
nor U20146 (N_20146,N_20062,N_20040);
and U20147 (N_20147,N_19925,N_19985);
or U20148 (N_20148,N_19851,N_19854);
and U20149 (N_20149,N_19894,N_19998);
nor U20150 (N_20150,N_19870,N_19941);
or U20151 (N_20151,N_20057,N_20016);
or U20152 (N_20152,N_20017,N_20029);
nor U20153 (N_20153,N_20095,N_20038);
xor U20154 (N_20154,N_20033,N_19827);
or U20155 (N_20155,N_19929,N_19989);
or U20156 (N_20156,N_19866,N_19955);
nor U20157 (N_20157,N_19890,N_19872);
nor U20158 (N_20158,N_20023,N_19984);
or U20159 (N_20159,N_20000,N_20066);
xnor U20160 (N_20160,N_20078,N_20086);
and U20161 (N_20161,N_19807,N_19983);
nand U20162 (N_20162,N_19834,N_19959);
and U20163 (N_20163,N_19863,N_19949);
and U20164 (N_20164,N_19848,N_20024);
nand U20165 (N_20165,N_20005,N_19951);
xor U20166 (N_20166,N_19841,N_20090);
xor U20167 (N_20167,N_20076,N_19885);
and U20168 (N_20168,N_19931,N_20051);
and U20169 (N_20169,N_19932,N_20001);
xnor U20170 (N_20170,N_19917,N_19873);
xor U20171 (N_20171,N_20071,N_19893);
nand U20172 (N_20172,N_20008,N_19956);
nor U20173 (N_20173,N_19812,N_20013);
and U20174 (N_20174,N_20094,N_20042);
nor U20175 (N_20175,N_19936,N_20026);
xnor U20176 (N_20176,N_20052,N_20045);
xor U20177 (N_20177,N_19857,N_19879);
xor U20178 (N_20178,N_19902,N_20025);
and U20179 (N_20179,N_20039,N_19937);
or U20180 (N_20180,N_20087,N_19960);
xnor U20181 (N_20181,N_19997,N_19846);
and U20182 (N_20182,N_20050,N_19911);
and U20183 (N_20183,N_20028,N_19887);
nand U20184 (N_20184,N_19856,N_19889);
or U20185 (N_20185,N_20044,N_19933);
or U20186 (N_20186,N_19868,N_19930);
nand U20187 (N_20187,N_19968,N_20085);
nor U20188 (N_20188,N_19888,N_19904);
nor U20189 (N_20189,N_20048,N_19831);
nand U20190 (N_20190,N_19871,N_19981);
xnor U20191 (N_20191,N_20070,N_19875);
or U20192 (N_20192,N_19828,N_19926);
and U20193 (N_20193,N_19836,N_19811);
xnor U20194 (N_20194,N_19877,N_19891);
nor U20195 (N_20195,N_20092,N_19859);
xor U20196 (N_20196,N_20034,N_20084);
or U20197 (N_20197,N_19958,N_20069);
and U20198 (N_20198,N_19928,N_20027);
nor U20199 (N_20199,N_19988,N_19838);
xor U20200 (N_20200,N_19922,N_19947);
xor U20201 (N_20201,N_19817,N_19961);
and U20202 (N_20202,N_19876,N_19886);
and U20203 (N_20203,N_19974,N_20060);
nand U20204 (N_20204,N_19916,N_19861);
nand U20205 (N_20205,N_20064,N_19952);
or U20206 (N_20206,N_20015,N_20010);
or U20207 (N_20207,N_19869,N_19969);
xnor U20208 (N_20208,N_20041,N_19880);
nand U20209 (N_20209,N_19972,N_20068);
xnor U20210 (N_20210,N_19977,N_20047);
or U20211 (N_20211,N_19821,N_19901);
nor U20212 (N_20212,N_19921,N_20067);
nand U20213 (N_20213,N_19953,N_19913);
and U20214 (N_20214,N_20098,N_20030);
xor U20215 (N_20215,N_20083,N_19943);
xnor U20216 (N_20216,N_19822,N_19830);
xor U20217 (N_20217,N_19923,N_20065);
xor U20218 (N_20218,N_20036,N_19801);
nor U20219 (N_20219,N_19814,N_19982);
and U20220 (N_20220,N_20059,N_19881);
xnor U20221 (N_20221,N_20035,N_20097);
or U20222 (N_20222,N_19826,N_19954);
nor U20223 (N_20223,N_20073,N_19910);
or U20224 (N_20224,N_20081,N_19878);
and U20225 (N_20225,N_20058,N_19897);
nand U20226 (N_20226,N_20080,N_20004);
nand U20227 (N_20227,N_19905,N_20089);
nand U20228 (N_20228,N_19963,N_19805);
or U20229 (N_20229,N_19950,N_19967);
xnor U20230 (N_20230,N_20002,N_19993);
or U20231 (N_20231,N_20019,N_20054);
xor U20232 (N_20232,N_19987,N_19860);
and U20233 (N_20233,N_19942,N_20063);
and U20234 (N_20234,N_19946,N_19809);
nor U20235 (N_20235,N_19842,N_20020);
xnor U20236 (N_20236,N_19957,N_19802);
and U20237 (N_20237,N_20082,N_19892);
or U20238 (N_20238,N_19944,N_19934);
and U20239 (N_20239,N_19994,N_19850);
or U20240 (N_20240,N_19895,N_19833);
and U20241 (N_20241,N_19918,N_20077);
or U20242 (N_20242,N_20046,N_19849);
xnor U20243 (N_20243,N_19975,N_19800);
nor U20244 (N_20244,N_19804,N_19815);
xor U20245 (N_20245,N_19966,N_19808);
nor U20246 (N_20246,N_19844,N_20032);
and U20247 (N_20247,N_19855,N_20018);
and U20248 (N_20248,N_19883,N_19938);
nor U20249 (N_20249,N_19853,N_20011);
and U20250 (N_20250,N_19963,N_19819);
or U20251 (N_20251,N_20089,N_19848);
xnor U20252 (N_20252,N_19997,N_19801);
nor U20253 (N_20253,N_19905,N_19809);
xnor U20254 (N_20254,N_20041,N_19821);
nor U20255 (N_20255,N_19814,N_19926);
and U20256 (N_20256,N_20083,N_20014);
and U20257 (N_20257,N_19821,N_20071);
and U20258 (N_20258,N_19831,N_19936);
nand U20259 (N_20259,N_20006,N_19868);
and U20260 (N_20260,N_20040,N_19980);
and U20261 (N_20261,N_20097,N_19849);
nand U20262 (N_20262,N_20040,N_19937);
or U20263 (N_20263,N_19847,N_20098);
or U20264 (N_20264,N_19830,N_20034);
nor U20265 (N_20265,N_19863,N_19807);
xnor U20266 (N_20266,N_19884,N_19849);
nor U20267 (N_20267,N_19943,N_19974);
or U20268 (N_20268,N_20092,N_20019);
and U20269 (N_20269,N_20087,N_20072);
xnor U20270 (N_20270,N_19964,N_19821);
nand U20271 (N_20271,N_19903,N_20060);
nand U20272 (N_20272,N_19901,N_19965);
or U20273 (N_20273,N_19942,N_19818);
or U20274 (N_20274,N_19972,N_20088);
xnor U20275 (N_20275,N_19864,N_19979);
nor U20276 (N_20276,N_19857,N_20050);
nor U20277 (N_20277,N_19963,N_19860);
nand U20278 (N_20278,N_19983,N_19906);
or U20279 (N_20279,N_19978,N_19991);
xnor U20280 (N_20280,N_19883,N_19892);
xor U20281 (N_20281,N_19822,N_19991);
and U20282 (N_20282,N_19873,N_19932);
nor U20283 (N_20283,N_19817,N_20007);
nor U20284 (N_20284,N_19903,N_20097);
nand U20285 (N_20285,N_19964,N_19873);
or U20286 (N_20286,N_19944,N_20092);
xor U20287 (N_20287,N_19884,N_20051);
nor U20288 (N_20288,N_20076,N_19958);
nor U20289 (N_20289,N_19883,N_19837);
nand U20290 (N_20290,N_20071,N_19919);
nor U20291 (N_20291,N_19900,N_19826);
or U20292 (N_20292,N_20033,N_20074);
and U20293 (N_20293,N_20044,N_19807);
and U20294 (N_20294,N_19888,N_19808);
or U20295 (N_20295,N_19803,N_19843);
xnor U20296 (N_20296,N_19861,N_20003);
or U20297 (N_20297,N_19858,N_20051);
nand U20298 (N_20298,N_20056,N_20079);
nor U20299 (N_20299,N_19846,N_19974);
and U20300 (N_20300,N_19851,N_20038);
nand U20301 (N_20301,N_20034,N_19878);
nand U20302 (N_20302,N_19877,N_19863);
xnor U20303 (N_20303,N_19931,N_19948);
nand U20304 (N_20304,N_19909,N_20090);
or U20305 (N_20305,N_19968,N_19981);
nand U20306 (N_20306,N_19952,N_19933);
nor U20307 (N_20307,N_19840,N_19891);
and U20308 (N_20308,N_20035,N_19983);
and U20309 (N_20309,N_19885,N_19974);
nand U20310 (N_20310,N_19939,N_19970);
or U20311 (N_20311,N_20097,N_19978);
nand U20312 (N_20312,N_19811,N_19950);
or U20313 (N_20313,N_19810,N_20095);
and U20314 (N_20314,N_19999,N_19912);
or U20315 (N_20315,N_19974,N_20031);
xnor U20316 (N_20316,N_20004,N_19886);
or U20317 (N_20317,N_19876,N_20011);
or U20318 (N_20318,N_20066,N_19877);
xor U20319 (N_20319,N_19867,N_19936);
xnor U20320 (N_20320,N_20029,N_19863);
nand U20321 (N_20321,N_19872,N_19907);
nand U20322 (N_20322,N_19928,N_20024);
nand U20323 (N_20323,N_19913,N_20082);
and U20324 (N_20324,N_19942,N_20007);
nand U20325 (N_20325,N_20046,N_20034);
or U20326 (N_20326,N_20039,N_20064);
and U20327 (N_20327,N_19998,N_19960);
nor U20328 (N_20328,N_19890,N_19919);
and U20329 (N_20329,N_19948,N_20025);
or U20330 (N_20330,N_19836,N_19969);
nor U20331 (N_20331,N_19825,N_20048);
xor U20332 (N_20332,N_19837,N_19945);
or U20333 (N_20333,N_19958,N_20065);
nor U20334 (N_20334,N_20076,N_19823);
nor U20335 (N_20335,N_20061,N_19993);
and U20336 (N_20336,N_20083,N_20035);
and U20337 (N_20337,N_19946,N_19971);
nor U20338 (N_20338,N_20018,N_19807);
nor U20339 (N_20339,N_19911,N_20001);
nor U20340 (N_20340,N_19969,N_19823);
nor U20341 (N_20341,N_19917,N_19941);
or U20342 (N_20342,N_19879,N_19902);
nand U20343 (N_20343,N_19808,N_19822);
xor U20344 (N_20344,N_19936,N_19915);
or U20345 (N_20345,N_20009,N_19801);
and U20346 (N_20346,N_19880,N_20071);
xor U20347 (N_20347,N_19825,N_20055);
or U20348 (N_20348,N_19894,N_19841);
nand U20349 (N_20349,N_20003,N_19977);
nor U20350 (N_20350,N_19847,N_20094);
nor U20351 (N_20351,N_19864,N_20067);
nand U20352 (N_20352,N_20071,N_19810);
and U20353 (N_20353,N_20071,N_19973);
and U20354 (N_20354,N_20016,N_19985);
nand U20355 (N_20355,N_19987,N_19831);
xnor U20356 (N_20356,N_19968,N_19971);
and U20357 (N_20357,N_20030,N_19854);
xor U20358 (N_20358,N_19850,N_19990);
xor U20359 (N_20359,N_19915,N_20089);
nor U20360 (N_20360,N_20011,N_20057);
nand U20361 (N_20361,N_20064,N_19985);
nand U20362 (N_20362,N_19863,N_19891);
nand U20363 (N_20363,N_19832,N_19807);
nand U20364 (N_20364,N_19847,N_20067);
nand U20365 (N_20365,N_19812,N_19887);
nor U20366 (N_20366,N_20092,N_20069);
xor U20367 (N_20367,N_19845,N_20054);
and U20368 (N_20368,N_19958,N_20056);
nor U20369 (N_20369,N_20006,N_19819);
and U20370 (N_20370,N_19890,N_19805);
xor U20371 (N_20371,N_19926,N_20064);
nand U20372 (N_20372,N_19835,N_19841);
or U20373 (N_20373,N_20003,N_19981);
xnor U20374 (N_20374,N_19891,N_19842);
nor U20375 (N_20375,N_20065,N_19980);
and U20376 (N_20376,N_19863,N_19961);
and U20377 (N_20377,N_19871,N_19914);
xnor U20378 (N_20378,N_19998,N_20035);
xnor U20379 (N_20379,N_19923,N_19834);
and U20380 (N_20380,N_19884,N_20066);
nand U20381 (N_20381,N_19933,N_19851);
and U20382 (N_20382,N_19891,N_20081);
or U20383 (N_20383,N_19805,N_20042);
xnor U20384 (N_20384,N_19904,N_19803);
nand U20385 (N_20385,N_19983,N_19814);
or U20386 (N_20386,N_20007,N_20097);
nor U20387 (N_20387,N_19962,N_19933);
nor U20388 (N_20388,N_19876,N_20093);
and U20389 (N_20389,N_20008,N_19982);
nand U20390 (N_20390,N_19934,N_20013);
xor U20391 (N_20391,N_20026,N_20038);
or U20392 (N_20392,N_19901,N_19954);
or U20393 (N_20393,N_20042,N_19927);
nor U20394 (N_20394,N_20006,N_19896);
nand U20395 (N_20395,N_19986,N_19847);
xor U20396 (N_20396,N_19904,N_19873);
or U20397 (N_20397,N_19844,N_20033);
xor U20398 (N_20398,N_20079,N_19845);
nand U20399 (N_20399,N_20021,N_20086);
nor U20400 (N_20400,N_20144,N_20110);
xnor U20401 (N_20401,N_20156,N_20148);
or U20402 (N_20402,N_20134,N_20123);
xor U20403 (N_20403,N_20168,N_20130);
nor U20404 (N_20404,N_20310,N_20145);
or U20405 (N_20405,N_20248,N_20389);
nor U20406 (N_20406,N_20299,N_20139);
or U20407 (N_20407,N_20220,N_20141);
or U20408 (N_20408,N_20377,N_20385);
xor U20409 (N_20409,N_20250,N_20395);
xor U20410 (N_20410,N_20300,N_20172);
or U20411 (N_20411,N_20323,N_20115);
or U20412 (N_20412,N_20266,N_20133);
and U20413 (N_20413,N_20313,N_20338);
nand U20414 (N_20414,N_20177,N_20382);
xnor U20415 (N_20415,N_20329,N_20128);
and U20416 (N_20416,N_20147,N_20278);
nor U20417 (N_20417,N_20324,N_20166);
nor U20418 (N_20418,N_20244,N_20143);
nand U20419 (N_20419,N_20142,N_20288);
xnor U20420 (N_20420,N_20174,N_20397);
and U20421 (N_20421,N_20202,N_20352);
nand U20422 (N_20422,N_20232,N_20112);
xnor U20423 (N_20423,N_20341,N_20225);
and U20424 (N_20424,N_20118,N_20107);
nand U20425 (N_20425,N_20277,N_20276);
nand U20426 (N_20426,N_20175,N_20303);
xor U20427 (N_20427,N_20321,N_20293);
xnor U20428 (N_20428,N_20355,N_20103);
and U20429 (N_20429,N_20196,N_20235);
nor U20430 (N_20430,N_20302,N_20108);
or U20431 (N_20431,N_20273,N_20146);
or U20432 (N_20432,N_20369,N_20219);
nor U20433 (N_20433,N_20383,N_20368);
nor U20434 (N_20434,N_20239,N_20131);
or U20435 (N_20435,N_20178,N_20218);
xor U20436 (N_20436,N_20325,N_20348);
nor U20437 (N_20437,N_20316,N_20376);
and U20438 (N_20438,N_20167,N_20330);
nand U20439 (N_20439,N_20217,N_20315);
nor U20440 (N_20440,N_20121,N_20204);
nand U20441 (N_20441,N_20185,N_20340);
xnor U20442 (N_20442,N_20200,N_20201);
nand U20443 (N_20443,N_20109,N_20301);
and U20444 (N_20444,N_20336,N_20349);
nand U20445 (N_20445,N_20291,N_20347);
and U20446 (N_20446,N_20159,N_20371);
and U20447 (N_20447,N_20228,N_20160);
nand U20448 (N_20448,N_20374,N_20149);
nor U20449 (N_20449,N_20394,N_20307);
or U20450 (N_20450,N_20203,N_20126);
or U20451 (N_20451,N_20208,N_20237);
nor U20452 (N_20452,N_20274,N_20164);
nor U20453 (N_20453,N_20272,N_20365);
and U20454 (N_20454,N_20192,N_20358);
xor U20455 (N_20455,N_20361,N_20205);
nor U20456 (N_20456,N_20271,N_20106);
nor U20457 (N_20457,N_20238,N_20363);
xnor U20458 (N_20458,N_20137,N_20360);
or U20459 (N_20459,N_20233,N_20226);
xor U20460 (N_20460,N_20269,N_20264);
or U20461 (N_20461,N_20114,N_20311);
nand U20462 (N_20462,N_20211,N_20122);
nand U20463 (N_20463,N_20342,N_20247);
or U20464 (N_20464,N_20251,N_20215);
and U20465 (N_20465,N_20157,N_20357);
nor U20466 (N_20466,N_20193,N_20210);
and U20467 (N_20467,N_20136,N_20209);
or U20468 (N_20468,N_20183,N_20152);
nor U20469 (N_20469,N_20381,N_20231);
nor U20470 (N_20470,N_20213,N_20378);
nand U20471 (N_20471,N_20154,N_20356);
or U20472 (N_20472,N_20370,N_20286);
nand U20473 (N_20473,N_20306,N_20281);
and U20474 (N_20474,N_20294,N_20290);
and U20475 (N_20475,N_20304,N_20359);
nand U20476 (N_20476,N_20197,N_20260);
and U20477 (N_20477,N_20198,N_20326);
xnor U20478 (N_20478,N_20339,N_20375);
and U20479 (N_20479,N_20259,N_20181);
and U20480 (N_20480,N_20116,N_20399);
and U20481 (N_20481,N_20379,N_20162);
or U20482 (N_20482,N_20182,N_20111);
and U20483 (N_20483,N_20275,N_20270);
or U20484 (N_20484,N_20367,N_20191);
and U20485 (N_20485,N_20305,N_20362);
xor U20486 (N_20486,N_20135,N_20100);
and U20487 (N_20487,N_20267,N_20265);
and U20488 (N_20488,N_20190,N_20240);
nand U20489 (N_20489,N_20222,N_20392);
and U20490 (N_20490,N_20245,N_20262);
and U20491 (N_20491,N_20129,N_20391);
nand U20492 (N_20492,N_20216,N_20343);
xnor U20493 (N_20493,N_20125,N_20322);
or U20494 (N_20494,N_20199,N_20320);
nand U20495 (N_20495,N_20180,N_20187);
nor U20496 (N_20496,N_20334,N_20295);
nor U20497 (N_20497,N_20366,N_20188);
nand U20498 (N_20498,N_20171,N_20354);
nor U20499 (N_20499,N_20227,N_20297);
xor U20500 (N_20500,N_20289,N_20184);
nor U20501 (N_20501,N_20331,N_20223);
or U20502 (N_20502,N_20353,N_20351);
and U20503 (N_20503,N_20345,N_20234);
or U20504 (N_20504,N_20332,N_20253);
and U20505 (N_20505,N_20241,N_20384);
or U20506 (N_20506,N_20169,N_20246);
nand U20507 (N_20507,N_20279,N_20396);
and U20508 (N_20508,N_20344,N_20195);
and U20509 (N_20509,N_20364,N_20132);
and U20510 (N_20510,N_20314,N_20257);
and U20511 (N_20511,N_20298,N_20102);
and U20512 (N_20512,N_20255,N_20229);
or U20513 (N_20513,N_20153,N_20138);
or U20514 (N_20514,N_20283,N_20280);
or U20515 (N_20515,N_20258,N_20101);
nor U20516 (N_20516,N_20249,N_20150);
and U20517 (N_20517,N_20388,N_20212);
nor U20518 (N_20518,N_20327,N_20312);
nand U20519 (N_20519,N_20221,N_20296);
or U20520 (N_20520,N_20256,N_20176);
xor U20521 (N_20521,N_20214,N_20165);
xnor U20522 (N_20522,N_20335,N_20104);
nor U20523 (N_20523,N_20242,N_20163);
nand U20524 (N_20524,N_20292,N_20346);
or U20525 (N_20525,N_20337,N_20170);
and U20526 (N_20526,N_20151,N_20398);
nand U20527 (N_20527,N_20386,N_20380);
nand U20528 (N_20528,N_20224,N_20207);
nor U20529 (N_20529,N_20252,N_20309);
nand U20530 (N_20530,N_20319,N_20284);
xor U20531 (N_20531,N_20124,N_20254);
or U20532 (N_20532,N_20393,N_20236);
nand U20533 (N_20533,N_20206,N_20119);
nor U20534 (N_20534,N_20179,N_20308);
nor U20535 (N_20535,N_20194,N_20390);
or U20536 (N_20536,N_20243,N_20350);
xnor U20537 (N_20537,N_20158,N_20263);
or U20538 (N_20538,N_20189,N_20117);
xor U20539 (N_20539,N_20155,N_20186);
and U20540 (N_20540,N_20127,N_20268);
or U20541 (N_20541,N_20373,N_20372);
and U20542 (N_20542,N_20140,N_20120);
and U20543 (N_20543,N_20333,N_20282);
nor U20544 (N_20544,N_20328,N_20261);
and U20545 (N_20545,N_20173,N_20230);
nand U20546 (N_20546,N_20113,N_20285);
nand U20547 (N_20547,N_20317,N_20387);
nand U20548 (N_20548,N_20287,N_20318);
or U20549 (N_20549,N_20105,N_20161);
or U20550 (N_20550,N_20150,N_20395);
xnor U20551 (N_20551,N_20247,N_20275);
and U20552 (N_20552,N_20349,N_20146);
and U20553 (N_20553,N_20395,N_20230);
nand U20554 (N_20554,N_20208,N_20212);
or U20555 (N_20555,N_20216,N_20266);
or U20556 (N_20556,N_20135,N_20365);
nand U20557 (N_20557,N_20114,N_20245);
nand U20558 (N_20558,N_20244,N_20275);
nand U20559 (N_20559,N_20380,N_20207);
and U20560 (N_20560,N_20189,N_20147);
or U20561 (N_20561,N_20190,N_20262);
nand U20562 (N_20562,N_20354,N_20382);
nand U20563 (N_20563,N_20167,N_20141);
xor U20564 (N_20564,N_20222,N_20238);
nand U20565 (N_20565,N_20399,N_20308);
or U20566 (N_20566,N_20310,N_20227);
nor U20567 (N_20567,N_20319,N_20360);
or U20568 (N_20568,N_20397,N_20301);
xor U20569 (N_20569,N_20189,N_20343);
xor U20570 (N_20570,N_20163,N_20259);
nand U20571 (N_20571,N_20290,N_20397);
nor U20572 (N_20572,N_20105,N_20173);
and U20573 (N_20573,N_20277,N_20255);
nor U20574 (N_20574,N_20244,N_20329);
nor U20575 (N_20575,N_20164,N_20314);
or U20576 (N_20576,N_20362,N_20178);
or U20577 (N_20577,N_20300,N_20379);
nand U20578 (N_20578,N_20329,N_20192);
xnor U20579 (N_20579,N_20327,N_20335);
nand U20580 (N_20580,N_20320,N_20302);
nor U20581 (N_20581,N_20165,N_20260);
and U20582 (N_20582,N_20286,N_20234);
nand U20583 (N_20583,N_20249,N_20361);
or U20584 (N_20584,N_20138,N_20166);
and U20585 (N_20585,N_20311,N_20221);
and U20586 (N_20586,N_20261,N_20370);
and U20587 (N_20587,N_20122,N_20249);
and U20588 (N_20588,N_20342,N_20250);
xor U20589 (N_20589,N_20185,N_20162);
nor U20590 (N_20590,N_20178,N_20230);
or U20591 (N_20591,N_20321,N_20178);
or U20592 (N_20592,N_20134,N_20225);
or U20593 (N_20593,N_20377,N_20125);
or U20594 (N_20594,N_20298,N_20181);
nand U20595 (N_20595,N_20136,N_20298);
and U20596 (N_20596,N_20259,N_20396);
xnor U20597 (N_20597,N_20357,N_20214);
or U20598 (N_20598,N_20162,N_20137);
xor U20599 (N_20599,N_20193,N_20100);
nand U20600 (N_20600,N_20100,N_20215);
and U20601 (N_20601,N_20383,N_20208);
xor U20602 (N_20602,N_20344,N_20220);
xor U20603 (N_20603,N_20161,N_20251);
and U20604 (N_20604,N_20390,N_20338);
nand U20605 (N_20605,N_20324,N_20302);
nand U20606 (N_20606,N_20226,N_20335);
and U20607 (N_20607,N_20123,N_20394);
nand U20608 (N_20608,N_20127,N_20182);
xnor U20609 (N_20609,N_20388,N_20140);
and U20610 (N_20610,N_20222,N_20371);
and U20611 (N_20611,N_20365,N_20201);
or U20612 (N_20612,N_20163,N_20299);
nor U20613 (N_20613,N_20267,N_20238);
and U20614 (N_20614,N_20161,N_20143);
or U20615 (N_20615,N_20221,N_20399);
xnor U20616 (N_20616,N_20207,N_20154);
or U20617 (N_20617,N_20106,N_20118);
or U20618 (N_20618,N_20151,N_20325);
and U20619 (N_20619,N_20135,N_20360);
xnor U20620 (N_20620,N_20301,N_20376);
nand U20621 (N_20621,N_20258,N_20360);
or U20622 (N_20622,N_20258,N_20154);
xor U20623 (N_20623,N_20178,N_20302);
xor U20624 (N_20624,N_20152,N_20241);
and U20625 (N_20625,N_20223,N_20125);
and U20626 (N_20626,N_20123,N_20372);
nor U20627 (N_20627,N_20261,N_20357);
or U20628 (N_20628,N_20112,N_20320);
nor U20629 (N_20629,N_20242,N_20245);
nor U20630 (N_20630,N_20230,N_20171);
nor U20631 (N_20631,N_20110,N_20284);
or U20632 (N_20632,N_20314,N_20376);
or U20633 (N_20633,N_20337,N_20220);
or U20634 (N_20634,N_20130,N_20333);
or U20635 (N_20635,N_20357,N_20243);
nor U20636 (N_20636,N_20356,N_20176);
xor U20637 (N_20637,N_20153,N_20189);
nand U20638 (N_20638,N_20149,N_20396);
or U20639 (N_20639,N_20378,N_20139);
or U20640 (N_20640,N_20237,N_20164);
or U20641 (N_20641,N_20374,N_20321);
nand U20642 (N_20642,N_20280,N_20285);
and U20643 (N_20643,N_20397,N_20183);
or U20644 (N_20644,N_20372,N_20176);
nand U20645 (N_20645,N_20228,N_20184);
nand U20646 (N_20646,N_20260,N_20155);
nand U20647 (N_20647,N_20260,N_20378);
and U20648 (N_20648,N_20210,N_20397);
nor U20649 (N_20649,N_20208,N_20342);
and U20650 (N_20650,N_20267,N_20222);
nand U20651 (N_20651,N_20285,N_20260);
xor U20652 (N_20652,N_20386,N_20249);
or U20653 (N_20653,N_20251,N_20378);
nand U20654 (N_20654,N_20356,N_20160);
xor U20655 (N_20655,N_20316,N_20251);
and U20656 (N_20656,N_20104,N_20196);
xor U20657 (N_20657,N_20277,N_20299);
xnor U20658 (N_20658,N_20344,N_20317);
xor U20659 (N_20659,N_20102,N_20264);
or U20660 (N_20660,N_20301,N_20270);
xnor U20661 (N_20661,N_20255,N_20181);
nor U20662 (N_20662,N_20343,N_20269);
and U20663 (N_20663,N_20383,N_20175);
and U20664 (N_20664,N_20231,N_20275);
and U20665 (N_20665,N_20262,N_20260);
or U20666 (N_20666,N_20283,N_20183);
xnor U20667 (N_20667,N_20224,N_20276);
nor U20668 (N_20668,N_20351,N_20242);
nor U20669 (N_20669,N_20338,N_20272);
nor U20670 (N_20670,N_20290,N_20193);
and U20671 (N_20671,N_20330,N_20149);
xnor U20672 (N_20672,N_20300,N_20370);
nor U20673 (N_20673,N_20290,N_20182);
nand U20674 (N_20674,N_20114,N_20220);
and U20675 (N_20675,N_20321,N_20163);
or U20676 (N_20676,N_20197,N_20370);
nor U20677 (N_20677,N_20263,N_20253);
and U20678 (N_20678,N_20396,N_20235);
xnor U20679 (N_20679,N_20234,N_20369);
or U20680 (N_20680,N_20110,N_20379);
or U20681 (N_20681,N_20152,N_20126);
or U20682 (N_20682,N_20129,N_20254);
and U20683 (N_20683,N_20358,N_20185);
nor U20684 (N_20684,N_20308,N_20280);
or U20685 (N_20685,N_20156,N_20396);
and U20686 (N_20686,N_20341,N_20113);
and U20687 (N_20687,N_20183,N_20166);
nor U20688 (N_20688,N_20226,N_20163);
and U20689 (N_20689,N_20116,N_20128);
and U20690 (N_20690,N_20151,N_20259);
nor U20691 (N_20691,N_20116,N_20266);
nand U20692 (N_20692,N_20316,N_20199);
or U20693 (N_20693,N_20339,N_20192);
nor U20694 (N_20694,N_20258,N_20277);
or U20695 (N_20695,N_20336,N_20170);
or U20696 (N_20696,N_20129,N_20131);
nor U20697 (N_20697,N_20115,N_20232);
or U20698 (N_20698,N_20299,N_20256);
xnor U20699 (N_20699,N_20171,N_20373);
or U20700 (N_20700,N_20444,N_20584);
nor U20701 (N_20701,N_20557,N_20497);
and U20702 (N_20702,N_20524,N_20676);
or U20703 (N_20703,N_20543,N_20457);
or U20704 (N_20704,N_20544,N_20468);
xnor U20705 (N_20705,N_20423,N_20510);
and U20706 (N_20706,N_20669,N_20417);
or U20707 (N_20707,N_20507,N_20445);
and U20708 (N_20708,N_20685,N_20469);
xnor U20709 (N_20709,N_20491,N_20449);
or U20710 (N_20710,N_20661,N_20547);
and U20711 (N_20711,N_20474,N_20562);
or U20712 (N_20712,N_20473,N_20634);
or U20713 (N_20713,N_20617,N_20426);
and U20714 (N_20714,N_20521,N_20421);
or U20715 (N_20715,N_20574,N_20528);
and U20716 (N_20716,N_20662,N_20682);
xor U20717 (N_20717,N_20680,N_20658);
nand U20718 (N_20718,N_20501,N_20597);
nor U20719 (N_20719,N_20433,N_20533);
or U20720 (N_20720,N_20509,N_20460);
nor U20721 (N_20721,N_20601,N_20690);
nor U20722 (N_20722,N_20465,N_20570);
nand U20723 (N_20723,N_20422,N_20590);
nand U20724 (N_20724,N_20477,N_20493);
and U20725 (N_20725,N_20630,N_20506);
nor U20726 (N_20726,N_20625,N_20560);
nor U20727 (N_20727,N_20627,N_20539);
and U20728 (N_20728,N_20600,N_20613);
nand U20729 (N_20729,N_20434,N_20559);
xnor U20730 (N_20730,N_20698,N_20548);
nand U20731 (N_20731,N_20579,N_20646);
and U20732 (N_20732,N_20565,N_20499);
nand U20733 (N_20733,N_20576,N_20692);
and U20734 (N_20734,N_20448,N_20500);
nor U20735 (N_20735,N_20492,N_20435);
and U20736 (N_20736,N_20631,N_20575);
or U20737 (N_20737,N_20628,N_20512);
xor U20738 (N_20738,N_20404,N_20656);
nand U20739 (N_20739,N_20487,N_20644);
xnor U20740 (N_20740,N_20667,N_20619);
nor U20741 (N_20741,N_20450,N_20593);
and U20742 (N_20742,N_20456,N_20504);
nor U20743 (N_20743,N_20623,N_20503);
and U20744 (N_20744,N_20502,N_20581);
and U20745 (N_20745,N_20616,N_20564);
nand U20746 (N_20746,N_20639,N_20679);
or U20747 (N_20747,N_20535,N_20563);
or U20748 (N_20748,N_20516,N_20476);
or U20749 (N_20749,N_20572,N_20606);
or U20750 (N_20750,N_20602,N_20546);
nor U20751 (N_20751,N_20532,N_20540);
and U20752 (N_20752,N_20596,N_20446);
xor U20753 (N_20753,N_20462,N_20478);
xnor U20754 (N_20754,N_20519,N_20635);
or U20755 (N_20755,N_20678,N_20674);
nand U20756 (N_20756,N_20459,N_20413);
xor U20757 (N_20757,N_20580,N_20489);
nor U20758 (N_20758,N_20551,N_20490);
or U20759 (N_20759,N_20406,N_20451);
xnor U20760 (N_20760,N_20699,N_20420);
xnor U20761 (N_20761,N_20569,N_20466);
nand U20762 (N_20762,N_20441,N_20675);
xor U20763 (N_20763,N_20668,N_20649);
nor U20764 (N_20764,N_20587,N_20481);
nand U20765 (N_20765,N_20607,N_20571);
and U20766 (N_20766,N_20670,N_20643);
and U20767 (N_20767,N_20431,N_20647);
nand U20768 (N_20768,N_20483,N_20472);
nand U20769 (N_20769,N_20482,N_20498);
nor U20770 (N_20770,N_20505,N_20583);
nand U20771 (N_20771,N_20517,N_20645);
nand U20772 (N_20772,N_20652,N_20427);
xnor U20773 (N_20773,N_20523,N_20626);
and U20774 (N_20774,N_20555,N_20620);
and U20775 (N_20775,N_20642,N_20567);
or U20776 (N_20776,N_20556,N_20454);
xor U20777 (N_20777,N_20479,N_20402);
or U20778 (N_20778,N_20621,N_20447);
or U20779 (N_20779,N_20530,N_20470);
and U20780 (N_20780,N_20688,N_20419);
nor U20781 (N_20781,N_20640,N_20424);
nor U20782 (N_20782,N_20654,N_20592);
nor U20783 (N_20783,N_20693,N_20561);
or U20784 (N_20784,N_20558,N_20549);
nand U20785 (N_20785,N_20467,N_20418);
xnor U20786 (N_20786,N_20629,N_20513);
or U20787 (N_20787,N_20614,N_20536);
and U20788 (N_20788,N_20514,N_20494);
nor U20789 (N_20789,N_20508,N_20538);
nand U20790 (N_20790,N_20541,N_20485);
xnor U20791 (N_20791,N_20672,N_20552);
and U20792 (N_20792,N_20610,N_20415);
and U20793 (N_20793,N_20689,N_20636);
nand U20794 (N_20794,N_20464,N_20573);
or U20795 (N_20795,N_20615,N_20432);
nand U20796 (N_20796,N_20648,N_20566);
or U20797 (N_20797,N_20577,N_20405);
or U20798 (N_20798,N_20442,N_20624);
or U20799 (N_20799,N_20681,N_20683);
or U20800 (N_20800,N_20458,N_20400);
nor U20801 (N_20801,N_20591,N_20438);
and U20802 (N_20802,N_20401,N_20641);
nand U20803 (N_20803,N_20436,N_20653);
and U20804 (N_20804,N_20638,N_20550);
and U20805 (N_20805,N_20463,N_20582);
xnor U20806 (N_20806,N_20537,N_20527);
nor U20807 (N_20807,N_20515,N_20443);
nand U20808 (N_20808,N_20429,N_20598);
and U20809 (N_20809,N_20471,N_20612);
nor U20810 (N_20810,N_20664,N_20694);
or U20811 (N_20811,N_20655,N_20665);
and U20812 (N_20812,N_20439,N_20531);
or U20813 (N_20813,N_20618,N_20659);
nand U20814 (N_20814,N_20409,N_20452);
nand U20815 (N_20815,N_20430,N_20486);
or U20816 (N_20816,N_20496,N_20604);
nand U20817 (N_20817,N_20633,N_20554);
nand U20818 (N_20818,N_20578,N_20608);
and U20819 (N_20819,N_20440,N_20522);
or U20820 (N_20820,N_20589,N_20545);
or U20821 (N_20821,N_20637,N_20416);
nand U20822 (N_20822,N_20553,N_20599);
nand U20823 (N_20823,N_20650,N_20412);
nand U20824 (N_20824,N_20594,N_20525);
or U20825 (N_20825,N_20526,N_20696);
and U20826 (N_20826,N_20407,N_20585);
or U20827 (N_20827,N_20603,N_20632);
or U20828 (N_20828,N_20660,N_20410);
or U20829 (N_20829,N_20488,N_20437);
or U20830 (N_20830,N_20691,N_20414);
nand U20831 (N_20831,N_20495,N_20666);
nor U20832 (N_20832,N_20511,N_20673);
xnor U20833 (N_20833,N_20697,N_20687);
or U20834 (N_20834,N_20542,N_20403);
and U20835 (N_20835,N_20671,N_20605);
xnor U20836 (N_20836,N_20611,N_20484);
and U20837 (N_20837,N_20518,N_20686);
xor U20838 (N_20838,N_20657,N_20408);
and U20839 (N_20839,N_20595,N_20651);
nand U20840 (N_20840,N_20695,N_20411);
nand U20841 (N_20841,N_20461,N_20588);
or U20842 (N_20842,N_20622,N_20534);
nand U20843 (N_20843,N_20529,N_20453);
xor U20844 (N_20844,N_20684,N_20609);
nor U20845 (N_20845,N_20425,N_20586);
or U20846 (N_20846,N_20455,N_20677);
and U20847 (N_20847,N_20480,N_20475);
xnor U20848 (N_20848,N_20663,N_20428);
and U20849 (N_20849,N_20568,N_20520);
and U20850 (N_20850,N_20402,N_20442);
nor U20851 (N_20851,N_20609,N_20629);
nand U20852 (N_20852,N_20621,N_20674);
xor U20853 (N_20853,N_20680,N_20607);
nor U20854 (N_20854,N_20628,N_20692);
or U20855 (N_20855,N_20643,N_20459);
or U20856 (N_20856,N_20570,N_20548);
and U20857 (N_20857,N_20429,N_20664);
and U20858 (N_20858,N_20549,N_20414);
or U20859 (N_20859,N_20461,N_20682);
nand U20860 (N_20860,N_20476,N_20416);
nor U20861 (N_20861,N_20535,N_20687);
nand U20862 (N_20862,N_20624,N_20645);
nand U20863 (N_20863,N_20498,N_20480);
xor U20864 (N_20864,N_20557,N_20498);
nand U20865 (N_20865,N_20666,N_20436);
nand U20866 (N_20866,N_20439,N_20604);
nand U20867 (N_20867,N_20448,N_20438);
xor U20868 (N_20868,N_20643,N_20409);
nand U20869 (N_20869,N_20634,N_20694);
xnor U20870 (N_20870,N_20649,N_20513);
or U20871 (N_20871,N_20564,N_20486);
xor U20872 (N_20872,N_20609,N_20513);
and U20873 (N_20873,N_20619,N_20439);
or U20874 (N_20874,N_20606,N_20549);
and U20875 (N_20875,N_20439,N_20668);
nand U20876 (N_20876,N_20499,N_20537);
xnor U20877 (N_20877,N_20669,N_20432);
nand U20878 (N_20878,N_20611,N_20487);
nand U20879 (N_20879,N_20601,N_20427);
nand U20880 (N_20880,N_20616,N_20458);
and U20881 (N_20881,N_20597,N_20585);
and U20882 (N_20882,N_20405,N_20517);
xor U20883 (N_20883,N_20475,N_20571);
or U20884 (N_20884,N_20560,N_20516);
xor U20885 (N_20885,N_20630,N_20520);
or U20886 (N_20886,N_20699,N_20666);
xnor U20887 (N_20887,N_20560,N_20577);
and U20888 (N_20888,N_20407,N_20638);
nor U20889 (N_20889,N_20607,N_20545);
xnor U20890 (N_20890,N_20437,N_20650);
nor U20891 (N_20891,N_20480,N_20597);
nand U20892 (N_20892,N_20473,N_20654);
and U20893 (N_20893,N_20455,N_20648);
nand U20894 (N_20894,N_20475,N_20565);
and U20895 (N_20895,N_20636,N_20474);
xor U20896 (N_20896,N_20621,N_20677);
nand U20897 (N_20897,N_20445,N_20682);
or U20898 (N_20898,N_20548,N_20697);
or U20899 (N_20899,N_20662,N_20545);
nor U20900 (N_20900,N_20433,N_20542);
nand U20901 (N_20901,N_20517,N_20430);
or U20902 (N_20902,N_20405,N_20447);
or U20903 (N_20903,N_20629,N_20684);
and U20904 (N_20904,N_20405,N_20672);
nand U20905 (N_20905,N_20487,N_20514);
nand U20906 (N_20906,N_20506,N_20414);
xnor U20907 (N_20907,N_20528,N_20515);
or U20908 (N_20908,N_20444,N_20616);
nor U20909 (N_20909,N_20444,N_20476);
xnor U20910 (N_20910,N_20424,N_20698);
and U20911 (N_20911,N_20477,N_20596);
xor U20912 (N_20912,N_20552,N_20414);
and U20913 (N_20913,N_20520,N_20579);
or U20914 (N_20914,N_20478,N_20604);
and U20915 (N_20915,N_20655,N_20674);
nand U20916 (N_20916,N_20556,N_20697);
and U20917 (N_20917,N_20483,N_20506);
nor U20918 (N_20918,N_20517,N_20577);
or U20919 (N_20919,N_20548,N_20533);
and U20920 (N_20920,N_20607,N_20543);
or U20921 (N_20921,N_20512,N_20578);
nor U20922 (N_20922,N_20679,N_20462);
xor U20923 (N_20923,N_20694,N_20472);
nand U20924 (N_20924,N_20655,N_20589);
xnor U20925 (N_20925,N_20615,N_20531);
nor U20926 (N_20926,N_20606,N_20628);
and U20927 (N_20927,N_20682,N_20608);
and U20928 (N_20928,N_20676,N_20663);
and U20929 (N_20929,N_20409,N_20639);
nor U20930 (N_20930,N_20595,N_20460);
xor U20931 (N_20931,N_20639,N_20508);
and U20932 (N_20932,N_20614,N_20479);
nand U20933 (N_20933,N_20690,N_20678);
and U20934 (N_20934,N_20514,N_20496);
nand U20935 (N_20935,N_20485,N_20472);
or U20936 (N_20936,N_20415,N_20526);
xnor U20937 (N_20937,N_20433,N_20569);
nand U20938 (N_20938,N_20496,N_20530);
and U20939 (N_20939,N_20675,N_20450);
or U20940 (N_20940,N_20439,N_20696);
xor U20941 (N_20941,N_20624,N_20427);
and U20942 (N_20942,N_20532,N_20511);
xnor U20943 (N_20943,N_20581,N_20548);
xor U20944 (N_20944,N_20571,N_20674);
or U20945 (N_20945,N_20676,N_20636);
or U20946 (N_20946,N_20490,N_20645);
and U20947 (N_20947,N_20545,N_20418);
xor U20948 (N_20948,N_20486,N_20586);
and U20949 (N_20949,N_20600,N_20449);
nand U20950 (N_20950,N_20463,N_20449);
and U20951 (N_20951,N_20493,N_20486);
nand U20952 (N_20952,N_20653,N_20512);
or U20953 (N_20953,N_20651,N_20407);
xor U20954 (N_20954,N_20529,N_20498);
xor U20955 (N_20955,N_20425,N_20487);
or U20956 (N_20956,N_20444,N_20606);
xor U20957 (N_20957,N_20566,N_20429);
or U20958 (N_20958,N_20450,N_20651);
and U20959 (N_20959,N_20446,N_20633);
nor U20960 (N_20960,N_20473,N_20515);
and U20961 (N_20961,N_20593,N_20662);
or U20962 (N_20962,N_20479,N_20491);
nor U20963 (N_20963,N_20404,N_20642);
xnor U20964 (N_20964,N_20473,N_20443);
nand U20965 (N_20965,N_20663,N_20660);
or U20966 (N_20966,N_20433,N_20628);
and U20967 (N_20967,N_20460,N_20468);
nor U20968 (N_20968,N_20548,N_20481);
and U20969 (N_20969,N_20687,N_20595);
nor U20970 (N_20970,N_20570,N_20554);
or U20971 (N_20971,N_20518,N_20533);
and U20972 (N_20972,N_20590,N_20401);
nor U20973 (N_20973,N_20655,N_20666);
nor U20974 (N_20974,N_20429,N_20630);
or U20975 (N_20975,N_20533,N_20531);
and U20976 (N_20976,N_20642,N_20670);
or U20977 (N_20977,N_20411,N_20434);
xnor U20978 (N_20978,N_20635,N_20673);
and U20979 (N_20979,N_20427,N_20694);
nand U20980 (N_20980,N_20566,N_20428);
xnor U20981 (N_20981,N_20592,N_20689);
xnor U20982 (N_20982,N_20686,N_20420);
nand U20983 (N_20983,N_20651,N_20658);
and U20984 (N_20984,N_20681,N_20475);
or U20985 (N_20985,N_20629,N_20491);
nand U20986 (N_20986,N_20458,N_20620);
nand U20987 (N_20987,N_20555,N_20475);
xnor U20988 (N_20988,N_20469,N_20408);
nor U20989 (N_20989,N_20546,N_20538);
nor U20990 (N_20990,N_20641,N_20500);
or U20991 (N_20991,N_20519,N_20416);
and U20992 (N_20992,N_20694,N_20558);
or U20993 (N_20993,N_20426,N_20481);
xor U20994 (N_20994,N_20550,N_20611);
xor U20995 (N_20995,N_20494,N_20546);
and U20996 (N_20996,N_20456,N_20410);
nand U20997 (N_20997,N_20648,N_20528);
and U20998 (N_20998,N_20541,N_20488);
nand U20999 (N_20999,N_20681,N_20449);
and U21000 (N_21000,N_20772,N_20864);
nand U21001 (N_21001,N_20958,N_20913);
nor U21002 (N_21002,N_20931,N_20823);
nand U21003 (N_21003,N_20767,N_20708);
nand U21004 (N_21004,N_20942,N_20833);
or U21005 (N_21005,N_20847,N_20905);
xor U21006 (N_21006,N_20946,N_20818);
and U21007 (N_21007,N_20828,N_20939);
and U21008 (N_21008,N_20790,N_20964);
and U21009 (N_21009,N_20992,N_20920);
xnor U21010 (N_21010,N_20716,N_20882);
nand U21011 (N_21011,N_20903,N_20901);
nand U21012 (N_21012,N_20706,N_20883);
xnor U21013 (N_21013,N_20921,N_20727);
or U21014 (N_21014,N_20947,N_20712);
xor U21015 (N_21015,N_20737,N_20938);
or U21016 (N_21016,N_20856,N_20777);
or U21017 (N_21017,N_20922,N_20820);
nor U21018 (N_21018,N_20956,N_20940);
or U21019 (N_21019,N_20733,N_20990);
nand U21020 (N_21020,N_20934,N_20861);
nand U21021 (N_21021,N_20775,N_20965);
xnor U21022 (N_21022,N_20951,N_20858);
or U21023 (N_21023,N_20899,N_20845);
xnor U21024 (N_21024,N_20766,N_20837);
xnor U21025 (N_21025,N_20738,N_20742);
xor U21026 (N_21026,N_20929,N_20937);
nand U21027 (N_21027,N_20853,N_20764);
xnor U21028 (N_21028,N_20840,N_20863);
nand U21029 (N_21029,N_20843,N_20980);
nor U21030 (N_21030,N_20898,N_20717);
and U21031 (N_21031,N_20709,N_20855);
nor U21032 (N_21032,N_20994,N_20746);
and U21033 (N_21033,N_20888,N_20740);
or U21034 (N_21034,N_20987,N_20978);
xnor U21035 (N_21035,N_20782,N_20897);
nand U21036 (N_21036,N_20741,N_20896);
xor U21037 (N_21037,N_20860,N_20735);
or U21038 (N_21038,N_20815,N_20752);
and U21039 (N_21039,N_20850,N_20874);
xor U21040 (N_21040,N_20841,N_20962);
nor U21041 (N_21041,N_20854,N_20989);
nor U21042 (N_21042,N_20731,N_20952);
nor U21043 (N_21043,N_20936,N_20801);
nor U21044 (N_21044,N_20813,N_20912);
and U21045 (N_21045,N_20832,N_20928);
or U21046 (N_21046,N_20759,N_20959);
and U21047 (N_21047,N_20814,N_20932);
or U21048 (N_21048,N_20799,N_20890);
and U21049 (N_21049,N_20982,N_20839);
and U21050 (N_21050,N_20793,N_20788);
nand U21051 (N_21051,N_20983,N_20852);
and U21052 (N_21052,N_20822,N_20809);
or U21053 (N_21053,N_20768,N_20779);
or U21054 (N_21054,N_20797,N_20902);
and U21055 (N_21055,N_20795,N_20900);
xnor U21056 (N_21056,N_20842,N_20804);
nor U21057 (N_21057,N_20872,N_20889);
nand U21058 (N_21058,N_20807,N_20953);
and U21059 (N_21059,N_20880,N_20873);
nor U21060 (N_21060,N_20784,N_20720);
nand U21061 (N_21061,N_20778,N_20836);
or U21062 (N_21062,N_20805,N_20957);
nand U21063 (N_21063,N_20857,N_20876);
or U21064 (N_21064,N_20995,N_20949);
nand U21065 (N_21065,N_20750,N_20985);
xor U21066 (N_21066,N_20714,N_20988);
nor U21067 (N_21067,N_20954,N_20713);
nor U21068 (N_21068,N_20948,N_20721);
nand U21069 (N_21069,N_20821,N_20844);
or U21070 (N_21070,N_20884,N_20803);
nor U21071 (N_21071,N_20838,N_20812);
nor U21072 (N_21072,N_20830,N_20894);
xor U21073 (N_21073,N_20925,N_20911);
xor U21074 (N_21074,N_20968,N_20941);
xnor U21075 (N_21075,N_20908,N_20751);
and U21076 (N_21076,N_20945,N_20825);
nand U21077 (N_21077,N_20966,N_20891);
and U21078 (N_21078,N_20715,N_20700);
nor U21079 (N_21079,N_20748,N_20736);
and U21080 (N_21080,N_20870,N_20927);
or U21081 (N_21081,N_20771,N_20950);
nand U21082 (N_21082,N_20878,N_20783);
or U21083 (N_21083,N_20917,N_20909);
and U21084 (N_21084,N_20986,N_20753);
xnor U21085 (N_21085,N_20892,N_20846);
or U21086 (N_21086,N_20745,N_20710);
and U21087 (N_21087,N_20919,N_20824);
xor U21088 (N_21088,N_20754,N_20749);
or U21089 (N_21089,N_20943,N_20722);
or U21090 (N_21090,N_20802,N_20904);
and U21091 (N_21091,N_20794,N_20976);
or U21092 (N_21092,N_20967,N_20791);
xnor U21093 (N_21093,N_20906,N_20895);
or U21094 (N_21094,N_20743,N_20955);
or U21095 (N_21095,N_20865,N_20819);
nor U21096 (N_21096,N_20868,N_20881);
nand U21097 (N_21097,N_20707,N_20762);
xnor U21098 (N_21098,N_20849,N_20998);
nand U21099 (N_21099,N_20765,N_20893);
nor U21100 (N_21100,N_20859,N_20918);
nand U21101 (N_21101,N_20826,N_20729);
and U21102 (N_21102,N_20773,N_20835);
nand U21103 (N_21103,N_20848,N_20792);
nand U21104 (N_21104,N_20725,N_20944);
nor U21105 (N_21105,N_20785,N_20798);
nand U21106 (N_21106,N_20973,N_20960);
nand U21107 (N_21107,N_20774,N_20997);
nand U21108 (N_21108,N_20879,N_20757);
and U21109 (N_21109,N_20730,N_20993);
nor U21110 (N_21110,N_20760,N_20703);
nand U21111 (N_21111,N_20974,N_20786);
nand U21112 (N_21112,N_20769,N_20963);
nand U21113 (N_21113,N_20796,N_20726);
nor U21114 (N_21114,N_20869,N_20755);
and U21115 (N_21115,N_20719,N_20728);
or U21116 (N_21116,N_20806,N_20744);
and U21117 (N_21117,N_20739,N_20977);
xnor U21118 (N_21118,N_20808,N_20885);
xnor U21119 (N_21119,N_20867,N_20810);
or U21120 (N_21120,N_20817,N_20776);
nor U21121 (N_21121,N_20981,N_20800);
nand U21122 (N_21122,N_20862,N_20770);
xnor U21123 (N_21123,N_20969,N_20789);
or U21124 (N_21124,N_20723,N_20984);
and U21125 (N_21125,N_20915,N_20831);
and U21126 (N_21126,N_20996,N_20875);
or U21127 (N_21127,N_20704,N_20702);
nand U21128 (N_21128,N_20761,N_20705);
nor U21129 (N_21129,N_20827,N_20907);
and U21130 (N_21130,N_20877,N_20734);
xnor U21131 (N_21131,N_20886,N_20756);
xnor U21132 (N_21132,N_20780,N_20758);
nand U21133 (N_21133,N_20711,N_20914);
nand U21134 (N_21134,N_20787,N_20871);
nor U21135 (N_21135,N_20834,N_20866);
nor U21136 (N_21136,N_20961,N_20935);
nor U21137 (N_21137,N_20732,N_20972);
or U21138 (N_21138,N_20975,N_20887);
and U21139 (N_21139,N_20910,N_20701);
nand U21140 (N_21140,N_20971,N_20718);
or U21141 (N_21141,N_20781,N_20923);
xnor U21142 (N_21142,N_20999,N_20811);
xnor U21143 (N_21143,N_20763,N_20851);
xnor U21144 (N_21144,N_20916,N_20724);
nand U21145 (N_21145,N_20816,N_20970);
nor U21146 (N_21146,N_20924,N_20930);
xnor U21147 (N_21147,N_20829,N_20979);
xnor U21148 (N_21148,N_20933,N_20926);
nor U21149 (N_21149,N_20747,N_20991);
nor U21150 (N_21150,N_20894,N_20827);
nand U21151 (N_21151,N_20835,N_20761);
nor U21152 (N_21152,N_20853,N_20936);
nand U21153 (N_21153,N_20724,N_20974);
nand U21154 (N_21154,N_20958,N_20886);
and U21155 (N_21155,N_20880,N_20885);
or U21156 (N_21156,N_20742,N_20973);
and U21157 (N_21157,N_20741,N_20956);
nand U21158 (N_21158,N_20802,N_20709);
xor U21159 (N_21159,N_20922,N_20918);
nor U21160 (N_21160,N_20796,N_20989);
and U21161 (N_21161,N_20758,N_20902);
nor U21162 (N_21162,N_20890,N_20711);
and U21163 (N_21163,N_20939,N_20989);
or U21164 (N_21164,N_20721,N_20828);
xnor U21165 (N_21165,N_20830,N_20777);
xor U21166 (N_21166,N_20945,N_20718);
nand U21167 (N_21167,N_20832,N_20775);
and U21168 (N_21168,N_20880,N_20817);
nor U21169 (N_21169,N_20802,N_20956);
or U21170 (N_21170,N_20952,N_20852);
nand U21171 (N_21171,N_20906,N_20882);
xnor U21172 (N_21172,N_20888,N_20704);
and U21173 (N_21173,N_20830,N_20992);
nand U21174 (N_21174,N_20940,N_20742);
nor U21175 (N_21175,N_20983,N_20938);
nor U21176 (N_21176,N_20899,N_20934);
nand U21177 (N_21177,N_20990,N_20851);
xor U21178 (N_21178,N_20825,N_20860);
nand U21179 (N_21179,N_20906,N_20987);
xnor U21180 (N_21180,N_20763,N_20732);
nor U21181 (N_21181,N_20991,N_20865);
xnor U21182 (N_21182,N_20789,N_20918);
or U21183 (N_21183,N_20734,N_20923);
or U21184 (N_21184,N_20701,N_20936);
nand U21185 (N_21185,N_20831,N_20754);
nor U21186 (N_21186,N_20965,N_20937);
and U21187 (N_21187,N_20889,N_20745);
nor U21188 (N_21188,N_20796,N_20949);
xnor U21189 (N_21189,N_20705,N_20716);
and U21190 (N_21190,N_20811,N_20731);
nor U21191 (N_21191,N_20732,N_20915);
nor U21192 (N_21192,N_20775,N_20870);
and U21193 (N_21193,N_20884,N_20933);
nand U21194 (N_21194,N_20888,N_20700);
and U21195 (N_21195,N_20764,N_20715);
and U21196 (N_21196,N_20793,N_20950);
nand U21197 (N_21197,N_20967,N_20781);
xor U21198 (N_21198,N_20938,N_20926);
xnor U21199 (N_21199,N_20998,N_20808);
and U21200 (N_21200,N_20843,N_20724);
xnor U21201 (N_21201,N_20804,N_20975);
and U21202 (N_21202,N_20728,N_20802);
nand U21203 (N_21203,N_20955,N_20924);
nor U21204 (N_21204,N_20863,N_20778);
nor U21205 (N_21205,N_20832,N_20892);
and U21206 (N_21206,N_20930,N_20846);
nand U21207 (N_21207,N_20863,N_20914);
nor U21208 (N_21208,N_20700,N_20843);
xor U21209 (N_21209,N_20937,N_20866);
xor U21210 (N_21210,N_20718,N_20746);
nor U21211 (N_21211,N_20999,N_20786);
or U21212 (N_21212,N_20920,N_20792);
nor U21213 (N_21213,N_20761,N_20771);
and U21214 (N_21214,N_20877,N_20708);
nor U21215 (N_21215,N_20983,N_20716);
and U21216 (N_21216,N_20873,N_20701);
or U21217 (N_21217,N_20946,N_20773);
xor U21218 (N_21218,N_20984,N_20806);
xor U21219 (N_21219,N_20845,N_20751);
or U21220 (N_21220,N_20832,N_20816);
and U21221 (N_21221,N_20939,N_20752);
or U21222 (N_21222,N_20936,N_20878);
nand U21223 (N_21223,N_20731,N_20981);
or U21224 (N_21224,N_20929,N_20720);
xnor U21225 (N_21225,N_20927,N_20824);
nor U21226 (N_21226,N_20960,N_20745);
nand U21227 (N_21227,N_20869,N_20924);
nor U21228 (N_21228,N_20963,N_20928);
nor U21229 (N_21229,N_20751,N_20746);
and U21230 (N_21230,N_20937,N_20804);
nand U21231 (N_21231,N_20887,N_20919);
and U21232 (N_21232,N_20747,N_20944);
and U21233 (N_21233,N_20864,N_20952);
nor U21234 (N_21234,N_20978,N_20786);
and U21235 (N_21235,N_20700,N_20731);
and U21236 (N_21236,N_20920,N_20919);
xnor U21237 (N_21237,N_20841,N_20939);
and U21238 (N_21238,N_20718,N_20969);
nand U21239 (N_21239,N_20852,N_20865);
xnor U21240 (N_21240,N_20816,N_20888);
and U21241 (N_21241,N_20894,N_20983);
or U21242 (N_21242,N_20732,N_20978);
nor U21243 (N_21243,N_20754,N_20740);
or U21244 (N_21244,N_20985,N_20924);
or U21245 (N_21245,N_20835,N_20749);
nor U21246 (N_21246,N_20790,N_20841);
or U21247 (N_21247,N_20876,N_20956);
xnor U21248 (N_21248,N_20779,N_20763);
xnor U21249 (N_21249,N_20847,N_20737);
xor U21250 (N_21250,N_20732,N_20953);
nand U21251 (N_21251,N_20718,N_20763);
xor U21252 (N_21252,N_20997,N_20765);
nor U21253 (N_21253,N_20836,N_20950);
nor U21254 (N_21254,N_20848,N_20827);
xnor U21255 (N_21255,N_20860,N_20822);
nand U21256 (N_21256,N_20924,N_20833);
nor U21257 (N_21257,N_20762,N_20722);
nand U21258 (N_21258,N_20920,N_20758);
xor U21259 (N_21259,N_20717,N_20988);
nand U21260 (N_21260,N_20760,N_20960);
or U21261 (N_21261,N_20700,N_20951);
xnor U21262 (N_21262,N_20772,N_20867);
and U21263 (N_21263,N_20773,N_20903);
and U21264 (N_21264,N_20923,N_20729);
xnor U21265 (N_21265,N_20826,N_20876);
nand U21266 (N_21266,N_20992,N_20922);
and U21267 (N_21267,N_20780,N_20995);
xor U21268 (N_21268,N_20897,N_20829);
nor U21269 (N_21269,N_20770,N_20980);
nor U21270 (N_21270,N_20735,N_20733);
nor U21271 (N_21271,N_20788,N_20868);
nor U21272 (N_21272,N_20704,N_20718);
nand U21273 (N_21273,N_20805,N_20806);
nand U21274 (N_21274,N_20965,N_20885);
or U21275 (N_21275,N_20944,N_20938);
or U21276 (N_21276,N_20788,N_20777);
or U21277 (N_21277,N_20988,N_20704);
nand U21278 (N_21278,N_20878,N_20724);
nor U21279 (N_21279,N_20858,N_20851);
nand U21280 (N_21280,N_20941,N_20926);
and U21281 (N_21281,N_20707,N_20844);
or U21282 (N_21282,N_20848,N_20861);
and U21283 (N_21283,N_20842,N_20776);
and U21284 (N_21284,N_20712,N_20792);
nand U21285 (N_21285,N_20772,N_20910);
and U21286 (N_21286,N_20849,N_20791);
nand U21287 (N_21287,N_20839,N_20827);
nand U21288 (N_21288,N_20923,N_20975);
nand U21289 (N_21289,N_20920,N_20908);
xor U21290 (N_21290,N_20877,N_20836);
and U21291 (N_21291,N_20827,N_20934);
nor U21292 (N_21292,N_20980,N_20853);
nor U21293 (N_21293,N_20737,N_20931);
xnor U21294 (N_21294,N_20785,N_20894);
nor U21295 (N_21295,N_20867,N_20925);
nand U21296 (N_21296,N_20922,N_20746);
and U21297 (N_21297,N_20809,N_20710);
nor U21298 (N_21298,N_20967,N_20977);
nand U21299 (N_21299,N_20715,N_20977);
nor U21300 (N_21300,N_21064,N_21043);
or U21301 (N_21301,N_21163,N_21146);
nor U21302 (N_21302,N_21049,N_21248);
and U21303 (N_21303,N_21228,N_21050);
and U21304 (N_21304,N_21100,N_21193);
and U21305 (N_21305,N_21125,N_21135);
or U21306 (N_21306,N_21218,N_21183);
or U21307 (N_21307,N_21151,N_21212);
nand U21308 (N_21308,N_21029,N_21264);
xnor U21309 (N_21309,N_21251,N_21214);
xor U21310 (N_21310,N_21116,N_21224);
or U21311 (N_21311,N_21281,N_21095);
nor U21312 (N_21312,N_21046,N_21237);
or U21313 (N_21313,N_21232,N_21053);
or U21314 (N_21314,N_21065,N_21241);
or U21315 (N_21315,N_21081,N_21140);
or U21316 (N_21316,N_21036,N_21270);
xor U21317 (N_21317,N_21035,N_21139);
xor U21318 (N_21318,N_21058,N_21013);
or U21319 (N_21319,N_21216,N_21072);
and U21320 (N_21320,N_21266,N_21278);
xor U21321 (N_21321,N_21179,N_21079);
or U21322 (N_21322,N_21026,N_21002);
xnor U21323 (N_21323,N_21090,N_21202);
nand U21324 (N_21324,N_21048,N_21108);
nor U21325 (N_21325,N_21290,N_21115);
nand U21326 (N_21326,N_21088,N_21102);
nor U21327 (N_21327,N_21205,N_21189);
or U21328 (N_21328,N_21167,N_21020);
nand U21329 (N_21329,N_21153,N_21156);
or U21330 (N_21330,N_21119,N_21110);
nor U21331 (N_21331,N_21068,N_21136);
or U21332 (N_21332,N_21015,N_21235);
or U21333 (N_21333,N_21221,N_21215);
nor U21334 (N_21334,N_21234,N_21148);
and U21335 (N_21335,N_21273,N_21150);
or U21336 (N_21336,N_21143,N_21096);
or U21337 (N_21337,N_21184,N_21052);
and U21338 (N_21338,N_21253,N_21134);
nand U21339 (N_21339,N_21256,N_21129);
xnor U21340 (N_21340,N_21120,N_21132);
and U21341 (N_21341,N_21194,N_21155);
nor U21342 (N_21342,N_21098,N_21008);
and U21343 (N_21343,N_21297,N_21169);
or U21344 (N_21344,N_21001,N_21229);
xor U21345 (N_21345,N_21201,N_21094);
xor U21346 (N_21346,N_21299,N_21041);
and U21347 (N_21347,N_21254,N_21018);
or U21348 (N_21348,N_21074,N_21076);
or U21349 (N_21349,N_21004,N_21069);
nor U21350 (N_21350,N_21240,N_21282);
or U21351 (N_21351,N_21027,N_21011);
nor U21352 (N_21352,N_21023,N_21181);
nor U21353 (N_21353,N_21138,N_21249);
and U21354 (N_21354,N_21044,N_21097);
and U21355 (N_21355,N_21296,N_21230);
xor U21356 (N_21356,N_21159,N_21010);
nand U21357 (N_21357,N_21186,N_21158);
or U21358 (N_21358,N_21293,N_21066);
or U21359 (N_21359,N_21091,N_21113);
nand U21360 (N_21360,N_21226,N_21089);
nand U21361 (N_21361,N_21219,N_21261);
xnor U21362 (N_21362,N_21280,N_21047);
nand U21363 (N_21363,N_21103,N_21170);
xnor U21364 (N_21364,N_21128,N_21242);
or U21365 (N_21365,N_21277,N_21187);
xnor U21366 (N_21366,N_21268,N_21217);
nor U21367 (N_21367,N_21177,N_21203);
nand U21368 (N_21368,N_21207,N_21198);
nor U21369 (N_21369,N_21284,N_21080);
nor U21370 (N_21370,N_21021,N_21180);
or U21371 (N_21371,N_21222,N_21298);
xnor U21372 (N_21372,N_21121,N_21022);
and U21373 (N_21373,N_21259,N_21061);
or U21374 (N_21374,N_21040,N_21037);
or U21375 (N_21375,N_21060,N_21250);
nand U21376 (N_21376,N_21006,N_21275);
nor U21377 (N_21377,N_21016,N_21105);
nor U21378 (N_21378,N_21019,N_21123);
nor U21379 (N_21379,N_21051,N_21032);
nor U21380 (N_21380,N_21034,N_21038);
xor U21381 (N_21381,N_21124,N_21126);
or U21382 (N_21382,N_21204,N_21272);
xor U21383 (N_21383,N_21276,N_21244);
or U21384 (N_21384,N_21283,N_21109);
or U21385 (N_21385,N_21185,N_21057);
xnor U21386 (N_21386,N_21030,N_21257);
nor U21387 (N_21387,N_21267,N_21028);
xnor U21388 (N_21388,N_21233,N_21182);
xor U21389 (N_21389,N_21070,N_21208);
and U21390 (N_21390,N_21117,N_21085);
or U21391 (N_21391,N_21188,N_21130);
nor U21392 (N_21392,N_21099,N_21114);
xnor U21393 (N_21393,N_21122,N_21104);
or U21394 (N_21394,N_21252,N_21292);
nand U21395 (N_21395,N_21017,N_21107);
nand U21396 (N_21396,N_21174,N_21192);
nand U21397 (N_21397,N_21054,N_21279);
or U21398 (N_21398,N_21166,N_21025);
nand U21399 (N_21399,N_21291,N_21031);
nand U21400 (N_21400,N_21213,N_21000);
or U21401 (N_21401,N_21196,N_21231);
nor U21402 (N_21402,N_21012,N_21220);
nand U21403 (N_21403,N_21144,N_21118);
xor U21404 (N_21404,N_21246,N_21199);
xor U21405 (N_21405,N_21077,N_21172);
xor U21406 (N_21406,N_21112,N_21161);
nor U21407 (N_21407,N_21045,N_21178);
or U21408 (N_21408,N_21067,N_21262);
or U21409 (N_21409,N_21271,N_21239);
nand U21410 (N_21410,N_21210,N_21195);
or U21411 (N_21411,N_21033,N_21288);
nor U21412 (N_21412,N_21269,N_21005);
nor U21413 (N_21413,N_21175,N_21131);
or U21414 (N_21414,N_21223,N_21236);
or U21415 (N_21415,N_21071,N_21092);
nand U21416 (N_21416,N_21168,N_21247);
xnor U21417 (N_21417,N_21075,N_21294);
nand U21418 (N_21418,N_21141,N_21062);
or U21419 (N_21419,N_21206,N_21289);
nand U21420 (N_21420,N_21164,N_21225);
xnor U21421 (N_21421,N_21211,N_21106);
or U21422 (N_21422,N_21014,N_21295);
or U21423 (N_21423,N_21173,N_21127);
and U21424 (N_21424,N_21083,N_21243);
nor U21425 (N_21425,N_21137,N_21165);
nor U21426 (N_21426,N_21154,N_21286);
and U21427 (N_21427,N_21078,N_21007);
xnor U21428 (N_21428,N_21260,N_21101);
xnor U21429 (N_21429,N_21059,N_21171);
or U21430 (N_21430,N_21227,N_21009);
nand U21431 (N_21431,N_21056,N_21149);
nor U21432 (N_21432,N_21082,N_21063);
nor U21433 (N_21433,N_21039,N_21209);
and U21434 (N_21434,N_21162,N_21160);
nand U21435 (N_21435,N_21258,N_21190);
nor U21436 (N_21436,N_21274,N_21073);
or U21437 (N_21437,N_21093,N_21263);
nor U21438 (N_21438,N_21142,N_21003);
or U21439 (N_21439,N_21197,N_21147);
nor U21440 (N_21440,N_21157,N_21176);
xnor U21441 (N_21441,N_21255,N_21084);
and U21442 (N_21442,N_21024,N_21191);
nor U21443 (N_21443,N_21245,N_21200);
or U21444 (N_21444,N_21086,N_21111);
xor U21445 (N_21445,N_21238,N_21042);
nor U21446 (N_21446,N_21145,N_21287);
nand U21447 (N_21447,N_21285,N_21055);
nor U21448 (N_21448,N_21265,N_21087);
or U21449 (N_21449,N_21152,N_21133);
xnor U21450 (N_21450,N_21256,N_21051);
or U21451 (N_21451,N_21185,N_21024);
nor U21452 (N_21452,N_21233,N_21058);
xor U21453 (N_21453,N_21294,N_21225);
and U21454 (N_21454,N_21115,N_21131);
nor U21455 (N_21455,N_21146,N_21189);
xnor U21456 (N_21456,N_21063,N_21288);
or U21457 (N_21457,N_21147,N_21207);
or U21458 (N_21458,N_21268,N_21263);
and U21459 (N_21459,N_21195,N_21038);
xor U21460 (N_21460,N_21181,N_21056);
nand U21461 (N_21461,N_21005,N_21291);
and U21462 (N_21462,N_21263,N_21028);
xnor U21463 (N_21463,N_21220,N_21236);
nand U21464 (N_21464,N_21233,N_21014);
or U21465 (N_21465,N_21190,N_21179);
nand U21466 (N_21466,N_21169,N_21023);
or U21467 (N_21467,N_21274,N_21270);
xnor U21468 (N_21468,N_21229,N_21281);
xnor U21469 (N_21469,N_21245,N_21028);
and U21470 (N_21470,N_21123,N_21078);
xnor U21471 (N_21471,N_21269,N_21292);
and U21472 (N_21472,N_21127,N_21291);
and U21473 (N_21473,N_21229,N_21138);
nor U21474 (N_21474,N_21287,N_21001);
or U21475 (N_21475,N_21160,N_21081);
nand U21476 (N_21476,N_21063,N_21205);
or U21477 (N_21477,N_21103,N_21181);
nor U21478 (N_21478,N_21102,N_21029);
or U21479 (N_21479,N_21240,N_21219);
xnor U21480 (N_21480,N_21122,N_21091);
and U21481 (N_21481,N_21291,N_21165);
and U21482 (N_21482,N_21059,N_21251);
or U21483 (N_21483,N_21051,N_21036);
or U21484 (N_21484,N_21115,N_21247);
nor U21485 (N_21485,N_21197,N_21194);
nor U21486 (N_21486,N_21126,N_21263);
xor U21487 (N_21487,N_21115,N_21172);
xnor U21488 (N_21488,N_21175,N_21287);
and U21489 (N_21489,N_21227,N_21000);
xnor U21490 (N_21490,N_21037,N_21252);
nand U21491 (N_21491,N_21043,N_21199);
nand U21492 (N_21492,N_21293,N_21011);
nand U21493 (N_21493,N_21062,N_21029);
and U21494 (N_21494,N_21203,N_21244);
nor U21495 (N_21495,N_21138,N_21292);
nand U21496 (N_21496,N_21233,N_21188);
nor U21497 (N_21497,N_21212,N_21012);
nand U21498 (N_21498,N_21039,N_21054);
nand U21499 (N_21499,N_21013,N_21229);
nor U21500 (N_21500,N_21247,N_21116);
and U21501 (N_21501,N_21193,N_21204);
nor U21502 (N_21502,N_21161,N_21016);
xor U21503 (N_21503,N_21085,N_21109);
nand U21504 (N_21504,N_21138,N_21031);
nor U21505 (N_21505,N_21250,N_21038);
and U21506 (N_21506,N_21042,N_21224);
nand U21507 (N_21507,N_21053,N_21046);
and U21508 (N_21508,N_21291,N_21223);
xor U21509 (N_21509,N_21243,N_21227);
xnor U21510 (N_21510,N_21228,N_21116);
or U21511 (N_21511,N_21274,N_21107);
nand U21512 (N_21512,N_21037,N_21189);
nor U21513 (N_21513,N_21231,N_21220);
or U21514 (N_21514,N_21290,N_21079);
and U21515 (N_21515,N_21286,N_21245);
or U21516 (N_21516,N_21225,N_21045);
or U21517 (N_21517,N_21232,N_21014);
nand U21518 (N_21518,N_21036,N_21063);
nor U21519 (N_21519,N_21038,N_21118);
nand U21520 (N_21520,N_21119,N_21282);
and U21521 (N_21521,N_21274,N_21064);
nor U21522 (N_21522,N_21053,N_21276);
or U21523 (N_21523,N_21149,N_21295);
nor U21524 (N_21524,N_21275,N_21055);
nor U21525 (N_21525,N_21005,N_21141);
nor U21526 (N_21526,N_21085,N_21179);
nor U21527 (N_21527,N_21101,N_21174);
nor U21528 (N_21528,N_21269,N_21086);
and U21529 (N_21529,N_21296,N_21179);
nand U21530 (N_21530,N_21284,N_21157);
and U21531 (N_21531,N_21115,N_21185);
xnor U21532 (N_21532,N_21235,N_21205);
xnor U21533 (N_21533,N_21172,N_21148);
nand U21534 (N_21534,N_21211,N_21049);
nand U21535 (N_21535,N_21183,N_21184);
and U21536 (N_21536,N_21285,N_21132);
and U21537 (N_21537,N_21081,N_21227);
nor U21538 (N_21538,N_21187,N_21121);
xor U21539 (N_21539,N_21228,N_21241);
nor U21540 (N_21540,N_21077,N_21123);
nand U21541 (N_21541,N_21297,N_21082);
nand U21542 (N_21542,N_21215,N_21033);
xnor U21543 (N_21543,N_21067,N_21174);
or U21544 (N_21544,N_21135,N_21267);
or U21545 (N_21545,N_21109,N_21120);
or U21546 (N_21546,N_21271,N_21210);
nand U21547 (N_21547,N_21085,N_21155);
and U21548 (N_21548,N_21040,N_21215);
or U21549 (N_21549,N_21040,N_21192);
nor U21550 (N_21550,N_21276,N_21164);
and U21551 (N_21551,N_21097,N_21045);
nor U21552 (N_21552,N_21244,N_21157);
and U21553 (N_21553,N_21225,N_21273);
and U21554 (N_21554,N_21158,N_21072);
nand U21555 (N_21555,N_21206,N_21068);
xnor U21556 (N_21556,N_21140,N_21200);
and U21557 (N_21557,N_21276,N_21292);
and U21558 (N_21558,N_21011,N_21058);
xor U21559 (N_21559,N_21219,N_21227);
or U21560 (N_21560,N_21250,N_21295);
nand U21561 (N_21561,N_21057,N_21250);
xnor U21562 (N_21562,N_21027,N_21293);
or U21563 (N_21563,N_21250,N_21163);
xnor U21564 (N_21564,N_21093,N_21267);
or U21565 (N_21565,N_21145,N_21117);
and U21566 (N_21566,N_21014,N_21261);
and U21567 (N_21567,N_21284,N_21007);
nor U21568 (N_21568,N_21246,N_21093);
nor U21569 (N_21569,N_21138,N_21052);
nor U21570 (N_21570,N_21169,N_21162);
nand U21571 (N_21571,N_21147,N_21086);
and U21572 (N_21572,N_21138,N_21063);
nor U21573 (N_21573,N_21297,N_21095);
and U21574 (N_21574,N_21275,N_21194);
xor U21575 (N_21575,N_21057,N_21213);
xnor U21576 (N_21576,N_21219,N_21074);
nor U21577 (N_21577,N_21031,N_21199);
nand U21578 (N_21578,N_21087,N_21201);
or U21579 (N_21579,N_21297,N_21096);
xor U21580 (N_21580,N_21253,N_21054);
nor U21581 (N_21581,N_21224,N_21187);
nand U21582 (N_21582,N_21115,N_21081);
and U21583 (N_21583,N_21247,N_21076);
nor U21584 (N_21584,N_21067,N_21124);
nand U21585 (N_21585,N_21190,N_21105);
nor U21586 (N_21586,N_21102,N_21040);
and U21587 (N_21587,N_21212,N_21240);
xor U21588 (N_21588,N_21184,N_21203);
nor U21589 (N_21589,N_21013,N_21252);
xnor U21590 (N_21590,N_21063,N_21256);
and U21591 (N_21591,N_21190,N_21088);
nor U21592 (N_21592,N_21122,N_21203);
nand U21593 (N_21593,N_21016,N_21076);
xnor U21594 (N_21594,N_21109,N_21219);
and U21595 (N_21595,N_21223,N_21232);
and U21596 (N_21596,N_21277,N_21142);
nand U21597 (N_21597,N_21078,N_21273);
xnor U21598 (N_21598,N_21015,N_21029);
or U21599 (N_21599,N_21202,N_21037);
nor U21600 (N_21600,N_21504,N_21554);
nand U21601 (N_21601,N_21572,N_21520);
nor U21602 (N_21602,N_21505,N_21467);
nand U21603 (N_21603,N_21486,N_21507);
nand U21604 (N_21604,N_21466,N_21359);
and U21605 (N_21605,N_21559,N_21409);
xor U21606 (N_21606,N_21301,N_21581);
and U21607 (N_21607,N_21365,N_21519);
nor U21608 (N_21608,N_21441,N_21338);
nor U21609 (N_21609,N_21378,N_21410);
nand U21610 (N_21610,N_21584,N_21318);
nand U21611 (N_21611,N_21588,N_21339);
nand U21612 (N_21612,N_21470,N_21597);
nand U21613 (N_21613,N_21328,N_21349);
and U21614 (N_21614,N_21502,N_21325);
nand U21615 (N_21615,N_21313,N_21333);
and U21616 (N_21616,N_21516,N_21380);
nand U21617 (N_21617,N_21457,N_21362);
nand U21618 (N_21618,N_21562,N_21364);
and U21619 (N_21619,N_21542,N_21398);
nand U21620 (N_21620,N_21553,N_21568);
nand U21621 (N_21621,N_21421,N_21548);
or U21622 (N_21622,N_21371,N_21435);
xor U21623 (N_21623,N_21425,N_21387);
xnor U21624 (N_21624,N_21352,N_21375);
and U21625 (N_21625,N_21503,N_21514);
and U21626 (N_21626,N_21443,N_21305);
and U21627 (N_21627,N_21575,N_21414);
and U21628 (N_21628,N_21307,N_21451);
and U21629 (N_21629,N_21423,N_21437);
nand U21630 (N_21630,N_21401,N_21513);
nand U21631 (N_21631,N_21476,N_21337);
and U21632 (N_21632,N_21388,N_21518);
xor U21633 (N_21633,N_21506,N_21406);
or U21634 (N_21634,N_21461,N_21422);
or U21635 (N_21635,N_21569,N_21356);
nor U21636 (N_21636,N_21453,N_21563);
or U21637 (N_21637,N_21442,N_21521);
or U21638 (N_21638,N_21404,N_21412);
xor U21639 (N_21639,N_21446,N_21590);
and U21640 (N_21640,N_21574,N_21386);
nor U21641 (N_21641,N_21493,N_21576);
nand U21642 (N_21642,N_21557,N_21529);
nand U21643 (N_21643,N_21447,N_21561);
or U21644 (N_21644,N_21471,N_21587);
and U21645 (N_21645,N_21340,N_21427);
xor U21646 (N_21646,N_21345,N_21434);
nand U21647 (N_21647,N_21302,N_21303);
or U21648 (N_21648,N_21577,N_21495);
nand U21649 (N_21649,N_21540,N_21396);
and U21650 (N_21650,N_21458,N_21330);
nor U21651 (N_21651,N_21573,N_21537);
and U21652 (N_21652,N_21402,N_21585);
nand U21653 (N_21653,N_21580,N_21530);
xor U21654 (N_21654,N_21323,N_21360);
or U21655 (N_21655,N_21450,N_21555);
nand U21656 (N_21656,N_21353,N_21405);
nor U21657 (N_21657,N_21547,N_21456);
or U21658 (N_21658,N_21515,N_21381);
nor U21659 (N_21659,N_21429,N_21361);
and U21660 (N_21660,N_21475,N_21312);
nor U21661 (N_21661,N_21327,N_21355);
or U21662 (N_21662,N_21477,N_21424);
or U21663 (N_21663,N_21489,N_21321);
nor U21664 (N_21664,N_21465,N_21481);
xnor U21665 (N_21665,N_21415,N_21319);
and U21666 (N_21666,N_21314,N_21463);
nand U21667 (N_21667,N_21394,N_21390);
or U21668 (N_21668,N_21374,N_21599);
nor U21669 (N_21669,N_21528,N_21532);
nor U21670 (N_21670,N_21464,N_21335);
xor U21671 (N_21671,N_21315,N_21354);
or U21672 (N_21672,N_21311,N_21370);
or U21673 (N_21673,N_21436,N_21510);
xor U21674 (N_21674,N_21449,N_21376);
nand U21675 (N_21675,N_21395,N_21309);
or U21676 (N_21676,N_21544,N_21543);
nor U21677 (N_21677,N_21462,N_21533);
nor U21678 (N_21678,N_21591,N_21480);
xnor U21679 (N_21679,N_21560,N_21500);
or U21680 (N_21680,N_21347,N_21306);
nor U21681 (N_21681,N_21369,N_21350);
and U21682 (N_21682,N_21433,N_21541);
nor U21683 (N_21683,N_21596,N_21346);
nand U21684 (N_21684,N_21391,N_21534);
or U21685 (N_21685,N_21400,N_21331);
xor U21686 (N_21686,N_21420,N_21320);
nand U21687 (N_21687,N_21417,N_21492);
nor U21688 (N_21688,N_21536,N_21334);
xnor U21689 (N_21689,N_21368,N_21566);
xor U21690 (N_21690,N_21324,N_21509);
xor U21691 (N_21691,N_21418,N_21316);
nor U21692 (N_21692,N_21598,N_21497);
nor U21693 (N_21693,N_21485,N_21539);
nor U21694 (N_21694,N_21508,N_21479);
or U21695 (N_21695,N_21348,N_21525);
xnor U21696 (N_21696,N_21571,N_21411);
xor U21697 (N_21697,N_21416,N_21379);
and U21698 (N_21698,N_21432,N_21531);
nor U21699 (N_21699,N_21392,N_21473);
nor U21700 (N_21700,N_21439,N_21428);
and U21701 (N_21701,N_21430,N_21490);
nand U21702 (N_21702,N_21455,N_21438);
xor U21703 (N_21703,N_21593,N_21579);
and U21704 (N_21704,N_21499,N_21389);
or U21705 (N_21705,N_21377,N_21511);
nand U21706 (N_21706,N_21484,N_21440);
nor U21707 (N_21707,N_21556,N_21565);
or U21708 (N_21708,N_21583,N_21413);
nand U21709 (N_21709,N_21383,N_21501);
and U21710 (N_21710,N_21472,N_21524);
nand U21711 (N_21711,N_21384,N_21397);
or U21712 (N_21712,N_21523,N_21512);
xnor U21713 (N_21713,N_21491,N_21342);
and U21714 (N_21714,N_21550,N_21460);
nand U21715 (N_21715,N_21341,N_21308);
xor U21716 (N_21716,N_21452,N_21578);
or U21717 (N_21717,N_21488,N_21545);
or U21718 (N_21718,N_21399,N_21496);
nor U21719 (N_21719,N_21592,N_21552);
xnor U21720 (N_21720,N_21549,N_21431);
or U21721 (N_21721,N_21445,N_21487);
nor U21722 (N_21722,N_21317,N_21336);
nand U21723 (N_21723,N_21459,N_21448);
or U21724 (N_21724,N_21344,N_21326);
nand U21725 (N_21725,N_21382,N_21332);
and U21726 (N_21726,N_21367,N_21403);
nand U21727 (N_21727,N_21351,N_21454);
or U21728 (N_21728,N_21498,N_21522);
nand U21729 (N_21729,N_21494,N_21564);
nor U21730 (N_21730,N_21551,N_21310);
nand U21731 (N_21731,N_21474,N_21546);
and U21732 (N_21732,N_21408,N_21586);
xor U21733 (N_21733,N_21426,N_21483);
or U21734 (N_21734,N_21594,N_21468);
xnor U21735 (N_21735,N_21357,N_21478);
or U21736 (N_21736,N_21300,N_21373);
and U21737 (N_21737,N_21358,N_21589);
or U21738 (N_21738,N_21393,N_21567);
nand U21739 (N_21739,N_21482,N_21535);
or U21740 (N_21740,N_21372,N_21385);
nand U21741 (N_21741,N_21407,N_21304);
nor U21742 (N_21742,N_21363,N_21595);
xor U21743 (N_21743,N_21469,N_21558);
xnor U21744 (N_21744,N_21366,N_21343);
xnor U21745 (N_21745,N_21444,N_21517);
nor U21746 (N_21746,N_21570,N_21527);
or U21747 (N_21747,N_21538,N_21329);
nand U21748 (N_21748,N_21526,N_21419);
nand U21749 (N_21749,N_21322,N_21582);
and U21750 (N_21750,N_21437,N_21497);
xor U21751 (N_21751,N_21544,N_21561);
nand U21752 (N_21752,N_21460,N_21462);
nand U21753 (N_21753,N_21412,N_21395);
nor U21754 (N_21754,N_21391,N_21462);
or U21755 (N_21755,N_21572,N_21433);
xor U21756 (N_21756,N_21555,N_21309);
nor U21757 (N_21757,N_21564,N_21589);
and U21758 (N_21758,N_21467,N_21431);
nand U21759 (N_21759,N_21392,N_21311);
nand U21760 (N_21760,N_21574,N_21360);
and U21761 (N_21761,N_21428,N_21599);
nand U21762 (N_21762,N_21545,N_21379);
or U21763 (N_21763,N_21453,N_21463);
and U21764 (N_21764,N_21459,N_21596);
xor U21765 (N_21765,N_21461,N_21495);
nand U21766 (N_21766,N_21422,N_21448);
nand U21767 (N_21767,N_21453,N_21415);
xnor U21768 (N_21768,N_21351,N_21325);
and U21769 (N_21769,N_21584,N_21524);
nand U21770 (N_21770,N_21574,N_21475);
and U21771 (N_21771,N_21361,N_21427);
or U21772 (N_21772,N_21359,N_21492);
nand U21773 (N_21773,N_21374,N_21451);
and U21774 (N_21774,N_21369,N_21360);
nor U21775 (N_21775,N_21365,N_21554);
nor U21776 (N_21776,N_21327,N_21344);
nor U21777 (N_21777,N_21530,N_21537);
xor U21778 (N_21778,N_21328,N_21543);
nand U21779 (N_21779,N_21330,N_21512);
and U21780 (N_21780,N_21389,N_21581);
and U21781 (N_21781,N_21587,N_21454);
nor U21782 (N_21782,N_21347,N_21389);
xor U21783 (N_21783,N_21563,N_21596);
or U21784 (N_21784,N_21365,N_21380);
nor U21785 (N_21785,N_21426,N_21450);
and U21786 (N_21786,N_21333,N_21525);
nand U21787 (N_21787,N_21476,N_21329);
xnor U21788 (N_21788,N_21588,N_21400);
nor U21789 (N_21789,N_21556,N_21420);
or U21790 (N_21790,N_21430,N_21308);
nand U21791 (N_21791,N_21508,N_21417);
nand U21792 (N_21792,N_21474,N_21595);
xor U21793 (N_21793,N_21583,N_21563);
and U21794 (N_21794,N_21301,N_21333);
nand U21795 (N_21795,N_21548,N_21332);
or U21796 (N_21796,N_21325,N_21345);
and U21797 (N_21797,N_21323,N_21337);
and U21798 (N_21798,N_21326,N_21425);
nand U21799 (N_21799,N_21412,N_21365);
xnor U21800 (N_21800,N_21423,N_21517);
nor U21801 (N_21801,N_21567,N_21525);
nand U21802 (N_21802,N_21375,N_21372);
or U21803 (N_21803,N_21515,N_21443);
or U21804 (N_21804,N_21413,N_21330);
nor U21805 (N_21805,N_21484,N_21441);
xor U21806 (N_21806,N_21590,N_21403);
xnor U21807 (N_21807,N_21388,N_21540);
or U21808 (N_21808,N_21456,N_21512);
xor U21809 (N_21809,N_21336,N_21459);
nand U21810 (N_21810,N_21533,N_21457);
and U21811 (N_21811,N_21408,N_21330);
nand U21812 (N_21812,N_21338,N_21332);
or U21813 (N_21813,N_21326,N_21474);
or U21814 (N_21814,N_21464,N_21578);
and U21815 (N_21815,N_21378,N_21371);
and U21816 (N_21816,N_21540,N_21534);
nand U21817 (N_21817,N_21512,N_21348);
xnor U21818 (N_21818,N_21443,N_21354);
or U21819 (N_21819,N_21451,N_21309);
or U21820 (N_21820,N_21312,N_21387);
xnor U21821 (N_21821,N_21477,N_21520);
nor U21822 (N_21822,N_21469,N_21384);
nor U21823 (N_21823,N_21377,N_21394);
nor U21824 (N_21824,N_21435,N_21427);
and U21825 (N_21825,N_21555,N_21391);
nand U21826 (N_21826,N_21448,N_21440);
xnor U21827 (N_21827,N_21477,N_21454);
xor U21828 (N_21828,N_21500,N_21383);
and U21829 (N_21829,N_21557,N_21379);
xnor U21830 (N_21830,N_21462,N_21321);
xnor U21831 (N_21831,N_21322,N_21323);
or U21832 (N_21832,N_21566,N_21413);
xnor U21833 (N_21833,N_21349,N_21582);
and U21834 (N_21834,N_21587,N_21442);
or U21835 (N_21835,N_21516,N_21405);
or U21836 (N_21836,N_21412,N_21564);
or U21837 (N_21837,N_21301,N_21416);
and U21838 (N_21838,N_21311,N_21593);
nand U21839 (N_21839,N_21492,N_21358);
or U21840 (N_21840,N_21377,N_21527);
and U21841 (N_21841,N_21489,N_21409);
xnor U21842 (N_21842,N_21520,N_21563);
or U21843 (N_21843,N_21514,N_21438);
nor U21844 (N_21844,N_21356,N_21312);
xnor U21845 (N_21845,N_21541,N_21423);
xor U21846 (N_21846,N_21391,N_21409);
xnor U21847 (N_21847,N_21411,N_21377);
nand U21848 (N_21848,N_21337,N_21472);
nor U21849 (N_21849,N_21343,N_21373);
xor U21850 (N_21850,N_21312,N_21319);
or U21851 (N_21851,N_21475,N_21400);
xor U21852 (N_21852,N_21381,N_21384);
and U21853 (N_21853,N_21355,N_21393);
or U21854 (N_21854,N_21536,N_21386);
nand U21855 (N_21855,N_21415,N_21526);
or U21856 (N_21856,N_21344,N_21385);
xnor U21857 (N_21857,N_21311,N_21506);
and U21858 (N_21858,N_21465,N_21526);
or U21859 (N_21859,N_21432,N_21308);
or U21860 (N_21860,N_21458,N_21586);
or U21861 (N_21861,N_21563,N_21523);
nor U21862 (N_21862,N_21336,N_21520);
nand U21863 (N_21863,N_21336,N_21458);
nor U21864 (N_21864,N_21421,N_21498);
nand U21865 (N_21865,N_21342,N_21324);
xnor U21866 (N_21866,N_21488,N_21315);
nor U21867 (N_21867,N_21333,N_21328);
and U21868 (N_21868,N_21334,N_21330);
and U21869 (N_21869,N_21480,N_21543);
xor U21870 (N_21870,N_21572,N_21589);
xnor U21871 (N_21871,N_21370,N_21522);
and U21872 (N_21872,N_21586,N_21385);
and U21873 (N_21873,N_21572,N_21498);
xor U21874 (N_21874,N_21309,N_21459);
nor U21875 (N_21875,N_21364,N_21582);
xor U21876 (N_21876,N_21422,N_21443);
nor U21877 (N_21877,N_21428,N_21319);
or U21878 (N_21878,N_21524,N_21593);
or U21879 (N_21879,N_21419,N_21565);
xnor U21880 (N_21880,N_21426,N_21507);
or U21881 (N_21881,N_21385,N_21306);
and U21882 (N_21882,N_21451,N_21329);
nand U21883 (N_21883,N_21482,N_21307);
and U21884 (N_21884,N_21343,N_21560);
xor U21885 (N_21885,N_21457,N_21524);
or U21886 (N_21886,N_21420,N_21346);
xnor U21887 (N_21887,N_21441,N_21485);
xor U21888 (N_21888,N_21326,N_21312);
or U21889 (N_21889,N_21543,N_21326);
xnor U21890 (N_21890,N_21376,N_21432);
and U21891 (N_21891,N_21556,N_21518);
xor U21892 (N_21892,N_21530,N_21467);
nor U21893 (N_21893,N_21451,N_21461);
xor U21894 (N_21894,N_21541,N_21596);
or U21895 (N_21895,N_21373,N_21442);
nand U21896 (N_21896,N_21464,N_21359);
and U21897 (N_21897,N_21547,N_21509);
and U21898 (N_21898,N_21404,N_21345);
or U21899 (N_21899,N_21488,N_21528);
or U21900 (N_21900,N_21818,N_21870);
xor U21901 (N_21901,N_21653,N_21754);
and U21902 (N_21902,N_21723,N_21770);
and U21903 (N_21903,N_21684,N_21657);
nand U21904 (N_21904,N_21862,N_21830);
nor U21905 (N_21905,N_21753,N_21732);
nand U21906 (N_21906,N_21806,N_21821);
nor U21907 (N_21907,N_21876,N_21882);
nor U21908 (N_21908,N_21796,N_21704);
nor U21909 (N_21909,N_21625,N_21603);
nand U21910 (N_21910,N_21757,N_21825);
nor U21911 (N_21911,N_21716,N_21655);
nand U21912 (N_21912,N_21823,N_21812);
nor U21913 (N_21913,N_21696,N_21744);
and U21914 (N_21914,N_21609,N_21700);
xnor U21915 (N_21915,N_21842,N_21802);
and U21916 (N_21916,N_21665,N_21675);
or U21917 (N_21917,N_21865,N_21797);
and U21918 (N_21918,N_21729,N_21750);
or U21919 (N_21919,N_21746,N_21861);
xor U21920 (N_21920,N_21889,N_21624);
or U21921 (N_21921,N_21883,N_21899);
xnor U21922 (N_21922,N_21714,N_21843);
and U21923 (N_21923,N_21793,N_21745);
nand U21924 (N_21924,N_21869,N_21715);
nor U21925 (N_21925,N_21637,N_21803);
nor U21926 (N_21926,N_21819,N_21814);
nor U21927 (N_21927,N_21709,N_21604);
nor U21928 (N_21928,N_21671,N_21766);
nand U21929 (N_21929,N_21602,N_21719);
or U21930 (N_21930,N_21670,N_21683);
nand U21931 (N_21931,N_21769,N_21779);
nor U21932 (N_21932,N_21826,N_21787);
or U21933 (N_21933,N_21789,N_21689);
nor U21934 (N_21934,N_21620,N_21771);
xnor U21935 (N_21935,N_21785,N_21833);
xor U21936 (N_21936,N_21688,N_21897);
xnor U21937 (N_21937,N_21698,N_21764);
xor U21938 (N_21938,N_21879,N_21840);
nor U21939 (N_21939,N_21672,N_21634);
nand U21940 (N_21940,N_21706,N_21780);
xnor U21941 (N_21941,N_21648,N_21893);
and U21942 (N_21942,N_21642,N_21791);
nor U21943 (N_21943,N_21852,N_21717);
nor U21944 (N_21944,N_21873,N_21762);
or U21945 (N_21945,N_21794,N_21828);
or U21946 (N_21946,N_21857,N_21761);
nand U21947 (N_21947,N_21649,N_21608);
or U21948 (N_21948,N_21886,N_21892);
nand U21949 (N_21949,N_21699,N_21816);
or U21950 (N_21950,N_21749,N_21752);
nand U21951 (N_21951,N_21827,N_21659);
nand U21952 (N_21952,N_21740,N_21663);
nor U21953 (N_21953,N_21838,N_21601);
and U21954 (N_21954,N_21645,N_21864);
and U21955 (N_21955,N_21713,N_21612);
xor U21956 (N_21956,N_21868,N_21845);
or U21957 (N_21957,N_21773,N_21777);
or U21958 (N_21958,N_21735,N_21631);
and U21959 (N_21959,N_21756,N_21619);
and U21960 (N_21960,N_21682,N_21686);
or U21961 (N_21961,N_21822,N_21772);
nor U21962 (N_21962,N_21703,N_21694);
nand U21963 (N_21963,N_21765,N_21859);
xnor U21964 (N_21964,N_21707,N_21844);
or U21965 (N_21965,N_21627,N_21669);
or U21966 (N_21966,N_21853,N_21606);
or U21967 (N_21967,N_21884,N_21691);
and U21968 (N_21968,N_21808,N_21721);
nand U21969 (N_21969,N_21712,N_21877);
xnor U21970 (N_21970,N_21759,N_21805);
or U21971 (N_21971,N_21635,N_21760);
xnor U21972 (N_21972,N_21734,N_21871);
xnor U21973 (N_21973,N_21741,N_21662);
nor U21974 (N_21974,N_21885,N_21829);
or U21975 (N_21975,N_21846,N_21632);
xnor U21976 (N_21976,N_21739,N_21701);
nand U21977 (N_21977,N_21654,N_21743);
nand U21978 (N_21978,N_21737,N_21863);
nor U21979 (N_21979,N_21668,N_21834);
xnor U21980 (N_21980,N_21693,N_21809);
and U21981 (N_21981,N_21730,N_21888);
xor U21982 (N_21982,N_21621,N_21849);
nand U21983 (N_21983,N_21810,N_21678);
or U21984 (N_21984,N_21775,N_21705);
or U21985 (N_21985,N_21898,N_21801);
or U21986 (N_21986,N_21799,N_21835);
xor U21987 (N_21987,N_21839,N_21613);
nand U21988 (N_21988,N_21788,N_21792);
and U21989 (N_21989,N_21643,N_21605);
xnor U21990 (N_21990,N_21628,N_21751);
xor U21991 (N_21991,N_21781,N_21674);
and U21992 (N_21992,N_21639,N_21646);
or U21993 (N_21993,N_21666,N_21687);
and U21994 (N_21994,N_21872,N_21807);
or U21995 (N_21995,N_21854,N_21633);
xnor U21996 (N_21996,N_21677,N_21733);
or U21997 (N_21997,N_21811,N_21774);
nand U21998 (N_21998,N_21820,N_21640);
or U21999 (N_21999,N_21630,N_21860);
or U22000 (N_22000,N_21790,N_21600);
and U22001 (N_22001,N_21736,N_21626);
nor U22002 (N_22002,N_21881,N_21664);
xor U22003 (N_22003,N_21875,N_21615);
or U22004 (N_22004,N_21644,N_21660);
nor U22005 (N_22005,N_21728,N_21692);
xnor U22006 (N_22006,N_21724,N_21798);
xnor U22007 (N_22007,N_21702,N_21891);
or U22008 (N_22008,N_21837,N_21786);
nor U22009 (N_22009,N_21848,N_21763);
and U22010 (N_22010,N_21855,N_21817);
and U22011 (N_22011,N_21618,N_21856);
nand U22012 (N_22012,N_21858,N_21718);
or U22013 (N_22013,N_21804,N_21758);
or U22014 (N_22014,N_21836,N_21795);
nand U22015 (N_22015,N_21607,N_21641);
xor U22016 (N_22016,N_21831,N_21647);
nor U22017 (N_22017,N_21614,N_21711);
xnor U22018 (N_22018,N_21710,N_21673);
and U22019 (N_22019,N_21866,N_21890);
or U22020 (N_22020,N_21824,N_21720);
or U22021 (N_22021,N_21747,N_21767);
nand U22022 (N_22022,N_21742,N_21726);
nor U22023 (N_22023,N_21629,N_21874);
nand U22024 (N_22024,N_21782,N_21776);
and U22025 (N_22025,N_21695,N_21887);
or U22026 (N_22026,N_21708,N_21611);
and U22027 (N_22027,N_21755,N_21690);
xnor U22028 (N_22028,N_21667,N_21880);
nand U22029 (N_22029,N_21878,N_21622);
xnor U22030 (N_22030,N_21894,N_21841);
xnor U22031 (N_22031,N_21800,N_21676);
or U22032 (N_22032,N_21813,N_21661);
nor U22033 (N_22033,N_21851,N_21697);
nor U22034 (N_22034,N_21748,N_21778);
nand U22035 (N_22035,N_21725,N_21658);
xnor U22036 (N_22036,N_21623,N_21896);
and U22037 (N_22037,N_21727,N_21616);
xnor U22038 (N_22038,N_21681,N_21679);
nand U22039 (N_22039,N_21650,N_21738);
nand U22040 (N_22040,N_21784,N_21636);
and U22041 (N_22041,N_21867,N_21815);
nand U22042 (N_22042,N_21847,N_21680);
xnor U22043 (N_22043,N_21895,N_21651);
and U22044 (N_22044,N_21685,N_21652);
nand U22045 (N_22045,N_21617,N_21832);
nand U22046 (N_22046,N_21731,N_21656);
nor U22047 (N_22047,N_21722,N_21610);
and U22048 (N_22048,N_21850,N_21783);
xor U22049 (N_22049,N_21768,N_21638);
xor U22050 (N_22050,N_21842,N_21662);
and U22051 (N_22051,N_21816,N_21639);
and U22052 (N_22052,N_21786,N_21724);
nor U22053 (N_22053,N_21808,N_21602);
and U22054 (N_22054,N_21707,N_21724);
nand U22055 (N_22055,N_21807,N_21890);
xnor U22056 (N_22056,N_21627,N_21821);
xnor U22057 (N_22057,N_21821,N_21803);
or U22058 (N_22058,N_21703,N_21776);
and U22059 (N_22059,N_21845,N_21622);
nand U22060 (N_22060,N_21680,N_21814);
nor U22061 (N_22061,N_21882,N_21640);
nand U22062 (N_22062,N_21826,N_21775);
or U22063 (N_22063,N_21801,N_21730);
nand U22064 (N_22064,N_21619,N_21882);
xor U22065 (N_22065,N_21651,N_21669);
and U22066 (N_22066,N_21614,N_21805);
or U22067 (N_22067,N_21625,N_21767);
or U22068 (N_22068,N_21887,N_21704);
xnor U22069 (N_22069,N_21607,N_21623);
and U22070 (N_22070,N_21639,N_21661);
xor U22071 (N_22071,N_21793,N_21732);
nand U22072 (N_22072,N_21882,N_21714);
nor U22073 (N_22073,N_21840,N_21779);
nor U22074 (N_22074,N_21668,N_21630);
xnor U22075 (N_22075,N_21673,N_21641);
nor U22076 (N_22076,N_21637,N_21687);
nand U22077 (N_22077,N_21881,N_21702);
xnor U22078 (N_22078,N_21652,N_21786);
or U22079 (N_22079,N_21748,N_21828);
nand U22080 (N_22080,N_21749,N_21661);
xor U22081 (N_22081,N_21813,N_21663);
nand U22082 (N_22082,N_21750,N_21609);
xor U22083 (N_22083,N_21694,N_21840);
xnor U22084 (N_22084,N_21768,N_21751);
xor U22085 (N_22085,N_21753,N_21641);
nand U22086 (N_22086,N_21686,N_21617);
nor U22087 (N_22087,N_21681,N_21706);
nor U22088 (N_22088,N_21616,N_21753);
xor U22089 (N_22089,N_21680,N_21649);
nor U22090 (N_22090,N_21721,N_21727);
nor U22091 (N_22091,N_21827,N_21761);
and U22092 (N_22092,N_21864,N_21656);
or U22093 (N_22093,N_21628,N_21813);
and U22094 (N_22094,N_21621,N_21609);
xnor U22095 (N_22095,N_21641,N_21612);
nand U22096 (N_22096,N_21773,N_21630);
nor U22097 (N_22097,N_21717,N_21778);
xor U22098 (N_22098,N_21617,N_21828);
nor U22099 (N_22099,N_21754,N_21644);
and U22100 (N_22100,N_21880,N_21827);
xnor U22101 (N_22101,N_21758,N_21653);
and U22102 (N_22102,N_21696,N_21606);
and U22103 (N_22103,N_21869,N_21662);
nand U22104 (N_22104,N_21782,N_21730);
nor U22105 (N_22105,N_21763,N_21775);
xor U22106 (N_22106,N_21632,N_21662);
or U22107 (N_22107,N_21623,N_21751);
or U22108 (N_22108,N_21674,N_21633);
nand U22109 (N_22109,N_21748,N_21855);
xnor U22110 (N_22110,N_21834,N_21755);
xnor U22111 (N_22111,N_21732,N_21858);
or U22112 (N_22112,N_21831,N_21627);
nor U22113 (N_22113,N_21642,N_21734);
xnor U22114 (N_22114,N_21688,N_21874);
and U22115 (N_22115,N_21634,N_21821);
or U22116 (N_22116,N_21862,N_21807);
xor U22117 (N_22117,N_21743,N_21704);
nor U22118 (N_22118,N_21763,N_21750);
or U22119 (N_22119,N_21860,N_21815);
nor U22120 (N_22120,N_21623,N_21815);
or U22121 (N_22121,N_21831,N_21836);
or U22122 (N_22122,N_21624,N_21766);
nand U22123 (N_22123,N_21810,N_21768);
xnor U22124 (N_22124,N_21605,N_21809);
xor U22125 (N_22125,N_21612,N_21614);
nor U22126 (N_22126,N_21884,N_21899);
xnor U22127 (N_22127,N_21824,N_21666);
nand U22128 (N_22128,N_21846,N_21793);
or U22129 (N_22129,N_21686,N_21833);
and U22130 (N_22130,N_21764,N_21760);
or U22131 (N_22131,N_21706,N_21752);
or U22132 (N_22132,N_21845,N_21696);
and U22133 (N_22133,N_21886,N_21648);
nand U22134 (N_22134,N_21852,N_21893);
nor U22135 (N_22135,N_21621,N_21748);
nor U22136 (N_22136,N_21690,N_21814);
and U22137 (N_22137,N_21802,N_21856);
nor U22138 (N_22138,N_21667,N_21640);
or U22139 (N_22139,N_21739,N_21698);
xor U22140 (N_22140,N_21745,N_21642);
nand U22141 (N_22141,N_21866,N_21614);
and U22142 (N_22142,N_21650,N_21614);
and U22143 (N_22143,N_21875,N_21746);
xor U22144 (N_22144,N_21673,N_21712);
xor U22145 (N_22145,N_21884,N_21821);
nor U22146 (N_22146,N_21810,N_21755);
or U22147 (N_22147,N_21794,N_21896);
xnor U22148 (N_22148,N_21793,N_21850);
xor U22149 (N_22149,N_21843,N_21647);
or U22150 (N_22150,N_21844,N_21609);
nor U22151 (N_22151,N_21832,N_21669);
or U22152 (N_22152,N_21854,N_21611);
xor U22153 (N_22153,N_21653,N_21813);
nor U22154 (N_22154,N_21653,N_21628);
or U22155 (N_22155,N_21776,N_21793);
and U22156 (N_22156,N_21757,N_21671);
nor U22157 (N_22157,N_21649,N_21875);
nor U22158 (N_22158,N_21663,N_21734);
xnor U22159 (N_22159,N_21833,N_21637);
xnor U22160 (N_22160,N_21781,N_21613);
xor U22161 (N_22161,N_21827,N_21707);
or U22162 (N_22162,N_21764,N_21697);
nand U22163 (N_22163,N_21770,N_21737);
nor U22164 (N_22164,N_21639,N_21720);
nor U22165 (N_22165,N_21812,N_21608);
nand U22166 (N_22166,N_21735,N_21869);
nand U22167 (N_22167,N_21647,N_21608);
and U22168 (N_22168,N_21834,N_21745);
or U22169 (N_22169,N_21790,N_21818);
nor U22170 (N_22170,N_21783,N_21732);
xnor U22171 (N_22171,N_21657,N_21835);
nand U22172 (N_22172,N_21756,N_21805);
nor U22173 (N_22173,N_21641,N_21601);
and U22174 (N_22174,N_21793,N_21861);
nor U22175 (N_22175,N_21600,N_21705);
nor U22176 (N_22176,N_21630,N_21678);
and U22177 (N_22177,N_21880,N_21619);
nand U22178 (N_22178,N_21783,N_21840);
nand U22179 (N_22179,N_21789,N_21608);
nor U22180 (N_22180,N_21829,N_21775);
nand U22181 (N_22181,N_21639,N_21883);
nor U22182 (N_22182,N_21664,N_21800);
nor U22183 (N_22183,N_21771,N_21805);
or U22184 (N_22184,N_21617,N_21830);
and U22185 (N_22185,N_21689,N_21696);
or U22186 (N_22186,N_21700,N_21860);
xnor U22187 (N_22187,N_21864,N_21665);
nand U22188 (N_22188,N_21788,N_21685);
nor U22189 (N_22189,N_21833,N_21850);
and U22190 (N_22190,N_21612,N_21693);
or U22191 (N_22191,N_21650,N_21791);
or U22192 (N_22192,N_21662,N_21862);
nand U22193 (N_22193,N_21827,N_21772);
and U22194 (N_22194,N_21751,N_21846);
nor U22195 (N_22195,N_21639,N_21834);
nor U22196 (N_22196,N_21880,N_21836);
and U22197 (N_22197,N_21772,N_21682);
and U22198 (N_22198,N_21605,N_21637);
and U22199 (N_22199,N_21750,N_21867);
nand U22200 (N_22200,N_22157,N_22015);
nand U22201 (N_22201,N_22140,N_22170);
xor U22202 (N_22202,N_22021,N_22127);
and U22203 (N_22203,N_21913,N_21929);
nor U22204 (N_22204,N_22044,N_21915);
and U22205 (N_22205,N_22019,N_21969);
xnor U22206 (N_22206,N_21903,N_21946);
nand U22207 (N_22207,N_22112,N_22158);
nor U22208 (N_22208,N_22133,N_22060);
nand U22209 (N_22209,N_21914,N_21908);
and U22210 (N_22210,N_22057,N_22121);
nand U22211 (N_22211,N_21965,N_22191);
and U22212 (N_22212,N_22146,N_22061);
or U22213 (N_22213,N_22055,N_21952);
or U22214 (N_22214,N_21987,N_22190);
or U22215 (N_22215,N_22045,N_22197);
nand U22216 (N_22216,N_22184,N_22004);
nand U22217 (N_22217,N_22056,N_22027);
and U22218 (N_22218,N_21958,N_22094);
nand U22219 (N_22219,N_22033,N_22043);
or U22220 (N_22220,N_22165,N_22042);
or U22221 (N_22221,N_22011,N_22059);
or U22222 (N_22222,N_22109,N_22012);
and U22223 (N_22223,N_21941,N_22030);
and U22224 (N_22224,N_22174,N_22028);
or U22225 (N_22225,N_22001,N_22072);
xnor U22226 (N_22226,N_21973,N_21954);
or U22227 (N_22227,N_22176,N_22107);
nor U22228 (N_22228,N_21905,N_21989);
nor U22229 (N_22229,N_22037,N_22089);
or U22230 (N_22230,N_22171,N_21967);
or U22231 (N_22231,N_22151,N_21962);
xor U22232 (N_22232,N_21988,N_22169);
or U22233 (N_22233,N_22187,N_22083);
nand U22234 (N_22234,N_22132,N_22068);
or U22235 (N_22235,N_21953,N_22147);
nor U22236 (N_22236,N_21975,N_22149);
or U22237 (N_22237,N_21966,N_22185);
and U22238 (N_22238,N_22102,N_21907);
nor U22239 (N_22239,N_22155,N_21947);
or U22240 (N_22240,N_22082,N_22078);
nor U22241 (N_22241,N_22017,N_22116);
and U22242 (N_22242,N_22054,N_22179);
xor U22243 (N_22243,N_22138,N_21925);
and U22244 (N_22244,N_21990,N_21995);
xnor U22245 (N_22245,N_21993,N_21920);
and U22246 (N_22246,N_22163,N_22036);
nor U22247 (N_22247,N_21950,N_21918);
or U22248 (N_22248,N_22098,N_22196);
nor U22249 (N_22249,N_21949,N_22070);
xor U22250 (N_22250,N_22175,N_22143);
xnor U22251 (N_22251,N_21960,N_22166);
nand U22252 (N_22252,N_22050,N_22020);
and U22253 (N_22253,N_22035,N_21961);
or U22254 (N_22254,N_21968,N_21938);
xnor U22255 (N_22255,N_22022,N_21921);
nor U22256 (N_22256,N_22073,N_22101);
or U22257 (N_22257,N_22077,N_22108);
nor U22258 (N_22258,N_21919,N_22096);
and U22259 (N_22259,N_22113,N_21999);
xor U22260 (N_22260,N_22154,N_22081);
nor U22261 (N_22261,N_21964,N_21963);
or U22262 (N_22262,N_22177,N_22016);
and U22263 (N_22263,N_22122,N_22168);
nand U22264 (N_22264,N_22131,N_21923);
and U22265 (N_22265,N_22142,N_21976);
or U22266 (N_22266,N_22007,N_21959);
xor U22267 (N_22267,N_22117,N_22195);
nand U22268 (N_22268,N_21992,N_22049);
nand U22269 (N_22269,N_22160,N_21981);
or U22270 (N_22270,N_22118,N_21942);
and U22271 (N_22271,N_22120,N_22128);
nand U22272 (N_22272,N_21974,N_22172);
and U22273 (N_22273,N_22023,N_22074);
and U22274 (N_22274,N_22080,N_22024);
nand U22275 (N_22275,N_22009,N_21932);
nand U22276 (N_22276,N_22193,N_22002);
nand U22277 (N_22277,N_22097,N_22075);
or U22278 (N_22278,N_21930,N_21998);
nand U22279 (N_22279,N_21948,N_21904);
nor U22280 (N_22280,N_22183,N_22090);
xor U22281 (N_22281,N_22085,N_22173);
and U22282 (N_22282,N_22014,N_22192);
nand U22283 (N_22283,N_22086,N_22052);
nor U22284 (N_22284,N_21957,N_22064);
xnor U22285 (N_22285,N_22129,N_22124);
xnor U22286 (N_22286,N_21979,N_22025);
or U22287 (N_22287,N_22111,N_22018);
nand U22288 (N_22288,N_22058,N_21980);
or U22289 (N_22289,N_22087,N_21902);
nand U22290 (N_22290,N_21943,N_22088);
nand U22291 (N_22291,N_22162,N_22032);
xor U22292 (N_22292,N_21922,N_22062);
and U22293 (N_22293,N_21917,N_22040);
nand U22294 (N_22294,N_22167,N_22008);
or U22295 (N_22295,N_22141,N_22152);
nand U22296 (N_22296,N_22110,N_22010);
and U22297 (N_22297,N_21935,N_22198);
or U22298 (N_22298,N_21984,N_21997);
and U22299 (N_22299,N_21916,N_22093);
or U22300 (N_22300,N_22106,N_21933);
and U22301 (N_22301,N_22076,N_21978);
and U22302 (N_22302,N_22051,N_21944);
nor U22303 (N_22303,N_21945,N_22123);
nor U22304 (N_22304,N_22006,N_21909);
nor U22305 (N_22305,N_22092,N_22194);
nand U22306 (N_22306,N_22039,N_21996);
nand U22307 (N_22307,N_22047,N_22199);
or U22308 (N_22308,N_22156,N_21986);
xor U22309 (N_22309,N_22150,N_22119);
nor U22310 (N_22310,N_22144,N_22139);
xnor U22311 (N_22311,N_22126,N_21972);
nand U22312 (N_22312,N_22099,N_22013);
and U22313 (N_22313,N_22063,N_22029);
nor U22314 (N_22314,N_22148,N_21924);
and U22315 (N_22315,N_22161,N_21906);
xnor U22316 (N_22316,N_22181,N_21994);
nor U22317 (N_22317,N_21926,N_22048);
nand U22318 (N_22318,N_21927,N_22104);
and U22319 (N_22319,N_22053,N_22135);
nor U22320 (N_22320,N_22178,N_22153);
or U22321 (N_22321,N_21956,N_22003);
xor U22322 (N_22322,N_21910,N_22031);
nor U22323 (N_22323,N_22065,N_22159);
and U22324 (N_22324,N_22134,N_22079);
or U22325 (N_22325,N_22069,N_21901);
nor U22326 (N_22326,N_22095,N_22038);
nor U22327 (N_22327,N_22034,N_21937);
or U22328 (N_22328,N_22005,N_22091);
xor U22329 (N_22329,N_21955,N_22041);
or U22330 (N_22330,N_22182,N_22000);
nand U22331 (N_22331,N_22188,N_22026);
xnor U22332 (N_22332,N_21991,N_22084);
and U22333 (N_22333,N_22103,N_21940);
and U22334 (N_22334,N_22136,N_21936);
xor U22335 (N_22335,N_22067,N_22046);
nor U22336 (N_22336,N_21985,N_22180);
nand U22337 (N_22337,N_21912,N_22189);
nand U22338 (N_22338,N_22125,N_21928);
or U22339 (N_22339,N_21970,N_22105);
nand U22340 (N_22340,N_21931,N_22186);
nand U22341 (N_22341,N_21977,N_22100);
or U22342 (N_22342,N_22130,N_21951);
nand U22343 (N_22343,N_22137,N_21983);
xor U22344 (N_22344,N_22114,N_21934);
nor U22345 (N_22345,N_22115,N_21982);
nand U22346 (N_22346,N_21900,N_22071);
or U22347 (N_22347,N_22145,N_22066);
and U22348 (N_22348,N_21911,N_21971);
nand U22349 (N_22349,N_21939,N_22164);
and U22350 (N_22350,N_22154,N_21980);
nand U22351 (N_22351,N_22163,N_21937);
and U22352 (N_22352,N_22059,N_22172);
nand U22353 (N_22353,N_21945,N_22036);
nand U22354 (N_22354,N_21990,N_22115);
and U22355 (N_22355,N_21947,N_22055);
nand U22356 (N_22356,N_21917,N_22137);
nor U22357 (N_22357,N_22081,N_22149);
nor U22358 (N_22358,N_22137,N_22136);
and U22359 (N_22359,N_22144,N_22044);
nor U22360 (N_22360,N_22026,N_22080);
or U22361 (N_22361,N_22166,N_22024);
nand U22362 (N_22362,N_22149,N_22037);
or U22363 (N_22363,N_21975,N_22167);
nand U22364 (N_22364,N_22000,N_21919);
xnor U22365 (N_22365,N_22018,N_21937);
or U22366 (N_22366,N_21936,N_22198);
and U22367 (N_22367,N_21942,N_21935);
nand U22368 (N_22368,N_22098,N_22189);
and U22369 (N_22369,N_22126,N_22182);
xnor U22370 (N_22370,N_21940,N_22186);
nand U22371 (N_22371,N_22143,N_22063);
xor U22372 (N_22372,N_21952,N_22049);
and U22373 (N_22373,N_22044,N_22077);
or U22374 (N_22374,N_22092,N_22060);
and U22375 (N_22375,N_22047,N_21963);
nand U22376 (N_22376,N_22074,N_22039);
nand U22377 (N_22377,N_22087,N_22145);
nor U22378 (N_22378,N_22036,N_22166);
nand U22379 (N_22379,N_21983,N_21986);
nor U22380 (N_22380,N_21917,N_22054);
and U22381 (N_22381,N_21959,N_21949);
nand U22382 (N_22382,N_21920,N_22152);
or U22383 (N_22383,N_22084,N_21993);
and U22384 (N_22384,N_22025,N_21928);
nand U22385 (N_22385,N_22077,N_21958);
nand U22386 (N_22386,N_21941,N_22113);
xnor U22387 (N_22387,N_21953,N_21975);
or U22388 (N_22388,N_22024,N_21913);
and U22389 (N_22389,N_22014,N_21969);
and U22390 (N_22390,N_21919,N_22089);
xor U22391 (N_22391,N_22123,N_21971);
xnor U22392 (N_22392,N_22057,N_22036);
nor U22393 (N_22393,N_22095,N_21994);
or U22394 (N_22394,N_22110,N_22067);
nor U22395 (N_22395,N_22055,N_22064);
or U22396 (N_22396,N_22003,N_22079);
nor U22397 (N_22397,N_21947,N_22019);
and U22398 (N_22398,N_21940,N_22059);
and U22399 (N_22399,N_22064,N_22057);
or U22400 (N_22400,N_22099,N_21944);
or U22401 (N_22401,N_22063,N_22049);
nand U22402 (N_22402,N_22195,N_21954);
or U22403 (N_22403,N_22028,N_22162);
nand U22404 (N_22404,N_21970,N_21919);
and U22405 (N_22405,N_22117,N_22182);
xnor U22406 (N_22406,N_22085,N_22083);
xnor U22407 (N_22407,N_21970,N_22075);
or U22408 (N_22408,N_22087,N_22194);
and U22409 (N_22409,N_22127,N_22087);
nor U22410 (N_22410,N_22183,N_21957);
and U22411 (N_22411,N_21907,N_22110);
or U22412 (N_22412,N_22062,N_22191);
nand U22413 (N_22413,N_21987,N_22000);
and U22414 (N_22414,N_21921,N_22082);
xnor U22415 (N_22415,N_22079,N_22183);
xnor U22416 (N_22416,N_22011,N_21904);
or U22417 (N_22417,N_22198,N_22000);
and U22418 (N_22418,N_22103,N_21975);
or U22419 (N_22419,N_22191,N_22116);
xor U22420 (N_22420,N_22026,N_22025);
or U22421 (N_22421,N_22128,N_22112);
nor U22422 (N_22422,N_21952,N_22009);
xor U22423 (N_22423,N_21969,N_22119);
or U22424 (N_22424,N_21977,N_22065);
nor U22425 (N_22425,N_22195,N_22173);
and U22426 (N_22426,N_22036,N_21939);
nand U22427 (N_22427,N_22049,N_22173);
xnor U22428 (N_22428,N_22087,N_21900);
xor U22429 (N_22429,N_22050,N_22024);
nand U22430 (N_22430,N_22076,N_22186);
nand U22431 (N_22431,N_21984,N_22185);
and U22432 (N_22432,N_21920,N_22136);
or U22433 (N_22433,N_21905,N_21940);
nand U22434 (N_22434,N_21934,N_21991);
xnor U22435 (N_22435,N_22013,N_22050);
nand U22436 (N_22436,N_21972,N_22051);
nand U22437 (N_22437,N_21954,N_21947);
xnor U22438 (N_22438,N_22176,N_21986);
and U22439 (N_22439,N_22182,N_22077);
or U22440 (N_22440,N_21977,N_21922);
or U22441 (N_22441,N_22001,N_21911);
nor U22442 (N_22442,N_21914,N_22000);
xnor U22443 (N_22443,N_22103,N_22116);
or U22444 (N_22444,N_21926,N_21984);
and U22445 (N_22445,N_21987,N_21943);
or U22446 (N_22446,N_21969,N_21994);
and U22447 (N_22447,N_22112,N_22159);
xor U22448 (N_22448,N_21963,N_21965);
or U22449 (N_22449,N_21959,N_21979);
nand U22450 (N_22450,N_21975,N_22108);
or U22451 (N_22451,N_21950,N_21928);
nand U22452 (N_22452,N_22193,N_22014);
and U22453 (N_22453,N_21939,N_22191);
xnor U22454 (N_22454,N_21912,N_22126);
nand U22455 (N_22455,N_22190,N_22025);
and U22456 (N_22456,N_22130,N_22187);
nand U22457 (N_22457,N_22033,N_21991);
xor U22458 (N_22458,N_21948,N_22038);
or U22459 (N_22459,N_22089,N_21945);
xnor U22460 (N_22460,N_22052,N_22183);
or U22461 (N_22461,N_21902,N_21988);
and U22462 (N_22462,N_22145,N_22048);
nor U22463 (N_22463,N_21960,N_22143);
xnor U22464 (N_22464,N_22045,N_22025);
and U22465 (N_22465,N_22083,N_22109);
nor U22466 (N_22466,N_22060,N_21901);
nand U22467 (N_22467,N_22094,N_21929);
nor U22468 (N_22468,N_22071,N_22096);
xnor U22469 (N_22469,N_22195,N_22033);
nor U22470 (N_22470,N_22192,N_21909);
and U22471 (N_22471,N_22073,N_21920);
and U22472 (N_22472,N_21943,N_22142);
xnor U22473 (N_22473,N_22093,N_22178);
and U22474 (N_22474,N_22140,N_22152);
nor U22475 (N_22475,N_21976,N_22008);
and U22476 (N_22476,N_22098,N_22157);
and U22477 (N_22477,N_22110,N_21964);
or U22478 (N_22478,N_21915,N_22038);
nor U22479 (N_22479,N_22134,N_21972);
nor U22480 (N_22480,N_22087,N_22134);
and U22481 (N_22481,N_22022,N_21918);
and U22482 (N_22482,N_22032,N_22150);
xnor U22483 (N_22483,N_21924,N_21965);
xnor U22484 (N_22484,N_22148,N_21900);
and U22485 (N_22485,N_22161,N_22177);
and U22486 (N_22486,N_21916,N_21922);
nor U22487 (N_22487,N_22023,N_21916);
and U22488 (N_22488,N_22117,N_22143);
xor U22489 (N_22489,N_21949,N_22144);
nor U22490 (N_22490,N_21955,N_22012);
nor U22491 (N_22491,N_22131,N_22199);
nand U22492 (N_22492,N_22115,N_22130);
xnor U22493 (N_22493,N_22077,N_21919);
nand U22494 (N_22494,N_21971,N_22015);
and U22495 (N_22495,N_22013,N_22002);
xnor U22496 (N_22496,N_21992,N_22027);
xor U22497 (N_22497,N_22139,N_21946);
nor U22498 (N_22498,N_21928,N_21925);
nor U22499 (N_22499,N_22076,N_22137);
xor U22500 (N_22500,N_22442,N_22393);
xor U22501 (N_22501,N_22455,N_22367);
nor U22502 (N_22502,N_22214,N_22239);
nor U22503 (N_22503,N_22238,N_22211);
and U22504 (N_22504,N_22449,N_22324);
nand U22505 (N_22505,N_22496,N_22227);
nor U22506 (N_22506,N_22423,N_22312);
nor U22507 (N_22507,N_22244,N_22419);
xnor U22508 (N_22508,N_22241,N_22350);
nand U22509 (N_22509,N_22413,N_22495);
nand U22510 (N_22510,N_22381,N_22399);
xnor U22511 (N_22511,N_22437,N_22360);
or U22512 (N_22512,N_22424,N_22438);
and U22513 (N_22513,N_22240,N_22222);
xor U22514 (N_22514,N_22451,N_22255);
or U22515 (N_22515,N_22204,N_22328);
nor U22516 (N_22516,N_22409,N_22300);
or U22517 (N_22517,N_22220,N_22411);
nor U22518 (N_22518,N_22349,N_22362);
nor U22519 (N_22519,N_22269,N_22200);
or U22520 (N_22520,N_22281,N_22448);
xor U22521 (N_22521,N_22470,N_22256);
nand U22522 (N_22522,N_22389,N_22237);
nor U22523 (N_22523,N_22418,N_22277);
nor U22524 (N_22524,N_22215,N_22473);
or U22525 (N_22525,N_22407,N_22479);
or U22526 (N_22526,N_22388,N_22357);
and U22527 (N_22527,N_22391,N_22314);
nor U22528 (N_22528,N_22494,N_22348);
nand U22529 (N_22529,N_22242,N_22316);
nor U22530 (N_22530,N_22375,N_22342);
nand U22531 (N_22531,N_22422,N_22201);
nor U22532 (N_22532,N_22321,N_22489);
and U22533 (N_22533,N_22370,N_22374);
and U22534 (N_22534,N_22283,N_22229);
or U22535 (N_22535,N_22304,N_22412);
nand U22536 (N_22536,N_22271,N_22355);
and U22537 (N_22537,N_22309,N_22208);
or U22538 (N_22538,N_22297,N_22352);
or U22539 (N_22539,N_22450,N_22341);
and U22540 (N_22540,N_22274,N_22447);
and U22541 (N_22541,N_22441,N_22464);
xnor U22542 (N_22542,N_22245,N_22457);
or U22543 (N_22543,N_22408,N_22383);
or U22544 (N_22544,N_22394,N_22462);
nand U22545 (N_22545,N_22280,N_22278);
xor U22546 (N_22546,N_22392,N_22395);
xor U22547 (N_22547,N_22497,N_22267);
nand U22548 (N_22548,N_22251,N_22458);
and U22549 (N_22549,N_22212,N_22445);
or U22550 (N_22550,N_22368,N_22253);
and U22551 (N_22551,N_22425,N_22326);
and U22552 (N_22552,N_22365,N_22460);
xnor U22553 (N_22553,N_22317,N_22226);
or U22554 (N_22554,N_22366,N_22285);
nand U22555 (N_22555,N_22259,N_22275);
or U22556 (N_22556,N_22296,N_22380);
xor U22557 (N_22557,N_22405,N_22354);
and U22558 (N_22558,N_22288,N_22223);
nor U22559 (N_22559,N_22213,N_22416);
nor U22560 (N_22560,N_22377,N_22345);
xnor U22561 (N_22561,N_22301,N_22382);
nand U22562 (N_22562,N_22439,N_22401);
nand U22563 (N_22563,N_22295,N_22268);
and U22564 (N_22564,N_22363,N_22263);
and U22565 (N_22565,N_22216,N_22276);
and U22566 (N_22566,N_22475,N_22347);
xor U22567 (N_22567,N_22225,N_22453);
or U22568 (N_22568,N_22335,N_22353);
xnor U22569 (N_22569,N_22284,N_22480);
and U22570 (N_22570,N_22444,N_22247);
xnor U22571 (N_22571,N_22429,N_22273);
nor U22572 (N_22572,N_22398,N_22266);
xnor U22573 (N_22573,N_22290,N_22310);
or U22574 (N_22574,N_22327,N_22210);
and U22575 (N_22575,N_22440,N_22435);
nand U22576 (N_22576,N_22339,N_22236);
xnor U22577 (N_22577,N_22232,N_22318);
nand U22578 (N_22578,N_22415,N_22390);
nand U22579 (N_22579,N_22228,N_22233);
and U22580 (N_22580,N_22414,N_22485);
xor U22581 (N_22581,N_22490,N_22396);
nor U22582 (N_22582,N_22336,N_22378);
nand U22583 (N_22583,N_22334,N_22434);
or U22584 (N_22584,N_22488,N_22474);
nand U22585 (N_22585,N_22358,N_22446);
nor U22586 (N_22586,N_22376,N_22231);
or U22587 (N_22587,N_22406,N_22230);
nand U22588 (N_22588,N_22385,N_22346);
nor U22589 (N_22589,N_22203,N_22491);
nand U22590 (N_22590,N_22478,N_22484);
xnor U22591 (N_22591,N_22384,N_22487);
and U22592 (N_22592,N_22282,N_22330);
xnor U22593 (N_22593,N_22302,N_22252);
nand U22594 (N_22594,N_22426,N_22387);
and U22595 (N_22595,N_22308,N_22481);
nand U22596 (N_22596,N_22218,N_22331);
nor U22597 (N_22597,N_22463,N_22270);
nand U22598 (N_22598,N_22454,N_22471);
xor U22599 (N_22599,N_22207,N_22224);
and U22600 (N_22600,N_22249,N_22493);
and U22601 (N_22601,N_22325,N_22306);
and U22602 (N_22602,N_22291,N_22329);
nand U22603 (N_22603,N_22206,N_22427);
nor U22604 (N_22604,N_22492,N_22322);
or U22605 (N_22605,N_22307,N_22344);
nor U22606 (N_22606,N_22472,N_22286);
and U22607 (N_22607,N_22430,N_22234);
or U22608 (N_22608,N_22258,N_22202);
or U22609 (N_22609,N_22293,N_22265);
nand U22610 (N_22610,N_22372,N_22257);
nand U22611 (N_22611,N_22219,N_22467);
nor U22612 (N_22612,N_22364,N_22343);
nor U22613 (N_22613,N_22410,N_22217);
nor U22614 (N_22614,N_22459,N_22313);
or U22615 (N_22615,N_22303,N_22315);
and U22616 (N_22616,N_22351,N_22452);
and U22617 (N_22617,N_22209,N_22298);
and U22618 (N_22618,N_22433,N_22456);
nand U22619 (N_22619,N_22420,N_22264);
xor U22620 (N_22620,N_22404,N_22221);
or U22621 (N_22621,N_22469,N_22333);
nand U22622 (N_22622,N_22243,N_22261);
xnor U22623 (N_22623,N_22468,N_22287);
or U22624 (N_22624,N_22292,N_22465);
nor U22625 (N_22625,N_22466,N_22337);
and U22626 (N_22626,N_22299,N_22386);
nor U22627 (N_22627,N_22379,N_22432);
xor U22628 (N_22628,N_22428,N_22235);
xnor U22629 (N_22629,N_22323,N_22338);
xnor U22630 (N_22630,N_22289,N_22483);
nor U22631 (N_22631,N_22402,N_22205);
and U22632 (N_22632,N_22248,N_22498);
and U22633 (N_22633,N_22340,N_22476);
nand U22634 (N_22634,N_22294,N_22260);
nor U22635 (N_22635,N_22279,N_22320);
xnor U22636 (N_22636,N_22369,N_22400);
nand U22637 (N_22637,N_22477,N_22431);
or U22638 (N_22638,N_22482,N_22443);
or U22639 (N_22639,N_22305,N_22250);
xor U22640 (N_22640,N_22311,N_22371);
nor U22641 (N_22641,N_22421,N_22246);
or U22642 (N_22642,N_22262,N_22373);
or U22643 (N_22643,N_22361,N_22486);
or U22644 (N_22644,N_22332,N_22356);
and U22645 (N_22645,N_22272,N_22499);
nand U22646 (N_22646,N_22436,N_22403);
nand U22647 (N_22647,N_22359,N_22254);
nor U22648 (N_22648,N_22397,N_22319);
and U22649 (N_22649,N_22461,N_22417);
xnor U22650 (N_22650,N_22226,N_22239);
and U22651 (N_22651,N_22259,N_22266);
nand U22652 (N_22652,N_22398,N_22343);
nand U22653 (N_22653,N_22420,N_22329);
nor U22654 (N_22654,N_22416,N_22462);
nor U22655 (N_22655,N_22285,N_22356);
or U22656 (N_22656,N_22319,N_22271);
and U22657 (N_22657,N_22232,N_22312);
xor U22658 (N_22658,N_22313,N_22277);
and U22659 (N_22659,N_22400,N_22472);
nand U22660 (N_22660,N_22441,N_22449);
nor U22661 (N_22661,N_22320,N_22422);
or U22662 (N_22662,N_22451,N_22213);
nor U22663 (N_22663,N_22229,N_22263);
xor U22664 (N_22664,N_22284,N_22275);
or U22665 (N_22665,N_22351,N_22222);
or U22666 (N_22666,N_22233,N_22217);
xor U22667 (N_22667,N_22243,N_22377);
or U22668 (N_22668,N_22334,N_22219);
xor U22669 (N_22669,N_22420,N_22245);
nor U22670 (N_22670,N_22297,N_22346);
nand U22671 (N_22671,N_22418,N_22311);
nand U22672 (N_22672,N_22375,N_22455);
nand U22673 (N_22673,N_22333,N_22455);
or U22674 (N_22674,N_22356,N_22385);
and U22675 (N_22675,N_22458,N_22377);
xnor U22676 (N_22676,N_22275,N_22216);
or U22677 (N_22677,N_22443,N_22402);
and U22678 (N_22678,N_22357,N_22271);
and U22679 (N_22679,N_22334,N_22373);
or U22680 (N_22680,N_22430,N_22224);
or U22681 (N_22681,N_22330,N_22496);
nand U22682 (N_22682,N_22258,N_22440);
or U22683 (N_22683,N_22256,N_22214);
xor U22684 (N_22684,N_22225,N_22264);
and U22685 (N_22685,N_22485,N_22223);
or U22686 (N_22686,N_22373,N_22280);
nand U22687 (N_22687,N_22473,N_22382);
xor U22688 (N_22688,N_22418,N_22330);
and U22689 (N_22689,N_22488,N_22201);
and U22690 (N_22690,N_22429,N_22372);
and U22691 (N_22691,N_22481,N_22479);
nand U22692 (N_22692,N_22379,N_22218);
nor U22693 (N_22693,N_22332,N_22447);
or U22694 (N_22694,N_22475,N_22414);
or U22695 (N_22695,N_22472,N_22275);
or U22696 (N_22696,N_22389,N_22234);
nor U22697 (N_22697,N_22422,N_22352);
or U22698 (N_22698,N_22485,N_22408);
nand U22699 (N_22699,N_22472,N_22291);
or U22700 (N_22700,N_22260,N_22406);
nand U22701 (N_22701,N_22400,N_22450);
or U22702 (N_22702,N_22463,N_22457);
nand U22703 (N_22703,N_22285,N_22217);
nand U22704 (N_22704,N_22287,N_22221);
or U22705 (N_22705,N_22436,N_22265);
and U22706 (N_22706,N_22307,N_22426);
or U22707 (N_22707,N_22302,N_22438);
nor U22708 (N_22708,N_22385,N_22230);
or U22709 (N_22709,N_22375,N_22448);
nand U22710 (N_22710,N_22286,N_22242);
nand U22711 (N_22711,N_22446,N_22241);
nor U22712 (N_22712,N_22226,N_22303);
nand U22713 (N_22713,N_22315,N_22486);
xor U22714 (N_22714,N_22397,N_22243);
and U22715 (N_22715,N_22219,N_22312);
xnor U22716 (N_22716,N_22388,N_22251);
xor U22717 (N_22717,N_22211,N_22458);
nand U22718 (N_22718,N_22229,N_22242);
nand U22719 (N_22719,N_22495,N_22305);
xnor U22720 (N_22720,N_22406,N_22468);
nand U22721 (N_22721,N_22378,N_22321);
nor U22722 (N_22722,N_22488,N_22344);
xnor U22723 (N_22723,N_22349,N_22291);
or U22724 (N_22724,N_22319,N_22223);
and U22725 (N_22725,N_22283,N_22307);
or U22726 (N_22726,N_22386,N_22284);
or U22727 (N_22727,N_22311,N_22381);
nand U22728 (N_22728,N_22251,N_22268);
nand U22729 (N_22729,N_22218,N_22476);
or U22730 (N_22730,N_22419,N_22371);
or U22731 (N_22731,N_22436,N_22314);
and U22732 (N_22732,N_22418,N_22299);
nor U22733 (N_22733,N_22377,N_22358);
nand U22734 (N_22734,N_22462,N_22405);
nor U22735 (N_22735,N_22444,N_22464);
or U22736 (N_22736,N_22281,N_22288);
xnor U22737 (N_22737,N_22218,N_22213);
nand U22738 (N_22738,N_22302,N_22419);
nand U22739 (N_22739,N_22497,N_22459);
nand U22740 (N_22740,N_22310,N_22449);
xor U22741 (N_22741,N_22263,N_22341);
or U22742 (N_22742,N_22470,N_22434);
xnor U22743 (N_22743,N_22451,N_22217);
and U22744 (N_22744,N_22400,N_22409);
nor U22745 (N_22745,N_22367,N_22443);
nor U22746 (N_22746,N_22359,N_22263);
xor U22747 (N_22747,N_22443,N_22262);
or U22748 (N_22748,N_22286,N_22456);
and U22749 (N_22749,N_22235,N_22265);
xnor U22750 (N_22750,N_22467,N_22335);
or U22751 (N_22751,N_22405,N_22409);
and U22752 (N_22752,N_22329,N_22258);
and U22753 (N_22753,N_22371,N_22397);
nor U22754 (N_22754,N_22378,N_22464);
nor U22755 (N_22755,N_22274,N_22208);
nand U22756 (N_22756,N_22371,N_22493);
nand U22757 (N_22757,N_22258,N_22430);
or U22758 (N_22758,N_22289,N_22401);
nor U22759 (N_22759,N_22383,N_22407);
xnor U22760 (N_22760,N_22218,N_22310);
and U22761 (N_22761,N_22479,N_22226);
or U22762 (N_22762,N_22447,N_22386);
and U22763 (N_22763,N_22450,N_22470);
nor U22764 (N_22764,N_22331,N_22252);
xor U22765 (N_22765,N_22256,N_22434);
nand U22766 (N_22766,N_22222,N_22393);
or U22767 (N_22767,N_22274,N_22449);
xor U22768 (N_22768,N_22424,N_22439);
or U22769 (N_22769,N_22328,N_22472);
or U22770 (N_22770,N_22370,N_22211);
xor U22771 (N_22771,N_22227,N_22389);
or U22772 (N_22772,N_22307,N_22302);
xor U22773 (N_22773,N_22418,N_22410);
nand U22774 (N_22774,N_22226,N_22436);
xor U22775 (N_22775,N_22346,N_22443);
or U22776 (N_22776,N_22342,N_22285);
or U22777 (N_22777,N_22268,N_22312);
xor U22778 (N_22778,N_22224,N_22362);
or U22779 (N_22779,N_22408,N_22488);
xnor U22780 (N_22780,N_22369,N_22373);
nand U22781 (N_22781,N_22254,N_22309);
xnor U22782 (N_22782,N_22318,N_22497);
xor U22783 (N_22783,N_22351,N_22472);
nand U22784 (N_22784,N_22409,N_22292);
or U22785 (N_22785,N_22360,N_22209);
xnor U22786 (N_22786,N_22445,N_22248);
and U22787 (N_22787,N_22436,N_22366);
nand U22788 (N_22788,N_22301,N_22410);
xnor U22789 (N_22789,N_22377,N_22298);
nor U22790 (N_22790,N_22259,N_22323);
nand U22791 (N_22791,N_22464,N_22216);
nand U22792 (N_22792,N_22229,N_22284);
or U22793 (N_22793,N_22216,N_22490);
nor U22794 (N_22794,N_22344,N_22294);
xor U22795 (N_22795,N_22372,N_22238);
nor U22796 (N_22796,N_22271,N_22488);
xnor U22797 (N_22797,N_22441,N_22253);
or U22798 (N_22798,N_22258,N_22295);
and U22799 (N_22799,N_22436,N_22481);
nor U22800 (N_22800,N_22799,N_22525);
nor U22801 (N_22801,N_22742,N_22548);
nand U22802 (N_22802,N_22730,N_22700);
or U22803 (N_22803,N_22566,N_22579);
and U22804 (N_22804,N_22638,N_22738);
xnor U22805 (N_22805,N_22612,N_22643);
xor U22806 (N_22806,N_22685,N_22555);
xnor U22807 (N_22807,N_22721,N_22636);
xnor U22808 (N_22808,N_22739,N_22796);
nand U22809 (N_22809,N_22637,N_22653);
nand U22810 (N_22810,N_22659,N_22564);
or U22811 (N_22811,N_22681,N_22722);
nand U22812 (N_22812,N_22593,N_22763);
and U22813 (N_22813,N_22765,N_22667);
nand U22814 (N_22814,N_22590,N_22628);
and U22815 (N_22815,N_22797,N_22517);
and U22816 (N_22816,N_22544,N_22584);
xnor U22817 (N_22817,N_22668,N_22600);
xnor U22818 (N_22818,N_22791,N_22563);
xor U22819 (N_22819,N_22666,N_22746);
xor U22820 (N_22820,N_22758,N_22654);
and U22821 (N_22821,N_22727,N_22714);
and U22822 (N_22822,N_22633,N_22516);
or U22823 (N_22823,N_22617,N_22629);
nand U22824 (N_22824,N_22520,N_22538);
nor U22825 (N_22825,N_22705,N_22616);
and U22826 (N_22826,N_22788,N_22677);
nor U22827 (N_22827,N_22503,N_22792);
and U22828 (N_22828,N_22754,N_22652);
and U22829 (N_22829,N_22787,N_22686);
nand U22830 (N_22830,N_22562,N_22726);
xor U22831 (N_22831,N_22508,N_22597);
and U22832 (N_22832,N_22540,N_22692);
nand U22833 (N_22833,N_22728,N_22783);
nand U22834 (N_22834,N_22559,N_22610);
and U22835 (N_22835,N_22789,N_22713);
xnor U22836 (N_22836,N_22602,N_22743);
and U22837 (N_22837,N_22711,N_22569);
and U22838 (N_22838,N_22546,N_22771);
nor U22839 (N_22839,N_22646,N_22755);
xnor U22840 (N_22840,N_22620,N_22524);
nand U22841 (N_22841,N_22550,N_22752);
nand U22842 (N_22842,N_22679,N_22775);
nand U22843 (N_22843,N_22515,N_22545);
or U22844 (N_22844,N_22644,N_22585);
and U22845 (N_22845,N_22782,N_22675);
nor U22846 (N_22846,N_22634,N_22757);
nand U22847 (N_22847,N_22619,N_22598);
or U22848 (N_22848,N_22660,N_22756);
or U22849 (N_22849,N_22504,N_22794);
or U22850 (N_22850,N_22766,N_22541);
or U22851 (N_22851,N_22767,N_22561);
xor U22852 (N_22852,N_22717,N_22753);
and U22853 (N_22853,N_22725,N_22583);
nand U22854 (N_22854,N_22680,N_22734);
nand U22855 (N_22855,N_22737,N_22672);
or U22856 (N_22856,N_22608,N_22501);
nor U22857 (N_22857,N_22655,N_22708);
or U22858 (N_22858,N_22648,N_22786);
and U22859 (N_22859,N_22502,N_22773);
nand U22860 (N_22860,N_22568,N_22749);
and U22861 (N_22861,N_22622,N_22693);
or U22862 (N_22862,N_22580,N_22500);
and U22863 (N_22863,N_22573,N_22718);
nand U22864 (N_22864,N_22735,N_22678);
xnor U22865 (N_22865,N_22631,N_22647);
and U22866 (N_22866,N_22689,N_22640);
or U22867 (N_22867,N_22720,N_22736);
or U22868 (N_22868,N_22798,N_22691);
or U22869 (N_22869,N_22704,N_22707);
nand U22870 (N_22870,N_22549,N_22527);
and U22871 (N_22871,N_22509,N_22529);
xor U22872 (N_22872,N_22582,N_22656);
and U22873 (N_22873,N_22532,N_22710);
nor U22874 (N_22874,N_22603,N_22599);
xor U22875 (N_22875,N_22591,N_22657);
or U22876 (N_22876,N_22696,N_22649);
nor U22877 (N_22877,N_22770,N_22577);
or U22878 (N_22878,N_22557,N_22729);
and U22879 (N_22879,N_22611,N_22699);
nand U22880 (N_22880,N_22543,N_22618);
nand U22881 (N_22881,N_22687,N_22776);
nand U22882 (N_22882,N_22639,N_22748);
or U22883 (N_22883,N_22663,N_22642);
nor U22884 (N_22884,N_22510,N_22690);
xor U22885 (N_22885,N_22784,N_22790);
nor U22886 (N_22886,N_22609,N_22522);
nor U22887 (N_22887,N_22741,N_22641);
nor U22888 (N_22888,N_22526,N_22523);
and U22889 (N_22889,N_22570,N_22669);
and U22890 (N_22890,N_22625,N_22706);
or U22891 (N_22891,N_22596,N_22665);
nor U22892 (N_22892,N_22607,N_22632);
or U22893 (N_22893,N_22751,N_22781);
and U22894 (N_22894,N_22740,N_22712);
and U22895 (N_22895,N_22682,N_22627);
and U22896 (N_22896,N_22605,N_22575);
nor U22897 (N_22897,N_22507,N_22701);
and U22898 (N_22898,N_22733,N_22785);
nor U22899 (N_22899,N_22521,N_22780);
nand U22900 (N_22900,N_22614,N_22547);
and U22901 (N_22901,N_22592,N_22558);
nor U22902 (N_22902,N_22724,N_22578);
and U22903 (N_22903,N_22531,N_22553);
xor U22904 (N_22904,N_22601,N_22537);
xor U22905 (N_22905,N_22512,N_22554);
or U22906 (N_22906,N_22698,N_22664);
nor U22907 (N_22907,N_22574,N_22565);
nand U22908 (N_22908,N_22506,N_22626);
xor U22909 (N_22909,N_22604,N_22572);
xnor U22910 (N_22910,N_22581,N_22688);
nand U22911 (N_22911,N_22650,N_22764);
and U22912 (N_22912,N_22772,N_22542);
xor U22913 (N_22913,N_22630,N_22793);
or U22914 (N_22914,N_22539,N_22697);
or U22915 (N_22915,N_22536,N_22645);
xnor U22916 (N_22916,N_22768,N_22779);
or U22917 (N_22917,N_22658,N_22662);
and U22918 (N_22918,N_22694,N_22513);
or U22919 (N_22919,N_22535,N_22673);
nand U22920 (N_22920,N_22519,N_22576);
and U22921 (N_22921,N_22530,N_22511);
nand U22922 (N_22922,N_22719,N_22774);
xor U22923 (N_22923,N_22777,N_22560);
xnor U22924 (N_22924,N_22514,N_22744);
nand U22925 (N_22925,N_22621,N_22551);
and U22926 (N_22926,N_22761,N_22571);
nor U22927 (N_22927,N_22683,N_22635);
or U22928 (N_22928,N_22586,N_22518);
or U22929 (N_22929,N_22651,N_22613);
and U22930 (N_22930,N_22588,N_22589);
nor U22931 (N_22931,N_22715,N_22623);
and U22932 (N_22932,N_22702,N_22606);
nor U22933 (N_22933,N_22661,N_22595);
nand U22934 (N_22934,N_22533,N_22674);
nand U22935 (N_22935,N_22624,N_22716);
xor U22936 (N_22936,N_22594,N_22778);
nand U22937 (N_22937,N_22723,N_22795);
nand U22938 (N_22938,N_22505,N_22671);
and U22939 (N_22939,N_22747,N_22684);
or U22940 (N_22940,N_22769,N_22760);
or U22941 (N_22941,N_22759,N_22709);
or U22942 (N_22942,N_22703,N_22615);
nand U22943 (N_22943,N_22732,N_22552);
nor U22944 (N_22944,N_22762,N_22731);
xor U22945 (N_22945,N_22556,N_22587);
xnor U22946 (N_22946,N_22750,N_22695);
or U22947 (N_22947,N_22670,N_22534);
xor U22948 (N_22948,N_22528,N_22676);
nand U22949 (N_22949,N_22745,N_22567);
or U22950 (N_22950,N_22616,N_22675);
and U22951 (N_22951,N_22560,N_22586);
nor U22952 (N_22952,N_22787,N_22768);
nor U22953 (N_22953,N_22780,N_22510);
and U22954 (N_22954,N_22781,N_22730);
and U22955 (N_22955,N_22712,N_22590);
and U22956 (N_22956,N_22725,N_22798);
nand U22957 (N_22957,N_22779,N_22757);
and U22958 (N_22958,N_22722,N_22789);
nor U22959 (N_22959,N_22761,N_22590);
nand U22960 (N_22960,N_22788,N_22578);
and U22961 (N_22961,N_22638,N_22778);
and U22962 (N_22962,N_22772,N_22655);
or U22963 (N_22963,N_22505,N_22552);
xor U22964 (N_22964,N_22795,N_22701);
nor U22965 (N_22965,N_22792,N_22506);
or U22966 (N_22966,N_22565,N_22755);
nand U22967 (N_22967,N_22776,N_22752);
xnor U22968 (N_22968,N_22542,N_22601);
and U22969 (N_22969,N_22799,N_22776);
nand U22970 (N_22970,N_22530,N_22549);
nand U22971 (N_22971,N_22503,N_22743);
nor U22972 (N_22972,N_22741,N_22765);
and U22973 (N_22973,N_22663,N_22558);
and U22974 (N_22974,N_22583,N_22545);
xor U22975 (N_22975,N_22757,N_22539);
or U22976 (N_22976,N_22751,N_22671);
and U22977 (N_22977,N_22587,N_22751);
xor U22978 (N_22978,N_22726,N_22572);
xor U22979 (N_22979,N_22759,N_22776);
and U22980 (N_22980,N_22534,N_22568);
xnor U22981 (N_22981,N_22557,N_22525);
nand U22982 (N_22982,N_22685,N_22786);
nor U22983 (N_22983,N_22759,N_22644);
nand U22984 (N_22984,N_22773,N_22587);
and U22985 (N_22985,N_22694,N_22762);
nand U22986 (N_22986,N_22713,N_22524);
nor U22987 (N_22987,N_22740,N_22588);
and U22988 (N_22988,N_22665,N_22759);
or U22989 (N_22989,N_22507,N_22558);
and U22990 (N_22990,N_22778,N_22728);
or U22991 (N_22991,N_22685,N_22622);
or U22992 (N_22992,N_22773,N_22788);
and U22993 (N_22993,N_22707,N_22505);
xnor U22994 (N_22994,N_22741,N_22624);
nand U22995 (N_22995,N_22655,N_22559);
nor U22996 (N_22996,N_22794,N_22532);
nand U22997 (N_22997,N_22764,N_22638);
nand U22998 (N_22998,N_22774,N_22748);
or U22999 (N_22999,N_22509,N_22527);
nand U23000 (N_23000,N_22720,N_22783);
nand U23001 (N_23001,N_22678,N_22563);
nor U23002 (N_23002,N_22798,N_22553);
and U23003 (N_23003,N_22669,N_22722);
and U23004 (N_23004,N_22633,N_22507);
xor U23005 (N_23005,N_22526,N_22572);
and U23006 (N_23006,N_22621,N_22631);
or U23007 (N_23007,N_22745,N_22523);
or U23008 (N_23008,N_22668,N_22579);
nor U23009 (N_23009,N_22683,N_22652);
nand U23010 (N_23010,N_22683,N_22772);
xnor U23011 (N_23011,N_22541,N_22608);
nor U23012 (N_23012,N_22687,N_22714);
or U23013 (N_23013,N_22748,N_22768);
xnor U23014 (N_23014,N_22631,N_22618);
or U23015 (N_23015,N_22633,N_22691);
nor U23016 (N_23016,N_22551,N_22754);
nand U23017 (N_23017,N_22525,N_22717);
xnor U23018 (N_23018,N_22633,N_22558);
and U23019 (N_23019,N_22593,N_22798);
or U23020 (N_23020,N_22717,N_22559);
nand U23021 (N_23021,N_22654,N_22583);
nor U23022 (N_23022,N_22725,N_22641);
nor U23023 (N_23023,N_22797,N_22574);
nand U23024 (N_23024,N_22791,N_22550);
and U23025 (N_23025,N_22653,N_22552);
nand U23026 (N_23026,N_22656,N_22635);
nand U23027 (N_23027,N_22628,N_22593);
and U23028 (N_23028,N_22524,N_22588);
or U23029 (N_23029,N_22687,N_22653);
nand U23030 (N_23030,N_22692,N_22605);
and U23031 (N_23031,N_22606,N_22581);
and U23032 (N_23032,N_22641,N_22696);
nor U23033 (N_23033,N_22780,N_22659);
and U23034 (N_23034,N_22564,N_22701);
and U23035 (N_23035,N_22638,N_22510);
and U23036 (N_23036,N_22517,N_22533);
nand U23037 (N_23037,N_22582,N_22786);
xnor U23038 (N_23038,N_22517,N_22638);
nor U23039 (N_23039,N_22515,N_22783);
or U23040 (N_23040,N_22585,N_22588);
xnor U23041 (N_23041,N_22515,N_22566);
nor U23042 (N_23042,N_22632,N_22686);
xnor U23043 (N_23043,N_22578,N_22596);
nand U23044 (N_23044,N_22604,N_22656);
nor U23045 (N_23045,N_22666,N_22596);
xor U23046 (N_23046,N_22597,N_22659);
or U23047 (N_23047,N_22668,N_22720);
xnor U23048 (N_23048,N_22579,N_22772);
xor U23049 (N_23049,N_22593,N_22569);
and U23050 (N_23050,N_22665,N_22671);
or U23051 (N_23051,N_22655,N_22741);
xor U23052 (N_23052,N_22789,N_22609);
xor U23053 (N_23053,N_22692,N_22539);
nor U23054 (N_23054,N_22604,N_22754);
xnor U23055 (N_23055,N_22753,N_22514);
and U23056 (N_23056,N_22791,N_22769);
and U23057 (N_23057,N_22557,N_22786);
nor U23058 (N_23058,N_22526,N_22586);
and U23059 (N_23059,N_22718,N_22526);
nor U23060 (N_23060,N_22777,N_22515);
xor U23061 (N_23061,N_22727,N_22524);
or U23062 (N_23062,N_22607,N_22619);
nand U23063 (N_23063,N_22616,N_22662);
and U23064 (N_23064,N_22784,N_22719);
xnor U23065 (N_23065,N_22753,N_22564);
and U23066 (N_23066,N_22685,N_22571);
nand U23067 (N_23067,N_22665,N_22757);
and U23068 (N_23068,N_22523,N_22564);
nand U23069 (N_23069,N_22769,N_22765);
or U23070 (N_23070,N_22791,N_22684);
and U23071 (N_23071,N_22709,N_22583);
nand U23072 (N_23072,N_22765,N_22548);
and U23073 (N_23073,N_22597,N_22540);
nand U23074 (N_23074,N_22510,N_22591);
nand U23075 (N_23075,N_22676,N_22661);
nand U23076 (N_23076,N_22520,N_22516);
and U23077 (N_23077,N_22656,N_22710);
nand U23078 (N_23078,N_22736,N_22781);
nand U23079 (N_23079,N_22501,N_22746);
nor U23080 (N_23080,N_22787,N_22640);
nand U23081 (N_23081,N_22534,N_22557);
xor U23082 (N_23082,N_22707,N_22764);
nor U23083 (N_23083,N_22579,N_22750);
nor U23084 (N_23084,N_22672,N_22744);
nor U23085 (N_23085,N_22519,N_22633);
or U23086 (N_23086,N_22707,N_22580);
nor U23087 (N_23087,N_22796,N_22680);
nand U23088 (N_23088,N_22776,N_22786);
xnor U23089 (N_23089,N_22601,N_22505);
and U23090 (N_23090,N_22609,N_22539);
or U23091 (N_23091,N_22607,N_22766);
nand U23092 (N_23092,N_22528,N_22583);
and U23093 (N_23093,N_22673,N_22720);
nor U23094 (N_23094,N_22548,N_22575);
and U23095 (N_23095,N_22616,N_22720);
xnor U23096 (N_23096,N_22588,N_22577);
nand U23097 (N_23097,N_22560,N_22684);
nor U23098 (N_23098,N_22562,N_22630);
nand U23099 (N_23099,N_22786,N_22525);
and U23100 (N_23100,N_22958,N_22933);
xnor U23101 (N_23101,N_22986,N_22938);
and U23102 (N_23102,N_23000,N_22898);
and U23103 (N_23103,N_22832,N_23086);
xnor U23104 (N_23104,N_23044,N_22939);
or U23105 (N_23105,N_22825,N_22871);
nor U23106 (N_23106,N_22922,N_22889);
or U23107 (N_23107,N_22847,N_22904);
or U23108 (N_23108,N_22801,N_22979);
or U23109 (N_23109,N_23068,N_22924);
xor U23110 (N_23110,N_22872,N_22823);
or U23111 (N_23111,N_22987,N_22921);
nor U23112 (N_23112,N_22900,N_23015);
nand U23113 (N_23113,N_22945,N_22960);
nand U23114 (N_23114,N_22976,N_23056);
nor U23115 (N_23115,N_22919,N_22994);
or U23116 (N_23116,N_22892,N_22881);
nand U23117 (N_23117,N_23058,N_22884);
xnor U23118 (N_23118,N_23007,N_22999);
and U23119 (N_23119,N_22967,N_22951);
and U23120 (N_23120,N_22948,N_22836);
and U23121 (N_23121,N_22842,N_22962);
xnor U23122 (N_23122,N_23064,N_22983);
nand U23123 (N_23123,N_23005,N_23006);
nor U23124 (N_23124,N_22895,N_22863);
and U23125 (N_23125,N_22966,N_22804);
and U23126 (N_23126,N_22981,N_22866);
and U23127 (N_23127,N_23085,N_22918);
nand U23128 (N_23128,N_22995,N_23089);
and U23129 (N_23129,N_22879,N_22899);
nor U23130 (N_23130,N_22998,N_22943);
nand U23131 (N_23131,N_23075,N_23011);
nand U23132 (N_23132,N_22838,N_22851);
nand U23133 (N_23133,N_22920,N_23087);
xnor U23134 (N_23134,N_22868,N_22839);
and U23135 (N_23135,N_23041,N_22810);
and U23136 (N_23136,N_22885,N_23072);
and U23137 (N_23137,N_22867,N_23012);
xnor U23138 (N_23138,N_22935,N_22852);
nor U23139 (N_23139,N_23029,N_23091);
or U23140 (N_23140,N_22860,N_22806);
nor U23141 (N_23141,N_22803,N_22854);
and U23142 (N_23142,N_23059,N_23039);
xor U23143 (N_23143,N_22876,N_23022);
nand U23144 (N_23144,N_22974,N_22934);
xnor U23145 (N_23145,N_23051,N_22993);
or U23146 (N_23146,N_23081,N_23098);
nand U23147 (N_23147,N_22901,N_23082);
and U23148 (N_23148,N_22843,N_22833);
or U23149 (N_23149,N_22941,N_22848);
xnor U23150 (N_23150,N_23099,N_22965);
xnor U23151 (N_23151,N_22950,N_22902);
and U23152 (N_23152,N_22942,N_23020);
nor U23153 (N_23153,N_22864,N_22980);
or U23154 (N_23154,N_22856,N_22984);
nand U23155 (N_23155,N_23001,N_23031);
or U23156 (N_23156,N_23066,N_22953);
and U23157 (N_23157,N_23071,N_23037);
nor U23158 (N_23158,N_22813,N_22946);
nor U23159 (N_23159,N_22831,N_22952);
or U23160 (N_23160,N_22858,N_22887);
and U23161 (N_23161,N_22862,N_22957);
nor U23162 (N_23162,N_23028,N_23009);
nor U23163 (N_23163,N_23014,N_22816);
or U23164 (N_23164,N_22956,N_22834);
and U23165 (N_23165,N_23035,N_23030);
and U23166 (N_23166,N_23010,N_23073);
nand U23167 (N_23167,N_22882,N_23033);
nand U23168 (N_23168,N_22971,N_22961);
nor U23169 (N_23169,N_22877,N_23084);
or U23170 (N_23170,N_22928,N_22857);
and U23171 (N_23171,N_22909,N_23062);
and U23172 (N_23172,N_22844,N_22869);
nand U23173 (N_23173,N_23003,N_22824);
xor U23174 (N_23174,N_22908,N_23026);
nor U23175 (N_23175,N_22988,N_23079);
or U23176 (N_23176,N_22989,N_23002);
nor U23177 (N_23177,N_22947,N_23097);
and U23178 (N_23178,N_22944,N_22954);
nand U23179 (N_23179,N_22968,N_22894);
nor U23180 (N_23180,N_22821,N_23050);
nand U23181 (N_23181,N_23018,N_22932);
xnor U23182 (N_23182,N_22923,N_22883);
nor U23183 (N_23183,N_22907,N_22893);
xnor U23184 (N_23184,N_23083,N_23040);
xor U23185 (N_23185,N_22875,N_22817);
nand U23186 (N_23186,N_23090,N_22859);
or U23187 (N_23187,N_22930,N_22814);
and U23188 (N_23188,N_22982,N_22916);
and U23189 (N_23189,N_23055,N_22931);
nand U23190 (N_23190,N_22914,N_23060);
nand U23191 (N_23191,N_22903,N_22978);
or U23192 (N_23192,N_22913,N_23063);
or U23193 (N_23193,N_23065,N_22815);
nand U23194 (N_23194,N_23076,N_22840);
or U23195 (N_23195,N_23027,N_22926);
nand U23196 (N_23196,N_23094,N_22853);
nand U23197 (N_23197,N_22972,N_22969);
nor U23198 (N_23198,N_22973,N_22874);
nor U23199 (N_23199,N_22997,N_22812);
or U23200 (N_23200,N_23088,N_23017);
nand U23201 (N_23201,N_22873,N_23046);
or U23202 (N_23202,N_23034,N_23008);
and U23203 (N_23203,N_22990,N_23057);
and U23204 (N_23204,N_22837,N_22925);
nor U23205 (N_23205,N_23021,N_22975);
nand U23206 (N_23206,N_22805,N_23048);
xnor U23207 (N_23207,N_22897,N_22829);
and U23208 (N_23208,N_22802,N_22964);
nor U23209 (N_23209,N_23042,N_23067);
xor U23210 (N_23210,N_22861,N_22917);
nor U23211 (N_23211,N_23053,N_23016);
nand U23212 (N_23212,N_22992,N_23023);
xor U23213 (N_23213,N_22955,N_22808);
and U23214 (N_23214,N_22828,N_22819);
nor U23215 (N_23215,N_22886,N_22830);
nand U23216 (N_23216,N_23074,N_22991);
xor U23217 (N_23217,N_23019,N_23092);
and U23218 (N_23218,N_23043,N_22940);
xor U23219 (N_23219,N_23025,N_22949);
nand U23220 (N_23220,N_23095,N_22985);
and U23221 (N_23221,N_22850,N_23049);
nor U23222 (N_23222,N_22927,N_22809);
nand U23223 (N_23223,N_22878,N_22977);
xnor U23224 (N_23224,N_22890,N_23038);
nor U23225 (N_23225,N_22963,N_22912);
and U23226 (N_23226,N_22905,N_22959);
nor U23227 (N_23227,N_23054,N_22929);
and U23228 (N_23228,N_22936,N_22915);
nand U23229 (N_23229,N_22800,N_23069);
nand U23230 (N_23230,N_22846,N_22937);
or U23231 (N_23231,N_23032,N_22911);
nor U23232 (N_23232,N_23078,N_22841);
xnor U23233 (N_23233,N_22906,N_22891);
or U23234 (N_23234,N_23096,N_23070);
and U23235 (N_23235,N_23080,N_23061);
nor U23236 (N_23236,N_23045,N_22896);
and U23237 (N_23237,N_23047,N_22849);
and U23238 (N_23238,N_22811,N_23077);
nand U23239 (N_23239,N_22910,N_22835);
xnor U23240 (N_23240,N_23013,N_23024);
xnor U23241 (N_23241,N_23036,N_22820);
nor U23242 (N_23242,N_22807,N_22845);
and U23243 (N_23243,N_22826,N_23093);
nand U23244 (N_23244,N_22880,N_22888);
nand U23245 (N_23245,N_22970,N_22865);
and U23246 (N_23246,N_22827,N_23004);
xnor U23247 (N_23247,N_22870,N_22855);
and U23248 (N_23248,N_23052,N_22818);
and U23249 (N_23249,N_22996,N_22822);
or U23250 (N_23250,N_22847,N_22996);
nor U23251 (N_23251,N_23049,N_22827);
or U23252 (N_23252,N_22992,N_22826);
or U23253 (N_23253,N_22879,N_22972);
or U23254 (N_23254,N_22998,N_23071);
nor U23255 (N_23255,N_22933,N_22936);
and U23256 (N_23256,N_23018,N_22909);
nand U23257 (N_23257,N_22806,N_23004);
xnor U23258 (N_23258,N_23099,N_22955);
and U23259 (N_23259,N_22899,N_23093);
xnor U23260 (N_23260,N_22889,N_22854);
nor U23261 (N_23261,N_23056,N_23075);
xnor U23262 (N_23262,N_22961,N_22972);
nand U23263 (N_23263,N_23054,N_23080);
xor U23264 (N_23264,N_23021,N_22805);
or U23265 (N_23265,N_22934,N_23008);
and U23266 (N_23266,N_22955,N_22967);
nand U23267 (N_23267,N_22843,N_22847);
and U23268 (N_23268,N_22954,N_22936);
nand U23269 (N_23269,N_22875,N_22833);
and U23270 (N_23270,N_22973,N_22803);
xnor U23271 (N_23271,N_23005,N_22881);
xor U23272 (N_23272,N_23054,N_22836);
xnor U23273 (N_23273,N_22956,N_22866);
xnor U23274 (N_23274,N_22870,N_23027);
and U23275 (N_23275,N_22819,N_22982);
nand U23276 (N_23276,N_22919,N_22998);
nor U23277 (N_23277,N_23069,N_22818);
xor U23278 (N_23278,N_23009,N_22880);
or U23279 (N_23279,N_23042,N_23034);
xnor U23280 (N_23280,N_22822,N_22922);
xnor U23281 (N_23281,N_22920,N_23079);
and U23282 (N_23282,N_22901,N_22922);
and U23283 (N_23283,N_22988,N_22831);
and U23284 (N_23284,N_22843,N_22961);
nand U23285 (N_23285,N_23045,N_22903);
nand U23286 (N_23286,N_23041,N_22976);
and U23287 (N_23287,N_22916,N_23014);
xnor U23288 (N_23288,N_22902,N_22841);
nand U23289 (N_23289,N_22882,N_23083);
nand U23290 (N_23290,N_23093,N_22874);
xor U23291 (N_23291,N_22871,N_23078);
and U23292 (N_23292,N_22987,N_22846);
or U23293 (N_23293,N_22882,N_22801);
xor U23294 (N_23294,N_22886,N_22945);
nor U23295 (N_23295,N_22853,N_22809);
nor U23296 (N_23296,N_22825,N_22920);
or U23297 (N_23297,N_22911,N_23019);
xnor U23298 (N_23298,N_23026,N_23006);
or U23299 (N_23299,N_23092,N_22895);
and U23300 (N_23300,N_22836,N_23032);
nor U23301 (N_23301,N_22920,N_22873);
or U23302 (N_23302,N_22842,N_22888);
nand U23303 (N_23303,N_22840,N_22986);
or U23304 (N_23304,N_23073,N_22866);
or U23305 (N_23305,N_22936,N_23022);
nor U23306 (N_23306,N_22919,N_22895);
xnor U23307 (N_23307,N_23098,N_23034);
and U23308 (N_23308,N_22905,N_22842);
nor U23309 (N_23309,N_22819,N_22919);
nand U23310 (N_23310,N_23035,N_22933);
xor U23311 (N_23311,N_22878,N_22963);
xnor U23312 (N_23312,N_22971,N_23034);
nor U23313 (N_23313,N_22847,N_23079);
nor U23314 (N_23314,N_22987,N_23053);
xnor U23315 (N_23315,N_22859,N_22875);
or U23316 (N_23316,N_22915,N_22944);
and U23317 (N_23317,N_23073,N_22809);
and U23318 (N_23318,N_22839,N_22912);
and U23319 (N_23319,N_23064,N_23075);
nand U23320 (N_23320,N_22863,N_22825);
xnor U23321 (N_23321,N_22908,N_22961);
and U23322 (N_23322,N_23034,N_23060);
and U23323 (N_23323,N_22841,N_23097);
and U23324 (N_23324,N_23067,N_22895);
nand U23325 (N_23325,N_23034,N_22829);
and U23326 (N_23326,N_22930,N_22819);
nand U23327 (N_23327,N_23020,N_22824);
or U23328 (N_23328,N_22806,N_22892);
or U23329 (N_23329,N_22910,N_22964);
nor U23330 (N_23330,N_22917,N_22879);
nand U23331 (N_23331,N_23065,N_22886);
xor U23332 (N_23332,N_22957,N_22800);
and U23333 (N_23333,N_22993,N_23082);
or U23334 (N_23334,N_23053,N_23036);
xnor U23335 (N_23335,N_22878,N_23003);
or U23336 (N_23336,N_22874,N_22805);
xnor U23337 (N_23337,N_22829,N_22836);
xor U23338 (N_23338,N_22801,N_22912);
or U23339 (N_23339,N_23083,N_22800);
and U23340 (N_23340,N_22940,N_23032);
nand U23341 (N_23341,N_23096,N_22827);
nand U23342 (N_23342,N_22877,N_23067);
or U23343 (N_23343,N_22982,N_22874);
nor U23344 (N_23344,N_22850,N_23077);
xnor U23345 (N_23345,N_23034,N_22839);
nand U23346 (N_23346,N_22913,N_22870);
and U23347 (N_23347,N_22927,N_22847);
nand U23348 (N_23348,N_22852,N_22988);
or U23349 (N_23349,N_22835,N_22809);
nor U23350 (N_23350,N_22923,N_23024);
nor U23351 (N_23351,N_22828,N_22823);
or U23352 (N_23352,N_22813,N_23022);
nand U23353 (N_23353,N_22943,N_22938);
nor U23354 (N_23354,N_22963,N_22919);
and U23355 (N_23355,N_22802,N_22963);
nand U23356 (N_23356,N_22888,N_22836);
and U23357 (N_23357,N_23022,N_22841);
and U23358 (N_23358,N_22913,N_22973);
and U23359 (N_23359,N_22804,N_23014);
or U23360 (N_23360,N_22977,N_23093);
and U23361 (N_23361,N_23008,N_23096);
or U23362 (N_23362,N_22887,N_22919);
or U23363 (N_23363,N_23006,N_22910);
xor U23364 (N_23364,N_22993,N_23000);
and U23365 (N_23365,N_22824,N_23077);
or U23366 (N_23366,N_22995,N_23086);
or U23367 (N_23367,N_23082,N_23041);
xnor U23368 (N_23368,N_22847,N_23072);
nand U23369 (N_23369,N_22964,N_23027);
or U23370 (N_23370,N_22842,N_23071);
and U23371 (N_23371,N_22855,N_23054);
nand U23372 (N_23372,N_22873,N_22836);
xnor U23373 (N_23373,N_22822,N_22917);
nor U23374 (N_23374,N_22928,N_22892);
nor U23375 (N_23375,N_22994,N_22804);
nor U23376 (N_23376,N_22893,N_22966);
and U23377 (N_23377,N_23050,N_23077);
nor U23378 (N_23378,N_22880,N_22905);
or U23379 (N_23379,N_22828,N_23012);
nand U23380 (N_23380,N_22813,N_23068);
nor U23381 (N_23381,N_23013,N_22888);
nand U23382 (N_23382,N_22951,N_22811);
xor U23383 (N_23383,N_22866,N_22835);
or U23384 (N_23384,N_22802,N_22973);
nor U23385 (N_23385,N_23026,N_23080);
xor U23386 (N_23386,N_22940,N_22997);
and U23387 (N_23387,N_22826,N_22946);
nor U23388 (N_23388,N_22933,N_22916);
xor U23389 (N_23389,N_22909,N_22824);
xnor U23390 (N_23390,N_22999,N_22900);
nor U23391 (N_23391,N_22853,N_22892);
and U23392 (N_23392,N_22824,N_22940);
nand U23393 (N_23393,N_22837,N_22851);
nor U23394 (N_23394,N_23000,N_22882);
nand U23395 (N_23395,N_23018,N_22813);
xor U23396 (N_23396,N_22933,N_23065);
xnor U23397 (N_23397,N_22918,N_22872);
nand U23398 (N_23398,N_23000,N_22809);
or U23399 (N_23399,N_23011,N_22874);
nand U23400 (N_23400,N_23335,N_23342);
and U23401 (N_23401,N_23229,N_23140);
and U23402 (N_23402,N_23111,N_23239);
xor U23403 (N_23403,N_23274,N_23112);
nand U23404 (N_23404,N_23398,N_23392);
and U23405 (N_23405,N_23197,N_23366);
nand U23406 (N_23406,N_23269,N_23250);
and U23407 (N_23407,N_23211,N_23288);
nand U23408 (N_23408,N_23178,N_23100);
or U23409 (N_23409,N_23322,N_23196);
nand U23410 (N_23410,N_23109,N_23209);
nand U23411 (N_23411,N_23117,N_23388);
nand U23412 (N_23412,N_23202,N_23205);
xnor U23413 (N_23413,N_23175,N_23304);
nor U23414 (N_23414,N_23358,N_23270);
nor U23415 (N_23415,N_23146,N_23360);
or U23416 (N_23416,N_23373,N_23198);
xnor U23417 (N_23417,N_23216,N_23259);
nor U23418 (N_23418,N_23253,N_23236);
or U23419 (N_23419,N_23218,N_23230);
nor U23420 (N_23420,N_23130,N_23351);
and U23421 (N_23421,N_23272,N_23164);
nor U23422 (N_23422,N_23354,N_23278);
nor U23423 (N_23423,N_23154,N_23357);
and U23424 (N_23424,N_23161,N_23371);
nor U23425 (N_23425,N_23310,N_23103);
nand U23426 (N_23426,N_23325,N_23138);
xnor U23427 (N_23427,N_23153,N_23247);
nand U23428 (N_23428,N_23150,N_23252);
nor U23429 (N_23429,N_23372,N_23382);
xor U23430 (N_23430,N_23330,N_23386);
nor U23431 (N_23431,N_23306,N_23381);
or U23432 (N_23432,N_23394,N_23170);
or U23433 (N_23433,N_23345,N_23350);
and U23434 (N_23434,N_23263,N_23167);
xor U23435 (N_23435,N_23148,N_23266);
nand U23436 (N_23436,N_23181,N_23344);
nor U23437 (N_23437,N_23273,N_23115);
xnor U23438 (N_23438,N_23258,N_23171);
nor U23439 (N_23439,N_23316,N_23141);
nand U23440 (N_23440,N_23353,N_23152);
nor U23441 (N_23441,N_23192,N_23346);
nor U23442 (N_23442,N_23245,N_23110);
nand U23443 (N_23443,N_23367,N_23318);
xnor U23444 (N_23444,N_23169,N_23241);
or U23445 (N_23445,N_23219,N_23231);
and U23446 (N_23446,N_23395,N_23389);
nand U23447 (N_23447,N_23213,N_23251);
nor U23448 (N_23448,N_23396,N_23340);
or U23449 (N_23449,N_23133,N_23280);
nand U23450 (N_23450,N_23299,N_23294);
xnor U23451 (N_23451,N_23285,N_23293);
nand U23452 (N_23452,N_23369,N_23162);
nand U23453 (N_23453,N_23297,N_23200);
nand U23454 (N_23454,N_23352,N_23127);
nand U23455 (N_23455,N_23276,N_23107);
nand U23456 (N_23456,N_23361,N_23208);
or U23457 (N_23457,N_23290,N_23317);
and U23458 (N_23458,N_23365,N_23159);
xnor U23459 (N_23459,N_23124,N_23101);
and U23460 (N_23460,N_23244,N_23234);
xnor U23461 (N_23461,N_23179,N_23256);
xnor U23462 (N_23462,N_23185,N_23217);
nand U23463 (N_23463,N_23207,N_23182);
nor U23464 (N_23464,N_23172,N_23116);
nand U23465 (N_23465,N_23158,N_23149);
nand U23466 (N_23466,N_23206,N_23260);
nand U23467 (N_23467,N_23289,N_23291);
nor U23468 (N_23468,N_23163,N_23257);
nor U23469 (N_23469,N_23343,N_23300);
or U23470 (N_23470,N_23254,N_23393);
or U23471 (N_23471,N_23368,N_23189);
and U23472 (N_23472,N_23199,N_23370);
nor U23473 (N_23473,N_23194,N_23377);
or U23474 (N_23474,N_23271,N_23337);
xnor U23475 (N_23475,N_23364,N_23120);
nand U23476 (N_23476,N_23186,N_23378);
xnor U23477 (N_23477,N_23312,N_23104);
nand U23478 (N_23478,N_23264,N_23336);
or U23479 (N_23479,N_23246,N_23320);
or U23480 (N_23480,N_23220,N_23242);
or U23481 (N_23481,N_23331,N_23145);
xor U23482 (N_23482,N_23321,N_23296);
nand U23483 (N_23483,N_23237,N_23379);
or U23484 (N_23484,N_23383,N_23298);
xor U23485 (N_23485,N_23166,N_23118);
nand U23486 (N_23486,N_23284,N_23349);
nand U23487 (N_23487,N_23384,N_23305);
xnor U23488 (N_23488,N_23238,N_23160);
or U23489 (N_23489,N_23249,N_23292);
xor U23490 (N_23490,N_23212,N_23108);
or U23491 (N_23491,N_23341,N_23123);
xnor U23492 (N_23492,N_23329,N_23232);
or U23493 (N_23493,N_23262,N_23201);
nand U23494 (N_23494,N_23286,N_23210);
and U23495 (N_23495,N_23225,N_23282);
and U23496 (N_23496,N_23319,N_23339);
nor U23497 (N_23497,N_23183,N_23326);
or U23498 (N_23498,N_23122,N_23314);
nand U23499 (N_23499,N_23307,N_23356);
nand U23500 (N_23500,N_23265,N_23151);
and U23501 (N_23501,N_23363,N_23390);
and U23502 (N_23502,N_23126,N_23177);
xnor U23503 (N_23503,N_23157,N_23303);
xnor U23504 (N_23504,N_23311,N_23195);
and U23505 (N_23505,N_23135,N_23333);
and U23506 (N_23506,N_23188,N_23180);
or U23507 (N_23507,N_23355,N_23334);
and U23508 (N_23508,N_23184,N_23332);
xor U23509 (N_23509,N_23248,N_23295);
or U23510 (N_23510,N_23128,N_23281);
xor U23511 (N_23511,N_23235,N_23338);
xor U23512 (N_23512,N_23144,N_23359);
nand U23513 (N_23513,N_23222,N_23376);
xor U23514 (N_23514,N_23191,N_23228);
nor U23515 (N_23515,N_23136,N_23309);
and U23516 (N_23516,N_23142,N_23137);
nor U23517 (N_23517,N_23113,N_23375);
nor U23518 (N_23518,N_23324,N_23121);
nor U23519 (N_23519,N_23374,N_23348);
xor U23520 (N_23520,N_23203,N_23156);
and U23521 (N_23521,N_23165,N_23214);
xor U23522 (N_23522,N_23131,N_23385);
or U23523 (N_23523,N_23347,N_23223);
nand U23524 (N_23524,N_23391,N_23174);
or U23525 (N_23525,N_23233,N_23129);
or U23526 (N_23526,N_23168,N_23275);
xnor U23527 (N_23527,N_23362,N_23106);
or U23528 (N_23528,N_23193,N_23308);
or U23529 (N_23529,N_23261,N_23102);
nor U23530 (N_23530,N_23173,N_23155);
nor U23531 (N_23531,N_23139,N_23397);
nor U23532 (N_23532,N_23190,N_23268);
nor U23533 (N_23533,N_23279,N_23125);
nand U23534 (N_23534,N_23302,N_23387);
xor U23535 (N_23535,N_23226,N_23328);
nor U23536 (N_23536,N_23119,N_23380);
and U23537 (N_23537,N_23277,N_23147);
nand U23538 (N_23538,N_23243,N_23204);
nor U23539 (N_23539,N_23215,N_23143);
or U23540 (N_23540,N_23327,N_23187);
and U23541 (N_23541,N_23176,N_23221);
nor U23542 (N_23542,N_23134,N_23313);
or U23543 (N_23543,N_23315,N_23114);
nand U23544 (N_23544,N_23105,N_23240);
and U23545 (N_23545,N_23132,N_23283);
xor U23546 (N_23546,N_23227,N_23301);
nor U23547 (N_23547,N_23323,N_23255);
and U23548 (N_23548,N_23287,N_23399);
nand U23549 (N_23549,N_23224,N_23267);
xnor U23550 (N_23550,N_23126,N_23106);
and U23551 (N_23551,N_23227,N_23394);
nand U23552 (N_23552,N_23210,N_23242);
nand U23553 (N_23553,N_23376,N_23295);
and U23554 (N_23554,N_23342,N_23248);
nand U23555 (N_23555,N_23266,N_23325);
xor U23556 (N_23556,N_23258,N_23248);
and U23557 (N_23557,N_23227,N_23199);
and U23558 (N_23558,N_23140,N_23368);
or U23559 (N_23559,N_23179,N_23292);
and U23560 (N_23560,N_23205,N_23367);
and U23561 (N_23561,N_23151,N_23350);
and U23562 (N_23562,N_23378,N_23198);
or U23563 (N_23563,N_23183,N_23126);
and U23564 (N_23564,N_23253,N_23304);
xor U23565 (N_23565,N_23124,N_23324);
and U23566 (N_23566,N_23368,N_23260);
nor U23567 (N_23567,N_23215,N_23281);
nor U23568 (N_23568,N_23324,N_23295);
nand U23569 (N_23569,N_23297,N_23396);
and U23570 (N_23570,N_23234,N_23263);
nand U23571 (N_23571,N_23146,N_23173);
xnor U23572 (N_23572,N_23221,N_23181);
nand U23573 (N_23573,N_23358,N_23170);
or U23574 (N_23574,N_23381,N_23242);
and U23575 (N_23575,N_23154,N_23205);
nand U23576 (N_23576,N_23387,N_23216);
and U23577 (N_23577,N_23339,N_23139);
xnor U23578 (N_23578,N_23164,N_23241);
xnor U23579 (N_23579,N_23110,N_23190);
or U23580 (N_23580,N_23299,N_23308);
nor U23581 (N_23581,N_23369,N_23146);
xnor U23582 (N_23582,N_23224,N_23377);
or U23583 (N_23583,N_23225,N_23270);
nor U23584 (N_23584,N_23322,N_23342);
xnor U23585 (N_23585,N_23323,N_23341);
and U23586 (N_23586,N_23304,N_23157);
and U23587 (N_23587,N_23194,N_23261);
and U23588 (N_23588,N_23116,N_23276);
and U23589 (N_23589,N_23222,N_23306);
and U23590 (N_23590,N_23113,N_23325);
nor U23591 (N_23591,N_23176,N_23287);
and U23592 (N_23592,N_23380,N_23162);
or U23593 (N_23593,N_23151,N_23148);
xnor U23594 (N_23594,N_23176,N_23128);
and U23595 (N_23595,N_23283,N_23345);
xnor U23596 (N_23596,N_23264,N_23152);
nand U23597 (N_23597,N_23197,N_23109);
or U23598 (N_23598,N_23330,N_23130);
or U23599 (N_23599,N_23245,N_23199);
nor U23600 (N_23600,N_23253,N_23346);
and U23601 (N_23601,N_23312,N_23361);
xnor U23602 (N_23602,N_23310,N_23349);
xnor U23603 (N_23603,N_23121,N_23396);
and U23604 (N_23604,N_23111,N_23374);
and U23605 (N_23605,N_23373,N_23346);
nor U23606 (N_23606,N_23216,N_23219);
nor U23607 (N_23607,N_23357,N_23307);
nor U23608 (N_23608,N_23273,N_23164);
nor U23609 (N_23609,N_23181,N_23264);
nand U23610 (N_23610,N_23256,N_23300);
nor U23611 (N_23611,N_23166,N_23362);
nor U23612 (N_23612,N_23195,N_23288);
xnor U23613 (N_23613,N_23211,N_23142);
nand U23614 (N_23614,N_23341,N_23214);
nand U23615 (N_23615,N_23275,N_23276);
xnor U23616 (N_23616,N_23225,N_23245);
xor U23617 (N_23617,N_23141,N_23176);
nand U23618 (N_23618,N_23193,N_23370);
and U23619 (N_23619,N_23207,N_23184);
xnor U23620 (N_23620,N_23299,N_23321);
nor U23621 (N_23621,N_23123,N_23338);
nor U23622 (N_23622,N_23116,N_23211);
nand U23623 (N_23623,N_23101,N_23356);
nand U23624 (N_23624,N_23274,N_23359);
and U23625 (N_23625,N_23328,N_23191);
xor U23626 (N_23626,N_23214,N_23259);
or U23627 (N_23627,N_23233,N_23108);
xnor U23628 (N_23628,N_23112,N_23119);
nor U23629 (N_23629,N_23370,N_23208);
and U23630 (N_23630,N_23313,N_23255);
nand U23631 (N_23631,N_23171,N_23277);
nand U23632 (N_23632,N_23372,N_23199);
and U23633 (N_23633,N_23243,N_23192);
and U23634 (N_23634,N_23327,N_23131);
nand U23635 (N_23635,N_23151,N_23163);
or U23636 (N_23636,N_23282,N_23132);
and U23637 (N_23637,N_23220,N_23237);
or U23638 (N_23638,N_23267,N_23387);
xnor U23639 (N_23639,N_23252,N_23303);
or U23640 (N_23640,N_23260,N_23322);
nor U23641 (N_23641,N_23122,N_23214);
and U23642 (N_23642,N_23185,N_23382);
nand U23643 (N_23643,N_23265,N_23291);
or U23644 (N_23644,N_23142,N_23135);
or U23645 (N_23645,N_23202,N_23159);
nand U23646 (N_23646,N_23353,N_23372);
or U23647 (N_23647,N_23289,N_23233);
xor U23648 (N_23648,N_23102,N_23310);
and U23649 (N_23649,N_23212,N_23160);
xor U23650 (N_23650,N_23164,N_23238);
or U23651 (N_23651,N_23240,N_23114);
or U23652 (N_23652,N_23132,N_23102);
or U23653 (N_23653,N_23222,N_23110);
xnor U23654 (N_23654,N_23362,N_23207);
nor U23655 (N_23655,N_23320,N_23277);
and U23656 (N_23656,N_23324,N_23399);
nor U23657 (N_23657,N_23261,N_23187);
nor U23658 (N_23658,N_23291,N_23110);
or U23659 (N_23659,N_23134,N_23341);
and U23660 (N_23660,N_23359,N_23282);
xnor U23661 (N_23661,N_23143,N_23210);
and U23662 (N_23662,N_23386,N_23147);
and U23663 (N_23663,N_23232,N_23304);
xor U23664 (N_23664,N_23218,N_23340);
xnor U23665 (N_23665,N_23357,N_23196);
or U23666 (N_23666,N_23225,N_23244);
or U23667 (N_23667,N_23391,N_23319);
nor U23668 (N_23668,N_23163,N_23344);
xor U23669 (N_23669,N_23187,N_23299);
nand U23670 (N_23670,N_23369,N_23144);
and U23671 (N_23671,N_23259,N_23298);
or U23672 (N_23672,N_23302,N_23208);
and U23673 (N_23673,N_23256,N_23374);
nor U23674 (N_23674,N_23113,N_23330);
xnor U23675 (N_23675,N_23233,N_23395);
nor U23676 (N_23676,N_23237,N_23330);
nor U23677 (N_23677,N_23311,N_23115);
nand U23678 (N_23678,N_23395,N_23305);
nor U23679 (N_23679,N_23393,N_23330);
nor U23680 (N_23680,N_23254,N_23126);
nand U23681 (N_23681,N_23124,N_23272);
nand U23682 (N_23682,N_23264,N_23387);
nand U23683 (N_23683,N_23207,N_23130);
nor U23684 (N_23684,N_23355,N_23122);
or U23685 (N_23685,N_23324,N_23211);
and U23686 (N_23686,N_23299,N_23174);
nand U23687 (N_23687,N_23241,N_23334);
and U23688 (N_23688,N_23341,N_23374);
and U23689 (N_23689,N_23286,N_23165);
and U23690 (N_23690,N_23256,N_23273);
nand U23691 (N_23691,N_23196,N_23296);
xor U23692 (N_23692,N_23206,N_23202);
or U23693 (N_23693,N_23342,N_23301);
and U23694 (N_23694,N_23254,N_23200);
nand U23695 (N_23695,N_23246,N_23399);
or U23696 (N_23696,N_23172,N_23290);
and U23697 (N_23697,N_23157,N_23195);
xor U23698 (N_23698,N_23224,N_23135);
nor U23699 (N_23699,N_23243,N_23157);
nor U23700 (N_23700,N_23517,N_23542);
nor U23701 (N_23701,N_23669,N_23643);
nor U23702 (N_23702,N_23597,N_23653);
xnor U23703 (N_23703,N_23459,N_23418);
xor U23704 (N_23704,N_23479,N_23514);
and U23705 (N_23705,N_23478,N_23591);
nand U23706 (N_23706,N_23681,N_23468);
nand U23707 (N_23707,N_23678,N_23499);
xor U23708 (N_23708,N_23620,N_23606);
and U23709 (N_23709,N_23648,N_23655);
xor U23710 (N_23710,N_23533,N_23439);
or U23711 (N_23711,N_23524,N_23460);
nor U23712 (N_23712,N_23414,N_23471);
or U23713 (N_23713,N_23550,N_23570);
or U23714 (N_23714,N_23527,N_23448);
and U23715 (N_23715,N_23497,N_23537);
nand U23716 (N_23716,N_23465,N_23472);
and U23717 (N_23717,N_23580,N_23635);
nor U23718 (N_23718,N_23561,N_23661);
or U23719 (N_23719,N_23658,N_23423);
nand U23720 (N_23720,N_23672,N_23470);
nand U23721 (N_23721,N_23541,N_23564);
and U23722 (N_23722,N_23500,N_23554);
nand U23723 (N_23723,N_23494,N_23599);
xor U23724 (N_23724,N_23419,N_23657);
or U23725 (N_23725,N_23464,N_23660);
or U23726 (N_23726,N_23697,N_23403);
xnor U23727 (N_23727,N_23602,N_23536);
xnor U23728 (N_23728,N_23574,N_23611);
xnor U23729 (N_23729,N_23692,N_23633);
nor U23730 (N_23730,N_23557,N_23639);
nand U23731 (N_23731,N_23670,N_23626);
and U23732 (N_23732,N_23452,N_23477);
nand U23733 (N_23733,N_23650,N_23445);
or U23734 (N_23734,N_23462,N_23590);
or U23735 (N_23735,N_23528,N_23690);
nand U23736 (N_23736,N_23566,N_23637);
or U23737 (N_23737,N_23677,N_23446);
nor U23738 (N_23738,N_23642,N_23401);
xnor U23739 (N_23739,N_23532,N_23507);
nor U23740 (N_23740,N_23604,N_23600);
or U23741 (N_23741,N_23505,N_23513);
or U23742 (N_23742,N_23493,N_23520);
xor U23743 (N_23743,N_23573,N_23529);
nand U23744 (N_23744,N_23640,N_23576);
nand U23745 (N_23745,N_23495,N_23461);
nor U23746 (N_23746,N_23556,N_23673);
nor U23747 (N_23747,N_23416,N_23417);
xor U23748 (N_23748,N_23649,N_23409);
nand U23749 (N_23749,N_23593,N_23422);
xnor U23750 (N_23750,N_23685,N_23453);
nor U23751 (N_23751,N_23689,N_23518);
xnor U23752 (N_23752,N_23562,N_23680);
xor U23753 (N_23753,N_23463,N_23488);
or U23754 (N_23754,N_23686,N_23696);
xnor U23755 (N_23755,N_23615,N_23695);
nand U23756 (N_23756,N_23492,N_23607);
and U23757 (N_23757,N_23683,N_23665);
nand U23758 (N_23758,N_23530,N_23592);
xnor U23759 (N_23759,N_23585,N_23552);
or U23760 (N_23760,N_23441,N_23630);
nor U23761 (N_23761,N_23456,N_23415);
or U23762 (N_23762,N_23578,N_23628);
nand U23763 (N_23763,N_23581,N_23589);
and U23764 (N_23764,N_23598,N_23410);
nand U23765 (N_23765,N_23601,N_23671);
nor U23766 (N_23766,N_23534,N_23612);
and U23767 (N_23767,N_23484,N_23688);
nand U23768 (N_23768,N_23525,N_23654);
xnor U23769 (N_23769,N_23547,N_23631);
and U23770 (N_23770,N_23496,N_23447);
nor U23771 (N_23771,N_23610,N_23627);
and U23772 (N_23772,N_23485,N_23539);
nor U23773 (N_23773,N_23467,N_23618);
nand U23774 (N_23774,N_23603,N_23641);
or U23775 (N_23775,N_23645,N_23408);
nand U23776 (N_23776,N_23569,N_23502);
or U23777 (N_23777,N_23511,N_23621);
or U23778 (N_23778,N_23568,N_23651);
xor U23779 (N_23779,N_23444,N_23668);
and U23780 (N_23780,N_23616,N_23503);
nor U23781 (N_23781,N_23634,N_23667);
nand U23782 (N_23782,N_23427,N_23519);
and U23783 (N_23783,N_23664,N_23451);
nand U23784 (N_23784,N_23424,N_23544);
xnor U23785 (N_23785,N_23659,N_23475);
nor U23786 (N_23786,N_23512,N_23636);
or U23787 (N_23787,N_23455,N_23624);
and U23788 (N_23788,N_23483,N_23553);
and U23789 (N_23789,N_23567,N_23571);
and U23790 (N_23790,N_23605,N_23619);
nand U23791 (N_23791,N_23489,N_23656);
xor U23792 (N_23792,N_23438,N_23443);
and U23793 (N_23793,N_23623,N_23476);
and U23794 (N_23794,N_23594,N_23579);
xor U23795 (N_23795,N_23449,N_23609);
nor U23796 (N_23796,N_23596,N_23587);
xor U23797 (N_23797,N_23560,N_23405);
or U23798 (N_23798,N_23515,N_23436);
and U23799 (N_23799,N_23586,N_23454);
nor U23800 (N_23800,N_23676,N_23508);
xnor U23801 (N_23801,N_23662,N_23501);
and U23802 (N_23802,N_23434,N_23558);
or U23803 (N_23803,N_23543,N_23450);
nand U23804 (N_23804,N_23506,N_23487);
or U23805 (N_23805,N_23458,N_23442);
nand U23806 (N_23806,N_23694,N_23563);
nor U23807 (N_23807,N_23420,N_23663);
or U23808 (N_23808,N_23666,N_23491);
nor U23809 (N_23809,N_23684,N_23437);
xnor U23810 (N_23810,N_23691,N_23582);
nor U23811 (N_23811,N_23429,N_23522);
or U23812 (N_23812,N_23466,N_23435);
nand U23813 (N_23813,N_23555,N_23486);
nor U23814 (N_23814,N_23440,N_23402);
nand U23815 (N_23815,N_23413,N_23652);
or U23816 (N_23816,N_23433,N_23632);
xnor U23817 (N_23817,N_23644,N_23546);
xnor U23818 (N_23818,N_23548,N_23469);
xnor U23819 (N_23819,N_23583,N_23474);
xor U23820 (N_23820,N_23457,N_23411);
or U23821 (N_23821,N_23584,N_23608);
or U23822 (N_23822,N_23516,N_23535);
nand U23823 (N_23823,N_23647,N_23498);
nand U23824 (N_23824,N_23577,N_23481);
nor U23825 (N_23825,N_23421,N_23509);
nand U23826 (N_23826,N_23698,N_23622);
and U23827 (N_23827,N_23595,N_23426);
nor U23828 (N_23828,N_23565,N_23490);
nor U23829 (N_23829,N_23693,N_23613);
or U23830 (N_23830,N_23406,N_23480);
and U23831 (N_23831,N_23521,N_23523);
nand U23832 (N_23832,N_23545,N_23614);
or U23833 (N_23833,N_23531,N_23588);
xnor U23834 (N_23834,N_23646,N_23538);
and U23835 (N_23835,N_23431,N_23404);
nand U23836 (N_23836,N_23625,N_23510);
xnor U23837 (N_23837,N_23412,N_23504);
or U23838 (N_23838,N_23428,N_23407);
and U23839 (N_23839,N_23617,N_23629);
nand U23840 (N_23840,N_23682,N_23674);
and U23841 (N_23841,N_23551,N_23540);
and U23842 (N_23842,N_23679,N_23675);
or U23843 (N_23843,N_23432,N_23699);
nor U23844 (N_23844,N_23473,N_23572);
and U23845 (N_23845,N_23549,N_23400);
nand U23846 (N_23846,N_23575,N_23482);
xor U23847 (N_23847,N_23687,N_23430);
nor U23848 (N_23848,N_23425,N_23559);
or U23849 (N_23849,N_23526,N_23638);
nor U23850 (N_23850,N_23464,N_23456);
or U23851 (N_23851,N_23554,N_23454);
nand U23852 (N_23852,N_23535,N_23453);
xnor U23853 (N_23853,N_23437,N_23687);
xnor U23854 (N_23854,N_23592,N_23487);
and U23855 (N_23855,N_23447,N_23412);
xnor U23856 (N_23856,N_23406,N_23657);
or U23857 (N_23857,N_23603,N_23525);
nor U23858 (N_23858,N_23546,N_23508);
or U23859 (N_23859,N_23475,N_23584);
nand U23860 (N_23860,N_23579,N_23539);
xnor U23861 (N_23861,N_23452,N_23486);
nand U23862 (N_23862,N_23661,N_23427);
xor U23863 (N_23863,N_23506,N_23533);
or U23864 (N_23864,N_23613,N_23639);
xor U23865 (N_23865,N_23593,N_23581);
xnor U23866 (N_23866,N_23687,N_23677);
and U23867 (N_23867,N_23688,N_23668);
and U23868 (N_23868,N_23488,N_23430);
xor U23869 (N_23869,N_23531,N_23695);
nor U23870 (N_23870,N_23545,N_23653);
nand U23871 (N_23871,N_23635,N_23522);
xor U23872 (N_23872,N_23649,N_23690);
and U23873 (N_23873,N_23661,N_23567);
nand U23874 (N_23874,N_23452,N_23690);
xor U23875 (N_23875,N_23636,N_23685);
nor U23876 (N_23876,N_23491,N_23410);
nand U23877 (N_23877,N_23644,N_23528);
or U23878 (N_23878,N_23582,N_23579);
or U23879 (N_23879,N_23638,N_23544);
and U23880 (N_23880,N_23669,N_23508);
or U23881 (N_23881,N_23648,N_23643);
xor U23882 (N_23882,N_23584,N_23620);
xor U23883 (N_23883,N_23638,N_23455);
nor U23884 (N_23884,N_23459,N_23496);
xor U23885 (N_23885,N_23693,N_23520);
xor U23886 (N_23886,N_23602,N_23490);
nand U23887 (N_23887,N_23478,N_23635);
nand U23888 (N_23888,N_23546,N_23600);
nand U23889 (N_23889,N_23698,N_23596);
xor U23890 (N_23890,N_23562,N_23534);
and U23891 (N_23891,N_23695,N_23624);
xnor U23892 (N_23892,N_23551,N_23626);
or U23893 (N_23893,N_23690,N_23509);
nand U23894 (N_23894,N_23670,N_23552);
or U23895 (N_23895,N_23501,N_23464);
or U23896 (N_23896,N_23591,N_23605);
nand U23897 (N_23897,N_23642,N_23489);
or U23898 (N_23898,N_23618,N_23671);
xnor U23899 (N_23899,N_23500,N_23646);
and U23900 (N_23900,N_23556,N_23662);
nor U23901 (N_23901,N_23672,N_23611);
nand U23902 (N_23902,N_23594,N_23492);
xnor U23903 (N_23903,N_23569,N_23521);
or U23904 (N_23904,N_23486,N_23519);
nand U23905 (N_23905,N_23571,N_23689);
or U23906 (N_23906,N_23499,N_23501);
xor U23907 (N_23907,N_23653,N_23667);
nand U23908 (N_23908,N_23511,N_23561);
nor U23909 (N_23909,N_23501,N_23659);
or U23910 (N_23910,N_23400,N_23528);
nand U23911 (N_23911,N_23536,N_23628);
and U23912 (N_23912,N_23560,N_23412);
and U23913 (N_23913,N_23625,N_23574);
or U23914 (N_23914,N_23695,N_23677);
xor U23915 (N_23915,N_23420,N_23482);
nand U23916 (N_23916,N_23547,N_23643);
xnor U23917 (N_23917,N_23441,N_23623);
xnor U23918 (N_23918,N_23450,N_23552);
xnor U23919 (N_23919,N_23686,N_23635);
or U23920 (N_23920,N_23606,N_23488);
and U23921 (N_23921,N_23467,N_23464);
or U23922 (N_23922,N_23432,N_23591);
and U23923 (N_23923,N_23612,N_23567);
nor U23924 (N_23924,N_23649,N_23534);
nor U23925 (N_23925,N_23525,N_23630);
xnor U23926 (N_23926,N_23641,N_23480);
xnor U23927 (N_23927,N_23443,N_23612);
and U23928 (N_23928,N_23639,N_23449);
nand U23929 (N_23929,N_23500,N_23447);
or U23930 (N_23930,N_23699,N_23513);
nor U23931 (N_23931,N_23516,N_23451);
or U23932 (N_23932,N_23487,N_23456);
nand U23933 (N_23933,N_23665,N_23668);
and U23934 (N_23934,N_23571,N_23630);
xnor U23935 (N_23935,N_23630,N_23508);
nand U23936 (N_23936,N_23671,N_23475);
and U23937 (N_23937,N_23605,N_23594);
and U23938 (N_23938,N_23632,N_23657);
and U23939 (N_23939,N_23622,N_23694);
nand U23940 (N_23940,N_23602,N_23589);
xnor U23941 (N_23941,N_23694,N_23400);
nand U23942 (N_23942,N_23597,N_23430);
nor U23943 (N_23943,N_23697,N_23533);
nor U23944 (N_23944,N_23665,N_23491);
and U23945 (N_23945,N_23544,N_23445);
and U23946 (N_23946,N_23634,N_23696);
and U23947 (N_23947,N_23553,N_23467);
or U23948 (N_23948,N_23423,N_23676);
xnor U23949 (N_23949,N_23458,N_23660);
and U23950 (N_23950,N_23680,N_23495);
and U23951 (N_23951,N_23695,N_23405);
nor U23952 (N_23952,N_23624,N_23589);
nand U23953 (N_23953,N_23693,N_23651);
nor U23954 (N_23954,N_23401,N_23658);
nor U23955 (N_23955,N_23481,N_23600);
nor U23956 (N_23956,N_23602,N_23624);
xor U23957 (N_23957,N_23659,N_23538);
or U23958 (N_23958,N_23566,N_23622);
nand U23959 (N_23959,N_23401,N_23499);
or U23960 (N_23960,N_23577,N_23601);
xnor U23961 (N_23961,N_23508,N_23469);
nor U23962 (N_23962,N_23553,N_23666);
xor U23963 (N_23963,N_23564,N_23694);
nor U23964 (N_23964,N_23682,N_23510);
nor U23965 (N_23965,N_23613,N_23566);
nand U23966 (N_23966,N_23498,N_23560);
xor U23967 (N_23967,N_23633,N_23694);
nor U23968 (N_23968,N_23602,N_23414);
or U23969 (N_23969,N_23457,N_23616);
and U23970 (N_23970,N_23675,N_23590);
and U23971 (N_23971,N_23576,N_23423);
xor U23972 (N_23972,N_23645,N_23685);
xor U23973 (N_23973,N_23538,N_23403);
nor U23974 (N_23974,N_23539,N_23493);
and U23975 (N_23975,N_23507,N_23550);
xor U23976 (N_23976,N_23674,N_23631);
xnor U23977 (N_23977,N_23430,N_23541);
or U23978 (N_23978,N_23483,N_23622);
and U23979 (N_23979,N_23689,N_23513);
and U23980 (N_23980,N_23508,N_23503);
nor U23981 (N_23981,N_23626,N_23517);
nand U23982 (N_23982,N_23542,N_23411);
nand U23983 (N_23983,N_23546,N_23609);
nor U23984 (N_23984,N_23469,N_23448);
nand U23985 (N_23985,N_23568,N_23509);
and U23986 (N_23986,N_23412,N_23431);
and U23987 (N_23987,N_23659,N_23468);
nand U23988 (N_23988,N_23457,N_23453);
and U23989 (N_23989,N_23676,N_23574);
or U23990 (N_23990,N_23583,N_23529);
nand U23991 (N_23991,N_23571,N_23626);
nor U23992 (N_23992,N_23411,N_23681);
and U23993 (N_23993,N_23556,N_23663);
and U23994 (N_23994,N_23487,N_23547);
nor U23995 (N_23995,N_23456,N_23461);
xnor U23996 (N_23996,N_23667,N_23561);
nor U23997 (N_23997,N_23680,N_23669);
nand U23998 (N_23998,N_23585,N_23413);
nor U23999 (N_23999,N_23445,N_23415);
xor U24000 (N_24000,N_23740,N_23803);
or U24001 (N_24001,N_23983,N_23701);
xnor U24002 (N_24002,N_23734,N_23984);
or U24003 (N_24003,N_23974,N_23884);
or U24004 (N_24004,N_23778,N_23970);
nand U24005 (N_24005,N_23855,N_23864);
and U24006 (N_24006,N_23877,N_23757);
or U24007 (N_24007,N_23949,N_23870);
xor U24008 (N_24008,N_23773,N_23898);
xnor U24009 (N_24009,N_23765,N_23736);
or U24010 (N_24010,N_23790,N_23913);
xnor U24011 (N_24011,N_23885,N_23986);
and U24012 (N_24012,N_23801,N_23707);
nand U24013 (N_24013,N_23872,N_23869);
or U24014 (N_24014,N_23795,N_23860);
nor U24015 (N_24015,N_23907,N_23867);
xnor U24016 (N_24016,N_23840,N_23964);
xor U24017 (N_24017,N_23873,N_23819);
or U24018 (N_24018,N_23771,N_23807);
nand U24019 (N_24019,N_23737,N_23813);
and U24020 (N_24020,N_23962,N_23838);
xor U24021 (N_24021,N_23766,N_23991);
and U24022 (N_24022,N_23826,N_23925);
xnor U24023 (N_24023,N_23879,N_23805);
or U24024 (N_24024,N_23893,N_23876);
nand U24025 (N_24025,N_23748,N_23997);
nor U24026 (N_24026,N_23727,N_23868);
and U24027 (N_24027,N_23921,N_23976);
nand U24028 (N_24028,N_23918,N_23897);
and U24029 (N_24029,N_23811,N_23782);
and U24030 (N_24030,N_23797,N_23927);
nor U24031 (N_24031,N_23961,N_23709);
nor U24032 (N_24032,N_23906,N_23895);
xor U24033 (N_24033,N_23746,N_23954);
nor U24034 (N_24034,N_23837,N_23752);
and U24035 (N_24035,N_23888,N_23963);
nor U24036 (N_24036,N_23761,N_23995);
nor U24037 (N_24037,N_23793,N_23874);
nand U24038 (N_24038,N_23772,N_23754);
nor U24039 (N_24039,N_23985,N_23948);
xor U24040 (N_24040,N_23785,N_23878);
and U24041 (N_24041,N_23816,N_23828);
or U24042 (N_24042,N_23940,N_23742);
nor U24043 (N_24043,N_23739,N_23971);
xnor U24044 (N_24044,N_23978,N_23892);
xnor U24045 (N_24045,N_23977,N_23990);
xor U24046 (N_24046,N_23706,N_23718);
nand U24047 (N_24047,N_23779,N_23777);
nand U24048 (N_24048,N_23967,N_23929);
nor U24049 (N_24049,N_23836,N_23800);
nor U24050 (N_24050,N_23731,N_23999);
xnor U24051 (N_24051,N_23809,N_23751);
or U24052 (N_24052,N_23883,N_23862);
or U24053 (N_24053,N_23786,N_23965);
nand U24054 (N_24054,N_23848,N_23743);
nor U24055 (N_24055,N_23762,N_23835);
or U24056 (N_24056,N_23760,N_23996);
and U24057 (N_24057,N_23723,N_23890);
nor U24058 (N_24058,N_23945,N_23871);
and U24059 (N_24059,N_23851,N_23825);
or U24060 (N_24060,N_23796,N_23924);
nor U24061 (N_24061,N_23946,N_23902);
nor U24062 (N_24062,N_23829,N_23725);
nor U24063 (N_24063,N_23810,N_23747);
nand U24064 (N_24064,N_23903,N_23756);
xor U24065 (N_24065,N_23802,N_23863);
and U24066 (N_24066,N_23833,N_23972);
xor U24067 (N_24067,N_23856,N_23959);
xnor U24068 (N_24068,N_23764,N_23899);
nand U24069 (N_24069,N_23719,N_23843);
and U24070 (N_24070,N_23915,N_23726);
nor U24071 (N_24071,N_23787,N_23794);
and U24072 (N_24072,N_23817,N_23744);
xnor U24073 (N_24073,N_23753,N_23944);
xnor U24074 (N_24074,N_23937,N_23889);
nand U24075 (N_24075,N_23712,N_23947);
nor U24076 (N_24076,N_23926,N_23939);
nor U24077 (N_24077,N_23784,N_23824);
nor U24078 (N_24078,N_23763,N_23839);
xor U24079 (N_24079,N_23846,N_23717);
or U24080 (N_24080,N_23881,N_23776);
nor U24081 (N_24081,N_23919,N_23716);
and U24082 (N_24082,N_23806,N_23820);
or U24083 (N_24083,N_23953,N_23988);
nand U24084 (N_24084,N_23982,N_23951);
or U24085 (N_24085,N_23956,N_23732);
nor U24086 (N_24086,N_23781,N_23722);
or U24087 (N_24087,N_23710,N_23729);
nand U24088 (N_24088,N_23823,N_23830);
or U24089 (N_24089,N_23981,N_23711);
and U24090 (N_24090,N_23832,N_23850);
nand U24091 (N_24091,N_23720,N_23882);
nand U24092 (N_24092,N_23822,N_23875);
nand U24093 (N_24093,N_23791,N_23755);
or U24094 (N_24094,N_23834,N_23941);
and U24095 (N_24095,N_23886,N_23758);
nor U24096 (N_24096,N_23935,N_23702);
nand U24097 (N_24097,N_23866,N_23842);
xor U24098 (N_24098,N_23943,N_23909);
xor U24099 (N_24099,N_23827,N_23708);
nor U24100 (N_24100,N_23960,N_23774);
nand U24101 (N_24101,N_23955,N_23923);
or U24102 (N_24102,N_23932,N_23704);
or U24103 (N_24103,N_23942,N_23914);
and U24104 (N_24104,N_23814,N_23703);
and U24105 (N_24105,N_23911,N_23894);
or U24106 (N_24106,N_23821,N_23713);
xor U24107 (N_24107,N_23730,N_23969);
or U24108 (N_24108,N_23783,N_23880);
and U24109 (N_24109,N_23841,N_23975);
xnor U24110 (N_24110,N_23788,N_23896);
and U24111 (N_24111,N_23768,N_23973);
or U24112 (N_24112,N_23859,N_23847);
xnor U24113 (N_24113,N_23815,N_23992);
and U24114 (N_24114,N_23950,N_23745);
nor U24115 (N_24115,N_23966,N_23714);
and U24116 (N_24116,N_23910,N_23922);
and U24117 (N_24117,N_23901,N_23994);
or U24118 (N_24118,N_23861,N_23987);
and U24119 (N_24119,N_23705,N_23968);
nand U24120 (N_24120,N_23769,N_23957);
nor U24121 (N_24121,N_23887,N_23952);
xnor U24122 (N_24122,N_23715,N_23905);
and U24123 (N_24123,N_23930,N_23993);
nor U24124 (N_24124,N_23989,N_23733);
or U24125 (N_24125,N_23917,N_23789);
or U24126 (N_24126,N_23928,N_23780);
or U24127 (N_24127,N_23858,N_23759);
nor U24128 (N_24128,N_23721,N_23738);
nor U24129 (N_24129,N_23775,N_23958);
xnor U24130 (N_24130,N_23857,N_23908);
and U24131 (N_24131,N_23916,N_23792);
and U24132 (N_24132,N_23931,N_23808);
nor U24133 (N_24133,N_23891,N_23920);
or U24134 (N_24134,N_23741,N_23998);
and U24135 (N_24135,N_23770,N_23804);
nand U24136 (N_24136,N_23865,N_23934);
xor U24137 (N_24137,N_23844,N_23980);
or U24138 (N_24138,N_23933,N_23724);
nand U24139 (N_24139,N_23936,N_23767);
and U24140 (N_24140,N_23900,N_23904);
nor U24141 (N_24141,N_23799,N_23818);
or U24142 (N_24142,N_23728,N_23912);
nor U24143 (N_24143,N_23979,N_23852);
nor U24144 (N_24144,N_23849,N_23845);
or U24145 (N_24145,N_23812,N_23853);
and U24146 (N_24146,N_23938,N_23735);
xor U24147 (N_24147,N_23854,N_23750);
and U24148 (N_24148,N_23700,N_23831);
and U24149 (N_24149,N_23749,N_23798);
xor U24150 (N_24150,N_23858,N_23937);
nand U24151 (N_24151,N_23832,N_23981);
nand U24152 (N_24152,N_23874,N_23937);
nor U24153 (N_24153,N_23725,N_23937);
nor U24154 (N_24154,N_23797,N_23790);
xor U24155 (N_24155,N_23803,N_23841);
nand U24156 (N_24156,N_23933,N_23767);
or U24157 (N_24157,N_23733,N_23980);
or U24158 (N_24158,N_23878,N_23752);
xor U24159 (N_24159,N_23794,N_23937);
or U24160 (N_24160,N_23710,N_23796);
nor U24161 (N_24161,N_23993,N_23785);
and U24162 (N_24162,N_23978,N_23972);
and U24163 (N_24163,N_23853,N_23891);
nand U24164 (N_24164,N_23747,N_23868);
or U24165 (N_24165,N_23776,N_23942);
nand U24166 (N_24166,N_23860,N_23977);
nor U24167 (N_24167,N_23897,N_23915);
or U24168 (N_24168,N_23848,N_23956);
nor U24169 (N_24169,N_23953,N_23976);
nor U24170 (N_24170,N_23772,N_23846);
and U24171 (N_24171,N_23966,N_23760);
nand U24172 (N_24172,N_23745,N_23995);
nand U24173 (N_24173,N_23835,N_23827);
xor U24174 (N_24174,N_23929,N_23820);
or U24175 (N_24175,N_23888,N_23951);
nor U24176 (N_24176,N_23896,N_23974);
xnor U24177 (N_24177,N_23838,N_23789);
nand U24178 (N_24178,N_23909,N_23880);
or U24179 (N_24179,N_23786,N_23962);
nor U24180 (N_24180,N_23885,N_23893);
nor U24181 (N_24181,N_23740,N_23973);
nand U24182 (N_24182,N_23856,N_23963);
and U24183 (N_24183,N_23777,N_23737);
nor U24184 (N_24184,N_23896,N_23813);
nor U24185 (N_24185,N_23830,N_23775);
or U24186 (N_24186,N_23832,N_23742);
nand U24187 (N_24187,N_23912,N_23704);
nor U24188 (N_24188,N_23954,N_23802);
or U24189 (N_24189,N_23871,N_23756);
and U24190 (N_24190,N_23884,N_23849);
nand U24191 (N_24191,N_23899,N_23811);
nand U24192 (N_24192,N_23922,N_23768);
and U24193 (N_24193,N_23946,N_23887);
and U24194 (N_24194,N_23856,N_23989);
nand U24195 (N_24195,N_23808,N_23748);
and U24196 (N_24196,N_23982,N_23946);
nand U24197 (N_24197,N_23963,N_23997);
and U24198 (N_24198,N_23982,N_23835);
or U24199 (N_24199,N_23764,N_23731);
nand U24200 (N_24200,N_23801,N_23962);
nand U24201 (N_24201,N_23778,N_23724);
nor U24202 (N_24202,N_23757,N_23859);
nor U24203 (N_24203,N_23811,N_23732);
and U24204 (N_24204,N_23909,N_23885);
xor U24205 (N_24205,N_23884,N_23778);
nand U24206 (N_24206,N_23849,N_23906);
xnor U24207 (N_24207,N_23795,N_23830);
nand U24208 (N_24208,N_23713,N_23903);
or U24209 (N_24209,N_23866,N_23825);
xor U24210 (N_24210,N_23777,N_23822);
or U24211 (N_24211,N_23719,N_23961);
nand U24212 (N_24212,N_23806,N_23942);
xnor U24213 (N_24213,N_23949,N_23792);
and U24214 (N_24214,N_23857,N_23707);
nor U24215 (N_24215,N_23890,N_23754);
and U24216 (N_24216,N_23725,N_23766);
nor U24217 (N_24217,N_23703,N_23878);
xor U24218 (N_24218,N_23846,N_23751);
or U24219 (N_24219,N_23793,N_23996);
nor U24220 (N_24220,N_23999,N_23893);
or U24221 (N_24221,N_23707,N_23824);
and U24222 (N_24222,N_23782,N_23930);
nor U24223 (N_24223,N_23726,N_23925);
or U24224 (N_24224,N_23977,N_23981);
nor U24225 (N_24225,N_23951,N_23953);
xor U24226 (N_24226,N_23709,N_23703);
xor U24227 (N_24227,N_23959,N_23770);
and U24228 (N_24228,N_23700,N_23994);
and U24229 (N_24229,N_23942,N_23832);
or U24230 (N_24230,N_23887,N_23758);
or U24231 (N_24231,N_23971,N_23877);
nand U24232 (N_24232,N_23709,N_23701);
and U24233 (N_24233,N_23738,N_23945);
nor U24234 (N_24234,N_23716,N_23809);
and U24235 (N_24235,N_23991,N_23746);
xor U24236 (N_24236,N_23893,N_23712);
nand U24237 (N_24237,N_23760,N_23794);
or U24238 (N_24238,N_23923,N_23815);
xnor U24239 (N_24239,N_23915,N_23753);
or U24240 (N_24240,N_23927,N_23881);
and U24241 (N_24241,N_23879,N_23900);
nor U24242 (N_24242,N_23853,N_23925);
and U24243 (N_24243,N_23908,N_23941);
nor U24244 (N_24244,N_23830,N_23881);
or U24245 (N_24245,N_23758,N_23778);
nand U24246 (N_24246,N_23838,N_23713);
or U24247 (N_24247,N_23847,N_23716);
or U24248 (N_24248,N_23743,N_23709);
nor U24249 (N_24249,N_23924,N_23740);
nor U24250 (N_24250,N_23895,N_23759);
xor U24251 (N_24251,N_23871,N_23720);
nand U24252 (N_24252,N_23742,N_23909);
nand U24253 (N_24253,N_23801,N_23888);
or U24254 (N_24254,N_23910,N_23736);
and U24255 (N_24255,N_23948,N_23954);
xnor U24256 (N_24256,N_23988,N_23838);
and U24257 (N_24257,N_23802,N_23902);
nor U24258 (N_24258,N_23907,N_23914);
nand U24259 (N_24259,N_23743,N_23726);
or U24260 (N_24260,N_23928,N_23750);
or U24261 (N_24261,N_23965,N_23885);
nand U24262 (N_24262,N_23915,N_23846);
and U24263 (N_24263,N_23831,N_23833);
nand U24264 (N_24264,N_23907,N_23729);
or U24265 (N_24265,N_23932,N_23789);
xnor U24266 (N_24266,N_23963,N_23829);
or U24267 (N_24267,N_23795,N_23907);
xnor U24268 (N_24268,N_23960,N_23741);
nor U24269 (N_24269,N_23800,N_23765);
or U24270 (N_24270,N_23808,N_23818);
nand U24271 (N_24271,N_23980,N_23707);
and U24272 (N_24272,N_23703,N_23788);
and U24273 (N_24273,N_23810,N_23843);
nor U24274 (N_24274,N_23825,N_23975);
or U24275 (N_24275,N_23928,N_23754);
xnor U24276 (N_24276,N_23906,N_23939);
or U24277 (N_24277,N_23747,N_23732);
xor U24278 (N_24278,N_23920,N_23860);
xnor U24279 (N_24279,N_23966,N_23794);
or U24280 (N_24280,N_23930,N_23938);
nor U24281 (N_24281,N_23873,N_23731);
nand U24282 (N_24282,N_23991,N_23931);
xnor U24283 (N_24283,N_23716,N_23788);
nand U24284 (N_24284,N_23973,N_23825);
and U24285 (N_24285,N_23720,N_23908);
xor U24286 (N_24286,N_23853,N_23849);
nand U24287 (N_24287,N_23944,N_23921);
nand U24288 (N_24288,N_23896,N_23749);
xnor U24289 (N_24289,N_23704,N_23991);
nand U24290 (N_24290,N_23888,N_23784);
or U24291 (N_24291,N_23930,N_23956);
and U24292 (N_24292,N_23760,N_23870);
xor U24293 (N_24293,N_23788,N_23874);
nor U24294 (N_24294,N_23893,N_23998);
and U24295 (N_24295,N_23915,N_23757);
nand U24296 (N_24296,N_23700,N_23789);
xnor U24297 (N_24297,N_23833,N_23803);
or U24298 (N_24298,N_23799,N_23786);
or U24299 (N_24299,N_23769,N_23798);
nand U24300 (N_24300,N_24135,N_24107);
nor U24301 (N_24301,N_24152,N_24227);
nand U24302 (N_24302,N_24178,N_24240);
nor U24303 (N_24303,N_24159,N_24224);
or U24304 (N_24304,N_24042,N_24198);
or U24305 (N_24305,N_24050,N_24272);
and U24306 (N_24306,N_24153,N_24235);
xnor U24307 (N_24307,N_24214,N_24186);
nor U24308 (N_24308,N_24265,N_24118);
nand U24309 (N_24309,N_24239,N_24248);
nor U24310 (N_24310,N_24018,N_24256);
or U24311 (N_24311,N_24076,N_24200);
and U24312 (N_24312,N_24146,N_24169);
nor U24313 (N_24313,N_24253,N_24195);
and U24314 (N_24314,N_24019,N_24001);
nor U24315 (N_24315,N_24049,N_24279);
nor U24316 (N_24316,N_24197,N_24267);
xor U24317 (N_24317,N_24184,N_24236);
and U24318 (N_24318,N_24137,N_24298);
nand U24319 (N_24319,N_24207,N_24048);
or U24320 (N_24320,N_24142,N_24055);
or U24321 (N_24321,N_24145,N_24120);
nor U24322 (N_24322,N_24000,N_24278);
or U24323 (N_24323,N_24147,N_24128);
xnor U24324 (N_24324,N_24160,N_24182);
nand U24325 (N_24325,N_24225,N_24201);
xnor U24326 (N_24326,N_24136,N_24038);
and U24327 (N_24327,N_24290,N_24172);
and U24328 (N_24328,N_24250,N_24068);
and U24329 (N_24329,N_24101,N_24177);
and U24330 (N_24330,N_24045,N_24295);
and U24331 (N_24331,N_24229,N_24228);
nor U24332 (N_24332,N_24154,N_24241);
nor U24333 (N_24333,N_24130,N_24085);
nor U24334 (N_24334,N_24148,N_24098);
xor U24335 (N_24335,N_24123,N_24007);
xnor U24336 (N_24336,N_24066,N_24131);
nand U24337 (N_24337,N_24299,N_24113);
nor U24338 (N_24338,N_24210,N_24183);
nor U24339 (N_24339,N_24175,N_24035);
xnor U24340 (N_24340,N_24108,N_24078);
nand U24341 (N_24341,N_24208,N_24282);
nand U24342 (N_24342,N_24296,N_24079);
nor U24343 (N_24343,N_24083,N_24029);
nor U24344 (N_24344,N_24074,N_24161);
xor U24345 (N_24345,N_24090,N_24285);
or U24346 (N_24346,N_24259,N_24163);
nor U24347 (N_24347,N_24185,N_24046);
nand U24348 (N_24348,N_24116,N_24139);
and U24349 (N_24349,N_24133,N_24180);
nand U24350 (N_24350,N_24275,N_24288);
or U24351 (N_24351,N_24039,N_24286);
or U24352 (N_24352,N_24077,N_24155);
or U24353 (N_24353,N_24121,N_24181);
xnor U24354 (N_24354,N_24191,N_24268);
or U24355 (N_24355,N_24105,N_24099);
and U24356 (N_24356,N_24162,N_24047);
xor U24357 (N_24357,N_24258,N_24244);
xor U24358 (N_24358,N_24003,N_24106);
nor U24359 (N_24359,N_24209,N_24218);
or U24360 (N_24360,N_24260,N_24254);
nand U24361 (N_24361,N_24251,N_24030);
xor U24362 (N_24362,N_24173,N_24100);
nand U24363 (N_24363,N_24102,N_24230);
xor U24364 (N_24364,N_24205,N_24084);
and U24365 (N_24365,N_24156,N_24151);
and U24366 (N_24366,N_24247,N_24203);
or U24367 (N_24367,N_24231,N_24283);
nand U24368 (N_24368,N_24052,N_24037);
or U24369 (N_24369,N_24273,N_24060);
xnor U24370 (N_24370,N_24005,N_24134);
nor U24371 (N_24371,N_24058,N_24202);
or U24372 (N_24372,N_24023,N_24174);
nand U24373 (N_24373,N_24071,N_24168);
xnor U24374 (N_24374,N_24011,N_24269);
and U24375 (N_24375,N_24122,N_24276);
and U24376 (N_24376,N_24036,N_24075);
xnor U24377 (N_24377,N_24192,N_24215);
xnor U24378 (N_24378,N_24041,N_24166);
nor U24379 (N_24379,N_24096,N_24149);
nor U24380 (N_24380,N_24264,N_24021);
xnor U24381 (N_24381,N_24196,N_24233);
xnor U24382 (N_24382,N_24089,N_24013);
or U24383 (N_24383,N_24063,N_24261);
and U24384 (N_24384,N_24243,N_24129);
nor U24385 (N_24385,N_24289,N_24004);
or U24386 (N_24386,N_24216,N_24064);
nor U24387 (N_24387,N_24073,N_24284);
and U24388 (N_24388,N_24187,N_24280);
or U24389 (N_24389,N_24132,N_24025);
nor U24390 (N_24390,N_24015,N_24238);
xor U24391 (N_24391,N_24176,N_24255);
nor U24392 (N_24392,N_24190,N_24138);
nor U24393 (N_24393,N_24008,N_24206);
xor U24394 (N_24394,N_24217,N_24006);
nor U24395 (N_24395,N_24092,N_24262);
nor U24396 (N_24396,N_24043,N_24067);
nor U24397 (N_24397,N_24212,N_24193);
and U24398 (N_24398,N_24062,N_24158);
or U24399 (N_24399,N_24213,N_24220);
nor U24400 (N_24400,N_24032,N_24110);
and U24401 (N_24401,N_24223,N_24252);
xnor U24402 (N_24402,N_24119,N_24144);
nor U24403 (N_24403,N_24002,N_24094);
or U24404 (N_24404,N_24140,N_24167);
and U24405 (N_24405,N_24103,N_24031);
and U24406 (N_24406,N_24081,N_24057);
or U24407 (N_24407,N_24127,N_24274);
nor U24408 (N_24408,N_24024,N_24059);
or U24409 (N_24409,N_24245,N_24281);
xnor U24410 (N_24410,N_24088,N_24044);
nand U24411 (N_24411,N_24234,N_24242);
and U24412 (N_24412,N_24141,N_24056);
or U24413 (N_24413,N_24271,N_24124);
nand U24414 (N_24414,N_24014,N_24199);
xnor U24415 (N_24415,N_24080,N_24297);
nor U24416 (N_24416,N_24222,N_24012);
nand U24417 (N_24417,N_24028,N_24194);
nand U24418 (N_24418,N_24189,N_24226);
nand U24419 (N_24419,N_24020,N_24086);
nand U24420 (N_24420,N_24017,N_24179);
and U24421 (N_24421,N_24069,N_24087);
nand U24422 (N_24422,N_24027,N_24070);
and U24423 (N_24423,N_24109,N_24026);
nand U24424 (N_24424,N_24010,N_24293);
nor U24425 (N_24425,N_24104,N_24266);
and U24426 (N_24426,N_24061,N_24034);
nand U24427 (N_24427,N_24082,N_24291);
or U24428 (N_24428,N_24022,N_24033);
xor U24429 (N_24429,N_24111,N_24170);
xor U24430 (N_24430,N_24115,N_24294);
xnor U24431 (N_24431,N_24117,N_24270);
and U24432 (N_24432,N_24072,N_24114);
and U24433 (N_24433,N_24065,N_24125);
nor U24434 (N_24434,N_24053,N_24143);
xnor U24435 (N_24435,N_24091,N_24292);
nor U24436 (N_24436,N_24237,N_24263);
nand U24437 (N_24437,N_24051,N_24204);
nor U24438 (N_24438,N_24171,N_24257);
nor U24439 (N_24439,N_24040,N_24157);
nor U24440 (N_24440,N_24097,N_24126);
nand U24441 (N_24441,N_24054,N_24219);
nand U24442 (N_24442,N_24221,N_24165);
nand U24443 (N_24443,N_24232,N_24009);
nand U24444 (N_24444,N_24211,N_24277);
nand U24445 (N_24445,N_24249,N_24112);
nand U24446 (N_24446,N_24188,N_24150);
xor U24447 (N_24447,N_24093,N_24016);
xnor U24448 (N_24448,N_24164,N_24246);
nor U24449 (N_24449,N_24287,N_24095);
xnor U24450 (N_24450,N_24297,N_24207);
nand U24451 (N_24451,N_24295,N_24037);
nand U24452 (N_24452,N_24034,N_24181);
and U24453 (N_24453,N_24089,N_24216);
nor U24454 (N_24454,N_24204,N_24156);
nand U24455 (N_24455,N_24181,N_24133);
or U24456 (N_24456,N_24116,N_24064);
nand U24457 (N_24457,N_24114,N_24206);
xnor U24458 (N_24458,N_24240,N_24201);
nand U24459 (N_24459,N_24281,N_24106);
nor U24460 (N_24460,N_24085,N_24020);
xor U24461 (N_24461,N_24178,N_24205);
xor U24462 (N_24462,N_24019,N_24150);
nand U24463 (N_24463,N_24046,N_24279);
xor U24464 (N_24464,N_24162,N_24259);
xor U24465 (N_24465,N_24290,N_24044);
or U24466 (N_24466,N_24196,N_24266);
nor U24467 (N_24467,N_24081,N_24281);
nand U24468 (N_24468,N_24209,N_24025);
and U24469 (N_24469,N_24109,N_24030);
nand U24470 (N_24470,N_24065,N_24258);
nor U24471 (N_24471,N_24181,N_24129);
nand U24472 (N_24472,N_24013,N_24256);
and U24473 (N_24473,N_24241,N_24047);
or U24474 (N_24474,N_24048,N_24238);
nor U24475 (N_24475,N_24173,N_24082);
nand U24476 (N_24476,N_24000,N_24107);
or U24477 (N_24477,N_24092,N_24005);
xnor U24478 (N_24478,N_24268,N_24068);
nand U24479 (N_24479,N_24251,N_24001);
and U24480 (N_24480,N_24000,N_24050);
and U24481 (N_24481,N_24040,N_24168);
nor U24482 (N_24482,N_24222,N_24238);
or U24483 (N_24483,N_24240,N_24236);
and U24484 (N_24484,N_24223,N_24010);
and U24485 (N_24485,N_24279,N_24030);
nor U24486 (N_24486,N_24252,N_24242);
nand U24487 (N_24487,N_24263,N_24002);
nor U24488 (N_24488,N_24177,N_24253);
nand U24489 (N_24489,N_24036,N_24261);
and U24490 (N_24490,N_24040,N_24274);
or U24491 (N_24491,N_24198,N_24120);
and U24492 (N_24492,N_24102,N_24251);
or U24493 (N_24493,N_24005,N_24073);
and U24494 (N_24494,N_24262,N_24068);
or U24495 (N_24495,N_24227,N_24106);
nand U24496 (N_24496,N_24294,N_24061);
nor U24497 (N_24497,N_24281,N_24291);
and U24498 (N_24498,N_24057,N_24105);
or U24499 (N_24499,N_24120,N_24278);
nand U24500 (N_24500,N_24004,N_24235);
xnor U24501 (N_24501,N_24266,N_24164);
xor U24502 (N_24502,N_24063,N_24108);
or U24503 (N_24503,N_24040,N_24020);
nor U24504 (N_24504,N_24123,N_24227);
nand U24505 (N_24505,N_24124,N_24075);
xnor U24506 (N_24506,N_24024,N_24006);
nor U24507 (N_24507,N_24209,N_24280);
nand U24508 (N_24508,N_24060,N_24186);
nand U24509 (N_24509,N_24174,N_24250);
nand U24510 (N_24510,N_24024,N_24042);
and U24511 (N_24511,N_24032,N_24299);
nor U24512 (N_24512,N_24179,N_24005);
nand U24513 (N_24513,N_24283,N_24031);
nor U24514 (N_24514,N_24000,N_24115);
xnor U24515 (N_24515,N_24119,N_24034);
nor U24516 (N_24516,N_24226,N_24059);
xor U24517 (N_24517,N_24254,N_24279);
or U24518 (N_24518,N_24139,N_24224);
xnor U24519 (N_24519,N_24177,N_24231);
nor U24520 (N_24520,N_24103,N_24196);
and U24521 (N_24521,N_24020,N_24064);
nor U24522 (N_24522,N_24014,N_24202);
and U24523 (N_24523,N_24017,N_24145);
nand U24524 (N_24524,N_24137,N_24193);
or U24525 (N_24525,N_24228,N_24026);
or U24526 (N_24526,N_24217,N_24157);
nand U24527 (N_24527,N_24118,N_24192);
xnor U24528 (N_24528,N_24150,N_24270);
or U24529 (N_24529,N_24051,N_24233);
xnor U24530 (N_24530,N_24091,N_24113);
and U24531 (N_24531,N_24021,N_24188);
or U24532 (N_24532,N_24250,N_24244);
nor U24533 (N_24533,N_24039,N_24294);
xor U24534 (N_24534,N_24077,N_24002);
nand U24535 (N_24535,N_24272,N_24150);
nand U24536 (N_24536,N_24213,N_24141);
and U24537 (N_24537,N_24183,N_24177);
or U24538 (N_24538,N_24102,N_24060);
or U24539 (N_24539,N_24263,N_24272);
and U24540 (N_24540,N_24037,N_24070);
or U24541 (N_24541,N_24266,N_24052);
nor U24542 (N_24542,N_24091,N_24034);
and U24543 (N_24543,N_24227,N_24069);
nand U24544 (N_24544,N_24093,N_24135);
nand U24545 (N_24545,N_24101,N_24017);
or U24546 (N_24546,N_24187,N_24285);
xor U24547 (N_24547,N_24159,N_24115);
and U24548 (N_24548,N_24095,N_24224);
or U24549 (N_24549,N_24086,N_24094);
xnor U24550 (N_24550,N_24229,N_24166);
and U24551 (N_24551,N_24128,N_24294);
nand U24552 (N_24552,N_24071,N_24079);
nor U24553 (N_24553,N_24159,N_24023);
xor U24554 (N_24554,N_24044,N_24195);
nand U24555 (N_24555,N_24256,N_24002);
nor U24556 (N_24556,N_24016,N_24175);
nand U24557 (N_24557,N_24226,N_24124);
nand U24558 (N_24558,N_24006,N_24058);
nor U24559 (N_24559,N_24011,N_24069);
nand U24560 (N_24560,N_24299,N_24048);
xnor U24561 (N_24561,N_24172,N_24049);
nor U24562 (N_24562,N_24240,N_24243);
xor U24563 (N_24563,N_24025,N_24110);
or U24564 (N_24564,N_24013,N_24122);
xor U24565 (N_24565,N_24099,N_24024);
nor U24566 (N_24566,N_24183,N_24144);
or U24567 (N_24567,N_24221,N_24166);
nand U24568 (N_24568,N_24147,N_24197);
nand U24569 (N_24569,N_24015,N_24052);
nand U24570 (N_24570,N_24038,N_24016);
nand U24571 (N_24571,N_24194,N_24169);
xnor U24572 (N_24572,N_24241,N_24223);
nand U24573 (N_24573,N_24183,N_24074);
and U24574 (N_24574,N_24164,N_24188);
nor U24575 (N_24575,N_24264,N_24016);
nor U24576 (N_24576,N_24257,N_24298);
or U24577 (N_24577,N_24238,N_24062);
nor U24578 (N_24578,N_24051,N_24012);
xor U24579 (N_24579,N_24269,N_24205);
xnor U24580 (N_24580,N_24251,N_24037);
or U24581 (N_24581,N_24068,N_24212);
or U24582 (N_24582,N_24260,N_24197);
xor U24583 (N_24583,N_24115,N_24256);
and U24584 (N_24584,N_24154,N_24111);
xnor U24585 (N_24585,N_24126,N_24294);
and U24586 (N_24586,N_24271,N_24062);
or U24587 (N_24587,N_24031,N_24112);
and U24588 (N_24588,N_24158,N_24145);
xor U24589 (N_24589,N_24105,N_24279);
nand U24590 (N_24590,N_24068,N_24147);
nand U24591 (N_24591,N_24175,N_24046);
and U24592 (N_24592,N_24246,N_24180);
or U24593 (N_24593,N_24263,N_24113);
and U24594 (N_24594,N_24214,N_24123);
xor U24595 (N_24595,N_24275,N_24106);
nor U24596 (N_24596,N_24255,N_24170);
or U24597 (N_24597,N_24253,N_24063);
nor U24598 (N_24598,N_24159,N_24069);
and U24599 (N_24599,N_24037,N_24260);
or U24600 (N_24600,N_24503,N_24302);
nand U24601 (N_24601,N_24515,N_24466);
or U24602 (N_24602,N_24598,N_24574);
and U24603 (N_24603,N_24569,N_24396);
nor U24604 (N_24604,N_24445,N_24392);
nor U24605 (N_24605,N_24481,N_24546);
nand U24606 (N_24606,N_24334,N_24349);
nand U24607 (N_24607,N_24456,N_24514);
and U24608 (N_24608,N_24372,N_24523);
xnor U24609 (N_24609,N_24439,N_24340);
xor U24610 (N_24610,N_24542,N_24432);
nand U24611 (N_24611,N_24560,N_24363);
and U24612 (N_24612,N_24527,N_24457);
nor U24613 (N_24613,N_24538,N_24433);
nand U24614 (N_24614,N_24468,N_24368);
xor U24615 (N_24615,N_24552,N_24477);
and U24616 (N_24616,N_24365,N_24380);
or U24617 (N_24617,N_24506,N_24354);
xor U24618 (N_24618,N_24545,N_24386);
nor U24619 (N_24619,N_24328,N_24597);
xnor U24620 (N_24620,N_24577,N_24572);
xor U24621 (N_24621,N_24374,N_24453);
nand U24622 (N_24622,N_24476,N_24424);
or U24623 (N_24623,N_24400,N_24504);
nand U24624 (N_24624,N_24492,N_24460);
nand U24625 (N_24625,N_24359,N_24357);
or U24626 (N_24626,N_24403,N_24406);
or U24627 (N_24627,N_24407,N_24384);
nor U24628 (N_24628,N_24440,N_24347);
nand U24629 (N_24629,N_24316,N_24423);
or U24630 (N_24630,N_24420,N_24304);
nor U24631 (N_24631,N_24570,N_24308);
nand U24632 (N_24632,N_24509,N_24511);
nor U24633 (N_24633,N_24534,N_24518);
nand U24634 (N_24634,N_24307,N_24490);
nor U24635 (N_24635,N_24376,N_24500);
nand U24636 (N_24636,N_24398,N_24556);
xnor U24637 (N_24637,N_24579,N_24554);
xor U24638 (N_24638,N_24418,N_24452);
and U24639 (N_24639,N_24459,N_24339);
nor U24640 (N_24640,N_24410,N_24350);
and U24641 (N_24641,N_24450,N_24564);
xnor U24642 (N_24642,N_24548,N_24411);
nor U24643 (N_24643,N_24348,N_24438);
nor U24644 (N_24644,N_24314,N_24487);
or U24645 (N_24645,N_24558,N_24409);
and U24646 (N_24646,N_24495,N_24342);
and U24647 (N_24647,N_24584,N_24362);
nor U24648 (N_24648,N_24448,N_24399);
nor U24649 (N_24649,N_24443,N_24371);
and U24650 (N_24650,N_24413,N_24532);
or U24651 (N_24651,N_24482,N_24581);
nand U24652 (N_24652,N_24563,N_24370);
xor U24653 (N_24653,N_24441,N_24303);
or U24654 (N_24654,N_24522,N_24306);
and U24655 (N_24655,N_24337,N_24344);
xor U24656 (N_24656,N_24305,N_24463);
and U24657 (N_24657,N_24589,N_24530);
xnor U24658 (N_24658,N_24402,N_24309);
or U24659 (N_24659,N_24341,N_24493);
or U24660 (N_24660,N_24462,N_24508);
nor U24661 (N_24661,N_24377,N_24507);
nand U24662 (N_24662,N_24580,N_24431);
xnor U24663 (N_24663,N_24549,N_24533);
and U24664 (N_24664,N_24395,N_24427);
or U24665 (N_24665,N_24381,N_24571);
xor U24666 (N_24666,N_24338,N_24486);
nor U24667 (N_24667,N_24329,N_24367);
or U24668 (N_24668,N_24578,N_24390);
nand U24669 (N_24669,N_24573,N_24575);
xnor U24670 (N_24670,N_24346,N_24461);
xnor U24671 (N_24671,N_24473,N_24586);
or U24672 (N_24672,N_24434,N_24378);
nand U24673 (N_24673,N_24470,N_24455);
xor U24674 (N_24674,N_24583,N_24414);
nor U24675 (N_24675,N_24393,N_24469);
or U24676 (N_24676,N_24526,N_24355);
and U24677 (N_24677,N_24385,N_24369);
nand U24678 (N_24678,N_24561,N_24528);
or U24679 (N_24679,N_24595,N_24480);
and U24680 (N_24680,N_24587,N_24336);
nand U24681 (N_24681,N_24512,N_24412);
and U24682 (N_24682,N_24557,N_24458);
xor U24683 (N_24683,N_24428,N_24590);
xnor U24684 (N_24684,N_24324,N_24425);
or U24685 (N_24685,N_24525,N_24536);
nor U24686 (N_24686,N_24405,N_24585);
xnor U24687 (N_24687,N_24352,N_24404);
and U24688 (N_24688,N_24547,N_24566);
or U24689 (N_24689,N_24442,N_24345);
or U24690 (N_24690,N_24332,N_24596);
xor U24691 (N_24691,N_24451,N_24543);
nor U24692 (N_24692,N_24373,N_24312);
xor U24693 (N_24693,N_24535,N_24421);
nor U24694 (N_24694,N_24498,N_24322);
nor U24695 (N_24695,N_24358,N_24464);
nor U24696 (N_24696,N_24553,N_24323);
or U24697 (N_24697,N_24517,N_24465);
or U24698 (N_24698,N_24388,N_24529);
or U24699 (N_24699,N_24300,N_24389);
xnor U24700 (N_24700,N_24568,N_24331);
nor U24701 (N_24701,N_24502,N_24576);
nor U24702 (N_24702,N_24524,N_24379);
nor U24703 (N_24703,N_24383,N_24429);
or U24704 (N_24704,N_24555,N_24397);
xor U24705 (N_24705,N_24335,N_24499);
nor U24706 (N_24706,N_24416,N_24483);
nor U24707 (N_24707,N_24419,N_24426);
and U24708 (N_24708,N_24479,N_24593);
nand U24709 (N_24709,N_24321,N_24550);
and U24710 (N_24710,N_24592,N_24594);
nor U24711 (N_24711,N_24531,N_24537);
or U24712 (N_24712,N_24494,N_24353);
nor U24713 (N_24713,N_24444,N_24467);
nand U24714 (N_24714,N_24565,N_24521);
nand U24715 (N_24715,N_24327,N_24520);
or U24716 (N_24716,N_24599,N_24505);
nor U24717 (N_24717,N_24484,N_24540);
or U24718 (N_24718,N_24516,N_24325);
nor U24719 (N_24719,N_24496,N_24510);
or U24720 (N_24720,N_24485,N_24366);
nand U24721 (N_24721,N_24311,N_24317);
nor U24722 (N_24722,N_24356,N_24401);
or U24723 (N_24723,N_24472,N_24360);
nand U24724 (N_24724,N_24582,N_24333);
or U24725 (N_24725,N_24539,N_24313);
nor U24726 (N_24726,N_24562,N_24422);
and U24727 (N_24727,N_24488,N_24320);
nand U24728 (N_24728,N_24437,N_24319);
xnor U24729 (N_24729,N_24567,N_24491);
nor U24730 (N_24730,N_24588,N_24559);
or U24731 (N_24731,N_24318,N_24454);
nor U24732 (N_24732,N_24301,N_24446);
nor U24733 (N_24733,N_24415,N_24361);
and U24734 (N_24734,N_24436,N_24375);
and U24735 (N_24735,N_24519,N_24343);
nand U24736 (N_24736,N_24501,N_24474);
and U24737 (N_24737,N_24326,N_24310);
and U24738 (N_24738,N_24351,N_24394);
nand U24739 (N_24739,N_24489,N_24478);
and U24740 (N_24740,N_24591,N_24497);
or U24741 (N_24741,N_24447,N_24382);
xor U24742 (N_24742,N_24513,N_24551);
nand U24743 (N_24743,N_24449,N_24391);
or U24744 (N_24744,N_24435,N_24364);
and U24745 (N_24745,N_24541,N_24475);
nand U24746 (N_24746,N_24417,N_24330);
and U24747 (N_24747,N_24315,N_24430);
or U24748 (N_24748,N_24387,N_24471);
and U24749 (N_24749,N_24408,N_24544);
nor U24750 (N_24750,N_24599,N_24344);
and U24751 (N_24751,N_24513,N_24440);
xnor U24752 (N_24752,N_24443,N_24413);
nand U24753 (N_24753,N_24397,N_24404);
or U24754 (N_24754,N_24584,N_24460);
nor U24755 (N_24755,N_24315,N_24495);
nor U24756 (N_24756,N_24521,N_24412);
nand U24757 (N_24757,N_24499,N_24416);
or U24758 (N_24758,N_24497,N_24422);
or U24759 (N_24759,N_24434,N_24335);
nor U24760 (N_24760,N_24520,N_24387);
nor U24761 (N_24761,N_24422,N_24549);
xor U24762 (N_24762,N_24368,N_24484);
nand U24763 (N_24763,N_24412,N_24336);
nor U24764 (N_24764,N_24473,N_24317);
nor U24765 (N_24765,N_24369,N_24597);
or U24766 (N_24766,N_24459,N_24306);
nor U24767 (N_24767,N_24379,N_24316);
and U24768 (N_24768,N_24432,N_24367);
and U24769 (N_24769,N_24486,N_24567);
nand U24770 (N_24770,N_24312,N_24396);
nand U24771 (N_24771,N_24523,N_24517);
and U24772 (N_24772,N_24591,N_24547);
or U24773 (N_24773,N_24342,N_24510);
xnor U24774 (N_24774,N_24315,N_24302);
and U24775 (N_24775,N_24392,N_24508);
and U24776 (N_24776,N_24597,N_24405);
nand U24777 (N_24777,N_24412,N_24456);
xor U24778 (N_24778,N_24575,N_24334);
nand U24779 (N_24779,N_24431,N_24597);
nor U24780 (N_24780,N_24392,N_24493);
xnor U24781 (N_24781,N_24510,N_24579);
nand U24782 (N_24782,N_24406,N_24350);
xor U24783 (N_24783,N_24488,N_24343);
nand U24784 (N_24784,N_24599,N_24393);
and U24785 (N_24785,N_24580,N_24484);
nand U24786 (N_24786,N_24457,N_24587);
nor U24787 (N_24787,N_24363,N_24553);
and U24788 (N_24788,N_24396,N_24321);
nand U24789 (N_24789,N_24352,N_24466);
nand U24790 (N_24790,N_24576,N_24499);
nand U24791 (N_24791,N_24593,N_24369);
or U24792 (N_24792,N_24552,N_24382);
nor U24793 (N_24793,N_24361,N_24380);
xor U24794 (N_24794,N_24315,N_24309);
nand U24795 (N_24795,N_24492,N_24307);
xnor U24796 (N_24796,N_24447,N_24310);
and U24797 (N_24797,N_24350,N_24599);
nand U24798 (N_24798,N_24323,N_24329);
or U24799 (N_24799,N_24391,N_24532);
xnor U24800 (N_24800,N_24445,N_24521);
nor U24801 (N_24801,N_24556,N_24562);
nor U24802 (N_24802,N_24429,N_24334);
xnor U24803 (N_24803,N_24321,N_24392);
nor U24804 (N_24804,N_24537,N_24512);
nand U24805 (N_24805,N_24413,N_24322);
xnor U24806 (N_24806,N_24381,N_24494);
nand U24807 (N_24807,N_24514,N_24530);
xnor U24808 (N_24808,N_24525,N_24330);
and U24809 (N_24809,N_24582,N_24383);
xor U24810 (N_24810,N_24483,N_24480);
xor U24811 (N_24811,N_24530,N_24317);
or U24812 (N_24812,N_24493,N_24501);
nor U24813 (N_24813,N_24488,N_24356);
or U24814 (N_24814,N_24318,N_24403);
xor U24815 (N_24815,N_24309,N_24342);
xnor U24816 (N_24816,N_24325,N_24395);
nor U24817 (N_24817,N_24320,N_24318);
nor U24818 (N_24818,N_24477,N_24546);
and U24819 (N_24819,N_24479,N_24422);
xor U24820 (N_24820,N_24425,N_24358);
xor U24821 (N_24821,N_24349,N_24379);
and U24822 (N_24822,N_24404,N_24556);
nor U24823 (N_24823,N_24522,N_24561);
nor U24824 (N_24824,N_24366,N_24591);
nand U24825 (N_24825,N_24491,N_24325);
or U24826 (N_24826,N_24534,N_24445);
xor U24827 (N_24827,N_24339,N_24301);
xor U24828 (N_24828,N_24560,N_24515);
and U24829 (N_24829,N_24417,N_24381);
nand U24830 (N_24830,N_24346,N_24424);
and U24831 (N_24831,N_24446,N_24443);
and U24832 (N_24832,N_24559,N_24310);
nand U24833 (N_24833,N_24362,N_24428);
or U24834 (N_24834,N_24543,N_24323);
and U24835 (N_24835,N_24471,N_24320);
or U24836 (N_24836,N_24579,N_24594);
xnor U24837 (N_24837,N_24398,N_24314);
xor U24838 (N_24838,N_24542,N_24325);
xnor U24839 (N_24839,N_24370,N_24447);
nor U24840 (N_24840,N_24408,N_24439);
nand U24841 (N_24841,N_24505,N_24303);
nand U24842 (N_24842,N_24582,N_24528);
nand U24843 (N_24843,N_24459,N_24572);
nor U24844 (N_24844,N_24312,N_24402);
nor U24845 (N_24845,N_24561,N_24544);
and U24846 (N_24846,N_24365,N_24452);
or U24847 (N_24847,N_24458,N_24336);
nand U24848 (N_24848,N_24578,N_24306);
nand U24849 (N_24849,N_24428,N_24430);
or U24850 (N_24850,N_24501,N_24382);
nand U24851 (N_24851,N_24468,N_24482);
xor U24852 (N_24852,N_24418,N_24506);
and U24853 (N_24853,N_24589,N_24394);
nand U24854 (N_24854,N_24563,N_24342);
nor U24855 (N_24855,N_24495,N_24482);
and U24856 (N_24856,N_24568,N_24377);
nor U24857 (N_24857,N_24479,N_24303);
nor U24858 (N_24858,N_24410,N_24476);
or U24859 (N_24859,N_24540,N_24476);
or U24860 (N_24860,N_24324,N_24451);
and U24861 (N_24861,N_24392,N_24317);
nand U24862 (N_24862,N_24387,N_24486);
and U24863 (N_24863,N_24455,N_24424);
and U24864 (N_24864,N_24478,N_24355);
or U24865 (N_24865,N_24579,N_24413);
xnor U24866 (N_24866,N_24578,N_24402);
nand U24867 (N_24867,N_24561,N_24341);
nor U24868 (N_24868,N_24309,N_24496);
and U24869 (N_24869,N_24439,N_24318);
nor U24870 (N_24870,N_24508,N_24594);
or U24871 (N_24871,N_24432,N_24459);
or U24872 (N_24872,N_24389,N_24375);
nor U24873 (N_24873,N_24594,N_24394);
nor U24874 (N_24874,N_24439,N_24525);
and U24875 (N_24875,N_24512,N_24323);
or U24876 (N_24876,N_24563,N_24432);
nor U24877 (N_24877,N_24589,N_24531);
nand U24878 (N_24878,N_24346,N_24438);
nor U24879 (N_24879,N_24403,N_24312);
xor U24880 (N_24880,N_24460,N_24359);
and U24881 (N_24881,N_24380,N_24385);
xor U24882 (N_24882,N_24445,N_24319);
and U24883 (N_24883,N_24412,N_24581);
or U24884 (N_24884,N_24476,N_24361);
or U24885 (N_24885,N_24462,N_24336);
or U24886 (N_24886,N_24314,N_24410);
or U24887 (N_24887,N_24448,N_24501);
or U24888 (N_24888,N_24552,N_24534);
nand U24889 (N_24889,N_24473,N_24320);
or U24890 (N_24890,N_24389,N_24482);
nor U24891 (N_24891,N_24582,N_24538);
and U24892 (N_24892,N_24424,N_24380);
and U24893 (N_24893,N_24398,N_24421);
or U24894 (N_24894,N_24495,N_24378);
xnor U24895 (N_24895,N_24577,N_24358);
and U24896 (N_24896,N_24376,N_24546);
and U24897 (N_24897,N_24488,N_24510);
and U24898 (N_24898,N_24497,N_24346);
or U24899 (N_24899,N_24357,N_24331);
or U24900 (N_24900,N_24621,N_24733);
and U24901 (N_24901,N_24685,N_24881);
nor U24902 (N_24902,N_24880,N_24724);
nand U24903 (N_24903,N_24776,N_24654);
nand U24904 (N_24904,N_24819,N_24703);
xnor U24905 (N_24905,N_24811,N_24648);
nand U24906 (N_24906,N_24879,N_24824);
xor U24907 (N_24907,N_24823,N_24647);
xor U24908 (N_24908,N_24661,N_24797);
nor U24909 (N_24909,N_24799,N_24759);
and U24910 (N_24910,N_24888,N_24731);
and U24911 (N_24911,N_24869,N_24637);
and U24912 (N_24912,N_24764,N_24610);
and U24913 (N_24913,N_24715,N_24625);
xor U24914 (N_24914,N_24605,N_24665);
nand U24915 (N_24915,N_24695,N_24690);
and U24916 (N_24916,N_24779,N_24747);
and U24917 (N_24917,N_24636,N_24650);
nor U24918 (N_24918,N_24868,N_24845);
or U24919 (N_24919,N_24633,N_24816);
xnor U24920 (N_24920,N_24886,N_24872);
and U24921 (N_24921,N_24600,N_24624);
or U24922 (N_24922,N_24667,N_24890);
nand U24923 (N_24923,N_24627,N_24607);
or U24924 (N_24924,N_24866,N_24889);
and U24925 (N_24925,N_24865,N_24662);
or U24926 (N_24926,N_24641,N_24856);
xor U24927 (N_24927,N_24660,N_24895);
nand U24928 (N_24928,N_24817,N_24773);
or U24929 (N_24929,N_24843,N_24796);
or U24930 (N_24930,N_24870,N_24707);
nor U24931 (N_24931,N_24739,N_24760);
nand U24932 (N_24932,N_24635,N_24602);
nor U24933 (N_24933,N_24896,N_24770);
nor U24934 (N_24934,N_24885,N_24812);
and U24935 (N_24935,N_24639,N_24678);
nand U24936 (N_24936,N_24780,N_24826);
xnor U24937 (N_24937,N_24728,N_24619);
or U24938 (N_24938,N_24882,N_24792);
xor U24939 (N_24939,N_24749,N_24814);
nand U24940 (N_24940,N_24751,N_24864);
and U24941 (N_24941,N_24734,N_24657);
and U24942 (N_24942,N_24804,N_24787);
nor U24943 (N_24943,N_24679,N_24850);
nand U24944 (N_24944,N_24626,N_24863);
nor U24945 (N_24945,N_24725,N_24651);
or U24946 (N_24946,N_24646,N_24709);
nand U24947 (N_24947,N_24744,N_24769);
xnor U24948 (N_24948,N_24653,N_24884);
nor U24949 (N_24949,N_24877,N_24673);
or U24950 (N_24950,N_24858,N_24839);
xnor U24951 (N_24951,N_24829,N_24798);
and U24952 (N_24952,N_24832,N_24887);
or U24953 (N_24953,N_24813,N_24748);
nand U24954 (N_24954,N_24701,N_24899);
and U24955 (N_24955,N_24846,N_24892);
nor U24956 (N_24956,N_24768,N_24743);
nor U24957 (N_24957,N_24807,N_24755);
nand U24958 (N_24958,N_24841,N_24805);
nor U24959 (N_24959,N_24615,N_24698);
nand U24960 (N_24960,N_24783,N_24855);
and U24961 (N_24961,N_24815,N_24758);
or U24962 (N_24962,N_24623,N_24831);
nor U24963 (N_24963,N_24828,N_24862);
or U24964 (N_24964,N_24871,N_24860);
or U24965 (N_24965,N_24849,N_24691);
nand U24966 (N_24966,N_24840,N_24613);
xor U24967 (N_24967,N_24774,N_24891);
xnor U24968 (N_24968,N_24794,N_24754);
nand U24969 (N_24969,N_24753,N_24622);
and U24970 (N_24970,N_24687,N_24677);
and U24971 (N_24971,N_24642,N_24717);
xnor U24972 (N_24972,N_24689,N_24767);
nor U24973 (N_24973,N_24874,N_24851);
or U24974 (N_24974,N_24752,N_24803);
nand U24975 (N_24975,N_24713,N_24785);
nand U24976 (N_24976,N_24762,N_24699);
nand U24977 (N_24977,N_24668,N_24740);
xor U24978 (N_24978,N_24810,N_24847);
nor U24979 (N_24979,N_24873,N_24655);
nor U24980 (N_24980,N_24837,N_24793);
nand U24981 (N_24981,N_24688,N_24848);
nor U24982 (N_24982,N_24852,N_24842);
xnor U24983 (N_24983,N_24620,N_24741);
or U24984 (N_24984,N_24737,N_24649);
or U24985 (N_24985,N_24763,N_24675);
and U24986 (N_24986,N_24696,N_24630);
xor U24987 (N_24987,N_24632,N_24683);
and U24988 (N_24988,N_24601,N_24612);
or U24989 (N_24989,N_24721,N_24634);
or U24990 (N_24990,N_24854,N_24761);
nand U24991 (N_24991,N_24844,N_24756);
xnor U24992 (N_24992,N_24676,N_24716);
or U24993 (N_24993,N_24827,N_24686);
and U24994 (N_24994,N_24789,N_24611);
and U24995 (N_24995,N_24857,N_24700);
nor U24996 (N_24996,N_24714,N_24784);
or U24997 (N_24997,N_24853,N_24712);
nand U24998 (N_24998,N_24818,N_24730);
and U24999 (N_24999,N_24684,N_24708);
nand U25000 (N_25000,N_24681,N_24656);
or U25001 (N_25001,N_24719,N_24875);
or U25002 (N_25002,N_24609,N_24859);
nor U25003 (N_25003,N_24736,N_24663);
and U25004 (N_25004,N_24788,N_24778);
xnor U25005 (N_25005,N_24883,N_24652);
nor U25006 (N_25006,N_24618,N_24772);
xnor U25007 (N_25007,N_24672,N_24617);
nand U25008 (N_25008,N_24838,N_24680);
and U25009 (N_25009,N_24729,N_24898);
or U25010 (N_25010,N_24834,N_24765);
and U25011 (N_25011,N_24745,N_24645);
nor U25012 (N_25012,N_24825,N_24629);
xor U25013 (N_25013,N_24746,N_24694);
nor U25014 (N_25014,N_24809,N_24658);
nand U25015 (N_25015,N_24718,N_24821);
or U25016 (N_25016,N_24790,N_24897);
nand U25017 (N_25017,N_24835,N_24836);
nor U25018 (N_25018,N_24893,N_24705);
nand U25019 (N_25019,N_24643,N_24781);
and U25020 (N_25020,N_24640,N_24861);
or U25021 (N_25021,N_24757,N_24666);
nor U25022 (N_25022,N_24750,N_24878);
and U25023 (N_25023,N_24723,N_24742);
and U25024 (N_25024,N_24771,N_24795);
xnor U25025 (N_25025,N_24604,N_24738);
xnor U25026 (N_25026,N_24766,N_24732);
or U25027 (N_25027,N_24659,N_24822);
nor U25028 (N_25028,N_24704,N_24735);
nor U25029 (N_25029,N_24692,N_24710);
or U25030 (N_25030,N_24867,N_24614);
nand U25031 (N_25031,N_24820,N_24894);
nand U25032 (N_25032,N_24801,N_24669);
xnor U25033 (N_25033,N_24786,N_24711);
nand U25034 (N_25034,N_24876,N_24808);
or U25035 (N_25035,N_24671,N_24830);
and U25036 (N_25036,N_24697,N_24616);
nor U25037 (N_25037,N_24706,N_24693);
xnor U25038 (N_25038,N_24702,N_24833);
nor U25039 (N_25039,N_24670,N_24727);
xnor U25040 (N_25040,N_24777,N_24631);
nand U25041 (N_25041,N_24806,N_24674);
nand U25042 (N_25042,N_24782,N_24628);
and U25043 (N_25043,N_24720,N_24606);
nor U25044 (N_25044,N_24603,N_24664);
nand U25045 (N_25045,N_24722,N_24638);
nor U25046 (N_25046,N_24608,N_24644);
and U25047 (N_25047,N_24791,N_24800);
xnor U25048 (N_25048,N_24775,N_24726);
xnor U25049 (N_25049,N_24682,N_24802);
or U25050 (N_25050,N_24873,N_24610);
nor U25051 (N_25051,N_24612,N_24791);
or U25052 (N_25052,N_24795,N_24648);
nor U25053 (N_25053,N_24715,N_24771);
nand U25054 (N_25054,N_24721,N_24724);
xnor U25055 (N_25055,N_24836,N_24844);
nor U25056 (N_25056,N_24805,N_24813);
nand U25057 (N_25057,N_24612,N_24622);
or U25058 (N_25058,N_24771,N_24762);
or U25059 (N_25059,N_24718,N_24799);
nand U25060 (N_25060,N_24725,N_24724);
or U25061 (N_25061,N_24773,N_24884);
xor U25062 (N_25062,N_24615,N_24660);
nor U25063 (N_25063,N_24666,N_24702);
xnor U25064 (N_25064,N_24837,N_24710);
and U25065 (N_25065,N_24660,N_24827);
or U25066 (N_25066,N_24636,N_24848);
and U25067 (N_25067,N_24852,N_24757);
or U25068 (N_25068,N_24772,N_24794);
xnor U25069 (N_25069,N_24869,N_24638);
nand U25070 (N_25070,N_24804,N_24892);
xor U25071 (N_25071,N_24707,N_24749);
xnor U25072 (N_25072,N_24670,N_24892);
or U25073 (N_25073,N_24605,N_24635);
or U25074 (N_25074,N_24720,N_24791);
nand U25075 (N_25075,N_24869,N_24784);
nand U25076 (N_25076,N_24837,N_24749);
nand U25077 (N_25077,N_24694,N_24877);
nand U25078 (N_25078,N_24676,N_24804);
xor U25079 (N_25079,N_24740,N_24607);
xor U25080 (N_25080,N_24614,N_24674);
nand U25081 (N_25081,N_24608,N_24814);
xor U25082 (N_25082,N_24684,N_24688);
or U25083 (N_25083,N_24753,N_24656);
or U25084 (N_25084,N_24846,N_24768);
and U25085 (N_25085,N_24887,N_24870);
and U25086 (N_25086,N_24648,N_24609);
xnor U25087 (N_25087,N_24804,N_24600);
nor U25088 (N_25088,N_24834,N_24692);
nand U25089 (N_25089,N_24877,N_24707);
nand U25090 (N_25090,N_24781,N_24822);
nand U25091 (N_25091,N_24885,N_24852);
xnor U25092 (N_25092,N_24733,N_24745);
nor U25093 (N_25093,N_24705,N_24880);
xnor U25094 (N_25094,N_24740,N_24857);
nand U25095 (N_25095,N_24705,N_24861);
nor U25096 (N_25096,N_24865,N_24681);
xnor U25097 (N_25097,N_24744,N_24614);
nor U25098 (N_25098,N_24723,N_24600);
and U25099 (N_25099,N_24709,N_24686);
nor U25100 (N_25100,N_24681,N_24809);
nand U25101 (N_25101,N_24710,N_24877);
xor U25102 (N_25102,N_24793,N_24702);
or U25103 (N_25103,N_24872,N_24899);
or U25104 (N_25104,N_24692,N_24687);
nand U25105 (N_25105,N_24712,N_24632);
nand U25106 (N_25106,N_24729,N_24623);
nor U25107 (N_25107,N_24685,N_24888);
nand U25108 (N_25108,N_24859,N_24631);
nand U25109 (N_25109,N_24772,N_24645);
nor U25110 (N_25110,N_24764,N_24746);
nand U25111 (N_25111,N_24880,N_24716);
nand U25112 (N_25112,N_24609,N_24776);
nor U25113 (N_25113,N_24686,N_24654);
xor U25114 (N_25114,N_24812,N_24632);
and U25115 (N_25115,N_24676,N_24611);
nand U25116 (N_25116,N_24622,N_24735);
and U25117 (N_25117,N_24695,N_24605);
nand U25118 (N_25118,N_24643,N_24713);
and U25119 (N_25119,N_24744,N_24727);
xor U25120 (N_25120,N_24854,N_24657);
xnor U25121 (N_25121,N_24614,N_24641);
and U25122 (N_25122,N_24700,N_24632);
nand U25123 (N_25123,N_24870,N_24743);
and U25124 (N_25124,N_24733,N_24701);
xnor U25125 (N_25125,N_24809,N_24882);
nor U25126 (N_25126,N_24722,N_24741);
nor U25127 (N_25127,N_24629,N_24787);
and U25128 (N_25128,N_24741,N_24768);
nand U25129 (N_25129,N_24770,N_24750);
nand U25130 (N_25130,N_24836,N_24623);
nor U25131 (N_25131,N_24657,N_24883);
xnor U25132 (N_25132,N_24710,N_24864);
nand U25133 (N_25133,N_24879,N_24846);
and U25134 (N_25134,N_24840,N_24624);
nor U25135 (N_25135,N_24667,N_24692);
nor U25136 (N_25136,N_24691,N_24662);
nor U25137 (N_25137,N_24786,N_24822);
nand U25138 (N_25138,N_24631,N_24898);
nand U25139 (N_25139,N_24622,N_24794);
nor U25140 (N_25140,N_24702,N_24831);
and U25141 (N_25141,N_24610,N_24828);
and U25142 (N_25142,N_24705,N_24653);
and U25143 (N_25143,N_24871,N_24897);
nand U25144 (N_25144,N_24735,N_24807);
xnor U25145 (N_25145,N_24643,N_24628);
xor U25146 (N_25146,N_24623,N_24783);
or U25147 (N_25147,N_24742,N_24695);
xor U25148 (N_25148,N_24644,N_24656);
xor U25149 (N_25149,N_24768,N_24807);
or U25150 (N_25150,N_24741,N_24650);
xnor U25151 (N_25151,N_24867,N_24649);
xnor U25152 (N_25152,N_24602,N_24705);
and U25153 (N_25153,N_24731,N_24892);
and U25154 (N_25154,N_24846,N_24857);
xnor U25155 (N_25155,N_24757,N_24706);
nor U25156 (N_25156,N_24611,N_24629);
nand U25157 (N_25157,N_24687,N_24666);
xor U25158 (N_25158,N_24671,N_24827);
nor U25159 (N_25159,N_24875,N_24674);
or U25160 (N_25160,N_24740,N_24765);
nand U25161 (N_25161,N_24735,N_24648);
and U25162 (N_25162,N_24747,N_24727);
xnor U25163 (N_25163,N_24600,N_24647);
xnor U25164 (N_25164,N_24712,N_24667);
nor U25165 (N_25165,N_24759,N_24769);
xnor U25166 (N_25166,N_24791,N_24701);
nor U25167 (N_25167,N_24787,N_24793);
and U25168 (N_25168,N_24878,N_24749);
nand U25169 (N_25169,N_24716,N_24779);
xnor U25170 (N_25170,N_24897,N_24646);
or U25171 (N_25171,N_24832,N_24623);
xnor U25172 (N_25172,N_24739,N_24847);
or U25173 (N_25173,N_24612,N_24733);
and U25174 (N_25174,N_24898,N_24836);
nand U25175 (N_25175,N_24606,N_24894);
nand U25176 (N_25176,N_24750,N_24631);
or U25177 (N_25177,N_24723,N_24631);
or U25178 (N_25178,N_24623,N_24635);
xnor U25179 (N_25179,N_24764,N_24693);
or U25180 (N_25180,N_24767,N_24633);
or U25181 (N_25181,N_24682,N_24612);
or U25182 (N_25182,N_24793,N_24681);
nand U25183 (N_25183,N_24797,N_24760);
nand U25184 (N_25184,N_24879,N_24757);
or U25185 (N_25185,N_24612,N_24774);
nand U25186 (N_25186,N_24722,N_24796);
and U25187 (N_25187,N_24823,N_24622);
xor U25188 (N_25188,N_24865,N_24877);
nand U25189 (N_25189,N_24833,N_24747);
and U25190 (N_25190,N_24859,N_24637);
or U25191 (N_25191,N_24736,N_24805);
and U25192 (N_25192,N_24680,N_24713);
nor U25193 (N_25193,N_24894,N_24721);
nand U25194 (N_25194,N_24896,N_24682);
nor U25195 (N_25195,N_24623,N_24611);
or U25196 (N_25196,N_24727,N_24708);
or U25197 (N_25197,N_24797,N_24871);
nor U25198 (N_25198,N_24837,N_24873);
nor U25199 (N_25199,N_24619,N_24857);
or U25200 (N_25200,N_25143,N_25038);
nor U25201 (N_25201,N_24949,N_25006);
or U25202 (N_25202,N_24975,N_25022);
nand U25203 (N_25203,N_25108,N_25020);
or U25204 (N_25204,N_24946,N_24916);
or U25205 (N_25205,N_25175,N_25054);
nand U25206 (N_25206,N_25059,N_25098);
and U25207 (N_25207,N_25080,N_25178);
and U25208 (N_25208,N_25104,N_24930);
xor U25209 (N_25209,N_25052,N_25088);
nand U25210 (N_25210,N_25172,N_25100);
xnor U25211 (N_25211,N_24910,N_25164);
nand U25212 (N_25212,N_24962,N_25153);
and U25213 (N_25213,N_24900,N_25189);
nor U25214 (N_25214,N_25049,N_25072);
xnor U25215 (N_25215,N_24904,N_25056);
and U25216 (N_25216,N_25169,N_25195);
nor U25217 (N_25217,N_24991,N_25018);
or U25218 (N_25218,N_24994,N_25176);
or U25219 (N_25219,N_24978,N_25087);
nand U25220 (N_25220,N_25057,N_25194);
and U25221 (N_25221,N_25086,N_24972);
or U25222 (N_25222,N_25065,N_25042);
nand U25223 (N_25223,N_24928,N_25013);
nand U25224 (N_25224,N_25003,N_24934);
and U25225 (N_25225,N_24971,N_24951);
xnor U25226 (N_25226,N_25117,N_25139);
nand U25227 (N_25227,N_24992,N_24931);
nand U25228 (N_25228,N_24985,N_25145);
or U25229 (N_25229,N_24909,N_25012);
nand U25230 (N_25230,N_25064,N_25029);
or U25231 (N_25231,N_24915,N_25190);
nor U25232 (N_25232,N_25127,N_25102);
nor U25233 (N_25233,N_25146,N_25103);
or U25234 (N_25234,N_24926,N_25083);
and U25235 (N_25235,N_24963,N_24917);
nand U25236 (N_25236,N_25024,N_25113);
xor U25237 (N_25237,N_25090,N_25135);
nand U25238 (N_25238,N_25151,N_24980);
nand U25239 (N_25239,N_25157,N_24990);
nor U25240 (N_25240,N_25063,N_25170);
xnor U25241 (N_25241,N_25046,N_25152);
or U25242 (N_25242,N_25133,N_24921);
or U25243 (N_25243,N_24936,N_25158);
nor U25244 (N_25244,N_25192,N_25047);
nor U25245 (N_25245,N_25036,N_25061);
nand U25246 (N_25246,N_25101,N_25082);
nor U25247 (N_25247,N_25150,N_25084);
or U25248 (N_25248,N_24922,N_25030);
nand U25249 (N_25249,N_25183,N_25159);
nand U25250 (N_25250,N_25193,N_25166);
nor U25251 (N_25251,N_25134,N_25004);
nor U25252 (N_25252,N_25031,N_25122);
xor U25253 (N_25253,N_25058,N_24970);
and U25254 (N_25254,N_24984,N_24913);
and U25255 (N_25255,N_25069,N_24997);
or U25256 (N_25256,N_25137,N_24943);
xnor U25257 (N_25257,N_25155,N_25026);
nand U25258 (N_25258,N_25132,N_25188);
nand U25259 (N_25259,N_24925,N_25111);
and U25260 (N_25260,N_25105,N_24924);
xor U25261 (N_25261,N_25180,N_25095);
and U25262 (N_25262,N_25125,N_25093);
and U25263 (N_25263,N_25162,N_25037);
or U25264 (N_25264,N_25089,N_25184);
or U25265 (N_25265,N_25067,N_24940);
nand U25266 (N_25266,N_25109,N_24906);
nor U25267 (N_25267,N_25051,N_24905);
xor U25268 (N_25268,N_25043,N_24976);
nand U25269 (N_25269,N_25110,N_25106);
or U25270 (N_25270,N_25199,N_24901);
xor U25271 (N_25271,N_24935,N_24929);
or U25272 (N_25272,N_25055,N_25039);
nor U25273 (N_25273,N_25021,N_24988);
xnor U25274 (N_25274,N_25015,N_24942);
or U25275 (N_25275,N_24989,N_24948);
nor U25276 (N_25276,N_25167,N_24950);
xor U25277 (N_25277,N_25077,N_25121);
nor U25278 (N_25278,N_25185,N_25142);
xnor U25279 (N_25279,N_25075,N_24974);
xnor U25280 (N_25280,N_25114,N_25023);
and U25281 (N_25281,N_25124,N_25187);
xnor U25282 (N_25282,N_25181,N_24961);
nor U25283 (N_25283,N_25073,N_24987);
nand U25284 (N_25284,N_25002,N_25070);
xor U25285 (N_25285,N_25144,N_24911);
and U25286 (N_25286,N_25034,N_25131);
nor U25287 (N_25287,N_25016,N_25148);
nor U25288 (N_25288,N_25094,N_24995);
nand U25289 (N_25289,N_25197,N_25160);
xor U25290 (N_25290,N_25091,N_24958);
nor U25291 (N_25291,N_24969,N_25040);
nor U25292 (N_25292,N_24902,N_24977);
or U25293 (N_25293,N_24933,N_25008);
or U25294 (N_25294,N_24998,N_25198);
or U25295 (N_25295,N_25182,N_25028);
or U25296 (N_25296,N_25156,N_25099);
nor U25297 (N_25297,N_25116,N_24945);
nor U25298 (N_25298,N_24966,N_25092);
or U25299 (N_25299,N_25071,N_25050);
xor U25300 (N_25300,N_25009,N_25096);
and U25301 (N_25301,N_25035,N_25032);
xor U25302 (N_25302,N_24954,N_25115);
nor U25303 (N_25303,N_25076,N_24912);
nand U25304 (N_25304,N_24944,N_24973);
or U25305 (N_25305,N_25000,N_25174);
xor U25306 (N_25306,N_25014,N_24956);
nand U25307 (N_25307,N_25112,N_25107);
xnor U25308 (N_25308,N_24947,N_24907);
nor U25309 (N_25309,N_24979,N_25141);
and U25310 (N_25310,N_25053,N_25097);
and U25311 (N_25311,N_25078,N_25007);
nor U25312 (N_25312,N_25027,N_24957);
nand U25313 (N_25313,N_25068,N_24952);
nor U25314 (N_25314,N_25130,N_24996);
or U25315 (N_25315,N_25079,N_25163);
and U25316 (N_25316,N_25129,N_24941);
nand U25317 (N_25317,N_25085,N_24932);
nor U25318 (N_25318,N_24960,N_24927);
nor U25319 (N_25319,N_25126,N_25177);
nand U25320 (N_25320,N_25001,N_24982);
nor U25321 (N_25321,N_24923,N_25168);
and U25322 (N_25322,N_25136,N_25123);
xnor U25323 (N_25323,N_25011,N_24999);
and U25324 (N_25324,N_25165,N_25048);
and U25325 (N_25325,N_25171,N_25149);
nor U25326 (N_25326,N_25119,N_24959);
or U25327 (N_25327,N_25140,N_25186);
nand U25328 (N_25328,N_25138,N_25196);
or U25329 (N_25329,N_25010,N_24918);
and U25330 (N_25330,N_25120,N_25066);
xor U25331 (N_25331,N_24968,N_24919);
nor U25332 (N_25332,N_25191,N_25044);
and U25333 (N_25333,N_24967,N_25173);
xor U25334 (N_25334,N_25161,N_25005);
or U25335 (N_25335,N_25045,N_25179);
nand U25336 (N_25336,N_25019,N_24993);
and U25337 (N_25337,N_24953,N_24955);
xor U25338 (N_25338,N_25154,N_24986);
or U25339 (N_25339,N_25147,N_25128);
xnor U25340 (N_25340,N_24903,N_24964);
nor U25341 (N_25341,N_25074,N_24920);
xnor U25342 (N_25342,N_24908,N_24914);
xor U25343 (N_25343,N_25033,N_25081);
nand U25344 (N_25344,N_25025,N_24939);
nor U25345 (N_25345,N_24965,N_25060);
nor U25346 (N_25346,N_24981,N_24937);
nor U25347 (N_25347,N_25062,N_24983);
nor U25348 (N_25348,N_25017,N_24938);
nand U25349 (N_25349,N_25041,N_25118);
nand U25350 (N_25350,N_25177,N_25134);
nand U25351 (N_25351,N_25110,N_25006);
nor U25352 (N_25352,N_25182,N_25136);
or U25353 (N_25353,N_25077,N_24940);
nand U25354 (N_25354,N_25135,N_25105);
xor U25355 (N_25355,N_25055,N_24962);
nand U25356 (N_25356,N_25030,N_25045);
and U25357 (N_25357,N_25028,N_25099);
and U25358 (N_25358,N_25018,N_24914);
and U25359 (N_25359,N_24999,N_24948);
nand U25360 (N_25360,N_25006,N_25127);
nor U25361 (N_25361,N_25142,N_25022);
xor U25362 (N_25362,N_25050,N_24945);
nand U25363 (N_25363,N_25086,N_25173);
nor U25364 (N_25364,N_25154,N_25006);
nand U25365 (N_25365,N_25026,N_25038);
xor U25366 (N_25366,N_25181,N_24954);
or U25367 (N_25367,N_25020,N_24996);
nand U25368 (N_25368,N_25115,N_24963);
and U25369 (N_25369,N_24981,N_25004);
xor U25370 (N_25370,N_25182,N_24997);
xor U25371 (N_25371,N_25038,N_24944);
nor U25372 (N_25372,N_25024,N_25173);
or U25373 (N_25373,N_25162,N_25196);
and U25374 (N_25374,N_25088,N_25076);
or U25375 (N_25375,N_25100,N_25070);
or U25376 (N_25376,N_25179,N_25177);
nand U25377 (N_25377,N_25070,N_25198);
nand U25378 (N_25378,N_24912,N_25041);
xor U25379 (N_25379,N_24982,N_25181);
or U25380 (N_25380,N_25107,N_25186);
and U25381 (N_25381,N_24956,N_24976);
or U25382 (N_25382,N_25098,N_25030);
nand U25383 (N_25383,N_25187,N_25038);
nand U25384 (N_25384,N_24907,N_24963);
or U25385 (N_25385,N_24913,N_25005);
nor U25386 (N_25386,N_24930,N_24926);
xor U25387 (N_25387,N_25052,N_24983);
nor U25388 (N_25388,N_25140,N_25180);
or U25389 (N_25389,N_25122,N_24960);
or U25390 (N_25390,N_25148,N_24967);
xnor U25391 (N_25391,N_25153,N_25176);
nand U25392 (N_25392,N_25078,N_25149);
xor U25393 (N_25393,N_25140,N_25090);
and U25394 (N_25394,N_25131,N_24953);
xor U25395 (N_25395,N_25010,N_24930);
xnor U25396 (N_25396,N_25036,N_25013);
or U25397 (N_25397,N_25058,N_24967);
nor U25398 (N_25398,N_25158,N_25124);
nor U25399 (N_25399,N_25063,N_25000);
and U25400 (N_25400,N_25050,N_25123);
nand U25401 (N_25401,N_24972,N_24934);
nor U25402 (N_25402,N_25101,N_24933);
and U25403 (N_25403,N_25041,N_25080);
and U25404 (N_25404,N_24913,N_25041);
xnor U25405 (N_25405,N_24929,N_25002);
nand U25406 (N_25406,N_25135,N_25016);
or U25407 (N_25407,N_25183,N_25104);
xnor U25408 (N_25408,N_24906,N_24949);
and U25409 (N_25409,N_24922,N_24955);
nand U25410 (N_25410,N_24952,N_25074);
nor U25411 (N_25411,N_25066,N_24980);
or U25412 (N_25412,N_25128,N_24962);
nor U25413 (N_25413,N_24956,N_24954);
nand U25414 (N_25414,N_24939,N_25096);
nand U25415 (N_25415,N_25144,N_25117);
xor U25416 (N_25416,N_25149,N_25061);
xnor U25417 (N_25417,N_24986,N_25077);
nand U25418 (N_25418,N_25026,N_24971);
xnor U25419 (N_25419,N_24986,N_25188);
nor U25420 (N_25420,N_24933,N_25052);
nor U25421 (N_25421,N_25143,N_24998);
nand U25422 (N_25422,N_25052,N_24955);
and U25423 (N_25423,N_24981,N_25044);
xor U25424 (N_25424,N_24936,N_24935);
nand U25425 (N_25425,N_25145,N_24984);
or U25426 (N_25426,N_25096,N_25010);
nand U25427 (N_25427,N_24905,N_24908);
xnor U25428 (N_25428,N_25113,N_25066);
nand U25429 (N_25429,N_25132,N_25100);
nand U25430 (N_25430,N_24952,N_25150);
xor U25431 (N_25431,N_24999,N_25082);
or U25432 (N_25432,N_24961,N_25121);
nor U25433 (N_25433,N_25009,N_24951);
xnor U25434 (N_25434,N_24965,N_24921);
or U25435 (N_25435,N_25145,N_25031);
or U25436 (N_25436,N_25173,N_25078);
or U25437 (N_25437,N_24952,N_24901);
xor U25438 (N_25438,N_24992,N_24947);
and U25439 (N_25439,N_25001,N_25117);
nand U25440 (N_25440,N_25066,N_25067);
and U25441 (N_25441,N_25046,N_24938);
nor U25442 (N_25442,N_25120,N_25155);
or U25443 (N_25443,N_24978,N_25064);
nor U25444 (N_25444,N_25166,N_25013);
or U25445 (N_25445,N_25186,N_25195);
or U25446 (N_25446,N_25148,N_25181);
and U25447 (N_25447,N_25045,N_24961);
and U25448 (N_25448,N_24939,N_25170);
or U25449 (N_25449,N_24928,N_25114);
or U25450 (N_25450,N_24974,N_25067);
and U25451 (N_25451,N_24906,N_25173);
and U25452 (N_25452,N_25052,N_25163);
and U25453 (N_25453,N_25101,N_25166);
nor U25454 (N_25454,N_25111,N_24910);
or U25455 (N_25455,N_25182,N_25133);
nor U25456 (N_25456,N_25194,N_24929);
xor U25457 (N_25457,N_24943,N_25158);
nand U25458 (N_25458,N_24987,N_25045);
nand U25459 (N_25459,N_25008,N_24925);
nand U25460 (N_25460,N_25124,N_24980);
and U25461 (N_25461,N_24933,N_25022);
nor U25462 (N_25462,N_25137,N_24907);
or U25463 (N_25463,N_25119,N_24994);
nor U25464 (N_25464,N_24959,N_25068);
xor U25465 (N_25465,N_24901,N_25109);
xnor U25466 (N_25466,N_25154,N_25076);
and U25467 (N_25467,N_25121,N_25046);
nor U25468 (N_25468,N_24955,N_25044);
xnor U25469 (N_25469,N_24970,N_25063);
or U25470 (N_25470,N_25129,N_25092);
and U25471 (N_25471,N_24982,N_25030);
nor U25472 (N_25472,N_24984,N_25029);
nand U25473 (N_25473,N_24990,N_25001);
nand U25474 (N_25474,N_25147,N_25078);
nand U25475 (N_25475,N_25156,N_24977);
and U25476 (N_25476,N_25156,N_24998);
nor U25477 (N_25477,N_25156,N_25166);
and U25478 (N_25478,N_25072,N_25047);
nor U25479 (N_25479,N_25133,N_24945);
or U25480 (N_25480,N_25169,N_24912);
and U25481 (N_25481,N_25123,N_25111);
nor U25482 (N_25482,N_25170,N_25012);
xor U25483 (N_25483,N_25032,N_24997);
nand U25484 (N_25484,N_25082,N_24937);
or U25485 (N_25485,N_24946,N_25007);
and U25486 (N_25486,N_25045,N_25017);
or U25487 (N_25487,N_25067,N_24939);
and U25488 (N_25488,N_24978,N_25106);
nor U25489 (N_25489,N_25070,N_25126);
and U25490 (N_25490,N_24924,N_25125);
nand U25491 (N_25491,N_25012,N_24903);
xor U25492 (N_25492,N_25188,N_25090);
xor U25493 (N_25493,N_25190,N_25046);
or U25494 (N_25494,N_24995,N_25142);
nor U25495 (N_25495,N_25157,N_24996);
and U25496 (N_25496,N_25127,N_24988);
and U25497 (N_25497,N_25147,N_24911);
nand U25498 (N_25498,N_24952,N_24912);
nand U25499 (N_25499,N_25066,N_25187);
nor U25500 (N_25500,N_25215,N_25311);
nand U25501 (N_25501,N_25297,N_25232);
and U25502 (N_25502,N_25286,N_25401);
or U25503 (N_25503,N_25205,N_25291);
xor U25504 (N_25504,N_25278,N_25436);
and U25505 (N_25505,N_25272,N_25496);
and U25506 (N_25506,N_25314,N_25387);
nand U25507 (N_25507,N_25200,N_25481);
nand U25508 (N_25508,N_25306,N_25470);
nand U25509 (N_25509,N_25270,N_25262);
or U25510 (N_25510,N_25488,N_25341);
nor U25511 (N_25511,N_25349,N_25449);
xor U25512 (N_25512,N_25428,N_25288);
nand U25513 (N_25513,N_25405,N_25203);
or U25514 (N_25514,N_25485,N_25279);
xnor U25515 (N_25515,N_25430,N_25337);
or U25516 (N_25516,N_25296,N_25440);
nand U25517 (N_25517,N_25421,N_25452);
nand U25518 (N_25518,N_25216,N_25475);
and U25519 (N_25519,N_25427,N_25357);
or U25520 (N_25520,N_25323,N_25395);
or U25521 (N_25521,N_25327,N_25422);
or U25522 (N_25522,N_25458,N_25444);
nor U25523 (N_25523,N_25378,N_25425);
nor U25524 (N_25524,N_25469,N_25487);
nand U25525 (N_25525,N_25313,N_25243);
xor U25526 (N_25526,N_25456,N_25301);
nor U25527 (N_25527,N_25354,N_25251);
nand U25528 (N_25528,N_25394,N_25379);
xor U25529 (N_25529,N_25446,N_25489);
and U25530 (N_25530,N_25256,N_25213);
or U25531 (N_25531,N_25237,N_25318);
or U25532 (N_25532,N_25331,N_25207);
nor U25533 (N_25533,N_25467,N_25273);
and U25534 (N_25534,N_25476,N_25375);
nand U25535 (N_25535,N_25201,N_25413);
or U25536 (N_25536,N_25265,N_25332);
and U25537 (N_25537,N_25439,N_25235);
or U25538 (N_25538,N_25453,N_25325);
xnor U25539 (N_25539,N_25420,N_25455);
nand U25540 (N_25540,N_25433,N_25477);
or U25541 (N_25541,N_25445,N_25239);
or U25542 (N_25542,N_25304,N_25385);
nand U25543 (N_25543,N_25204,N_25267);
nor U25544 (N_25544,N_25495,N_25217);
nor U25545 (N_25545,N_25211,N_25463);
and U25546 (N_25546,N_25490,N_25339);
or U25547 (N_25547,N_25462,N_25340);
nand U25548 (N_25548,N_25457,N_25284);
xnor U25549 (N_25549,N_25404,N_25266);
or U25550 (N_25550,N_25491,N_25231);
nor U25551 (N_25551,N_25329,N_25402);
and U25552 (N_25552,N_25434,N_25408);
xor U25553 (N_25553,N_25330,N_25376);
nand U25554 (N_25554,N_25257,N_25416);
and U25555 (N_25555,N_25355,N_25423);
xnor U25556 (N_25556,N_25233,N_25419);
nand U25557 (N_25557,N_25388,N_25308);
and U25558 (N_25558,N_25362,N_25206);
or U25559 (N_25559,N_25335,N_25365);
and U25560 (N_25560,N_25292,N_25260);
nor U25561 (N_25561,N_25380,N_25263);
xor U25562 (N_25562,N_25482,N_25367);
nand U25563 (N_25563,N_25303,N_25336);
or U25564 (N_25564,N_25448,N_25438);
and U25565 (N_25565,N_25221,N_25472);
xnor U25566 (N_25566,N_25363,N_25460);
nor U25567 (N_25567,N_25351,N_25499);
xor U25568 (N_25568,N_25236,N_25223);
or U25569 (N_25569,N_25412,N_25400);
nor U25570 (N_25570,N_25242,N_25326);
xnor U25571 (N_25571,N_25373,N_25210);
nand U25572 (N_25572,N_25299,N_25361);
nor U25573 (N_25573,N_25358,N_25240);
xnor U25574 (N_25574,N_25259,N_25426);
nand U25575 (N_25575,N_25468,N_25442);
and U25576 (N_25576,N_25268,N_25399);
nor U25577 (N_25577,N_25238,N_25281);
and U25578 (N_25578,N_25390,N_25492);
or U25579 (N_25579,N_25316,N_25271);
nand U25580 (N_25580,N_25209,N_25411);
nand U25581 (N_25581,N_25391,N_25437);
xor U25582 (N_25582,N_25319,N_25451);
or U25583 (N_25583,N_25396,N_25300);
xor U25584 (N_25584,N_25359,N_25377);
nand U25585 (N_25585,N_25353,N_25498);
nor U25586 (N_25586,N_25474,N_25224);
nor U25587 (N_25587,N_25334,N_25494);
and U25588 (N_25588,N_25246,N_25429);
or U25589 (N_25589,N_25285,N_25274);
xor U25590 (N_25590,N_25454,N_25352);
nor U25591 (N_25591,N_25407,N_25372);
or U25592 (N_25592,N_25219,N_25346);
nor U25593 (N_25593,N_25280,N_25295);
and U25594 (N_25594,N_25253,N_25366);
nor U25595 (N_25595,N_25381,N_25418);
or U25596 (N_25596,N_25447,N_25321);
nand U25597 (N_25597,N_25409,N_25208);
nand U25598 (N_25598,N_25461,N_25249);
and U25599 (N_25599,N_25302,N_25483);
xnor U25600 (N_25600,N_25252,N_25275);
nand U25601 (N_25601,N_25393,N_25320);
nand U25602 (N_25602,N_25383,N_25410);
xor U25603 (N_25603,N_25220,N_25225);
nor U25604 (N_25604,N_25269,N_25342);
nand U25605 (N_25605,N_25392,N_25347);
or U25606 (N_25606,N_25244,N_25228);
or U25607 (N_25607,N_25480,N_25368);
and U25608 (N_25608,N_25384,N_25431);
or U25609 (N_25609,N_25283,N_25360);
nor U25610 (N_25610,N_25369,N_25493);
or U25611 (N_25611,N_25374,N_25382);
xnor U25612 (N_25612,N_25294,N_25417);
and U25613 (N_25613,N_25486,N_25307);
or U25614 (N_25614,N_25234,N_25287);
or U25615 (N_25615,N_25214,N_25333);
nand U25616 (N_25616,N_25450,N_25276);
nor U25617 (N_25617,N_25471,N_25344);
xnor U25618 (N_25618,N_25356,N_25350);
nor U25619 (N_25619,N_25415,N_25254);
nor U25620 (N_25620,N_25226,N_25250);
or U25621 (N_25621,N_25441,N_25218);
xnor U25622 (N_25622,N_25345,N_25258);
and U25623 (N_25623,N_25465,N_25466);
xor U25624 (N_25624,N_25277,N_25290);
and U25625 (N_25625,N_25328,N_25222);
xnor U25626 (N_25626,N_25473,N_25424);
nand U25627 (N_25627,N_25371,N_25484);
and U25628 (N_25628,N_25264,N_25298);
xnor U25629 (N_25629,N_25310,N_25245);
nor U25630 (N_25630,N_25343,N_25293);
or U25631 (N_25631,N_25212,N_25414);
xor U25632 (N_25632,N_25247,N_25435);
nor U25633 (N_25633,N_25282,N_25348);
xnor U25634 (N_25634,N_25432,N_25230);
nor U25635 (N_25635,N_25406,N_25497);
nor U25636 (N_25636,N_25464,N_25317);
and U25637 (N_25637,N_25309,N_25386);
and U25638 (N_25638,N_25248,N_25338);
xnor U25639 (N_25639,N_25324,N_25202);
nor U25640 (N_25640,N_25241,N_25315);
and U25641 (N_25641,N_25459,N_25479);
nand U25642 (N_25642,N_25370,N_25255);
nor U25643 (N_25643,N_25364,N_25322);
xor U25644 (N_25644,N_25403,N_25227);
xnor U25645 (N_25645,N_25389,N_25478);
and U25646 (N_25646,N_25312,N_25261);
nand U25647 (N_25647,N_25398,N_25397);
nand U25648 (N_25648,N_25443,N_25229);
nand U25649 (N_25649,N_25305,N_25289);
nor U25650 (N_25650,N_25237,N_25294);
and U25651 (N_25651,N_25291,N_25308);
nor U25652 (N_25652,N_25201,N_25489);
or U25653 (N_25653,N_25390,N_25215);
nand U25654 (N_25654,N_25239,N_25485);
and U25655 (N_25655,N_25409,N_25359);
xnor U25656 (N_25656,N_25311,N_25455);
or U25657 (N_25657,N_25383,N_25235);
and U25658 (N_25658,N_25473,N_25395);
xor U25659 (N_25659,N_25321,N_25426);
nand U25660 (N_25660,N_25438,N_25398);
or U25661 (N_25661,N_25347,N_25352);
and U25662 (N_25662,N_25495,N_25486);
nand U25663 (N_25663,N_25444,N_25308);
and U25664 (N_25664,N_25375,N_25298);
nor U25665 (N_25665,N_25244,N_25279);
xor U25666 (N_25666,N_25379,N_25240);
and U25667 (N_25667,N_25253,N_25352);
nor U25668 (N_25668,N_25332,N_25425);
nand U25669 (N_25669,N_25243,N_25324);
xnor U25670 (N_25670,N_25459,N_25449);
or U25671 (N_25671,N_25420,N_25252);
nor U25672 (N_25672,N_25315,N_25406);
nor U25673 (N_25673,N_25239,N_25470);
or U25674 (N_25674,N_25439,N_25405);
nor U25675 (N_25675,N_25222,N_25449);
xnor U25676 (N_25676,N_25377,N_25282);
nand U25677 (N_25677,N_25366,N_25494);
or U25678 (N_25678,N_25361,N_25259);
xor U25679 (N_25679,N_25271,N_25201);
and U25680 (N_25680,N_25418,N_25250);
nor U25681 (N_25681,N_25405,N_25315);
nor U25682 (N_25682,N_25271,N_25392);
nor U25683 (N_25683,N_25464,N_25427);
xnor U25684 (N_25684,N_25267,N_25335);
xor U25685 (N_25685,N_25209,N_25279);
or U25686 (N_25686,N_25229,N_25449);
nor U25687 (N_25687,N_25414,N_25403);
xor U25688 (N_25688,N_25367,N_25263);
xor U25689 (N_25689,N_25419,N_25384);
xnor U25690 (N_25690,N_25351,N_25263);
and U25691 (N_25691,N_25346,N_25226);
or U25692 (N_25692,N_25360,N_25253);
xnor U25693 (N_25693,N_25449,N_25291);
nor U25694 (N_25694,N_25260,N_25426);
or U25695 (N_25695,N_25498,N_25451);
nand U25696 (N_25696,N_25472,N_25259);
or U25697 (N_25697,N_25207,N_25432);
nor U25698 (N_25698,N_25316,N_25429);
xor U25699 (N_25699,N_25382,N_25321);
or U25700 (N_25700,N_25264,N_25225);
and U25701 (N_25701,N_25341,N_25407);
or U25702 (N_25702,N_25231,N_25388);
nor U25703 (N_25703,N_25469,N_25402);
nand U25704 (N_25704,N_25344,N_25200);
nand U25705 (N_25705,N_25413,N_25433);
and U25706 (N_25706,N_25467,N_25217);
and U25707 (N_25707,N_25488,N_25268);
and U25708 (N_25708,N_25214,N_25390);
nand U25709 (N_25709,N_25283,N_25387);
or U25710 (N_25710,N_25223,N_25273);
nor U25711 (N_25711,N_25412,N_25209);
nor U25712 (N_25712,N_25354,N_25381);
or U25713 (N_25713,N_25302,N_25317);
nand U25714 (N_25714,N_25481,N_25400);
nor U25715 (N_25715,N_25499,N_25221);
xor U25716 (N_25716,N_25398,N_25420);
and U25717 (N_25717,N_25430,N_25299);
and U25718 (N_25718,N_25352,N_25218);
nor U25719 (N_25719,N_25385,N_25241);
nor U25720 (N_25720,N_25232,N_25360);
or U25721 (N_25721,N_25346,N_25345);
or U25722 (N_25722,N_25467,N_25412);
nor U25723 (N_25723,N_25235,N_25452);
and U25724 (N_25724,N_25327,N_25467);
nand U25725 (N_25725,N_25472,N_25443);
or U25726 (N_25726,N_25301,N_25232);
xnor U25727 (N_25727,N_25433,N_25328);
nand U25728 (N_25728,N_25453,N_25481);
or U25729 (N_25729,N_25471,N_25390);
xor U25730 (N_25730,N_25205,N_25457);
or U25731 (N_25731,N_25324,N_25323);
xor U25732 (N_25732,N_25335,N_25350);
nand U25733 (N_25733,N_25277,N_25281);
nor U25734 (N_25734,N_25430,N_25359);
or U25735 (N_25735,N_25341,N_25280);
xor U25736 (N_25736,N_25244,N_25221);
nor U25737 (N_25737,N_25257,N_25230);
xnor U25738 (N_25738,N_25274,N_25333);
xnor U25739 (N_25739,N_25245,N_25384);
or U25740 (N_25740,N_25317,N_25413);
nor U25741 (N_25741,N_25447,N_25341);
nor U25742 (N_25742,N_25479,N_25480);
and U25743 (N_25743,N_25461,N_25266);
or U25744 (N_25744,N_25338,N_25386);
and U25745 (N_25745,N_25260,N_25354);
and U25746 (N_25746,N_25427,N_25234);
nor U25747 (N_25747,N_25309,N_25221);
nand U25748 (N_25748,N_25237,N_25465);
nor U25749 (N_25749,N_25302,N_25438);
and U25750 (N_25750,N_25394,N_25468);
nand U25751 (N_25751,N_25317,N_25206);
nor U25752 (N_25752,N_25240,N_25258);
and U25753 (N_25753,N_25488,N_25400);
nor U25754 (N_25754,N_25224,N_25446);
nand U25755 (N_25755,N_25365,N_25481);
and U25756 (N_25756,N_25339,N_25402);
xor U25757 (N_25757,N_25359,N_25239);
or U25758 (N_25758,N_25301,N_25351);
or U25759 (N_25759,N_25219,N_25280);
xnor U25760 (N_25760,N_25309,N_25259);
xor U25761 (N_25761,N_25248,N_25305);
xnor U25762 (N_25762,N_25246,N_25398);
and U25763 (N_25763,N_25285,N_25428);
nor U25764 (N_25764,N_25289,N_25301);
and U25765 (N_25765,N_25442,N_25451);
and U25766 (N_25766,N_25497,N_25375);
xnor U25767 (N_25767,N_25293,N_25449);
nand U25768 (N_25768,N_25315,N_25208);
nor U25769 (N_25769,N_25463,N_25418);
or U25770 (N_25770,N_25395,N_25347);
and U25771 (N_25771,N_25465,N_25418);
and U25772 (N_25772,N_25428,N_25383);
and U25773 (N_25773,N_25345,N_25211);
nand U25774 (N_25774,N_25267,N_25289);
nor U25775 (N_25775,N_25303,N_25364);
xor U25776 (N_25776,N_25377,N_25445);
and U25777 (N_25777,N_25344,N_25300);
nor U25778 (N_25778,N_25359,N_25316);
nor U25779 (N_25779,N_25281,N_25466);
and U25780 (N_25780,N_25360,N_25486);
or U25781 (N_25781,N_25495,N_25423);
xor U25782 (N_25782,N_25490,N_25302);
and U25783 (N_25783,N_25211,N_25443);
or U25784 (N_25784,N_25237,N_25415);
xnor U25785 (N_25785,N_25365,N_25387);
nor U25786 (N_25786,N_25441,N_25231);
and U25787 (N_25787,N_25249,N_25479);
or U25788 (N_25788,N_25250,N_25241);
or U25789 (N_25789,N_25406,N_25235);
nand U25790 (N_25790,N_25219,N_25494);
or U25791 (N_25791,N_25252,N_25416);
xor U25792 (N_25792,N_25414,N_25492);
xnor U25793 (N_25793,N_25352,N_25405);
and U25794 (N_25794,N_25208,N_25299);
nand U25795 (N_25795,N_25321,N_25264);
and U25796 (N_25796,N_25371,N_25226);
and U25797 (N_25797,N_25262,N_25390);
nand U25798 (N_25798,N_25236,N_25278);
nand U25799 (N_25799,N_25240,N_25443);
or U25800 (N_25800,N_25605,N_25666);
nor U25801 (N_25801,N_25656,N_25718);
and U25802 (N_25802,N_25751,N_25600);
nand U25803 (N_25803,N_25717,N_25722);
or U25804 (N_25804,N_25681,N_25588);
xor U25805 (N_25805,N_25632,N_25532);
and U25806 (N_25806,N_25533,N_25747);
and U25807 (N_25807,N_25553,N_25797);
or U25808 (N_25808,N_25640,N_25779);
and U25809 (N_25809,N_25740,N_25522);
nand U25810 (N_25810,N_25508,N_25595);
nor U25811 (N_25811,N_25592,N_25556);
xnor U25812 (N_25812,N_25540,N_25650);
or U25813 (N_25813,N_25596,N_25619);
nand U25814 (N_25814,N_25559,N_25750);
nand U25815 (N_25815,N_25663,N_25597);
nor U25816 (N_25816,N_25539,N_25795);
nor U25817 (N_25817,N_25628,N_25626);
xnor U25818 (N_25818,N_25798,N_25775);
nor U25819 (N_25819,N_25618,N_25791);
and U25820 (N_25820,N_25564,N_25664);
nand U25821 (N_25821,N_25571,N_25748);
and U25822 (N_25822,N_25721,N_25506);
xor U25823 (N_25823,N_25661,N_25771);
or U25824 (N_25824,N_25613,N_25727);
nand U25825 (N_25825,N_25544,N_25547);
or U25826 (N_25826,N_25677,N_25786);
nor U25827 (N_25827,N_25662,N_25774);
or U25828 (N_25828,N_25711,N_25504);
nor U25829 (N_25829,N_25624,N_25788);
and U25830 (N_25830,N_25629,N_25693);
xor U25831 (N_25831,N_25582,N_25524);
nand U25832 (N_25832,N_25610,N_25554);
and U25833 (N_25833,N_25581,N_25646);
nor U25834 (N_25834,N_25660,N_25599);
and U25835 (N_25835,N_25578,N_25704);
nor U25836 (N_25836,N_25555,N_25793);
xnor U25837 (N_25837,N_25604,N_25558);
or U25838 (N_25838,N_25667,N_25754);
nor U25839 (N_25839,N_25591,N_25515);
or U25840 (N_25840,N_25616,N_25799);
nand U25841 (N_25841,N_25606,N_25525);
nor U25842 (N_25842,N_25659,N_25587);
nand U25843 (N_25843,N_25636,N_25520);
xor U25844 (N_25844,N_25701,N_25691);
and U25845 (N_25845,N_25777,N_25784);
nand U25846 (N_25846,N_25523,N_25541);
and U25847 (N_25847,N_25538,N_25696);
and U25848 (N_25848,N_25514,N_25526);
and U25849 (N_25849,N_25509,N_25676);
nand U25850 (N_25850,N_25776,N_25537);
nor U25851 (N_25851,N_25735,N_25726);
xor U25852 (N_25852,N_25723,N_25651);
or U25853 (N_25853,N_25607,N_25741);
xor U25854 (N_25854,N_25633,N_25725);
nand U25855 (N_25855,N_25694,N_25787);
or U25856 (N_25856,N_25762,N_25529);
nor U25857 (N_25857,N_25713,N_25567);
xnor U25858 (N_25858,N_25637,N_25627);
or U25859 (N_25859,N_25521,N_25589);
nor U25860 (N_25860,N_25579,N_25729);
nor U25861 (N_25861,N_25570,N_25734);
nor U25862 (N_25862,N_25736,N_25692);
or U25863 (N_25863,N_25766,N_25643);
nor U25864 (N_25864,N_25615,N_25732);
and U25865 (N_25865,N_25642,N_25789);
xnor U25866 (N_25866,N_25511,N_25796);
and U25867 (N_25867,N_25699,N_25546);
or U25868 (N_25868,N_25623,N_25565);
xor U25869 (N_25869,N_25697,N_25782);
and U25870 (N_25870,N_25769,N_25534);
nand U25871 (N_25871,N_25630,N_25738);
and U25872 (N_25872,N_25505,N_25703);
nand U25873 (N_25873,N_25728,N_25608);
and U25874 (N_25874,N_25654,N_25742);
nor U25875 (N_25875,N_25535,N_25683);
nand U25876 (N_25876,N_25707,N_25513);
or U25877 (N_25877,N_25719,N_25601);
nand U25878 (N_25878,N_25781,N_25716);
nor U25879 (N_25879,N_25647,N_25528);
nor U25880 (N_25880,N_25543,N_25580);
and U25881 (N_25881,N_25739,N_25687);
and U25882 (N_25882,N_25550,N_25764);
and U25883 (N_25883,N_25686,N_25552);
nor U25884 (N_25884,N_25503,N_25785);
or U25885 (N_25885,N_25756,N_25737);
nand U25886 (N_25886,N_25745,N_25573);
or U25887 (N_25887,N_25689,N_25566);
and U25888 (N_25888,N_25645,N_25631);
nor U25889 (N_25889,N_25768,N_25690);
nor U25890 (N_25890,N_25792,N_25670);
nand U25891 (N_25891,N_25702,N_25622);
or U25892 (N_25892,N_25593,N_25617);
nor U25893 (N_25893,N_25545,N_25575);
nand U25894 (N_25894,N_25744,N_25765);
or U25895 (N_25895,N_25767,N_25510);
or U25896 (N_25896,N_25583,N_25772);
and U25897 (N_25897,N_25652,N_25603);
nor U25898 (N_25898,N_25758,N_25743);
xor U25899 (N_25899,N_25568,N_25698);
nor U25900 (N_25900,N_25594,N_25609);
xnor U25901 (N_25901,N_25679,N_25598);
xor U25902 (N_25902,N_25653,N_25574);
nor U25903 (N_25903,N_25770,N_25635);
xnor U25904 (N_25904,N_25516,N_25531);
nand U25905 (N_25905,N_25576,N_25731);
and U25906 (N_25906,N_25527,N_25695);
xnor U25907 (N_25907,N_25519,N_25644);
and U25908 (N_25908,N_25730,N_25753);
or U25909 (N_25909,N_25548,N_25733);
or U25910 (N_25910,N_25557,N_25562);
or U25911 (N_25911,N_25705,N_25649);
nand U25912 (N_25912,N_25572,N_25639);
nor U25913 (N_25913,N_25678,N_25755);
and U25914 (N_25914,N_25673,N_25684);
or U25915 (N_25915,N_25634,N_25648);
and U25916 (N_25916,N_25674,N_25563);
or U25917 (N_25917,N_25586,N_25790);
and U25918 (N_25918,N_25680,N_25773);
xor U25919 (N_25919,N_25657,N_25668);
or U25920 (N_25920,N_25507,N_25706);
xnor U25921 (N_25921,N_25746,N_25512);
nand U25922 (N_25922,N_25763,N_25569);
or U25923 (N_25923,N_25672,N_25602);
and U25924 (N_25924,N_25549,N_25708);
nand U25925 (N_25925,N_25783,N_25518);
or U25926 (N_25926,N_25658,N_25502);
and U25927 (N_25927,N_25712,N_25584);
xnor U25928 (N_25928,N_25590,N_25778);
nand U25929 (N_25929,N_25709,N_25641);
nor U25930 (N_25930,N_25757,N_25625);
nand U25931 (N_25931,N_25585,N_25577);
or U25932 (N_25932,N_25685,N_25655);
nand U25933 (N_25933,N_25714,N_25682);
nand U25934 (N_25934,N_25560,N_25749);
nor U25935 (N_25935,N_25611,N_25638);
nor U25936 (N_25936,N_25551,N_25780);
nand U25937 (N_25937,N_25621,N_25501);
nor U25938 (N_25938,N_25710,N_25752);
nand U25939 (N_25939,N_25669,N_25620);
xnor U25940 (N_25940,N_25760,N_25724);
or U25941 (N_25941,N_25500,N_25536);
xor U25942 (N_25942,N_25517,N_25688);
nand U25943 (N_25943,N_25759,N_25675);
nor U25944 (N_25944,N_25612,N_25542);
and U25945 (N_25945,N_25761,N_25700);
nand U25946 (N_25946,N_25561,N_25614);
nand U25947 (N_25947,N_25671,N_25715);
or U25948 (N_25948,N_25794,N_25530);
nor U25949 (N_25949,N_25665,N_25720);
nor U25950 (N_25950,N_25702,N_25516);
nor U25951 (N_25951,N_25705,N_25622);
xnor U25952 (N_25952,N_25575,N_25690);
xor U25953 (N_25953,N_25547,N_25771);
xor U25954 (N_25954,N_25735,N_25794);
nor U25955 (N_25955,N_25543,N_25582);
and U25956 (N_25956,N_25770,N_25624);
nor U25957 (N_25957,N_25616,N_25586);
nand U25958 (N_25958,N_25666,N_25512);
nand U25959 (N_25959,N_25750,N_25659);
xnor U25960 (N_25960,N_25693,N_25746);
xor U25961 (N_25961,N_25746,N_25638);
and U25962 (N_25962,N_25581,N_25558);
or U25963 (N_25963,N_25539,N_25701);
nor U25964 (N_25964,N_25553,N_25572);
and U25965 (N_25965,N_25592,N_25612);
or U25966 (N_25966,N_25622,N_25601);
nand U25967 (N_25967,N_25789,N_25582);
nand U25968 (N_25968,N_25505,N_25565);
nand U25969 (N_25969,N_25595,N_25692);
nor U25970 (N_25970,N_25656,N_25672);
xnor U25971 (N_25971,N_25517,N_25666);
nor U25972 (N_25972,N_25657,N_25601);
nand U25973 (N_25973,N_25556,N_25648);
nor U25974 (N_25974,N_25734,N_25772);
xnor U25975 (N_25975,N_25616,N_25549);
and U25976 (N_25976,N_25629,N_25799);
xnor U25977 (N_25977,N_25502,N_25709);
nor U25978 (N_25978,N_25501,N_25714);
nand U25979 (N_25979,N_25610,N_25791);
nand U25980 (N_25980,N_25560,N_25548);
and U25981 (N_25981,N_25523,N_25598);
nor U25982 (N_25982,N_25658,N_25571);
nand U25983 (N_25983,N_25784,N_25755);
or U25984 (N_25984,N_25701,N_25785);
nor U25985 (N_25985,N_25644,N_25669);
xnor U25986 (N_25986,N_25676,N_25606);
or U25987 (N_25987,N_25775,N_25534);
nand U25988 (N_25988,N_25727,N_25737);
or U25989 (N_25989,N_25641,N_25529);
or U25990 (N_25990,N_25546,N_25789);
and U25991 (N_25991,N_25662,N_25740);
xor U25992 (N_25992,N_25786,N_25631);
and U25993 (N_25993,N_25650,N_25717);
and U25994 (N_25994,N_25606,N_25545);
and U25995 (N_25995,N_25682,N_25795);
xnor U25996 (N_25996,N_25546,N_25713);
or U25997 (N_25997,N_25538,N_25746);
nor U25998 (N_25998,N_25600,N_25596);
nand U25999 (N_25999,N_25785,N_25547);
nor U26000 (N_26000,N_25596,N_25565);
or U26001 (N_26001,N_25565,N_25797);
and U26002 (N_26002,N_25755,N_25555);
xnor U26003 (N_26003,N_25551,N_25776);
nand U26004 (N_26004,N_25610,N_25503);
nor U26005 (N_26005,N_25516,N_25676);
nor U26006 (N_26006,N_25503,N_25587);
or U26007 (N_26007,N_25501,N_25569);
and U26008 (N_26008,N_25611,N_25665);
and U26009 (N_26009,N_25666,N_25796);
or U26010 (N_26010,N_25580,N_25631);
or U26011 (N_26011,N_25675,N_25799);
or U26012 (N_26012,N_25710,N_25659);
xnor U26013 (N_26013,N_25540,N_25571);
and U26014 (N_26014,N_25511,N_25619);
nand U26015 (N_26015,N_25689,N_25570);
and U26016 (N_26016,N_25753,N_25557);
xnor U26017 (N_26017,N_25664,N_25750);
nand U26018 (N_26018,N_25588,N_25648);
or U26019 (N_26019,N_25519,N_25704);
nor U26020 (N_26020,N_25646,N_25670);
and U26021 (N_26021,N_25676,N_25599);
and U26022 (N_26022,N_25570,N_25610);
nor U26023 (N_26023,N_25517,N_25667);
xnor U26024 (N_26024,N_25662,N_25681);
nand U26025 (N_26025,N_25744,N_25530);
nor U26026 (N_26026,N_25714,N_25794);
nand U26027 (N_26027,N_25731,N_25584);
xnor U26028 (N_26028,N_25688,N_25510);
and U26029 (N_26029,N_25773,N_25737);
nor U26030 (N_26030,N_25674,N_25722);
and U26031 (N_26031,N_25522,N_25743);
or U26032 (N_26032,N_25560,N_25612);
xnor U26033 (N_26033,N_25781,N_25770);
xor U26034 (N_26034,N_25584,N_25575);
nand U26035 (N_26035,N_25541,N_25668);
nor U26036 (N_26036,N_25774,N_25691);
or U26037 (N_26037,N_25756,N_25588);
and U26038 (N_26038,N_25537,N_25662);
nor U26039 (N_26039,N_25631,N_25551);
and U26040 (N_26040,N_25501,N_25575);
nor U26041 (N_26041,N_25690,N_25547);
nor U26042 (N_26042,N_25773,N_25579);
nand U26043 (N_26043,N_25643,N_25745);
nand U26044 (N_26044,N_25624,N_25512);
nand U26045 (N_26045,N_25761,N_25782);
xor U26046 (N_26046,N_25524,N_25748);
nor U26047 (N_26047,N_25667,N_25619);
xor U26048 (N_26048,N_25585,N_25505);
or U26049 (N_26049,N_25736,N_25596);
xnor U26050 (N_26050,N_25768,N_25628);
and U26051 (N_26051,N_25712,N_25645);
and U26052 (N_26052,N_25529,N_25549);
and U26053 (N_26053,N_25788,N_25660);
nand U26054 (N_26054,N_25656,N_25658);
and U26055 (N_26055,N_25620,N_25521);
xnor U26056 (N_26056,N_25602,N_25647);
xor U26057 (N_26057,N_25732,N_25694);
xnor U26058 (N_26058,N_25634,N_25753);
and U26059 (N_26059,N_25516,N_25550);
or U26060 (N_26060,N_25628,N_25698);
and U26061 (N_26061,N_25724,N_25529);
nand U26062 (N_26062,N_25667,N_25510);
or U26063 (N_26063,N_25772,N_25754);
nand U26064 (N_26064,N_25746,N_25647);
xnor U26065 (N_26065,N_25687,N_25787);
nor U26066 (N_26066,N_25706,N_25550);
xnor U26067 (N_26067,N_25660,N_25756);
nor U26068 (N_26068,N_25776,N_25707);
and U26069 (N_26069,N_25606,N_25799);
nor U26070 (N_26070,N_25676,N_25678);
nand U26071 (N_26071,N_25524,N_25502);
xnor U26072 (N_26072,N_25669,N_25522);
nor U26073 (N_26073,N_25626,N_25505);
nand U26074 (N_26074,N_25751,N_25671);
nor U26075 (N_26075,N_25597,N_25557);
nand U26076 (N_26076,N_25785,N_25736);
xor U26077 (N_26077,N_25517,N_25786);
or U26078 (N_26078,N_25729,N_25503);
nor U26079 (N_26079,N_25750,N_25629);
or U26080 (N_26080,N_25722,N_25618);
xor U26081 (N_26081,N_25774,N_25766);
or U26082 (N_26082,N_25606,N_25514);
or U26083 (N_26083,N_25731,N_25755);
nor U26084 (N_26084,N_25730,N_25749);
xor U26085 (N_26085,N_25564,N_25615);
and U26086 (N_26086,N_25677,N_25567);
nand U26087 (N_26087,N_25578,N_25749);
or U26088 (N_26088,N_25798,N_25598);
or U26089 (N_26089,N_25589,N_25684);
nand U26090 (N_26090,N_25526,N_25797);
nand U26091 (N_26091,N_25713,N_25630);
and U26092 (N_26092,N_25762,N_25718);
or U26093 (N_26093,N_25504,N_25648);
nor U26094 (N_26094,N_25772,N_25675);
or U26095 (N_26095,N_25756,N_25635);
or U26096 (N_26096,N_25769,N_25551);
or U26097 (N_26097,N_25735,N_25533);
and U26098 (N_26098,N_25594,N_25777);
nand U26099 (N_26099,N_25696,N_25738);
xnor U26100 (N_26100,N_25837,N_25849);
nand U26101 (N_26101,N_25805,N_25903);
or U26102 (N_26102,N_25911,N_26009);
nand U26103 (N_26103,N_25986,N_25948);
and U26104 (N_26104,N_25852,N_25895);
or U26105 (N_26105,N_25821,N_25887);
nand U26106 (N_26106,N_25932,N_26053);
or U26107 (N_26107,N_25970,N_26082);
nand U26108 (N_26108,N_25961,N_25865);
nor U26109 (N_26109,N_26097,N_25872);
nor U26110 (N_26110,N_25934,N_25889);
nor U26111 (N_26111,N_25954,N_25910);
or U26112 (N_26112,N_25938,N_25807);
xnor U26113 (N_26113,N_25834,N_26014);
nor U26114 (N_26114,N_26029,N_25946);
nor U26115 (N_26115,N_25836,N_26032);
xor U26116 (N_26116,N_26078,N_25839);
nand U26117 (N_26117,N_25907,N_26060);
and U26118 (N_26118,N_25802,N_26070);
or U26119 (N_26119,N_25814,N_25813);
nor U26120 (N_26120,N_25994,N_26054);
nor U26121 (N_26121,N_25921,N_25806);
or U26122 (N_26122,N_25990,N_26081);
nor U26123 (N_26123,N_26061,N_25929);
xor U26124 (N_26124,N_25902,N_26089);
nand U26125 (N_26125,N_25982,N_26044);
xor U26126 (N_26126,N_25819,N_25888);
or U26127 (N_26127,N_25906,N_26091);
nor U26128 (N_26128,N_25965,N_25912);
or U26129 (N_26129,N_26028,N_25876);
xor U26130 (N_26130,N_26072,N_25960);
xnor U26131 (N_26131,N_25857,N_25815);
xor U26132 (N_26132,N_26008,N_25896);
nor U26133 (N_26133,N_26007,N_25962);
and U26134 (N_26134,N_25866,N_25973);
or U26135 (N_26135,N_25809,N_25920);
xor U26136 (N_26136,N_26083,N_25883);
nand U26137 (N_26137,N_25974,N_25999);
xnor U26138 (N_26138,N_25812,N_26079);
nand U26139 (N_26139,N_25848,N_25928);
nand U26140 (N_26140,N_26017,N_26036);
and U26141 (N_26141,N_25996,N_26074);
nand U26142 (N_26142,N_26006,N_25873);
xnor U26143 (N_26143,N_26095,N_26080);
nand U26144 (N_26144,N_26016,N_25984);
or U26145 (N_26145,N_26076,N_25987);
and U26146 (N_26146,N_25803,N_25882);
or U26147 (N_26147,N_25890,N_26033);
or U26148 (N_26148,N_25952,N_25944);
or U26149 (N_26149,N_25869,N_25936);
or U26150 (N_26150,N_25955,N_25884);
xor U26151 (N_26151,N_25918,N_25931);
nor U26152 (N_26152,N_25824,N_25957);
and U26153 (N_26153,N_25855,N_25941);
or U26154 (N_26154,N_26042,N_25816);
nand U26155 (N_26155,N_26005,N_25843);
nand U26156 (N_26156,N_25977,N_25923);
and U26157 (N_26157,N_26013,N_25831);
and U26158 (N_26158,N_26031,N_25879);
xnor U26159 (N_26159,N_26075,N_26030);
nor U26160 (N_26160,N_26049,N_25917);
or U26161 (N_26161,N_25959,N_26077);
nand U26162 (N_26162,N_26055,N_25886);
xor U26163 (N_26163,N_25925,N_25997);
nand U26164 (N_26164,N_26073,N_26010);
nand U26165 (N_26165,N_25945,N_26026);
nand U26166 (N_26166,N_25844,N_25893);
and U26167 (N_26167,N_25968,N_25826);
xnor U26168 (N_26168,N_25840,N_25971);
nor U26169 (N_26169,N_26067,N_26063);
and U26170 (N_26170,N_26022,N_25989);
xor U26171 (N_26171,N_25998,N_26001);
or U26172 (N_26172,N_25897,N_25940);
xnor U26173 (N_26173,N_26045,N_26098);
nor U26174 (N_26174,N_25991,N_26069);
and U26175 (N_26175,N_26037,N_25822);
and U26176 (N_26176,N_25862,N_26048);
and U26177 (N_26177,N_25851,N_25800);
xnor U26178 (N_26178,N_25874,N_25963);
xnor U26179 (N_26179,N_25995,N_26056);
xnor U26180 (N_26180,N_25828,N_26065);
or U26181 (N_26181,N_25801,N_25992);
xor U26182 (N_26182,N_25908,N_26025);
and U26183 (N_26183,N_25900,N_25892);
or U26184 (N_26184,N_26066,N_25985);
xnor U26185 (N_26185,N_25924,N_25956);
and U26186 (N_26186,N_25943,N_26086);
and U26187 (N_26187,N_25972,N_25919);
nor U26188 (N_26188,N_26062,N_26015);
nand U26189 (N_26189,N_25958,N_25850);
or U26190 (N_26190,N_26004,N_25841);
or U26191 (N_26191,N_26059,N_26003);
xor U26192 (N_26192,N_25926,N_25953);
or U26193 (N_26193,N_25845,N_25808);
nand U26194 (N_26194,N_25823,N_26002);
nor U26195 (N_26195,N_25878,N_25975);
or U26196 (N_26196,N_26018,N_25993);
nand U26197 (N_26197,N_25939,N_26041);
xor U26198 (N_26198,N_25885,N_25859);
or U26199 (N_26199,N_25820,N_25863);
and U26200 (N_26200,N_25942,N_25905);
xor U26201 (N_26201,N_25930,N_26027);
or U26202 (N_26202,N_26057,N_26052);
nand U26203 (N_26203,N_26051,N_25909);
and U26204 (N_26204,N_25833,N_25964);
xor U26205 (N_26205,N_25898,N_26085);
or U26206 (N_26206,N_26039,N_26047);
or U26207 (N_26207,N_26096,N_26064);
xor U26208 (N_26208,N_26050,N_26068);
nand U26209 (N_26209,N_26021,N_26012);
and U26210 (N_26210,N_25829,N_26000);
or U26211 (N_26211,N_25842,N_25935);
nor U26212 (N_26212,N_25933,N_25978);
or U26213 (N_26213,N_25853,N_26034);
nand U26214 (N_26214,N_25913,N_25832);
or U26215 (N_26215,N_26092,N_26023);
or U26216 (N_26216,N_26087,N_26035);
xnor U26217 (N_26217,N_25838,N_26084);
nor U26218 (N_26218,N_25868,N_25811);
nor U26219 (N_26219,N_25915,N_25875);
nand U26220 (N_26220,N_25976,N_25904);
nor U26221 (N_26221,N_26011,N_25827);
or U26222 (N_26222,N_25818,N_26090);
nand U26223 (N_26223,N_25856,N_25881);
and U26224 (N_26224,N_25810,N_25969);
nand U26225 (N_26225,N_25817,N_25830);
xor U26226 (N_26226,N_25846,N_25922);
and U26227 (N_26227,N_26038,N_25804);
nand U26228 (N_26228,N_26040,N_26020);
nor U26229 (N_26229,N_25966,N_26093);
nand U26230 (N_26230,N_25860,N_25835);
nand U26231 (N_26231,N_25891,N_25979);
xnor U26232 (N_26232,N_25854,N_25825);
or U26233 (N_26233,N_26046,N_25864);
or U26234 (N_26234,N_25867,N_25901);
xor U26235 (N_26235,N_26043,N_25988);
and U26236 (N_26236,N_25947,N_26071);
nand U26237 (N_26237,N_25847,N_25899);
or U26238 (N_26238,N_25877,N_25861);
xor U26239 (N_26239,N_25937,N_26058);
xnor U26240 (N_26240,N_25927,N_25981);
or U26241 (N_26241,N_25871,N_26088);
or U26242 (N_26242,N_25894,N_26019);
or U26243 (N_26243,N_26094,N_25914);
nand U26244 (N_26244,N_25870,N_25916);
and U26245 (N_26245,N_25949,N_26099);
xnor U26246 (N_26246,N_25951,N_25983);
xnor U26247 (N_26247,N_26024,N_25967);
or U26248 (N_26248,N_25880,N_25858);
nand U26249 (N_26249,N_25980,N_25950);
and U26250 (N_26250,N_25924,N_26098);
and U26251 (N_26251,N_25888,N_25960);
and U26252 (N_26252,N_25940,N_25813);
and U26253 (N_26253,N_25944,N_25807);
nand U26254 (N_26254,N_26068,N_25909);
nor U26255 (N_26255,N_25841,N_25967);
and U26256 (N_26256,N_26099,N_26078);
xor U26257 (N_26257,N_25986,N_25858);
xnor U26258 (N_26258,N_26071,N_26046);
nor U26259 (N_26259,N_26004,N_25887);
and U26260 (N_26260,N_25833,N_26032);
and U26261 (N_26261,N_26090,N_26049);
nand U26262 (N_26262,N_25956,N_25804);
nor U26263 (N_26263,N_26039,N_26093);
or U26264 (N_26264,N_26070,N_25841);
and U26265 (N_26265,N_25820,N_26055);
nor U26266 (N_26266,N_26016,N_25962);
or U26267 (N_26267,N_25858,N_26034);
and U26268 (N_26268,N_25845,N_26044);
and U26269 (N_26269,N_25946,N_25860);
nand U26270 (N_26270,N_25829,N_25854);
or U26271 (N_26271,N_25845,N_26066);
nand U26272 (N_26272,N_25971,N_25884);
and U26273 (N_26273,N_26065,N_25943);
and U26274 (N_26274,N_26035,N_25971);
or U26275 (N_26275,N_26008,N_25931);
xnor U26276 (N_26276,N_26047,N_26058);
or U26277 (N_26277,N_25895,N_25937);
nor U26278 (N_26278,N_25998,N_25968);
and U26279 (N_26279,N_26048,N_25982);
nand U26280 (N_26280,N_26073,N_26011);
or U26281 (N_26281,N_26052,N_26040);
nor U26282 (N_26282,N_26006,N_25808);
or U26283 (N_26283,N_25846,N_25911);
and U26284 (N_26284,N_25998,N_26016);
nand U26285 (N_26285,N_25884,N_25987);
or U26286 (N_26286,N_25983,N_25859);
or U26287 (N_26287,N_26094,N_25982);
nor U26288 (N_26288,N_25911,N_25946);
nand U26289 (N_26289,N_25839,N_25860);
xnor U26290 (N_26290,N_26081,N_25982);
or U26291 (N_26291,N_26048,N_26015);
or U26292 (N_26292,N_26042,N_25838);
or U26293 (N_26293,N_25991,N_25846);
xnor U26294 (N_26294,N_26013,N_25903);
xnor U26295 (N_26295,N_25954,N_26052);
nand U26296 (N_26296,N_26088,N_25999);
and U26297 (N_26297,N_26023,N_25838);
nand U26298 (N_26298,N_26077,N_25923);
xor U26299 (N_26299,N_25937,N_26057);
nor U26300 (N_26300,N_26051,N_26073);
or U26301 (N_26301,N_25951,N_26009);
or U26302 (N_26302,N_26022,N_25887);
or U26303 (N_26303,N_25948,N_26029);
or U26304 (N_26304,N_26048,N_25850);
xor U26305 (N_26305,N_25849,N_25843);
xor U26306 (N_26306,N_25862,N_25949);
nor U26307 (N_26307,N_25813,N_25877);
nor U26308 (N_26308,N_25969,N_25877);
nor U26309 (N_26309,N_25806,N_25853);
or U26310 (N_26310,N_25885,N_25923);
or U26311 (N_26311,N_25948,N_25899);
and U26312 (N_26312,N_25852,N_26051);
nor U26313 (N_26313,N_25872,N_26073);
nand U26314 (N_26314,N_25889,N_25858);
and U26315 (N_26315,N_25848,N_26084);
and U26316 (N_26316,N_26041,N_25931);
xnor U26317 (N_26317,N_25877,N_26028);
and U26318 (N_26318,N_26090,N_25845);
or U26319 (N_26319,N_26073,N_25977);
nor U26320 (N_26320,N_25816,N_25983);
or U26321 (N_26321,N_25825,N_25850);
nor U26322 (N_26322,N_25986,N_26015);
or U26323 (N_26323,N_26090,N_26027);
nor U26324 (N_26324,N_26057,N_26030);
nand U26325 (N_26325,N_25813,N_25812);
or U26326 (N_26326,N_25950,N_26010);
or U26327 (N_26327,N_26047,N_25807);
nor U26328 (N_26328,N_25879,N_25806);
and U26329 (N_26329,N_25910,N_25932);
or U26330 (N_26330,N_25994,N_25936);
nor U26331 (N_26331,N_26064,N_25979);
nor U26332 (N_26332,N_26079,N_25997);
nand U26333 (N_26333,N_25917,N_25833);
and U26334 (N_26334,N_25849,N_25804);
xor U26335 (N_26335,N_25819,N_26096);
and U26336 (N_26336,N_25806,N_26067);
xnor U26337 (N_26337,N_25957,N_25986);
or U26338 (N_26338,N_25944,N_25898);
xor U26339 (N_26339,N_25989,N_26037);
and U26340 (N_26340,N_25814,N_25972);
and U26341 (N_26341,N_26001,N_25853);
and U26342 (N_26342,N_25806,N_25823);
nor U26343 (N_26343,N_25886,N_26089);
xnor U26344 (N_26344,N_25862,N_25997);
or U26345 (N_26345,N_26068,N_25996);
or U26346 (N_26346,N_25800,N_26016);
nand U26347 (N_26347,N_25897,N_26017);
xnor U26348 (N_26348,N_25880,N_26023);
nand U26349 (N_26349,N_25877,N_25837);
or U26350 (N_26350,N_25841,N_26071);
and U26351 (N_26351,N_25957,N_26067);
nor U26352 (N_26352,N_25923,N_25875);
xnor U26353 (N_26353,N_25941,N_26085);
nand U26354 (N_26354,N_26085,N_25830);
nand U26355 (N_26355,N_25885,N_25823);
xor U26356 (N_26356,N_26079,N_25900);
xnor U26357 (N_26357,N_25946,N_26005);
or U26358 (N_26358,N_25977,N_26094);
nor U26359 (N_26359,N_26011,N_25934);
and U26360 (N_26360,N_26099,N_25910);
nor U26361 (N_26361,N_26066,N_25819);
or U26362 (N_26362,N_25938,N_25861);
or U26363 (N_26363,N_25955,N_25831);
and U26364 (N_26364,N_25927,N_25853);
nand U26365 (N_26365,N_26009,N_25840);
xor U26366 (N_26366,N_25824,N_25908);
xnor U26367 (N_26367,N_25911,N_25931);
nand U26368 (N_26368,N_26029,N_26021);
or U26369 (N_26369,N_25889,N_26096);
and U26370 (N_26370,N_25852,N_26039);
nor U26371 (N_26371,N_26002,N_25941);
or U26372 (N_26372,N_25850,N_25844);
and U26373 (N_26373,N_25883,N_25962);
nand U26374 (N_26374,N_26060,N_25981);
nor U26375 (N_26375,N_26063,N_25812);
and U26376 (N_26376,N_25981,N_25809);
and U26377 (N_26377,N_26050,N_26078);
nor U26378 (N_26378,N_25968,N_26004);
nand U26379 (N_26379,N_26086,N_25848);
or U26380 (N_26380,N_25864,N_25903);
nand U26381 (N_26381,N_25991,N_25921);
xnor U26382 (N_26382,N_25912,N_25977);
nand U26383 (N_26383,N_25835,N_26014);
and U26384 (N_26384,N_25829,N_25942);
or U26385 (N_26385,N_25950,N_25909);
and U26386 (N_26386,N_26051,N_25903);
or U26387 (N_26387,N_25954,N_25961);
and U26388 (N_26388,N_25971,N_25821);
xnor U26389 (N_26389,N_25842,N_25888);
nor U26390 (N_26390,N_25806,N_25810);
and U26391 (N_26391,N_25993,N_26014);
nor U26392 (N_26392,N_25936,N_25860);
nor U26393 (N_26393,N_26016,N_26071);
and U26394 (N_26394,N_25884,N_26035);
xor U26395 (N_26395,N_26038,N_25831);
nand U26396 (N_26396,N_26069,N_26024);
nor U26397 (N_26397,N_25827,N_25888);
nand U26398 (N_26398,N_25834,N_26058);
nor U26399 (N_26399,N_25963,N_25828);
xor U26400 (N_26400,N_26394,N_26242);
or U26401 (N_26401,N_26211,N_26370);
xor U26402 (N_26402,N_26160,N_26356);
nand U26403 (N_26403,N_26338,N_26215);
nand U26404 (N_26404,N_26247,N_26167);
nor U26405 (N_26405,N_26298,N_26210);
and U26406 (N_26406,N_26220,N_26339);
nor U26407 (N_26407,N_26152,N_26107);
xnor U26408 (N_26408,N_26119,N_26349);
or U26409 (N_26409,N_26116,N_26188);
xor U26410 (N_26410,N_26301,N_26348);
nand U26411 (N_26411,N_26121,N_26154);
nor U26412 (N_26412,N_26227,N_26129);
xor U26413 (N_26413,N_26282,N_26318);
nor U26414 (N_26414,N_26281,N_26104);
or U26415 (N_26415,N_26223,N_26102);
nand U26416 (N_26416,N_26390,N_26324);
or U26417 (N_26417,N_26212,N_26312);
nand U26418 (N_26418,N_26257,N_26326);
nand U26419 (N_26419,N_26249,N_26355);
nor U26420 (N_26420,N_26105,N_26137);
or U26421 (N_26421,N_26191,N_26114);
xnor U26422 (N_26422,N_26368,N_26149);
or U26423 (N_26423,N_26169,N_26251);
nor U26424 (N_26424,N_26381,N_26189);
nand U26425 (N_26425,N_26192,N_26358);
or U26426 (N_26426,N_26289,N_26205);
nor U26427 (N_26427,N_26385,N_26245);
and U26428 (N_26428,N_26311,N_26101);
xor U26429 (N_26429,N_26106,N_26214);
xnor U26430 (N_26430,N_26202,N_26283);
and U26431 (N_26431,N_26391,N_26206);
nor U26432 (N_26432,N_26269,N_26388);
nor U26433 (N_26433,N_26193,N_26310);
xor U26434 (N_26434,N_26316,N_26138);
nand U26435 (N_26435,N_26153,N_26264);
nand U26436 (N_26436,N_26239,N_26127);
or U26437 (N_26437,N_26181,N_26284);
nor U26438 (N_26438,N_26134,N_26243);
and U26439 (N_26439,N_26201,N_26131);
or U26440 (N_26440,N_26235,N_26158);
nor U26441 (N_26441,N_26250,N_26241);
xnor U26442 (N_26442,N_26331,N_26323);
xor U26443 (N_26443,N_26178,N_26186);
nor U26444 (N_26444,N_26360,N_26343);
and U26445 (N_26445,N_26329,N_26170);
nand U26446 (N_26446,N_26307,N_26268);
nor U26447 (N_26447,N_26180,N_26387);
or U26448 (N_26448,N_26353,N_26165);
xnor U26449 (N_26449,N_26159,N_26258);
xnor U26450 (N_26450,N_26109,N_26386);
and U26451 (N_26451,N_26150,N_26143);
nor U26452 (N_26452,N_26144,N_26313);
and U26453 (N_26453,N_26200,N_26110);
and U26454 (N_26454,N_26148,N_26304);
or U26455 (N_26455,N_26383,N_26330);
nand U26456 (N_26456,N_26378,N_26182);
nor U26457 (N_26457,N_26382,N_26184);
and U26458 (N_26458,N_26261,N_26233);
nor U26459 (N_26459,N_26364,N_26190);
xor U26460 (N_26460,N_26221,N_26285);
nand U26461 (N_26461,N_26142,N_26279);
nand U26462 (N_26462,N_26232,N_26396);
and U26463 (N_26463,N_26111,N_26224);
xnor U26464 (N_26464,N_26248,N_26197);
nor U26465 (N_26465,N_26240,N_26260);
nand U26466 (N_26466,N_26273,N_26128);
or U26467 (N_26467,N_26293,N_26136);
and U26468 (N_26468,N_26300,N_26347);
nor U26469 (N_26469,N_26276,N_26125);
and U26470 (N_26470,N_26229,N_26103);
nor U26471 (N_26471,N_26183,N_26267);
nor U26472 (N_26472,N_26342,N_26113);
and U26473 (N_26473,N_26203,N_26328);
nand U26474 (N_26474,N_26296,N_26286);
or U26475 (N_26475,N_26132,N_26108);
xor U26476 (N_26476,N_26333,N_26213);
nand U26477 (N_26477,N_26288,N_26246);
and U26478 (N_26478,N_26222,N_26265);
or U26479 (N_26479,N_26195,N_26367);
and U26480 (N_26480,N_26164,N_26147);
nand U26481 (N_26481,N_26397,N_26256);
or U26482 (N_26482,N_26322,N_26187);
xnor U26483 (N_26483,N_26295,N_26292);
xor U26484 (N_26484,N_26399,N_26126);
xor U26485 (N_26485,N_26179,N_26340);
nor U26486 (N_26486,N_26146,N_26274);
nand U26487 (N_26487,N_26327,N_26277);
nor U26488 (N_26488,N_26299,N_26365);
nor U26489 (N_26489,N_26162,N_26303);
nand U26490 (N_26490,N_26287,N_26357);
nand U26491 (N_26491,N_26384,N_26314);
and U26492 (N_26492,N_26325,N_26225);
or U26493 (N_26493,N_26361,N_26395);
or U26494 (N_26494,N_26175,N_26275);
nand U26495 (N_26495,N_26228,N_26157);
nor U26496 (N_26496,N_26135,N_26259);
nor U26497 (N_26497,N_26374,N_26163);
nand U26498 (N_26498,N_26117,N_26317);
nand U26499 (N_26499,N_26230,N_26161);
nand U26500 (N_26500,N_26253,N_26234);
or U26501 (N_26501,N_26209,N_26139);
nor U26502 (N_26502,N_26363,N_26392);
nand U26503 (N_26503,N_26315,N_26100);
and U26504 (N_26504,N_26321,N_26271);
nor U26505 (N_26505,N_26375,N_26306);
or U26506 (N_26506,N_26231,N_26112);
nor U26507 (N_26507,N_26207,N_26155);
and U26508 (N_26508,N_26236,N_26254);
nand U26509 (N_26509,N_26308,N_26359);
nor U26510 (N_26510,N_26172,N_26166);
nand U26511 (N_26511,N_26196,N_26297);
xnor U26512 (N_26512,N_26145,N_26290);
and U26513 (N_26513,N_26335,N_26336);
nor U26514 (N_26514,N_26217,N_26118);
xor U26515 (N_26515,N_26177,N_26173);
xor U26516 (N_26516,N_26244,N_26341);
nor U26517 (N_26517,N_26218,N_26130);
nand U26518 (N_26518,N_26369,N_26302);
nor U26519 (N_26519,N_26332,N_26352);
or U26520 (N_26520,N_26263,N_26262);
and U26521 (N_26521,N_26174,N_26171);
nor U26522 (N_26522,N_26372,N_26305);
or U26523 (N_26523,N_26123,N_26389);
xnor U26524 (N_26524,N_26270,N_26376);
xnor U26525 (N_26525,N_26226,N_26362);
and U26526 (N_26526,N_26278,N_26140);
or U26527 (N_26527,N_26194,N_26350);
and U26528 (N_26528,N_26345,N_26237);
and U26529 (N_26529,N_26373,N_26219);
or U26530 (N_26530,N_26133,N_26141);
xor U26531 (N_26531,N_26354,N_26122);
xor U26532 (N_26532,N_26344,N_26309);
nor U26533 (N_26533,N_26156,N_26379);
and U26534 (N_26534,N_26346,N_26371);
or U26535 (N_26535,N_26204,N_26272);
or U26536 (N_26536,N_26294,N_26208);
xor U26537 (N_26537,N_26377,N_26238);
and U26538 (N_26538,N_26334,N_26124);
and U26539 (N_26539,N_26216,N_26319);
xnor U26540 (N_26540,N_26120,N_26176);
or U26541 (N_26541,N_26115,N_26398);
xnor U26542 (N_26542,N_26393,N_26280);
nor U26543 (N_26543,N_26252,N_26351);
xor U26544 (N_26544,N_26151,N_26366);
and U26545 (N_26545,N_26291,N_26168);
nor U26546 (N_26546,N_26198,N_26199);
nor U26547 (N_26547,N_26337,N_26185);
or U26548 (N_26548,N_26380,N_26320);
xnor U26549 (N_26549,N_26266,N_26255);
and U26550 (N_26550,N_26116,N_26324);
nand U26551 (N_26551,N_26160,N_26315);
nor U26552 (N_26552,N_26269,N_26225);
nand U26553 (N_26553,N_26383,N_26343);
or U26554 (N_26554,N_26120,N_26225);
and U26555 (N_26555,N_26278,N_26202);
or U26556 (N_26556,N_26279,N_26161);
and U26557 (N_26557,N_26158,N_26279);
and U26558 (N_26558,N_26270,N_26150);
nor U26559 (N_26559,N_26396,N_26327);
nand U26560 (N_26560,N_26345,N_26143);
or U26561 (N_26561,N_26126,N_26274);
nor U26562 (N_26562,N_26392,N_26316);
xor U26563 (N_26563,N_26230,N_26332);
nor U26564 (N_26564,N_26170,N_26253);
and U26565 (N_26565,N_26373,N_26227);
xnor U26566 (N_26566,N_26385,N_26201);
xor U26567 (N_26567,N_26265,N_26233);
and U26568 (N_26568,N_26305,N_26203);
nor U26569 (N_26569,N_26254,N_26198);
or U26570 (N_26570,N_26200,N_26133);
or U26571 (N_26571,N_26318,N_26256);
or U26572 (N_26572,N_26285,N_26280);
nand U26573 (N_26573,N_26133,N_26219);
nor U26574 (N_26574,N_26248,N_26305);
nand U26575 (N_26575,N_26396,N_26347);
and U26576 (N_26576,N_26151,N_26329);
xor U26577 (N_26577,N_26166,N_26375);
or U26578 (N_26578,N_26250,N_26146);
nand U26579 (N_26579,N_26338,N_26186);
and U26580 (N_26580,N_26273,N_26152);
nor U26581 (N_26581,N_26107,N_26264);
or U26582 (N_26582,N_26303,N_26261);
nor U26583 (N_26583,N_26382,N_26124);
xnor U26584 (N_26584,N_26348,N_26364);
or U26585 (N_26585,N_26231,N_26242);
nor U26586 (N_26586,N_26359,N_26298);
nor U26587 (N_26587,N_26164,N_26149);
nand U26588 (N_26588,N_26381,N_26145);
nand U26589 (N_26589,N_26213,N_26373);
and U26590 (N_26590,N_26115,N_26247);
nor U26591 (N_26591,N_26354,N_26345);
or U26592 (N_26592,N_26397,N_26175);
xnor U26593 (N_26593,N_26219,N_26113);
nor U26594 (N_26594,N_26223,N_26167);
or U26595 (N_26595,N_26305,N_26304);
nand U26596 (N_26596,N_26365,N_26202);
and U26597 (N_26597,N_26186,N_26332);
and U26598 (N_26598,N_26266,N_26123);
nor U26599 (N_26599,N_26273,N_26193);
or U26600 (N_26600,N_26309,N_26220);
nor U26601 (N_26601,N_26343,N_26332);
xor U26602 (N_26602,N_26152,N_26149);
nor U26603 (N_26603,N_26244,N_26335);
nor U26604 (N_26604,N_26242,N_26144);
nand U26605 (N_26605,N_26145,N_26307);
nor U26606 (N_26606,N_26300,N_26370);
xor U26607 (N_26607,N_26160,N_26300);
xnor U26608 (N_26608,N_26392,N_26347);
and U26609 (N_26609,N_26314,N_26232);
xor U26610 (N_26610,N_26300,N_26288);
nand U26611 (N_26611,N_26107,N_26251);
xnor U26612 (N_26612,N_26160,N_26343);
or U26613 (N_26613,N_26338,N_26310);
and U26614 (N_26614,N_26296,N_26394);
nor U26615 (N_26615,N_26366,N_26354);
and U26616 (N_26616,N_26191,N_26346);
and U26617 (N_26617,N_26317,N_26397);
or U26618 (N_26618,N_26135,N_26181);
or U26619 (N_26619,N_26355,N_26233);
and U26620 (N_26620,N_26181,N_26361);
or U26621 (N_26621,N_26384,N_26142);
xor U26622 (N_26622,N_26368,N_26306);
and U26623 (N_26623,N_26296,N_26268);
or U26624 (N_26624,N_26126,N_26184);
or U26625 (N_26625,N_26331,N_26215);
nor U26626 (N_26626,N_26253,N_26326);
nand U26627 (N_26627,N_26221,N_26399);
nand U26628 (N_26628,N_26162,N_26290);
xor U26629 (N_26629,N_26315,N_26366);
nor U26630 (N_26630,N_26283,N_26393);
xor U26631 (N_26631,N_26309,N_26324);
nor U26632 (N_26632,N_26222,N_26396);
nand U26633 (N_26633,N_26300,N_26201);
xnor U26634 (N_26634,N_26224,N_26211);
nand U26635 (N_26635,N_26382,N_26262);
nor U26636 (N_26636,N_26246,N_26248);
nor U26637 (N_26637,N_26243,N_26229);
nor U26638 (N_26638,N_26359,N_26192);
or U26639 (N_26639,N_26139,N_26258);
nor U26640 (N_26640,N_26380,N_26134);
nand U26641 (N_26641,N_26213,N_26202);
and U26642 (N_26642,N_26359,N_26299);
nor U26643 (N_26643,N_26172,N_26197);
nand U26644 (N_26644,N_26152,N_26350);
xnor U26645 (N_26645,N_26253,N_26240);
or U26646 (N_26646,N_26206,N_26296);
xor U26647 (N_26647,N_26338,N_26321);
nor U26648 (N_26648,N_26269,N_26323);
nor U26649 (N_26649,N_26192,N_26325);
and U26650 (N_26650,N_26243,N_26373);
or U26651 (N_26651,N_26339,N_26234);
or U26652 (N_26652,N_26260,N_26123);
nor U26653 (N_26653,N_26165,N_26214);
and U26654 (N_26654,N_26216,N_26208);
xor U26655 (N_26655,N_26371,N_26110);
nor U26656 (N_26656,N_26389,N_26252);
nor U26657 (N_26657,N_26191,N_26289);
and U26658 (N_26658,N_26278,N_26376);
and U26659 (N_26659,N_26203,N_26109);
xor U26660 (N_26660,N_26319,N_26106);
xor U26661 (N_26661,N_26370,N_26330);
nand U26662 (N_26662,N_26180,N_26242);
xor U26663 (N_26663,N_26158,N_26147);
nor U26664 (N_26664,N_26187,N_26213);
nor U26665 (N_26665,N_26152,N_26110);
nand U26666 (N_26666,N_26267,N_26278);
xor U26667 (N_26667,N_26278,N_26119);
nor U26668 (N_26668,N_26293,N_26122);
and U26669 (N_26669,N_26268,N_26227);
or U26670 (N_26670,N_26137,N_26169);
xor U26671 (N_26671,N_26368,N_26120);
and U26672 (N_26672,N_26276,N_26121);
or U26673 (N_26673,N_26338,N_26217);
nand U26674 (N_26674,N_26118,N_26330);
nand U26675 (N_26675,N_26239,N_26282);
nor U26676 (N_26676,N_26216,N_26196);
nor U26677 (N_26677,N_26308,N_26325);
nor U26678 (N_26678,N_26316,N_26115);
nor U26679 (N_26679,N_26178,N_26136);
and U26680 (N_26680,N_26202,N_26226);
xor U26681 (N_26681,N_26362,N_26224);
and U26682 (N_26682,N_26393,N_26246);
xor U26683 (N_26683,N_26164,N_26195);
xnor U26684 (N_26684,N_26348,N_26217);
and U26685 (N_26685,N_26230,N_26357);
xor U26686 (N_26686,N_26220,N_26293);
nand U26687 (N_26687,N_26138,N_26339);
xor U26688 (N_26688,N_26387,N_26329);
xor U26689 (N_26689,N_26334,N_26317);
xor U26690 (N_26690,N_26121,N_26379);
nor U26691 (N_26691,N_26252,N_26190);
nand U26692 (N_26692,N_26299,N_26337);
and U26693 (N_26693,N_26350,N_26111);
or U26694 (N_26694,N_26265,N_26284);
nor U26695 (N_26695,N_26158,N_26209);
xnor U26696 (N_26696,N_26135,N_26291);
xnor U26697 (N_26697,N_26302,N_26196);
nand U26698 (N_26698,N_26351,N_26364);
nand U26699 (N_26699,N_26396,N_26395);
nand U26700 (N_26700,N_26517,N_26644);
and U26701 (N_26701,N_26491,N_26555);
xor U26702 (N_26702,N_26636,N_26525);
nand U26703 (N_26703,N_26419,N_26582);
xor U26704 (N_26704,N_26679,N_26569);
and U26705 (N_26705,N_26489,N_26461);
nor U26706 (N_26706,N_26691,N_26473);
nor U26707 (N_26707,N_26623,N_26523);
nand U26708 (N_26708,N_26513,N_26552);
nor U26709 (N_26709,N_26572,N_26422);
nor U26710 (N_26710,N_26418,N_26652);
nor U26711 (N_26711,N_26527,N_26415);
nand U26712 (N_26712,N_26465,N_26635);
nor U26713 (N_26713,N_26414,N_26588);
or U26714 (N_26714,N_26684,N_26509);
and U26715 (N_26715,N_26524,N_26455);
nand U26716 (N_26716,N_26549,N_26657);
or U26717 (N_26717,N_26618,N_26435);
xnor U26718 (N_26718,N_26602,N_26590);
nor U26719 (N_26719,N_26551,N_26463);
and U26720 (N_26720,N_26685,N_26406);
xor U26721 (N_26721,N_26655,N_26411);
xor U26722 (N_26722,N_26468,N_26457);
xor U26723 (N_26723,N_26470,N_26682);
and U26724 (N_26724,N_26615,N_26674);
xor U26725 (N_26725,N_26614,N_26548);
and U26726 (N_26726,N_26550,N_26454);
xor U26727 (N_26727,N_26677,N_26649);
or U26728 (N_26728,N_26420,N_26532);
or U26729 (N_26729,N_26646,N_26488);
and U26730 (N_26730,N_26421,N_26449);
xnor U26731 (N_26731,N_26499,N_26651);
or U26732 (N_26732,N_26570,N_26562);
or U26733 (N_26733,N_26583,N_26669);
nor U26734 (N_26734,N_26514,N_26633);
or U26735 (N_26735,N_26664,N_26497);
and U26736 (N_26736,N_26428,N_26687);
nor U26737 (N_26737,N_26476,N_26621);
nand U26738 (N_26738,N_26441,N_26486);
or U26739 (N_26739,N_26510,N_26451);
or U26740 (N_26740,N_26412,N_26403);
xnor U26741 (N_26741,N_26547,N_26681);
nand U26742 (N_26742,N_26650,N_26540);
and U26743 (N_26743,N_26627,N_26689);
nor U26744 (N_26744,N_26626,N_26611);
or U26745 (N_26745,N_26672,N_26542);
nor U26746 (N_26746,N_26563,N_26640);
and U26747 (N_26747,N_26595,N_26661);
xor U26748 (N_26748,N_26612,N_26413);
xnor U26749 (N_26749,N_26605,N_26586);
or U26750 (N_26750,N_26654,N_26637);
or U26751 (N_26751,N_26566,N_26668);
xnor U26752 (N_26752,N_26530,N_26622);
xor U26753 (N_26753,N_26466,N_26696);
or U26754 (N_26754,N_26653,N_26608);
and U26755 (N_26755,N_26643,N_26495);
and U26756 (N_26756,N_26528,N_26577);
or U26757 (N_26757,N_26401,N_26629);
and U26758 (N_26758,N_26581,N_26545);
xnor U26759 (N_26759,N_26444,N_26579);
or U26760 (N_26760,N_26560,N_26477);
nor U26761 (N_26761,N_26610,N_26553);
nand U26762 (N_26762,N_26592,N_26625);
nor U26763 (N_26763,N_26447,N_26405);
or U26764 (N_26764,N_26459,N_26506);
nand U26765 (N_26765,N_26460,N_26603);
and U26766 (N_26766,N_26537,N_26434);
and U26767 (N_26767,N_26500,N_26693);
nor U26768 (N_26768,N_26526,N_26642);
xor U26769 (N_26769,N_26539,N_26516);
or U26770 (N_26770,N_26452,N_26698);
xnor U26771 (N_26771,N_26648,N_26599);
and U26772 (N_26772,N_26502,N_26670);
or U26773 (N_26773,N_26515,N_26416);
nand U26774 (N_26774,N_26624,N_26439);
xnor U26775 (N_26775,N_26462,N_26641);
and U26776 (N_26776,N_26666,N_26609);
xor U26777 (N_26777,N_26505,N_26658);
or U26778 (N_26778,N_26587,N_26492);
or U26779 (N_26779,N_26559,N_26408);
xnor U26780 (N_26780,N_26593,N_26596);
nor U26781 (N_26781,N_26518,N_26409);
xor U26782 (N_26782,N_26519,N_26688);
xnor U26783 (N_26783,N_26564,N_26487);
or U26784 (N_26784,N_26673,N_26494);
xor U26785 (N_26785,N_26675,N_26561);
or U26786 (N_26786,N_26480,N_26432);
nand U26787 (N_26787,N_26680,N_26425);
nand U26788 (N_26788,N_26508,N_26558);
nor U26789 (N_26789,N_26667,N_26531);
or U26790 (N_26790,N_26472,N_26427);
nor U26791 (N_26791,N_26576,N_26503);
nor U26792 (N_26792,N_26541,N_26628);
and U26793 (N_26793,N_26662,N_26474);
nand U26794 (N_26794,N_26529,N_26695);
nand U26795 (N_26795,N_26630,N_26458);
or U26796 (N_26796,N_26607,N_26543);
xor U26797 (N_26797,N_26694,N_26521);
xnor U26798 (N_26798,N_26456,N_26511);
nand U26799 (N_26799,N_26634,N_26501);
and U26800 (N_26800,N_26546,N_26520);
and U26801 (N_26801,N_26697,N_26591);
or U26802 (N_26802,N_26571,N_26533);
nor U26803 (N_26803,N_26482,N_26446);
xor U26804 (N_26804,N_26601,N_26426);
xor U26805 (N_26805,N_26600,N_26638);
or U26806 (N_26806,N_26589,N_26443);
or U26807 (N_26807,N_26423,N_26678);
nor U26808 (N_26808,N_26479,N_26554);
nor U26809 (N_26809,N_26619,N_26557);
nand U26810 (N_26810,N_26597,N_26660);
xnor U26811 (N_26811,N_26690,N_26617);
xor U26812 (N_26812,N_26665,N_26431);
xor U26813 (N_26813,N_26437,N_26464);
xnor U26814 (N_26814,N_26481,N_26407);
and U26815 (N_26815,N_26498,N_26645);
nor U26816 (N_26816,N_26534,N_26632);
nand U26817 (N_26817,N_26469,N_26453);
and U26818 (N_26818,N_26556,N_26402);
xnor U26819 (N_26819,N_26671,N_26433);
nor U26820 (N_26820,N_26659,N_26536);
or U26821 (N_26821,N_26400,N_26493);
nand U26822 (N_26822,N_26538,N_26484);
nor U26823 (N_26823,N_26568,N_26440);
nand U26824 (N_26824,N_26496,N_26410);
xor U26825 (N_26825,N_26584,N_26567);
nand U26826 (N_26826,N_26699,N_26580);
or U26827 (N_26827,N_26471,N_26686);
or U26828 (N_26828,N_26573,N_26448);
xor U26829 (N_26829,N_26475,N_26535);
nor U26830 (N_26830,N_26504,N_26598);
and U26831 (N_26831,N_26613,N_26574);
xor U26832 (N_26832,N_26544,N_26442);
and U26833 (N_26833,N_26450,N_26483);
nor U26834 (N_26834,N_26436,N_26676);
nor U26835 (N_26835,N_26417,N_26692);
or U26836 (N_26836,N_26620,N_26522);
xor U26837 (N_26837,N_26445,N_26478);
xnor U26838 (N_26838,N_26467,N_26438);
and U26839 (N_26839,N_26578,N_26663);
and U26840 (N_26840,N_26656,N_26585);
xor U26841 (N_26841,N_26631,N_26683);
and U26842 (N_26842,N_26604,N_26647);
nand U26843 (N_26843,N_26616,N_26507);
or U26844 (N_26844,N_26424,N_26404);
and U26845 (N_26845,N_26606,N_26512);
and U26846 (N_26846,N_26565,N_26430);
nor U26847 (N_26847,N_26490,N_26485);
xor U26848 (N_26848,N_26429,N_26639);
nand U26849 (N_26849,N_26594,N_26575);
xor U26850 (N_26850,N_26473,N_26536);
xnor U26851 (N_26851,N_26637,N_26545);
and U26852 (N_26852,N_26601,N_26544);
nor U26853 (N_26853,N_26407,N_26500);
or U26854 (N_26854,N_26608,N_26635);
and U26855 (N_26855,N_26609,N_26482);
nor U26856 (N_26856,N_26544,N_26531);
xor U26857 (N_26857,N_26569,N_26435);
and U26858 (N_26858,N_26420,N_26578);
or U26859 (N_26859,N_26612,N_26469);
and U26860 (N_26860,N_26635,N_26695);
or U26861 (N_26861,N_26565,N_26529);
or U26862 (N_26862,N_26690,N_26610);
xnor U26863 (N_26863,N_26615,N_26477);
xor U26864 (N_26864,N_26496,N_26633);
nor U26865 (N_26865,N_26459,N_26440);
or U26866 (N_26866,N_26613,N_26673);
xor U26867 (N_26867,N_26581,N_26551);
nor U26868 (N_26868,N_26601,N_26600);
xor U26869 (N_26869,N_26694,N_26594);
or U26870 (N_26870,N_26442,N_26597);
nor U26871 (N_26871,N_26606,N_26684);
nor U26872 (N_26872,N_26490,N_26515);
or U26873 (N_26873,N_26486,N_26687);
and U26874 (N_26874,N_26579,N_26601);
xor U26875 (N_26875,N_26466,N_26607);
nor U26876 (N_26876,N_26409,N_26605);
and U26877 (N_26877,N_26474,N_26470);
nand U26878 (N_26878,N_26455,N_26551);
nor U26879 (N_26879,N_26623,N_26669);
nand U26880 (N_26880,N_26437,N_26420);
or U26881 (N_26881,N_26417,N_26642);
nand U26882 (N_26882,N_26449,N_26436);
or U26883 (N_26883,N_26491,N_26696);
xor U26884 (N_26884,N_26614,N_26542);
and U26885 (N_26885,N_26571,N_26424);
xnor U26886 (N_26886,N_26551,N_26676);
and U26887 (N_26887,N_26618,N_26678);
and U26888 (N_26888,N_26475,N_26456);
or U26889 (N_26889,N_26498,N_26443);
or U26890 (N_26890,N_26557,N_26498);
nor U26891 (N_26891,N_26633,N_26521);
nor U26892 (N_26892,N_26426,N_26592);
nor U26893 (N_26893,N_26514,N_26677);
nand U26894 (N_26894,N_26682,N_26556);
nand U26895 (N_26895,N_26610,N_26509);
and U26896 (N_26896,N_26515,N_26624);
and U26897 (N_26897,N_26514,N_26593);
or U26898 (N_26898,N_26576,N_26529);
nor U26899 (N_26899,N_26684,N_26489);
nand U26900 (N_26900,N_26456,N_26462);
and U26901 (N_26901,N_26491,N_26512);
and U26902 (N_26902,N_26596,N_26470);
nand U26903 (N_26903,N_26490,N_26683);
nand U26904 (N_26904,N_26435,N_26500);
or U26905 (N_26905,N_26562,N_26621);
xnor U26906 (N_26906,N_26585,N_26689);
nor U26907 (N_26907,N_26418,N_26637);
and U26908 (N_26908,N_26508,N_26425);
and U26909 (N_26909,N_26470,N_26458);
xnor U26910 (N_26910,N_26696,N_26564);
and U26911 (N_26911,N_26569,N_26481);
nor U26912 (N_26912,N_26483,N_26443);
nor U26913 (N_26913,N_26491,N_26563);
nor U26914 (N_26914,N_26522,N_26547);
and U26915 (N_26915,N_26467,N_26430);
and U26916 (N_26916,N_26606,N_26553);
or U26917 (N_26917,N_26663,N_26528);
and U26918 (N_26918,N_26504,N_26499);
or U26919 (N_26919,N_26451,N_26664);
nor U26920 (N_26920,N_26516,N_26520);
xnor U26921 (N_26921,N_26559,N_26627);
and U26922 (N_26922,N_26562,N_26417);
nor U26923 (N_26923,N_26634,N_26532);
nand U26924 (N_26924,N_26666,N_26491);
and U26925 (N_26925,N_26641,N_26624);
nand U26926 (N_26926,N_26632,N_26476);
nor U26927 (N_26927,N_26521,N_26499);
nor U26928 (N_26928,N_26400,N_26486);
and U26929 (N_26929,N_26674,N_26509);
nor U26930 (N_26930,N_26663,N_26635);
and U26931 (N_26931,N_26694,N_26546);
or U26932 (N_26932,N_26558,N_26650);
and U26933 (N_26933,N_26492,N_26643);
nand U26934 (N_26934,N_26456,N_26449);
and U26935 (N_26935,N_26513,N_26601);
and U26936 (N_26936,N_26414,N_26423);
and U26937 (N_26937,N_26499,N_26531);
nor U26938 (N_26938,N_26430,N_26687);
or U26939 (N_26939,N_26602,N_26565);
nand U26940 (N_26940,N_26559,N_26635);
and U26941 (N_26941,N_26400,N_26580);
nand U26942 (N_26942,N_26593,N_26501);
or U26943 (N_26943,N_26401,N_26669);
xor U26944 (N_26944,N_26645,N_26594);
and U26945 (N_26945,N_26512,N_26480);
or U26946 (N_26946,N_26517,N_26409);
and U26947 (N_26947,N_26640,N_26507);
nor U26948 (N_26948,N_26497,N_26493);
nor U26949 (N_26949,N_26538,N_26643);
xor U26950 (N_26950,N_26597,N_26650);
xnor U26951 (N_26951,N_26401,N_26566);
and U26952 (N_26952,N_26513,N_26662);
and U26953 (N_26953,N_26609,N_26527);
and U26954 (N_26954,N_26636,N_26495);
and U26955 (N_26955,N_26662,N_26480);
nand U26956 (N_26956,N_26685,N_26496);
nand U26957 (N_26957,N_26665,N_26522);
nand U26958 (N_26958,N_26573,N_26411);
and U26959 (N_26959,N_26505,N_26429);
or U26960 (N_26960,N_26682,N_26573);
or U26961 (N_26961,N_26408,N_26667);
and U26962 (N_26962,N_26480,N_26639);
or U26963 (N_26963,N_26592,N_26656);
or U26964 (N_26964,N_26433,N_26585);
nor U26965 (N_26965,N_26609,N_26573);
nor U26966 (N_26966,N_26653,N_26688);
xor U26967 (N_26967,N_26461,N_26567);
nor U26968 (N_26968,N_26488,N_26638);
and U26969 (N_26969,N_26649,N_26494);
nor U26970 (N_26970,N_26416,N_26689);
xnor U26971 (N_26971,N_26495,N_26469);
and U26972 (N_26972,N_26409,N_26681);
or U26973 (N_26973,N_26592,N_26650);
nor U26974 (N_26974,N_26501,N_26699);
or U26975 (N_26975,N_26424,N_26553);
or U26976 (N_26976,N_26470,N_26497);
nor U26977 (N_26977,N_26451,N_26607);
or U26978 (N_26978,N_26453,N_26665);
xor U26979 (N_26979,N_26533,N_26532);
nor U26980 (N_26980,N_26542,N_26557);
and U26981 (N_26981,N_26693,N_26480);
nand U26982 (N_26982,N_26497,N_26628);
xor U26983 (N_26983,N_26548,N_26557);
nor U26984 (N_26984,N_26685,N_26445);
and U26985 (N_26985,N_26424,N_26494);
or U26986 (N_26986,N_26608,N_26539);
nor U26987 (N_26987,N_26685,N_26643);
and U26988 (N_26988,N_26631,N_26429);
or U26989 (N_26989,N_26692,N_26607);
nor U26990 (N_26990,N_26419,N_26489);
nor U26991 (N_26991,N_26670,N_26469);
or U26992 (N_26992,N_26505,N_26420);
nand U26993 (N_26993,N_26586,N_26574);
xor U26994 (N_26994,N_26440,N_26453);
xor U26995 (N_26995,N_26488,N_26402);
nand U26996 (N_26996,N_26492,N_26548);
or U26997 (N_26997,N_26676,N_26444);
and U26998 (N_26998,N_26688,N_26594);
nor U26999 (N_26999,N_26452,N_26686);
and U27000 (N_27000,N_26901,N_26728);
or U27001 (N_27001,N_26951,N_26965);
and U27002 (N_27002,N_26733,N_26744);
and U27003 (N_27003,N_26860,N_26754);
and U27004 (N_27004,N_26748,N_26961);
or U27005 (N_27005,N_26762,N_26861);
and U27006 (N_27006,N_26954,N_26752);
xnor U27007 (N_27007,N_26932,N_26827);
or U27008 (N_27008,N_26843,N_26848);
nand U27009 (N_27009,N_26970,N_26996);
and U27010 (N_27010,N_26765,N_26830);
xor U27011 (N_27011,N_26947,N_26873);
nand U27012 (N_27012,N_26889,N_26858);
and U27013 (N_27013,N_26824,N_26972);
nand U27014 (N_27014,N_26891,N_26711);
nand U27015 (N_27015,N_26902,N_26914);
xnor U27016 (N_27016,N_26832,N_26903);
nand U27017 (N_27017,N_26995,N_26915);
nand U27018 (N_27018,N_26899,N_26785);
and U27019 (N_27019,N_26989,N_26809);
nand U27020 (N_27020,N_26781,N_26878);
xor U27021 (N_27021,N_26880,N_26730);
nand U27022 (N_27022,N_26774,N_26775);
nand U27023 (N_27023,N_26896,N_26799);
or U27024 (N_27024,N_26857,N_26723);
xnor U27025 (N_27025,N_26934,N_26950);
xnor U27026 (N_27026,N_26712,N_26983);
and U27027 (N_27027,N_26740,N_26713);
nor U27028 (N_27028,N_26945,N_26842);
xnor U27029 (N_27029,N_26869,N_26962);
nor U27030 (N_27030,N_26955,N_26791);
and U27031 (N_27031,N_26750,N_26795);
and U27032 (N_27032,N_26836,N_26770);
and U27033 (N_27033,N_26816,N_26909);
or U27034 (N_27034,N_26751,N_26802);
xnor U27035 (N_27035,N_26956,N_26724);
nand U27036 (N_27036,N_26773,N_26870);
nand U27037 (N_27037,N_26818,N_26786);
xor U27038 (N_27038,N_26892,N_26801);
nor U27039 (N_27039,N_26737,N_26722);
nor U27040 (N_27040,N_26831,N_26828);
nand U27041 (N_27041,N_26839,N_26783);
or U27042 (N_27042,N_26888,N_26700);
or U27043 (N_27043,N_26803,N_26985);
xnor U27044 (N_27044,N_26881,N_26953);
nand U27045 (N_27045,N_26859,N_26813);
or U27046 (N_27046,N_26979,N_26905);
nand U27047 (N_27047,N_26727,N_26731);
and U27048 (N_27048,N_26709,N_26768);
and U27049 (N_27049,N_26797,N_26837);
nand U27050 (N_27050,N_26850,N_26755);
and U27051 (N_27051,N_26845,N_26933);
nand U27052 (N_27052,N_26841,N_26912);
xor U27053 (N_27053,N_26810,N_26868);
xor U27054 (N_27054,N_26876,N_26884);
xnor U27055 (N_27055,N_26997,N_26968);
nor U27056 (N_27056,N_26817,N_26964);
and U27057 (N_27057,N_26906,N_26782);
or U27058 (N_27058,N_26990,N_26793);
xnor U27059 (N_27059,N_26745,N_26986);
and U27060 (N_27060,N_26998,N_26946);
xor U27061 (N_27061,N_26812,N_26917);
and U27062 (N_27062,N_26913,N_26936);
and U27063 (N_27063,N_26920,N_26777);
nand U27064 (N_27064,N_26833,N_26931);
and U27065 (N_27065,N_26764,N_26710);
xor U27066 (N_27066,N_26800,N_26838);
nand U27067 (N_27067,N_26821,N_26924);
nand U27068 (N_27068,N_26872,N_26987);
xnor U27069 (N_27069,N_26829,N_26811);
nand U27070 (N_27070,N_26703,N_26941);
nand U27071 (N_27071,N_26999,N_26796);
or U27072 (N_27072,N_26840,N_26957);
nor U27073 (N_27073,N_26792,N_26760);
or U27074 (N_27074,N_26784,N_26788);
xor U27075 (N_27075,N_26992,N_26980);
nand U27076 (N_27076,N_26994,N_26942);
xor U27077 (N_27077,N_26704,N_26926);
xor U27078 (N_27078,N_26823,N_26893);
and U27079 (N_27079,N_26807,N_26826);
nand U27080 (N_27080,N_26966,N_26715);
nand U27081 (N_27081,N_26875,N_26835);
and U27082 (N_27082,N_26767,N_26778);
xnor U27083 (N_27083,N_26769,N_26798);
xnor U27084 (N_27084,N_26976,N_26794);
or U27085 (N_27085,N_26834,N_26789);
nand U27086 (N_27086,N_26776,N_26981);
or U27087 (N_27087,N_26927,N_26805);
and U27088 (N_27088,N_26705,N_26988);
nand U27089 (N_27089,N_26758,N_26959);
nand U27090 (N_27090,N_26761,N_26707);
xnor U27091 (N_27091,N_26895,N_26719);
nand U27092 (N_27092,N_26701,N_26787);
nor U27093 (N_27093,N_26772,N_26949);
nor U27094 (N_27094,N_26874,N_26919);
or U27095 (N_27095,N_26819,N_26766);
and U27096 (N_27096,N_26739,N_26900);
xor U27097 (N_27097,N_26929,N_26897);
nor U27098 (N_27098,N_26944,N_26885);
nor U27099 (N_27099,N_26814,N_26721);
nor U27100 (N_27100,N_26939,N_26883);
and U27101 (N_27101,N_26882,N_26967);
xnor U27102 (N_27102,N_26851,N_26726);
nand U27103 (N_27103,N_26943,N_26742);
nand U27104 (N_27104,N_26863,N_26925);
and U27105 (N_27105,N_26763,N_26984);
nor U27106 (N_27106,N_26736,N_26973);
or U27107 (N_27107,N_26923,N_26908);
and U27108 (N_27108,N_26844,N_26907);
xnor U27109 (N_27109,N_26911,N_26928);
and U27110 (N_27110,N_26779,N_26978);
or U27111 (N_27111,N_26993,N_26977);
nor U27112 (N_27112,N_26771,N_26846);
and U27113 (N_27113,N_26852,N_26938);
xnor U27114 (N_27114,N_26756,N_26922);
and U27115 (N_27115,N_26804,N_26935);
nor U27116 (N_27116,N_26747,N_26790);
nor U27117 (N_27117,N_26865,N_26847);
nor U27118 (N_27118,N_26720,N_26749);
nand U27119 (N_27119,N_26971,N_26741);
or U27120 (N_27120,N_26717,N_26743);
and U27121 (N_27121,N_26871,N_26963);
nand U27122 (N_27122,N_26725,N_26822);
xor U27123 (N_27123,N_26759,N_26930);
or U27124 (N_27124,N_26849,N_26853);
nand U27125 (N_27125,N_26887,N_26702);
nor U27126 (N_27126,N_26815,N_26916);
or U27127 (N_27127,N_26854,N_26921);
nand U27128 (N_27128,N_26952,N_26877);
or U27129 (N_27129,N_26808,N_26714);
and U27130 (N_27130,N_26886,N_26856);
nor U27131 (N_27131,N_26937,N_26940);
nor U27132 (N_27132,N_26948,N_26820);
nor U27133 (N_27133,N_26974,N_26862);
nand U27134 (N_27134,N_26780,N_26910);
and U27135 (N_27135,N_26904,N_26894);
nor U27136 (N_27136,N_26866,N_26982);
nand U27137 (N_27137,N_26729,N_26706);
or U27138 (N_27138,N_26890,N_26975);
xor U27139 (N_27139,N_26806,N_26879);
nor U27140 (N_27140,N_26738,N_26718);
nor U27141 (N_27141,N_26969,N_26734);
and U27142 (N_27142,N_26991,N_26753);
nand U27143 (N_27143,N_26716,N_26746);
or U27144 (N_27144,N_26825,N_26918);
and U27145 (N_27145,N_26855,N_26867);
and U27146 (N_27146,N_26735,N_26757);
nand U27147 (N_27147,N_26898,N_26958);
xnor U27148 (N_27148,N_26708,N_26864);
xor U27149 (N_27149,N_26960,N_26732);
nor U27150 (N_27150,N_26802,N_26876);
nor U27151 (N_27151,N_26869,N_26989);
or U27152 (N_27152,N_26812,N_26817);
nor U27153 (N_27153,N_26767,N_26970);
or U27154 (N_27154,N_26963,N_26791);
nor U27155 (N_27155,N_26958,N_26930);
and U27156 (N_27156,N_26991,N_26700);
and U27157 (N_27157,N_26892,N_26894);
xnor U27158 (N_27158,N_26883,N_26875);
xor U27159 (N_27159,N_26937,N_26830);
nand U27160 (N_27160,N_26818,N_26759);
nor U27161 (N_27161,N_26797,N_26826);
xor U27162 (N_27162,N_26968,N_26793);
xnor U27163 (N_27163,N_26857,N_26970);
xor U27164 (N_27164,N_26935,N_26997);
nor U27165 (N_27165,N_26981,N_26914);
and U27166 (N_27166,N_26810,N_26726);
nand U27167 (N_27167,N_26845,N_26909);
and U27168 (N_27168,N_26740,N_26925);
or U27169 (N_27169,N_26830,N_26952);
xnor U27170 (N_27170,N_26994,N_26880);
xor U27171 (N_27171,N_26983,N_26998);
xnor U27172 (N_27172,N_26967,N_26897);
nand U27173 (N_27173,N_26879,N_26924);
or U27174 (N_27174,N_26905,N_26779);
or U27175 (N_27175,N_26914,N_26758);
or U27176 (N_27176,N_26885,N_26752);
or U27177 (N_27177,N_26933,N_26758);
and U27178 (N_27178,N_26898,N_26983);
xor U27179 (N_27179,N_26787,N_26747);
nand U27180 (N_27180,N_26871,N_26958);
xor U27181 (N_27181,N_26719,N_26718);
and U27182 (N_27182,N_26857,N_26975);
xnor U27183 (N_27183,N_26900,N_26825);
xor U27184 (N_27184,N_26743,N_26776);
nor U27185 (N_27185,N_26713,N_26986);
and U27186 (N_27186,N_26990,N_26863);
or U27187 (N_27187,N_26703,N_26731);
or U27188 (N_27188,N_26704,N_26978);
nand U27189 (N_27189,N_26964,N_26998);
xnor U27190 (N_27190,N_26967,N_26837);
and U27191 (N_27191,N_26712,N_26819);
nand U27192 (N_27192,N_26923,N_26912);
and U27193 (N_27193,N_26753,N_26949);
or U27194 (N_27194,N_26879,N_26854);
nor U27195 (N_27195,N_26747,N_26724);
nor U27196 (N_27196,N_26921,N_26820);
and U27197 (N_27197,N_26845,N_26744);
or U27198 (N_27198,N_26792,N_26991);
nand U27199 (N_27199,N_26912,N_26949);
nand U27200 (N_27200,N_26721,N_26775);
xnor U27201 (N_27201,N_26836,N_26971);
or U27202 (N_27202,N_26781,N_26958);
xnor U27203 (N_27203,N_26781,N_26732);
or U27204 (N_27204,N_26932,N_26934);
xor U27205 (N_27205,N_26751,N_26768);
nor U27206 (N_27206,N_26882,N_26822);
and U27207 (N_27207,N_26758,N_26969);
or U27208 (N_27208,N_26733,N_26994);
or U27209 (N_27209,N_26873,N_26983);
xor U27210 (N_27210,N_26805,N_26912);
or U27211 (N_27211,N_26903,N_26706);
and U27212 (N_27212,N_26867,N_26823);
xnor U27213 (N_27213,N_26978,N_26902);
or U27214 (N_27214,N_26758,N_26810);
and U27215 (N_27215,N_26794,N_26986);
nand U27216 (N_27216,N_26848,N_26928);
nor U27217 (N_27217,N_26757,N_26781);
xnor U27218 (N_27218,N_26931,N_26726);
and U27219 (N_27219,N_26702,N_26733);
nor U27220 (N_27220,N_26774,N_26894);
and U27221 (N_27221,N_26703,N_26997);
nor U27222 (N_27222,N_26773,N_26931);
and U27223 (N_27223,N_26991,N_26926);
nand U27224 (N_27224,N_26918,N_26966);
nand U27225 (N_27225,N_26713,N_26962);
xnor U27226 (N_27226,N_26761,N_26944);
nor U27227 (N_27227,N_26817,N_26869);
and U27228 (N_27228,N_26924,N_26803);
nand U27229 (N_27229,N_26773,N_26782);
and U27230 (N_27230,N_26964,N_26811);
and U27231 (N_27231,N_26794,N_26885);
nand U27232 (N_27232,N_26783,N_26896);
or U27233 (N_27233,N_26726,N_26911);
xor U27234 (N_27234,N_26942,N_26956);
or U27235 (N_27235,N_26878,N_26735);
and U27236 (N_27236,N_26826,N_26760);
nand U27237 (N_27237,N_26743,N_26943);
xor U27238 (N_27238,N_26802,N_26948);
nor U27239 (N_27239,N_26968,N_26967);
or U27240 (N_27240,N_26894,N_26929);
and U27241 (N_27241,N_26772,N_26785);
or U27242 (N_27242,N_26711,N_26948);
or U27243 (N_27243,N_26876,N_26992);
nor U27244 (N_27244,N_26742,N_26856);
and U27245 (N_27245,N_26765,N_26758);
and U27246 (N_27246,N_26900,N_26774);
or U27247 (N_27247,N_26795,N_26820);
or U27248 (N_27248,N_26852,N_26986);
xor U27249 (N_27249,N_26883,N_26889);
nor U27250 (N_27250,N_26854,N_26981);
xor U27251 (N_27251,N_26865,N_26893);
nor U27252 (N_27252,N_26729,N_26801);
xor U27253 (N_27253,N_26982,N_26809);
nand U27254 (N_27254,N_26806,N_26787);
and U27255 (N_27255,N_26978,N_26864);
nor U27256 (N_27256,N_26717,N_26849);
nor U27257 (N_27257,N_26776,N_26786);
nand U27258 (N_27258,N_26794,N_26841);
or U27259 (N_27259,N_26910,N_26937);
nand U27260 (N_27260,N_26943,N_26824);
and U27261 (N_27261,N_26871,N_26746);
or U27262 (N_27262,N_26764,N_26779);
xnor U27263 (N_27263,N_26817,N_26804);
nor U27264 (N_27264,N_26930,N_26836);
nand U27265 (N_27265,N_26852,N_26988);
or U27266 (N_27266,N_26816,N_26947);
nor U27267 (N_27267,N_26754,N_26838);
nor U27268 (N_27268,N_26928,N_26929);
nor U27269 (N_27269,N_26900,N_26811);
xor U27270 (N_27270,N_26736,N_26725);
nor U27271 (N_27271,N_26892,N_26987);
and U27272 (N_27272,N_26930,N_26989);
nand U27273 (N_27273,N_26973,N_26999);
nand U27274 (N_27274,N_26921,N_26940);
or U27275 (N_27275,N_26894,N_26920);
and U27276 (N_27276,N_26842,N_26933);
nor U27277 (N_27277,N_26765,N_26950);
nor U27278 (N_27278,N_26744,N_26906);
or U27279 (N_27279,N_26996,N_26902);
nor U27280 (N_27280,N_26803,N_26765);
xor U27281 (N_27281,N_26767,N_26993);
nand U27282 (N_27282,N_26706,N_26913);
or U27283 (N_27283,N_26735,N_26807);
or U27284 (N_27284,N_26777,N_26993);
nand U27285 (N_27285,N_26966,N_26861);
nor U27286 (N_27286,N_26832,N_26990);
or U27287 (N_27287,N_26972,N_26768);
nand U27288 (N_27288,N_26951,N_26834);
nand U27289 (N_27289,N_26712,N_26953);
and U27290 (N_27290,N_26919,N_26750);
nand U27291 (N_27291,N_26749,N_26836);
nor U27292 (N_27292,N_26776,N_26775);
or U27293 (N_27293,N_26847,N_26925);
or U27294 (N_27294,N_26753,N_26767);
xnor U27295 (N_27295,N_26773,N_26924);
xnor U27296 (N_27296,N_26818,N_26829);
or U27297 (N_27297,N_26858,N_26724);
nor U27298 (N_27298,N_26755,N_26865);
or U27299 (N_27299,N_26731,N_26863);
nor U27300 (N_27300,N_27094,N_27059);
nand U27301 (N_27301,N_27234,N_27281);
nor U27302 (N_27302,N_27152,N_27247);
and U27303 (N_27303,N_27033,N_27040);
nand U27304 (N_27304,N_27085,N_27295);
nand U27305 (N_27305,N_27170,N_27187);
and U27306 (N_27306,N_27294,N_27105);
nand U27307 (N_27307,N_27007,N_27060);
or U27308 (N_27308,N_27173,N_27006);
nand U27309 (N_27309,N_27136,N_27038);
nor U27310 (N_27310,N_27264,N_27076);
nor U27311 (N_27311,N_27122,N_27071);
xor U27312 (N_27312,N_27270,N_27055);
nand U27313 (N_27313,N_27080,N_27192);
nand U27314 (N_27314,N_27057,N_27127);
xor U27315 (N_27315,N_27074,N_27256);
xor U27316 (N_27316,N_27140,N_27248);
nand U27317 (N_27317,N_27068,N_27037);
and U27318 (N_27318,N_27276,N_27265);
nor U27319 (N_27319,N_27114,N_27117);
and U27320 (N_27320,N_27126,N_27023);
and U27321 (N_27321,N_27175,N_27253);
nor U27322 (N_27322,N_27069,N_27027);
xnor U27323 (N_27323,N_27290,N_27277);
nand U27324 (N_27324,N_27077,N_27049);
nand U27325 (N_27325,N_27082,N_27211);
xnor U27326 (N_27326,N_27092,N_27054);
or U27327 (N_27327,N_27284,N_27153);
xor U27328 (N_27328,N_27031,N_27177);
nand U27329 (N_27329,N_27016,N_27106);
nor U27330 (N_27330,N_27017,N_27018);
nor U27331 (N_27331,N_27202,N_27228);
nor U27332 (N_27332,N_27204,N_27189);
xnor U27333 (N_27333,N_27195,N_27024);
or U27334 (N_27334,N_27095,N_27123);
xnor U27335 (N_27335,N_27199,N_27169);
xnor U27336 (N_27336,N_27112,N_27081);
nor U27337 (N_27337,N_27252,N_27121);
nor U27338 (N_27338,N_27010,N_27046);
nand U27339 (N_27339,N_27050,N_27083);
and U27340 (N_27340,N_27188,N_27184);
or U27341 (N_27341,N_27125,N_27233);
nor U27342 (N_27342,N_27174,N_27014);
nor U27343 (N_27343,N_27020,N_27269);
nand U27344 (N_27344,N_27097,N_27251);
xor U27345 (N_27345,N_27065,N_27198);
nor U27346 (N_27346,N_27282,N_27047);
xnor U27347 (N_27347,N_27259,N_27229);
nand U27348 (N_27348,N_27176,N_27021);
xnor U27349 (N_27349,N_27255,N_27186);
or U27350 (N_27350,N_27292,N_27289);
nor U27351 (N_27351,N_27171,N_27058);
nand U27352 (N_27352,N_27216,N_27206);
xor U27353 (N_27353,N_27182,N_27203);
and U27354 (N_27354,N_27181,N_27263);
nor U27355 (N_27355,N_27141,N_27053);
nor U27356 (N_27356,N_27146,N_27167);
and U27357 (N_27357,N_27242,N_27110);
nand U27358 (N_27358,N_27113,N_27096);
nor U27359 (N_27359,N_27185,N_27279);
nor U27360 (N_27360,N_27004,N_27222);
and U27361 (N_27361,N_27257,N_27147);
xnor U27362 (N_27362,N_27268,N_27145);
xor U27363 (N_27363,N_27226,N_27118);
and U27364 (N_27364,N_27267,N_27196);
xor U27365 (N_27365,N_27034,N_27197);
xnor U27366 (N_27366,N_27298,N_27039);
nor U27367 (N_27367,N_27030,N_27193);
nand U27368 (N_27368,N_27164,N_27012);
or U27369 (N_27369,N_27026,N_27142);
nand U27370 (N_27370,N_27154,N_27208);
nor U27371 (N_27371,N_27210,N_27029);
and U27372 (N_27372,N_27161,N_27091);
nand U27373 (N_27373,N_27078,N_27099);
nor U27374 (N_27374,N_27205,N_27201);
xnor U27375 (N_27375,N_27104,N_27019);
or U27376 (N_27376,N_27261,N_27166);
and U27377 (N_27377,N_27278,N_27093);
nand U27378 (N_27378,N_27235,N_27219);
or U27379 (N_27379,N_27108,N_27138);
and U27380 (N_27380,N_27134,N_27063);
nor U27381 (N_27381,N_27243,N_27254);
or U27382 (N_27382,N_27137,N_27089);
nand U27383 (N_27383,N_27086,N_27246);
and U27384 (N_27384,N_27200,N_27139);
xor U27385 (N_27385,N_27172,N_27266);
nor U27386 (N_27386,N_27035,N_27079);
and U27387 (N_27387,N_27143,N_27133);
nand U27388 (N_27388,N_27052,N_27214);
nand U27389 (N_27389,N_27045,N_27003);
nor U27390 (N_27390,N_27232,N_27191);
nand U27391 (N_27391,N_27013,N_27131);
and U27392 (N_27392,N_27245,N_27250);
nand U27393 (N_27393,N_27275,N_27107);
xnor U27394 (N_27394,N_27230,N_27215);
xnor U27395 (N_27395,N_27130,N_27075);
and U27396 (N_27396,N_27151,N_27036);
nand U27397 (N_27397,N_27119,N_27299);
nor U27398 (N_27398,N_27042,N_27044);
nand U27399 (N_27399,N_27217,N_27120);
nand U27400 (N_27400,N_27218,N_27001);
nor U27401 (N_27401,N_27209,N_27280);
and U27402 (N_27402,N_27238,N_27159);
nor U27403 (N_27403,N_27090,N_27148);
nand U27404 (N_27404,N_27150,N_27272);
nor U27405 (N_27405,N_27223,N_27240);
nor U27406 (N_27406,N_27260,N_27132);
or U27407 (N_27407,N_27098,N_27157);
and U27408 (N_27408,N_27072,N_27149);
nor U27409 (N_27409,N_27194,N_27244);
xor U27410 (N_27410,N_27015,N_27236);
or U27411 (N_27411,N_27051,N_27220);
xor U27412 (N_27412,N_27274,N_27032);
nand U27413 (N_27413,N_27178,N_27124);
and U27414 (N_27414,N_27022,N_27162);
and U27415 (N_27415,N_27158,N_27287);
and U27416 (N_27416,N_27064,N_27286);
nand U27417 (N_27417,N_27135,N_27258);
nor U27418 (N_27418,N_27009,N_27271);
or U27419 (N_27419,N_27283,N_27180);
and U27420 (N_27420,N_27115,N_27011);
xnor U27421 (N_27421,N_27102,N_27116);
and U27422 (N_27422,N_27297,N_27043);
or U27423 (N_27423,N_27103,N_27179);
xor U27424 (N_27424,N_27101,N_27084);
or U27425 (N_27425,N_27109,N_27025);
nand U27426 (N_27426,N_27156,N_27067);
nand U27427 (N_27427,N_27061,N_27183);
nor U27428 (N_27428,N_27100,N_27190);
or U27429 (N_27429,N_27227,N_27213);
or U27430 (N_27430,N_27088,N_27262);
and U27431 (N_27431,N_27212,N_27241);
xor U27432 (N_27432,N_27000,N_27066);
nor U27433 (N_27433,N_27207,N_27168);
nand U27434 (N_27434,N_27165,N_27041);
nor U27435 (N_27435,N_27249,N_27163);
xor U27436 (N_27436,N_27160,N_27073);
xnor U27437 (N_27437,N_27285,N_27062);
xor U27438 (N_27438,N_27239,N_27111);
or U27439 (N_27439,N_27056,N_27128);
nand U27440 (N_27440,N_27293,N_27002);
and U27441 (N_27441,N_27291,N_27005);
nand U27442 (N_27442,N_27070,N_27155);
or U27443 (N_27443,N_27224,N_27273);
xor U27444 (N_27444,N_27225,N_27048);
nor U27445 (N_27445,N_27221,N_27087);
or U27446 (N_27446,N_27288,N_27231);
or U27447 (N_27447,N_27144,N_27028);
or U27448 (N_27448,N_27237,N_27296);
or U27449 (N_27449,N_27008,N_27129);
and U27450 (N_27450,N_27032,N_27113);
nor U27451 (N_27451,N_27256,N_27197);
nand U27452 (N_27452,N_27051,N_27095);
nor U27453 (N_27453,N_27155,N_27078);
xnor U27454 (N_27454,N_27000,N_27268);
xnor U27455 (N_27455,N_27000,N_27197);
nand U27456 (N_27456,N_27083,N_27241);
xor U27457 (N_27457,N_27214,N_27228);
xnor U27458 (N_27458,N_27009,N_27229);
nand U27459 (N_27459,N_27203,N_27110);
xor U27460 (N_27460,N_27168,N_27291);
or U27461 (N_27461,N_27020,N_27006);
nor U27462 (N_27462,N_27208,N_27159);
nand U27463 (N_27463,N_27062,N_27086);
nand U27464 (N_27464,N_27012,N_27245);
and U27465 (N_27465,N_27260,N_27051);
and U27466 (N_27466,N_27193,N_27228);
nor U27467 (N_27467,N_27263,N_27106);
or U27468 (N_27468,N_27130,N_27013);
nand U27469 (N_27469,N_27186,N_27153);
nand U27470 (N_27470,N_27007,N_27018);
nor U27471 (N_27471,N_27079,N_27112);
nor U27472 (N_27472,N_27054,N_27286);
and U27473 (N_27473,N_27025,N_27104);
xnor U27474 (N_27474,N_27045,N_27061);
and U27475 (N_27475,N_27186,N_27168);
xnor U27476 (N_27476,N_27226,N_27289);
nor U27477 (N_27477,N_27008,N_27109);
xor U27478 (N_27478,N_27296,N_27131);
nor U27479 (N_27479,N_27198,N_27016);
xnor U27480 (N_27480,N_27015,N_27089);
or U27481 (N_27481,N_27149,N_27075);
and U27482 (N_27482,N_27176,N_27147);
or U27483 (N_27483,N_27101,N_27186);
xnor U27484 (N_27484,N_27135,N_27196);
xor U27485 (N_27485,N_27109,N_27056);
and U27486 (N_27486,N_27269,N_27073);
nor U27487 (N_27487,N_27068,N_27218);
or U27488 (N_27488,N_27107,N_27039);
nor U27489 (N_27489,N_27180,N_27177);
xnor U27490 (N_27490,N_27022,N_27119);
or U27491 (N_27491,N_27211,N_27083);
xnor U27492 (N_27492,N_27192,N_27111);
nor U27493 (N_27493,N_27142,N_27179);
nor U27494 (N_27494,N_27083,N_27058);
or U27495 (N_27495,N_27227,N_27277);
nor U27496 (N_27496,N_27097,N_27074);
xor U27497 (N_27497,N_27287,N_27242);
and U27498 (N_27498,N_27147,N_27130);
xnor U27499 (N_27499,N_27219,N_27212);
or U27500 (N_27500,N_27035,N_27117);
or U27501 (N_27501,N_27294,N_27217);
xnor U27502 (N_27502,N_27282,N_27070);
and U27503 (N_27503,N_27139,N_27266);
nor U27504 (N_27504,N_27052,N_27135);
and U27505 (N_27505,N_27182,N_27051);
nor U27506 (N_27506,N_27246,N_27259);
or U27507 (N_27507,N_27121,N_27164);
xor U27508 (N_27508,N_27230,N_27070);
or U27509 (N_27509,N_27138,N_27244);
xnor U27510 (N_27510,N_27267,N_27150);
xor U27511 (N_27511,N_27212,N_27151);
nand U27512 (N_27512,N_27004,N_27228);
nand U27513 (N_27513,N_27232,N_27285);
or U27514 (N_27514,N_27004,N_27029);
nand U27515 (N_27515,N_27144,N_27141);
xnor U27516 (N_27516,N_27281,N_27289);
and U27517 (N_27517,N_27046,N_27168);
xnor U27518 (N_27518,N_27105,N_27229);
and U27519 (N_27519,N_27266,N_27071);
nor U27520 (N_27520,N_27047,N_27064);
and U27521 (N_27521,N_27037,N_27263);
or U27522 (N_27522,N_27156,N_27109);
nor U27523 (N_27523,N_27138,N_27186);
or U27524 (N_27524,N_27236,N_27071);
nor U27525 (N_27525,N_27269,N_27192);
nor U27526 (N_27526,N_27065,N_27113);
nor U27527 (N_27527,N_27056,N_27255);
or U27528 (N_27528,N_27071,N_27173);
or U27529 (N_27529,N_27054,N_27124);
or U27530 (N_27530,N_27209,N_27163);
xor U27531 (N_27531,N_27278,N_27049);
and U27532 (N_27532,N_27244,N_27055);
xnor U27533 (N_27533,N_27252,N_27022);
nor U27534 (N_27534,N_27088,N_27175);
and U27535 (N_27535,N_27099,N_27032);
and U27536 (N_27536,N_27220,N_27027);
nor U27537 (N_27537,N_27193,N_27200);
nand U27538 (N_27538,N_27251,N_27129);
nor U27539 (N_27539,N_27196,N_27259);
xor U27540 (N_27540,N_27162,N_27223);
xor U27541 (N_27541,N_27284,N_27009);
nand U27542 (N_27542,N_27191,N_27153);
nor U27543 (N_27543,N_27199,N_27108);
and U27544 (N_27544,N_27289,N_27145);
and U27545 (N_27545,N_27298,N_27020);
or U27546 (N_27546,N_27160,N_27288);
or U27547 (N_27547,N_27212,N_27159);
and U27548 (N_27548,N_27191,N_27082);
nand U27549 (N_27549,N_27043,N_27030);
nor U27550 (N_27550,N_27208,N_27182);
or U27551 (N_27551,N_27266,N_27149);
and U27552 (N_27552,N_27087,N_27110);
and U27553 (N_27553,N_27037,N_27113);
and U27554 (N_27554,N_27080,N_27150);
nor U27555 (N_27555,N_27092,N_27299);
or U27556 (N_27556,N_27147,N_27161);
nor U27557 (N_27557,N_27122,N_27266);
xnor U27558 (N_27558,N_27202,N_27081);
and U27559 (N_27559,N_27246,N_27110);
xnor U27560 (N_27560,N_27285,N_27071);
xor U27561 (N_27561,N_27212,N_27235);
nand U27562 (N_27562,N_27254,N_27269);
xnor U27563 (N_27563,N_27039,N_27035);
and U27564 (N_27564,N_27249,N_27165);
nand U27565 (N_27565,N_27024,N_27292);
nor U27566 (N_27566,N_27184,N_27251);
or U27567 (N_27567,N_27080,N_27149);
nand U27568 (N_27568,N_27279,N_27002);
nand U27569 (N_27569,N_27159,N_27148);
and U27570 (N_27570,N_27282,N_27223);
nor U27571 (N_27571,N_27161,N_27110);
nand U27572 (N_27572,N_27067,N_27114);
or U27573 (N_27573,N_27100,N_27049);
and U27574 (N_27574,N_27292,N_27164);
nor U27575 (N_27575,N_27066,N_27255);
or U27576 (N_27576,N_27001,N_27125);
nand U27577 (N_27577,N_27048,N_27090);
xnor U27578 (N_27578,N_27141,N_27152);
nand U27579 (N_27579,N_27109,N_27114);
nand U27580 (N_27580,N_27071,N_27160);
nor U27581 (N_27581,N_27226,N_27252);
or U27582 (N_27582,N_27221,N_27157);
or U27583 (N_27583,N_27143,N_27238);
xor U27584 (N_27584,N_27221,N_27254);
xnor U27585 (N_27585,N_27101,N_27032);
and U27586 (N_27586,N_27100,N_27115);
nand U27587 (N_27587,N_27079,N_27191);
and U27588 (N_27588,N_27164,N_27074);
xnor U27589 (N_27589,N_27047,N_27100);
and U27590 (N_27590,N_27202,N_27014);
xor U27591 (N_27591,N_27299,N_27097);
xnor U27592 (N_27592,N_27012,N_27023);
nor U27593 (N_27593,N_27283,N_27155);
nand U27594 (N_27594,N_27254,N_27281);
xnor U27595 (N_27595,N_27181,N_27098);
nand U27596 (N_27596,N_27013,N_27180);
or U27597 (N_27597,N_27086,N_27031);
xnor U27598 (N_27598,N_27045,N_27225);
xor U27599 (N_27599,N_27024,N_27127);
or U27600 (N_27600,N_27591,N_27589);
xor U27601 (N_27601,N_27315,N_27458);
nor U27602 (N_27602,N_27433,N_27376);
nor U27603 (N_27603,N_27587,N_27511);
and U27604 (N_27604,N_27588,N_27412);
and U27605 (N_27605,N_27534,N_27408);
or U27606 (N_27606,N_27371,N_27465);
nor U27607 (N_27607,N_27528,N_27475);
xnor U27608 (N_27608,N_27393,N_27339);
nand U27609 (N_27609,N_27426,N_27554);
xnor U27610 (N_27610,N_27402,N_27468);
nor U27611 (N_27611,N_27449,N_27574);
or U27612 (N_27612,N_27301,N_27398);
xor U27613 (N_27613,N_27538,N_27300);
and U27614 (N_27614,N_27441,N_27355);
or U27615 (N_27615,N_27537,N_27503);
and U27616 (N_27616,N_27413,N_27362);
nor U27617 (N_27617,N_27377,N_27466);
nand U27618 (N_27618,N_27473,N_27430);
nor U27619 (N_27619,N_27566,N_27526);
and U27620 (N_27620,N_27508,N_27460);
or U27621 (N_27621,N_27354,N_27521);
or U27622 (N_27622,N_27437,N_27352);
or U27623 (N_27623,N_27399,N_27327);
nor U27624 (N_27624,N_27461,N_27389);
xor U27625 (N_27625,N_27310,N_27516);
or U27626 (N_27626,N_27386,N_27410);
xor U27627 (N_27627,N_27541,N_27559);
nand U27628 (N_27628,N_27557,N_27494);
nor U27629 (N_27629,N_27435,N_27498);
xor U27630 (N_27630,N_27328,N_27418);
nor U27631 (N_27631,N_27324,N_27406);
nand U27632 (N_27632,N_27302,N_27414);
nand U27633 (N_27633,N_27507,N_27488);
xor U27634 (N_27634,N_27467,N_27542);
nor U27635 (N_27635,N_27540,N_27431);
and U27636 (N_27636,N_27471,N_27490);
and U27637 (N_27637,N_27429,N_27489);
nand U27638 (N_27638,N_27423,N_27319);
or U27639 (N_27639,N_27351,N_27492);
or U27640 (N_27640,N_27580,N_27312);
nand U27641 (N_27641,N_27530,N_27479);
or U27642 (N_27642,N_27365,N_27305);
xnor U27643 (N_27643,N_27487,N_27350);
and U27644 (N_27644,N_27316,N_27575);
nand U27645 (N_27645,N_27384,N_27563);
xnor U27646 (N_27646,N_27546,N_27484);
nand U27647 (N_27647,N_27582,N_27560);
nand U27648 (N_27648,N_27367,N_27331);
xor U27649 (N_27649,N_27512,N_27445);
or U27650 (N_27650,N_27422,N_27564);
xor U27651 (N_27651,N_27486,N_27529);
xnor U27652 (N_27652,N_27405,N_27366);
and U27653 (N_27653,N_27364,N_27347);
nand U27654 (N_27654,N_27514,N_27353);
nor U27655 (N_27655,N_27522,N_27325);
xnor U27656 (N_27656,N_27556,N_27388);
or U27657 (N_27657,N_27450,N_27524);
or U27658 (N_27658,N_27535,N_27593);
nor U27659 (N_27659,N_27361,N_27455);
nand U27660 (N_27660,N_27439,N_27480);
and U27661 (N_27661,N_27572,N_27309);
nand U27662 (N_27662,N_27571,N_27539);
and U27663 (N_27663,N_27357,N_27320);
and U27664 (N_27664,N_27417,N_27520);
xor U27665 (N_27665,N_27323,N_27509);
nor U27666 (N_27666,N_27373,N_27493);
and U27667 (N_27667,N_27341,N_27579);
nor U27668 (N_27668,N_27532,N_27395);
and U27669 (N_27669,N_27573,N_27510);
or U27670 (N_27670,N_27337,N_27311);
xnor U27671 (N_27671,N_27472,N_27531);
and U27672 (N_27672,N_27330,N_27444);
xnor U27673 (N_27673,N_27419,N_27329);
and U27674 (N_27674,N_27313,N_27491);
xor U27675 (N_27675,N_27519,N_27454);
nor U27676 (N_27676,N_27442,N_27533);
xor U27677 (N_27677,N_27499,N_27436);
or U27678 (N_27678,N_27322,N_27482);
and U27679 (N_27679,N_27504,N_27334);
nor U27680 (N_27680,N_27427,N_27581);
xnor U27681 (N_27681,N_27432,N_27382);
nand U27682 (N_27682,N_27396,N_27409);
and U27683 (N_27683,N_27375,N_27415);
xnor U27684 (N_27684,N_27567,N_27505);
and U27685 (N_27685,N_27372,N_27391);
nor U27686 (N_27686,N_27363,N_27565);
nor U27687 (N_27687,N_27333,N_27321);
or U27688 (N_27688,N_27558,N_27477);
and U27689 (N_27689,N_27578,N_27304);
nor U27690 (N_27690,N_27407,N_27478);
or U27691 (N_27691,N_27378,N_27336);
nand U27692 (N_27692,N_27576,N_27545);
nor U27693 (N_27693,N_27446,N_27344);
and U27694 (N_27694,N_27317,N_27544);
and U27695 (N_27695,N_27392,N_27451);
or U27696 (N_27696,N_27411,N_27595);
nand U27697 (N_27697,N_27335,N_27561);
or U27698 (N_27698,N_27424,N_27463);
nand U27699 (N_27699,N_27585,N_27456);
nand U27700 (N_27700,N_27551,N_27577);
or U27701 (N_27701,N_27549,N_27469);
or U27702 (N_27702,N_27345,N_27448);
xnor U27703 (N_27703,N_27440,N_27387);
nor U27704 (N_27704,N_27497,N_27379);
xor U27705 (N_27705,N_27599,N_27525);
or U27706 (N_27706,N_27552,N_27425);
xor U27707 (N_27707,N_27598,N_27584);
nand U27708 (N_27708,N_27453,N_27555);
nand U27709 (N_27709,N_27416,N_27306);
nand U27710 (N_27710,N_27326,N_27483);
and U27711 (N_27711,N_27459,N_27346);
nand U27712 (N_27712,N_27536,N_27586);
nor U27713 (N_27713,N_27338,N_27421);
nand U27714 (N_27714,N_27447,N_27308);
nand U27715 (N_27715,N_27369,N_27506);
nor U27716 (N_27716,N_27348,N_27597);
or U27717 (N_27717,N_27462,N_27527);
xor U27718 (N_27718,N_27457,N_27358);
and U27719 (N_27719,N_27548,N_27394);
and U27720 (N_27720,N_27403,N_27370);
nor U27721 (N_27721,N_27502,N_27594);
or U27722 (N_27722,N_27428,N_27332);
and U27723 (N_27723,N_27474,N_27340);
xor U27724 (N_27724,N_27314,N_27356);
xnor U27725 (N_27725,N_27553,N_27464);
or U27726 (N_27726,N_27523,N_27481);
xor U27727 (N_27727,N_27596,N_27381);
or U27728 (N_27728,N_27496,N_27400);
nor U27729 (N_27729,N_27443,N_27349);
xor U27730 (N_27730,N_27303,N_27390);
nand U27731 (N_27731,N_27495,N_27360);
nor U27732 (N_27732,N_27383,N_27374);
xnor U27733 (N_27733,N_27385,N_27452);
or U27734 (N_27734,N_27401,N_27515);
xor U27735 (N_27735,N_27517,N_27501);
and U27736 (N_27736,N_27420,N_27434);
xnor U27737 (N_27737,N_27318,N_27476);
or U27738 (N_27738,N_27543,N_27380);
xnor U27739 (N_27739,N_27485,N_27359);
and U27740 (N_27740,N_27397,N_27562);
nand U27741 (N_27741,N_27438,N_27568);
or U27742 (N_27742,N_27570,N_27550);
xor U27743 (N_27743,N_27547,N_27569);
nand U27744 (N_27744,N_27583,N_27592);
xnor U27745 (N_27745,N_27368,N_27470);
and U27746 (N_27746,N_27404,N_27342);
xor U27747 (N_27747,N_27343,N_27307);
or U27748 (N_27748,N_27513,N_27500);
or U27749 (N_27749,N_27590,N_27518);
nand U27750 (N_27750,N_27370,N_27318);
nand U27751 (N_27751,N_27467,N_27396);
nor U27752 (N_27752,N_27578,N_27400);
xnor U27753 (N_27753,N_27457,N_27520);
xor U27754 (N_27754,N_27393,N_27446);
and U27755 (N_27755,N_27500,N_27330);
nand U27756 (N_27756,N_27506,N_27376);
or U27757 (N_27757,N_27573,N_27367);
nand U27758 (N_27758,N_27574,N_27370);
and U27759 (N_27759,N_27513,N_27305);
nor U27760 (N_27760,N_27462,N_27312);
xor U27761 (N_27761,N_27364,N_27307);
and U27762 (N_27762,N_27343,N_27326);
and U27763 (N_27763,N_27494,N_27548);
xnor U27764 (N_27764,N_27534,N_27562);
or U27765 (N_27765,N_27373,N_27581);
nand U27766 (N_27766,N_27533,N_27335);
and U27767 (N_27767,N_27497,N_27397);
and U27768 (N_27768,N_27328,N_27535);
xor U27769 (N_27769,N_27494,N_27430);
nor U27770 (N_27770,N_27599,N_27566);
nor U27771 (N_27771,N_27578,N_27444);
or U27772 (N_27772,N_27488,N_27585);
or U27773 (N_27773,N_27521,N_27497);
and U27774 (N_27774,N_27543,N_27578);
nand U27775 (N_27775,N_27594,N_27496);
xor U27776 (N_27776,N_27529,N_27565);
or U27777 (N_27777,N_27573,N_27421);
nand U27778 (N_27778,N_27426,N_27568);
nand U27779 (N_27779,N_27583,N_27420);
or U27780 (N_27780,N_27461,N_27480);
xor U27781 (N_27781,N_27587,N_27585);
or U27782 (N_27782,N_27310,N_27417);
xnor U27783 (N_27783,N_27563,N_27426);
nor U27784 (N_27784,N_27428,N_27441);
and U27785 (N_27785,N_27580,N_27506);
xnor U27786 (N_27786,N_27399,N_27344);
and U27787 (N_27787,N_27591,N_27515);
xnor U27788 (N_27788,N_27373,N_27466);
or U27789 (N_27789,N_27597,N_27391);
and U27790 (N_27790,N_27350,N_27390);
or U27791 (N_27791,N_27364,N_27542);
nand U27792 (N_27792,N_27454,N_27387);
nand U27793 (N_27793,N_27426,N_27475);
and U27794 (N_27794,N_27493,N_27584);
nor U27795 (N_27795,N_27311,N_27408);
xor U27796 (N_27796,N_27307,N_27377);
or U27797 (N_27797,N_27561,N_27592);
or U27798 (N_27798,N_27546,N_27464);
nor U27799 (N_27799,N_27573,N_27490);
nor U27800 (N_27800,N_27570,N_27502);
xor U27801 (N_27801,N_27488,N_27451);
or U27802 (N_27802,N_27365,N_27381);
xor U27803 (N_27803,N_27406,N_27387);
nor U27804 (N_27804,N_27589,N_27312);
or U27805 (N_27805,N_27399,N_27547);
xnor U27806 (N_27806,N_27543,N_27523);
and U27807 (N_27807,N_27353,N_27535);
nor U27808 (N_27808,N_27575,N_27369);
nor U27809 (N_27809,N_27521,N_27372);
xor U27810 (N_27810,N_27359,N_27497);
and U27811 (N_27811,N_27336,N_27545);
and U27812 (N_27812,N_27340,N_27320);
or U27813 (N_27813,N_27421,N_27561);
nor U27814 (N_27814,N_27392,N_27334);
or U27815 (N_27815,N_27581,N_27587);
nor U27816 (N_27816,N_27462,N_27589);
nand U27817 (N_27817,N_27403,N_27558);
or U27818 (N_27818,N_27415,N_27417);
and U27819 (N_27819,N_27372,N_27397);
and U27820 (N_27820,N_27303,N_27476);
and U27821 (N_27821,N_27378,N_27430);
nand U27822 (N_27822,N_27317,N_27474);
nand U27823 (N_27823,N_27317,N_27326);
nor U27824 (N_27824,N_27586,N_27524);
nor U27825 (N_27825,N_27413,N_27561);
and U27826 (N_27826,N_27389,N_27459);
and U27827 (N_27827,N_27359,N_27457);
xnor U27828 (N_27828,N_27306,N_27582);
nor U27829 (N_27829,N_27464,N_27420);
or U27830 (N_27830,N_27429,N_27534);
xnor U27831 (N_27831,N_27530,N_27470);
or U27832 (N_27832,N_27583,N_27314);
xnor U27833 (N_27833,N_27560,N_27546);
and U27834 (N_27834,N_27544,N_27369);
nor U27835 (N_27835,N_27547,N_27479);
and U27836 (N_27836,N_27589,N_27557);
nor U27837 (N_27837,N_27304,N_27510);
xnor U27838 (N_27838,N_27388,N_27305);
nor U27839 (N_27839,N_27578,N_27374);
and U27840 (N_27840,N_27327,N_27564);
and U27841 (N_27841,N_27479,N_27525);
nand U27842 (N_27842,N_27406,N_27557);
and U27843 (N_27843,N_27515,N_27442);
xnor U27844 (N_27844,N_27412,N_27553);
nand U27845 (N_27845,N_27529,N_27547);
nand U27846 (N_27846,N_27494,N_27329);
or U27847 (N_27847,N_27318,N_27423);
nor U27848 (N_27848,N_27324,N_27530);
xnor U27849 (N_27849,N_27470,N_27465);
xor U27850 (N_27850,N_27447,N_27415);
xnor U27851 (N_27851,N_27448,N_27581);
and U27852 (N_27852,N_27465,N_27360);
or U27853 (N_27853,N_27527,N_27383);
nor U27854 (N_27854,N_27533,N_27515);
or U27855 (N_27855,N_27459,N_27419);
or U27856 (N_27856,N_27437,N_27409);
and U27857 (N_27857,N_27462,N_27339);
and U27858 (N_27858,N_27389,N_27574);
xor U27859 (N_27859,N_27542,N_27533);
or U27860 (N_27860,N_27504,N_27353);
nor U27861 (N_27861,N_27444,N_27583);
xor U27862 (N_27862,N_27351,N_27553);
or U27863 (N_27863,N_27523,N_27310);
nor U27864 (N_27864,N_27316,N_27514);
or U27865 (N_27865,N_27571,N_27372);
nor U27866 (N_27866,N_27343,N_27563);
xnor U27867 (N_27867,N_27433,N_27362);
or U27868 (N_27868,N_27315,N_27335);
and U27869 (N_27869,N_27357,N_27381);
nand U27870 (N_27870,N_27357,N_27378);
and U27871 (N_27871,N_27371,N_27341);
or U27872 (N_27872,N_27589,N_27317);
xor U27873 (N_27873,N_27322,N_27384);
or U27874 (N_27874,N_27462,N_27457);
xor U27875 (N_27875,N_27573,N_27426);
xor U27876 (N_27876,N_27371,N_27478);
and U27877 (N_27877,N_27481,N_27446);
and U27878 (N_27878,N_27582,N_27371);
xnor U27879 (N_27879,N_27366,N_27427);
nand U27880 (N_27880,N_27591,N_27576);
nor U27881 (N_27881,N_27313,N_27544);
nor U27882 (N_27882,N_27355,N_27566);
nand U27883 (N_27883,N_27483,N_27593);
nand U27884 (N_27884,N_27529,N_27533);
nor U27885 (N_27885,N_27595,N_27441);
nand U27886 (N_27886,N_27314,N_27315);
nand U27887 (N_27887,N_27522,N_27486);
xor U27888 (N_27888,N_27402,N_27517);
nor U27889 (N_27889,N_27338,N_27320);
and U27890 (N_27890,N_27306,N_27362);
or U27891 (N_27891,N_27575,N_27435);
nand U27892 (N_27892,N_27597,N_27408);
xor U27893 (N_27893,N_27337,N_27548);
nor U27894 (N_27894,N_27475,N_27581);
nor U27895 (N_27895,N_27472,N_27504);
nand U27896 (N_27896,N_27305,N_27543);
and U27897 (N_27897,N_27362,N_27313);
xnor U27898 (N_27898,N_27344,N_27530);
or U27899 (N_27899,N_27470,N_27418);
nand U27900 (N_27900,N_27781,N_27870);
xnor U27901 (N_27901,N_27701,N_27688);
nand U27902 (N_27902,N_27761,N_27643);
xor U27903 (N_27903,N_27635,N_27673);
xor U27904 (N_27904,N_27824,N_27841);
xnor U27905 (N_27905,N_27835,N_27763);
and U27906 (N_27906,N_27878,N_27850);
xnor U27907 (N_27907,N_27668,N_27745);
xor U27908 (N_27908,N_27788,N_27853);
nand U27909 (N_27909,N_27806,N_27722);
nor U27910 (N_27910,N_27672,N_27778);
xor U27911 (N_27911,N_27783,N_27713);
nor U27912 (N_27912,N_27621,N_27796);
or U27913 (N_27913,N_27691,N_27771);
and U27914 (N_27914,N_27830,N_27848);
xor U27915 (N_27915,N_27801,N_27708);
or U27916 (N_27916,N_27724,N_27653);
nor U27917 (N_27917,N_27802,N_27856);
xnor U27918 (N_27918,N_27782,N_27623);
and U27919 (N_27919,N_27604,N_27819);
and U27920 (N_27920,N_27727,N_27644);
nand U27921 (N_27921,N_27666,N_27662);
nor U27922 (N_27922,N_27756,N_27613);
and U27923 (N_27923,N_27891,N_27833);
or U27924 (N_27924,N_27669,N_27791);
xor U27925 (N_27925,N_27754,N_27732);
and U27926 (N_27926,N_27695,N_27849);
xnor U27927 (N_27927,N_27725,N_27839);
xnor U27928 (N_27928,N_27871,N_27785);
nor U27929 (N_27929,N_27620,N_27651);
xor U27930 (N_27930,N_27847,N_27881);
nand U27931 (N_27931,N_27731,N_27883);
nand U27932 (N_27932,N_27720,N_27654);
nand U27933 (N_27933,N_27652,N_27838);
nor U27934 (N_27934,N_27696,N_27612);
nor U27935 (N_27935,N_27834,N_27657);
xnor U27936 (N_27936,N_27705,N_27809);
and U27937 (N_27937,N_27775,N_27733);
nor U27938 (N_27938,N_27624,N_27893);
and U27939 (N_27939,N_27677,N_27712);
nand U27940 (N_27940,N_27715,N_27619);
nor U27941 (N_27941,N_27854,N_27752);
and U27942 (N_27942,N_27670,N_27676);
nor U27943 (N_27943,N_27884,N_27741);
nand U27944 (N_27944,N_27898,N_27719);
nor U27945 (N_27945,N_27642,N_27821);
nand U27946 (N_27946,N_27865,N_27875);
or U27947 (N_27947,N_27611,N_27879);
or U27948 (N_27948,N_27675,N_27660);
nor U27949 (N_27949,N_27664,N_27795);
nor U27950 (N_27950,N_27774,N_27681);
or U27951 (N_27951,N_27858,N_27707);
nand U27952 (N_27952,N_27726,N_27855);
xor U27953 (N_27953,N_27603,N_27790);
nor U27954 (N_27954,N_27646,N_27869);
nor U27955 (N_27955,N_27814,N_27810);
or U27956 (N_27956,N_27873,N_27617);
or U27957 (N_27957,N_27844,N_27818);
and U27958 (N_27958,N_27888,N_27805);
nand U27959 (N_27959,N_27812,N_27655);
nand U27960 (N_27960,N_27671,N_27689);
xnor U27961 (N_27961,N_27773,N_27697);
xnor U27962 (N_27962,N_27863,N_27736);
and U27963 (N_27963,N_27823,N_27700);
nand U27964 (N_27964,N_27784,N_27626);
and U27965 (N_27965,N_27717,N_27772);
or U27966 (N_27966,N_27886,N_27614);
nor U27967 (N_27967,N_27765,N_27827);
xor U27968 (N_27968,N_27792,N_27767);
or U27969 (N_27969,N_27716,N_27890);
and U27970 (N_27970,N_27851,N_27889);
or U27971 (N_27971,N_27740,N_27702);
xor U27972 (N_27972,N_27859,N_27641);
or U27973 (N_27973,N_27692,N_27721);
nand U27974 (N_27974,N_27777,N_27887);
nor U27975 (N_27975,N_27897,N_27825);
nand U27976 (N_27976,N_27629,N_27882);
nand U27977 (N_27977,N_27729,N_27768);
and U27978 (N_27978,N_27800,N_27780);
nand U27979 (N_27979,N_27822,N_27728);
nand U27980 (N_27980,N_27826,N_27816);
nand U27981 (N_27981,N_27694,N_27684);
nand U27982 (N_27982,N_27896,N_27658);
nand U27983 (N_27983,N_27811,N_27867);
and U27984 (N_27984,N_27638,N_27723);
or U27985 (N_27985,N_27757,N_27759);
and U27986 (N_27986,N_27633,N_27840);
nand U27987 (N_27987,N_27743,N_27747);
nand U27988 (N_27988,N_27742,N_27864);
xor U27989 (N_27989,N_27861,N_27832);
nor U27990 (N_27990,N_27685,N_27710);
xnor U27991 (N_27991,N_27665,N_27857);
nor U27992 (N_27992,N_27750,N_27899);
nor U27993 (N_27993,N_27607,N_27770);
or U27994 (N_27994,N_27845,N_27630);
xor U27995 (N_27995,N_27815,N_27711);
nand U27996 (N_27996,N_27866,N_27687);
nand U27997 (N_27997,N_27779,N_27628);
and U27998 (N_27998,N_27730,N_27753);
and U27999 (N_27999,N_27808,N_27735);
nand U28000 (N_28000,N_27714,N_27877);
xor U28001 (N_28001,N_27709,N_27659);
and U28002 (N_28002,N_27600,N_27804);
or U28003 (N_28003,N_27634,N_27766);
and U28004 (N_28004,N_27656,N_27895);
and U28005 (N_28005,N_27680,N_27699);
nor U28006 (N_28006,N_27648,N_27616);
or U28007 (N_28007,N_27606,N_27762);
nand U28008 (N_28008,N_27737,N_27706);
xor U28009 (N_28009,N_27609,N_27682);
xnor U28010 (N_28010,N_27748,N_27751);
xor U28011 (N_28011,N_27860,N_27894);
xnor U28012 (N_28012,N_27637,N_27787);
or U28013 (N_28013,N_27610,N_27837);
and U28014 (N_28014,N_27789,N_27836);
xnor U28015 (N_28015,N_27885,N_27813);
nand U28016 (N_28016,N_27661,N_27876);
nand U28017 (N_28017,N_27663,N_27797);
xnor U28018 (N_28018,N_27640,N_27718);
nor U28019 (N_28019,N_27880,N_27843);
xor U28020 (N_28020,N_27817,N_27686);
or U28021 (N_28021,N_27807,N_27868);
xor U28022 (N_28022,N_27639,N_27872);
nor U28023 (N_28023,N_27678,N_27829);
nand U28024 (N_28024,N_27622,N_27650);
nor U28025 (N_28025,N_27769,N_27862);
nor U28026 (N_28026,N_27679,N_27828);
nor U28027 (N_28027,N_27803,N_27793);
or U28028 (N_28028,N_27625,N_27704);
or U28029 (N_28029,N_27649,N_27794);
and U28030 (N_28030,N_27798,N_27601);
nand U28031 (N_28031,N_27647,N_27786);
and U28032 (N_28032,N_27674,N_27820);
or U28033 (N_28033,N_27636,N_27605);
nor U28034 (N_28034,N_27739,N_27631);
or U28035 (N_28035,N_27618,N_27755);
xor U28036 (N_28036,N_27892,N_27690);
nand U28037 (N_28037,N_27738,N_27608);
nor U28038 (N_28038,N_27632,N_27683);
or U28039 (N_28039,N_27667,N_27746);
nor U28040 (N_28040,N_27760,N_27602);
and U28041 (N_28041,N_27627,N_27831);
or U28042 (N_28042,N_27749,N_27842);
nand U28043 (N_28043,N_27693,N_27874);
and U28044 (N_28044,N_27776,N_27615);
and U28045 (N_28045,N_27758,N_27734);
and U28046 (N_28046,N_27764,N_27799);
and U28047 (N_28047,N_27852,N_27744);
xor U28048 (N_28048,N_27703,N_27645);
and U28049 (N_28049,N_27698,N_27846);
and U28050 (N_28050,N_27845,N_27835);
nand U28051 (N_28051,N_27794,N_27808);
nor U28052 (N_28052,N_27669,N_27891);
nor U28053 (N_28053,N_27818,N_27757);
and U28054 (N_28054,N_27675,N_27843);
xnor U28055 (N_28055,N_27764,N_27700);
or U28056 (N_28056,N_27787,N_27816);
or U28057 (N_28057,N_27678,N_27689);
nor U28058 (N_28058,N_27771,N_27688);
and U28059 (N_28059,N_27638,N_27680);
or U28060 (N_28060,N_27874,N_27798);
or U28061 (N_28061,N_27605,N_27863);
or U28062 (N_28062,N_27714,N_27678);
and U28063 (N_28063,N_27728,N_27852);
nand U28064 (N_28064,N_27623,N_27707);
xor U28065 (N_28065,N_27850,N_27822);
and U28066 (N_28066,N_27880,N_27689);
or U28067 (N_28067,N_27844,N_27761);
xor U28068 (N_28068,N_27619,N_27695);
or U28069 (N_28069,N_27771,N_27753);
xor U28070 (N_28070,N_27659,N_27892);
and U28071 (N_28071,N_27623,N_27771);
nand U28072 (N_28072,N_27747,N_27885);
nor U28073 (N_28073,N_27863,N_27809);
xor U28074 (N_28074,N_27832,N_27764);
or U28075 (N_28075,N_27716,N_27641);
or U28076 (N_28076,N_27613,N_27662);
nor U28077 (N_28077,N_27725,N_27674);
or U28078 (N_28078,N_27864,N_27892);
xnor U28079 (N_28079,N_27871,N_27836);
nand U28080 (N_28080,N_27858,N_27788);
nor U28081 (N_28081,N_27773,N_27750);
xor U28082 (N_28082,N_27868,N_27797);
nand U28083 (N_28083,N_27718,N_27765);
and U28084 (N_28084,N_27709,N_27712);
and U28085 (N_28085,N_27807,N_27808);
nand U28086 (N_28086,N_27698,N_27616);
nor U28087 (N_28087,N_27675,N_27629);
nand U28088 (N_28088,N_27616,N_27822);
and U28089 (N_28089,N_27854,N_27707);
and U28090 (N_28090,N_27895,N_27799);
nand U28091 (N_28091,N_27605,N_27815);
xnor U28092 (N_28092,N_27763,N_27667);
and U28093 (N_28093,N_27845,N_27798);
and U28094 (N_28094,N_27756,N_27847);
xnor U28095 (N_28095,N_27725,N_27842);
nor U28096 (N_28096,N_27876,N_27875);
nand U28097 (N_28097,N_27767,N_27672);
xor U28098 (N_28098,N_27841,N_27779);
nor U28099 (N_28099,N_27801,N_27825);
and U28100 (N_28100,N_27851,N_27887);
xnor U28101 (N_28101,N_27699,N_27721);
nor U28102 (N_28102,N_27870,N_27775);
nor U28103 (N_28103,N_27875,N_27651);
xor U28104 (N_28104,N_27658,N_27789);
and U28105 (N_28105,N_27891,N_27787);
xnor U28106 (N_28106,N_27776,N_27740);
and U28107 (N_28107,N_27709,N_27775);
xnor U28108 (N_28108,N_27833,N_27679);
or U28109 (N_28109,N_27838,N_27628);
xor U28110 (N_28110,N_27897,N_27727);
xor U28111 (N_28111,N_27668,N_27672);
xor U28112 (N_28112,N_27853,N_27676);
and U28113 (N_28113,N_27798,N_27722);
nand U28114 (N_28114,N_27643,N_27776);
nand U28115 (N_28115,N_27825,N_27639);
or U28116 (N_28116,N_27746,N_27629);
or U28117 (N_28117,N_27869,N_27859);
nor U28118 (N_28118,N_27782,N_27635);
nor U28119 (N_28119,N_27882,N_27659);
xor U28120 (N_28120,N_27876,N_27894);
or U28121 (N_28121,N_27787,N_27814);
nand U28122 (N_28122,N_27698,N_27841);
xor U28123 (N_28123,N_27676,N_27784);
and U28124 (N_28124,N_27849,N_27876);
nor U28125 (N_28125,N_27680,N_27732);
nor U28126 (N_28126,N_27884,N_27620);
or U28127 (N_28127,N_27753,N_27635);
nor U28128 (N_28128,N_27609,N_27615);
or U28129 (N_28129,N_27897,N_27720);
nor U28130 (N_28130,N_27841,N_27850);
xor U28131 (N_28131,N_27729,N_27681);
and U28132 (N_28132,N_27882,N_27867);
or U28133 (N_28133,N_27702,N_27805);
xnor U28134 (N_28134,N_27645,N_27679);
or U28135 (N_28135,N_27764,N_27744);
xnor U28136 (N_28136,N_27676,N_27890);
nand U28137 (N_28137,N_27693,N_27824);
xor U28138 (N_28138,N_27815,N_27663);
nor U28139 (N_28139,N_27722,N_27648);
or U28140 (N_28140,N_27833,N_27613);
and U28141 (N_28141,N_27637,N_27706);
or U28142 (N_28142,N_27717,N_27710);
and U28143 (N_28143,N_27645,N_27807);
xor U28144 (N_28144,N_27868,N_27741);
or U28145 (N_28145,N_27717,N_27721);
and U28146 (N_28146,N_27815,N_27799);
xor U28147 (N_28147,N_27849,N_27642);
or U28148 (N_28148,N_27602,N_27813);
and U28149 (N_28149,N_27696,N_27634);
or U28150 (N_28150,N_27846,N_27605);
or U28151 (N_28151,N_27709,N_27667);
nand U28152 (N_28152,N_27782,N_27836);
or U28153 (N_28153,N_27705,N_27723);
nor U28154 (N_28154,N_27611,N_27692);
or U28155 (N_28155,N_27848,N_27757);
xor U28156 (N_28156,N_27664,N_27741);
nand U28157 (N_28157,N_27864,N_27670);
nor U28158 (N_28158,N_27821,N_27730);
or U28159 (N_28159,N_27877,N_27775);
and U28160 (N_28160,N_27667,N_27722);
xnor U28161 (N_28161,N_27770,N_27815);
nor U28162 (N_28162,N_27895,N_27750);
nand U28163 (N_28163,N_27660,N_27729);
and U28164 (N_28164,N_27718,N_27620);
xor U28165 (N_28165,N_27673,N_27757);
nand U28166 (N_28166,N_27677,N_27636);
xor U28167 (N_28167,N_27884,N_27817);
nor U28168 (N_28168,N_27680,N_27869);
xnor U28169 (N_28169,N_27847,N_27786);
or U28170 (N_28170,N_27781,N_27832);
or U28171 (N_28171,N_27871,N_27658);
or U28172 (N_28172,N_27765,N_27799);
xor U28173 (N_28173,N_27849,N_27791);
nand U28174 (N_28174,N_27639,N_27758);
or U28175 (N_28175,N_27631,N_27795);
nand U28176 (N_28176,N_27634,N_27764);
nor U28177 (N_28177,N_27750,N_27761);
and U28178 (N_28178,N_27669,N_27663);
and U28179 (N_28179,N_27864,N_27778);
nand U28180 (N_28180,N_27849,N_27808);
and U28181 (N_28181,N_27853,N_27777);
and U28182 (N_28182,N_27852,N_27771);
nand U28183 (N_28183,N_27784,N_27722);
nor U28184 (N_28184,N_27840,N_27834);
xnor U28185 (N_28185,N_27798,N_27833);
nor U28186 (N_28186,N_27876,N_27784);
nor U28187 (N_28187,N_27613,N_27634);
nand U28188 (N_28188,N_27826,N_27815);
or U28189 (N_28189,N_27759,N_27690);
nor U28190 (N_28190,N_27881,N_27813);
nor U28191 (N_28191,N_27746,N_27780);
or U28192 (N_28192,N_27605,N_27682);
and U28193 (N_28193,N_27691,N_27867);
nand U28194 (N_28194,N_27725,N_27792);
nor U28195 (N_28195,N_27835,N_27757);
or U28196 (N_28196,N_27845,N_27754);
nand U28197 (N_28197,N_27780,N_27733);
nor U28198 (N_28198,N_27741,N_27718);
or U28199 (N_28199,N_27830,N_27693);
nor U28200 (N_28200,N_27952,N_28027);
nand U28201 (N_28201,N_28025,N_28109);
nor U28202 (N_28202,N_28007,N_28023);
xor U28203 (N_28203,N_28028,N_28032);
or U28204 (N_28204,N_28014,N_27905);
and U28205 (N_28205,N_27901,N_28111);
xor U28206 (N_28206,N_28022,N_28103);
nand U28207 (N_28207,N_28038,N_27948);
nor U28208 (N_28208,N_27924,N_28070);
nand U28209 (N_28209,N_28015,N_28130);
or U28210 (N_28210,N_27959,N_28180);
nand U28211 (N_28211,N_28040,N_27983);
xnor U28212 (N_28212,N_28145,N_28066);
and U28213 (N_28213,N_28039,N_28123);
xor U28214 (N_28214,N_27975,N_27943);
nor U28215 (N_28215,N_27917,N_28030);
or U28216 (N_28216,N_28065,N_28047);
nand U28217 (N_28217,N_27945,N_28078);
and U28218 (N_28218,N_28165,N_27962);
nor U28219 (N_28219,N_27911,N_28019);
xnor U28220 (N_28220,N_28149,N_28160);
nor U28221 (N_28221,N_27978,N_27989);
nor U28222 (N_28222,N_28024,N_28035);
nor U28223 (N_28223,N_27906,N_27964);
and U28224 (N_28224,N_28068,N_27953);
nor U28225 (N_28225,N_28143,N_27907);
nand U28226 (N_28226,N_28094,N_27944);
nand U28227 (N_28227,N_28042,N_27908);
or U28228 (N_28228,N_28077,N_28079);
or U28229 (N_28229,N_27980,N_28091);
and U28230 (N_28230,N_28110,N_27995);
xor U28231 (N_28231,N_28080,N_28159);
xnor U28232 (N_28232,N_28041,N_28045);
and U28233 (N_28233,N_27925,N_28097);
or U28234 (N_28234,N_28146,N_28153);
nand U28235 (N_28235,N_27913,N_28193);
nor U28236 (N_28236,N_27984,N_28168);
and U28237 (N_28237,N_27967,N_28063);
nor U28238 (N_28238,N_27970,N_28029);
nor U28239 (N_28239,N_28190,N_28105);
and U28240 (N_28240,N_28088,N_27932);
nor U28241 (N_28241,N_28128,N_28085);
nand U28242 (N_28242,N_28102,N_28112);
nor U28243 (N_28243,N_28171,N_28107);
nor U28244 (N_28244,N_28004,N_28099);
nor U28245 (N_28245,N_28170,N_28185);
nor U28246 (N_28246,N_27926,N_27902);
nand U28247 (N_28247,N_28139,N_28134);
nand U28248 (N_28248,N_28126,N_28129);
or U28249 (N_28249,N_27957,N_27950);
or U28250 (N_28250,N_28184,N_28183);
nand U28251 (N_28251,N_27935,N_28148);
nand U28252 (N_28252,N_28158,N_27921);
or U28253 (N_28253,N_28064,N_27938);
nor U28254 (N_28254,N_28003,N_28167);
or U28255 (N_28255,N_28127,N_27992);
or U28256 (N_28256,N_28000,N_27934);
xnor U28257 (N_28257,N_28006,N_27949);
nor U28258 (N_28258,N_28072,N_28096);
and U28259 (N_28259,N_27955,N_28012);
or U28260 (N_28260,N_28187,N_27968);
and U28261 (N_28261,N_28192,N_27918);
and U28262 (N_28262,N_28002,N_27920);
or U28263 (N_28263,N_27903,N_28043);
xor U28264 (N_28264,N_28033,N_27993);
or U28265 (N_28265,N_28087,N_27928);
nand U28266 (N_28266,N_28073,N_28114);
and U28267 (N_28267,N_28131,N_28052);
nand U28268 (N_28268,N_28051,N_27933);
xnor U28269 (N_28269,N_28150,N_28074);
xor U28270 (N_28270,N_27974,N_28186);
nor U28271 (N_28271,N_28049,N_28095);
or U28272 (N_28272,N_28081,N_27971);
and U28273 (N_28273,N_28163,N_28198);
and U28274 (N_28274,N_28058,N_27936);
xor U28275 (N_28275,N_27998,N_28036);
and U28276 (N_28276,N_27991,N_28119);
nor U28277 (N_28277,N_28031,N_27958);
xnor U28278 (N_28278,N_27951,N_28141);
nand U28279 (N_28279,N_27900,N_28108);
or U28280 (N_28280,N_28116,N_27994);
nor U28281 (N_28281,N_28005,N_28197);
nand U28282 (N_28282,N_28071,N_28155);
or U28283 (N_28283,N_27966,N_28057);
xor U28284 (N_28284,N_28182,N_27904);
xnor U28285 (N_28285,N_28067,N_28164);
xor U28286 (N_28286,N_28194,N_27999);
or U28287 (N_28287,N_28137,N_27987);
nand U28288 (N_28288,N_28044,N_28083);
xor U28289 (N_28289,N_27946,N_28136);
nand U28290 (N_28290,N_28152,N_28021);
nand U28291 (N_28291,N_28177,N_28157);
and U28292 (N_28292,N_28001,N_27961);
and U28293 (N_28293,N_27963,N_28151);
or U28294 (N_28294,N_27915,N_28069);
and U28295 (N_28295,N_28196,N_27929);
nand U28296 (N_28296,N_28054,N_28018);
nand U28297 (N_28297,N_28037,N_28135);
xor U28298 (N_28298,N_27965,N_28181);
and U28299 (N_28299,N_28059,N_28173);
and U28300 (N_28300,N_28133,N_28162);
nand U28301 (N_28301,N_27954,N_27981);
or U28302 (N_28302,N_27912,N_27947);
and U28303 (N_28303,N_28060,N_28176);
xnor U28304 (N_28304,N_27990,N_28115);
xor U28305 (N_28305,N_28138,N_28104);
nor U28306 (N_28306,N_27914,N_27973);
and U28307 (N_28307,N_28161,N_27956);
and U28308 (N_28308,N_28156,N_28062);
xor U28309 (N_28309,N_28122,N_28199);
or U28310 (N_28310,N_28113,N_28172);
and U28311 (N_28311,N_27927,N_28098);
or U28312 (N_28312,N_28166,N_28120);
nor U28313 (N_28313,N_28092,N_28191);
and U28314 (N_28314,N_28169,N_28121);
or U28315 (N_28315,N_27996,N_28034);
nand U28316 (N_28316,N_28179,N_27982);
nand U28317 (N_28317,N_27969,N_27960);
nor U28318 (N_28318,N_27942,N_28125);
nand U28319 (N_28319,N_28011,N_28013);
nor U28320 (N_28320,N_27988,N_28178);
or U28321 (N_28321,N_27976,N_28140);
nand U28322 (N_28322,N_27977,N_27922);
and U28323 (N_28323,N_28106,N_27940);
nand U28324 (N_28324,N_27972,N_27939);
nand U28325 (N_28325,N_27997,N_28188);
and U28326 (N_28326,N_28147,N_27979);
or U28327 (N_28327,N_28053,N_28195);
and U28328 (N_28328,N_28086,N_28082);
and U28329 (N_28329,N_28089,N_28117);
nor U28330 (N_28330,N_27986,N_28189);
and U28331 (N_28331,N_27937,N_28061);
nand U28332 (N_28332,N_28076,N_28016);
nor U28333 (N_28333,N_28075,N_27909);
xor U28334 (N_28334,N_28010,N_28100);
and U28335 (N_28335,N_28084,N_28090);
and U28336 (N_28336,N_28118,N_27923);
xor U28337 (N_28337,N_28009,N_28056);
and U28338 (N_28338,N_28132,N_28017);
and U28339 (N_28339,N_27916,N_28055);
nand U28340 (N_28340,N_27985,N_27931);
nor U28341 (N_28341,N_28154,N_28093);
nor U28342 (N_28342,N_28124,N_28174);
nand U28343 (N_28343,N_28048,N_27941);
or U28344 (N_28344,N_27930,N_28050);
and U28345 (N_28345,N_27919,N_28142);
xor U28346 (N_28346,N_28026,N_28046);
or U28347 (N_28347,N_27910,N_28175);
xnor U28348 (N_28348,N_28101,N_28008);
and U28349 (N_28349,N_28144,N_28020);
or U28350 (N_28350,N_28146,N_27911);
and U28351 (N_28351,N_28063,N_27933);
and U28352 (N_28352,N_28003,N_27959);
and U28353 (N_28353,N_28026,N_28077);
or U28354 (N_28354,N_28074,N_28196);
or U28355 (N_28355,N_28169,N_27966);
xor U28356 (N_28356,N_27986,N_28195);
nor U28357 (N_28357,N_27921,N_27903);
nand U28358 (N_28358,N_28111,N_28050);
or U28359 (N_28359,N_28189,N_28139);
and U28360 (N_28360,N_28152,N_27970);
xnor U28361 (N_28361,N_28096,N_28008);
and U28362 (N_28362,N_28112,N_28190);
and U28363 (N_28363,N_28134,N_28152);
or U28364 (N_28364,N_27959,N_27915);
nand U28365 (N_28365,N_28080,N_28177);
and U28366 (N_28366,N_28067,N_28104);
nor U28367 (N_28367,N_28155,N_28046);
and U28368 (N_28368,N_27955,N_27947);
or U28369 (N_28369,N_28084,N_28103);
or U28370 (N_28370,N_28090,N_28065);
xnor U28371 (N_28371,N_28134,N_28176);
nor U28372 (N_28372,N_28101,N_28086);
or U28373 (N_28373,N_27935,N_28061);
nand U28374 (N_28374,N_27931,N_28179);
xnor U28375 (N_28375,N_27991,N_28018);
or U28376 (N_28376,N_28160,N_28084);
xnor U28377 (N_28377,N_27996,N_28036);
xor U28378 (N_28378,N_27984,N_28039);
and U28379 (N_28379,N_28118,N_27919);
nand U28380 (N_28380,N_28096,N_27913);
xnor U28381 (N_28381,N_28030,N_28042);
or U28382 (N_28382,N_28070,N_28182);
or U28383 (N_28383,N_28155,N_27976);
and U28384 (N_28384,N_28086,N_28105);
or U28385 (N_28385,N_27974,N_28150);
xor U28386 (N_28386,N_28181,N_28144);
nor U28387 (N_28387,N_27929,N_28098);
nand U28388 (N_28388,N_28075,N_27930);
or U28389 (N_28389,N_28162,N_28152);
xor U28390 (N_28390,N_28171,N_27987);
xnor U28391 (N_28391,N_27956,N_27969);
xor U28392 (N_28392,N_28184,N_28017);
xnor U28393 (N_28393,N_28054,N_27916);
nor U28394 (N_28394,N_27969,N_28160);
and U28395 (N_28395,N_28090,N_28119);
or U28396 (N_28396,N_28005,N_28088);
xor U28397 (N_28397,N_27917,N_28096);
nand U28398 (N_28398,N_27924,N_28129);
xnor U28399 (N_28399,N_28069,N_28084);
nand U28400 (N_28400,N_27922,N_28181);
xor U28401 (N_28401,N_28054,N_28181);
nor U28402 (N_28402,N_28078,N_28121);
nand U28403 (N_28403,N_28125,N_27907);
xor U28404 (N_28404,N_28016,N_28085);
or U28405 (N_28405,N_27931,N_28018);
nor U28406 (N_28406,N_28193,N_28187);
nor U28407 (N_28407,N_27916,N_28016);
xor U28408 (N_28408,N_28070,N_28023);
nor U28409 (N_28409,N_28036,N_27937);
or U28410 (N_28410,N_28097,N_28152);
xnor U28411 (N_28411,N_28122,N_27938);
or U28412 (N_28412,N_28060,N_27905);
xnor U28413 (N_28413,N_27985,N_28047);
nor U28414 (N_28414,N_27917,N_28018);
nor U28415 (N_28415,N_28060,N_27902);
nor U28416 (N_28416,N_28109,N_28194);
xnor U28417 (N_28417,N_27964,N_28128);
xor U28418 (N_28418,N_28187,N_28157);
and U28419 (N_28419,N_28186,N_28181);
and U28420 (N_28420,N_27936,N_27943);
or U28421 (N_28421,N_28000,N_28048);
nand U28422 (N_28422,N_28183,N_27935);
nand U28423 (N_28423,N_28069,N_27991);
xor U28424 (N_28424,N_28016,N_28130);
and U28425 (N_28425,N_28163,N_28030);
or U28426 (N_28426,N_28122,N_27995);
and U28427 (N_28427,N_27969,N_28104);
xnor U28428 (N_28428,N_28176,N_28064);
or U28429 (N_28429,N_28163,N_28194);
or U28430 (N_28430,N_28047,N_27900);
nor U28431 (N_28431,N_28039,N_28037);
xnor U28432 (N_28432,N_28140,N_27906);
nor U28433 (N_28433,N_28137,N_27969);
nand U28434 (N_28434,N_28016,N_27977);
and U28435 (N_28435,N_28009,N_28151);
nor U28436 (N_28436,N_27970,N_28052);
and U28437 (N_28437,N_27915,N_27981);
or U28438 (N_28438,N_27986,N_28127);
and U28439 (N_28439,N_27916,N_27997);
and U28440 (N_28440,N_27901,N_28150);
and U28441 (N_28441,N_28112,N_28040);
nand U28442 (N_28442,N_28133,N_28170);
nor U28443 (N_28443,N_28175,N_27976);
or U28444 (N_28444,N_27937,N_28180);
and U28445 (N_28445,N_27904,N_28107);
or U28446 (N_28446,N_28111,N_28064);
nor U28447 (N_28447,N_28182,N_28135);
nor U28448 (N_28448,N_28006,N_28192);
xor U28449 (N_28449,N_27928,N_28061);
nand U28450 (N_28450,N_28194,N_27903);
nand U28451 (N_28451,N_27907,N_27995);
xnor U28452 (N_28452,N_28138,N_27904);
or U28453 (N_28453,N_28028,N_28042);
nor U28454 (N_28454,N_27968,N_28071);
xor U28455 (N_28455,N_27953,N_28156);
and U28456 (N_28456,N_28029,N_28089);
nor U28457 (N_28457,N_28099,N_27956);
or U28458 (N_28458,N_28198,N_27976);
and U28459 (N_28459,N_28119,N_27913);
or U28460 (N_28460,N_28187,N_28185);
or U28461 (N_28461,N_28186,N_28183);
xor U28462 (N_28462,N_27903,N_28161);
and U28463 (N_28463,N_28168,N_28024);
nor U28464 (N_28464,N_27912,N_28052);
or U28465 (N_28465,N_28136,N_27966);
xor U28466 (N_28466,N_27927,N_28178);
xor U28467 (N_28467,N_28073,N_27964);
or U28468 (N_28468,N_28010,N_28189);
nor U28469 (N_28469,N_27908,N_28050);
or U28470 (N_28470,N_28058,N_27938);
nand U28471 (N_28471,N_27943,N_27988);
and U28472 (N_28472,N_27917,N_28054);
nand U28473 (N_28473,N_28171,N_28173);
or U28474 (N_28474,N_28059,N_28150);
or U28475 (N_28475,N_28104,N_27944);
or U28476 (N_28476,N_28182,N_28056);
and U28477 (N_28477,N_28146,N_27991);
nor U28478 (N_28478,N_28089,N_28077);
or U28479 (N_28479,N_28061,N_28020);
xnor U28480 (N_28480,N_28175,N_28131);
nor U28481 (N_28481,N_28147,N_27938);
and U28482 (N_28482,N_27915,N_27922);
or U28483 (N_28483,N_27908,N_28170);
and U28484 (N_28484,N_27932,N_28198);
nor U28485 (N_28485,N_27987,N_27919);
and U28486 (N_28486,N_28150,N_28012);
and U28487 (N_28487,N_28111,N_28140);
or U28488 (N_28488,N_28090,N_27978);
nor U28489 (N_28489,N_27902,N_28161);
and U28490 (N_28490,N_27963,N_28048);
and U28491 (N_28491,N_27919,N_27961);
or U28492 (N_28492,N_27926,N_28179);
nor U28493 (N_28493,N_28038,N_28124);
nor U28494 (N_28494,N_27921,N_28195);
nor U28495 (N_28495,N_28149,N_28012);
and U28496 (N_28496,N_28170,N_27902);
nor U28497 (N_28497,N_27903,N_28064);
nor U28498 (N_28498,N_28002,N_28144);
xnor U28499 (N_28499,N_28147,N_28120);
nand U28500 (N_28500,N_28432,N_28479);
xnor U28501 (N_28501,N_28212,N_28335);
or U28502 (N_28502,N_28390,N_28323);
and U28503 (N_28503,N_28333,N_28473);
xor U28504 (N_28504,N_28281,N_28382);
xnor U28505 (N_28505,N_28404,N_28318);
or U28506 (N_28506,N_28406,N_28225);
nand U28507 (N_28507,N_28283,N_28465);
and U28508 (N_28508,N_28210,N_28476);
xor U28509 (N_28509,N_28410,N_28280);
or U28510 (N_28510,N_28240,N_28299);
or U28511 (N_28511,N_28391,N_28327);
nand U28512 (N_28512,N_28450,N_28360);
and U28513 (N_28513,N_28493,N_28379);
xor U28514 (N_28514,N_28427,N_28289);
or U28515 (N_28515,N_28329,N_28262);
or U28516 (N_28516,N_28405,N_28436);
or U28517 (N_28517,N_28231,N_28317);
xnor U28518 (N_28518,N_28429,N_28492);
xor U28519 (N_28519,N_28264,N_28208);
or U28520 (N_28520,N_28319,N_28266);
and U28521 (N_28521,N_28467,N_28250);
or U28522 (N_28522,N_28246,N_28394);
nor U28523 (N_28523,N_28237,N_28292);
or U28524 (N_28524,N_28257,N_28336);
nor U28525 (N_28525,N_28373,N_28234);
xor U28526 (N_28526,N_28206,N_28337);
or U28527 (N_28527,N_28407,N_28412);
or U28528 (N_28528,N_28422,N_28290);
xnor U28529 (N_28529,N_28346,N_28236);
and U28530 (N_28530,N_28483,N_28277);
xnor U28531 (N_28531,N_28420,N_28453);
or U28532 (N_28532,N_28487,N_28307);
or U28533 (N_28533,N_28214,N_28330);
or U28534 (N_28534,N_28293,N_28460);
nand U28535 (N_28535,N_28204,N_28273);
and U28536 (N_28536,N_28238,N_28400);
or U28537 (N_28537,N_28315,N_28464);
or U28538 (N_28538,N_28279,N_28253);
xor U28539 (N_28539,N_28377,N_28261);
or U28540 (N_28540,N_28286,N_28217);
or U28541 (N_28541,N_28259,N_28452);
nor U28542 (N_28542,N_28345,N_28303);
xor U28543 (N_28543,N_28269,N_28369);
xnor U28544 (N_28544,N_28457,N_28439);
nand U28545 (N_28545,N_28472,N_28278);
and U28546 (N_28546,N_28320,N_28497);
xnor U28547 (N_28547,N_28362,N_28386);
nor U28548 (N_28548,N_28267,N_28252);
nor U28549 (N_28549,N_28351,N_28263);
and U28550 (N_28550,N_28301,N_28475);
nor U28551 (N_28551,N_28437,N_28489);
or U28552 (N_28552,N_28353,N_28372);
and U28553 (N_28553,N_28371,N_28341);
or U28554 (N_28554,N_28331,N_28496);
xor U28555 (N_28555,N_28350,N_28284);
xor U28556 (N_28556,N_28398,N_28477);
nand U28557 (N_28557,N_28348,N_28367);
or U28558 (N_28558,N_28478,N_28222);
and U28559 (N_28559,N_28241,N_28393);
or U28560 (N_28560,N_28224,N_28219);
or U28561 (N_28561,N_28349,N_28211);
xnor U28562 (N_28562,N_28430,N_28499);
xor U28563 (N_28563,N_28368,N_28326);
nor U28564 (N_28564,N_28365,N_28202);
and U28565 (N_28565,N_28215,N_28313);
xnor U28566 (N_28566,N_28358,N_28311);
nor U28567 (N_28567,N_28409,N_28359);
or U28568 (N_28568,N_28414,N_28232);
or U28569 (N_28569,N_28288,N_28426);
and U28570 (N_28570,N_28287,N_28374);
xor U28571 (N_28571,N_28469,N_28227);
or U28572 (N_28572,N_28399,N_28322);
nand U28573 (N_28573,N_28347,N_28271);
nor U28574 (N_28574,N_28383,N_28364);
xor U28575 (N_28575,N_28380,N_28291);
or U28576 (N_28576,N_28239,N_28396);
nor U28577 (N_28577,N_28375,N_28223);
or U28578 (N_28578,N_28471,N_28443);
and U28579 (N_28579,N_28352,N_28378);
or U28580 (N_28580,N_28235,N_28424);
and U28581 (N_28581,N_28421,N_28423);
and U28582 (N_28582,N_28242,N_28397);
nand U28583 (N_28583,N_28230,N_28446);
nor U28584 (N_28584,N_28310,N_28296);
and U28585 (N_28585,N_28454,N_28334);
nor U28586 (N_28586,N_28229,N_28248);
and U28587 (N_28587,N_28247,N_28300);
nor U28588 (N_28588,N_28495,N_28249);
nor U28589 (N_28589,N_28302,N_28415);
or U28590 (N_28590,N_28297,N_28314);
xnor U28591 (N_28591,N_28474,N_28440);
or U28592 (N_28592,N_28370,N_28306);
and U28593 (N_28593,N_28416,N_28468);
xnor U28594 (N_28594,N_28403,N_28265);
nand U28595 (N_28595,N_28305,N_28216);
or U28596 (N_28596,N_28482,N_28339);
xor U28597 (N_28597,N_28389,N_28402);
and U28598 (N_28598,N_28332,N_28419);
nand U28599 (N_28599,N_28376,N_28308);
xnor U28600 (N_28600,N_28254,N_28411);
xor U28601 (N_28601,N_28226,N_28243);
nor U28602 (N_28602,N_28295,N_28221);
xnor U28603 (N_28603,N_28498,N_28438);
nor U28604 (N_28604,N_28434,N_28385);
and U28605 (N_28605,N_28459,N_28228);
nor U28606 (N_28606,N_28325,N_28316);
nor U28607 (N_28607,N_28418,N_28340);
or U28608 (N_28608,N_28282,N_28260);
nand U28609 (N_28609,N_28285,N_28363);
nor U28610 (N_28610,N_28309,N_28491);
xor U28611 (N_28611,N_28494,N_28381);
nor U28612 (N_28612,N_28444,N_28251);
and U28613 (N_28613,N_28484,N_28490);
or U28614 (N_28614,N_28463,N_28481);
xor U28615 (N_28615,N_28449,N_28357);
nor U28616 (N_28616,N_28312,N_28205);
or U28617 (N_28617,N_28486,N_28244);
nand U28618 (N_28618,N_28321,N_28213);
and U28619 (N_28619,N_28387,N_28425);
nand U28620 (N_28620,N_28344,N_28388);
nand U28621 (N_28621,N_28220,N_28270);
or U28622 (N_28622,N_28445,N_28488);
and U28623 (N_28623,N_28200,N_28417);
nand U28624 (N_28624,N_28408,N_28354);
nand U28625 (N_28625,N_28442,N_28451);
and U28626 (N_28626,N_28461,N_28218);
nand U28627 (N_28627,N_28343,N_28361);
nor U28628 (N_28628,N_28274,N_28462);
nand U28629 (N_28629,N_28441,N_28392);
xor U28630 (N_28630,N_28276,N_28428);
nand U28631 (N_28631,N_28395,N_28455);
nand U28632 (N_28632,N_28431,N_28456);
and U28633 (N_28633,N_28401,N_28366);
nand U28634 (N_28634,N_28485,N_28324);
nor U28635 (N_28635,N_28245,N_28413);
nand U28636 (N_28636,N_28338,N_28470);
nor U28637 (N_28637,N_28304,N_28203);
and U28638 (N_28638,N_28272,N_28384);
or U28639 (N_28639,N_28233,N_28255);
or U28640 (N_28640,N_28356,N_28207);
or U28641 (N_28641,N_28342,N_28201);
xor U28642 (N_28642,N_28258,N_28458);
xor U28643 (N_28643,N_28268,N_28433);
nand U28644 (N_28644,N_28298,N_28466);
xor U28645 (N_28645,N_28328,N_28275);
and U28646 (N_28646,N_28256,N_28355);
nand U28647 (N_28647,N_28447,N_28209);
nand U28648 (N_28648,N_28435,N_28448);
and U28649 (N_28649,N_28294,N_28480);
or U28650 (N_28650,N_28315,N_28484);
nand U28651 (N_28651,N_28309,N_28341);
nor U28652 (N_28652,N_28312,N_28256);
nand U28653 (N_28653,N_28428,N_28483);
and U28654 (N_28654,N_28490,N_28315);
nor U28655 (N_28655,N_28448,N_28493);
nor U28656 (N_28656,N_28461,N_28387);
nand U28657 (N_28657,N_28378,N_28304);
xor U28658 (N_28658,N_28434,N_28245);
or U28659 (N_28659,N_28333,N_28339);
nand U28660 (N_28660,N_28248,N_28249);
nor U28661 (N_28661,N_28450,N_28406);
and U28662 (N_28662,N_28388,N_28296);
nand U28663 (N_28663,N_28326,N_28284);
nand U28664 (N_28664,N_28473,N_28489);
or U28665 (N_28665,N_28399,N_28482);
nor U28666 (N_28666,N_28225,N_28430);
nand U28667 (N_28667,N_28484,N_28408);
nand U28668 (N_28668,N_28237,N_28305);
xnor U28669 (N_28669,N_28251,N_28221);
and U28670 (N_28670,N_28242,N_28443);
xnor U28671 (N_28671,N_28217,N_28391);
xor U28672 (N_28672,N_28340,N_28262);
xnor U28673 (N_28673,N_28409,N_28287);
nand U28674 (N_28674,N_28258,N_28397);
and U28675 (N_28675,N_28299,N_28280);
and U28676 (N_28676,N_28357,N_28486);
or U28677 (N_28677,N_28206,N_28279);
nand U28678 (N_28678,N_28334,N_28330);
or U28679 (N_28679,N_28292,N_28475);
nand U28680 (N_28680,N_28300,N_28301);
xor U28681 (N_28681,N_28397,N_28408);
or U28682 (N_28682,N_28305,N_28272);
or U28683 (N_28683,N_28331,N_28440);
or U28684 (N_28684,N_28441,N_28318);
nor U28685 (N_28685,N_28280,N_28281);
nand U28686 (N_28686,N_28445,N_28271);
or U28687 (N_28687,N_28365,N_28314);
xor U28688 (N_28688,N_28346,N_28482);
nand U28689 (N_28689,N_28324,N_28398);
or U28690 (N_28690,N_28268,N_28320);
nor U28691 (N_28691,N_28394,N_28238);
and U28692 (N_28692,N_28222,N_28305);
xnor U28693 (N_28693,N_28207,N_28490);
xor U28694 (N_28694,N_28409,N_28310);
or U28695 (N_28695,N_28363,N_28256);
and U28696 (N_28696,N_28296,N_28280);
xnor U28697 (N_28697,N_28481,N_28430);
xnor U28698 (N_28698,N_28256,N_28373);
xor U28699 (N_28699,N_28489,N_28287);
or U28700 (N_28700,N_28382,N_28200);
nor U28701 (N_28701,N_28234,N_28316);
and U28702 (N_28702,N_28267,N_28362);
nor U28703 (N_28703,N_28333,N_28443);
xnor U28704 (N_28704,N_28218,N_28466);
and U28705 (N_28705,N_28303,N_28411);
xor U28706 (N_28706,N_28277,N_28403);
nand U28707 (N_28707,N_28329,N_28291);
nor U28708 (N_28708,N_28421,N_28262);
and U28709 (N_28709,N_28256,N_28220);
nor U28710 (N_28710,N_28342,N_28395);
or U28711 (N_28711,N_28474,N_28429);
nor U28712 (N_28712,N_28205,N_28411);
xnor U28713 (N_28713,N_28454,N_28491);
or U28714 (N_28714,N_28336,N_28397);
and U28715 (N_28715,N_28251,N_28377);
nand U28716 (N_28716,N_28304,N_28243);
or U28717 (N_28717,N_28238,N_28352);
and U28718 (N_28718,N_28225,N_28317);
and U28719 (N_28719,N_28239,N_28449);
and U28720 (N_28720,N_28283,N_28268);
and U28721 (N_28721,N_28268,N_28406);
or U28722 (N_28722,N_28356,N_28358);
or U28723 (N_28723,N_28201,N_28484);
nand U28724 (N_28724,N_28309,N_28213);
nand U28725 (N_28725,N_28490,N_28299);
and U28726 (N_28726,N_28393,N_28304);
xor U28727 (N_28727,N_28358,N_28350);
and U28728 (N_28728,N_28408,N_28347);
and U28729 (N_28729,N_28204,N_28360);
xnor U28730 (N_28730,N_28202,N_28430);
and U28731 (N_28731,N_28492,N_28461);
xnor U28732 (N_28732,N_28262,N_28367);
or U28733 (N_28733,N_28388,N_28241);
nand U28734 (N_28734,N_28296,N_28484);
or U28735 (N_28735,N_28262,N_28447);
nor U28736 (N_28736,N_28356,N_28216);
and U28737 (N_28737,N_28286,N_28309);
nand U28738 (N_28738,N_28294,N_28419);
or U28739 (N_28739,N_28223,N_28445);
xnor U28740 (N_28740,N_28249,N_28237);
and U28741 (N_28741,N_28454,N_28426);
and U28742 (N_28742,N_28224,N_28427);
or U28743 (N_28743,N_28478,N_28423);
nor U28744 (N_28744,N_28237,N_28200);
or U28745 (N_28745,N_28216,N_28467);
nor U28746 (N_28746,N_28339,N_28362);
or U28747 (N_28747,N_28302,N_28323);
and U28748 (N_28748,N_28261,N_28283);
and U28749 (N_28749,N_28334,N_28372);
and U28750 (N_28750,N_28307,N_28454);
and U28751 (N_28751,N_28391,N_28442);
or U28752 (N_28752,N_28206,N_28218);
nand U28753 (N_28753,N_28378,N_28450);
xnor U28754 (N_28754,N_28451,N_28343);
xor U28755 (N_28755,N_28412,N_28429);
nor U28756 (N_28756,N_28387,N_28337);
xor U28757 (N_28757,N_28397,N_28256);
nor U28758 (N_28758,N_28210,N_28300);
or U28759 (N_28759,N_28483,N_28367);
nand U28760 (N_28760,N_28494,N_28378);
nor U28761 (N_28761,N_28436,N_28469);
nand U28762 (N_28762,N_28306,N_28223);
and U28763 (N_28763,N_28450,N_28493);
and U28764 (N_28764,N_28436,N_28401);
or U28765 (N_28765,N_28401,N_28494);
xor U28766 (N_28766,N_28287,N_28248);
xor U28767 (N_28767,N_28412,N_28295);
nand U28768 (N_28768,N_28481,N_28312);
or U28769 (N_28769,N_28400,N_28473);
and U28770 (N_28770,N_28287,N_28251);
and U28771 (N_28771,N_28474,N_28491);
nor U28772 (N_28772,N_28422,N_28359);
and U28773 (N_28773,N_28442,N_28294);
xnor U28774 (N_28774,N_28231,N_28220);
xor U28775 (N_28775,N_28248,N_28237);
xor U28776 (N_28776,N_28212,N_28210);
xor U28777 (N_28777,N_28444,N_28322);
xor U28778 (N_28778,N_28267,N_28359);
xor U28779 (N_28779,N_28245,N_28341);
xnor U28780 (N_28780,N_28259,N_28329);
and U28781 (N_28781,N_28291,N_28341);
and U28782 (N_28782,N_28219,N_28485);
or U28783 (N_28783,N_28234,N_28278);
and U28784 (N_28784,N_28315,N_28252);
nor U28785 (N_28785,N_28238,N_28362);
xor U28786 (N_28786,N_28374,N_28323);
and U28787 (N_28787,N_28455,N_28414);
and U28788 (N_28788,N_28337,N_28324);
xnor U28789 (N_28789,N_28246,N_28368);
nor U28790 (N_28790,N_28234,N_28416);
and U28791 (N_28791,N_28317,N_28436);
nand U28792 (N_28792,N_28338,N_28239);
and U28793 (N_28793,N_28306,N_28488);
nand U28794 (N_28794,N_28388,N_28417);
nor U28795 (N_28795,N_28438,N_28415);
xor U28796 (N_28796,N_28280,N_28440);
or U28797 (N_28797,N_28297,N_28368);
and U28798 (N_28798,N_28271,N_28381);
and U28799 (N_28799,N_28464,N_28471);
xor U28800 (N_28800,N_28622,N_28545);
xor U28801 (N_28801,N_28778,N_28530);
and U28802 (N_28802,N_28548,N_28603);
and U28803 (N_28803,N_28678,N_28735);
nand U28804 (N_28804,N_28777,N_28713);
nor U28805 (N_28805,N_28514,N_28567);
and U28806 (N_28806,N_28590,N_28529);
or U28807 (N_28807,N_28652,N_28788);
nor U28808 (N_28808,N_28647,N_28748);
nand U28809 (N_28809,N_28554,N_28502);
and U28810 (N_28810,N_28673,N_28628);
or U28811 (N_28811,N_28779,N_28753);
nor U28812 (N_28812,N_28527,N_28614);
nor U28813 (N_28813,N_28761,N_28686);
or U28814 (N_28814,N_28704,N_28729);
and U28815 (N_28815,N_28575,N_28679);
xnor U28816 (N_28816,N_28602,N_28598);
nand U28817 (N_28817,N_28798,N_28608);
xor U28818 (N_28818,N_28595,N_28724);
and U28819 (N_28819,N_28773,N_28671);
xnor U28820 (N_28820,N_28692,N_28662);
and U28821 (N_28821,N_28523,N_28743);
xnor U28822 (N_28822,N_28585,N_28593);
nor U28823 (N_28823,N_28746,N_28645);
xnor U28824 (N_28824,N_28549,N_28659);
and U28825 (N_28825,N_28552,N_28584);
nor U28826 (N_28826,N_28640,N_28758);
nor U28827 (N_28827,N_28651,N_28543);
xor U28828 (N_28828,N_28555,N_28566);
and U28829 (N_28829,N_28714,N_28736);
xor U28830 (N_28830,N_28781,N_28635);
nand U28831 (N_28831,N_28701,N_28546);
nand U28832 (N_28832,N_28702,N_28630);
xor U28833 (N_28833,N_28790,N_28558);
and U28834 (N_28834,N_28741,N_28646);
and U28835 (N_28835,N_28601,N_28663);
xor U28836 (N_28836,N_28518,N_28520);
nand U28837 (N_28837,N_28634,N_28687);
xnor U28838 (N_28838,N_28670,N_28507);
xor U28839 (N_28839,N_28697,N_28793);
nand U28840 (N_28840,N_28577,N_28787);
and U28841 (N_28841,N_28740,N_28528);
and U28842 (N_28842,N_28755,N_28609);
and U28843 (N_28843,N_28587,N_28706);
and U28844 (N_28844,N_28572,N_28547);
or U28845 (N_28845,N_28606,N_28531);
nor U28846 (N_28846,N_28696,N_28565);
or U28847 (N_28847,N_28725,N_28750);
nor U28848 (N_28848,N_28654,N_28717);
and U28849 (N_28849,N_28756,N_28580);
or U28850 (N_28850,N_28629,N_28532);
or U28851 (N_28851,N_28541,N_28691);
and U28852 (N_28852,N_28737,N_28785);
or U28853 (N_28853,N_28642,N_28749);
nand U28854 (N_28854,N_28765,N_28672);
nor U28855 (N_28855,N_28666,N_28700);
and U28856 (N_28856,N_28684,N_28723);
nor U28857 (N_28857,N_28738,N_28711);
and U28858 (N_28858,N_28718,N_28557);
or U28859 (N_28859,N_28513,N_28762);
nor U28860 (N_28860,N_28660,N_28665);
or U28861 (N_28861,N_28551,N_28699);
nand U28862 (N_28862,N_28721,N_28703);
xnor U28863 (N_28863,N_28770,N_28739);
xnor U28864 (N_28864,N_28681,N_28568);
or U28865 (N_28865,N_28767,N_28742);
nor U28866 (N_28866,N_28669,N_28559);
nor U28867 (N_28867,N_28799,N_28538);
nand U28868 (N_28868,N_28553,N_28764);
xor U28869 (N_28869,N_28616,N_28540);
and U28870 (N_28870,N_28759,N_28641);
nor U28871 (N_28871,N_28727,N_28754);
and U28872 (N_28872,N_28607,N_28683);
and U28873 (N_28873,N_28775,N_28732);
or U28874 (N_28874,N_28535,N_28617);
or U28875 (N_28875,N_28690,N_28680);
or U28876 (N_28876,N_28644,N_28637);
nor U28877 (N_28877,N_28612,N_28534);
nand U28878 (N_28878,N_28772,N_28620);
nor U28879 (N_28879,N_28694,N_28632);
and U28880 (N_28880,N_28599,N_28618);
xor U28881 (N_28881,N_28658,N_28794);
nor U28882 (N_28882,N_28589,N_28720);
xnor U28883 (N_28883,N_28796,N_28615);
and U28884 (N_28884,N_28771,N_28763);
xnor U28885 (N_28885,N_28563,N_28578);
nand U28886 (N_28886,N_28581,N_28592);
nor U28887 (N_28887,N_28569,N_28560);
xor U28888 (N_28888,N_28537,N_28708);
xnor U28889 (N_28889,N_28521,N_28757);
and U28890 (N_28890,N_28769,N_28509);
or U28891 (N_28891,N_28733,N_28611);
xor U28892 (N_28892,N_28685,N_28657);
or U28893 (N_28893,N_28744,N_28522);
xnor U28894 (N_28894,N_28656,N_28621);
and U28895 (N_28895,N_28655,N_28536);
nand U28896 (N_28896,N_28613,N_28550);
and U28897 (N_28897,N_28639,N_28505);
nor U28898 (N_28898,N_28675,N_28719);
nor U28899 (N_28899,N_28517,N_28664);
nand U28900 (N_28900,N_28501,N_28582);
xor U28901 (N_28901,N_28605,N_28650);
and U28902 (N_28902,N_28734,N_28689);
xnor U28903 (N_28903,N_28712,N_28705);
or U28904 (N_28904,N_28722,N_28782);
nor U28905 (N_28905,N_28516,N_28574);
nand U28906 (N_28906,N_28631,N_28667);
xor U28907 (N_28907,N_28795,N_28648);
nand U28908 (N_28908,N_28676,N_28751);
nand U28909 (N_28909,N_28625,N_28682);
nor U28910 (N_28910,N_28564,N_28780);
xnor U28911 (N_28911,N_28627,N_28730);
nor U28912 (N_28912,N_28524,N_28544);
nor U28913 (N_28913,N_28789,N_28745);
xnor U28914 (N_28914,N_28797,N_28594);
nand U28915 (N_28915,N_28623,N_28500);
xnor U28916 (N_28916,N_28525,N_28556);
nand U28917 (N_28917,N_28512,N_28597);
xor U28918 (N_28918,N_28511,N_28503);
xnor U28919 (N_28919,N_28693,N_28573);
nand U28920 (N_28920,N_28508,N_28510);
and U28921 (N_28921,N_28731,N_28760);
xor U28922 (N_28922,N_28792,N_28583);
nor U28923 (N_28923,N_28636,N_28591);
and U28924 (N_28924,N_28728,N_28533);
and U28925 (N_28925,N_28783,N_28526);
and U28926 (N_28926,N_28698,N_28649);
nor U28927 (N_28927,N_28677,N_28576);
xor U28928 (N_28928,N_28643,N_28786);
nand U28929 (N_28929,N_28709,N_28716);
nand U28930 (N_28930,N_28776,N_28561);
and U28931 (N_28931,N_28726,N_28571);
nor U28932 (N_28932,N_28619,N_28715);
nand U28933 (N_28933,N_28504,N_28768);
nor U28934 (N_28934,N_28752,N_28707);
xor U28935 (N_28935,N_28633,N_28661);
nor U28936 (N_28936,N_28674,N_28610);
nor U28937 (N_28937,N_28586,N_28653);
and U28938 (N_28938,N_28791,N_28766);
or U28939 (N_28939,N_28539,N_28695);
and U28940 (N_28940,N_28668,N_28604);
nor U28941 (N_28941,N_28579,N_28638);
and U28942 (N_28942,N_28596,N_28626);
nor U28943 (N_28943,N_28519,N_28774);
and U28944 (N_28944,N_28688,N_28710);
nand U28945 (N_28945,N_28747,N_28784);
nand U28946 (N_28946,N_28624,N_28600);
nor U28947 (N_28947,N_28515,N_28588);
nor U28948 (N_28948,N_28570,N_28562);
nor U28949 (N_28949,N_28542,N_28506);
nand U28950 (N_28950,N_28697,N_28673);
and U28951 (N_28951,N_28670,N_28577);
or U28952 (N_28952,N_28641,N_28738);
or U28953 (N_28953,N_28508,N_28751);
nor U28954 (N_28954,N_28592,N_28562);
and U28955 (N_28955,N_28525,N_28631);
xnor U28956 (N_28956,N_28648,N_28684);
or U28957 (N_28957,N_28645,N_28798);
nor U28958 (N_28958,N_28601,N_28636);
xor U28959 (N_28959,N_28632,N_28582);
nand U28960 (N_28960,N_28671,N_28509);
nor U28961 (N_28961,N_28712,N_28754);
nor U28962 (N_28962,N_28670,N_28631);
xor U28963 (N_28963,N_28639,N_28588);
and U28964 (N_28964,N_28640,N_28614);
or U28965 (N_28965,N_28508,N_28585);
or U28966 (N_28966,N_28563,N_28733);
nand U28967 (N_28967,N_28615,N_28522);
or U28968 (N_28968,N_28778,N_28679);
and U28969 (N_28969,N_28708,N_28618);
or U28970 (N_28970,N_28783,N_28768);
nand U28971 (N_28971,N_28636,N_28681);
nand U28972 (N_28972,N_28509,N_28796);
or U28973 (N_28973,N_28732,N_28755);
and U28974 (N_28974,N_28588,N_28794);
nand U28975 (N_28975,N_28533,N_28657);
or U28976 (N_28976,N_28617,N_28587);
or U28977 (N_28977,N_28613,N_28542);
xor U28978 (N_28978,N_28587,N_28687);
nand U28979 (N_28979,N_28786,N_28515);
and U28980 (N_28980,N_28667,N_28650);
nor U28981 (N_28981,N_28714,N_28537);
and U28982 (N_28982,N_28512,N_28534);
nand U28983 (N_28983,N_28721,N_28706);
nor U28984 (N_28984,N_28684,N_28785);
nand U28985 (N_28985,N_28745,N_28626);
or U28986 (N_28986,N_28793,N_28629);
nand U28987 (N_28987,N_28679,N_28779);
and U28988 (N_28988,N_28719,N_28630);
or U28989 (N_28989,N_28589,N_28718);
and U28990 (N_28990,N_28715,N_28725);
or U28991 (N_28991,N_28514,N_28794);
xnor U28992 (N_28992,N_28719,N_28723);
xnor U28993 (N_28993,N_28761,N_28793);
nor U28994 (N_28994,N_28500,N_28568);
nand U28995 (N_28995,N_28527,N_28749);
nor U28996 (N_28996,N_28799,N_28709);
xnor U28997 (N_28997,N_28678,N_28756);
nor U28998 (N_28998,N_28553,N_28627);
and U28999 (N_28999,N_28514,N_28608);
nor U29000 (N_29000,N_28663,N_28590);
or U29001 (N_29001,N_28592,N_28616);
and U29002 (N_29002,N_28717,N_28665);
or U29003 (N_29003,N_28672,N_28692);
nor U29004 (N_29004,N_28560,N_28597);
and U29005 (N_29005,N_28507,N_28702);
nor U29006 (N_29006,N_28734,N_28554);
xnor U29007 (N_29007,N_28701,N_28577);
xor U29008 (N_29008,N_28617,N_28683);
xnor U29009 (N_29009,N_28621,N_28629);
nand U29010 (N_29010,N_28602,N_28676);
xnor U29011 (N_29011,N_28603,N_28708);
xor U29012 (N_29012,N_28644,N_28623);
nor U29013 (N_29013,N_28677,N_28580);
or U29014 (N_29014,N_28778,N_28522);
or U29015 (N_29015,N_28645,N_28664);
or U29016 (N_29016,N_28702,N_28748);
nor U29017 (N_29017,N_28564,N_28591);
nor U29018 (N_29018,N_28619,N_28610);
and U29019 (N_29019,N_28641,N_28655);
nand U29020 (N_29020,N_28685,N_28537);
nand U29021 (N_29021,N_28646,N_28728);
and U29022 (N_29022,N_28538,N_28750);
xor U29023 (N_29023,N_28594,N_28630);
nor U29024 (N_29024,N_28778,N_28630);
nand U29025 (N_29025,N_28503,N_28722);
and U29026 (N_29026,N_28613,N_28590);
or U29027 (N_29027,N_28580,N_28562);
nor U29028 (N_29028,N_28626,N_28792);
xor U29029 (N_29029,N_28603,N_28532);
nor U29030 (N_29030,N_28632,N_28721);
or U29031 (N_29031,N_28774,N_28582);
or U29032 (N_29032,N_28560,N_28712);
xor U29033 (N_29033,N_28559,N_28713);
nand U29034 (N_29034,N_28522,N_28738);
nand U29035 (N_29035,N_28580,N_28767);
nand U29036 (N_29036,N_28763,N_28736);
xor U29037 (N_29037,N_28750,N_28508);
nand U29038 (N_29038,N_28682,N_28705);
nor U29039 (N_29039,N_28714,N_28767);
nor U29040 (N_29040,N_28665,N_28785);
and U29041 (N_29041,N_28615,N_28609);
nand U29042 (N_29042,N_28544,N_28647);
and U29043 (N_29043,N_28653,N_28505);
nor U29044 (N_29044,N_28578,N_28657);
nor U29045 (N_29045,N_28785,N_28644);
xor U29046 (N_29046,N_28570,N_28608);
nand U29047 (N_29047,N_28690,N_28513);
or U29048 (N_29048,N_28587,N_28701);
nor U29049 (N_29049,N_28677,N_28734);
xor U29050 (N_29050,N_28553,N_28779);
nand U29051 (N_29051,N_28718,N_28602);
and U29052 (N_29052,N_28732,N_28563);
nor U29053 (N_29053,N_28591,N_28671);
xor U29054 (N_29054,N_28596,N_28654);
nor U29055 (N_29055,N_28733,N_28728);
or U29056 (N_29056,N_28711,N_28746);
xnor U29057 (N_29057,N_28762,N_28528);
or U29058 (N_29058,N_28743,N_28602);
nor U29059 (N_29059,N_28673,N_28506);
xnor U29060 (N_29060,N_28751,N_28660);
and U29061 (N_29061,N_28581,N_28641);
xnor U29062 (N_29062,N_28616,N_28797);
nor U29063 (N_29063,N_28575,N_28770);
xnor U29064 (N_29064,N_28735,N_28519);
nand U29065 (N_29065,N_28690,N_28595);
and U29066 (N_29066,N_28573,N_28718);
xor U29067 (N_29067,N_28715,N_28512);
xnor U29068 (N_29068,N_28583,N_28601);
or U29069 (N_29069,N_28761,N_28757);
nor U29070 (N_29070,N_28782,N_28681);
and U29071 (N_29071,N_28673,N_28589);
nand U29072 (N_29072,N_28554,N_28692);
and U29073 (N_29073,N_28623,N_28697);
xor U29074 (N_29074,N_28568,N_28668);
nand U29075 (N_29075,N_28744,N_28722);
and U29076 (N_29076,N_28520,N_28638);
nand U29077 (N_29077,N_28511,N_28794);
nor U29078 (N_29078,N_28585,N_28715);
xnor U29079 (N_29079,N_28605,N_28777);
and U29080 (N_29080,N_28751,N_28784);
xnor U29081 (N_29081,N_28619,N_28545);
nor U29082 (N_29082,N_28770,N_28556);
or U29083 (N_29083,N_28506,N_28697);
or U29084 (N_29084,N_28648,N_28528);
xnor U29085 (N_29085,N_28778,N_28545);
or U29086 (N_29086,N_28581,N_28643);
nor U29087 (N_29087,N_28611,N_28559);
or U29088 (N_29088,N_28694,N_28671);
nand U29089 (N_29089,N_28674,N_28766);
nor U29090 (N_29090,N_28550,N_28541);
or U29091 (N_29091,N_28769,N_28683);
nand U29092 (N_29092,N_28745,N_28553);
nor U29093 (N_29093,N_28647,N_28595);
xor U29094 (N_29094,N_28765,N_28547);
xnor U29095 (N_29095,N_28738,N_28591);
nand U29096 (N_29096,N_28570,N_28671);
nor U29097 (N_29097,N_28559,N_28665);
nor U29098 (N_29098,N_28558,N_28656);
nor U29099 (N_29099,N_28726,N_28527);
and U29100 (N_29100,N_28981,N_28911);
or U29101 (N_29101,N_28824,N_28982);
xnor U29102 (N_29102,N_28857,N_29029);
nor U29103 (N_29103,N_28984,N_28933);
or U29104 (N_29104,N_28927,N_28854);
or U29105 (N_29105,N_29051,N_29088);
nor U29106 (N_29106,N_28940,N_28871);
and U29107 (N_29107,N_29013,N_29095);
and U29108 (N_29108,N_28802,N_28990);
and U29109 (N_29109,N_29005,N_28936);
xor U29110 (N_29110,N_28809,N_28860);
and U29111 (N_29111,N_28995,N_28926);
nand U29112 (N_29112,N_28829,N_29050);
nand U29113 (N_29113,N_28916,N_29001);
nand U29114 (N_29114,N_28856,N_29081);
nor U29115 (N_29115,N_29073,N_29086);
nand U29116 (N_29116,N_28839,N_28954);
nand U29117 (N_29117,N_29010,N_28876);
or U29118 (N_29118,N_29057,N_29084);
and U29119 (N_29119,N_29056,N_28855);
nand U29120 (N_29120,N_29036,N_28844);
nor U29121 (N_29121,N_28810,N_28974);
nor U29122 (N_29122,N_29011,N_28814);
nor U29123 (N_29123,N_29049,N_28953);
nor U29124 (N_29124,N_29037,N_29031);
and U29125 (N_29125,N_28813,N_29039);
and U29126 (N_29126,N_29090,N_28828);
and U29127 (N_29127,N_28945,N_29038);
and U29128 (N_29128,N_28869,N_28837);
and U29129 (N_29129,N_28921,N_28887);
and U29130 (N_29130,N_28867,N_28820);
nor U29131 (N_29131,N_29042,N_28840);
nand U29132 (N_29132,N_28868,N_28834);
nor U29133 (N_29133,N_28909,N_28955);
and U29134 (N_29134,N_28967,N_28944);
and U29135 (N_29135,N_28975,N_29076);
and U29136 (N_29136,N_29070,N_29082);
nor U29137 (N_29137,N_29053,N_28920);
and U29138 (N_29138,N_28965,N_28932);
nand U29139 (N_29139,N_28978,N_28893);
xor U29140 (N_29140,N_28947,N_29069);
and U29141 (N_29141,N_28922,N_28847);
xor U29142 (N_29142,N_28859,N_29022);
xnor U29143 (N_29143,N_28956,N_28819);
nand U29144 (N_29144,N_29033,N_28845);
and U29145 (N_29145,N_28822,N_29058);
or U29146 (N_29146,N_29000,N_28923);
and U29147 (N_29147,N_29020,N_28960);
or U29148 (N_29148,N_28852,N_29028);
nand U29149 (N_29149,N_28880,N_29087);
and U29150 (N_29150,N_28864,N_28905);
nand U29151 (N_29151,N_29024,N_29016);
nand U29152 (N_29152,N_28818,N_28898);
or U29153 (N_29153,N_28918,N_28963);
nand U29154 (N_29154,N_28830,N_28806);
nand U29155 (N_29155,N_28997,N_28891);
and U29156 (N_29156,N_28889,N_28924);
and U29157 (N_29157,N_29059,N_28966);
or U29158 (N_29158,N_28968,N_28913);
xor U29159 (N_29159,N_28842,N_29097);
or U29160 (N_29160,N_29054,N_28989);
or U29161 (N_29161,N_29092,N_28900);
nand U29162 (N_29162,N_28964,N_29080);
and U29163 (N_29163,N_28914,N_28912);
nor U29164 (N_29164,N_28878,N_28804);
nand U29165 (N_29165,N_28831,N_29052);
nor U29166 (N_29166,N_28972,N_29014);
or U29167 (N_29167,N_29089,N_28985);
and U29168 (N_29168,N_28938,N_28904);
nand U29169 (N_29169,N_28925,N_29019);
and U29170 (N_29170,N_29021,N_28872);
nor U29171 (N_29171,N_29012,N_28890);
xnor U29172 (N_29172,N_28858,N_28883);
and U29173 (N_29173,N_28902,N_28976);
and U29174 (N_29174,N_28882,N_28992);
nand U29175 (N_29175,N_29018,N_28884);
xnor U29176 (N_29176,N_28915,N_29096);
and U29177 (N_29177,N_28942,N_28870);
xor U29178 (N_29178,N_28962,N_29035);
nand U29179 (N_29179,N_28812,N_28841);
or U29180 (N_29180,N_28811,N_28941);
or U29181 (N_29181,N_29060,N_28881);
and U29182 (N_29182,N_29025,N_29030);
or U29183 (N_29183,N_28886,N_28817);
and U29184 (N_29184,N_28983,N_29015);
nand U29185 (N_29185,N_28934,N_28980);
or U29186 (N_29186,N_28903,N_28987);
xor U29187 (N_29187,N_28959,N_28977);
nand U29188 (N_29188,N_28986,N_28907);
and U29189 (N_29189,N_29072,N_28815);
nand U29190 (N_29190,N_28800,N_28952);
nor U29191 (N_29191,N_28879,N_29006);
and U29192 (N_29192,N_28849,N_28994);
xor U29193 (N_29193,N_29002,N_28998);
or U29194 (N_29194,N_29047,N_28825);
nor U29195 (N_29195,N_28930,N_29027);
xor U29196 (N_29196,N_29045,N_29009);
nand U29197 (N_29197,N_28931,N_29066);
or U29198 (N_29198,N_28897,N_28894);
nand U29199 (N_29199,N_28950,N_28993);
or U29200 (N_29200,N_29078,N_29041);
nor U29201 (N_29201,N_29093,N_29046);
and U29202 (N_29202,N_28832,N_29068);
nor U29203 (N_29203,N_28835,N_28957);
and U29204 (N_29204,N_29094,N_28973);
nor U29205 (N_29205,N_28979,N_29064);
nor U29206 (N_29206,N_28850,N_28969);
nor U29207 (N_29207,N_28875,N_28958);
and U29208 (N_29208,N_28826,N_28991);
and U29209 (N_29209,N_28853,N_28838);
and U29210 (N_29210,N_28816,N_28877);
xor U29211 (N_29211,N_28805,N_29075);
nor U29212 (N_29212,N_28821,N_29007);
xnor U29213 (N_29213,N_28873,N_28843);
nand U29214 (N_29214,N_29043,N_28865);
and U29215 (N_29215,N_29003,N_29062);
nor U29216 (N_29216,N_28901,N_28919);
nor U29217 (N_29217,N_28949,N_28892);
nor U29218 (N_29218,N_29004,N_29044);
nor U29219 (N_29219,N_28971,N_28863);
or U29220 (N_29220,N_28861,N_29099);
or U29221 (N_29221,N_29063,N_28929);
xor U29222 (N_29222,N_28937,N_28895);
or U29223 (N_29223,N_29055,N_28948);
xnor U29224 (N_29224,N_28803,N_28808);
xor U29225 (N_29225,N_29061,N_28908);
nand U29226 (N_29226,N_28848,N_29083);
or U29227 (N_29227,N_29048,N_29091);
xnor U29228 (N_29228,N_28935,N_28833);
nor U29229 (N_29229,N_29074,N_29077);
or U29230 (N_29230,N_29079,N_29026);
xnor U29231 (N_29231,N_29065,N_28874);
nor U29232 (N_29232,N_28823,N_28851);
or U29233 (N_29233,N_28896,N_29023);
nand U29234 (N_29234,N_28917,N_28862);
or U29235 (N_29235,N_28999,N_29085);
and U29236 (N_29236,N_28988,N_28807);
or U29237 (N_29237,N_28885,N_28866);
nand U29238 (N_29238,N_28951,N_28899);
nor U29239 (N_29239,N_28939,N_28801);
and U29240 (N_29240,N_28946,N_29034);
nand U29241 (N_29241,N_29017,N_28827);
nor U29242 (N_29242,N_29032,N_28910);
nor U29243 (N_29243,N_28836,N_28846);
or U29244 (N_29244,N_29040,N_29067);
nor U29245 (N_29245,N_28928,N_28906);
xnor U29246 (N_29246,N_28970,N_28996);
nor U29247 (N_29247,N_29071,N_28961);
and U29248 (N_29248,N_28943,N_29098);
nand U29249 (N_29249,N_29008,N_28888);
nand U29250 (N_29250,N_28825,N_28863);
and U29251 (N_29251,N_28860,N_29004);
nand U29252 (N_29252,N_28979,N_29081);
xnor U29253 (N_29253,N_28879,N_28942);
or U29254 (N_29254,N_28995,N_28835);
and U29255 (N_29255,N_29040,N_28854);
or U29256 (N_29256,N_28981,N_29042);
nand U29257 (N_29257,N_29018,N_28868);
or U29258 (N_29258,N_29094,N_29036);
or U29259 (N_29259,N_29035,N_28952);
or U29260 (N_29260,N_28939,N_28933);
xnor U29261 (N_29261,N_28931,N_28949);
nor U29262 (N_29262,N_28908,N_28965);
nand U29263 (N_29263,N_28826,N_28996);
nor U29264 (N_29264,N_28978,N_28955);
or U29265 (N_29265,N_28915,N_28958);
or U29266 (N_29266,N_28906,N_29096);
or U29267 (N_29267,N_28874,N_28966);
nor U29268 (N_29268,N_28935,N_29062);
and U29269 (N_29269,N_29063,N_29076);
nor U29270 (N_29270,N_28877,N_28991);
nor U29271 (N_29271,N_28952,N_28823);
nor U29272 (N_29272,N_28994,N_28855);
nor U29273 (N_29273,N_28971,N_28801);
xnor U29274 (N_29274,N_28951,N_29052);
xor U29275 (N_29275,N_29004,N_29042);
xnor U29276 (N_29276,N_28839,N_28870);
xnor U29277 (N_29277,N_29010,N_28908);
nor U29278 (N_29278,N_29041,N_29037);
nand U29279 (N_29279,N_29091,N_29075);
xor U29280 (N_29280,N_28897,N_28882);
nand U29281 (N_29281,N_28975,N_29011);
nor U29282 (N_29282,N_28891,N_29019);
or U29283 (N_29283,N_28895,N_28833);
or U29284 (N_29284,N_28868,N_28983);
and U29285 (N_29285,N_28849,N_28909);
or U29286 (N_29286,N_29089,N_29017);
nand U29287 (N_29287,N_28875,N_28866);
xor U29288 (N_29288,N_28988,N_28817);
nand U29289 (N_29289,N_29051,N_28898);
and U29290 (N_29290,N_29065,N_28932);
nand U29291 (N_29291,N_28922,N_29093);
or U29292 (N_29292,N_29085,N_28995);
nand U29293 (N_29293,N_29016,N_28993);
and U29294 (N_29294,N_29048,N_28967);
or U29295 (N_29295,N_28895,N_29003);
nand U29296 (N_29296,N_28844,N_28962);
xnor U29297 (N_29297,N_28821,N_29023);
and U29298 (N_29298,N_29020,N_29096);
xor U29299 (N_29299,N_28807,N_29081);
or U29300 (N_29300,N_29011,N_28905);
or U29301 (N_29301,N_29028,N_29024);
and U29302 (N_29302,N_29032,N_28960);
xor U29303 (N_29303,N_29086,N_28973);
and U29304 (N_29304,N_29086,N_28925);
nand U29305 (N_29305,N_28914,N_28959);
nand U29306 (N_29306,N_28915,N_29085);
nor U29307 (N_29307,N_28829,N_28929);
nand U29308 (N_29308,N_28821,N_28895);
nand U29309 (N_29309,N_29080,N_28872);
nor U29310 (N_29310,N_29027,N_29075);
or U29311 (N_29311,N_28932,N_28848);
nor U29312 (N_29312,N_28955,N_28854);
nor U29313 (N_29313,N_29068,N_28904);
or U29314 (N_29314,N_28837,N_28884);
nand U29315 (N_29315,N_28876,N_29082);
xor U29316 (N_29316,N_28838,N_28803);
and U29317 (N_29317,N_28833,N_28995);
and U29318 (N_29318,N_28816,N_28957);
nand U29319 (N_29319,N_28828,N_28904);
nand U29320 (N_29320,N_28965,N_28895);
xnor U29321 (N_29321,N_28882,N_28986);
nor U29322 (N_29322,N_29028,N_28949);
nor U29323 (N_29323,N_28904,N_29035);
xor U29324 (N_29324,N_29076,N_28836);
nor U29325 (N_29325,N_29007,N_29083);
nor U29326 (N_29326,N_28954,N_29093);
or U29327 (N_29327,N_29033,N_28834);
nand U29328 (N_29328,N_28999,N_28921);
xor U29329 (N_29329,N_29077,N_28955);
or U29330 (N_29330,N_28877,N_28828);
xnor U29331 (N_29331,N_28998,N_28987);
and U29332 (N_29332,N_28942,N_28969);
nor U29333 (N_29333,N_28993,N_28888);
nor U29334 (N_29334,N_28827,N_28999);
or U29335 (N_29335,N_28813,N_29028);
nand U29336 (N_29336,N_29080,N_28835);
nand U29337 (N_29337,N_28994,N_29077);
nor U29338 (N_29338,N_29039,N_28804);
or U29339 (N_29339,N_28803,N_29043);
nand U29340 (N_29340,N_29055,N_29068);
nor U29341 (N_29341,N_28880,N_29061);
xor U29342 (N_29342,N_29039,N_29052);
xnor U29343 (N_29343,N_29067,N_28889);
nor U29344 (N_29344,N_28843,N_28963);
nor U29345 (N_29345,N_28941,N_28877);
nor U29346 (N_29346,N_28923,N_28809);
xnor U29347 (N_29347,N_29023,N_29079);
and U29348 (N_29348,N_28974,N_28845);
xor U29349 (N_29349,N_29057,N_28826);
xnor U29350 (N_29350,N_28929,N_29099);
and U29351 (N_29351,N_29015,N_28936);
nand U29352 (N_29352,N_29071,N_28880);
and U29353 (N_29353,N_28804,N_28801);
nand U29354 (N_29354,N_28818,N_29011);
and U29355 (N_29355,N_29054,N_28916);
and U29356 (N_29356,N_28823,N_29043);
nor U29357 (N_29357,N_28910,N_28948);
or U29358 (N_29358,N_29043,N_28834);
or U29359 (N_29359,N_28805,N_29016);
or U29360 (N_29360,N_28930,N_28956);
and U29361 (N_29361,N_29095,N_28980);
xor U29362 (N_29362,N_29056,N_28944);
nor U29363 (N_29363,N_28924,N_29030);
and U29364 (N_29364,N_28844,N_28856);
nand U29365 (N_29365,N_28933,N_28916);
nand U29366 (N_29366,N_29057,N_29048);
nor U29367 (N_29367,N_29043,N_28804);
nor U29368 (N_29368,N_28869,N_28946);
xor U29369 (N_29369,N_29008,N_28997);
or U29370 (N_29370,N_29041,N_28907);
nand U29371 (N_29371,N_28880,N_28808);
nand U29372 (N_29372,N_29043,N_29057);
nand U29373 (N_29373,N_29083,N_28893);
nor U29374 (N_29374,N_28872,N_28828);
xnor U29375 (N_29375,N_28932,N_29082);
xnor U29376 (N_29376,N_28844,N_28996);
and U29377 (N_29377,N_29060,N_28961);
and U29378 (N_29378,N_28872,N_28829);
or U29379 (N_29379,N_28896,N_28846);
and U29380 (N_29380,N_28923,N_28819);
nor U29381 (N_29381,N_29000,N_28908);
xor U29382 (N_29382,N_29041,N_28931);
nor U29383 (N_29383,N_28854,N_28889);
or U29384 (N_29384,N_28877,N_29032);
xor U29385 (N_29385,N_28982,N_28818);
xor U29386 (N_29386,N_29083,N_28836);
nor U29387 (N_29387,N_28915,N_28847);
nor U29388 (N_29388,N_28950,N_29022);
and U29389 (N_29389,N_28934,N_28801);
nor U29390 (N_29390,N_28918,N_29095);
nand U29391 (N_29391,N_28928,N_28979);
nand U29392 (N_29392,N_29054,N_29050);
xnor U29393 (N_29393,N_28958,N_28858);
nor U29394 (N_29394,N_29022,N_29014);
or U29395 (N_29395,N_28918,N_28845);
nand U29396 (N_29396,N_28874,N_28897);
nor U29397 (N_29397,N_29095,N_29097);
nor U29398 (N_29398,N_29065,N_28916);
nor U29399 (N_29399,N_28924,N_28890);
nor U29400 (N_29400,N_29311,N_29324);
nand U29401 (N_29401,N_29159,N_29138);
nor U29402 (N_29402,N_29209,N_29183);
nor U29403 (N_29403,N_29127,N_29297);
and U29404 (N_29404,N_29397,N_29139);
or U29405 (N_29405,N_29181,N_29117);
or U29406 (N_29406,N_29275,N_29145);
and U29407 (N_29407,N_29102,N_29298);
xor U29408 (N_29408,N_29351,N_29168);
xnor U29409 (N_29409,N_29252,N_29326);
nor U29410 (N_29410,N_29287,N_29355);
or U29411 (N_29411,N_29151,N_29122);
and U29412 (N_29412,N_29106,N_29233);
or U29413 (N_29413,N_29308,N_29246);
nand U29414 (N_29414,N_29382,N_29156);
or U29415 (N_29415,N_29202,N_29273);
nor U29416 (N_29416,N_29339,N_29258);
xor U29417 (N_29417,N_29388,N_29132);
nand U29418 (N_29418,N_29242,N_29303);
xnor U29419 (N_29419,N_29200,N_29197);
and U29420 (N_29420,N_29364,N_29315);
nand U29421 (N_29421,N_29111,N_29280);
or U29422 (N_29422,N_29128,N_29229);
xor U29423 (N_29423,N_29161,N_29206);
nand U29424 (N_29424,N_29332,N_29396);
or U29425 (N_29425,N_29329,N_29187);
and U29426 (N_29426,N_29283,N_29194);
nor U29427 (N_29427,N_29386,N_29336);
nand U29428 (N_29428,N_29251,N_29387);
and U29429 (N_29429,N_29141,N_29208);
and U29430 (N_29430,N_29193,N_29333);
xnor U29431 (N_29431,N_29366,N_29293);
nand U29432 (N_29432,N_29214,N_29266);
nand U29433 (N_29433,N_29392,N_29325);
xor U29434 (N_29434,N_29395,N_29112);
nand U29435 (N_29435,N_29224,N_29152);
xor U29436 (N_29436,N_29317,N_29256);
nor U29437 (N_29437,N_29399,N_29365);
nor U29438 (N_29438,N_29144,N_29162);
and U29439 (N_29439,N_29270,N_29278);
or U29440 (N_29440,N_29157,N_29116);
nand U29441 (N_29441,N_29158,N_29346);
xnor U29442 (N_29442,N_29115,N_29340);
xnor U29443 (N_29443,N_29153,N_29222);
nor U29444 (N_29444,N_29105,N_29100);
nor U29445 (N_29445,N_29221,N_29369);
nand U29446 (N_29446,N_29248,N_29295);
and U29447 (N_29447,N_29334,N_29367);
and U29448 (N_29448,N_29368,N_29140);
xor U29449 (N_29449,N_29265,N_29204);
xnor U29450 (N_29450,N_29330,N_29241);
xor U29451 (N_29451,N_29288,N_29338);
or U29452 (N_29452,N_29376,N_29189);
or U29453 (N_29453,N_29166,N_29307);
or U29454 (N_29454,N_29123,N_29378);
nand U29455 (N_29455,N_29199,N_29302);
xnor U29456 (N_29456,N_29321,N_29306);
nor U29457 (N_29457,N_29104,N_29174);
or U29458 (N_29458,N_29154,N_29380);
and U29459 (N_29459,N_29149,N_29212);
or U29460 (N_29460,N_29309,N_29289);
nor U29461 (N_29461,N_29356,N_29377);
and U29462 (N_29462,N_29205,N_29103);
or U29463 (N_29463,N_29391,N_29147);
or U29464 (N_29464,N_29284,N_29237);
or U29465 (N_29465,N_29171,N_29260);
or U29466 (N_29466,N_29163,N_29195);
nand U29467 (N_29467,N_29286,N_29322);
or U29468 (N_29468,N_29245,N_29375);
xor U29469 (N_29469,N_29381,N_29108);
or U29470 (N_29470,N_29394,N_29259);
and U29471 (N_29471,N_29169,N_29190);
and U29472 (N_29472,N_29337,N_29316);
nand U29473 (N_29473,N_29213,N_29341);
and U29474 (N_29474,N_29335,N_29384);
nor U29475 (N_29475,N_29276,N_29107);
nor U29476 (N_29476,N_29314,N_29211);
and U29477 (N_29477,N_29185,N_29347);
or U29478 (N_29478,N_29285,N_29320);
nor U29479 (N_29479,N_29191,N_29274);
nand U29480 (N_29480,N_29217,N_29305);
and U29481 (N_29481,N_29370,N_29360);
nor U29482 (N_29482,N_29349,N_29198);
and U29483 (N_29483,N_29186,N_29167);
nor U29484 (N_29484,N_29264,N_29216);
nand U29485 (N_29485,N_29113,N_29210);
nand U29486 (N_29486,N_29226,N_29249);
nor U29487 (N_29487,N_29268,N_29160);
nand U29488 (N_29488,N_29121,N_29318);
and U29489 (N_29489,N_29379,N_29371);
and U29490 (N_29490,N_29150,N_29155);
nand U29491 (N_29491,N_29331,N_29136);
or U29492 (N_29492,N_29133,N_29184);
nand U29493 (N_29493,N_29130,N_29119);
and U29494 (N_29494,N_29243,N_29227);
and U29495 (N_29495,N_29291,N_29219);
and U29496 (N_29496,N_29148,N_29247);
or U29497 (N_29497,N_29277,N_29345);
nor U29498 (N_29498,N_29348,N_29281);
or U29499 (N_29499,N_29129,N_29196);
xor U29500 (N_29500,N_29207,N_29257);
or U29501 (N_29501,N_29238,N_29301);
xnor U29502 (N_29502,N_29310,N_29393);
xnor U29503 (N_29503,N_29269,N_29101);
xnor U29504 (N_29504,N_29353,N_29383);
xor U29505 (N_29505,N_29173,N_29352);
nand U29506 (N_29506,N_29262,N_29267);
xor U29507 (N_29507,N_29299,N_29358);
and U29508 (N_29508,N_29176,N_29240);
and U29509 (N_29509,N_29296,N_29385);
and U29510 (N_29510,N_29126,N_29361);
or U29511 (N_29511,N_29110,N_29244);
and U29512 (N_29512,N_29327,N_29342);
nand U29513 (N_29513,N_29373,N_29343);
xnor U29514 (N_29514,N_29182,N_29137);
nand U29515 (N_29515,N_29263,N_29319);
or U29516 (N_29516,N_29225,N_29254);
and U29517 (N_29517,N_29362,N_29218);
nor U29518 (N_29518,N_29118,N_29304);
or U29519 (N_29519,N_29372,N_29312);
nand U29520 (N_29520,N_29175,N_29374);
or U29521 (N_29521,N_29313,N_29239);
nor U29522 (N_29522,N_29255,N_29170);
nor U29523 (N_29523,N_29178,N_29201);
or U29524 (N_29524,N_29228,N_29142);
or U29525 (N_29525,N_29294,N_29165);
nand U29526 (N_29526,N_29253,N_29220);
nand U29527 (N_29527,N_29344,N_29215);
and U29528 (N_29528,N_29230,N_29179);
nand U29529 (N_29529,N_29250,N_29120);
or U29530 (N_29530,N_29134,N_29292);
xor U29531 (N_29531,N_29146,N_29143);
and U29532 (N_29532,N_29272,N_29235);
or U29533 (N_29533,N_29223,N_29164);
nor U29534 (N_29534,N_29135,N_29300);
and U29535 (N_29535,N_29180,N_29357);
and U29536 (N_29536,N_29236,N_29203);
or U29537 (N_29537,N_29398,N_29131);
or U29538 (N_29538,N_29323,N_29192);
nor U29539 (N_29539,N_29109,N_29125);
nand U29540 (N_29540,N_29363,N_29354);
nand U29541 (N_29541,N_29177,N_29271);
xor U29542 (N_29542,N_29390,N_29328);
nand U29543 (N_29543,N_29350,N_29290);
nand U29544 (N_29544,N_29261,N_29282);
or U29545 (N_29545,N_29124,N_29114);
xnor U29546 (N_29546,N_29234,N_29232);
or U29547 (N_29547,N_29279,N_29389);
or U29548 (N_29548,N_29231,N_29188);
nor U29549 (N_29549,N_29359,N_29172);
xnor U29550 (N_29550,N_29114,N_29326);
or U29551 (N_29551,N_29323,N_29128);
or U29552 (N_29552,N_29141,N_29253);
xor U29553 (N_29553,N_29341,N_29337);
nand U29554 (N_29554,N_29126,N_29268);
nand U29555 (N_29555,N_29392,N_29380);
or U29556 (N_29556,N_29334,N_29116);
nor U29557 (N_29557,N_29286,N_29300);
and U29558 (N_29558,N_29196,N_29354);
or U29559 (N_29559,N_29155,N_29148);
xor U29560 (N_29560,N_29166,N_29226);
nor U29561 (N_29561,N_29264,N_29328);
xnor U29562 (N_29562,N_29107,N_29182);
or U29563 (N_29563,N_29255,N_29335);
xor U29564 (N_29564,N_29292,N_29226);
or U29565 (N_29565,N_29298,N_29339);
and U29566 (N_29566,N_29370,N_29275);
and U29567 (N_29567,N_29246,N_29104);
nand U29568 (N_29568,N_29364,N_29131);
xor U29569 (N_29569,N_29309,N_29189);
nor U29570 (N_29570,N_29170,N_29267);
or U29571 (N_29571,N_29275,N_29346);
and U29572 (N_29572,N_29281,N_29280);
xor U29573 (N_29573,N_29327,N_29258);
or U29574 (N_29574,N_29213,N_29275);
or U29575 (N_29575,N_29333,N_29340);
nor U29576 (N_29576,N_29169,N_29330);
nor U29577 (N_29577,N_29124,N_29169);
or U29578 (N_29578,N_29217,N_29139);
xnor U29579 (N_29579,N_29249,N_29395);
xnor U29580 (N_29580,N_29100,N_29190);
or U29581 (N_29581,N_29382,N_29101);
nor U29582 (N_29582,N_29214,N_29182);
and U29583 (N_29583,N_29355,N_29382);
nor U29584 (N_29584,N_29185,N_29121);
and U29585 (N_29585,N_29319,N_29251);
and U29586 (N_29586,N_29350,N_29110);
nor U29587 (N_29587,N_29366,N_29348);
or U29588 (N_29588,N_29148,N_29200);
and U29589 (N_29589,N_29304,N_29296);
nand U29590 (N_29590,N_29392,N_29298);
nand U29591 (N_29591,N_29129,N_29252);
and U29592 (N_29592,N_29234,N_29101);
and U29593 (N_29593,N_29126,N_29260);
xor U29594 (N_29594,N_29332,N_29222);
and U29595 (N_29595,N_29361,N_29150);
xnor U29596 (N_29596,N_29118,N_29276);
or U29597 (N_29597,N_29369,N_29155);
nor U29598 (N_29598,N_29201,N_29224);
xnor U29599 (N_29599,N_29183,N_29358);
and U29600 (N_29600,N_29156,N_29110);
xnor U29601 (N_29601,N_29321,N_29179);
nor U29602 (N_29602,N_29335,N_29303);
or U29603 (N_29603,N_29250,N_29227);
or U29604 (N_29604,N_29354,N_29192);
xnor U29605 (N_29605,N_29172,N_29230);
nor U29606 (N_29606,N_29178,N_29229);
and U29607 (N_29607,N_29277,N_29112);
nand U29608 (N_29608,N_29190,N_29136);
xnor U29609 (N_29609,N_29392,N_29176);
nand U29610 (N_29610,N_29286,N_29166);
or U29611 (N_29611,N_29129,N_29201);
xor U29612 (N_29612,N_29393,N_29229);
xnor U29613 (N_29613,N_29355,N_29176);
xnor U29614 (N_29614,N_29338,N_29284);
xnor U29615 (N_29615,N_29359,N_29106);
nor U29616 (N_29616,N_29374,N_29293);
nand U29617 (N_29617,N_29378,N_29379);
and U29618 (N_29618,N_29115,N_29308);
xnor U29619 (N_29619,N_29298,N_29346);
nor U29620 (N_29620,N_29388,N_29168);
xor U29621 (N_29621,N_29380,N_29376);
xor U29622 (N_29622,N_29191,N_29111);
or U29623 (N_29623,N_29376,N_29213);
or U29624 (N_29624,N_29176,N_29204);
nand U29625 (N_29625,N_29277,N_29363);
nand U29626 (N_29626,N_29332,N_29303);
xor U29627 (N_29627,N_29119,N_29246);
or U29628 (N_29628,N_29175,N_29170);
xnor U29629 (N_29629,N_29209,N_29185);
and U29630 (N_29630,N_29390,N_29381);
or U29631 (N_29631,N_29319,N_29303);
xor U29632 (N_29632,N_29372,N_29130);
and U29633 (N_29633,N_29113,N_29303);
or U29634 (N_29634,N_29339,N_29285);
and U29635 (N_29635,N_29339,N_29287);
nand U29636 (N_29636,N_29134,N_29271);
xor U29637 (N_29637,N_29194,N_29237);
or U29638 (N_29638,N_29226,N_29196);
and U29639 (N_29639,N_29280,N_29314);
xnor U29640 (N_29640,N_29268,N_29173);
xnor U29641 (N_29641,N_29351,N_29262);
xor U29642 (N_29642,N_29315,N_29270);
nor U29643 (N_29643,N_29361,N_29173);
xor U29644 (N_29644,N_29187,N_29242);
and U29645 (N_29645,N_29253,N_29294);
nand U29646 (N_29646,N_29277,N_29250);
and U29647 (N_29647,N_29326,N_29240);
or U29648 (N_29648,N_29126,N_29141);
or U29649 (N_29649,N_29211,N_29267);
and U29650 (N_29650,N_29257,N_29186);
nor U29651 (N_29651,N_29331,N_29262);
and U29652 (N_29652,N_29216,N_29156);
nand U29653 (N_29653,N_29170,N_29106);
and U29654 (N_29654,N_29139,N_29228);
xnor U29655 (N_29655,N_29377,N_29206);
xor U29656 (N_29656,N_29266,N_29376);
or U29657 (N_29657,N_29144,N_29283);
nand U29658 (N_29658,N_29143,N_29296);
nand U29659 (N_29659,N_29149,N_29127);
nor U29660 (N_29660,N_29177,N_29145);
nand U29661 (N_29661,N_29249,N_29193);
nand U29662 (N_29662,N_29211,N_29379);
xor U29663 (N_29663,N_29311,N_29262);
xnor U29664 (N_29664,N_29376,N_29172);
xor U29665 (N_29665,N_29344,N_29185);
or U29666 (N_29666,N_29146,N_29337);
nand U29667 (N_29667,N_29369,N_29343);
nor U29668 (N_29668,N_29282,N_29253);
nand U29669 (N_29669,N_29287,N_29123);
nand U29670 (N_29670,N_29319,N_29253);
nand U29671 (N_29671,N_29380,N_29290);
nand U29672 (N_29672,N_29381,N_29113);
nor U29673 (N_29673,N_29261,N_29320);
nand U29674 (N_29674,N_29389,N_29216);
nand U29675 (N_29675,N_29322,N_29164);
nor U29676 (N_29676,N_29356,N_29123);
nand U29677 (N_29677,N_29288,N_29340);
nand U29678 (N_29678,N_29221,N_29269);
and U29679 (N_29679,N_29245,N_29394);
and U29680 (N_29680,N_29338,N_29178);
nor U29681 (N_29681,N_29329,N_29326);
and U29682 (N_29682,N_29165,N_29172);
and U29683 (N_29683,N_29323,N_29393);
or U29684 (N_29684,N_29249,N_29385);
nor U29685 (N_29685,N_29300,N_29352);
nor U29686 (N_29686,N_29312,N_29226);
nor U29687 (N_29687,N_29363,N_29375);
or U29688 (N_29688,N_29189,N_29357);
or U29689 (N_29689,N_29268,N_29119);
xor U29690 (N_29690,N_29327,N_29103);
or U29691 (N_29691,N_29157,N_29177);
nand U29692 (N_29692,N_29277,N_29171);
xor U29693 (N_29693,N_29126,N_29389);
and U29694 (N_29694,N_29383,N_29190);
nor U29695 (N_29695,N_29190,N_29292);
nor U29696 (N_29696,N_29389,N_29341);
and U29697 (N_29697,N_29243,N_29145);
nand U29698 (N_29698,N_29360,N_29297);
xnor U29699 (N_29699,N_29205,N_29319);
nor U29700 (N_29700,N_29667,N_29564);
and U29701 (N_29701,N_29660,N_29690);
nand U29702 (N_29702,N_29466,N_29481);
and U29703 (N_29703,N_29599,N_29537);
nor U29704 (N_29704,N_29426,N_29516);
or U29705 (N_29705,N_29566,N_29402);
or U29706 (N_29706,N_29651,N_29683);
nand U29707 (N_29707,N_29561,N_29530);
nor U29708 (N_29708,N_29477,N_29638);
xnor U29709 (N_29709,N_29512,N_29440);
and U29710 (N_29710,N_29511,N_29431);
and U29711 (N_29711,N_29586,N_29665);
and U29712 (N_29712,N_29614,N_29653);
nor U29713 (N_29713,N_29626,N_29613);
nand U29714 (N_29714,N_29585,N_29423);
nor U29715 (N_29715,N_29538,N_29501);
xnor U29716 (N_29716,N_29528,N_29699);
nor U29717 (N_29717,N_29598,N_29607);
nand U29718 (N_29718,N_29438,N_29546);
or U29719 (N_29719,N_29458,N_29587);
nand U29720 (N_29720,N_29502,N_29418);
xnor U29721 (N_29721,N_29403,N_29694);
xor U29722 (N_29722,N_29487,N_29539);
nand U29723 (N_29723,N_29689,N_29496);
and U29724 (N_29724,N_29497,N_29636);
nor U29725 (N_29725,N_29474,N_29483);
nor U29726 (N_29726,N_29644,N_29556);
nand U29727 (N_29727,N_29411,N_29577);
nand U29728 (N_29728,N_29602,N_29562);
or U29729 (N_29729,N_29567,N_29643);
xor U29730 (N_29730,N_29685,N_29439);
xor U29731 (N_29731,N_29475,N_29434);
or U29732 (N_29732,N_29415,N_29491);
nor U29733 (N_29733,N_29473,N_29414);
and U29734 (N_29734,N_29633,N_29432);
and U29735 (N_29735,N_29507,N_29449);
nor U29736 (N_29736,N_29547,N_29428);
nor U29737 (N_29737,N_29533,N_29489);
nor U29738 (N_29738,N_29608,N_29605);
xor U29739 (N_29739,N_29529,N_29583);
xor U29740 (N_29740,N_29488,N_29435);
nor U29741 (N_29741,N_29593,N_29408);
and U29742 (N_29742,N_29629,N_29563);
nand U29743 (N_29743,N_29551,N_29464);
or U29744 (N_29744,N_29407,N_29601);
xnor U29745 (N_29745,N_29559,N_29553);
nand U29746 (N_29746,N_29430,N_29612);
nor U29747 (N_29747,N_29641,N_29446);
xor U29748 (N_29748,N_29632,N_29600);
and U29749 (N_29749,N_29517,N_29575);
or U29750 (N_29750,N_29549,N_29630);
nor U29751 (N_29751,N_29558,N_29445);
or U29752 (N_29752,N_29659,N_29437);
and U29753 (N_29753,N_29621,N_29588);
nor U29754 (N_29754,N_29603,N_29480);
nand U29755 (N_29755,N_29425,N_29527);
and U29756 (N_29756,N_29436,N_29670);
or U29757 (N_29757,N_29451,N_29554);
nor U29758 (N_29758,N_29625,N_29617);
nand U29759 (N_29759,N_29574,N_29655);
nor U29760 (N_29760,N_29597,N_29518);
and U29761 (N_29761,N_29461,N_29457);
nor U29762 (N_29762,N_29637,N_29526);
xor U29763 (N_29763,N_29623,N_29687);
or U29764 (N_29764,N_29634,N_29628);
nor U29765 (N_29765,N_29419,N_29532);
or U29766 (N_29766,N_29521,N_29669);
xor U29767 (N_29767,N_29478,N_29500);
and U29768 (N_29768,N_29460,N_29698);
nand U29769 (N_29769,N_29677,N_29544);
or U29770 (N_29770,N_29592,N_29609);
nand U29771 (N_29771,N_29424,N_29686);
nand U29772 (N_29772,N_29443,N_29666);
and U29773 (N_29773,N_29467,N_29557);
xor U29774 (N_29774,N_29627,N_29681);
nand U29775 (N_29775,N_29565,N_29406);
and U29776 (N_29776,N_29472,N_29486);
and U29777 (N_29777,N_29676,N_29657);
xnor U29778 (N_29778,N_29450,N_29688);
and U29779 (N_29779,N_29479,N_29535);
and U29780 (N_29780,N_29648,N_29620);
or U29781 (N_29781,N_29662,N_29646);
or U29782 (N_29782,N_29661,N_29695);
nand U29783 (N_29783,N_29409,N_29570);
xnor U29784 (N_29784,N_29606,N_29456);
and U29785 (N_29785,N_29624,N_29484);
or U29786 (N_29786,N_29691,N_29581);
or U29787 (N_29787,N_29519,N_29673);
nor U29788 (N_29788,N_29668,N_29639);
or U29789 (N_29789,N_29468,N_29444);
nand U29790 (N_29790,N_29679,N_29550);
nand U29791 (N_29791,N_29524,N_29604);
or U29792 (N_29792,N_29469,N_29654);
nor U29793 (N_29793,N_29494,N_29642);
and U29794 (N_29794,N_29455,N_29692);
xnor U29795 (N_29795,N_29442,N_29522);
and U29796 (N_29796,N_29459,N_29454);
or U29797 (N_29797,N_29647,N_29552);
and U29798 (N_29798,N_29515,N_29576);
xnor U29799 (N_29799,N_29578,N_29584);
xor U29800 (N_29800,N_29693,N_29568);
nor U29801 (N_29801,N_29509,N_29674);
xor U29802 (N_29802,N_29678,N_29572);
xnor U29803 (N_29803,N_29635,N_29548);
nor U29804 (N_29804,N_29672,N_29611);
xor U29805 (N_29805,N_29560,N_29416);
or U29806 (N_29806,N_29463,N_29405);
and U29807 (N_29807,N_29596,N_29429);
nor U29808 (N_29808,N_29680,N_29619);
nand U29809 (N_29809,N_29671,N_29421);
nor U29810 (N_29810,N_29555,N_29675);
xnor U29811 (N_29811,N_29525,N_29656);
nand U29812 (N_29812,N_29697,N_29401);
or U29813 (N_29813,N_29582,N_29490);
and U29814 (N_29814,N_29536,N_29573);
xnor U29815 (N_29815,N_29513,N_29470);
nor U29816 (N_29816,N_29652,N_29493);
xnor U29817 (N_29817,N_29492,N_29508);
or U29818 (N_29818,N_29400,N_29417);
xnor U29819 (N_29819,N_29412,N_29594);
xor U29820 (N_29820,N_29545,N_29413);
nor U29821 (N_29821,N_29618,N_29523);
and U29822 (N_29822,N_29616,N_29540);
xor U29823 (N_29823,N_29453,N_29542);
and U29824 (N_29824,N_29591,N_29441);
xor U29825 (N_29825,N_29541,N_29471);
or U29826 (N_29826,N_29543,N_29645);
nor U29827 (N_29827,N_29682,N_29448);
and U29828 (N_29828,N_29498,N_29571);
xor U29829 (N_29829,N_29465,N_29505);
nand U29830 (N_29830,N_29520,N_29595);
and U29831 (N_29831,N_29531,N_29514);
nor U29832 (N_29832,N_29610,N_29485);
and U29833 (N_29833,N_29650,N_29649);
nor U29834 (N_29834,N_29534,N_29663);
and U29835 (N_29835,N_29499,N_29410);
nor U29836 (N_29836,N_29482,N_29658);
nor U29837 (N_29837,N_29615,N_29569);
xnor U29838 (N_29838,N_29447,N_29684);
and U29839 (N_29839,N_29622,N_29404);
nand U29840 (N_29840,N_29579,N_29580);
or U29841 (N_29841,N_29631,N_29504);
or U29842 (N_29842,N_29420,N_29510);
or U29843 (N_29843,N_29476,N_29589);
xor U29844 (N_29844,N_29664,N_29506);
nand U29845 (N_29845,N_29422,N_29427);
or U29846 (N_29846,N_29452,N_29503);
nand U29847 (N_29847,N_29640,N_29462);
nand U29848 (N_29848,N_29433,N_29590);
or U29849 (N_29849,N_29495,N_29696);
nand U29850 (N_29850,N_29507,N_29565);
nand U29851 (N_29851,N_29405,N_29623);
xor U29852 (N_29852,N_29647,N_29672);
xor U29853 (N_29853,N_29621,N_29591);
xnor U29854 (N_29854,N_29625,N_29464);
xor U29855 (N_29855,N_29630,N_29593);
and U29856 (N_29856,N_29485,N_29650);
xor U29857 (N_29857,N_29554,N_29547);
or U29858 (N_29858,N_29407,N_29543);
nor U29859 (N_29859,N_29661,N_29407);
and U29860 (N_29860,N_29643,N_29587);
nor U29861 (N_29861,N_29438,N_29515);
nand U29862 (N_29862,N_29639,N_29623);
nand U29863 (N_29863,N_29695,N_29556);
nand U29864 (N_29864,N_29622,N_29616);
xnor U29865 (N_29865,N_29534,N_29492);
nor U29866 (N_29866,N_29445,N_29585);
and U29867 (N_29867,N_29638,N_29445);
nor U29868 (N_29868,N_29618,N_29625);
or U29869 (N_29869,N_29585,N_29513);
nand U29870 (N_29870,N_29611,N_29558);
and U29871 (N_29871,N_29681,N_29519);
nand U29872 (N_29872,N_29680,N_29539);
nand U29873 (N_29873,N_29635,N_29674);
and U29874 (N_29874,N_29533,N_29483);
nor U29875 (N_29875,N_29452,N_29524);
nor U29876 (N_29876,N_29497,N_29552);
nor U29877 (N_29877,N_29428,N_29413);
and U29878 (N_29878,N_29628,N_29521);
nor U29879 (N_29879,N_29452,N_29692);
nor U29880 (N_29880,N_29465,N_29668);
or U29881 (N_29881,N_29478,N_29661);
xnor U29882 (N_29882,N_29404,N_29478);
nor U29883 (N_29883,N_29481,N_29433);
nor U29884 (N_29884,N_29629,N_29555);
nand U29885 (N_29885,N_29494,N_29459);
nor U29886 (N_29886,N_29402,N_29604);
nor U29887 (N_29887,N_29504,N_29538);
or U29888 (N_29888,N_29400,N_29538);
or U29889 (N_29889,N_29546,N_29663);
or U29890 (N_29890,N_29626,N_29452);
xor U29891 (N_29891,N_29575,N_29516);
nor U29892 (N_29892,N_29657,N_29605);
nor U29893 (N_29893,N_29457,N_29491);
and U29894 (N_29894,N_29691,N_29584);
nand U29895 (N_29895,N_29693,N_29683);
xor U29896 (N_29896,N_29446,N_29510);
and U29897 (N_29897,N_29404,N_29558);
or U29898 (N_29898,N_29427,N_29437);
and U29899 (N_29899,N_29695,N_29528);
or U29900 (N_29900,N_29559,N_29540);
nand U29901 (N_29901,N_29499,N_29463);
xor U29902 (N_29902,N_29615,N_29666);
or U29903 (N_29903,N_29652,N_29415);
nand U29904 (N_29904,N_29596,N_29699);
nor U29905 (N_29905,N_29405,N_29499);
and U29906 (N_29906,N_29570,N_29464);
or U29907 (N_29907,N_29460,N_29628);
or U29908 (N_29908,N_29585,N_29598);
nor U29909 (N_29909,N_29580,N_29633);
nor U29910 (N_29910,N_29613,N_29671);
or U29911 (N_29911,N_29577,N_29604);
and U29912 (N_29912,N_29565,N_29592);
xor U29913 (N_29913,N_29416,N_29647);
xnor U29914 (N_29914,N_29684,N_29449);
nand U29915 (N_29915,N_29542,N_29617);
and U29916 (N_29916,N_29468,N_29569);
nor U29917 (N_29917,N_29500,N_29609);
nand U29918 (N_29918,N_29676,N_29408);
and U29919 (N_29919,N_29485,N_29675);
xnor U29920 (N_29920,N_29489,N_29459);
nand U29921 (N_29921,N_29624,N_29421);
nand U29922 (N_29922,N_29605,N_29494);
and U29923 (N_29923,N_29529,N_29661);
nor U29924 (N_29924,N_29405,N_29445);
or U29925 (N_29925,N_29493,N_29600);
and U29926 (N_29926,N_29578,N_29615);
and U29927 (N_29927,N_29586,N_29476);
nor U29928 (N_29928,N_29585,N_29687);
or U29929 (N_29929,N_29680,N_29693);
xor U29930 (N_29930,N_29526,N_29569);
or U29931 (N_29931,N_29598,N_29446);
nor U29932 (N_29932,N_29494,N_29530);
and U29933 (N_29933,N_29541,N_29436);
xnor U29934 (N_29934,N_29477,N_29416);
nand U29935 (N_29935,N_29611,N_29685);
nor U29936 (N_29936,N_29418,N_29669);
xnor U29937 (N_29937,N_29586,N_29424);
nand U29938 (N_29938,N_29578,N_29477);
nand U29939 (N_29939,N_29634,N_29578);
nor U29940 (N_29940,N_29473,N_29477);
or U29941 (N_29941,N_29552,N_29566);
nor U29942 (N_29942,N_29640,N_29502);
and U29943 (N_29943,N_29685,N_29407);
and U29944 (N_29944,N_29412,N_29541);
nand U29945 (N_29945,N_29547,N_29594);
or U29946 (N_29946,N_29584,N_29479);
nand U29947 (N_29947,N_29621,N_29489);
and U29948 (N_29948,N_29514,N_29416);
xnor U29949 (N_29949,N_29432,N_29526);
nor U29950 (N_29950,N_29558,N_29628);
xor U29951 (N_29951,N_29615,N_29598);
nor U29952 (N_29952,N_29585,N_29694);
or U29953 (N_29953,N_29522,N_29463);
xnor U29954 (N_29954,N_29501,N_29420);
or U29955 (N_29955,N_29632,N_29661);
or U29956 (N_29956,N_29619,N_29435);
nor U29957 (N_29957,N_29558,N_29525);
nand U29958 (N_29958,N_29634,N_29657);
nor U29959 (N_29959,N_29454,N_29418);
xnor U29960 (N_29960,N_29603,N_29696);
xnor U29961 (N_29961,N_29657,N_29407);
nor U29962 (N_29962,N_29438,N_29446);
nor U29963 (N_29963,N_29450,N_29645);
or U29964 (N_29964,N_29580,N_29413);
and U29965 (N_29965,N_29583,N_29587);
nor U29966 (N_29966,N_29634,N_29664);
nor U29967 (N_29967,N_29557,N_29611);
nor U29968 (N_29968,N_29583,N_29656);
nor U29969 (N_29969,N_29506,N_29428);
nor U29970 (N_29970,N_29413,N_29631);
xor U29971 (N_29971,N_29520,N_29627);
and U29972 (N_29972,N_29544,N_29480);
nor U29973 (N_29973,N_29579,N_29545);
xnor U29974 (N_29974,N_29490,N_29407);
nand U29975 (N_29975,N_29500,N_29560);
or U29976 (N_29976,N_29600,N_29587);
nand U29977 (N_29977,N_29675,N_29690);
nand U29978 (N_29978,N_29479,N_29598);
nand U29979 (N_29979,N_29415,N_29578);
nor U29980 (N_29980,N_29515,N_29464);
or U29981 (N_29981,N_29576,N_29656);
and U29982 (N_29982,N_29421,N_29645);
xnor U29983 (N_29983,N_29667,N_29569);
and U29984 (N_29984,N_29578,N_29489);
or U29985 (N_29985,N_29573,N_29513);
or U29986 (N_29986,N_29543,N_29662);
nor U29987 (N_29987,N_29628,N_29685);
nand U29988 (N_29988,N_29528,N_29535);
nand U29989 (N_29989,N_29660,N_29494);
nand U29990 (N_29990,N_29590,N_29489);
nor U29991 (N_29991,N_29416,N_29450);
xor U29992 (N_29992,N_29460,N_29615);
nor U29993 (N_29993,N_29408,N_29477);
and U29994 (N_29994,N_29657,N_29675);
nand U29995 (N_29995,N_29673,N_29537);
and U29996 (N_29996,N_29407,N_29561);
nand U29997 (N_29997,N_29636,N_29625);
or U29998 (N_29998,N_29681,N_29453);
and U29999 (N_29999,N_29489,N_29457);
nor UO_0 (O_0,N_29704,N_29944);
or UO_1 (O_1,N_29731,N_29709);
nand UO_2 (O_2,N_29844,N_29925);
xnor UO_3 (O_3,N_29833,N_29788);
nand UO_4 (O_4,N_29960,N_29762);
or UO_5 (O_5,N_29958,N_29931);
nor UO_6 (O_6,N_29780,N_29943);
or UO_7 (O_7,N_29898,N_29813);
nor UO_8 (O_8,N_29779,N_29798);
nor UO_9 (O_9,N_29755,N_29908);
xor UO_10 (O_10,N_29849,N_29860);
nor UO_11 (O_11,N_29838,N_29975);
and UO_12 (O_12,N_29842,N_29711);
and UO_13 (O_13,N_29982,N_29806);
and UO_14 (O_14,N_29758,N_29893);
or UO_15 (O_15,N_29812,N_29829);
or UO_16 (O_16,N_29950,N_29822);
nand UO_17 (O_17,N_29754,N_29906);
nand UO_18 (O_18,N_29912,N_29937);
nor UO_19 (O_19,N_29753,N_29840);
and UO_20 (O_20,N_29811,N_29948);
xor UO_21 (O_21,N_29719,N_29782);
xor UO_22 (O_22,N_29993,N_29740);
nand UO_23 (O_23,N_29778,N_29884);
and UO_24 (O_24,N_29909,N_29761);
nor UO_25 (O_25,N_29752,N_29737);
xnor UO_26 (O_26,N_29888,N_29859);
or UO_27 (O_27,N_29972,N_29919);
or UO_28 (O_28,N_29872,N_29820);
nand UO_29 (O_29,N_29726,N_29878);
nand UO_30 (O_30,N_29828,N_29765);
or UO_31 (O_31,N_29789,N_29713);
nand UO_32 (O_32,N_29890,N_29799);
xor UO_33 (O_33,N_29866,N_29999);
nand UO_34 (O_34,N_29924,N_29824);
xor UO_35 (O_35,N_29864,N_29868);
and UO_36 (O_36,N_29902,N_29804);
nor UO_37 (O_37,N_29932,N_29876);
xor UO_38 (O_38,N_29959,N_29730);
or UO_39 (O_39,N_29980,N_29724);
nand UO_40 (O_40,N_29708,N_29803);
nor UO_41 (O_41,N_29873,N_29769);
nand UO_42 (O_42,N_29836,N_29775);
nand UO_43 (O_43,N_29794,N_29962);
and UO_44 (O_44,N_29831,N_29827);
and UO_45 (O_45,N_29776,N_29875);
and UO_46 (O_46,N_29718,N_29716);
nand UO_47 (O_47,N_29736,N_29870);
nor UO_48 (O_48,N_29747,N_29855);
nor UO_49 (O_49,N_29979,N_29749);
nor UO_50 (O_50,N_29700,N_29945);
xnor UO_51 (O_51,N_29871,N_29946);
nor UO_52 (O_52,N_29973,N_29841);
or UO_53 (O_53,N_29926,N_29990);
xor UO_54 (O_54,N_29942,N_29797);
and UO_55 (O_55,N_29725,N_29986);
nand UO_56 (O_56,N_29846,N_29913);
nand UO_57 (O_57,N_29966,N_29857);
nor UO_58 (O_58,N_29714,N_29783);
xor UO_59 (O_59,N_29819,N_29886);
nor UO_60 (O_60,N_29941,N_29947);
nand UO_61 (O_61,N_29810,N_29781);
and UO_62 (O_62,N_29892,N_29717);
nand UO_63 (O_63,N_29984,N_29832);
xnor UO_64 (O_64,N_29922,N_29742);
nor UO_65 (O_65,N_29764,N_29785);
and UO_66 (O_66,N_29883,N_29865);
nor UO_67 (O_67,N_29706,N_29994);
nand UO_68 (O_68,N_29701,N_29996);
and UO_69 (O_69,N_29748,N_29795);
nor UO_70 (O_70,N_29796,N_29915);
nor UO_71 (O_71,N_29957,N_29792);
xor UO_72 (O_72,N_29703,N_29746);
xor UO_73 (O_73,N_29777,N_29790);
and UO_74 (O_74,N_29858,N_29715);
or UO_75 (O_75,N_29933,N_29851);
and UO_76 (O_76,N_29720,N_29784);
or UO_77 (O_77,N_29768,N_29970);
nor UO_78 (O_78,N_29904,N_29787);
nor UO_79 (O_79,N_29914,N_29817);
nor UO_80 (O_80,N_29856,N_29953);
and UO_81 (O_81,N_29826,N_29741);
and UO_82 (O_82,N_29900,N_29918);
and UO_83 (O_83,N_29845,N_29995);
xor UO_84 (O_84,N_29901,N_29939);
nand UO_85 (O_85,N_29981,N_29951);
nand UO_86 (O_86,N_29916,N_29874);
nand UO_87 (O_87,N_29744,N_29862);
or UO_88 (O_88,N_29809,N_29882);
or UO_89 (O_89,N_29802,N_29920);
nor UO_90 (O_90,N_29805,N_29935);
or UO_91 (O_91,N_29707,N_29843);
or UO_92 (O_92,N_29773,N_29881);
and UO_93 (O_93,N_29879,N_29863);
and UO_94 (O_94,N_29997,N_29978);
xor UO_95 (O_95,N_29905,N_29968);
xnor UO_96 (O_96,N_29825,N_29771);
xnor UO_97 (O_97,N_29967,N_29899);
and UO_98 (O_98,N_29848,N_29814);
or UO_99 (O_99,N_29961,N_29772);
xor UO_100 (O_100,N_29989,N_29954);
nor UO_101 (O_101,N_29853,N_29751);
nor UO_102 (O_102,N_29963,N_29885);
nand UO_103 (O_103,N_29894,N_29743);
nand UO_104 (O_104,N_29940,N_29921);
xnor UO_105 (O_105,N_29891,N_29910);
xnor UO_106 (O_106,N_29750,N_29949);
xor UO_107 (O_107,N_29930,N_29735);
nand UO_108 (O_108,N_29733,N_29985);
xnor UO_109 (O_109,N_29971,N_29834);
xnor UO_110 (O_110,N_29767,N_29964);
xor UO_111 (O_111,N_29739,N_29721);
or UO_112 (O_112,N_29821,N_29887);
and UO_113 (O_113,N_29911,N_29992);
and UO_114 (O_114,N_29705,N_29710);
or UO_115 (O_115,N_29734,N_29880);
nor UO_116 (O_116,N_29974,N_29877);
or UO_117 (O_117,N_29786,N_29907);
or UO_118 (O_118,N_29729,N_29889);
and UO_119 (O_119,N_29850,N_29998);
nor UO_120 (O_120,N_29854,N_29759);
nor UO_121 (O_121,N_29929,N_29738);
nand UO_122 (O_122,N_29861,N_29756);
nor UO_123 (O_123,N_29923,N_29983);
and UO_124 (O_124,N_29955,N_29988);
nor UO_125 (O_125,N_29732,N_29969);
nor UO_126 (O_126,N_29774,N_29852);
and UO_127 (O_127,N_29897,N_29800);
nand UO_128 (O_128,N_29928,N_29895);
and UO_129 (O_129,N_29818,N_29938);
nor UO_130 (O_130,N_29917,N_29793);
or UO_131 (O_131,N_29896,N_29965);
xor UO_132 (O_132,N_29815,N_29847);
nand UO_133 (O_133,N_29760,N_29727);
xnor UO_134 (O_134,N_29956,N_29839);
xnor UO_135 (O_135,N_29816,N_29757);
or UO_136 (O_136,N_29952,N_29987);
xnor UO_137 (O_137,N_29791,N_29977);
nand UO_138 (O_138,N_29903,N_29976);
or UO_139 (O_139,N_29770,N_29807);
or UO_140 (O_140,N_29991,N_29823);
nand UO_141 (O_141,N_29869,N_29934);
and UO_142 (O_142,N_29723,N_29830);
xnor UO_143 (O_143,N_29763,N_29712);
and UO_144 (O_144,N_29722,N_29728);
or UO_145 (O_145,N_29702,N_29808);
and UO_146 (O_146,N_29835,N_29936);
and UO_147 (O_147,N_29837,N_29745);
and UO_148 (O_148,N_29801,N_29927);
nor UO_149 (O_149,N_29766,N_29867);
xnor UO_150 (O_150,N_29801,N_29859);
or UO_151 (O_151,N_29983,N_29847);
xnor UO_152 (O_152,N_29868,N_29878);
nor UO_153 (O_153,N_29901,N_29765);
or UO_154 (O_154,N_29773,N_29987);
nand UO_155 (O_155,N_29710,N_29860);
nor UO_156 (O_156,N_29713,N_29996);
nand UO_157 (O_157,N_29993,N_29896);
or UO_158 (O_158,N_29957,N_29845);
or UO_159 (O_159,N_29838,N_29764);
nand UO_160 (O_160,N_29717,N_29858);
nor UO_161 (O_161,N_29940,N_29838);
and UO_162 (O_162,N_29933,N_29756);
nor UO_163 (O_163,N_29852,N_29930);
and UO_164 (O_164,N_29872,N_29814);
and UO_165 (O_165,N_29804,N_29769);
xor UO_166 (O_166,N_29831,N_29731);
or UO_167 (O_167,N_29906,N_29842);
or UO_168 (O_168,N_29720,N_29796);
xnor UO_169 (O_169,N_29903,N_29798);
nor UO_170 (O_170,N_29816,N_29802);
nand UO_171 (O_171,N_29858,N_29745);
or UO_172 (O_172,N_29946,N_29718);
or UO_173 (O_173,N_29722,N_29910);
and UO_174 (O_174,N_29950,N_29761);
and UO_175 (O_175,N_29810,N_29808);
and UO_176 (O_176,N_29738,N_29793);
or UO_177 (O_177,N_29975,N_29951);
or UO_178 (O_178,N_29963,N_29736);
and UO_179 (O_179,N_29948,N_29816);
and UO_180 (O_180,N_29808,N_29863);
or UO_181 (O_181,N_29731,N_29857);
and UO_182 (O_182,N_29765,N_29989);
nor UO_183 (O_183,N_29942,N_29847);
nand UO_184 (O_184,N_29864,N_29808);
and UO_185 (O_185,N_29806,N_29719);
nand UO_186 (O_186,N_29719,N_29785);
or UO_187 (O_187,N_29915,N_29788);
or UO_188 (O_188,N_29945,N_29882);
nor UO_189 (O_189,N_29919,N_29797);
nand UO_190 (O_190,N_29978,N_29981);
nor UO_191 (O_191,N_29794,N_29810);
xnor UO_192 (O_192,N_29966,N_29852);
or UO_193 (O_193,N_29965,N_29932);
and UO_194 (O_194,N_29856,N_29723);
nor UO_195 (O_195,N_29959,N_29840);
or UO_196 (O_196,N_29919,N_29944);
or UO_197 (O_197,N_29705,N_29962);
nor UO_198 (O_198,N_29914,N_29860);
and UO_199 (O_199,N_29866,N_29949);
and UO_200 (O_200,N_29800,N_29730);
nor UO_201 (O_201,N_29712,N_29982);
or UO_202 (O_202,N_29981,N_29854);
and UO_203 (O_203,N_29974,N_29847);
nor UO_204 (O_204,N_29764,N_29703);
and UO_205 (O_205,N_29757,N_29913);
xor UO_206 (O_206,N_29920,N_29875);
nor UO_207 (O_207,N_29765,N_29972);
nand UO_208 (O_208,N_29908,N_29973);
xor UO_209 (O_209,N_29756,N_29702);
or UO_210 (O_210,N_29859,N_29786);
or UO_211 (O_211,N_29804,N_29833);
xnor UO_212 (O_212,N_29919,N_29828);
and UO_213 (O_213,N_29728,N_29700);
and UO_214 (O_214,N_29876,N_29848);
and UO_215 (O_215,N_29860,N_29811);
or UO_216 (O_216,N_29885,N_29868);
nand UO_217 (O_217,N_29851,N_29958);
nor UO_218 (O_218,N_29735,N_29801);
nor UO_219 (O_219,N_29719,N_29957);
xnor UO_220 (O_220,N_29934,N_29935);
and UO_221 (O_221,N_29920,N_29899);
or UO_222 (O_222,N_29914,N_29877);
xor UO_223 (O_223,N_29702,N_29739);
nand UO_224 (O_224,N_29991,N_29779);
nand UO_225 (O_225,N_29917,N_29704);
and UO_226 (O_226,N_29715,N_29855);
nor UO_227 (O_227,N_29972,N_29922);
nand UO_228 (O_228,N_29819,N_29991);
xor UO_229 (O_229,N_29892,N_29804);
nor UO_230 (O_230,N_29729,N_29969);
or UO_231 (O_231,N_29842,N_29912);
nand UO_232 (O_232,N_29735,N_29780);
and UO_233 (O_233,N_29849,N_29955);
and UO_234 (O_234,N_29782,N_29863);
nor UO_235 (O_235,N_29785,N_29789);
nor UO_236 (O_236,N_29893,N_29870);
nor UO_237 (O_237,N_29934,N_29854);
nor UO_238 (O_238,N_29822,N_29723);
and UO_239 (O_239,N_29953,N_29841);
or UO_240 (O_240,N_29916,N_29990);
nand UO_241 (O_241,N_29991,N_29787);
nand UO_242 (O_242,N_29971,N_29794);
nor UO_243 (O_243,N_29768,N_29832);
xor UO_244 (O_244,N_29995,N_29983);
or UO_245 (O_245,N_29738,N_29797);
nor UO_246 (O_246,N_29748,N_29716);
nand UO_247 (O_247,N_29775,N_29728);
and UO_248 (O_248,N_29774,N_29835);
or UO_249 (O_249,N_29738,N_29866);
or UO_250 (O_250,N_29864,N_29993);
nand UO_251 (O_251,N_29977,N_29913);
nand UO_252 (O_252,N_29977,N_29898);
nor UO_253 (O_253,N_29821,N_29977);
xnor UO_254 (O_254,N_29947,N_29780);
xor UO_255 (O_255,N_29743,N_29773);
or UO_256 (O_256,N_29803,N_29990);
xor UO_257 (O_257,N_29893,N_29809);
xor UO_258 (O_258,N_29862,N_29998);
xor UO_259 (O_259,N_29939,N_29832);
nand UO_260 (O_260,N_29986,N_29811);
nand UO_261 (O_261,N_29736,N_29706);
nand UO_262 (O_262,N_29726,N_29894);
and UO_263 (O_263,N_29929,N_29906);
and UO_264 (O_264,N_29960,N_29963);
nor UO_265 (O_265,N_29715,N_29711);
or UO_266 (O_266,N_29707,N_29766);
nor UO_267 (O_267,N_29814,N_29818);
xor UO_268 (O_268,N_29765,N_29797);
nor UO_269 (O_269,N_29745,N_29945);
and UO_270 (O_270,N_29788,N_29920);
nor UO_271 (O_271,N_29754,N_29872);
and UO_272 (O_272,N_29735,N_29977);
and UO_273 (O_273,N_29800,N_29915);
or UO_274 (O_274,N_29779,N_29980);
nor UO_275 (O_275,N_29831,N_29713);
and UO_276 (O_276,N_29978,N_29761);
and UO_277 (O_277,N_29780,N_29727);
xor UO_278 (O_278,N_29901,N_29710);
nand UO_279 (O_279,N_29812,N_29736);
nor UO_280 (O_280,N_29943,N_29927);
nor UO_281 (O_281,N_29952,N_29827);
nand UO_282 (O_282,N_29922,N_29830);
xor UO_283 (O_283,N_29756,N_29916);
nand UO_284 (O_284,N_29988,N_29879);
nor UO_285 (O_285,N_29900,N_29917);
nor UO_286 (O_286,N_29844,N_29833);
xor UO_287 (O_287,N_29937,N_29714);
nand UO_288 (O_288,N_29761,N_29714);
and UO_289 (O_289,N_29843,N_29887);
nor UO_290 (O_290,N_29928,N_29943);
and UO_291 (O_291,N_29898,N_29938);
nand UO_292 (O_292,N_29847,N_29931);
nor UO_293 (O_293,N_29939,N_29732);
xnor UO_294 (O_294,N_29899,N_29909);
xnor UO_295 (O_295,N_29796,N_29957);
xnor UO_296 (O_296,N_29878,N_29947);
or UO_297 (O_297,N_29839,N_29818);
xnor UO_298 (O_298,N_29825,N_29716);
and UO_299 (O_299,N_29940,N_29780);
nand UO_300 (O_300,N_29935,N_29850);
xor UO_301 (O_301,N_29804,N_29956);
and UO_302 (O_302,N_29885,N_29719);
xnor UO_303 (O_303,N_29871,N_29773);
and UO_304 (O_304,N_29748,N_29722);
or UO_305 (O_305,N_29970,N_29724);
nor UO_306 (O_306,N_29716,N_29973);
and UO_307 (O_307,N_29998,N_29788);
nor UO_308 (O_308,N_29755,N_29918);
and UO_309 (O_309,N_29885,N_29863);
and UO_310 (O_310,N_29738,N_29732);
or UO_311 (O_311,N_29989,N_29754);
and UO_312 (O_312,N_29931,N_29896);
and UO_313 (O_313,N_29926,N_29721);
or UO_314 (O_314,N_29809,N_29834);
or UO_315 (O_315,N_29741,N_29849);
or UO_316 (O_316,N_29982,N_29846);
xnor UO_317 (O_317,N_29860,N_29852);
or UO_318 (O_318,N_29939,N_29903);
and UO_319 (O_319,N_29830,N_29990);
or UO_320 (O_320,N_29775,N_29866);
or UO_321 (O_321,N_29917,N_29872);
and UO_322 (O_322,N_29719,N_29833);
or UO_323 (O_323,N_29895,N_29833);
nor UO_324 (O_324,N_29864,N_29877);
and UO_325 (O_325,N_29778,N_29732);
nand UO_326 (O_326,N_29761,N_29764);
nand UO_327 (O_327,N_29986,N_29871);
and UO_328 (O_328,N_29966,N_29740);
nor UO_329 (O_329,N_29823,N_29775);
and UO_330 (O_330,N_29977,N_29808);
or UO_331 (O_331,N_29988,N_29976);
nor UO_332 (O_332,N_29750,N_29734);
and UO_333 (O_333,N_29989,N_29922);
or UO_334 (O_334,N_29870,N_29954);
or UO_335 (O_335,N_29989,N_29942);
xnor UO_336 (O_336,N_29895,N_29890);
nor UO_337 (O_337,N_29912,N_29897);
nand UO_338 (O_338,N_29986,N_29915);
nand UO_339 (O_339,N_29754,N_29700);
and UO_340 (O_340,N_29779,N_29753);
nand UO_341 (O_341,N_29855,N_29871);
and UO_342 (O_342,N_29814,N_29877);
xnor UO_343 (O_343,N_29787,N_29722);
and UO_344 (O_344,N_29731,N_29701);
and UO_345 (O_345,N_29917,N_29953);
or UO_346 (O_346,N_29763,N_29981);
xnor UO_347 (O_347,N_29878,N_29742);
xnor UO_348 (O_348,N_29804,N_29938);
nand UO_349 (O_349,N_29860,N_29832);
and UO_350 (O_350,N_29791,N_29869);
xnor UO_351 (O_351,N_29951,N_29865);
xor UO_352 (O_352,N_29878,N_29705);
nor UO_353 (O_353,N_29971,N_29923);
nand UO_354 (O_354,N_29983,N_29967);
xor UO_355 (O_355,N_29785,N_29753);
nand UO_356 (O_356,N_29771,N_29977);
nor UO_357 (O_357,N_29799,N_29943);
or UO_358 (O_358,N_29701,N_29995);
and UO_359 (O_359,N_29857,N_29793);
nor UO_360 (O_360,N_29952,N_29851);
xor UO_361 (O_361,N_29964,N_29911);
or UO_362 (O_362,N_29947,N_29844);
nor UO_363 (O_363,N_29939,N_29934);
and UO_364 (O_364,N_29814,N_29825);
nor UO_365 (O_365,N_29782,N_29803);
or UO_366 (O_366,N_29848,N_29942);
xnor UO_367 (O_367,N_29841,N_29942);
xor UO_368 (O_368,N_29984,N_29882);
nor UO_369 (O_369,N_29722,N_29977);
or UO_370 (O_370,N_29749,N_29956);
nor UO_371 (O_371,N_29825,N_29752);
nand UO_372 (O_372,N_29790,N_29805);
nor UO_373 (O_373,N_29760,N_29834);
nand UO_374 (O_374,N_29908,N_29914);
xor UO_375 (O_375,N_29997,N_29825);
and UO_376 (O_376,N_29707,N_29929);
nor UO_377 (O_377,N_29998,N_29869);
and UO_378 (O_378,N_29790,N_29990);
or UO_379 (O_379,N_29893,N_29726);
nand UO_380 (O_380,N_29874,N_29726);
or UO_381 (O_381,N_29977,N_29803);
or UO_382 (O_382,N_29759,N_29897);
and UO_383 (O_383,N_29746,N_29819);
nand UO_384 (O_384,N_29983,N_29896);
nand UO_385 (O_385,N_29709,N_29782);
or UO_386 (O_386,N_29955,N_29954);
nand UO_387 (O_387,N_29901,N_29832);
xor UO_388 (O_388,N_29870,N_29940);
or UO_389 (O_389,N_29705,N_29733);
or UO_390 (O_390,N_29965,N_29845);
nor UO_391 (O_391,N_29701,N_29781);
nor UO_392 (O_392,N_29795,N_29902);
xor UO_393 (O_393,N_29970,N_29995);
xnor UO_394 (O_394,N_29700,N_29805);
nand UO_395 (O_395,N_29747,N_29981);
nand UO_396 (O_396,N_29854,N_29722);
nand UO_397 (O_397,N_29728,N_29901);
xor UO_398 (O_398,N_29985,N_29713);
nor UO_399 (O_399,N_29819,N_29930);
nand UO_400 (O_400,N_29706,N_29861);
and UO_401 (O_401,N_29815,N_29785);
xnor UO_402 (O_402,N_29808,N_29849);
and UO_403 (O_403,N_29773,N_29994);
and UO_404 (O_404,N_29936,N_29932);
and UO_405 (O_405,N_29978,N_29949);
nor UO_406 (O_406,N_29946,N_29712);
or UO_407 (O_407,N_29865,N_29939);
xor UO_408 (O_408,N_29845,N_29945);
or UO_409 (O_409,N_29858,N_29881);
or UO_410 (O_410,N_29747,N_29826);
or UO_411 (O_411,N_29945,N_29980);
and UO_412 (O_412,N_29756,N_29873);
or UO_413 (O_413,N_29948,N_29792);
nand UO_414 (O_414,N_29917,N_29857);
nor UO_415 (O_415,N_29848,N_29962);
nor UO_416 (O_416,N_29859,N_29717);
or UO_417 (O_417,N_29738,N_29850);
or UO_418 (O_418,N_29932,N_29822);
nor UO_419 (O_419,N_29996,N_29774);
or UO_420 (O_420,N_29845,N_29747);
and UO_421 (O_421,N_29730,N_29734);
and UO_422 (O_422,N_29795,N_29772);
xnor UO_423 (O_423,N_29963,N_29715);
or UO_424 (O_424,N_29951,N_29791);
xor UO_425 (O_425,N_29954,N_29826);
xnor UO_426 (O_426,N_29956,N_29713);
and UO_427 (O_427,N_29900,N_29701);
or UO_428 (O_428,N_29702,N_29834);
nor UO_429 (O_429,N_29884,N_29768);
or UO_430 (O_430,N_29764,N_29927);
and UO_431 (O_431,N_29915,N_29855);
xor UO_432 (O_432,N_29818,N_29861);
nand UO_433 (O_433,N_29784,N_29755);
and UO_434 (O_434,N_29842,N_29941);
and UO_435 (O_435,N_29856,N_29963);
xor UO_436 (O_436,N_29827,N_29826);
nand UO_437 (O_437,N_29849,N_29884);
nor UO_438 (O_438,N_29858,N_29723);
xor UO_439 (O_439,N_29967,N_29869);
xor UO_440 (O_440,N_29907,N_29998);
nor UO_441 (O_441,N_29960,N_29922);
nor UO_442 (O_442,N_29909,N_29778);
and UO_443 (O_443,N_29806,N_29906);
and UO_444 (O_444,N_29890,N_29914);
and UO_445 (O_445,N_29896,N_29806);
nand UO_446 (O_446,N_29750,N_29849);
and UO_447 (O_447,N_29831,N_29789);
nor UO_448 (O_448,N_29713,N_29810);
xnor UO_449 (O_449,N_29781,N_29988);
xnor UO_450 (O_450,N_29794,N_29891);
or UO_451 (O_451,N_29932,N_29927);
nor UO_452 (O_452,N_29782,N_29843);
nand UO_453 (O_453,N_29989,N_29843);
or UO_454 (O_454,N_29824,N_29826);
or UO_455 (O_455,N_29857,N_29724);
and UO_456 (O_456,N_29711,N_29815);
nand UO_457 (O_457,N_29964,N_29806);
or UO_458 (O_458,N_29878,N_29930);
xor UO_459 (O_459,N_29772,N_29784);
or UO_460 (O_460,N_29762,N_29908);
or UO_461 (O_461,N_29800,N_29795);
xnor UO_462 (O_462,N_29869,N_29948);
and UO_463 (O_463,N_29974,N_29776);
xnor UO_464 (O_464,N_29831,N_29808);
nand UO_465 (O_465,N_29907,N_29752);
or UO_466 (O_466,N_29714,N_29817);
nand UO_467 (O_467,N_29732,N_29957);
nor UO_468 (O_468,N_29846,N_29709);
nand UO_469 (O_469,N_29799,N_29708);
xnor UO_470 (O_470,N_29907,N_29928);
nor UO_471 (O_471,N_29742,N_29975);
nand UO_472 (O_472,N_29947,N_29894);
or UO_473 (O_473,N_29840,N_29905);
nand UO_474 (O_474,N_29714,N_29727);
xor UO_475 (O_475,N_29772,N_29767);
or UO_476 (O_476,N_29808,N_29820);
nand UO_477 (O_477,N_29743,N_29724);
and UO_478 (O_478,N_29955,N_29990);
or UO_479 (O_479,N_29803,N_29925);
nand UO_480 (O_480,N_29859,N_29705);
nand UO_481 (O_481,N_29759,N_29894);
nand UO_482 (O_482,N_29912,N_29821);
nand UO_483 (O_483,N_29968,N_29753);
nand UO_484 (O_484,N_29870,N_29714);
nor UO_485 (O_485,N_29844,N_29877);
nand UO_486 (O_486,N_29907,N_29929);
or UO_487 (O_487,N_29942,N_29897);
nor UO_488 (O_488,N_29821,N_29730);
and UO_489 (O_489,N_29874,N_29952);
and UO_490 (O_490,N_29847,N_29949);
and UO_491 (O_491,N_29713,N_29995);
and UO_492 (O_492,N_29745,N_29965);
nand UO_493 (O_493,N_29891,N_29877);
and UO_494 (O_494,N_29717,N_29702);
nand UO_495 (O_495,N_29795,N_29904);
and UO_496 (O_496,N_29740,N_29841);
nor UO_497 (O_497,N_29812,N_29820);
or UO_498 (O_498,N_29705,N_29813);
or UO_499 (O_499,N_29871,N_29896);
nor UO_500 (O_500,N_29919,N_29867);
nor UO_501 (O_501,N_29901,N_29872);
xor UO_502 (O_502,N_29926,N_29880);
xnor UO_503 (O_503,N_29756,N_29815);
nand UO_504 (O_504,N_29994,N_29735);
or UO_505 (O_505,N_29927,N_29939);
xor UO_506 (O_506,N_29796,N_29848);
and UO_507 (O_507,N_29929,N_29729);
or UO_508 (O_508,N_29890,N_29748);
and UO_509 (O_509,N_29733,N_29791);
nor UO_510 (O_510,N_29751,N_29918);
nor UO_511 (O_511,N_29876,N_29788);
nor UO_512 (O_512,N_29741,N_29728);
nor UO_513 (O_513,N_29983,N_29956);
and UO_514 (O_514,N_29913,N_29876);
xnor UO_515 (O_515,N_29726,N_29748);
xnor UO_516 (O_516,N_29891,N_29977);
and UO_517 (O_517,N_29951,N_29992);
nand UO_518 (O_518,N_29794,N_29929);
and UO_519 (O_519,N_29912,N_29928);
xnor UO_520 (O_520,N_29843,N_29723);
and UO_521 (O_521,N_29871,N_29977);
or UO_522 (O_522,N_29788,N_29898);
or UO_523 (O_523,N_29898,N_29868);
xnor UO_524 (O_524,N_29902,N_29843);
or UO_525 (O_525,N_29807,N_29880);
nand UO_526 (O_526,N_29843,N_29954);
and UO_527 (O_527,N_29937,N_29996);
xnor UO_528 (O_528,N_29854,N_29985);
nand UO_529 (O_529,N_29987,N_29957);
nor UO_530 (O_530,N_29952,N_29924);
nor UO_531 (O_531,N_29886,N_29807);
nor UO_532 (O_532,N_29909,N_29750);
nor UO_533 (O_533,N_29878,N_29938);
or UO_534 (O_534,N_29871,N_29851);
or UO_535 (O_535,N_29938,N_29925);
nor UO_536 (O_536,N_29858,N_29887);
nand UO_537 (O_537,N_29837,N_29715);
nor UO_538 (O_538,N_29971,N_29884);
nor UO_539 (O_539,N_29800,N_29804);
nand UO_540 (O_540,N_29792,N_29807);
or UO_541 (O_541,N_29931,N_29992);
or UO_542 (O_542,N_29706,N_29742);
or UO_543 (O_543,N_29721,N_29876);
or UO_544 (O_544,N_29881,N_29862);
or UO_545 (O_545,N_29708,N_29974);
or UO_546 (O_546,N_29824,N_29771);
nor UO_547 (O_547,N_29769,N_29850);
and UO_548 (O_548,N_29868,N_29881);
nand UO_549 (O_549,N_29797,N_29715);
and UO_550 (O_550,N_29764,N_29780);
nand UO_551 (O_551,N_29908,N_29834);
nand UO_552 (O_552,N_29782,N_29922);
or UO_553 (O_553,N_29762,N_29754);
nor UO_554 (O_554,N_29774,N_29946);
nand UO_555 (O_555,N_29998,N_29837);
and UO_556 (O_556,N_29857,N_29848);
and UO_557 (O_557,N_29706,N_29883);
nand UO_558 (O_558,N_29939,N_29771);
or UO_559 (O_559,N_29757,N_29730);
or UO_560 (O_560,N_29865,N_29905);
nor UO_561 (O_561,N_29898,N_29761);
and UO_562 (O_562,N_29960,N_29975);
nor UO_563 (O_563,N_29832,N_29941);
nand UO_564 (O_564,N_29841,N_29882);
nor UO_565 (O_565,N_29709,N_29903);
and UO_566 (O_566,N_29756,N_29996);
or UO_567 (O_567,N_29711,N_29953);
nand UO_568 (O_568,N_29954,N_29848);
or UO_569 (O_569,N_29820,N_29952);
and UO_570 (O_570,N_29910,N_29816);
nor UO_571 (O_571,N_29953,N_29846);
nand UO_572 (O_572,N_29876,N_29837);
xnor UO_573 (O_573,N_29789,N_29704);
nor UO_574 (O_574,N_29903,N_29979);
nor UO_575 (O_575,N_29758,N_29792);
or UO_576 (O_576,N_29782,N_29969);
xor UO_577 (O_577,N_29998,N_29796);
or UO_578 (O_578,N_29893,N_29983);
nand UO_579 (O_579,N_29733,N_29702);
nor UO_580 (O_580,N_29786,N_29718);
nor UO_581 (O_581,N_29941,N_29705);
and UO_582 (O_582,N_29921,N_29932);
nor UO_583 (O_583,N_29918,N_29773);
nand UO_584 (O_584,N_29762,N_29746);
or UO_585 (O_585,N_29703,N_29931);
xnor UO_586 (O_586,N_29843,N_29998);
xor UO_587 (O_587,N_29985,N_29772);
nor UO_588 (O_588,N_29722,N_29997);
and UO_589 (O_589,N_29964,N_29932);
or UO_590 (O_590,N_29962,N_29877);
or UO_591 (O_591,N_29876,N_29944);
nand UO_592 (O_592,N_29829,N_29713);
nand UO_593 (O_593,N_29968,N_29770);
xnor UO_594 (O_594,N_29777,N_29765);
xor UO_595 (O_595,N_29738,N_29781);
nand UO_596 (O_596,N_29753,N_29951);
nor UO_597 (O_597,N_29840,N_29862);
nand UO_598 (O_598,N_29823,N_29875);
and UO_599 (O_599,N_29854,N_29778);
nand UO_600 (O_600,N_29773,N_29944);
nor UO_601 (O_601,N_29910,N_29740);
or UO_602 (O_602,N_29743,N_29909);
and UO_603 (O_603,N_29798,N_29799);
xor UO_604 (O_604,N_29737,N_29805);
and UO_605 (O_605,N_29794,N_29935);
nand UO_606 (O_606,N_29866,N_29867);
nand UO_607 (O_607,N_29963,N_29753);
or UO_608 (O_608,N_29922,N_29894);
xor UO_609 (O_609,N_29902,N_29891);
nor UO_610 (O_610,N_29961,N_29729);
nor UO_611 (O_611,N_29971,N_29906);
nand UO_612 (O_612,N_29788,N_29827);
and UO_613 (O_613,N_29772,N_29769);
or UO_614 (O_614,N_29912,N_29975);
and UO_615 (O_615,N_29929,N_29715);
or UO_616 (O_616,N_29743,N_29842);
nor UO_617 (O_617,N_29891,N_29784);
nor UO_618 (O_618,N_29874,N_29739);
xnor UO_619 (O_619,N_29822,N_29826);
nor UO_620 (O_620,N_29932,N_29835);
or UO_621 (O_621,N_29929,N_29991);
xnor UO_622 (O_622,N_29866,N_29900);
or UO_623 (O_623,N_29874,N_29868);
or UO_624 (O_624,N_29731,N_29844);
or UO_625 (O_625,N_29889,N_29888);
or UO_626 (O_626,N_29919,N_29898);
or UO_627 (O_627,N_29868,N_29816);
or UO_628 (O_628,N_29956,N_29760);
nor UO_629 (O_629,N_29855,N_29884);
nor UO_630 (O_630,N_29934,N_29864);
and UO_631 (O_631,N_29921,N_29799);
and UO_632 (O_632,N_29802,N_29706);
xor UO_633 (O_633,N_29852,N_29936);
nor UO_634 (O_634,N_29858,N_29975);
nor UO_635 (O_635,N_29842,N_29997);
nand UO_636 (O_636,N_29777,N_29921);
nand UO_637 (O_637,N_29793,N_29790);
xnor UO_638 (O_638,N_29940,N_29881);
nand UO_639 (O_639,N_29995,N_29762);
xnor UO_640 (O_640,N_29872,N_29813);
or UO_641 (O_641,N_29885,N_29750);
and UO_642 (O_642,N_29770,N_29862);
and UO_643 (O_643,N_29933,N_29716);
nor UO_644 (O_644,N_29823,N_29970);
xnor UO_645 (O_645,N_29972,N_29981);
xnor UO_646 (O_646,N_29920,N_29827);
or UO_647 (O_647,N_29850,N_29786);
nor UO_648 (O_648,N_29823,N_29891);
nor UO_649 (O_649,N_29731,N_29752);
nand UO_650 (O_650,N_29914,N_29955);
nand UO_651 (O_651,N_29928,N_29847);
and UO_652 (O_652,N_29711,N_29724);
xor UO_653 (O_653,N_29778,N_29890);
and UO_654 (O_654,N_29817,N_29801);
or UO_655 (O_655,N_29808,N_29884);
nand UO_656 (O_656,N_29789,N_29968);
and UO_657 (O_657,N_29790,N_29742);
xnor UO_658 (O_658,N_29918,N_29799);
xnor UO_659 (O_659,N_29748,N_29827);
xnor UO_660 (O_660,N_29879,N_29894);
nor UO_661 (O_661,N_29977,N_29750);
or UO_662 (O_662,N_29874,N_29736);
and UO_663 (O_663,N_29944,N_29815);
or UO_664 (O_664,N_29861,N_29870);
or UO_665 (O_665,N_29968,N_29728);
and UO_666 (O_666,N_29772,N_29990);
nor UO_667 (O_667,N_29949,N_29852);
xnor UO_668 (O_668,N_29994,N_29710);
nor UO_669 (O_669,N_29945,N_29772);
and UO_670 (O_670,N_29701,N_29929);
and UO_671 (O_671,N_29775,N_29799);
and UO_672 (O_672,N_29892,N_29807);
nor UO_673 (O_673,N_29894,N_29891);
nor UO_674 (O_674,N_29829,N_29860);
nor UO_675 (O_675,N_29946,N_29924);
xnor UO_676 (O_676,N_29727,N_29813);
nand UO_677 (O_677,N_29802,N_29767);
nor UO_678 (O_678,N_29966,N_29755);
and UO_679 (O_679,N_29805,N_29836);
nand UO_680 (O_680,N_29712,N_29920);
nor UO_681 (O_681,N_29857,N_29739);
and UO_682 (O_682,N_29735,N_29830);
nand UO_683 (O_683,N_29730,N_29802);
or UO_684 (O_684,N_29937,N_29755);
and UO_685 (O_685,N_29997,N_29737);
xnor UO_686 (O_686,N_29827,N_29823);
xnor UO_687 (O_687,N_29812,N_29822);
and UO_688 (O_688,N_29840,N_29974);
nand UO_689 (O_689,N_29779,N_29748);
xnor UO_690 (O_690,N_29930,N_29706);
xnor UO_691 (O_691,N_29869,N_29925);
and UO_692 (O_692,N_29914,N_29850);
and UO_693 (O_693,N_29983,N_29864);
nor UO_694 (O_694,N_29776,N_29817);
and UO_695 (O_695,N_29914,N_29905);
or UO_696 (O_696,N_29939,N_29918);
or UO_697 (O_697,N_29858,N_29754);
or UO_698 (O_698,N_29822,N_29730);
and UO_699 (O_699,N_29706,N_29817);
xnor UO_700 (O_700,N_29973,N_29799);
and UO_701 (O_701,N_29843,N_29959);
nand UO_702 (O_702,N_29981,N_29949);
nor UO_703 (O_703,N_29976,N_29874);
nand UO_704 (O_704,N_29840,N_29846);
nor UO_705 (O_705,N_29820,N_29815);
nor UO_706 (O_706,N_29735,N_29729);
xor UO_707 (O_707,N_29954,N_29951);
nand UO_708 (O_708,N_29904,N_29763);
xor UO_709 (O_709,N_29759,N_29776);
nor UO_710 (O_710,N_29703,N_29769);
xor UO_711 (O_711,N_29826,N_29866);
nand UO_712 (O_712,N_29862,N_29738);
xnor UO_713 (O_713,N_29860,N_29788);
xor UO_714 (O_714,N_29810,N_29787);
xnor UO_715 (O_715,N_29930,N_29705);
nor UO_716 (O_716,N_29948,N_29804);
or UO_717 (O_717,N_29855,N_29996);
nand UO_718 (O_718,N_29751,N_29950);
nor UO_719 (O_719,N_29717,N_29928);
nand UO_720 (O_720,N_29905,N_29951);
and UO_721 (O_721,N_29915,N_29824);
nand UO_722 (O_722,N_29972,N_29812);
xnor UO_723 (O_723,N_29798,N_29899);
nand UO_724 (O_724,N_29736,N_29884);
or UO_725 (O_725,N_29879,N_29848);
xor UO_726 (O_726,N_29917,N_29893);
nor UO_727 (O_727,N_29888,N_29770);
or UO_728 (O_728,N_29842,N_29781);
xor UO_729 (O_729,N_29975,N_29752);
xnor UO_730 (O_730,N_29965,N_29835);
xor UO_731 (O_731,N_29822,N_29746);
or UO_732 (O_732,N_29920,N_29893);
nand UO_733 (O_733,N_29961,N_29842);
and UO_734 (O_734,N_29840,N_29773);
and UO_735 (O_735,N_29767,N_29949);
nor UO_736 (O_736,N_29813,N_29759);
and UO_737 (O_737,N_29917,N_29815);
nor UO_738 (O_738,N_29778,N_29948);
and UO_739 (O_739,N_29843,N_29762);
xnor UO_740 (O_740,N_29920,N_29757);
and UO_741 (O_741,N_29812,N_29920);
and UO_742 (O_742,N_29746,N_29975);
and UO_743 (O_743,N_29923,N_29710);
xnor UO_744 (O_744,N_29894,N_29930);
and UO_745 (O_745,N_29890,N_29949);
and UO_746 (O_746,N_29835,N_29756);
nor UO_747 (O_747,N_29710,N_29769);
nand UO_748 (O_748,N_29743,N_29720);
or UO_749 (O_749,N_29943,N_29883);
nor UO_750 (O_750,N_29930,N_29814);
or UO_751 (O_751,N_29750,N_29844);
nand UO_752 (O_752,N_29747,N_29960);
nor UO_753 (O_753,N_29940,N_29990);
and UO_754 (O_754,N_29768,N_29876);
and UO_755 (O_755,N_29779,N_29966);
xor UO_756 (O_756,N_29802,N_29919);
nand UO_757 (O_757,N_29920,N_29832);
nand UO_758 (O_758,N_29914,N_29779);
and UO_759 (O_759,N_29874,N_29773);
nor UO_760 (O_760,N_29873,N_29941);
nor UO_761 (O_761,N_29860,N_29963);
and UO_762 (O_762,N_29815,N_29732);
xnor UO_763 (O_763,N_29752,N_29864);
nand UO_764 (O_764,N_29907,N_29804);
and UO_765 (O_765,N_29897,N_29741);
xnor UO_766 (O_766,N_29771,N_29912);
xnor UO_767 (O_767,N_29942,N_29727);
nor UO_768 (O_768,N_29953,N_29807);
xnor UO_769 (O_769,N_29965,N_29921);
nor UO_770 (O_770,N_29933,N_29889);
nand UO_771 (O_771,N_29746,N_29976);
xor UO_772 (O_772,N_29957,N_29816);
nand UO_773 (O_773,N_29983,N_29860);
nand UO_774 (O_774,N_29748,N_29970);
nor UO_775 (O_775,N_29988,N_29875);
or UO_776 (O_776,N_29860,N_29793);
xnor UO_777 (O_777,N_29761,N_29947);
and UO_778 (O_778,N_29812,N_29705);
or UO_779 (O_779,N_29740,N_29721);
xnor UO_780 (O_780,N_29867,N_29873);
xor UO_781 (O_781,N_29984,N_29952);
and UO_782 (O_782,N_29733,N_29958);
nand UO_783 (O_783,N_29965,N_29721);
nand UO_784 (O_784,N_29885,N_29996);
nor UO_785 (O_785,N_29886,N_29963);
nor UO_786 (O_786,N_29924,N_29722);
and UO_787 (O_787,N_29820,N_29836);
nand UO_788 (O_788,N_29825,N_29987);
nand UO_789 (O_789,N_29988,N_29821);
nor UO_790 (O_790,N_29983,N_29856);
nor UO_791 (O_791,N_29888,N_29764);
nand UO_792 (O_792,N_29812,N_29922);
or UO_793 (O_793,N_29743,N_29916);
or UO_794 (O_794,N_29927,N_29969);
nand UO_795 (O_795,N_29706,N_29984);
or UO_796 (O_796,N_29868,N_29929);
or UO_797 (O_797,N_29710,N_29770);
xor UO_798 (O_798,N_29771,N_29911);
xor UO_799 (O_799,N_29709,N_29712);
nand UO_800 (O_800,N_29710,N_29963);
xnor UO_801 (O_801,N_29957,N_29836);
xnor UO_802 (O_802,N_29735,N_29940);
and UO_803 (O_803,N_29788,N_29906);
and UO_804 (O_804,N_29719,N_29998);
and UO_805 (O_805,N_29966,N_29911);
nand UO_806 (O_806,N_29848,N_29806);
and UO_807 (O_807,N_29995,N_29803);
or UO_808 (O_808,N_29932,N_29875);
xor UO_809 (O_809,N_29935,N_29965);
and UO_810 (O_810,N_29747,N_29912);
nor UO_811 (O_811,N_29989,N_29957);
and UO_812 (O_812,N_29843,N_29962);
nand UO_813 (O_813,N_29746,N_29962);
and UO_814 (O_814,N_29705,N_29796);
xor UO_815 (O_815,N_29722,N_29881);
nor UO_816 (O_816,N_29833,N_29821);
or UO_817 (O_817,N_29914,N_29799);
xor UO_818 (O_818,N_29909,N_29718);
xor UO_819 (O_819,N_29804,N_29771);
or UO_820 (O_820,N_29721,N_29786);
nand UO_821 (O_821,N_29911,N_29934);
and UO_822 (O_822,N_29764,N_29788);
and UO_823 (O_823,N_29950,N_29858);
nor UO_824 (O_824,N_29702,N_29809);
nor UO_825 (O_825,N_29807,N_29959);
or UO_826 (O_826,N_29883,N_29745);
xnor UO_827 (O_827,N_29995,N_29825);
xnor UO_828 (O_828,N_29766,N_29776);
xnor UO_829 (O_829,N_29723,N_29847);
and UO_830 (O_830,N_29854,N_29756);
xor UO_831 (O_831,N_29862,N_29980);
and UO_832 (O_832,N_29788,N_29951);
or UO_833 (O_833,N_29982,N_29753);
nor UO_834 (O_834,N_29728,N_29768);
and UO_835 (O_835,N_29926,N_29774);
nor UO_836 (O_836,N_29730,N_29852);
nor UO_837 (O_837,N_29770,N_29925);
nor UO_838 (O_838,N_29817,N_29904);
nand UO_839 (O_839,N_29825,N_29971);
and UO_840 (O_840,N_29833,N_29742);
and UO_841 (O_841,N_29709,N_29974);
xor UO_842 (O_842,N_29800,N_29901);
or UO_843 (O_843,N_29704,N_29962);
or UO_844 (O_844,N_29938,N_29852);
xor UO_845 (O_845,N_29938,N_29814);
nand UO_846 (O_846,N_29820,N_29921);
xnor UO_847 (O_847,N_29701,N_29708);
xor UO_848 (O_848,N_29990,N_29902);
and UO_849 (O_849,N_29964,N_29883);
or UO_850 (O_850,N_29979,N_29808);
nor UO_851 (O_851,N_29820,N_29971);
xor UO_852 (O_852,N_29856,N_29911);
and UO_853 (O_853,N_29870,N_29992);
and UO_854 (O_854,N_29838,N_29725);
or UO_855 (O_855,N_29843,N_29788);
nor UO_856 (O_856,N_29771,N_29941);
xor UO_857 (O_857,N_29804,N_29789);
and UO_858 (O_858,N_29706,N_29871);
nand UO_859 (O_859,N_29808,N_29969);
or UO_860 (O_860,N_29790,N_29959);
nand UO_861 (O_861,N_29913,N_29721);
nor UO_862 (O_862,N_29734,N_29869);
nor UO_863 (O_863,N_29953,N_29721);
and UO_864 (O_864,N_29866,N_29816);
xor UO_865 (O_865,N_29925,N_29754);
nor UO_866 (O_866,N_29828,N_29963);
and UO_867 (O_867,N_29871,N_29988);
nor UO_868 (O_868,N_29804,N_29744);
xnor UO_869 (O_869,N_29973,N_29807);
nor UO_870 (O_870,N_29929,N_29824);
xor UO_871 (O_871,N_29979,N_29977);
nor UO_872 (O_872,N_29727,N_29902);
or UO_873 (O_873,N_29880,N_29906);
xor UO_874 (O_874,N_29954,N_29705);
nand UO_875 (O_875,N_29954,N_29869);
nand UO_876 (O_876,N_29880,N_29905);
and UO_877 (O_877,N_29721,N_29796);
nor UO_878 (O_878,N_29939,N_29899);
and UO_879 (O_879,N_29755,N_29960);
nand UO_880 (O_880,N_29913,N_29804);
or UO_881 (O_881,N_29764,N_29859);
and UO_882 (O_882,N_29790,N_29713);
xor UO_883 (O_883,N_29911,N_29958);
nand UO_884 (O_884,N_29724,N_29745);
nand UO_885 (O_885,N_29811,N_29872);
nor UO_886 (O_886,N_29712,N_29737);
nor UO_887 (O_887,N_29765,N_29830);
xor UO_888 (O_888,N_29933,N_29840);
nor UO_889 (O_889,N_29937,N_29789);
or UO_890 (O_890,N_29915,N_29913);
or UO_891 (O_891,N_29821,N_29940);
and UO_892 (O_892,N_29956,N_29811);
or UO_893 (O_893,N_29776,N_29816);
and UO_894 (O_894,N_29791,N_29904);
xnor UO_895 (O_895,N_29736,N_29735);
nor UO_896 (O_896,N_29729,N_29881);
nand UO_897 (O_897,N_29844,N_29933);
or UO_898 (O_898,N_29729,N_29915);
or UO_899 (O_899,N_29806,N_29722);
nand UO_900 (O_900,N_29855,N_29778);
and UO_901 (O_901,N_29916,N_29999);
and UO_902 (O_902,N_29817,N_29805);
or UO_903 (O_903,N_29751,N_29937);
xnor UO_904 (O_904,N_29805,N_29971);
nand UO_905 (O_905,N_29849,N_29752);
xor UO_906 (O_906,N_29759,N_29994);
nand UO_907 (O_907,N_29961,N_29797);
and UO_908 (O_908,N_29827,N_29885);
nand UO_909 (O_909,N_29750,N_29946);
xnor UO_910 (O_910,N_29709,N_29916);
nand UO_911 (O_911,N_29891,N_29801);
and UO_912 (O_912,N_29751,N_29928);
nor UO_913 (O_913,N_29920,N_29828);
nand UO_914 (O_914,N_29898,N_29787);
and UO_915 (O_915,N_29847,N_29906);
or UO_916 (O_916,N_29987,N_29889);
nand UO_917 (O_917,N_29725,N_29782);
xnor UO_918 (O_918,N_29914,N_29846);
nand UO_919 (O_919,N_29912,N_29715);
xor UO_920 (O_920,N_29827,N_29939);
nor UO_921 (O_921,N_29920,N_29992);
nand UO_922 (O_922,N_29985,N_29864);
nand UO_923 (O_923,N_29899,N_29755);
nand UO_924 (O_924,N_29946,N_29925);
or UO_925 (O_925,N_29851,N_29870);
or UO_926 (O_926,N_29742,N_29837);
or UO_927 (O_927,N_29808,N_29704);
or UO_928 (O_928,N_29838,N_29700);
nand UO_929 (O_929,N_29935,N_29861);
nor UO_930 (O_930,N_29958,N_29814);
and UO_931 (O_931,N_29866,N_29878);
nor UO_932 (O_932,N_29916,N_29864);
nand UO_933 (O_933,N_29811,N_29749);
or UO_934 (O_934,N_29750,N_29724);
or UO_935 (O_935,N_29786,N_29926);
nand UO_936 (O_936,N_29876,N_29751);
nand UO_937 (O_937,N_29899,N_29803);
and UO_938 (O_938,N_29885,N_29758);
nand UO_939 (O_939,N_29950,N_29724);
and UO_940 (O_940,N_29930,N_29864);
xnor UO_941 (O_941,N_29833,N_29842);
xnor UO_942 (O_942,N_29841,N_29971);
xor UO_943 (O_943,N_29784,N_29952);
or UO_944 (O_944,N_29771,N_29997);
and UO_945 (O_945,N_29903,N_29850);
and UO_946 (O_946,N_29745,N_29931);
and UO_947 (O_947,N_29973,N_29752);
or UO_948 (O_948,N_29716,N_29703);
and UO_949 (O_949,N_29990,N_29900);
nand UO_950 (O_950,N_29885,N_29979);
nor UO_951 (O_951,N_29970,N_29877);
or UO_952 (O_952,N_29754,N_29999);
nand UO_953 (O_953,N_29952,N_29772);
nand UO_954 (O_954,N_29870,N_29982);
xor UO_955 (O_955,N_29948,N_29747);
nor UO_956 (O_956,N_29720,N_29828);
nand UO_957 (O_957,N_29971,N_29827);
and UO_958 (O_958,N_29897,N_29731);
xnor UO_959 (O_959,N_29719,N_29950);
xor UO_960 (O_960,N_29730,N_29909);
xnor UO_961 (O_961,N_29778,N_29746);
or UO_962 (O_962,N_29860,N_29993);
xor UO_963 (O_963,N_29871,N_29771);
and UO_964 (O_964,N_29966,N_29965);
or UO_965 (O_965,N_29820,N_29731);
nor UO_966 (O_966,N_29831,N_29848);
nand UO_967 (O_967,N_29922,N_29788);
nand UO_968 (O_968,N_29744,N_29746);
or UO_969 (O_969,N_29711,N_29855);
nor UO_970 (O_970,N_29792,N_29719);
and UO_971 (O_971,N_29930,N_29958);
or UO_972 (O_972,N_29777,N_29945);
xnor UO_973 (O_973,N_29927,N_29810);
and UO_974 (O_974,N_29933,N_29706);
or UO_975 (O_975,N_29826,N_29701);
xnor UO_976 (O_976,N_29997,N_29766);
xor UO_977 (O_977,N_29705,N_29909);
nor UO_978 (O_978,N_29866,N_29899);
xnor UO_979 (O_979,N_29957,N_29932);
or UO_980 (O_980,N_29911,N_29768);
nor UO_981 (O_981,N_29997,N_29913);
nor UO_982 (O_982,N_29861,N_29933);
and UO_983 (O_983,N_29959,N_29861);
and UO_984 (O_984,N_29988,N_29985);
or UO_985 (O_985,N_29843,N_29758);
nand UO_986 (O_986,N_29809,N_29963);
xnor UO_987 (O_987,N_29880,N_29762);
xor UO_988 (O_988,N_29932,N_29796);
xor UO_989 (O_989,N_29855,N_29852);
nand UO_990 (O_990,N_29890,N_29867);
nor UO_991 (O_991,N_29857,N_29845);
and UO_992 (O_992,N_29838,N_29826);
or UO_993 (O_993,N_29721,N_29942);
nand UO_994 (O_994,N_29811,N_29929);
and UO_995 (O_995,N_29938,N_29776);
xor UO_996 (O_996,N_29839,N_29947);
xor UO_997 (O_997,N_29878,N_29881);
nor UO_998 (O_998,N_29909,N_29789);
nor UO_999 (O_999,N_29826,N_29781);
or UO_1000 (O_1000,N_29968,N_29861);
or UO_1001 (O_1001,N_29861,N_29956);
xor UO_1002 (O_1002,N_29844,N_29797);
and UO_1003 (O_1003,N_29825,N_29883);
or UO_1004 (O_1004,N_29705,N_29926);
nand UO_1005 (O_1005,N_29875,N_29903);
xor UO_1006 (O_1006,N_29774,N_29791);
nand UO_1007 (O_1007,N_29890,N_29779);
nor UO_1008 (O_1008,N_29809,N_29940);
xnor UO_1009 (O_1009,N_29913,N_29725);
nand UO_1010 (O_1010,N_29704,N_29991);
and UO_1011 (O_1011,N_29707,N_29821);
xnor UO_1012 (O_1012,N_29764,N_29747);
or UO_1013 (O_1013,N_29792,N_29741);
and UO_1014 (O_1014,N_29802,N_29759);
or UO_1015 (O_1015,N_29975,N_29920);
xnor UO_1016 (O_1016,N_29888,N_29811);
and UO_1017 (O_1017,N_29902,N_29748);
and UO_1018 (O_1018,N_29870,N_29826);
and UO_1019 (O_1019,N_29924,N_29875);
xnor UO_1020 (O_1020,N_29907,N_29932);
xnor UO_1021 (O_1021,N_29810,N_29830);
xor UO_1022 (O_1022,N_29846,N_29996);
nor UO_1023 (O_1023,N_29999,N_29907);
or UO_1024 (O_1024,N_29875,N_29797);
nand UO_1025 (O_1025,N_29896,N_29894);
xnor UO_1026 (O_1026,N_29923,N_29929);
nor UO_1027 (O_1027,N_29751,N_29934);
xor UO_1028 (O_1028,N_29747,N_29770);
nor UO_1029 (O_1029,N_29895,N_29867);
and UO_1030 (O_1030,N_29721,N_29707);
nor UO_1031 (O_1031,N_29730,N_29715);
or UO_1032 (O_1032,N_29925,N_29719);
xnor UO_1033 (O_1033,N_29948,N_29899);
xor UO_1034 (O_1034,N_29908,N_29772);
nor UO_1035 (O_1035,N_29769,N_29882);
and UO_1036 (O_1036,N_29889,N_29823);
and UO_1037 (O_1037,N_29907,N_29849);
or UO_1038 (O_1038,N_29933,N_29994);
nand UO_1039 (O_1039,N_29947,N_29881);
xor UO_1040 (O_1040,N_29943,N_29734);
and UO_1041 (O_1041,N_29898,N_29818);
and UO_1042 (O_1042,N_29791,N_29784);
nor UO_1043 (O_1043,N_29822,N_29711);
or UO_1044 (O_1044,N_29991,N_29943);
and UO_1045 (O_1045,N_29930,N_29754);
and UO_1046 (O_1046,N_29815,N_29722);
or UO_1047 (O_1047,N_29905,N_29860);
xor UO_1048 (O_1048,N_29999,N_29968);
nor UO_1049 (O_1049,N_29970,N_29757);
or UO_1050 (O_1050,N_29718,N_29840);
or UO_1051 (O_1051,N_29923,N_29774);
and UO_1052 (O_1052,N_29872,N_29818);
or UO_1053 (O_1053,N_29910,N_29925);
xnor UO_1054 (O_1054,N_29770,N_29784);
nor UO_1055 (O_1055,N_29714,N_29813);
nor UO_1056 (O_1056,N_29778,N_29816);
or UO_1057 (O_1057,N_29733,N_29853);
xnor UO_1058 (O_1058,N_29891,N_29919);
or UO_1059 (O_1059,N_29755,N_29847);
or UO_1060 (O_1060,N_29761,N_29782);
nand UO_1061 (O_1061,N_29829,N_29960);
or UO_1062 (O_1062,N_29840,N_29882);
nand UO_1063 (O_1063,N_29925,N_29780);
nand UO_1064 (O_1064,N_29885,N_29927);
nand UO_1065 (O_1065,N_29881,N_29822);
xnor UO_1066 (O_1066,N_29722,N_29756);
nor UO_1067 (O_1067,N_29706,N_29925);
nand UO_1068 (O_1068,N_29900,N_29963);
and UO_1069 (O_1069,N_29838,N_29935);
and UO_1070 (O_1070,N_29741,N_29818);
nand UO_1071 (O_1071,N_29822,N_29888);
and UO_1072 (O_1072,N_29889,N_29876);
nand UO_1073 (O_1073,N_29926,N_29907);
nand UO_1074 (O_1074,N_29874,N_29899);
nor UO_1075 (O_1075,N_29940,N_29980);
nand UO_1076 (O_1076,N_29720,N_29777);
and UO_1077 (O_1077,N_29884,N_29984);
nand UO_1078 (O_1078,N_29811,N_29884);
nor UO_1079 (O_1079,N_29887,N_29938);
nand UO_1080 (O_1080,N_29702,N_29811);
xor UO_1081 (O_1081,N_29926,N_29711);
xnor UO_1082 (O_1082,N_29886,N_29995);
and UO_1083 (O_1083,N_29897,N_29921);
nand UO_1084 (O_1084,N_29799,N_29786);
nand UO_1085 (O_1085,N_29769,N_29756);
nand UO_1086 (O_1086,N_29800,N_29765);
nand UO_1087 (O_1087,N_29725,N_29875);
and UO_1088 (O_1088,N_29967,N_29939);
nand UO_1089 (O_1089,N_29960,N_29901);
or UO_1090 (O_1090,N_29826,N_29889);
nor UO_1091 (O_1091,N_29816,N_29806);
xor UO_1092 (O_1092,N_29892,N_29720);
xnor UO_1093 (O_1093,N_29992,N_29859);
xnor UO_1094 (O_1094,N_29771,N_29759);
and UO_1095 (O_1095,N_29825,N_29797);
and UO_1096 (O_1096,N_29709,N_29828);
and UO_1097 (O_1097,N_29860,N_29728);
and UO_1098 (O_1098,N_29704,N_29803);
or UO_1099 (O_1099,N_29866,N_29917);
nand UO_1100 (O_1100,N_29745,N_29825);
xor UO_1101 (O_1101,N_29880,N_29805);
nand UO_1102 (O_1102,N_29955,N_29706);
or UO_1103 (O_1103,N_29998,N_29780);
xnor UO_1104 (O_1104,N_29889,N_29731);
nor UO_1105 (O_1105,N_29810,N_29785);
or UO_1106 (O_1106,N_29712,N_29743);
nand UO_1107 (O_1107,N_29958,N_29761);
or UO_1108 (O_1108,N_29716,N_29731);
or UO_1109 (O_1109,N_29855,N_29929);
nand UO_1110 (O_1110,N_29805,N_29711);
xor UO_1111 (O_1111,N_29914,N_29820);
nand UO_1112 (O_1112,N_29937,N_29706);
xnor UO_1113 (O_1113,N_29745,N_29817);
nor UO_1114 (O_1114,N_29970,N_29834);
nand UO_1115 (O_1115,N_29960,N_29976);
and UO_1116 (O_1116,N_29757,N_29906);
or UO_1117 (O_1117,N_29768,N_29757);
nor UO_1118 (O_1118,N_29971,N_29704);
or UO_1119 (O_1119,N_29862,N_29794);
nor UO_1120 (O_1120,N_29842,N_29998);
xnor UO_1121 (O_1121,N_29775,N_29817);
nand UO_1122 (O_1122,N_29960,N_29923);
and UO_1123 (O_1123,N_29866,N_29881);
nor UO_1124 (O_1124,N_29934,N_29913);
or UO_1125 (O_1125,N_29956,N_29894);
xnor UO_1126 (O_1126,N_29820,N_29824);
or UO_1127 (O_1127,N_29895,N_29796);
and UO_1128 (O_1128,N_29855,N_29845);
nor UO_1129 (O_1129,N_29975,N_29879);
nand UO_1130 (O_1130,N_29854,N_29828);
and UO_1131 (O_1131,N_29902,N_29897);
nor UO_1132 (O_1132,N_29868,N_29775);
xor UO_1133 (O_1133,N_29960,N_29827);
nand UO_1134 (O_1134,N_29919,N_29956);
nor UO_1135 (O_1135,N_29712,N_29809);
nand UO_1136 (O_1136,N_29961,N_29710);
and UO_1137 (O_1137,N_29928,N_29854);
and UO_1138 (O_1138,N_29921,N_29760);
nand UO_1139 (O_1139,N_29947,N_29926);
nor UO_1140 (O_1140,N_29936,N_29949);
xnor UO_1141 (O_1141,N_29781,N_29887);
or UO_1142 (O_1142,N_29747,N_29755);
nand UO_1143 (O_1143,N_29708,N_29918);
nor UO_1144 (O_1144,N_29777,N_29968);
and UO_1145 (O_1145,N_29926,N_29822);
and UO_1146 (O_1146,N_29719,N_29857);
nor UO_1147 (O_1147,N_29937,N_29998);
or UO_1148 (O_1148,N_29831,N_29753);
xor UO_1149 (O_1149,N_29878,N_29762);
nor UO_1150 (O_1150,N_29939,N_29770);
nand UO_1151 (O_1151,N_29751,N_29828);
and UO_1152 (O_1152,N_29847,N_29722);
or UO_1153 (O_1153,N_29799,N_29836);
nor UO_1154 (O_1154,N_29993,N_29881);
or UO_1155 (O_1155,N_29993,N_29923);
nand UO_1156 (O_1156,N_29863,N_29767);
or UO_1157 (O_1157,N_29871,N_29736);
and UO_1158 (O_1158,N_29807,N_29736);
nor UO_1159 (O_1159,N_29733,N_29738);
xnor UO_1160 (O_1160,N_29742,N_29897);
nor UO_1161 (O_1161,N_29748,N_29796);
or UO_1162 (O_1162,N_29968,N_29939);
nand UO_1163 (O_1163,N_29948,N_29887);
xor UO_1164 (O_1164,N_29857,N_29840);
xnor UO_1165 (O_1165,N_29778,N_29830);
or UO_1166 (O_1166,N_29900,N_29736);
or UO_1167 (O_1167,N_29984,N_29906);
nand UO_1168 (O_1168,N_29752,N_29848);
nor UO_1169 (O_1169,N_29981,N_29773);
and UO_1170 (O_1170,N_29773,N_29952);
and UO_1171 (O_1171,N_29938,N_29945);
nor UO_1172 (O_1172,N_29883,N_29725);
or UO_1173 (O_1173,N_29928,N_29734);
xnor UO_1174 (O_1174,N_29775,N_29846);
or UO_1175 (O_1175,N_29969,N_29755);
nand UO_1176 (O_1176,N_29987,N_29923);
xnor UO_1177 (O_1177,N_29955,N_29937);
nor UO_1178 (O_1178,N_29910,N_29727);
nor UO_1179 (O_1179,N_29996,N_29835);
xnor UO_1180 (O_1180,N_29862,N_29735);
and UO_1181 (O_1181,N_29989,N_29805);
nand UO_1182 (O_1182,N_29957,N_29800);
or UO_1183 (O_1183,N_29832,N_29949);
or UO_1184 (O_1184,N_29734,N_29938);
nand UO_1185 (O_1185,N_29784,N_29701);
xor UO_1186 (O_1186,N_29808,N_29751);
nand UO_1187 (O_1187,N_29777,N_29793);
xor UO_1188 (O_1188,N_29946,N_29832);
and UO_1189 (O_1189,N_29969,N_29877);
and UO_1190 (O_1190,N_29820,N_29746);
nand UO_1191 (O_1191,N_29873,N_29887);
nor UO_1192 (O_1192,N_29970,N_29847);
and UO_1193 (O_1193,N_29825,N_29869);
or UO_1194 (O_1194,N_29808,N_29996);
and UO_1195 (O_1195,N_29700,N_29887);
xor UO_1196 (O_1196,N_29948,N_29710);
xnor UO_1197 (O_1197,N_29788,N_29832);
nand UO_1198 (O_1198,N_29977,N_29856);
and UO_1199 (O_1199,N_29760,N_29908);
nor UO_1200 (O_1200,N_29703,N_29842);
nand UO_1201 (O_1201,N_29908,N_29841);
xnor UO_1202 (O_1202,N_29861,N_29821);
and UO_1203 (O_1203,N_29903,N_29972);
nand UO_1204 (O_1204,N_29921,N_29915);
and UO_1205 (O_1205,N_29737,N_29727);
or UO_1206 (O_1206,N_29794,N_29722);
nand UO_1207 (O_1207,N_29913,N_29864);
or UO_1208 (O_1208,N_29798,N_29865);
nand UO_1209 (O_1209,N_29866,N_29779);
nand UO_1210 (O_1210,N_29700,N_29858);
nor UO_1211 (O_1211,N_29882,N_29953);
nand UO_1212 (O_1212,N_29903,N_29800);
nor UO_1213 (O_1213,N_29810,N_29835);
nor UO_1214 (O_1214,N_29951,N_29793);
xnor UO_1215 (O_1215,N_29713,N_29915);
nor UO_1216 (O_1216,N_29918,N_29843);
or UO_1217 (O_1217,N_29766,N_29715);
nor UO_1218 (O_1218,N_29827,N_29731);
and UO_1219 (O_1219,N_29834,N_29847);
or UO_1220 (O_1220,N_29937,N_29877);
nand UO_1221 (O_1221,N_29853,N_29752);
xor UO_1222 (O_1222,N_29792,N_29927);
xor UO_1223 (O_1223,N_29938,N_29914);
or UO_1224 (O_1224,N_29818,N_29711);
nor UO_1225 (O_1225,N_29876,N_29799);
and UO_1226 (O_1226,N_29827,N_29924);
xor UO_1227 (O_1227,N_29819,N_29931);
xnor UO_1228 (O_1228,N_29833,N_29721);
nand UO_1229 (O_1229,N_29927,N_29754);
nand UO_1230 (O_1230,N_29949,N_29814);
nand UO_1231 (O_1231,N_29859,N_29896);
xor UO_1232 (O_1232,N_29705,N_29811);
nor UO_1233 (O_1233,N_29996,N_29857);
nand UO_1234 (O_1234,N_29812,N_29776);
or UO_1235 (O_1235,N_29900,N_29780);
or UO_1236 (O_1236,N_29757,N_29822);
xor UO_1237 (O_1237,N_29744,N_29963);
and UO_1238 (O_1238,N_29809,N_29704);
nand UO_1239 (O_1239,N_29776,N_29741);
nor UO_1240 (O_1240,N_29869,N_29796);
xnor UO_1241 (O_1241,N_29881,N_29912);
or UO_1242 (O_1242,N_29773,N_29707);
nor UO_1243 (O_1243,N_29734,N_29949);
nand UO_1244 (O_1244,N_29995,N_29930);
and UO_1245 (O_1245,N_29962,N_29709);
xnor UO_1246 (O_1246,N_29747,N_29950);
nand UO_1247 (O_1247,N_29832,N_29708);
or UO_1248 (O_1248,N_29754,N_29940);
nand UO_1249 (O_1249,N_29910,N_29956);
xor UO_1250 (O_1250,N_29867,N_29796);
and UO_1251 (O_1251,N_29873,N_29964);
xor UO_1252 (O_1252,N_29921,N_29830);
xor UO_1253 (O_1253,N_29802,N_29757);
or UO_1254 (O_1254,N_29797,N_29716);
nor UO_1255 (O_1255,N_29812,N_29892);
or UO_1256 (O_1256,N_29978,N_29862);
or UO_1257 (O_1257,N_29780,N_29849);
xnor UO_1258 (O_1258,N_29985,N_29904);
xnor UO_1259 (O_1259,N_29944,N_29787);
xnor UO_1260 (O_1260,N_29950,N_29739);
and UO_1261 (O_1261,N_29764,N_29857);
or UO_1262 (O_1262,N_29890,N_29945);
or UO_1263 (O_1263,N_29956,N_29809);
or UO_1264 (O_1264,N_29986,N_29747);
and UO_1265 (O_1265,N_29842,N_29737);
nand UO_1266 (O_1266,N_29789,N_29920);
nor UO_1267 (O_1267,N_29869,N_29821);
nor UO_1268 (O_1268,N_29769,N_29783);
xor UO_1269 (O_1269,N_29968,N_29794);
nand UO_1270 (O_1270,N_29861,N_29942);
nand UO_1271 (O_1271,N_29883,N_29803);
xor UO_1272 (O_1272,N_29757,N_29977);
and UO_1273 (O_1273,N_29945,N_29883);
and UO_1274 (O_1274,N_29835,N_29970);
nor UO_1275 (O_1275,N_29870,N_29799);
xor UO_1276 (O_1276,N_29732,N_29962);
and UO_1277 (O_1277,N_29810,N_29777);
or UO_1278 (O_1278,N_29953,N_29724);
or UO_1279 (O_1279,N_29823,N_29904);
xor UO_1280 (O_1280,N_29978,N_29944);
or UO_1281 (O_1281,N_29895,N_29915);
and UO_1282 (O_1282,N_29721,N_29844);
or UO_1283 (O_1283,N_29930,N_29804);
nor UO_1284 (O_1284,N_29978,N_29959);
nor UO_1285 (O_1285,N_29919,N_29990);
nand UO_1286 (O_1286,N_29720,N_29805);
nand UO_1287 (O_1287,N_29827,N_29710);
or UO_1288 (O_1288,N_29755,N_29721);
and UO_1289 (O_1289,N_29732,N_29745);
and UO_1290 (O_1290,N_29841,N_29737);
and UO_1291 (O_1291,N_29799,N_29879);
nand UO_1292 (O_1292,N_29785,N_29911);
nor UO_1293 (O_1293,N_29984,N_29988);
nor UO_1294 (O_1294,N_29933,N_29748);
nand UO_1295 (O_1295,N_29720,N_29935);
nand UO_1296 (O_1296,N_29798,N_29816);
nor UO_1297 (O_1297,N_29750,N_29998);
nor UO_1298 (O_1298,N_29841,N_29845);
or UO_1299 (O_1299,N_29992,N_29886);
nand UO_1300 (O_1300,N_29828,N_29964);
nor UO_1301 (O_1301,N_29743,N_29756);
and UO_1302 (O_1302,N_29982,N_29709);
nand UO_1303 (O_1303,N_29712,N_29815);
nand UO_1304 (O_1304,N_29938,N_29939);
and UO_1305 (O_1305,N_29877,N_29727);
or UO_1306 (O_1306,N_29733,N_29742);
nor UO_1307 (O_1307,N_29727,N_29818);
xor UO_1308 (O_1308,N_29860,N_29761);
nand UO_1309 (O_1309,N_29767,N_29927);
xor UO_1310 (O_1310,N_29732,N_29838);
or UO_1311 (O_1311,N_29712,N_29925);
xnor UO_1312 (O_1312,N_29989,N_29702);
nand UO_1313 (O_1313,N_29742,N_29991);
or UO_1314 (O_1314,N_29962,N_29984);
xor UO_1315 (O_1315,N_29873,N_29973);
nor UO_1316 (O_1316,N_29808,N_29973);
nand UO_1317 (O_1317,N_29960,N_29911);
and UO_1318 (O_1318,N_29866,N_29943);
and UO_1319 (O_1319,N_29876,N_29929);
nor UO_1320 (O_1320,N_29874,N_29845);
nor UO_1321 (O_1321,N_29730,N_29890);
nand UO_1322 (O_1322,N_29908,N_29730);
xnor UO_1323 (O_1323,N_29805,N_29999);
xnor UO_1324 (O_1324,N_29842,N_29965);
or UO_1325 (O_1325,N_29903,N_29717);
or UO_1326 (O_1326,N_29709,N_29821);
or UO_1327 (O_1327,N_29893,N_29832);
xnor UO_1328 (O_1328,N_29804,N_29862);
or UO_1329 (O_1329,N_29921,N_29972);
xor UO_1330 (O_1330,N_29958,N_29712);
nor UO_1331 (O_1331,N_29957,N_29917);
nand UO_1332 (O_1332,N_29989,N_29893);
nor UO_1333 (O_1333,N_29816,N_29745);
and UO_1334 (O_1334,N_29950,N_29725);
and UO_1335 (O_1335,N_29834,N_29832);
and UO_1336 (O_1336,N_29860,N_29799);
nor UO_1337 (O_1337,N_29794,N_29978);
nand UO_1338 (O_1338,N_29967,N_29931);
nand UO_1339 (O_1339,N_29857,N_29981);
nand UO_1340 (O_1340,N_29843,N_29732);
xnor UO_1341 (O_1341,N_29734,N_29700);
or UO_1342 (O_1342,N_29855,N_29933);
and UO_1343 (O_1343,N_29875,N_29816);
nand UO_1344 (O_1344,N_29739,N_29941);
xnor UO_1345 (O_1345,N_29768,N_29983);
or UO_1346 (O_1346,N_29757,N_29972);
or UO_1347 (O_1347,N_29759,N_29934);
and UO_1348 (O_1348,N_29889,N_29875);
xor UO_1349 (O_1349,N_29739,N_29960);
nand UO_1350 (O_1350,N_29926,N_29969);
nand UO_1351 (O_1351,N_29924,N_29819);
nor UO_1352 (O_1352,N_29736,N_29714);
nand UO_1353 (O_1353,N_29752,N_29972);
or UO_1354 (O_1354,N_29731,N_29843);
or UO_1355 (O_1355,N_29723,N_29809);
nand UO_1356 (O_1356,N_29836,N_29793);
or UO_1357 (O_1357,N_29913,N_29853);
xnor UO_1358 (O_1358,N_29832,N_29816);
nor UO_1359 (O_1359,N_29897,N_29841);
nand UO_1360 (O_1360,N_29792,N_29864);
or UO_1361 (O_1361,N_29930,N_29990);
nor UO_1362 (O_1362,N_29816,N_29917);
or UO_1363 (O_1363,N_29950,N_29799);
nor UO_1364 (O_1364,N_29974,N_29764);
nand UO_1365 (O_1365,N_29846,N_29938);
xnor UO_1366 (O_1366,N_29775,N_29737);
nor UO_1367 (O_1367,N_29994,N_29717);
or UO_1368 (O_1368,N_29727,N_29826);
xor UO_1369 (O_1369,N_29965,N_29752);
xor UO_1370 (O_1370,N_29930,N_29947);
nand UO_1371 (O_1371,N_29859,N_29773);
xnor UO_1372 (O_1372,N_29752,N_29937);
and UO_1373 (O_1373,N_29861,N_29740);
nor UO_1374 (O_1374,N_29707,N_29878);
nand UO_1375 (O_1375,N_29960,N_29991);
and UO_1376 (O_1376,N_29738,N_29792);
nand UO_1377 (O_1377,N_29761,N_29840);
and UO_1378 (O_1378,N_29806,N_29926);
or UO_1379 (O_1379,N_29872,N_29784);
nor UO_1380 (O_1380,N_29752,N_29923);
nand UO_1381 (O_1381,N_29896,N_29732);
xor UO_1382 (O_1382,N_29789,N_29827);
and UO_1383 (O_1383,N_29776,N_29964);
nand UO_1384 (O_1384,N_29853,N_29770);
nor UO_1385 (O_1385,N_29992,N_29954);
nor UO_1386 (O_1386,N_29999,N_29817);
and UO_1387 (O_1387,N_29811,N_29893);
or UO_1388 (O_1388,N_29786,N_29988);
nand UO_1389 (O_1389,N_29931,N_29977);
nor UO_1390 (O_1390,N_29797,N_29827);
or UO_1391 (O_1391,N_29886,N_29984);
or UO_1392 (O_1392,N_29801,N_29748);
and UO_1393 (O_1393,N_29827,N_29963);
and UO_1394 (O_1394,N_29914,N_29927);
nor UO_1395 (O_1395,N_29751,N_29875);
nand UO_1396 (O_1396,N_29784,N_29793);
nand UO_1397 (O_1397,N_29922,N_29860);
and UO_1398 (O_1398,N_29795,N_29920);
nor UO_1399 (O_1399,N_29904,N_29755);
xnor UO_1400 (O_1400,N_29885,N_29920);
xnor UO_1401 (O_1401,N_29761,N_29833);
nor UO_1402 (O_1402,N_29768,N_29759);
or UO_1403 (O_1403,N_29895,N_29839);
nor UO_1404 (O_1404,N_29788,N_29705);
and UO_1405 (O_1405,N_29821,N_29745);
nor UO_1406 (O_1406,N_29777,N_29898);
and UO_1407 (O_1407,N_29980,N_29962);
or UO_1408 (O_1408,N_29822,N_29724);
or UO_1409 (O_1409,N_29842,N_29887);
nand UO_1410 (O_1410,N_29784,N_29782);
and UO_1411 (O_1411,N_29981,N_29725);
and UO_1412 (O_1412,N_29830,N_29905);
xor UO_1413 (O_1413,N_29919,N_29976);
nand UO_1414 (O_1414,N_29919,N_29973);
or UO_1415 (O_1415,N_29761,N_29746);
xor UO_1416 (O_1416,N_29924,N_29988);
xor UO_1417 (O_1417,N_29759,N_29988);
xnor UO_1418 (O_1418,N_29984,N_29931);
or UO_1419 (O_1419,N_29846,N_29990);
and UO_1420 (O_1420,N_29965,N_29936);
or UO_1421 (O_1421,N_29982,N_29748);
or UO_1422 (O_1422,N_29972,N_29802);
xnor UO_1423 (O_1423,N_29877,N_29806);
nor UO_1424 (O_1424,N_29864,N_29865);
xnor UO_1425 (O_1425,N_29834,N_29926);
and UO_1426 (O_1426,N_29747,N_29706);
nand UO_1427 (O_1427,N_29877,N_29846);
nand UO_1428 (O_1428,N_29841,N_29960);
and UO_1429 (O_1429,N_29772,N_29745);
nor UO_1430 (O_1430,N_29827,N_29870);
nand UO_1431 (O_1431,N_29952,N_29995);
nand UO_1432 (O_1432,N_29708,N_29946);
nand UO_1433 (O_1433,N_29990,N_29795);
nand UO_1434 (O_1434,N_29872,N_29805);
nand UO_1435 (O_1435,N_29931,N_29836);
xor UO_1436 (O_1436,N_29731,N_29733);
xnor UO_1437 (O_1437,N_29908,N_29962);
or UO_1438 (O_1438,N_29900,N_29786);
and UO_1439 (O_1439,N_29967,N_29725);
or UO_1440 (O_1440,N_29927,N_29886);
nor UO_1441 (O_1441,N_29749,N_29981);
and UO_1442 (O_1442,N_29878,N_29918);
xor UO_1443 (O_1443,N_29835,N_29907);
nor UO_1444 (O_1444,N_29999,N_29867);
nand UO_1445 (O_1445,N_29746,N_29747);
xor UO_1446 (O_1446,N_29903,N_29992);
and UO_1447 (O_1447,N_29707,N_29916);
or UO_1448 (O_1448,N_29950,N_29741);
nand UO_1449 (O_1449,N_29982,N_29784);
and UO_1450 (O_1450,N_29923,N_29842);
nand UO_1451 (O_1451,N_29753,N_29934);
nor UO_1452 (O_1452,N_29924,N_29821);
nor UO_1453 (O_1453,N_29712,N_29779);
or UO_1454 (O_1454,N_29976,N_29959);
or UO_1455 (O_1455,N_29732,N_29948);
xor UO_1456 (O_1456,N_29989,N_29743);
nand UO_1457 (O_1457,N_29806,N_29975);
nand UO_1458 (O_1458,N_29805,N_29799);
nor UO_1459 (O_1459,N_29742,N_29824);
or UO_1460 (O_1460,N_29950,N_29881);
or UO_1461 (O_1461,N_29702,N_29898);
nor UO_1462 (O_1462,N_29708,N_29926);
nand UO_1463 (O_1463,N_29992,N_29932);
nor UO_1464 (O_1464,N_29858,N_29923);
or UO_1465 (O_1465,N_29723,N_29850);
or UO_1466 (O_1466,N_29951,N_29962);
nor UO_1467 (O_1467,N_29943,N_29879);
nand UO_1468 (O_1468,N_29863,N_29950);
xnor UO_1469 (O_1469,N_29703,N_29722);
nand UO_1470 (O_1470,N_29727,N_29933);
nand UO_1471 (O_1471,N_29707,N_29962);
and UO_1472 (O_1472,N_29782,N_29933);
xor UO_1473 (O_1473,N_29861,N_29906);
or UO_1474 (O_1474,N_29885,N_29899);
nor UO_1475 (O_1475,N_29771,N_29967);
nor UO_1476 (O_1476,N_29827,N_29925);
or UO_1477 (O_1477,N_29956,N_29942);
nor UO_1478 (O_1478,N_29887,N_29706);
nand UO_1479 (O_1479,N_29923,N_29922);
nor UO_1480 (O_1480,N_29737,N_29941);
nor UO_1481 (O_1481,N_29702,N_29987);
xor UO_1482 (O_1482,N_29795,N_29992);
xor UO_1483 (O_1483,N_29870,N_29889);
and UO_1484 (O_1484,N_29894,N_29753);
nor UO_1485 (O_1485,N_29715,N_29894);
nor UO_1486 (O_1486,N_29820,N_29780);
and UO_1487 (O_1487,N_29935,N_29979);
xor UO_1488 (O_1488,N_29863,N_29823);
or UO_1489 (O_1489,N_29727,N_29710);
nor UO_1490 (O_1490,N_29715,N_29810);
xnor UO_1491 (O_1491,N_29800,N_29721);
or UO_1492 (O_1492,N_29880,N_29984);
nor UO_1493 (O_1493,N_29769,N_29786);
xor UO_1494 (O_1494,N_29856,N_29822);
or UO_1495 (O_1495,N_29894,N_29869);
nor UO_1496 (O_1496,N_29884,N_29958);
or UO_1497 (O_1497,N_29973,N_29797);
xnor UO_1498 (O_1498,N_29989,N_29896);
nand UO_1499 (O_1499,N_29705,N_29863);
and UO_1500 (O_1500,N_29910,N_29924);
nor UO_1501 (O_1501,N_29759,N_29797);
xor UO_1502 (O_1502,N_29958,N_29987);
and UO_1503 (O_1503,N_29973,N_29784);
xnor UO_1504 (O_1504,N_29789,N_29952);
nor UO_1505 (O_1505,N_29919,N_29963);
nor UO_1506 (O_1506,N_29788,N_29869);
or UO_1507 (O_1507,N_29900,N_29745);
or UO_1508 (O_1508,N_29768,N_29725);
nor UO_1509 (O_1509,N_29863,N_29795);
xor UO_1510 (O_1510,N_29961,N_29824);
xnor UO_1511 (O_1511,N_29741,N_29880);
nand UO_1512 (O_1512,N_29962,N_29808);
and UO_1513 (O_1513,N_29806,N_29900);
nand UO_1514 (O_1514,N_29972,N_29727);
or UO_1515 (O_1515,N_29839,N_29760);
and UO_1516 (O_1516,N_29979,N_29999);
nand UO_1517 (O_1517,N_29826,N_29716);
nand UO_1518 (O_1518,N_29731,N_29708);
nor UO_1519 (O_1519,N_29905,N_29718);
nand UO_1520 (O_1520,N_29734,N_29813);
and UO_1521 (O_1521,N_29744,N_29904);
nand UO_1522 (O_1522,N_29932,N_29747);
xor UO_1523 (O_1523,N_29746,N_29953);
nor UO_1524 (O_1524,N_29893,N_29710);
or UO_1525 (O_1525,N_29999,N_29719);
nand UO_1526 (O_1526,N_29796,N_29733);
nor UO_1527 (O_1527,N_29707,N_29744);
nand UO_1528 (O_1528,N_29859,N_29925);
or UO_1529 (O_1529,N_29723,N_29811);
or UO_1530 (O_1530,N_29847,N_29853);
xnor UO_1531 (O_1531,N_29731,N_29961);
or UO_1532 (O_1532,N_29749,N_29908);
and UO_1533 (O_1533,N_29726,N_29708);
or UO_1534 (O_1534,N_29786,N_29717);
nand UO_1535 (O_1535,N_29859,N_29849);
nand UO_1536 (O_1536,N_29798,N_29936);
nor UO_1537 (O_1537,N_29706,N_29737);
or UO_1538 (O_1538,N_29984,N_29881);
xnor UO_1539 (O_1539,N_29956,N_29793);
and UO_1540 (O_1540,N_29752,N_29732);
xor UO_1541 (O_1541,N_29969,N_29707);
nand UO_1542 (O_1542,N_29789,N_29974);
or UO_1543 (O_1543,N_29954,N_29991);
nand UO_1544 (O_1544,N_29962,N_29933);
nor UO_1545 (O_1545,N_29938,N_29807);
nand UO_1546 (O_1546,N_29958,N_29726);
and UO_1547 (O_1547,N_29936,N_29857);
nor UO_1548 (O_1548,N_29854,N_29733);
or UO_1549 (O_1549,N_29758,N_29700);
xor UO_1550 (O_1550,N_29703,N_29925);
and UO_1551 (O_1551,N_29756,N_29733);
nand UO_1552 (O_1552,N_29898,N_29904);
or UO_1553 (O_1553,N_29840,N_29764);
and UO_1554 (O_1554,N_29984,N_29973);
and UO_1555 (O_1555,N_29704,N_29737);
or UO_1556 (O_1556,N_29725,N_29859);
nor UO_1557 (O_1557,N_29752,N_29869);
nand UO_1558 (O_1558,N_29725,N_29738);
and UO_1559 (O_1559,N_29851,N_29786);
nor UO_1560 (O_1560,N_29706,N_29906);
nand UO_1561 (O_1561,N_29838,N_29710);
or UO_1562 (O_1562,N_29746,N_29834);
or UO_1563 (O_1563,N_29792,N_29793);
nor UO_1564 (O_1564,N_29986,N_29930);
xnor UO_1565 (O_1565,N_29908,N_29818);
nor UO_1566 (O_1566,N_29791,N_29745);
nand UO_1567 (O_1567,N_29745,N_29885);
and UO_1568 (O_1568,N_29954,N_29892);
nor UO_1569 (O_1569,N_29797,N_29725);
nand UO_1570 (O_1570,N_29935,N_29716);
or UO_1571 (O_1571,N_29893,N_29929);
and UO_1572 (O_1572,N_29735,N_29885);
nor UO_1573 (O_1573,N_29838,N_29963);
or UO_1574 (O_1574,N_29911,N_29978);
nor UO_1575 (O_1575,N_29714,N_29710);
or UO_1576 (O_1576,N_29845,N_29870);
or UO_1577 (O_1577,N_29984,N_29815);
or UO_1578 (O_1578,N_29775,N_29878);
nand UO_1579 (O_1579,N_29951,N_29782);
xor UO_1580 (O_1580,N_29734,N_29937);
xnor UO_1581 (O_1581,N_29703,N_29872);
xor UO_1582 (O_1582,N_29990,N_29905);
xor UO_1583 (O_1583,N_29805,N_29859);
nand UO_1584 (O_1584,N_29776,N_29910);
or UO_1585 (O_1585,N_29741,N_29835);
nand UO_1586 (O_1586,N_29762,N_29987);
and UO_1587 (O_1587,N_29775,N_29800);
xor UO_1588 (O_1588,N_29820,N_29969);
nor UO_1589 (O_1589,N_29956,N_29725);
and UO_1590 (O_1590,N_29935,N_29718);
nor UO_1591 (O_1591,N_29740,N_29874);
or UO_1592 (O_1592,N_29783,N_29896);
nand UO_1593 (O_1593,N_29931,N_29923);
and UO_1594 (O_1594,N_29754,N_29728);
nand UO_1595 (O_1595,N_29703,N_29780);
or UO_1596 (O_1596,N_29992,N_29865);
nor UO_1597 (O_1597,N_29769,N_29795);
and UO_1598 (O_1598,N_29845,N_29946);
nand UO_1599 (O_1599,N_29941,N_29945);
or UO_1600 (O_1600,N_29975,N_29835);
nor UO_1601 (O_1601,N_29706,N_29981);
or UO_1602 (O_1602,N_29782,N_29889);
or UO_1603 (O_1603,N_29768,N_29952);
and UO_1604 (O_1604,N_29983,N_29992);
and UO_1605 (O_1605,N_29731,N_29907);
nand UO_1606 (O_1606,N_29785,N_29749);
and UO_1607 (O_1607,N_29959,N_29889);
nor UO_1608 (O_1608,N_29997,N_29936);
xor UO_1609 (O_1609,N_29828,N_29804);
and UO_1610 (O_1610,N_29872,N_29946);
nand UO_1611 (O_1611,N_29988,N_29900);
xor UO_1612 (O_1612,N_29787,N_29900);
and UO_1613 (O_1613,N_29760,N_29951);
nand UO_1614 (O_1614,N_29808,N_29789);
nor UO_1615 (O_1615,N_29758,N_29935);
nor UO_1616 (O_1616,N_29779,N_29842);
and UO_1617 (O_1617,N_29741,N_29964);
or UO_1618 (O_1618,N_29758,N_29823);
nand UO_1619 (O_1619,N_29852,N_29929);
nand UO_1620 (O_1620,N_29865,N_29955);
and UO_1621 (O_1621,N_29920,N_29755);
or UO_1622 (O_1622,N_29951,N_29799);
or UO_1623 (O_1623,N_29912,N_29730);
nand UO_1624 (O_1624,N_29865,N_29902);
and UO_1625 (O_1625,N_29869,N_29841);
nand UO_1626 (O_1626,N_29924,N_29939);
nor UO_1627 (O_1627,N_29907,N_29883);
and UO_1628 (O_1628,N_29860,N_29736);
or UO_1629 (O_1629,N_29754,N_29845);
nand UO_1630 (O_1630,N_29963,N_29732);
nand UO_1631 (O_1631,N_29742,N_29908);
nand UO_1632 (O_1632,N_29777,N_29998);
and UO_1633 (O_1633,N_29748,N_29900);
nor UO_1634 (O_1634,N_29959,N_29798);
or UO_1635 (O_1635,N_29962,N_29928);
xnor UO_1636 (O_1636,N_29898,N_29728);
xnor UO_1637 (O_1637,N_29903,N_29960);
nand UO_1638 (O_1638,N_29846,N_29921);
and UO_1639 (O_1639,N_29749,N_29741);
or UO_1640 (O_1640,N_29872,N_29965);
xor UO_1641 (O_1641,N_29840,N_29704);
nor UO_1642 (O_1642,N_29921,N_29724);
and UO_1643 (O_1643,N_29795,N_29744);
nand UO_1644 (O_1644,N_29893,N_29761);
xor UO_1645 (O_1645,N_29808,N_29785);
and UO_1646 (O_1646,N_29754,N_29898);
nand UO_1647 (O_1647,N_29734,N_29837);
nand UO_1648 (O_1648,N_29834,N_29952);
nor UO_1649 (O_1649,N_29875,N_29850);
nand UO_1650 (O_1650,N_29752,N_29718);
xor UO_1651 (O_1651,N_29813,N_29858);
nor UO_1652 (O_1652,N_29707,N_29975);
nand UO_1653 (O_1653,N_29722,N_29863);
nand UO_1654 (O_1654,N_29827,N_29754);
and UO_1655 (O_1655,N_29943,N_29969);
nand UO_1656 (O_1656,N_29772,N_29843);
and UO_1657 (O_1657,N_29732,N_29828);
xor UO_1658 (O_1658,N_29893,N_29712);
nor UO_1659 (O_1659,N_29802,N_29821);
nor UO_1660 (O_1660,N_29920,N_29811);
xnor UO_1661 (O_1661,N_29917,N_29713);
nor UO_1662 (O_1662,N_29743,N_29824);
nand UO_1663 (O_1663,N_29804,N_29765);
nor UO_1664 (O_1664,N_29852,N_29909);
and UO_1665 (O_1665,N_29890,N_29928);
and UO_1666 (O_1666,N_29711,N_29945);
or UO_1667 (O_1667,N_29882,N_29967);
nand UO_1668 (O_1668,N_29736,N_29837);
or UO_1669 (O_1669,N_29813,N_29916);
and UO_1670 (O_1670,N_29974,N_29898);
or UO_1671 (O_1671,N_29745,N_29818);
or UO_1672 (O_1672,N_29969,N_29768);
nor UO_1673 (O_1673,N_29868,N_29989);
or UO_1674 (O_1674,N_29867,N_29833);
xnor UO_1675 (O_1675,N_29785,N_29868);
or UO_1676 (O_1676,N_29729,N_29817);
nor UO_1677 (O_1677,N_29925,N_29985);
nand UO_1678 (O_1678,N_29722,N_29901);
xor UO_1679 (O_1679,N_29731,N_29779);
nand UO_1680 (O_1680,N_29924,N_29855);
and UO_1681 (O_1681,N_29995,N_29968);
nand UO_1682 (O_1682,N_29999,N_29803);
nand UO_1683 (O_1683,N_29703,N_29862);
nor UO_1684 (O_1684,N_29825,N_29964);
and UO_1685 (O_1685,N_29924,N_29756);
nand UO_1686 (O_1686,N_29839,N_29766);
xor UO_1687 (O_1687,N_29901,N_29966);
nand UO_1688 (O_1688,N_29992,N_29991);
or UO_1689 (O_1689,N_29875,N_29819);
nand UO_1690 (O_1690,N_29947,N_29855);
or UO_1691 (O_1691,N_29846,N_29779);
xnor UO_1692 (O_1692,N_29841,N_29978);
xnor UO_1693 (O_1693,N_29862,N_29786);
and UO_1694 (O_1694,N_29760,N_29835);
or UO_1695 (O_1695,N_29935,N_29911);
nor UO_1696 (O_1696,N_29859,N_29889);
nor UO_1697 (O_1697,N_29847,N_29867);
nand UO_1698 (O_1698,N_29708,N_29861);
nand UO_1699 (O_1699,N_29873,N_29930);
nor UO_1700 (O_1700,N_29906,N_29843);
and UO_1701 (O_1701,N_29774,N_29784);
nor UO_1702 (O_1702,N_29794,N_29987);
or UO_1703 (O_1703,N_29998,N_29935);
nor UO_1704 (O_1704,N_29711,N_29706);
and UO_1705 (O_1705,N_29971,N_29946);
nand UO_1706 (O_1706,N_29711,N_29765);
and UO_1707 (O_1707,N_29986,N_29731);
nor UO_1708 (O_1708,N_29921,N_29904);
nor UO_1709 (O_1709,N_29805,N_29838);
nor UO_1710 (O_1710,N_29812,N_29966);
or UO_1711 (O_1711,N_29882,N_29929);
xor UO_1712 (O_1712,N_29844,N_29937);
xnor UO_1713 (O_1713,N_29982,N_29844);
or UO_1714 (O_1714,N_29775,N_29874);
nor UO_1715 (O_1715,N_29758,N_29755);
or UO_1716 (O_1716,N_29834,N_29798);
nor UO_1717 (O_1717,N_29797,N_29842);
nand UO_1718 (O_1718,N_29847,N_29854);
or UO_1719 (O_1719,N_29968,N_29824);
xnor UO_1720 (O_1720,N_29956,N_29958);
nor UO_1721 (O_1721,N_29889,N_29864);
and UO_1722 (O_1722,N_29825,N_29835);
nor UO_1723 (O_1723,N_29946,N_29919);
xnor UO_1724 (O_1724,N_29914,N_29849);
or UO_1725 (O_1725,N_29838,N_29702);
nor UO_1726 (O_1726,N_29997,N_29711);
or UO_1727 (O_1727,N_29837,N_29719);
nand UO_1728 (O_1728,N_29902,N_29869);
nand UO_1729 (O_1729,N_29867,N_29807);
or UO_1730 (O_1730,N_29831,N_29864);
xnor UO_1731 (O_1731,N_29812,N_29817);
or UO_1732 (O_1732,N_29815,N_29755);
nor UO_1733 (O_1733,N_29817,N_29827);
or UO_1734 (O_1734,N_29764,N_29936);
xor UO_1735 (O_1735,N_29836,N_29777);
nor UO_1736 (O_1736,N_29908,N_29767);
nor UO_1737 (O_1737,N_29849,N_29994);
and UO_1738 (O_1738,N_29830,N_29899);
and UO_1739 (O_1739,N_29901,N_29786);
and UO_1740 (O_1740,N_29803,N_29965);
and UO_1741 (O_1741,N_29839,N_29865);
or UO_1742 (O_1742,N_29916,N_29846);
xor UO_1743 (O_1743,N_29926,N_29804);
nor UO_1744 (O_1744,N_29773,N_29885);
or UO_1745 (O_1745,N_29744,N_29893);
nand UO_1746 (O_1746,N_29708,N_29728);
or UO_1747 (O_1747,N_29987,N_29868);
xor UO_1748 (O_1748,N_29764,N_29804);
nand UO_1749 (O_1749,N_29714,N_29995);
xor UO_1750 (O_1750,N_29940,N_29880);
nor UO_1751 (O_1751,N_29771,N_29900);
and UO_1752 (O_1752,N_29723,N_29898);
xor UO_1753 (O_1753,N_29919,N_29924);
xor UO_1754 (O_1754,N_29917,N_29756);
nor UO_1755 (O_1755,N_29751,N_29945);
and UO_1756 (O_1756,N_29711,N_29960);
nor UO_1757 (O_1757,N_29718,N_29944);
nand UO_1758 (O_1758,N_29863,N_29748);
xnor UO_1759 (O_1759,N_29754,N_29946);
and UO_1760 (O_1760,N_29881,N_29934);
nand UO_1761 (O_1761,N_29998,N_29756);
and UO_1762 (O_1762,N_29735,N_29941);
and UO_1763 (O_1763,N_29915,N_29901);
or UO_1764 (O_1764,N_29829,N_29810);
or UO_1765 (O_1765,N_29987,N_29907);
and UO_1766 (O_1766,N_29754,N_29910);
nor UO_1767 (O_1767,N_29991,N_29709);
or UO_1768 (O_1768,N_29811,N_29941);
or UO_1769 (O_1769,N_29944,N_29762);
xor UO_1770 (O_1770,N_29771,N_29920);
nor UO_1771 (O_1771,N_29704,N_29827);
xnor UO_1772 (O_1772,N_29839,N_29968);
xor UO_1773 (O_1773,N_29745,N_29967);
xor UO_1774 (O_1774,N_29852,N_29814);
nand UO_1775 (O_1775,N_29968,N_29991);
xnor UO_1776 (O_1776,N_29976,N_29766);
or UO_1777 (O_1777,N_29959,N_29935);
xnor UO_1778 (O_1778,N_29931,N_29869);
and UO_1779 (O_1779,N_29997,N_29910);
nand UO_1780 (O_1780,N_29783,N_29868);
and UO_1781 (O_1781,N_29762,N_29863);
and UO_1782 (O_1782,N_29982,N_29954);
nor UO_1783 (O_1783,N_29706,N_29758);
and UO_1784 (O_1784,N_29957,N_29995);
or UO_1785 (O_1785,N_29841,N_29928);
xor UO_1786 (O_1786,N_29713,N_29838);
nor UO_1787 (O_1787,N_29920,N_29958);
nor UO_1788 (O_1788,N_29901,N_29820);
nor UO_1789 (O_1789,N_29759,N_29852);
xor UO_1790 (O_1790,N_29707,N_29944);
nand UO_1791 (O_1791,N_29854,N_29975);
nor UO_1792 (O_1792,N_29966,N_29828);
nor UO_1793 (O_1793,N_29815,N_29824);
nand UO_1794 (O_1794,N_29978,N_29868);
or UO_1795 (O_1795,N_29776,N_29888);
nor UO_1796 (O_1796,N_29795,N_29976);
xor UO_1797 (O_1797,N_29737,N_29859);
or UO_1798 (O_1798,N_29801,N_29971);
xnor UO_1799 (O_1799,N_29730,N_29936);
xor UO_1800 (O_1800,N_29928,N_29746);
or UO_1801 (O_1801,N_29999,N_29875);
xnor UO_1802 (O_1802,N_29718,N_29704);
and UO_1803 (O_1803,N_29780,N_29973);
or UO_1804 (O_1804,N_29911,N_29830);
or UO_1805 (O_1805,N_29708,N_29887);
and UO_1806 (O_1806,N_29804,N_29993);
nor UO_1807 (O_1807,N_29746,N_29858);
nand UO_1808 (O_1808,N_29994,N_29877);
and UO_1809 (O_1809,N_29865,N_29845);
or UO_1810 (O_1810,N_29746,N_29797);
nor UO_1811 (O_1811,N_29962,N_29971);
nand UO_1812 (O_1812,N_29860,N_29936);
nand UO_1813 (O_1813,N_29832,N_29780);
or UO_1814 (O_1814,N_29886,N_29761);
nor UO_1815 (O_1815,N_29851,N_29837);
nor UO_1816 (O_1816,N_29814,N_29751);
or UO_1817 (O_1817,N_29969,N_29861);
nand UO_1818 (O_1818,N_29860,N_29883);
xnor UO_1819 (O_1819,N_29797,N_29997);
and UO_1820 (O_1820,N_29928,N_29882);
or UO_1821 (O_1821,N_29881,N_29919);
nor UO_1822 (O_1822,N_29765,N_29926);
nor UO_1823 (O_1823,N_29703,N_29785);
nor UO_1824 (O_1824,N_29852,N_29822);
and UO_1825 (O_1825,N_29833,N_29830);
nand UO_1826 (O_1826,N_29846,N_29825);
nor UO_1827 (O_1827,N_29731,N_29778);
or UO_1828 (O_1828,N_29766,N_29943);
nand UO_1829 (O_1829,N_29919,N_29795);
xor UO_1830 (O_1830,N_29742,N_29881);
nor UO_1831 (O_1831,N_29744,N_29724);
and UO_1832 (O_1832,N_29801,N_29978);
or UO_1833 (O_1833,N_29971,N_29808);
and UO_1834 (O_1834,N_29808,N_29836);
xnor UO_1835 (O_1835,N_29710,N_29884);
or UO_1836 (O_1836,N_29937,N_29951);
and UO_1837 (O_1837,N_29848,N_29996);
and UO_1838 (O_1838,N_29774,N_29956);
xnor UO_1839 (O_1839,N_29786,N_29745);
xnor UO_1840 (O_1840,N_29953,N_29894);
nand UO_1841 (O_1841,N_29714,N_29815);
xnor UO_1842 (O_1842,N_29891,N_29763);
xor UO_1843 (O_1843,N_29875,N_29786);
xnor UO_1844 (O_1844,N_29966,N_29712);
nor UO_1845 (O_1845,N_29894,N_29833);
or UO_1846 (O_1846,N_29794,N_29955);
nand UO_1847 (O_1847,N_29746,N_29855);
nor UO_1848 (O_1848,N_29818,N_29999);
xnor UO_1849 (O_1849,N_29736,N_29912);
nor UO_1850 (O_1850,N_29951,N_29765);
and UO_1851 (O_1851,N_29831,N_29948);
xor UO_1852 (O_1852,N_29718,N_29788);
nor UO_1853 (O_1853,N_29787,N_29943);
nand UO_1854 (O_1854,N_29853,N_29883);
nand UO_1855 (O_1855,N_29947,N_29964);
xor UO_1856 (O_1856,N_29876,N_29871);
xor UO_1857 (O_1857,N_29972,N_29847);
xnor UO_1858 (O_1858,N_29977,N_29709);
or UO_1859 (O_1859,N_29891,N_29982);
or UO_1860 (O_1860,N_29751,N_29988);
or UO_1861 (O_1861,N_29762,N_29751);
or UO_1862 (O_1862,N_29813,N_29980);
nor UO_1863 (O_1863,N_29915,N_29791);
nand UO_1864 (O_1864,N_29786,N_29703);
nor UO_1865 (O_1865,N_29938,N_29800);
nor UO_1866 (O_1866,N_29721,N_29917);
and UO_1867 (O_1867,N_29859,N_29795);
nor UO_1868 (O_1868,N_29838,N_29897);
and UO_1869 (O_1869,N_29831,N_29966);
and UO_1870 (O_1870,N_29984,N_29969);
or UO_1871 (O_1871,N_29792,N_29887);
or UO_1872 (O_1872,N_29736,N_29788);
and UO_1873 (O_1873,N_29979,N_29848);
nor UO_1874 (O_1874,N_29777,N_29818);
or UO_1875 (O_1875,N_29944,N_29845);
nand UO_1876 (O_1876,N_29768,N_29847);
or UO_1877 (O_1877,N_29980,N_29732);
or UO_1878 (O_1878,N_29850,N_29967);
and UO_1879 (O_1879,N_29776,N_29726);
nand UO_1880 (O_1880,N_29892,N_29817);
nand UO_1881 (O_1881,N_29979,N_29919);
nand UO_1882 (O_1882,N_29981,N_29735);
or UO_1883 (O_1883,N_29732,N_29940);
xnor UO_1884 (O_1884,N_29793,N_29964);
xor UO_1885 (O_1885,N_29905,N_29719);
nand UO_1886 (O_1886,N_29799,N_29899);
nand UO_1887 (O_1887,N_29908,N_29980);
and UO_1888 (O_1888,N_29850,N_29729);
or UO_1889 (O_1889,N_29934,N_29977);
and UO_1890 (O_1890,N_29901,N_29889);
nor UO_1891 (O_1891,N_29771,N_29793);
nor UO_1892 (O_1892,N_29772,N_29958);
and UO_1893 (O_1893,N_29928,N_29992);
xor UO_1894 (O_1894,N_29914,N_29954);
xor UO_1895 (O_1895,N_29945,N_29755);
nand UO_1896 (O_1896,N_29791,N_29981);
or UO_1897 (O_1897,N_29957,N_29737);
or UO_1898 (O_1898,N_29707,N_29826);
or UO_1899 (O_1899,N_29987,N_29748);
and UO_1900 (O_1900,N_29778,N_29785);
nor UO_1901 (O_1901,N_29867,N_29915);
nor UO_1902 (O_1902,N_29850,N_29855);
or UO_1903 (O_1903,N_29724,N_29901);
nand UO_1904 (O_1904,N_29894,N_29826);
xnor UO_1905 (O_1905,N_29822,N_29729);
nor UO_1906 (O_1906,N_29759,N_29905);
or UO_1907 (O_1907,N_29945,N_29795);
or UO_1908 (O_1908,N_29727,N_29940);
nand UO_1909 (O_1909,N_29787,N_29901);
nand UO_1910 (O_1910,N_29730,N_29843);
nand UO_1911 (O_1911,N_29978,N_29731);
or UO_1912 (O_1912,N_29928,N_29863);
and UO_1913 (O_1913,N_29741,N_29839);
nor UO_1914 (O_1914,N_29959,N_29847);
or UO_1915 (O_1915,N_29715,N_29820);
nor UO_1916 (O_1916,N_29739,N_29711);
and UO_1917 (O_1917,N_29922,N_29707);
xor UO_1918 (O_1918,N_29840,N_29953);
nor UO_1919 (O_1919,N_29796,N_29987);
nor UO_1920 (O_1920,N_29763,N_29948);
and UO_1921 (O_1921,N_29757,N_29764);
xnor UO_1922 (O_1922,N_29830,N_29913);
or UO_1923 (O_1923,N_29914,N_29730);
xor UO_1924 (O_1924,N_29820,N_29743);
or UO_1925 (O_1925,N_29887,N_29953);
or UO_1926 (O_1926,N_29824,N_29720);
xor UO_1927 (O_1927,N_29759,N_29973);
xor UO_1928 (O_1928,N_29786,N_29824);
and UO_1929 (O_1929,N_29917,N_29874);
nor UO_1930 (O_1930,N_29860,N_29911);
or UO_1931 (O_1931,N_29918,N_29793);
nor UO_1932 (O_1932,N_29882,N_29894);
xor UO_1933 (O_1933,N_29916,N_29885);
nor UO_1934 (O_1934,N_29758,N_29752);
or UO_1935 (O_1935,N_29974,N_29868);
and UO_1936 (O_1936,N_29708,N_29864);
nand UO_1937 (O_1937,N_29976,N_29827);
nor UO_1938 (O_1938,N_29716,N_29857);
nand UO_1939 (O_1939,N_29733,N_29865);
nand UO_1940 (O_1940,N_29989,N_29757);
nand UO_1941 (O_1941,N_29978,N_29765);
xor UO_1942 (O_1942,N_29752,N_29930);
and UO_1943 (O_1943,N_29721,N_29794);
nand UO_1944 (O_1944,N_29894,N_29748);
nand UO_1945 (O_1945,N_29722,N_29874);
nand UO_1946 (O_1946,N_29855,N_29946);
and UO_1947 (O_1947,N_29969,N_29944);
nor UO_1948 (O_1948,N_29840,N_29834);
xor UO_1949 (O_1949,N_29780,N_29799);
xnor UO_1950 (O_1950,N_29840,N_29870);
nor UO_1951 (O_1951,N_29826,N_29927);
nand UO_1952 (O_1952,N_29793,N_29842);
nand UO_1953 (O_1953,N_29703,N_29772);
and UO_1954 (O_1954,N_29866,N_29822);
xor UO_1955 (O_1955,N_29831,N_29904);
or UO_1956 (O_1956,N_29929,N_29817);
and UO_1957 (O_1957,N_29981,N_29793);
and UO_1958 (O_1958,N_29974,N_29906);
or UO_1959 (O_1959,N_29818,N_29842);
or UO_1960 (O_1960,N_29909,N_29936);
nand UO_1961 (O_1961,N_29837,N_29788);
and UO_1962 (O_1962,N_29923,N_29939);
nand UO_1963 (O_1963,N_29914,N_29702);
or UO_1964 (O_1964,N_29857,N_29915);
and UO_1965 (O_1965,N_29706,N_29704);
or UO_1966 (O_1966,N_29726,N_29859);
nor UO_1967 (O_1967,N_29776,N_29948);
or UO_1968 (O_1968,N_29831,N_29846);
nor UO_1969 (O_1969,N_29787,N_29998);
nand UO_1970 (O_1970,N_29706,N_29733);
and UO_1971 (O_1971,N_29981,N_29976);
and UO_1972 (O_1972,N_29880,N_29952);
nand UO_1973 (O_1973,N_29827,N_29820);
or UO_1974 (O_1974,N_29849,N_29725);
xnor UO_1975 (O_1975,N_29820,N_29729);
or UO_1976 (O_1976,N_29741,N_29762);
nor UO_1977 (O_1977,N_29944,N_29975);
and UO_1978 (O_1978,N_29769,N_29994);
and UO_1979 (O_1979,N_29772,N_29891);
xor UO_1980 (O_1980,N_29963,N_29985);
xnor UO_1981 (O_1981,N_29712,N_29916);
or UO_1982 (O_1982,N_29884,N_29866);
xnor UO_1983 (O_1983,N_29724,N_29747);
nand UO_1984 (O_1984,N_29775,N_29786);
nand UO_1985 (O_1985,N_29803,N_29746);
nand UO_1986 (O_1986,N_29996,N_29751);
and UO_1987 (O_1987,N_29787,N_29989);
or UO_1988 (O_1988,N_29746,N_29765);
nand UO_1989 (O_1989,N_29939,N_29782);
nor UO_1990 (O_1990,N_29857,N_29947);
xnor UO_1991 (O_1991,N_29905,N_29890);
and UO_1992 (O_1992,N_29968,N_29962);
or UO_1993 (O_1993,N_29790,N_29717);
nor UO_1994 (O_1994,N_29775,N_29832);
nor UO_1995 (O_1995,N_29703,N_29954);
xor UO_1996 (O_1996,N_29810,N_29798);
nand UO_1997 (O_1997,N_29763,N_29958);
nor UO_1998 (O_1998,N_29906,N_29787);
and UO_1999 (O_1999,N_29991,N_29963);
nand UO_2000 (O_2000,N_29943,N_29948);
nand UO_2001 (O_2001,N_29726,N_29900);
xnor UO_2002 (O_2002,N_29975,N_29810);
or UO_2003 (O_2003,N_29971,N_29864);
nor UO_2004 (O_2004,N_29712,N_29805);
nand UO_2005 (O_2005,N_29779,N_29929);
or UO_2006 (O_2006,N_29922,N_29953);
xnor UO_2007 (O_2007,N_29804,N_29893);
nor UO_2008 (O_2008,N_29955,N_29833);
or UO_2009 (O_2009,N_29733,N_29953);
or UO_2010 (O_2010,N_29743,N_29986);
nor UO_2011 (O_2011,N_29879,N_29833);
xnor UO_2012 (O_2012,N_29718,N_29941);
nand UO_2013 (O_2013,N_29930,N_29739);
nand UO_2014 (O_2014,N_29853,N_29833);
and UO_2015 (O_2015,N_29923,N_29709);
xnor UO_2016 (O_2016,N_29908,N_29931);
xnor UO_2017 (O_2017,N_29864,N_29861);
nor UO_2018 (O_2018,N_29997,N_29955);
and UO_2019 (O_2019,N_29752,N_29709);
xnor UO_2020 (O_2020,N_29902,N_29974);
or UO_2021 (O_2021,N_29751,N_29779);
nand UO_2022 (O_2022,N_29776,N_29923);
and UO_2023 (O_2023,N_29803,N_29824);
or UO_2024 (O_2024,N_29948,N_29775);
nor UO_2025 (O_2025,N_29734,N_29965);
and UO_2026 (O_2026,N_29742,N_29721);
nand UO_2027 (O_2027,N_29736,N_29861);
and UO_2028 (O_2028,N_29986,N_29951);
or UO_2029 (O_2029,N_29980,N_29832);
or UO_2030 (O_2030,N_29732,N_29958);
nor UO_2031 (O_2031,N_29901,N_29941);
and UO_2032 (O_2032,N_29922,N_29947);
or UO_2033 (O_2033,N_29927,N_29840);
xor UO_2034 (O_2034,N_29934,N_29891);
nor UO_2035 (O_2035,N_29871,N_29704);
or UO_2036 (O_2036,N_29928,N_29806);
nand UO_2037 (O_2037,N_29734,N_29827);
nand UO_2038 (O_2038,N_29990,N_29831);
or UO_2039 (O_2039,N_29924,N_29789);
nor UO_2040 (O_2040,N_29760,N_29810);
xor UO_2041 (O_2041,N_29859,N_29946);
nor UO_2042 (O_2042,N_29905,N_29995);
or UO_2043 (O_2043,N_29945,N_29793);
or UO_2044 (O_2044,N_29902,N_29754);
nor UO_2045 (O_2045,N_29939,N_29830);
xnor UO_2046 (O_2046,N_29858,N_29713);
and UO_2047 (O_2047,N_29914,N_29865);
or UO_2048 (O_2048,N_29798,N_29839);
or UO_2049 (O_2049,N_29935,N_29887);
or UO_2050 (O_2050,N_29789,N_29705);
and UO_2051 (O_2051,N_29854,N_29776);
and UO_2052 (O_2052,N_29901,N_29809);
and UO_2053 (O_2053,N_29702,N_29700);
and UO_2054 (O_2054,N_29892,N_29729);
xnor UO_2055 (O_2055,N_29844,N_29849);
xor UO_2056 (O_2056,N_29739,N_29821);
or UO_2057 (O_2057,N_29926,N_29953);
and UO_2058 (O_2058,N_29967,N_29816);
xor UO_2059 (O_2059,N_29851,N_29803);
nor UO_2060 (O_2060,N_29770,N_29967);
nor UO_2061 (O_2061,N_29721,N_29893);
xor UO_2062 (O_2062,N_29892,N_29893);
and UO_2063 (O_2063,N_29865,N_29949);
nand UO_2064 (O_2064,N_29960,N_29723);
or UO_2065 (O_2065,N_29913,N_29956);
or UO_2066 (O_2066,N_29838,N_29844);
and UO_2067 (O_2067,N_29745,N_29723);
xor UO_2068 (O_2068,N_29865,N_29787);
and UO_2069 (O_2069,N_29824,N_29979);
and UO_2070 (O_2070,N_29883,N_29843);
nand UO_2071 (O_2071,N_29850,N_29803);
nand UO_2072 (O_2072,N_29870,N_29884);
nor UO_2073 (O_2073,N_29750,N_29785);
or UO_2074 (O_2074,N_29775,N_29942);
nor UO_2075 (O_2075,N_29953,N_29874);
nor UO_2076 (O_2076,N_29802,N_29833);
nand UO_2077 (O_2077,N_29815,N_29877);
nand UO_2078 (O_2078,N_29735,N_29883);
and UO_2079 (O_2079,N_29971,N_29701);
or UO_2080 (O_2080,N_29704,N_29949);
nor UO_2081 (O_2081,N_29891,N_29863);
xnor UO_2082 (O_2082,N_29903,N_29712);
nand UO_2083 (O_2083,N_29991,N_29860);
and UO_2084 (O_2084,N_29979,N_29766);
and UO_2085 (O_2085,N_29701,N_29909);
and UO_2086 (O_2086,N_29829,N_29721);
nand UO_2087 (O_2087,N_29928,N_29934);
nand UO_2088 (O_2088,N_29767,N_29931);
xor UO_2089 (O_2089,N_29876,N_29920);
nor UO_2090 (O_2090,N_29868,N_29788);
xnor UO_2091 (O_2091,N_29844,N_29786);
nand UO_2092 (O_2092,N_29937,N_29898);
nor UO_2093 (O_2093,N_29721,N_29894);
nand UO_2094 (O_2094,N_29910,N_29880);
xor UO_2095 (O_2095,N_29790,N_29737);
nor UO_2096 (O_2096,N_29922,N_29771);
nor UO_2097 (O_2097,N_29967,N_29889);
xnor UO_2098 (O_2098,N_29832,N_29753);
xor UO_2099 (O_2099,N_29746,N_29837);
nand UO_2100 (O_2100,N_29887,N_29707);
and UO_2101 (O_2101,N_29775,N_29824);
and UO_2102 (O_2102,N_29921,N_29762);
nand UO_2103 (O_2103,N_29988,N_29713);
nand UO_2104 (O_2104,N_29852,N_29719);
or UO_2105 (O_2105,N_29848,N_29738);
nor UO_2106 (O_2106,N_29829,N_29847);
xnor UO_2107 (O_2107,N_29826,N_29739);
or UO_2108 (O_2108,N_29830,N_29874);
xor UO_2109 (O_2109,N_29712,N_29731);
or UO_2110 (O_2110,N_29773,N_29719);
nand UO_2111 (O_2111,N_29884,N_29719);
and UO_2112 (O_2112,N_29915,N_29951);
xnor UO_2113 (O_2113,N_29949,N_29950);
xor UO_2114 (O_2114,N_29792,N_29785);
xnor UO_2115 (O_2115,N_29910,N_29719);
nor UO_2116 (O_2116,N_29808,N_29846);
and UO_2117 (O_2117,N_29948,N_29823);
nor UO_2118 (O_2118,N_29783,N_29832);
and UO_2119 (O_2119,N_29857,N_29785);
nand UO_2120 (O_2120,N_29775,N_29715);
and UO_2121 (O_2121,N_29924,N_29711);
and UO_2122 (O_2122,N_29768,N_29924);
xnor UO_2123 (O_2123,N_29809,N_29973);
nand UO_2124 (O_2124,N_29781,N_29995);
or UO_2125 (O_2125,N_29987,N_29978);
nor UO_2126 (O_2126,N_29777,N_29797);
or UO_2127 (O_2127,N_29845,N_29987);
nand UO_2128 (O_2128,N_29916,N_29870);
xor UO_2129 (O_2129,N_29854,N_29875);
or UO_2130 (O_2130,N_29759,N_29936);
nand UO_2131 (O_2131,N_29859,N_29996);
or UO_2132 (O_2132,N_29700,N_29949);
or UO_2133 (O_2133,N_29954,N_29702);
nand UO_2134 (O_2134,N_29781,N_29968);
or UO_2135 (O_2135,N_29856,N_29968);
and UO_2136 (O_2136,N_29815,N_29750);
nor UO_2137 (O_2137,N_29941,N_29772);
or UO_2138 (O_2138,N_29816,N_29729);
xnor UO_2139 (O_2139,N_29846,N_29827);
or UO_2140 (O_2140,N_29996,N_29975);
nand UO_2141 (O_2141,N_29853,N_29788);
and UO_2142 (O_2142,N_29890,N_29846);
nand UO_2143 (O_2143,N_29825,N_29816);
xnor UO_2144 (O_2144,N_29843,N_29756);
or UO_2145 (O_2145,N_29854,N_29888);
nor UO_2146 (O_2146,N_29920,N_29952);
and UO_2147 (O_2147,N_29755,N_29831);
and UO_2148 (O_2148,N_29951,N_29883);
nor UO_2149 (O_2149,N_29826,N_29839);
or UO_2150 (O_2150,N_29905,N_29904);
nand UO_2151 (O_2151,N_29709,N_29726);
nand UO_2152 (O_2152,N_29835,N_29779);
nand UO_2153 (O_2153,N_29866,N_29780);
nand UO_2154 (O_2154,N_29844,N_29754);
and UO_2155 (O_2155,N_29888,N_29821);
xnor UO_2156 (O_2156,N_29736,N_29846);
and UO_2157 (O_2157,N_29703,N_29895);
xnor UO_2158 (O_2158,N_29838,N_29717);
and UO_2159 (O_2159,N_29853,N_29852);
xnor UO_2160 (O_2160,N_29754,N_29830);
nand UO_2161 (O_2161,N_29734,N_29717);
nand UO_2162 (O_2162,N_29943,N_29744);
and UO_2163 (O_2163,N_29924,N_29834);
nor UO_2164 (O_2164,N_29968,N_29976);
or UO_2165 (O_2165,N_29874,N_29994);
xor UO_2166 (O_2166,N_29715,N_29731);
or UO_2167 (O_2167,N_29957,N_29992);
or UO_2168 (O_2168,N_29841,N_29939);
nand UO_2169 (O_2169,N_29993,N_29908);
or UO_2170 (O_2170,N_29772,N_29838);
nand UO_2171 (O_2171,N_29716,N_29766);
xnor UO_2172 (O_2172,N_29993,N_29769);
nand UO_2173 (O_2173,N_29890,N_29754);
xnor UO_2174 (O_2174,N_29882,N_29872);
nor UO_2175 (O_2175,N_29941,N_29850);
and UO_2176 (O_2176,N_29734,N_29922);
and UO_2177 (O_2177,N_29840,N_29906);
or UO_2178 (O_2178,N_29814,N_29882);
nand UO_2179 (O_2179,N_29953,N_29811);
xnor UO_2180 (O_2180,N_29700,N_29722);
nand UO_2181 (O_2181,N_29801,N_29819);
and UO_2182 (O_2182,N_29715,N_29987);
nand UO_2183 (O_2183,N_29956,N_29798);
nor UO_2184 (O_2184,N_29830,N_29757);
or UO_2185 (O_2185,N_29729,N_29861);
nor UO_2186 (O_2186,N_29894,N_29814);
xor UO_2187 (O_2187,N_29956,N_29865);
xor UO_2188 (O_2188,N_29734,N_29984);
nand UO_2189 (O_2189,N_29898,N_29958);
nor UO_2190 (O_2190,N_29709,N_29955);
and UO_2191 (O_2191,N_29909,N_29719);
nor UO_2192 (O_2192,N_29972,N_29700);
nand UO_2193 (O_2193,N_29863,N_29956);
nor UO_2194 (O_2194,N_29929,N_29985);
xnor UO_2195 (O_2195,N_29982,N_29823);
or UO_2196 (O_2196,N_29836,N_29832);
xnor UO_2197 (O_2197,N_29701,N_29922);
or UO_2198 (O_2198,N_29827,N_29701);
xnor UO_2199 (O_2199,N_29807,N_29774);
nor UO_2200 (O_2200,N_29955,N_29974);
and UO_2201 (O_2201,N_29882,N_29733);
and UO_2202 (O_2202,N_29712,N_29850);
nor UO_2203 (O_2203,N_29809,N_29770);
or UO_2204 (O_2204,N_29983,N_29921);
nand UO_2205 (O_2205,N_29727,N_29741);
and UO_2206 (O_2206,N_29974,N_29891);
nand UO_2207 (O_2207,N_29810,N_29957);
and UO_2208 (O_2208,N_29792,N_29799);
or UO_2209 (O_2209,N_29968,N_29934);
and UO_2210 (O_2210,N_29872,N_29743);
nand UO_2211 (O_2211,N_29786,N_29849);
xnor UO_2212 (O_2212,N_29704,N_29893);
or UO_2213 (O_2213,N_29810,N_29813);
nor UO_2214 (O_2214,N_29899,N_29882);
and UO_2215 (O_2215,N_29824,N_29928);
nand UO_2216 (O_2216,N_29852,N_29743);
nand UO_2217 (O_2217,N_29700,N_29983);
and UO_2218 (O_2218,N_29748,N_29908);
or UO_2219 (O_2219,N_29952,N_29801);
or UO_2220 (O_2220,N_29960,N_29819);
or UO_2221 (O_2221,N_29896,N_29704);
nor UO_2222 (O_2222,N_29712,N_29759);
nor UO_2223 (O_2223,N_29914,N_29763);
or UO_2224 (O_2224,N_29964,N_29925);
or UO_2225 (O_2225,N_29704,N_29796);
nand UO_2226 (O_2226,N_29758,N_29857);
and UO_2227 (O_2227,N_29923,N_29702);
or UO_2228 (O_2228,N_29816,N_29973);
or UO_2229 (O_2229,N_29807,N_29818);
and UO_2230 (O_2230,N_29808,N_29806);
xor UO_2231 (O_2231,N_29975,N_29702);
nand UO_2232 (O_2232,N_29904,N_29736);
nor UO_2233 (O_2233,N_29893,N_29778);
nand UO_2234 (O_2234,N_29722,N_29941);
xnor UO_2235 (O_2235,N_29989,N_29944);
or UO_2236 (O_2236,N_29939,N_29974);
xnor UO_2237 (O_2237,N_29715,N_29823);
nor UO_2238 (O_2238,N_29757,N_29889);
nand UO_2239 (O_2239,N_29880,N_29859);
or UO_2240 (O_2240,N_29996,N_29969);
nand UO_2241 (O_2241,N_29713,N_29922);
nand UO_2242 (O_2242,N_29914,N_29937);
and UO_2243 (O_2243,N_29782,N_29763);
xnor UO_2244 (O_2244,N_29928,N_29718);
and UO_2245 (O_2245,N_29983,N_29782);
nand UO_2246 (O_2246,N_29988,N_29925);
or UO_2247 (O_2247,N_29804,N_29802);
and UO_2248 (O_2248,N_29958,N_29868);
xnor UO_2249 (O_2249,N_29816,N_29873);
nand UO_2250 (O_2250,N_29898,N_29934);
and UO_2251 (O_2251,N_29952,N_29731);
or UO_2252 (O_2252,N_29809,N_29816);
or UO_2253 (O_2253,N_29910,N_29783);
xor UO_2254 (O_2254,N_29971,N_29839);
xor UO_2255 (O_2255,N_29814,N_29844);
nor UO_2256 (O_2256,N_29819,N_29968);
nor UO_2257 (O_2257,N_29751,N_29880);
nor UO_2258 (O_2258,N_29815,N_29764);
nand UO_2259 (O_2259,N_29987,N_29900);
nor UO_2260 (O_2260,N_29847,N_29917);
nor UO_2261 (O_2261,N_29806,N_29811);
nor UO_2262 (O_2262,N_29889,N_29777);
or UO_2263 (O_2263,N_29822,N_29916);
xnor UO_2264 (O_2264,N_29797,N_29869);
or UO_2265 (O_2265,N_29808,N_29906);
xnor UO_2266 (O_2266,N_29924,N_29726);
or UO_2267 (O_2267,N_29924,N_29701);
and UO_2268 (O_2268,N_29801,N_29918);
nand UO_2269 (O_2269,N_29800,N_29746);
xor UO_2270 (O_2270,N_29826,N_29901);
nand UO_2271 (O_2271,N_29804,N_29735);
nor UO_2272 (O_2272,N_29832,N_29763);
or UO_2273 (O_2273,N_29754,N_29901);
nand UO_2274 (O_2274,N_29953,N_29705);
nor UO_2275 (O_2275,N_29983,N_29898);
nor UO_2276 (O_2276,N_29812,N_29702);
or UO_2277 (O_2277,N_29865,N_29976);
xnor UO_2278 (O_2278,N_29908,N_29991);
and UO_2279 (O_2279,N_29766,N_29799);
or UO_2280 (O_2280,N_29801,N_29767);
nand UO_2281 (O_2281,N_29823,N_29842);
nor UO_2282 (O_2282,N_29863,N_29709);
and UO_2283 (O_2283,N_29740,N_29777);
xor UO_2284 (O_2284,N_29861,N_29820);
and UO_2285 (O_2285,N_29945,N_29819);
and UO_2286 (O_2286,N_29834,N_29967);
nand UO_2287 (O_2287,N_29776,N_29880);
xnor UO_2288 (O_2288,N_29988,N_29731);
nand UO_2289 (O_2289,N_29963,N_29787);
nand UO_2290 (O_2290,N_29866,N_29894);
nand UO_2291 (O_2291,N_29792,N_29725);
nand UO_2292 (O_2292,N_29844,N_29987);
or UO_2293 (O_2293,N_29769,N_29732);
nor UO_2294 (O_2294,N_29960,N_29914);
or UO_2295 (O_2295,N_29872,N_29919);
xnor UO_2296 (O_2296,N_29896,N_29909);
and UO_2297 (O_2297,N_29701,N_29864);
xnor UO_2298 (O_2298,N_29944,N_29949);
xnor UO_2299 (O_2299,N_29961,N_29706);
and UO_2300 (O_2300,N_29778,N_29849);
or UO_2301 (O_2301,N_29965,N_29700);
nand UO_2302 (O_2302,N_29873,N_29927);
nor UO_2303 (O_2303,N_29899,N_29746);
or UO_2304 (O_2304,N_29712,N_29883);
nor UO_2305 (O_2305,N_29746,N_29880);
nor UO_2306 (O_2306,N_29809,N_29864);
xnor UO_2307 (O_2307,N_29723,N_29917);
or UO_2308 (O_2308,N_29862,N_29748);
nand UO_2309 (O_2309,N_29717,N_29738);
and UO_2310 (O_2310,N_29924,N_29740);
or UO_2311 (O_2311,N_29810,N_29968);
or UO_2312 (O_2312,N_29964,N_29770);
and UO_2313 (O_2313,N_29903,N_29944);
xor UO_2314 (O_2314,N_29708,N_29870);
nand UO_2315 (O_2315,N_29723,N_29845);
or UO_2316 (O_2316,N_29851,N_29922);
nand UO_2317 (O_2317,N_29782,N_29821);
or UO_2318 (O_2318,N_29713,N_29901);
or UO_2319 (O_2319,N_29792,N_29888);
or UO_2320 (O_2320,N_29857,N_29782);
and UO_2321 (O_2321,N_29983,N_29773);
xor UO_2322 (O_2322,N_29724,N_29995);
and UO_2323 (O_2323,N_29923,N_29798);
nand UO_2324 (O_2324,N_29818,N_29701);
nand UO_2325 (O_2325,N_29879,N_29792);
nand UO_2326 (O_2326,N_29817,N_29894);
or UO_2327 (O_2327,N_29886,N_29812);
and UO_2328 (O_2328,N_29707,N_29934);
nand UO_2329 (O_2329,N_29899,N_29801);
nor UO_2330 (O_2330,N_29776,N_29929);
or UO_2331 (O_2331,N_29943,N_29978);
xor UO_2332 (O_2332,N_29841,N_29701);
or UO_2333 (O_2333,N_29818,N_29998);
or UO_2334 (O_2334,N_29771,N_29961);
nor UO_2335 (O_2335,N_29884,N_29952);
and UO_2336 (O_2336,N_29796,N_29798);
nand UO_2337 (O_2337,N_29906,N_29777);
xor UO_2338 (O_2338,N_29938,N_29935);
or UO_2339 (O_2339,N_29844,N_29823);
nor UO_2340 (O_2340,N_29942,N_29952);
xor UO_2341 (O_2341,N_29888,N_29814);
xnor UO_2342 (O_2342,N_29773,N_29735);
nand UO_2343 (O_2343,N_29771,N_29943);
xor UO_2344 (O_2344,N_29761,N_29756);
nor UO_2345 (O_2345,N_29870,N_29905);
and UO_2346 (O_2346,N_29891,N_29836);
and UO_2347 (O_2347,N_29895,N_29861);
xnor UO_2348 (O_2348,N_29752,N_29792);
nor UO_2349 (O_2349,N_29801,N_29911);
or UO_2350 (O_2350,N_29783,N_29883);
or UO_2351 (O_2351,N_29946,N_29911);
xor UO_2352 (O_2352,N_29943,N_29940);
nor UO_2353 (O_2353,N_29858,N_29960);
nand UO_2354 (O_2354,N_29861,N_29721);
nor UO_2355 (O_2355,N_29779,N_29982);
xor UO_2356 (O_2356,N_29983,N_29948);
and UO_2357 (O_2357,N_29975,N_29928);
xor UO_2358 (O_2358,N_29781,N_29712);
xor UO_2359 (O_2359,N_29860,N_29767);
and UO_2360 (O_2360,N_29961,N_29955);
or UO_2361 (O_2361,N_29707,N_29784);
or UO_2362 (O_2362,N_29996,N_29834);
and UO_2363 (O_2363,N_29828,N_29982);
nor UO_2364 (O_2364,N_29720,N_29943);
xor UO_2365 (O_2365,N_29812,N_29921);
or UO_2366 (O_2366,N_29798,N_29744);
or UO_2367 (O_2367,N_29755,N_29915);
or UO_2368 (O_2368,N_29892,N_29919);
nor UO_2369 (O_2369,N_29960,N_29749);
xor UO_2370 (O_2370,N_29794,N_29777);
nand UO_2371 (O_2371,N_29795,N_29824);
nor UO_2372 (O_2372,N_29816,N_29884);
and UO_2373 (O_2373,N_29986,N_29994);
or UO_2374 (O_2374,N_29803,N_29751);
nand UO_2375 (O_2375,N_29703,N_29882);
and UO_2376 (O_2376,N_29928,N_29813);
nand UO_2377 (O_2377,N_29712,N_29706);
nor UO_2378 (O_2378,N_29823,N_29782);
xor UO_2379 (O_2379,N_29706,N_29810);
and UO_2380 (O_2380,N_29860,N_29787);
and UO_2381 (O_2381,N_29976,N_29907);
nand UO_2382 (O_2382,N_29765,N_29983);
or UO_2383 (O_2383,N_29715,N_29913);
and UO_2384 (O_2384,N_29969,N_29932);
and UO_2385 (O_2385,N_29891,N_29955);
nor UO_2386 (O_2386,N_29878,N_29812);
nand UO_2387 (O_2387,N_29917,N_29935);
nand UO_2388 (O_2388,N_29789,N_29814);
and UO_2389 (O_2389,N_29704,N_29998);
xnor UO_2390 (O_2390,N_29726,N_29952);
or UO_2391 (O_2391,N_29840,N_29751);
nand UO_2392 (O_2392,N_29893,N_29912);
xor UO_2393 (O_2393,N_29988,N_29918);
or UO_2394 (O_2394,N_29815,N_29990);
nor UO_2395 (O_2395,N_29863,N_29831);
and UO_2396 (O_2396,N_29856,N_29773);
nand UO_2397 (O_2397,N_29743,N_29832);
nor UO_2398 (O_2398,N_29729,N_29818);
nand UO_2399 (O_2399,N_29922,N_29936);
xnor UO_2400 (O_2400,N_29891,N_29725);
or UO_2401 (O_2401,N_29874,N_29755);
or UO_2402 (O_2402,N_29871,N_29875);
nor UO_2403 (O_2403,N_29805,N_29770);
or UO_2404 (O_2404,N_29718,N_29831);
nor UO_2405 (O_2405,N_29846,N_29863);
nand UO_2406 (O_2406,N_29714,N_29878);
or UO_2407 (O_2407,N_29834,N_29731);
xor UO_2408 (O_2408,N_29802,N_29829);
and UO_2409 (O_2409,N_29909,N_29923);
or UO_2410 (O_2410,N_29754,N_29723);
nor UO_2411 (O_2411,N_29958,N_29985);
and UO_2412 (O_2412,N_29802,N_29935);
and UO_2413 (O_2413,N_29918,N_29961);
nor UO_2414 (O_2414,N_29777,N_29939);
nand UO_2415 (O_2415,N_29750,N_29854);
nand UO_2416 (O_2416,N_29725,N_29965);
nor UO_2417 (O_2417,N_29864,N_29836);
nor UO_2418 (O_2418,N_29719,N_29899);
nor UO_2419 (O_2419,N_29796,N_29862);
or UO_2420 (O_2420,N_29832,N_29817);
or UO_2421 (O_2421,N_29802,N_29813);
or UO_2422 (O_2422,N_29962,N_29896);
nor UO_2423 (O_2423,N_29952,N_29713);
nor UO_2424 (O_2424,N_29911,N_29955);
or UO_2425 (O_2425,N_29929,N_29983);
xnor UO_2426 (O_2426,N_29811,N_29851);
xor UO_2427 (O_2427,N_29999,N_29753);
xor UO_2428 (O_2428,N_29808,N_29815);
nand UO_2429 (O_2429,N_29909,N_29707);
nand UO_2430 (O_2430,N_29894,N_29982);
xor UO_2431 (O_2431,N_29756,N_29710);
nand UO_2432 (O_2432,N_29954,N_29816);
nor UO_2433 (O_2433,N_29901,N_29989);
xnor UO_2434 (O_2434,N_29978,N_29961);
xnor UO_2435 (O_2435,N_29703,N_29905);
or UO_2436 (O_2436,N_29832,N_29808);
nor UO_2437 (O_2437,N_29740,N_29884);
or UO_2438 (O_2438,N_29834,N_29868);
or UO_2439 (O_2439,N_29855,N_29792);
nor UO_2440 (O_2440,N_29944,N_29795);
and UO_2441 (O_2441,N_29907,N_29757);
nor UO_2442 (O_2442,N_29966,N_29903);
nand UO_2443 (O_2443,N_29782,N_29898);
xnor UO_2444 (O_2444,N_29710,N_29799);
and UO_2445 (O_2445,N_29899,N_29918);
nand UO_2446 (O_2446,N_29759,N_29713);
nor UO_2447 (O_2447,N_29757,N_29951);
nand UO_2448 (O_2448,N_29915,N_29925);
nand UO_2449 (O_2449,N_29910,N_29921);
nand UO_2450 (O_2450,N_29927,N_29949);
and UO_2451 (O_2451,N_29961,N_29766);
or UO_2452 (O_2452,N_29713,N_29981);
or UO_2453 (O_2453,N_29707,N_29950);
and UO_2454 (O_2454,N_29878,N_29819);
and UO_2455 (O_2455,N_29873,N_29729);
nand UO_2456 (O_2456,N_29829,N_29779);
and UO_2457 (O_2457,N_29822,N_29937);
or UO_2458 (O_2458,N_29899,N_29987);
or UO_2459 (O_2459,N_29887,N_29862);
and UO_2460 (O_2460,N_29728,N_29855);
and UO_2461 (O_2461,N_29894,N_29745);
nand UO_2462 (O_2462,N_29943,N_29848);
xnor UO_2463 (O_2463,N_29805,N_29740);
or UO_2464 (O_2464,N_29768,N_29848);
nand UO_2465 (O_2465,N_29805,N_29984);
or UO_2466 (O_2466,N_29943,N_29913);
and UO_2467 (O_2467,N_29930,N_29725);
or UO_2468 (O_2468,N_29945,N_29804);
xnor UO_2469 (O_2469,N_29763,N_29962);
xnor UO_2470 (O_2470,N_29705,N_29996);
or UO_2471 (O_2471,N_29728,N_29751);
nor UO_2472 (O_2472,N_29860,N_29977);
nor UO_2473 (O_2473,N_29927,N_29946);
and UO_2474 (O_2474,N_29811,N_29981);
and UO_2475 (O_2475,N_29998,N_29726);
xnor UO_2476 (O_2476,N_29809,N_29719);
or UO_2477 (O_2477,N_29997,N_29717);
nor UO_2478 (O_2478,N_29990,N_29833);
and UO_2479 (O_2479,N_29712,N_29765);
and UO_2480 (O_2480,N_29912,N_29918);
or UO_2481 (O_2481,N_29904,N_29834);
xnor UO_2482 (O_2482,N_29844,N_29738);
xor UO_2483 (O_2483,N_29721,N_29853);
and UO_2484 (O_2484,N_29967,N_29738);
xor UO_2485 (O_2485,N_29760,N_29982);
nor UO_2486 (O_2486,N_29860,N_29797);
and UO_2487 (O_2487,N_29747,N_29823);
nand UO_2488 (O_2488,N_29726,N_29825);
nor UO_2489 (O_2489,N_29763,N_29866);
nand UO_2490 (O_2490,N_29709,N_29795);
and UO_2491 (O_2491,N_29961,N_29707);
nand UO_2492 (O_2492,N_29737,N_29868);
nand UO_2493 (O_2493,N_29988,N_29863);
xnor UO_2494 (O_2494,N_29830,N_29746);
nand UO_2495 (O_2495,N_29763,N_29820);
or UO_2496 (O_2496,N_29960,N_29805);
and UO_2497 (O_2497,N_29806,N_29955);
xor UO_2498 (O_2498,N_29853,N_29934);
xor UO_2499 (O_2499,N_29937,N_29793);
nand UO_2500 (O_2500,N_29716,N_29990);
nand UO_2501 (O_2501,N_29881,N_29875);
and UO_2502 (O_2502,N_29989,N_29735);
nor UO_2503 (O_2503,N_29929,N_29870);
nand UO_2504 (O_2504,N_29732,N_29704);
and UO_2505 (O_2505,N_29901,N_29926);
nand UO_2506 (O_2506,N_29785,N_29910);
nor UO_2507 (O_2507,N_29889,N_29992);
xor UO_2508 (O_2508,N_29887,N_29976);
xor UO_2509 (O_2509,N_29936,N_29966);
xnor UO_2510 (O_2510,N_29726,N_29735);
nor UO_2511 (O_2511,N_29735,N_29794);
nand UO_2512 (O_2512,N_29962,N_29929);
or UO_2513 (O_2513,N_29844,N_29842);
nand UO_2514 (O_2514,N_29877,N_29915);
nand UO_2515 (O_2515,N_29774,N_29883);
xnor UO_2516 (O_2516,N_29852,N_29854);
nand UO_2517 (O_2517,N_29710,N_29707);
xnor UO_2518 (O_2518,N_29724,N_29709);
or UO_2519 (O_2519,N_29970,N_29986);
xor UO_2520 (O_2520,N_29834,N_29960);
nor UO_2521 (O_2521,N_29702,N_29919);
and UO_2522 (O_2522,N_29930,N_29906);
and UO_2523 (O_2523,N_29772,N_29753);
nor UO_2524 (O_2524,N_29788,N_29980);
and UO_2525 (O_2525,N_29744,N_29933);
and UO_2526 (O_2526,N_29960,N_29897);
and UO_2527 (O_2527,N_29792,N_29876);
or UO_2528 (O_2528,N_29714,N_29908);
xor UO_2529 (O_2529,N_29900,N_29907);
nor UO_2530 (O_2530,N_29924,N_29942);
and UO_2531 (O_2531,N_29845,N_29705);
and UO_2532 (O_2532,N_29739,N_29830);
xnor UO_2533 (O_2533,N_29777,N_29774);
nor UO_2534 (O_2534,N_29734,N_29903);
nand UO_2535 (O_2535,N_29732,N_29711);
xnor UO_2536 (O_2536,N_29789,N_29884);
or UO_2537 (O_2537,N_29767,N_29732);
or UO_2538 (O_2538,N_29817,N_29853);
or UO_2539 (O_2539,N_29739,N_29953);
nand UO_2540 (O_2540,N_29818,N_29730);
or UO_2541 (O_2541,N_29947,N_29866);
and UO_2542 (O_2542,N_29774,N_29799);
and UO_2543 (O_2543,N_29732,N_29701);
and UO_2544 (O_2544,N_29860,N_29955);
nor UO_2545 (O_2545,N_29758,N_29732);
xor UO_2546 (O_2546,N_29990,N_29865);
and UO_2547 (O_2547,N_29969,N_29863);
and UO_2548 (O_2548,N_29955,N_29884);
and UO_2549 (O_2549,N_29863,N_29938);
nand UO_2550 (O_2550,N_29853,N_29767);
nand UO_2551 (O_2551,N_29740,N_29746);
and UO_2552 (O_2552,N_29842,N_29846);
nand UO_2553 (O_2553,N_29997,N_29943);
or UO_2554 (O_2554,N_29993,N_29914);
nand UO_2555 (O_2555,N_29946,N_29849);
or UO_2556 (O_2556,N_29984,N_29890);
or UO_2557 (O_2557,N_29750,N_29824);
nand UO_2558 (O_2558,N_29902,N_29708);
or UO_2559 (O_2559,N_29799,N_29746);
nand UO_2560 (O_2560,N_29870,N_29760);
and UO_2561 (O_2561,N_29779,N_29711);
nand UO_2562 (O_2562,N_29833,N_29976);
or UO_2563 (O_2563,N_29780,N_29718);
nand UO_2564 (O_2564,N_29829,N_29715);
xor UO_2565 (O_2565,N_29725,N_29711);
nand UO_2566 (O_2566,N_29804,N_29991);
xor UO_2567 (O_2567,N_29967,N_29937);
nor UO_2568 (O_2568,N_29847,N_29890);
and UO_2569 (O_2569,N_29775,N_29730);
nand UO_2570 (O_2570,N_29880,N_29815);
nand UO_2571 (O_2571,N_29889,N_29820);
nor UO_2572 (O_2572,N_29922,N_29736);
and UO_2573 (O_2573,N_29923,N_29944);
xnor UO_2574 (O_2574,N_29896,N_29814);
nand UO_2575 (O_2575,N_29920,N_29865);
nor UO_2576 (O_2576,N_29751,N_29776);
or UO_2577 (O_2577,N_29836,N_29934);
or UO_2578 (O_2578,N_29750,N_29926);
nor UO_2579 (O_2579,N_29745,N_29765);
and UO_2580 (O_2580,N_29890,N_29700);
or UO_2581 (O_2581,N_29908,N_29804);
nand UO_2582 (O_2582,N_29833,N_29820);
nand UO_2583 (O_2583,N_29859,N_29803);
xor UO_2584 (O_2584,N_29874,N_29836);
xnor UO_2585 (O_2585,N_29826,N_29814);
nor UO_2586 (O_2586,N_29799,N_29714);
nor UO_2587 (O_2587,N_29926,N_29891);
or UO_2588 (O_2588,N_29963,N_29935);
or UO_2589 (O_2589,N_29886,N_29922);
and UO_2590 (O_2590,N_29703,N_29910);
xor UO_2591 (O_2591,N_29974,N_29733);
or UO_2592 (O_2592,N_29852,N_29953);
or UO_2593 (O_2593,N_29700,N_29798);
and UO_2594 (O_2594,N_29744,N_29763);
nand UO_2595 (O_2595,N_29811,N_29908);
and UO_2596 (O_2596,N_29759,N_29868);
and UO_2597 (O_2597,N_29768,N_29777);
nand UO_2598 (O_2598,N_29999,N_29930);
xnor UO_2599 (O_2599,N_29710,N_29818);
or UO_2600 (O_2600,N_29998,N_29940);
and UO_2601 (O_2601,N_29715,N_29892);
or UO_2602 (O_2602,N_29995,N_29749);
xor UO_2603 (O_2603,N_29811,N_29979);
nor UO_2604 (O_2604,N_29762,N_29899);
nor UO_2605 (O_2605,N_29764,N_29712);
xor UO_2606 (O_2606,N_29943,N_29912);
and UO_2607 (O_2607,N_29997,N_29989);
and UO_2608 (O_2608,N_29767,N_29798);
and UO_2609 (O_2609,N_29986,N_29897);
nand UO_2610 (O_2610,N_29817,N_29913);
xnor UO_2611 (O_2611,N_29998,N_29724);
or UO_2612 (O_2612,N_29881,N_29753);
nor UO_2613 (O_2613,N_29875,N_29945);
xor UO_2614 (O_2614,N_29946,N_29744);
or UO_2615 (O_2615,N_29925,N_29913);
xnor UO_2616 (O_2616,N_29833,N_29856);
xor UO_2617 (O_2617,N_29909,N_29790);
xnor UO_2618 (O_2618,N_29797,N_29779);
nor UO_2619 (O_2619,N_29885,N_29834);
nor UO_2620 (O_2620,N_29983,N_29908);
and UO_2621 (O_2621,N_29718,N_29816);
nor UO_2622 (O_2622,N_29796,N_29731);
or UO_2623 (O_2623,N_29814,N_29868);
nor UO_2624 (O_2624,N_29805,N_29759);
and UO_2625 (O_2625,N_29863,N_29992);
and UO_2626 (O_2626,N_29735,N_29974);
nand UO_2627 (O_2627,N_29807,N_29893);
xor UO_2628 (O_2628,N_29907,N_29908);
nand UO_2629 (O_2629,N_29800,N_29828);
xnor UO_2630 (O_2630,N_29898,N_29909);
and UO_2631 (O_2631,N_29889,N_29926);
and UO_2632 (O_2632,N_29773,N_29774);
nand UO_2633 (O_2633,N_29848,N_29867);
and UO_2634 (O_2634,N_29819,N_29774);
xnor UO_2635 (O_2635,N_29732,N_29763);
nor UO_2636 (O_2636,N_29736,N_29960);
or UO_2637 (O_2637,N_29733,N_29779);
nand UO_2638 (O_2638,N_29845,N_29958);
nor UO_2639 (O_2639,N_29799,N_29718);
nor UO_2640 (O_2640,N_29929,N_29890);
or UO_2641 (O_2641,N_29980,N_29953);
or UO_2642 (O_2642,N_29750,N_29873);
nand UO_2643 (O_2643,N_29971,N_29789);
or UO_2644 (O_2644,N_29701,N_29723);
xor UO_2645 (O_2645,N_29962,N_29776);
and UO_2646 (O_2646,N_29767,N_29758);
and UO_2647 (O_2647,N_29963,N_29965);
nor UO_2648 (O_2648,N_29787,N_29940);
nor UO_2649 (O_2649,N_29782,N_29938);
and UO_2650 (O_2650,N_29809,N_29776);
and UO_2651 (O_2651,N_29981,N_29877);
xor UO_2652 (O_2652,N_29700,N_29841);
nor UO_2653 (O_2653,N_29989,N_29751);
nand UO_2654 (O_2654,N_29816,N_29984);
or UO_2655 (O_2655,N_29796,N_29898);
nand UO_2656 (O_2656,N_29905,N_29913);
nor UO_2657 (O_2657,N_29800,N_29837);
or UO_2658 (O_2658,N_29913,N_29739);
nor UO_2659 (O_2659,N_29933,N_29749);
nand UO_2660 (O_2660,N_29770,N_29890);
xor UO_2661 (O_2661,N_29964,N_29843);
nand UO_2662 (O_2662,N_29771,N_29748);
nand UO_2663 (O_2663,N_29859,N_29858);
nor UO_2664 (O_2664,N_29854,N_29944);
or UO_2665 (O_2665,N_29818,N_29736);
nor UO_2666 (O_2666,N_29844,N_29712);
nor UO_2667 (O_2667,N_29952,N_29734);
nand UO_2668 (O_2668,N_29982,N_29960);
and UO_2669 (O_2669,N_29882,N_29895);
xnor UO_2670 (O_2670,N_29928,N_29785);
and UO_2671 (O_2671,N_29858,N_29712);
xor UO_2672 (O_2672,N_29898,N_29936);
or UO_2673 (O_2673,N_29932,N_29882);
nor UO_2674 (O_2674,N_29806,N_29823);
and UO_2675 (O_2675,N_29756,N_29772);
nor UO_2676 (O_2676,N_29920,N_29929);
xor UO_2677 (O_2677,N_29858,N_29857);
nor UO_2678 (O_2678,N_29926,N_29739);
and UO_2679 (O_2679,N_29885,N_29888);
and UO_2680 (O_2680,N_29977,N_29759);
xor UO_2681 (O_2681,N_29809,N_29854);
xor UO_2682 (O_2682,N_29754,N_29752);
nand UO_2683 (O_2683,N_29966,N_29797);
nor UO_2684 (O_2684,N_29876,N_29782);
and UO_2685 (O_2685,N_29783,N_29746);
xnor UO_2686 (O_2686,N_29850,N_29937);
and UO_2687 (O_2687,N_29710,N_29782);
or UO_2688 (O_2688,N_29999,N_29976);
nand UO_2689 (O_2689,N_29780,N_29802);
xor UO_2690 (O_2690,N_29727,N_29938);
nand UO_2691 (O_2691,N_29706,N_29734);
and UO_2692 (O_2692,N_29811,N_29996);
nor UO_2693 (O_2693,N_29912,N_29935);
nor UO_2694 (O_2694,N_29919,N_29713);
nor UO_2695 (O_2695,N_29758,N_29899);
or UO_2696 (O_2696,N_29985,N_29821);
nand UO_2697 (O_2697,N_29856,N_29865);
nor UO_2698 (O_2698,N_29774,N_29857);
xnor UO_2699 (O_2699,N_29896,N_29836);
and UO_2700 (O_2700,N_29766,N_29751);
nand UO_2701 (O_2701,N_29908,N_29888);
nor UO_2702 (O_2702,N_29922,N_29855);
nand UO_2703 (O_2703,N_29770,N_29971);
and UO_2704 (O_2704,N_29726,N_29871);
nor UO_2705 (O_2705,N_29855,N_29911);
xor UO_2706 (O_2706,N_29885,N_29766);
and UO_2707 (O_2707,N_29807,N_29845);
nor UO_2708 (O_2708,N_29810,N_29900);
nand UO_2709 (O_2709,N_29841,N_29926);
xor UO_2710 (O_2710,N_29957,N_29908);
nor UO_2711 (O_2711,N_29893,N_29844);
or UO_2712 (O_2712,N_29711,N_29793);
nor UO_2713 (O_2713,N_29861,N_29774);
nor UO_2714 (O_2714,N_29802,N_29741);
xnor UO_2715 (O_2715,N_29941,N_29851);
or UO_2716 (O_2716,N_29986,N_29730);
xnor UO_2717 (O_2717,N_29833,N_29817);
xnor UO_2718 (O_2718,N_29818,N_29747);
nor UO_2719 (O_2719,N_29816,N_29999);
xnor UO_2720 (O_2720,N_29852,N_29713);
and UO_2721 (O_2721,N_29786,N_29833);
nor UO_2722 (O_2722,N_29994,N_29753);
and UO_2723 (O_2723,N_29953,N_29969);
nor UO_2724 (O_2724,N_29965,N_29792);
nand UO_2725 (O_2725,N_29750,N_29995);
or UO_2726 (O_2726,N_29967,N_29706);
xor UO_2727 (O_2727,N_29840,N_29713);
or UO_2728 (O_2728,N_29898,N_29753);
or UO_2729 (O_2729,N_29983,N_29876);
or UO_2730 (O_2730,N_29966,N_29933);
and UO_2731 (O_2731,N_29998,N_29925);
xnor UO_2732 (O_2732,N_29817,N_29969);
or UO_2733 (O_2733,N_29855,N_29714);
or UO_2734 (O_2734,N_29836,N_29961);
nand UO_2735 (O_2735,N_29920,N_29932);
nand UO_2736 (O_2736,N_29742,N_29782);
nor UO_2737 (O_2737,N_29965,N_29944);
xor UO_2738 (O_2738,N_29788,N_29774);
or UO_2739 (O_2739,N_29933,N_29703);
xnor UO_2740 (O_2740,N_29819,N_29721);
or UO_2741 (O_2741,N_29918,N_29945);
nand UO_2742 (O_2742,N_29914,N_29771);
or UO_2743 (O_2743,N_29978,N_29972);
nor UO_2744 (O_2744,N_29808,N_29872);
nand UO_2745 (O_2745,N_29716,N_29717);
xnor UO_2746 (O_2746,N_29904,N_29994);
and UO_2747 (O_2747,N_29906,N_29877);
nand UO_2748 (O_2748,N_29888,N_29817);
and UO_2749 (O_2749,N_29786,N_29985);
xnor UO_2750 (O_2750,N_29924,N_29985);
nor UO_2751 (O_2751,N_29821,N_29794);
nand UO_2752 (O_2752,N_29882,N_29721);
or UO_2753 (O_2753,N_29730,N_29897);
xor UO_2754 (O_2754,N_29881,N_29814);
or UO_2755 (O_2755,N_29713,N_29786);
and UO_2756 (O_2756,N_29983,N_29842);
or UO_2757 (O_2757,N_29872,N_29970);
nor UO_2758 (O_2758,N_29946,N_29779);
or UO_2759 (O_2759,N_29760,N_29877);
nor UO_2760 (O_2760,N_29906,N_29992);
nand UO_2761 (O_2761,N_29982,N_29961);
or UO_2762 (O_2762,N_29842,N_29917);
nor UO_2763 (O_2763,N_29994,N_29866);
and UO_2764 (O_2764,N_29930,N_29812);
nor UO_2765 (O_2765,N_29708,N_29936);
nand UO_2766 (O_2766,N_29941,N_29724);
xnor UO_2767 (O_2767,N_29928,N_29742);
and UO_2768 (O_2768,N_29926,N_29770);
or UO_2769 (O_2769,N_29896,N_29745);
nand UO_2770 (O_2770,N_29767,N_29718);
or UO_2771 (O_2771,N_29815,N_29930);
nor UO_2772 (O_2772,N_29821,N_29765);
and UO_2773 (O_2773,N_29928,N_29918);
or UO_2774 (O_2774,N_29726,N_29717);
and UO_2775 (O_2775,N_29795,N_29897);
nor UO_2776 (O_2776,N_29828,N_29864);
nor UO_2777 (O_2777,N_29954,N_29777);
nor UO_2778 (O_2778,N_29935,N_29910);
xor UO_2779 (O_2779,N_29818,N_29820);
nand UO_2780 (O_2780,N_29968,N_29896);
and UO_2781 (O_2781,N_29934,N_29967);
or UO_2782 (O_2782,N_29718,N_29878);
nor UO_2783 (O_2783,N_29784,N_29830);
and UO_2784 (O_2784,N_29880,N_29709);
xnor UO_2785 (O_2785,N_29712,N_29879);
and UO_2786 (O_2786,N_29909,N_29974);
and UO_2787 (O_2787,N_29956,N_29961);
nor UO_2788 (O_2788,N_29842,N_29708);
and UO_2789 (O_2789,N_29748,N_29821);
nor UO_2790 (O_2790,N_29863,N_29912);
or UO_2791 (O_2791,N_29728,N_29793);
and UO_2792 (O_2792,N_29701,N_29787);
xor UO_2793 (O_2793,N_29966,N_29809);
nand UO_2794 (O_2794,N_29700,N_29857);
xor UO_2795 (O_2795,N_29937,N_29981);
and UO_2796 (O_2796,N_29958,N_29877);
nor UO_2797 (O_2797,N_29838,N_29927);
xnor UO_2798 (O_2798,N_29845,N_29858);
or UO_2799 (O_2799,N_29739,N_29816);
and UO_2800 (O_2800,N_29927,N_29923);
xnor UO_2801 (O_2801,N_29832,N_29906);
nor UO_2802 (O_2802,N_29709,N_29898);
xnor UO_2803 (O_2803,N_29986,N_29983);
nand UO_2804 (O_2804,N_29850,N_29871);
nand UO_2805 (O_2805,N_29947,N_29890);
or UO_2806 (O_2806,N_29954,N_29751);
or UO_2807 (O_2807,N_29773,N_29897);
xnor UO_2808 (O_2808,N_29857,N_29958);
or UO_2809 (O_2809,N_29846,N_29950);
nand UO_2810 (O_2810,N_29991,N_29732);
nor UO_2811 (O_2811,N_29870,N_29746);
and UO_2812 (O_2812,N_29957,N_29701);
nand UO_2813 (O_2813,N_29938,N_29712);
xor UO_2814 (O_2814,N_29974,N_29760);
nor UO_2815 (O_2815,N_29703,N_29807);
and UO_2816 (O_2816,N_29848,N_29899);
xor UO_2817 (O_2817,N_29828,N_29922);
xor UO_2818 (O_2818,N_29813,N_29941);
nor UO_2819 (O_2819,N_29981,N_29804);
and UO_2820 (O_2820,N_29708,N_29981);
and UO_2821 (O_2821,N_29706,N_29926);
nor UO_2822 (O_2822,N_29711,N_29849);
and UO_2823 (O_2823,N_29718,N_29986);
or UO_2824 (O_2824,N_29866,N_29964);
or UO_2825 (O_2825,N_29960,N_29812);
nor UO_2826 (O_2826,N_29997,N_29897);
nor UO_2827 (O_2827,N_29865,N_29740);
xnor UO_2828 (O_2828,N_29892,N_29700);
xor UO_2829 (O_2829,N_29970,N_29796);
nor UO_2830 (O_2830,N_29797,N_29934);
nor UO_2831 (O_2831,N_29821,N_29828);
xnor UO_2832 (O_2832,N_29805,N_29934);
nand UO_2833 (O_2833,N_29861,N_29887);
nor UO_2834 (O_2834,N_29913,N_29769);
nand UO_2835 (O_2835,N_29735,N_29754);
or UO_2836 (O_2836,N_29862,N_29897);
and UO_2837 (O_2837,N_29791,N_29748);
xor UO_2838 (O_2838,N_29946,N_29906);
nor UO_2839 (O_2839,N_29817,N_29882);
and UO_2840 (O_2840,N_29913,N_29782);
xnor UO_2841 (O_2841,N_29971,N_29757);
or UO_2842 (O_2842,N_29738,N_29977);
and UO_2843 (O_2843,N_29702,N_29864);
nand UO_2844 (O_2844,N_29720,N_29854);
or UO_2845 (O_2845,N_29772,N_29818);
nor UO_2846 (O_2846,N_29974,N_29748);
xor UO_2847 (O_2847,N_29970,N_29873);
and UO_2848 (O_2848,N_29979,N_29797);
or UO_2849 (O_2849,N_29924,N_29865);
or UO_2850 (O_2850,N_29995,N_29855);
and UO_2851 (O_2851,N_29952,N_29719);
nor UO_2852 (O_2852,N_29981,N_29800);
and UO_2853 (O_2853,N_29896,N_29864);
nor UO_2854 (O_2854,N_29954,N_29936);
nand UO_2855 (O_2855,N_29964,N_29839);
or UO_2856 (O_2856,N_29739,N_29776);
xor UO_2857 (O_2857,N_29835,N_29877);
xor UO_2858 (O_2858,N_29969,N_29986);
or UO_2859 (O_2859,N_29712,N_29751);
or UO_2860 (O_2860,N_29987,N_29874);
or UO_2861 (O_2861,N_29701,N_29931);
and UO_2862 (O_2862,N_29922,N_29804);
or UO_2863 (O_2863,N_29753,N_29720);
nand UO_2864 (O_2864,N_29760,N_29965);
nor UO_2865 (O_2865,N_29982,N_29969);
xnor UO_2866 (O_2866,N_29747,N_29966);
nor UO_2867 (O_2867,N_29857,N_29824);
nor UO_2868 (O_2868,N_29811,N_29824);
nor UO_2869 (O_2869,N_29960,N_29926);
or UO_2870 (O_2870,N_29720,N_29965);
xor UO_2871 (O_2871,N_29858,N_29980);
nand UO_2872 (O_2872,N_29744,N_29952);
xnor UO_2873 (O_2873,N_29944,N_29846);
and UO_2874 (O_2874,N_29877,N_29837);
nand UO_2875 (O_2875,N_29904,N_29771);
or UO_2876 (O_2876,N_29926,N_29737);
xor UO_2877 (O_2877,N_29914,N_29741);
nand UO_2878 (O_2878,N_29844,N_29938);
and UO_2879 (O_2879,N_29889,N_29829);
xnor UO_2880 (O_2880,N_29782,N_29914);
and UO_2881 (O_2881,N_29845,N_29950);
and UO_2882 (O_2882,N_29858,N_29914);
xor UO_2883 (O_2883,N_29716,N_29802);
xnor UO_2884 (O_2884,N_29968,N_29805);
or UO_2885 (O_2885,N_29805,N_29902);
nand UO_2886 (O_2886,N_29930,N_29828);
and UO_2887 (O_2887,N_29867,N_29878);
and UO_2888 (O_2888,N_29725,N_29842);
or UO_2889 (O_2889,N_29831,N_29956);
xnor UO_2890 (O_2890,N_29957,N_29788);
or UO_2891 (O_2891,N_29881,N_29863);
nand UO_2892 (O_2892,N_29785,N_29950);
xor UO_2893 (O_2893,N_29891,N_29959);
nor UO_2894 (O_2894,N_29806,N_29707);
and UO_2895 (O_2895,N_29874,N_29919);
or UO_2896 (O_2896,N_29758,N_29805);
xnor UO_2897 (O_2897,N_29848,N_29860);
nor UO_2898 (O_2898,N_29910,N_29770);
nand UO_2899 (O_2899,N_29826,N_29710);
xnor UO_2900 (O_2900,N_29726,N_29920);
and UO_2901 (O_2901,N_29902,N_29740);
nor UO_2902 (O_2902,N_29717,N_29948);
nor UO_2903 (O_2903,N_29746,N_29755);
xnor UO_2904 (O_2904,N_29747,N_29847);
xor UO_2905 (O_2905,N_29799,N_29748);
and UO_2906 (O_2906,N_29854,N_29744);
nor UO_2907 (O_2907,N_29843,N_29975);
or UO_2908 (O_2908,N_29730,N_29974);
and UO_2909 (O_2909,N_29995,N_29734);
nand UO_2910 (O_2910,N_29903,N_29970);
nand UO_2911 (O_2911,N_29958,N_29713);
and UO_2912 (O_2912,N_29906,N_29701);
and UO_2913 (O_2913,N_29701,N_29811);
nand UO_2914 (O_2914,N_29834,N_29831);
nor UO_2915 (O_2915,N_29799,N_29827);
nand UO_2916 (O_2916,N_29766,N_29718);
nand UO_2917 (O_2917,N_29808,N_29782);
or UO_2918 (O_2918,N_29721,N_29944);
nor UO_2919 (O_2919,N_29916,N_29897);
nor UO_2920 (O_2920,N_29834,N_29875);
nand UO_2921 (O_2921,N_29871,N_29826);
xnor UO_2922 (O_2922,N_29943,N_29914);
and UO_2923 (O_2923,N_29975,N_29856);
nand UO_2924 (O_2924,N_29810,N_29793);
or UO_2925 (O_2925,N_29727,N_29701);
and UO_2926 (O_2926,N_29934,N_29900);
and UO_2927 (O_2927,N_29746,N_29963);
and UO_2928 (O_2928,N_29779,N_29806);
xnor UO_2929 (O_2929,N_29723,N_29772);
nor UO_2930 (O_2930,N_29916,N_29894);
nor UO_2931 (O_2931,N_29703,N_29788);
nor UO_2932 (O_2932,N_29730,N_29973);
nor UO_2933 (O_2933,N_29807,N_29868);
or UO_2934 (O_2934,N_29848,N_29919);
nand UO_2935 (O_2935,N_29915,N_29952);
and UO_2936 (O_2936,N_29714,N_29899);
and UO_2937 (O_2937,N_29939,N_29980);
nand UO_2938 (O_2938,N_29705,N_29849);
and UO_2939 (O_2939,N_29919,N_29975);
xor UO_2940 (O_2940,N_29882,N_29920);
xnor UO_2941 (O_2941,N_29915,N_29865);
or UO_2942 (O_2942,N_29890,N_29818);
nand UO_2943 (O_2943,N_29804,N_29897);
and UO_2944 (O_2944,N_29953,N_29860);
nor UO_2945 (O_2945,N_29870,N_29725);
or UO_2946 (O_2946,N_29970,N_29944);
nor UO_2947 (O_2947,N_29753,N_29940);
nor UO_2948 (O_2948,N_29821,N_29964);
nor UO_2949 (O_2949,N_29797,N_29984);
nor UO_2950 (O_2950,N_29951,N_29728);
or UO_2951 (O_2951,N_29854,N_29908);
nor UO_2952 (O_2952,N_29822,N_29770);
nor UO_2953 (O_2953,N_29850,N_29808);
or UO_2954 (O_2954,N_29701,N_29799);
xor UO_2955 (O_2955,N_29786,N_29891);
xor UO_2956 (O_2956,N_29714,N_29888);
and UO_2957 (O_2957,N_29756,N_29913);
and UO_2958 (O_2958,N_29906,N_29889);
and UO_2959 (O_2959,N_29990,N_29826);
xor UO_2960 (O_2960,N_29977,N_29737);
nand UO_2961 (O_2961,N_29822,N_29792);
nor UO_2962 (O_2962,N_29826,N_29946);
nand UO_2963 (O_2963,N_29967,N_29963);
or UO_2964 (O_2964,N_29943,N_29992);
xnor UO_2965 (O_2965,N_29817,N_29941);
and UO_2966 (O_2966,N_29969,N_29826);
and UO_2967 (O_2967,N_29797,N_29892);
nand UO_2968 (O_2968,N_29889,N_29995);
or UO_2969 (O_2969,N_29909,N_29704);
or UO_2970 (O_2970,N_29830,N_29918);
and UO_2971 (O_2971,N_29791,N_29953);
or UO_2972 (O_2972,N_29795,N_29823);
and UO_2973 (O_2973,N_29886,N_29725);
nor UO_2974 (O_2974,N_29700,N_29745);
nand UO_2975 (O_2975,N_29770,N_29800);
or UO_2976 (O_2976,N_29925,N_29714);
and UO_2977 (O_2977,N_29732,N_29844);
or UO_2978 (O_2978,N_29972,N_29851);
or UO_2979 (O_2979,N_29890,N_29980);
and UO_2980 (O_2980,N_29742,N_29997);
and UO_2981 (O_2981,N_29703,N_29953);
nor UO_2982 (O_2982,N_29779,N_29967);
or UO_2983 (O_2983,N_29778,N_29908);
and UO_2984 (O_2984,N_29928,N_29732);
nand UO_2985 (O_2985,N_29929,N_29869);
nor UO_2986 (O_2986,N_29804,N_29734);
or UO_2987 (O_2987,N_29840,N_29721);
nand UO_2988 (O_2988,N_29979,N_29922);
and UO_2989 (O_2989,N_29998,N_29895);
and UO_2990 (O_2990,N_29809,N_29725);
and UO_2991 (O_2991,N_29840,N_29901);
nand UO_2992 (O_2992,N_29985,N_29836);
and UO_2993 (O_2993,N_29889,N_29900);
and UO_2994 (O_2994,N_29890,N_29825);
xor UO_2995 (O_2995,N_29723,N_29746);
xor UO_2996 (O_2996,N_29953,N_29700);
nand UO_2997 (O_2997,N_29812,N_29785);
nor UO_2998 (O_2998,N_29754,N_29953);
and UO_2999 (O_2999,N_29935,N_29859);
nor UO_3000 (O_3000,N_29875,N_29980);
nand UO_3001 (O_3001,N_29911,N_29704);
nand UO_3002 (O_3002,N_29714,N_29828);
nor UO_3003 (O_3003,N_29758,N_29862);
nor UO_3004 (O_3004,N_29987,N_29792);
nand UO_3005 (O_3005,N_29910,N_29915);
and UO_3006 (O_3006,N_29977,N_29993);
and UO_3007 (O_3007,N_29815,N_29835);
or UO_3008 (O_3008,N_29896,N_29757);
or UO_3009 (O_3009,N_29951,N_29790);
and UO_3010 (O_3010,N_29815,N_29830);
nand UO_3011 (O_3011,N_29756,N_29770);
xnor UO_3012 (O_3012,N_29951,N_29816);
and UO_3013 (O_3013,N_29848,N_29939);
nand UO_3014 (O_3014,N_29820,N_29829);
xor UO_3015 (O_3015,N_29988,N_29700);
nand UO_3016 (O_3016,N_29856,N_29711);
nand UO_3017 (O_3017,N_29841,N_29814);
or UO_3018 (O_3018,N_29998,N_29817);
or UO_3019 (O_3019,N_29777,N_29803);
nor UO_3020 (O_3020,N_29742,N_29998);
nand UO_3021 (O_3021,N_29841,N_29803);
nor UO_3022 (O_3022,N_29957,N_29843);
xor UO_3023 (O_3023,N_29945,N_29993);
nand UO_3024 (O_3024,N_29856,N_29889);
nor UO_3025 (O_3025,N_29859,N_29879);
nor UO_3026 (O_3026,N_29854,N_29986);
xnor UO_3027 (O_3027,N_29834,N_29751);
nand UO_3028 (O_3028,N_29791,N_29990);
nor UO_3029 (O_3029,N_29749,N_29736);
and UO_3030 (O_3030,N_29907,N_29702);
or UO_3031 (O_3031,N_29740,N_29941);
nand UO_3032 (O_3032,N_29715,N_29849);
nor UO_3033 (O_3033,N_29970,N_29954);
xor UO_3034 (O_3034,N_29703,N_29789);
or UO_3035 (O_3035,N_29855,N_29706);
xor UO_3036 (O_3036,N_29703,N_29748);
or UO_3037 (O_3037,N_29972,N_29797);
nand UO_3038 (O_3038,N_29968,N_29945);
nand UO_3039 (O_3039,N_29996,N_29769);
and UO_3040 (O_3040,N_29836,N_29842);
nand UO_3041 (O_3041,N_29847,N_29799);
nand UO_3042 (O_3042,N_29904,N_29986);
nor UO_3043 (O_3043,N_29941,N_29912);
nand UO_3044 (O_3044,N_29863,N_29995);
nor UO_3045 (O_3045,N_29770,N_29781);
nand UO_3046 (O_3046,N_29705,N_29943);
or UO_3047 (O_3047,N_29729,N_29838);
or UO_3048 (O_3048,N_29798,N_29826);
nand UO_3049 (O_3049,N_29810,N_29952);
and UO_3050 (O_3050,N_29760,N_29936);
or UO_3051 (O_3051,N_29923,N_29869);
nand UO_3052 (O_3052,N_29915,N_29919);
and UO_3053 (O_3053,N_29985,N_29749);
or UO_3054 (O_3054,N_29975,N_29782);
or UO_3055 (O_3055,N_29920,N_29895);
xor UO_3056 (O_3056,N_29985,N_29739);
or UO_3057 (O_3057,N_29806,N_29752);
and UO_3058 (O_3058,N_29701,N_29914);
nor UO_3059 (O_3059,N_29946,N_29701);
xnor UO_3060 (O_3060,N_29957,N_29993);
nand UO_3061 (O_3061,N_29961,N_29988);
and UO_3062 (O_3062,N_29763,N_29813);
or UO_3063 (O_3063,N_29877,N_29711);
and UO_3064 (O_3064,N_29739,N_29885);
nor UO_3065 (O_3065,N_29815,N_29725);
and UO_3066 (O_3066,N_29908,N_29700);
nand UO_3067 (O_3067,N_29802,N_29762);
or UO_3068 (O_3068,N_29925,N_29858);
nand UO_3069 (O_3069,N_29715,N_29978);
xnor UO_3070 (O_3070,N_29741,N_29777);
xor UO_3071 (O_3071,N_29761,N_29726);
xnor UO_3072 (O_3072,N_29971,N_29702);
or UO_3073 (O_3073,N_29891,N_29952);
nand UO_3074 (O_3074,N_29965,N_29909);
or UO_3075 (O_3075,N_29903,N_29761);
nor UO_3076 (O_3076,N_29890,N_29908);
or UO_3077 (O_3077,N_29755,N_29756);
xor UO_3078 (O_3078,N_29832,N_29701);
and UO_3079 (O_3079,N_29792,N_29994);
xnor UO_3080 (O_3080,N_29919,N_29968);
and UO_3081 (O_3081,N_29769,N_29730);
or UO_3082 (O_3082,N_29988,N_29915);
and UO_3083 (O_3083,N_29738,N_29708);
or UO_3084 (O_3084,N_29994,N_29843);
nand UO_3085 (O_3085,N_29857,N_29707);
xor UO_3086 (O_3086,N_29850,N_29858);
nand UO_3087 (O_3087,N_29767,N_29739);
and UO_3088 (O_3088,N_29717,N_29905);
nor UO_3089 (O_3089,N_29833,N_29960);
xor UO_3090 (O_3090,N_29943,N_29798);
nor UO_3091 (O_3091,N_29822,N_29968);
and UO_3092 (O_3092,N_29987,N_29875);
and UO_3093 (O_3093,N_29731,N_29777);
nor UO_3094 (O_3094,N_29764,N_29884);
or UO_3095 (O_3095,N_29916,N_29746);
xnor UO_3096 (O_3096,N_29825,N_29859);
or UO_3097 (O_3097,N_29969,N_29773);
nand UO_3098 (O_3098,N_29972,N_29914);
and UO_3099 (O_3099,N_29836,N_29703);
or UO_3100 (O_3100,N_29744,N_29947);
and UO_3101 (O_3101,N_29825,N_29931);
xor UO_3102 (O_3102,N_29984,N_29916);
nor UO_3103 (O_3103,N_29781,N_29964);
xor UO_3104 (O_3104,N_29783,N_29863);
nand UO_3105 (O_3105,N_29787,N_29705);
xnor UO_3106 (O_3106,N_29805,N_29858);
xnor UO_3107 (O_3107,N_29700,N_29884);
nand UO_3108 (O_3108,N_29900,N_29951);
xnor UO_3109 (O_3109,N_29897,N_29785);
and UO_3110 (O_3110,N_29832,N_29952);
xor UO_3111 (O_3111,N_29958,N_29894);
nand UO_3112 (O_3112,N_29823,N_29940);
xor UO_3113 (O_3113,N_29916,N_29833);
nor UO_3114 (O_3114,N_29997,N_29875);
and UO_3115 (O_3115,N_29735,N_29943);
xnor UO_3116 (O_3116,N_29823,N_29966);
and UO_3117 (O_3117,N_29979,N_29970);
nand UO_3118 (O_3118,N_29783,N_29965);
and UO_3119 (O_3119,N_29811,N_29938);
xnor UO_3120 (O_3120,N_29826,N_29895);
xnor UO_3121 (O_3121,N_29773,N_29784);
nor UO_3122 (O_3122,N_29993,N_29739);
nand UO_3123 (O_3123,N_29866,N_29875);
and UO_3124 (O_3124,N_29749,N_29784);
nand UO_3125 (O_3125,N_29784,N_29804);
nor UO_3126 (O_3126,N_29700,N_29768);
nand UO_3127 (O_3127,N_29975,N_29873);
and UO_3128 (O_3128,N_29855,N_29864);
and UO_3129 (O_3129,N_29765,N_29761);
xor UO_3130 (O_3130,N_29877,N_29817);
xor UO_3131 (O_3131,N_29737,N_29857);
and UO_3132 (O_3132,N_29921,N_29847);
or UO_3133 (O_3133,N_29917,N_29725);
or UO_3134 (O_3134,N_29745,N_29802);
nand UO_3135 (O_3135,N_29871,N_29724);
nand UO_3136 (O_3136,N_29932,N_29811);
or UO_3137 (O_3137,N_29923,N_29811);
or UO_3138 (O_3138,N_29913,N_29810);
and UO_3139 (O_3139,N_29740,N_29725);
xnor UO_3140 (O_3140,N_29931,N_29774);
nand UO_3141 (O_3141,N_29746,N_29733);
xnor UO_3142 (O_3142,N_29974,N_29794);
nand UO_3143 (O_3143,N_29912,N_29871);
and UO_3144 (O_3144,N_29719,N_29765);
and UO_3145 (O_3145,N_29922,N_29821);
and UO_3146 (O_3146,N_29730,N_29747);
and UO_3147 (O_3147,N_29784,N_29799);
or UO_3148 (O_3148,N_29772,N_29781);
or UO_3149 (O_3149,N_29937,N_29975);
or UO_3150 (O_3150,N_29767,N_29943);
and UO_3151 (O_3151,N_29883,N_29875);
or UO_3152 (O_3152,N_29869,N_29703);
nor UO_3153 (O_3153,N_29992,N_29766);
xnor UO_3154 (O_3154,N_29902,N_29774);
nand UO_3155 (O_3155,N_29876,N_29956);
xnor UO_3156 (O_3156,N_29932,N_29954);
nand UO_3157 (O_3157,N_29928,N_29794);
nor UO_3158 (O_3158,N_29935,N_29986);
and UO_3159 (O_3159,N_29750,N_29768);
nand UO_3160 (O_3160,N_29868,N_29945);
nor UO_3161 (O_3161,N_29919,N_29788);
xor UO_3162 (O_3162,N_29858,N_29792);
or UO_3163 (O_3163,N_29803,N_29879);
xnor UO_3164 (O_3164,N_29807,N_29819);
nand UO_3165 (O_3165,N_29945,N_29838);
or UO_3166 (O_3166,N_29757,N_29811);
nor UO_3167 (O_3167,N_29894,N_29920);
or UO_3168 (O_3168,N_29998,N_29905);
nor UO_3169 (O_3169,N_29826,N_29970);
xor UO_3170 (O_3170,N_29921,N_29889);
xor UO_3171 (O_3171,N_29868,N_29830);
or UO_3172 (O_3172,N_29774,N_29932);
xnor UO_3173 (O_3173,N_29776,N_29705);
nand UO_3174 (O_3174,N_29767,N_29972);
nand UO_3175 (O_3175,N_29899,N_29917);
and UO_3176 (O_3176,N_29739,N_29814);
and UO_3177 (O_3177,N_29925,N_29713);
or UO_3178 (O_3178,N_29876,N_29927);
nor UO_3179 (O_3179,N_29801,N_29916);
nor UO_3180 (O_3180,N_29922,N_29848);
or UO_3181 (O_3181,N_29914,N_29870);
nand UO_3182 (O_3182,N_29886,N_29944);
xor UO_3183 (O_3183,N_29927,N_29851);
xnor UO_3184 (O_3184,N_29978,N_29983);
nor UO_3185 (O_3185,N_29920,N_29951);
nor UO_3186 (O_3186,N_29960,N_29722);
and UO_3187 (O_3187,N_29757,N_29803);
nor UO_3188 (O_3188,N_29755,N_29819);
xor UO_3189 (O_3189,N_29784,N_29865);
nand UO_3190 (O_3190,N_29971,N_29706);
nand UO_3191 (O_3191,N_29983,N_29756);
xnor UO_3192 (O_3192,N_29778,N_29745);
nand UO_3193 (O_3193,N_29735,N_29807);
or UO_3194 (O_3194,N_29930,N_29866);
nand UO_3195 (O_3195,N_29815,N_29977);
xnor UO_3196 (O_3196,N_29969,N_29783);
nor UO_3197 (O_3197,N_29920,N_29859);
and UO_3198 (O_3198,N_29705,N_29718);
or UO_3199 (O_3199,N_29721,N_29880);
or UO_3200 (O_3200,N_29816,N_29978);
or UO_3201 (O_3201,N_29781,N_29905);
or UO_3202 (O_3202,N_29948,N_29728);
and UO_3203 (O_3203,N_29952,N_29990);
and UO_3204 (O_3204,N_29930,N_29925);
and UO_3205 (O_3205,N_29769,N_29775);
or UO_3206 (O_3206,N_29757,N_29785);
or UO_3207 (O_3207,N_29814,N_29756);
and UO_3208 (O_3208,N_29991,N_29914);
and UO_3209 (O_3209,N_29826,N_29890);
and UO_3210 (O_3210,N_29937,N_29815);
nand UO_3211 (O_3211,N_29776,N_29728);
xnor UO_3212 (O_3212,N_29973,N_29904);
nand UO_3213 (O_3213,N_29839,N_29900);
xor UO_3214 (O_3214,N_29709,N_29819);
nand UO_3215 (O_3215,N_29744,N_29844);
xor UO_3216 (O_3216,N_29795,N_29766);
xor UO_3217 (O_3217,N_29939,N_29985);
xnor UO_3218 (O_3218,N_29964,N_29819);
and UO_3219 (O_3219,N_29705,N_29914);
xnor UO_3220 (O_3220,N_29919,N_29964);
nor UO_3221 (O_3221,N_29826,N_29844);
xor UO_3222 (O_3222,N_29753,N_29933);
nor UO_3223 (O_3223,N_29721,N_29736);
nand UO_3224 (O_3224,N_29873,N_29810);
or UO_3225 (O_3225,N_29832,N_29943);
and UO_3226 (O_3226,N_29867,N_29989);
and UO_3227 (O_3227,N_29884,N_29923);
and UO_3228 (O_3228,N_29945,N_29708);
nor UO_3229 (O_3229,N_29873,N_29832);
and UO_3230 (O_3230,N_29756,N_29945);
xnor UO_3231 (O_3231,N_29791,N_29833);
and UO_3232 (O_3232,N_29705,N_29904);
nor UO_3233 (O_3233,N_29880,N_29858);
nand UO_3234 (O_3234,N_29856,N_29731);
and UO_3235 (O_3235,N_29915,N_29807);
xnor UO_3236 (O_3236,N_29709,N_29789);
or UO_3237 (O_3237,N_29822,N_29939);
and UO_3238 (O_3238,N_29873,N_29939);
or UO_3239 (O_3239,N_29922,N_29889);
nor UO_3240 (O_3240,N_29903,N_29988);
or UO_3241 (O_3241,N_29808,N_29723);
nand UO_3242 (O_3242,N_29808,N_29925);
or UO_3243 (O_3243,N_29831,N_29768);
xor UO_3244 (O_3244,N_29928,N_29917);
and UO_3245 (O_3245,N_29935,N_29903);
and UO_3246 (O_3246,N_29814,N_29807);
or UO_3247 (O_3247,N_29907,N_29792);
or UO_3248 (O_3248,N_29851,N_29873);
and UO_3249 (O_3249,N_29906,N_29987);
or UO_3250 (O_3250,N_29787,N_29897);
xor UO_3251 (O_3251,N_29980,N_29895);
nand UO_3252 (O_3252,N_29789,N_29736);
nand UO_3253 (O_3253,N_29714,N_29974);
and UO_3254 (O_3254,N_29830,N_29993);
nor UO_3255 (O_3255,N_29862,N_29898);
or UO_3256 (O_3256,N_29857,N_29808);
or UO_3257 (O_3257,N_29738,N_29962);
or UO_3258 (O_3258,N_29972,N_29745);
nor UO_3259 (O_3259,N_29798,N_29789);
nor UO_3260 (O_3260,N_29731,N_29926);
nor UO_3261 (O_3261,N_29923,N_29875);
nand UO_3262 (O_3262,N_29863,N_29752);
or UO_3263 (O_3263,N_29729,N_29795);
and UO_3264 (O_3264,N_29786,N_29856);
and UO_3265 (O_3265,N_29743,N_29900);
xor UO_3266 (O_3266,N_29705,N_29700);
xor UO_3267 (O_3267,N_29883,N_29780);
nand UO_3268 (O_3268,N_29819,N_29916);
nor UO_3269 (O_3269,N_29806,N_29749);
xnor UO_3270 (O_3270,N_29946,N_29992);
nand UO_3271 (O_3271,N_29706,N_29858);
nor UO_3272 (O_3272,N_29769,N_29856);
and UO_3273 (O_3273,N_29990,N_29747);
nand UO_3274 (O_3274,N_29903,N_29720);
nand UO_3275 (O_3275,N_29932,N_29738);
and UO_3276 (O_3276,N_29909,N_29739);
and UO_3277 (O_3277,N_29826,N_29705);
and UO_3278 (O_3278,N_29828,N_29938);
xor UO_3279 (O_3279,N_29739,N_29898);
or UO_3280 (O_3280,N_29744,N_29732);
or UO_3281 (O_3281,N_29798,N_29843);
nand UO_3282 (O_3282,N_29881,N_29992);
nor UO_3283 (O_3283,N_29735,N_29837);
nand UO_3284 (O_3284,N_29787,N_29895);
nor UO_3285 (O_3285,N_29993,N_29839);
nor UO_3286 (O_3286,N_29778,N_29748);
nand UO_3287 (O_3287,N_29897,N_29792);
nand UO_3288 (O_3288,N_29857,N_29863);
and UO_3289 (O_3289,N_29836,N_29915);
and UO_3290 (O_3290,N_29701,N_29853);
or UO_3291 (O_3291,N_29981,N_29942);
nor UO_3292 (O_3292,N_29846,N_29816);
nand UO_3293 (O_3293,N_29837,N_29748);
nand UO_3294 (O_3294,N_29747,N_29842);
or UO_3295 (O_3295,N_29786,N_29768);
nor UO_3296 (O_3296,N_29886,N_29781);
and UO_3297 (O_3297,N_29933,N_29785);
and UO_3298 (O_3298,N_29866,N_29792);
nor UO_3299 (O_3299,N_29797,N_29754);
nand UO_3300 (O_3300,N_29862,N_29973);
or UO_3301 (O_3301,N_29795,N_29980);
or UO_3302 (O_3302,N_29766,N_29706);
xnor UO_3303 (O_3303,N_29741,N_29742);
or UO_3304 (O_3304,N_29899,N_29726);
or UO_3305 (O_3305,N_29873,N_29995);
and UO_3306 (O_3306,N_29962,N_29972);
or UO_3307 (O_3307,N_29842,N_29934);
xor UO_3308 (O_3308,N_29778,N_29721);
and UO_3309 (O_3309,N_29793,N_29940);
nand UO_3310 (O_3310,N_29701,N_29758);
and UO_3311 (O_3311,N_29828,N_29791);
or UO_3312 (O_3312,N_29708,N_29775);
or UO_3313 (O_3313,N_29805,N_29898);
nand UO_3314 (O_3314,N_29847,N_29956);
or UO_3315 (O_3315,N_29802,N_29845);
xor UO_3316 (O_3316,N_29806,N_29916);
xnor UO_3317 (O_3317,N_29882,N_29864);
and UO_3318 (O_3318,N_29981,N_29960);
xnor UO_3319 (O_3319,N_29817,N_29899);
nor UO_3320 (O_3320,N_29821,N_29839);
nor UO_3321 (O_3321,N_29820,N_29981);
xor UO_3322 (O_3322,N_29947,N_29869);
and UO_3323 (O_3323,N_29913,N_29720);
xnor UO_3324 (O_3324,N_29819,N_29951);
nor UO_3325 (O_3325,N_29892,N_29724);
xor UO_3326 (O_3326,N_29950,N_29752);
or UO_3327 (O_3327,N_29988,N_29853);
xnor UO_3328 (O_3328,N_29932,N_29794);
and UO_3329 (O_3329,N_29898,N_29948);
xor UO_3330 (O_3330,N_29871,N_29707);
nor UO_3331 (O_3331,N_29830,N_29935);
and UO_3332 (O_3332,N_29763,N_29807);
xor UO_3333 (O_3333,N_29773,N_29968);
xnor UO_3334 (O_3334,N_29763,N_29930);
nand UO_3335 (O_3335,N_29858,N_29833);
xnor UO_3336 (O_3336,N_29903,N_29994);
or UO_3337 (O_3337,N_29847,N_29842);
nand UO_3338 (O_3338,N_29783,N_29782);
nand UO_3339 (O_3339,N_29999,N_29793);
or UO_3340 (O_3340,N_29998,N_29956);
nor UO_3341 (O_3341,N_29727,N_29966);
nor UO_3342 (O_3342,N_29800,N_29844);
or UO_3343 (O_3343,N_29947,N_29793);
nand UO_3344 (O_3344,N_29894,N_29716);
and UO_3345 (O_3345,N_29881,N_29916);
or UO_3346 (O_3346,N_29897,N_29703);
and UO_3347 (O_3347,N_29817,N_29768);
nand UO_3348 (O_3348,N_29947,N_29997);
and UO_3349 (O_3349,N_29841,N_29850);
nand UO_3350 (O_3350,N_29779,N_29777);
or UO_3351 (O_3351,N_29801,N_29832);
and UO_3352 (O_3352,N_29750,N_29841);
nor UO_3353 (O_3353,N_29828,N_29810);
nor UO_3354 (O_3354,N_29832,N_29824);
nor UO_3355 (O_3355,N_29840,N_29976);
nor UO_3356 (O_3356,N_29874,N_29805);
nand UO_3357 (O_3357,N_29914,N_29801);
nor UO_3358 (O_3358,N_29865,N_29944);
or UO_3359 (O_3359,N_29980,N_29859);
xor UO_3360 (O_3360,N_29940,N_29767);
and UO_3361 (O_3361,N_29712,N_29825);
nor UO_3362 (O_3362,N_29886,N_29782);
and UO_3363 (O_3363,N_29707,N_29891);
nand UO_3364 (O_3364,N_29956,N_29952);
nor UO_3365 (O_3365,N_29798,N_29860);
and UO_3366 (O_3366,N_29708,N_29781);
nor UO_3367 (O_3367,N_29992,N_29962);
or UO_3368 (O_3368,N_29992,N_29923);
nand UO_3369 (O_3369,N_29802,N_29999);
and UO_3370 (O_3370,N_29954,N_29983);
xor UO_3371 (O_3371,N_29956,N_29990);
nand UO_3372 (O_3372,N_29927,N_29706);
and UO_3373 (O_3373,N_29910,N_29949);
and UO_3374 (O_3374,N_29838,N_29860);
xor UO_3375 (O_3375,N_29960,N_29808);
and UO_3376 (O_3376,N_29843,N_29840);
nand UO_3377 (O_3377,N_29860,N_29929);
or UO_3378 (O_3378,N_29807,N_29849);
nand UO_3379 (O_3379,N_29796,N_29961);
xnor UO_3380 (O_3380,N_29765,N_29730);
nor UO_3381 (O_3381,N_29964,N_29922);
nand UO_3382 (O_3382,N_29934,N_29708);
nor UO_3383 (O_3383,N_29719,N_29791);
nor UO_3384 (O_3384,N_29826,N_29837);
xor UO_3385 (O_3385,N_29747,N_29757);
and UO_3386 (O_3386,N_29862,N_29950);
nor UO_3387 (O_3387,N_29884,N_29905);
nor UO_3388 (O_3388,N_29744,N_29964);
and UO_3389 (O_3389,N_29845,N_29741);
and UO_3390 (O_3390,N_29964,N_29747);
and UO_3391 (O_3391,N_29888,N_29790);
xnor UO_3392 (O_3392,N_29724,N_29981);
and UO_3393 (O_3393,N_29875,N_29814);
nor UO_3394 (O_3394,N_29793,N_29781);
nand UO_3395 (O_3395,N_29759,N_29924);
xnor UO_3396 (O_3396,N_29951,N_29868);
and UO_3397 (O_3397,N_29918,N_29976);
nand UO_3398 (O_3398,N_29999,N_29756);
and UO_3399 (O_3399,N_29949,N_29762);
nor UO_3400 (O_3400,N_29846,N_29994);
xor UO_3401 (O_3401,N_29707,N_29949);
and UO_3402 (O_3402,N_29850,N_29921);
nor UO_3403 (O_3403,N_29851,N_29936);
or UO_3404 (O_3404,N_29920,N_29903);
or UO_3405 (O_3405,N_29905,N_29803);
and UO_3406 (O_3406,N_29900,N_29972);
nor UO_3407 (O_3407,N_29714,N_29905);
and UO_3408 (O_3408,N_29792,N_29751);
nand UO_3409 (O_3409,N_29865,N_29743);
nor UO_3410 (O_3410,N_29779,N_29945);
or UO_3411 (O_3411,N_29705,N_29942);
or UO_3412 (O_3412,N_29838,N_29907);
xnor UO_3413 (O_3413,N_29700,N_29821);
nor UO_3414 (O_3414,N_29980,N_29888);
xnor UO_3415 (O_3415,N_29956,N_29794);
or UO_3416 (O_3416,N_29819,N_29928);
or UO_3417 (O_3417,N_29967,N_29753);
nand UO_3418 (O_3418,N_29803,N_29926);
xnor UO_3419 (O_3419,N_29928,N_29884);
nand UO_3420 (O_3420,N_29709,N_29930);
nor UO_3421 (O_3421,N_29787,N_29717);
xnor UO_3422 (O_3422,N_29938,N_29987);
and UO_3423 (O_3423,N_29704,N_29735);
and UO_3424 (O_3424,N_29904,N_29947);
nor UO_3425 (O_3425,N_29984,N_29798);
nand UO_3426 (O_3426,N_29741,N_29772);
or UO_3427 (O_3427,N_29809,N_29821);
or UO_3428 (O_3428,N_29958,N_29910);
and UO_3429 (O_3429,N_29752,N_29746);
or UO_3430 (O_3430,N_29827,N_29795);
and UO_3431 (O_3431,N_29981,N_29994);
xnor UO_3432 (O_3432,N_29794,N_29813);
and UO_3433 (O_3433,N_29968,N_29879);
xnor UO_3434 (O_3434,N_29967,N_29733);
xnor UO_3435 (O_3435,N_29828,N_29761);
nand UO_3436 (O_3436,N_29701,N_29937);
nand UO_3437 (O_3437,N_29795,N_29983);
xor UO_3438 (O_3438,N_29796,N_29824);
and UO_3439 (O_3439,N_29787,N_29730);
nand UO_3440 (O_3440,N_29752,N_29716);
and UO_3441 (O_3441,N_29906,N_29846);
and UO_3442 (O_3442,N_29945,N_29943);
or UO_3443 (O_3443,N_29862,N_29864);
and UO_3444 (O_3444,N_29970,N_29947);
or UO_3445 (O_3445,N_29728,N_29755);
nor UO_3446 (O_3446,N_29746,N_29785);
xor UO_3447 (O_3447,N_29962,N_29863);
xor UO_3448 (O_3448,N_29844,N_29778);
and UO_3449 (O_3449,N_29733,N_29729);
nor UO_3450 (O_3450,N_29757,N_29832);
nor UO_3451 (O_3451,N_29932,N_29863);
xor UO_3452 (O_3452,N_29813,N_29748);
nand UO_3453 (O_3453,N_29905,N_29733);
or UO_3454 (O_3454,N_29825,N_29921);
nor UO_3455 (O_3455,N_29725,N_29982);
xor UO_3456 (O_3456,N_29830,N_29734);
or UO_3457 (O_3457,N_29918,N_29786);
xor UO_3458 (O_3458,N_29941,N_29793);
xnor UO_3459 (O_3459,N_29887,N_29875);
and UO_3460 (O_3460,N_29966,N_29958);
nor UO_3461 (O_3461,N_29988,N_29891);
nor UO_3462 (O_3462,N_29798,N_29948);
xnor UO_3463 (O_3463,N_29830,N_29945);
nand UO_3464 (O_3464,N_29985,N_29969);
or UO_3465 (O_3465,N_29897,N_29991);
xor UO_3466 (O_3466,N_29715,N_29806);
or UO_3467 (O_3467,N_29939,N_29784);
xnor UO_3468 (O_3468,N_29949,N_29924);
or UO_3469 (O_3469,N_29817,N_29923);
or UO_3470 (O_3470,N_29872,N_29993);
nand UO_3471 (O_3471,N_29720,N_29879);
nand UO_3472 (O_3472,N_29996,N_29878);
nand UO_3473 (O_3473,N_29912,N_29812);
nand UO_3474 (O_3474,N_29790,N_29808);
xor UO_3475 (O_3475,N_29731,N_29774);
xnor UO_3476 (O_3476,N_29764,N_29756);
and UO_3477 (O_3477,N_29728,N_29786);
or UO_3478 (O_3478,N_29986,N_29956);
xnor UO_3479 (O_3479,N_29914,N_29904);
xor UO_3480 (O_3480,N_29964,N_29791);
xor UO_3481 (O_3481,N_29795,N_29805);
or UO_3482 (O_3482,N_29704,N_29801);
nand UO_3483 (O_3483,N_29899,N_29892);
xor UO_3484 (O_3484,N_29909,N_29731);
and UO_3485 (O_3485,N_29711,N_29958);
nor UO_3486 (O_3486,N_29750,N_29868);
nand UO_3487 (O_3487,N_29940,N_29736);
or UO_3488 (O_3488,N_29758,N_29750);
nand UO_3489 (O_3489,N_29845,N_29890);
nand UO_3490 (O_3490,N_29915,N_29884);
and UO_3491 (O_3491,N_29862,N_29737);
nand UO_3492 (O_3492,N_29785,N_29942);
xor UO_3493 (O_3493,N_29729,N_29707);
or UO_3494 (O_3494,N_29700,N_29900);
and UO_3495 (O_3495,N_29750,N_29723);
nand UO_3496 (O_3496,N_29834,N_29837);
or UO_3497 (O_3497,N_29956,N_29742);
nand UO_3498 (O_3498,N_29931,N_29823);
nor UO_3499 (O_3499,N_29825,N_29913);
endmodule