module basic_5000_50000_5000_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_1878,In_3667);
or U1 (N_1,In_1849,In_2771);
nor U2 (N_2,In_4304,In_2755);
xor U3 (N_3,In_587,In_1828);
or U4 (N_4,In_1498,In_1099);
nand U5 (N_5,In_2608,In_1385);
nand U6 (N_6,In_1596,In_2480);
nand U7 (N_7,In_228,In_4837);
and U8 (N_8,In_2019,In_2494);
xor U9 (N_9,In_681,In_1838);
and U10 (N_10,In_875,In_2651);
and U11 (N_11,In_2601,In_4801);
nor U12 (N_12,In_4977,In_1757);
nand U13 (N_13,In_3375,In_3705);
nand U14 (N_14,In_1217,In_3245);
and U15 (N_15,In_3811,In_3880);
nand U16 (N_16,In_2655,In_2818);
nor U17 (N_17,In_840,In_4385);
and U18 (N_18,In_2979,In_4283);
and U19 (N_19,In_4622,In_4880);
or U20 (N_20,In_77,In_816);
or U21 (N_21,In_4399,In_2069);
nand U22 (N_22,In_4642,In_3308);
and U23 (N_23,In_2567,In_1968);
or U24 (N_24,In_2799,In_3043);
xnor U25 (N_25,In_1910,In_1004);
and U26 (N_26,In_1130,In_219);
nor U27 (N_27,In_1325,In_3801);
xnor U28 (N_28,In_1037,In_3474);
nand U29 (N_29,In_289,In_2718);
or U30 (N_30,In_4634,In_2883);
and U31 (N_31,In_2556,In_3925);
or U32 (N_32,In_4697,In_2203);
and U33 (N_33,In_99,In_567);
nand U34 (N_34,In_1943,In_276);
xnor U35 (N_35,In_4962,In_2274);
nand U36 (N_36,In_4007,In_4965);
nor U37 (N_37,In_1327,In_286);
xnor U38 (N_38,In_2352,In_1495);
or U39 (N_39,In_4479,In_621);
or U40 (N_40,In_3789,In_2198);
nor U41 (N_41,In_3357,In_995);
or U42 (N_42,In_3143,In_373);
xor U43 (N_43,In_796,In_4332);
and U44 (N_44,In_4469,In_2275);
nand U45 (N_45,In_3414,In_3389);
xor U46 (N_46,In_2028,In_1461);
nand U47 (N_47,In_4955,In_882);
nand U48 (N_48,In_196,In_476);
xnor U49 (N_49,In_1155,In_2781);
nor U50 (N_50,In_3084,In_2967);
nor U51 (N_51,In_1803,In_3348);
and U52 (N_52,In_3196,In_4257);
nor U53 (N_53,In_2416,In_3118);
nor U54 (N_54,In_3525,In_4519);
nand U55 (N_55,In_1510,In_1659);
nand U56 (N_56,In_2642,In_2266);
or U57 (N_57,In_4898,In_3826);
nor U58 (N_58,In_1378,In_2331);
and U59 (N_59,In_4023,In_4848);
nor U60 (N_60,In_1096,In_4030);
and U61 (N_61,In_1295,In_160);
nor U62 (N_62,In_392,In_605);
nor U63 (N_63,In_2242,In_3640);
nor U64 (N_64,In_1359,In_1913);
nor U65 (N_65,In_4849,In_4989);
or U66 (N_66,In_1916,In_4777);
xnor U67 (N_67,In_3516,In_3066);
xnor U68 (N_68,In_3695,In_2269);
and U69 (N_69,In_1529,In_4814);
and U70 (N_70,In_1591,In_4281);
nand U71 (N_71,In_3148,In_830);
nor U72 (N_72,In_2904,In_2670);
nand U73 (N_73,In_246,In_2102);
xnor U74 (N_74,In_439,In_3601);
nor U75 (N_75,In_907,In_3162);
xor U76 (N_76,In_3096,In_3339);
nand U77 (N_77,In_1297,In_4466);
or U78 (N_78,In_1886,In_3736);
or U79 (N_79,In_4176,In_258);
xor U80 (N_80,In_2957,In_2168);
and U81 (N_81,In_4610,In_4957);
nand U82 (N_82,In_2522,In_4318);
or U83 (N_83,In_4127,In_179);
nor U84 (N_84,In_1314,In_856);
and U85 (N_85,In_1984,In_2424);
nor U86 (N_86,In_4653,In_1507);
or U87 (N_87,In_1613,In_2592);
xnor U88 (N_88,In_1225,In_2074);
or U89 (N_89,In_4278,In_1435);
xor U90 (N_90,In_1407,In_2199);
and U91 (N_91,In_3488,In_1856);
and U92 (N_92,In_4891,In_4431);
xnor U93 (N_93,In_3007,In_1186);
nor U94 (N_94,In_2508,In_3663);
xnor U95 (N_95,In_1470,In_2138);
and U96 (N_96,In_2065,In_2495);
or U97 (N_97,In_2305,In_2082);
and U98 (N_98,In_2417,In_2772);
xor U99 (N_99,In_3476,In_4755);
nor U100 (N_100,In_2941,In_3427);
and U101 (N_101,In_4081,In_287);
and U102 (N_102,In_4565,In_44);
nand U103 (N_103,In_1287,In_1253);
nor U104 (N_104,In_530,In_1997);
xor U105 (N_105,In_154,In_661);
xnor U106 (N_106,In_4163,In_4548);
or U107 (N_107,In_1112,In_1722);
nand U108 (N_108,In_2693,In_4295);
nand U109 (N_109,In_1940,In_515);
or U110 (N_110,In_2440,In_3662);
and U111 (N_111,In_3964,In_2989);
and U112 (N_112,In_1201,In_3278);
xor U113 (N_113,In_2031,In_2895);
nand U114 (N_114,In_788,In_2842);
xnor U115 (N_115,In_2722,In_2034);
or U116 (N_116,In_2920,In_3631);
nor U117 (N_117,In_2600,In_3721);
nor U118 (N_118,In_2081,In_4672);
or U119 (N_119,In_249,In_4150);
nand U120 (N_120,In_3937,In_2506);
or U121 (N_121,In_3932,In_52);
and U122 (N_122,In_1340,In_1215);
nor U123 (N_123,In_4243,In_1169);
nand U124 (N_124,In_731,In_3412);
and U125 (N_125,In_4834,In_4794);
nand U126 (N_126,In_4074,In_2071);
nor U127 (N_127,In_4069,In_19);
or U128 (N_128,In_4252,In_1417);
nor U129 (N_129,In_3553,In_2149);
nand U130 (N_130,In_1009,In_1812);
and U131 (N_131,In_526,In_187);
xnor U132 (N_132,In_2857,In_2590);
or U133 (N_133,In_3251,In_2134);
xor U134 (N_134,In_3680,In_1714);
and U135 (N_135,In_3701,In_1232);
nor U136 (N_136,In_808,In_3696);
nand U137 (N_137,In_2917,In_1059);
xor U138 (N_138,In_1847,In_1612);
nor U139 (N_139,In_1787,In_4893);
nor U140 (N_140,In_3673,In_4836);
and U141 (N_141,In_4174,In_2067);
nand U142 (N_142,In_2903,In_3693);
or U143 (N_143,In_4482,In_520);
nand U144 (N_144,In_4047,In_4364);
nor U145 (N_145,In_3861,In_1729);
and U146 (N_146,In_541,In_400);
xnor U147 (N_147,In_775,In_2461);
nand U148 (N_148,In_3407,In_1411);
nor U149 (N_149,In_2797,In_1527);
nand U150 (N_150,In_3181,In_4013);
or U151 (N_151,In_4547,In_4494);
nand U152 (N_152,In_1116,In_4550);
nor U153 (N_153,In_1026,In_989);
and U154 (N_154,In_1924,In_3108);
nand U155 (N_155,In_1049,In_2684);
nor U156 (N_156,In_1542,In_1804);
and U157 (N_157,In_1513,In_1479);
or U158 (N_158,In_2083,In_4490);
and U159 (N_159,In_1036,In_4055);
nand U160 (N_160,In_4157,In_1746);
nor U161 (N_161,In_4630,In_4667);
or U162 (N_162,In_199,In_4656);
or U163 (N_163,In_1980,In_719);
xnor U164 (N_164,In_1947,In_545);
xnor U165 (N_165,In_3697,In_291);
nand U166 (N_166,In_416,In_387);
and U167 (N_167,In_3421,In_2481);
and U168 (N_168,In_3097,In_2535);
nor U169 (N_169,In_3018,In_1660);
or U170 (N_170,In_3253,In_2927);
xor U171 (N_171,In_3161,In_3552);
nor U172 (N_172,In_2202,In_2001);
and U173 (N_173,In_3828,In_2714);
and U174 (N_174,In_4995,In_3615);
or U175 (N_175,In_4128,In_1248);
xnor U176 (N_176,In_1742,In_4707);
xnor U177 (N_177,In_3294,In_4838);
xor U178 (N_178,In_354,In_4102);
and U179 (N_179,In_2749,In_3838);
xor U180 (N_180,In_4981,In_3408);
nor U181 (N_181,In_4476,In_4756);
nor U182 (N_182,In_3677,In_2819);
nand U183 (N_183,In_1089,In_634);
nand U184 (N_184,In_4588,In_894);
and U185 (N_185,In_4120,In_474);
and U186 (N_186,In_3060,In_1354);
nand U187 (N_187,In_2326,In_3757);
or U188 (N_188,In_3603,In_2365);
xnor U189 (N_189,In_1029,In_2958);
nor U190 (N_190,In_2251,In_1117);
nor U191 (N_191,In_4964,In_1556);
and U192 (N_192,In_3052,In_1971);
nor U193 (N_193,In_1552,In_2848);
and U194 (N_194,In_4910,In_27);
nor U195 (N_195,In_4640,In_665);
or U196 (N_196,In_2291,In_1467);
nand U197 (N_197,In_1097,In_4865);
nand U198 (N_198,In_4419,In_2725);
nand U199 (N_199,In_1324,In_2969);
xnor U200 (N_200,In_2187,In_1296);
xor U201 (N_201,In_1268,In_3495);
nor U202 (N_202,In_14,In_1921);
nand U203 (N_203,In_2690,In_4031);
nor U204 (N_204,In_4601,In_1727);
or U205 (N_205,In_3458,In_3071);
or U206 (N_206,In_3596,In_2041);
nor U207 (N_207,In_1170,In_4587);
xnor U208 (N_208,In_4813,In_4961);
nor U209 (N_209,In_247,In_4740);
xor U210 (N_210,In_4038,In_4341);
xnor U211 (N_211,In_1011,In_2555);
nand U212 (N_212,In_3630,In_643);
xnor U213 (N_213,In_57,In_1469);
xnor U214 (N_214,In_304,In_2003);
xnor U215 (N_215,In_1840,In_2058);
or U216 (N_216,In_571,In_2196);
nand U217 (N_217,In_3415,In_2699);
or U218 (N_218,In_217,In_3600);
nand U219 (N_219,In_3765,In_3208);
nor U220 (N_220,In_747,In_2817);
nor U221 (N_221,In_2175,In_3716);
and U222 (N_222,In_3742,In_4238);
nor U223 (N_223,In_2356,In_4478);
nand U224 (N_224,In_3286,In_3768);
xnor U225 (N_225,In_4311,In_4406);
xnor U226 (N_226,In_4641,In_2265);
nor U227 (N_227,In_2496,In_3247);
nor U228 (N_228,In_1264,In_1643);
and U229 (N_229,In_4573,In_1677);
nor U230 (N_230,In_3921,In_1432);
xnor U231 (N_231,In_4284,In_4182);
nor U232 (N_232,In_557,In_277);
or U233 (N_233,In_2271,In_2829);
nand U234 (N_234,In_8,In_2197);
nand U235 (N_235,In_1014,In_3902);
or U236 (N_236,In_782,In_1731);
xor U237 (N_237,In_4762,In_1740);
xnor U238 (N_238,In_3766,In_1959);
xnor U239 (N_239,In_2446,In_2195);
xor U240 (N_240,In_803,In_3349);
or U241 (N_241,In_4008,In_1717);
or U242 (N_242,In_4189,In_3436);
and U243 (N_243,In_1292,In_2816);
and U244 (N_244,In_1871,In_85);
nand U245 (N_245,In_2994,In_461);
and U246 (N_246,In_4557,In_3085);
nand U247 (N_247,In_1082,In_3026);
nor U248 (N_248,In_2936,In_1647);
and U249 (N_249,In_2382,In_2914);
and U250 (N_250,In_3409,In_74);
and U251 (N_251,In_2307,In_2243);
nor U252 (N_252,In_4978,In_426);
nand U253 (N_253,In_3632,In_384);
nand U254 (N_254,In_4061,In_3590);
nor U255 (N_255,In_432,In_3588);
nand U256 (N_256,In_3992,In_532);
and U257 (N_257,In_910,In_2836);
and U258 (N_258,In_4546,In_1023);
nor U259 (N_259,In_2475,In_2574);
nor U260 (N_260,In_3301,In_29);
or U261 (N_261,In_4106,In_702);
or U262 (N_262,In_2838,In_4649);
nand U263 (N_263,In_4843,In_838);
nor U264 (N_264,In_4844,In_4448);
nand U265 (N_265,In_2673,In_1310);
xor U266 (N_266,In_2039,In_1188);
xnor U267 (N_267,In_4138,In_3848);
nor U268 (N_268,In_4231,In_748);
and U269 (N_269,In_2701,In_4433);
nand U270 (N_270,In_807,In_2204);
nand U271 (N_271,In_2768,In_1171);
nand U272 (N_272,In_4054,In_1987);
nor U273 (N_273,In_4405,In_3190);
nor U274 (N_274,In_1543,In_519);
or U275 (N_275,In_2934,In_1339);
nand U276 (N_276,In_3452,In_477);
xor U277 (N_277,In_1930,In_4867);
or U278 (N_278,In_2521,In_608);
nand U279 (N_279,In_2993,In_1439);
nor U280 (N_280,In_877,In_3237);
xor U281 (N_281,In_1883,In_4280);
and U282 (N_282,In_1544,In_1805);
xnor U283 (N_283,In_3512,In_862);
and U284 (N_284,In_1967,In_4036);
xor U285 (N_285,In_4552,In_592);
and U286 (N_286,In_926,In_2120);
or U287 (N_287,In_4040,In_4320);
and U288 (N_288,In_2695,In_177);
or U289 (N_289,In_656,In_4168);
nand U290 (N_290,In_1960,In_4888);
nor U291 (N_291,In_3967,In_2519);
or U292 (N_292,In_4875,In_3400);
or U293 (N_293,In_2793,In_2996);
nor U294 (N_294,In_793,In_1276);
xnor U295 (N_295,In_3129,In_2944);
nand U296 (N_296,In_3907,In_1460);
and U297 (N_297,In_2933,In_261);
xnor U298 (N_298,In_4410,In_3679);
and U299 (N_299,In_535,In_1021);
nor U300 (N_300,In_2908,In_4742);
nand U301 (N_301,In_1972,In_2249);
nor U302 (N_302,In_2036,In_264);
or U303 (N_303,In_3000,In_2860);
or U304 (N_304,In_1751,In_2975);
or U305 (N_305,In_1762,In_4387);
xor U306 (N_306,In_1299,In_1394);
or U307 (N_307,In_341,In_745);
xor U308 (N_308,In_306,In_851);
and U309 (N_309,In_4868,In_3713);
xor U310 (N_310,In_4738,In_577);
nand U311 (N_311,In_904,In_1792);
and U312 (N_312,In_3947,In_4839);
nand U313 (N_313,In_2663,In_231);
nand U314 (N_314,In_2640,In_2825);
nand U315 (N_315,In_837,In_3669);
nand U316 (N_316,In_110,In_4741);
nand U317 (N_317,In_2541,In_4704);
nor U318 (N_318,In_4874,In_4415);
xnor U319 (N_319,In_978,In_42);
xnor U320 (N_320,In_2431,In_568);
xnor U321 (N_321,In_106,In_2516);
xor U322 (N_322,In_227,In_1005);
or U323 (N_323,In_3223,In_4358);
xnor U324 (N_324,In_4713,In_3371);
xor U325 (N_325,In_134,In_1111);
nand U326 (N_326,In_2486,In_4063);
nand U327 (N_327,In_2313,In_1649);
and U328 (N_328,In_3973,In_772);
xnor U329 (N_329,In_4970,In_3058);
nor U330 (N_330,In_2828,In_2612);
and U331 (N_331,In_4711,In_4663);
xor U332 (N_332,In_2561,In_1744);
nor U333 (N_333,In_1455,In_2792);
xnor U334 (N_334,In_590,In_240);
and U335 (N_335,In_3618,In_1351);
xnor U336 (N_336,In_879,In_3345);
xor U337 (N_337,In_2151,In_1842);
or U338 (N_338,In_3138,In_794);
or U339 (N_339,In_4924,In_714);
and U340 (N_340,In_3908,In_3782);
or U341 (N_341,In_3137,In_2208);
nand U342 (N_342,In_4728,In_4011);
or U343 (N_343,In_3112,In_3905);
and U344 (N_344,In_2657,In_4993);
or U345 (N_345,In_2005,In_3124);
nand U346 (N_346,In_302,In_997);
or U347 (N_347,In_630,In_1568);
nor U348 (N_348,In_3526,In_1535);
or U349 (N_349,In_774,In_1136);
or U350 (N_350,In_3086,In_3134);
xnor U351 (N_351,In_269,In_1050);
nand U352 (N_352,In_3582,In_581);
xnor U353 (N_353,In_327,In_4527);
and U354 (N_354,In_2008,In_3314);
xor U355 (N_355,In_3873,In_667);
xnor U356 (N_356,In_1286,In_3792);
nand U357 (N_357,In_1316,In_971);
nor U358 (N_358,In_644,In_1410);
or U359 (N_359,In_3323,In_4733);
nand U360 (N_360,In_3635,In_1690);
nand U361 (N_361,In_1114,In_2672);
nor U362 (N_362,In_3924,In_1379);
xnor U363 (N_363,In_144,In_4473);
nand U364 (N_364,In_1140,In_1970);
nand U365 (N_365,In_1309,In_3226);
xnor U366 (N_366,In_692,In_3886);
or U367 (N_367,In_1713,In_3222);
or U368 (N_368,In_493,In_455);
nand U369 (N_369,In_4599,In_3668);
or U370 (N_370,In_2193,In_2434);
nor U371 (N_371,In_1570,In_1476);
and U372 (N_372,In_2630,In_361);
nor U373 (N_373,In_1244,In_3579);
and U374 (N_374,In_863,In_2072);
or U375 (N_375,In_60,In_2215);
and U376 (N_376,In_4833,In_1464);
xnor U377 (N_377,In_2056,In_4354);
and U378 (N_378,In_1388,In_1912);
and U379 (N_379,In_3100,In_3778);
and U380 (N_380,In_3738,In_1598);
nor U381 (N_381,In_460,In_4229);
nand U382 (N_382,In_1433,In_1782);
nand U383 (N_383,In_3916,In_622);
xor U384 (N_384,In_4223,In_1844);
or U385 (N_385,In_3897,In_260);
nor U386 (N_386,In_3280,In_2871);
and U387 (N_387,In_4935,In_1794);
nand U388 (N_388,In_2614,In_4461);
nor U389 (N_389,In_2378,In_386);
and U390 (N_390,In_4067,In_108);
nand U391 (N_391,In_1154,In_4805);
nand U392 (N_392,In_3344,In_2066);
xor U393 (N_393,In_4621,In_3611);
or U394 (N_394,In_2984,In_572);
xor U395 (N_395,In_1166,In_4438);
nor U396 (N_396,In_509,In_4421);
xor U397 (N_397,In_3187,In_171);
or U398 (N_398,In_2604,In_751);
xnor U399 (N_399,In_4381,In_3035);
xnor U400 (N_400,In_4045,In_358);
or U401 (N_401,In_2032,In_1159);
xnor U402 (N_402,In_3426,In_3004);
xor U403 (N_403,In_4692,In_290);
or U404 (N_404,In_4840,In_1375);
nand U405 (N_405,In_4504,In_16);
and U406 (N_406,In_4949,In_165);
xnor U407 (N_407,In_3794,In_2394);
and U408 (N_408,In_917,In_3325);
xor U409 (N_409,In_4152,In_2551);
nand U410 (N_410,In_2272,In_3609);
nand U411 (N_411,In_2209,In_4617);
and U412 (N_412,In_4598,In_3377);
nor U413 (N_413,In_948,In_4361);
xor U414 (N_414,In_405,In_2846);
nand U415 (N_415,In_4224,In_1035);
xnor U416 (N_416,In_482,In_4449);
and U417 (N_417,In_2018,In_197);
nand U418 (N_418,In_1928,In_2851);
or U419 (N_419,In_1954,In_4563);
xor U420 (N_420,In_3616,In_3926);
nand U421 (N_421,In_3199,In_3013);
nand U422 (N_422,In_4474,In_4065);
and U423 (N_423,In_3728,In_2740);
and U424 (N_424,In_2518,In_3572);
xor U425 (N_425,In_3985,In_2063);
and U426 (N_426,In_857,In_3293);
and U427 (N_427,In_3062,In_4727);
nand U428 (N_428,In_4165,In_2925);
xor U429 (N_429,In_2361,In_1307);
or U430 (N_430,In_4968,In_2862);
and U431 (N_431,In_3670,In_220);
nand U432 (N_432,In_4513,In_984);
and U433 (N_433,In_1173,In_4409);
nor U434 (N_434,In_1926,In_4235);
nand U435 (N_435,In_2660,In_4091);
xor U436 (N_436,In_1989,In_3978);
and U437 (N_437,In_4453,In_2023);
and U438 (N_438,In_1092,In_4976);
and U439 (N_439,In_2977,In_4791);
xor U440 (N_440,In_4966,In_394);
xor U441 (N_441,In_4319,In_2284);
nand U442 (N_442,In_820,In_4650);
and U443 (N_443,In_484,In_2497);
and U444 (N_444,In_4933,In_376);
or U445 (N_445,In_229,In_3581);
and U446 (N_446,In_1144,In_194);
nor U447 (N_447,In_421,In_4633);
and U448 (N_448,In_2912,In_161);
or U449 (N_449,In_3087,In_67);
nand U450 (N_450,In_563,In_4618);
or U451 (N_451,In_3896,In_3246);
xnor U452 (N_452,In_3063,In_2509);
nor U453 (N_453,In_3597,In_4435);
nor U454 (N_454,In_2626,In_1353);
nor U455 (N_455,In_1666,In_4129);
nand U456 (N_456,In_2968,In_653);
xor U457 (N_457,In_2691,In_1839);
or U458 (N_458,In_3959,In_2805);
xnor U459 (N_459,In_2552,In_2295);
or U460 (N_460,In_312,In_2387);
nand U461 (N_461,In_3987,In_4259);
xor U462 (N_462,In_3403,In_1637);
nor U463 (N_463,In_3473,In_888);
and U464 (N_464,In_3858,In_3069);
and U465 (N_465,In_2955,In_897);
nand U466 (N_466,In_2739,In_1703);
and U467 (N_467,In_2164,In_3444);
or U468 (N_468,In_4746,In_4032);
xor U469 (N_469,In_1621,In_2629);
nor U470 (N_470,In_424,In_4930);
and U471 (N_471,In_4105,In_4486);
and U472 (N_472,In_1860,In_4472);
nor U473 (N_473,In_1755,In_4908);
or U474 (N_474,In_2776,In_3217);
or U475 (N_475,In_250,In_723);
nor U476 (N_476,In_4190,In_2304);
nor U477 (N_477,In_3456,In_4114);
nand U478 (N_478,In_2240,In_1094);
nand U479 (N_479,In_1277,In_912);
xor U480 (N_480,In_4901,In_4487);
and U481 (N_481,In_3274,In_4247);
nand U482 (N_482,In_4544,In_2207);
and U483 (N_483,In_2800,In_4439);
and U484 (N_484,In_4651,In_678);
nand U485 (N_485,In_2401,In_4359);
or U486 (N_486,In_2948,In_1846);
and U487 (N_487,In_3236,In_497);
or U488 (N_488,In_3117,In_4580);
nor U489 (N_489,In_2465,In_4953);
nand U490 (N_490,In_1420,In_2153);
xnor U491 (N_491,In_3003,In_680);
and U492 (N_492,In_944,In_3991);
nand U493 (N_493,In_3258,In_611);
nor U494 (N_494,In_4059,In_3);
xnor U495 (N_495,In_3619,In_1457);
or U496 (N_496,In_1605,In_3518);
nand U497 (N_497,In_740,In_1587);
or U498 (N_498,In_4842,In_3528);
nand U499 (N_499,In_3745,In_3350);
or U500 (N_500,In_2375,In_709);
nor U501 (N_501,In_1737,In_2594);
nand U502 (N_502,In_1734,In_960);
or U503 (N_503,In_4907,In_4180);
xnor U504 (N_504,In_4139,In_4185);
nand U505 (N_505,In_4161,In_764);
or U506 (N_506,In_321,In_726);
nand U507 (N_507,In_4988,In_884);
and U508 (N_508,In_2595,In_706);
or U509 (N_509,In_3149,In_4787);
and U510 (N_510,In_4915,In_4503);
xnor U511 (N_511,In_4770,In_1199);
xor U512 (N_512,In_690,In_1172);
or U513 (N_513,In_2390,In_4456);
xor U514 (N_514,In_4362,In_2888);
and U515 (N_515,In_3881,In_3057);
nand U516 (N_516,In_131,In_1266);
xor U517 (N_517,In_1484,In_657);
or U518 (N_518,In_654,In_4179);
xor U519 (N_519,In_3306,In_1083);
and U520 (N_520,In_2473,In_4208);
and U521 (N_521,In_619,In_4920);
xor U522 (N_522,In_2582,In_452);
nand U523 (N_523,In_4928,In_2514);
or U524 (N_524,In_2170,In_2892);
xor U525 (N_525,In_325,In_4083);
and U526 (N_526,In_4313,In_4312);
and U527 (N_527,In_4917,In_1235);
nor U528 (N_528,In_603,In_2338);
nor U529 (N_529,In_4535,In_2444);
nand U530 (N_530,In_735,In_3634);
xnor U531 (N_531,In_4115,In_4261);
nor U532 (N_532,In_575,In_4670);
and U533 (N_533,In_2852,In_4589);
nand U534 (N_534,In_486,In_434);
xnor U535 (N_535,In_1257,In_357);
nor U536 (N_536,In_1098,In_4586);
xnor U537 (N_537,In_3731,In_4810);
or U538 (N_538,In_3092,In_4710);
nand U539 (N_539,In_3479,In_4351);
nand U540 (N_540,In_2517,In_3169);
nor U541 (N_541,In_230,In_3102);
or U542 (N_542,In_3744,In_213);
or U543 (N_543,In_2369,In_3692);
nor U544 (N_544,In_2744,In_3021);
nand U545 (N_545,In_3051,In_1152);
nor U546 (N_546,In_243,In_1270);
nor U547 (N_547,In_2729,In_4467);
nand U548 (N_548,In_2254,In_1584);
or U549 (N_549,In_1157,In_3397);
and U550 (N_550,In_1739,In_4365);
nor U551 (N_551,In_2129,In_2589);
and U552 (N_552,In_3707,In_3006);
nand U553 (N_553,In_2650,In_3812);
xnor U554 (N_554,In_1304,In_1977);
or U555 (N_555,In_238,In_3012);
and U556 (N_556,In_3229,In_4611);
nor U557 (N_557,In_3014,In_3598);
xnor U558 (N_558,In_2115,In_896);
or U559 (N_559,In_3520,In_4356);
xnor U560 (N_560,In_1141,In_1866);
and U561 (N_561,In_1053,In_2459);
nor U562 (N_562,In_1331,In_977);
and U563 (N_563,In_3856,In_3111);
xor U564 (N_564,In_1738,In_3356);
or U565 (N_565,In_1848,In_3753);
xor U566 (N_566,In_4822,In_2119);
nand U567 (N_567,In_4355,In_61);
or U568 (N_568,In_3220,In_2389);
nor U569 (N_569,In_4443,In_2088);
nor U570 (N_570,In_1891,In_821);
and U571 (N_571,In_1601,In_4072);
or U572 (N_572,In_4170,In_1403);
nand U573 (N_573,In_2747,In_1750);
nor U574 (N_574,In_4784,In_3515);
and U575 (N_575,In_3871,In_4346);
xor U576 (N_576,In_2731,In_328);
or U577 (N_577,In_4967,In_534);
and U578 (N_578,In_1333,In_1530);
or U579 (N_579,In_3064,In_2907);
or U580 (N_580,In_3370,In_4014);
nand U581 (N_581,In_98,In_1390);
nor U582 (N_582,In_963,In_1193);
xor U583 (N_583,In_2239,In_518);
nor U584 (N_584,In_921,In_4488);
nand U585 (N_585,In_203,In_766);
or U586 (N_586,In_3131,In_3889);
xnor U587 (N_587,In_1687,In_4460);
nor U588 (N_588,In_2024,In_2613);
or U589 (N_589,In_4682,In_1313);
and U590 (N_590,In_4614,In_852);
or U591 (N_591,In_2794,In_2874);
nor U592 (N_592,In_2406,In_4673);
nand U593 (N_593,In_3799,In_2137);
nor U594 (N_594,In_1102,In_3901);
or U595 (N_595,In_3949,In_4269);
nand U596 (N_596,In_33,In_2477);
and U597 (N_597,In_4206,In_781);
xor U598 (N_598,In_2371,In_942);
nand U599 (N_599,In_2346,In_4070);
or U600 (N_600,In_3746,In_3829);
xor U601 (N_601,In_483,In_2839);
or U602 (N_602,In_1653,In_3001);
and U603 (N_603,In_880,In_1681);
nand U604 (N_604,In_2384,In_1768);
or U605 (N_605,In_2457,In_3309);
nand U606 (N_606,In_3050,In_1877);
or U607 (N_607,In_2915,In_720);
nor U608 (N_608,In_3646,In_1718);
nor U609 (N_609,In_4302,In_1575);
nor U610 (N_610,In_905,In_3960);
nor U611 (N_611,In_4432,In_1969);
and U612 (N_612,In_3622,In_1948);
xnor U613 (N_613,In_4,In_3360);
xnor U614 (N_614,In_1624,In_2533);
xnor U615 (N_615,In_732,In_4897);
nor U616 (N_616,In_2246,In_4134);
nand U617 (N_617,In_2333,In_2649);
and U618 (N_618,In_73,In_920);
xnor U619 (N_619,In_1400,In_4383);
xor U620 (N_620,In_348,In_3029);
nand U621 (N_621,In_1824,In_1110);
and U622 (N_622,In_2035,In_4236);
and U623 (N_623,In_898,In_4905);
or U624 (N_624,In_324,In_3689);
nand U625 (N_625,In_3365,In_718);
nor U626 (N_626,In_2743,In_828);
or U627 (N_627,In_1652,In_3353);
nor U628 (N_628,In_2281,In_2694);
or U629 (N_629,In_3712,In_3890);
xnor U630 (N_630,In_4085,In_1066);
xnor U631 (N_631,In_2728,In_2620);
nor U632 (N_632,In_418,In_1175);
and U633 (N_633,In_4244,In_1146);
xnor U634 (N_634,In_2220,In_3885);
xnor U635 (N_635,In_1808,In_1436);
nor U636 (N_636,In_1429,In_2675);
nand U637 (N_637,In_2230,In_582);
xor U638 (N_638,In_2261,In_2114);
nand U639 (N_639,In_679,In_3990);
or U640 (N_640,In_204,In_3095);
and U641 (N_641,In_234,In_4815);
nand U642 (N_642,In_1902,In_599);
nor U643 (N_643,In_3384,In_4218);
nand U644 (N_644,In_4952,In_2403);
nor U645 (N_645,In_3849,In_4363);
nand U646 (N_646,In_2645,In_337);
xnor U647 (N_647,In_1245,In_3591);
nor U648 (N_648,In_183,In_1710);
nand U649 (N_649,In_3104,In_2906);
nor U650 (N_650,In_4852,In_3997);
nor U651 (N_651,In_3032,In_1164);
and U652 (N_652,In_2837,In_2456);
nor U653 (N_653,In_3592,In_861);
and U654 (N_654,In_1419,In_1567);
and U655 (N_655,In_4246,In_3542);
xnor U656 (N_656,In_283,In_1240);
nand U657 (N_657,In_303,In_2531);
xnor U658 (N_658,In_3912,In_4334);
nor U659 (N_659,In_1865,In_1486);
and U660 (N_660,In_1747,In_3428);
and U661 (N_661,In_1641,In_4143);
nor U662 (N_662,In_3678,In_1079);
xor U663 (N_663,In_961,In_3396);
nor U664 (N_664,In_2344,In_1462);
and U665 (N_665,In_4858,In_4360);
nor U666 (N_666,In_1763,In_4973);
and U667 (N_667,In_3613,In_4027);
nand U668 (N_668,In_538,In_343);
nor U669 (N_669,In_3948,In_664);
nor U670 (N_670,In_4863,In_3113);
nor U671 (N_671,In_4561,In_2940);
nor U672 (N_672,In_3654,In_1368);
or U673 (N_673,In_666,In_3103);
nand U674 (N_674,In_4199,In_3037);
xnor U675 (N_675,In_4832,In_4198);
or U676 (N_676,In_397,In_999);
and U677 (N_677,In_2117,In_1143);
xor U678 (N_678,In_2247,In_860);
xnor U679 (N_679,In_2182,In_629);
or U680 (N_680,In_2931,In_4938);
nand U681 (N_681,In_892,In_408);
nand U682 (N_682,In_2053,In_4958);
and U683 (N_683,In_2831,In_3127);
nor U684 (N_684,In_2515,In_602);
xnor U685 (N_685,In_1771,In_4595);
nor U686 (N_686,In_4109,In_4209);
nor U687 (N_687,In_1564,In_1603);
nand U688 (N_688,In_4389,In_1508);
nand U689 (N_689,In_4394,In_4270);
and U690 (N_690,In_212,In_4657);
nand U691 (N_691,In_4173,In_235);
and U692 (N_692,In_1657,In_1291);
nor U693 (N_693,In_3672,In_4288);
nand U694 (N_694,In_3993,In_4142);
and U695 (N_695,In_876,In_539);
and U696 (N_696,In_84,In_3477);
nor U697 (N_697,In_1492,In_1854);
nor U698 (N_698,In_831,In_686);
xnor U699 (N_699,In_2964,In_3288);
nand U700 (N_700,In_2998,In_2709);
and U701 (N_701,In_1867,In_4644);
xnor U702 (N_702,In_143,In_1936);
xor U703 (N_703,In_4783,In_118);
nor U704 (N_704,In_1179,In_2586);
nor U705 (N_705,In_347,In_3784);
and U706 (N_706,In_2652,In_3438);
or U707 (N_707,In_739,In_2727);
or U708 (N_708,In_262,In_2922);
xor U709 (N_709,In_4164,In_558);
xnor U710 (N_710,In_1810,In_4441);
and U711 (N_711,In_923,In_1951);
or U712 (N_712,In_2503,In_2241);
nand U713 (N_713,In_596,In_37);
nor U714 (N_714,In_336,In_1664);
nand U715 (N_715,In_1337,In_4103);
or U716 (N_716,In_546,In_724);
xor U717 (N_717,In_924,In_1870);
xor U718 (N_718,In_1372,In_4331);
and U719 (N_719,In_2617,In_2894);
xor U720 (N_720,In_40,In_3393);
or U721 (N_721,In_3292,In_2499);
and U722 (N_722,In_936,In_3940);
nand U723 (N_723,In_407,In_4699);
or U724 (N_724,In_2073,In_1748);
nand U725 (N_725,In_701,In_865);
and U726 (N_726,In_4825,In_2025);
and U727 (N_727,In_4207,In_1896);
or U728 (N_728,In_1855,In_2529);
and U729 (N_729,In_3653,In_4094);
nand U730 (N_730,In_2588,In_338);
xnor U731 (N_731,In_296,In_4220);
xor U732 (N_732,In_940,In_3777);
nor U733 (N_733,In_3042,In_1373);
nor U734 (N_734,In_979,In_991);
nor U735 (N_735,In_3401,In_1837);
xnor U736 (N_736,In_906,In_913);
nand U737 (N_737,In_4562,In_4725);
and U738 (N_738,In_3211,In_4526);
or U739 (N_739,In_560,In_3935);
xnor U740 (N_740,In_1480,In_1906);
nand U741 (N_741,In_996,In_259);
nor U742 (N_742,In_3150,In_4172);
and U743 (N_743,In_364,In_4912);
xnor U744 (N_744,In_3823,In_3787);
nand U745 (N_745,In_3531,In_1452);
and U746 (N_746,In_4638,In_502);
nor U747 (N_747,In_2256,In_2680);
xor U748 (N_748,In_2091,In_4217);
or U749 (N_749,In_3242,In_2428);
xor U750 (N_750,In_3998,In_2659);
or U751 (N_751,In_4821,In_2606);
nand U752 (N_752,In_3756,In_1730);
or U753 (N_753,In_2277,In_4340);
nand U754 (N_754,In_773,In_3442);
xor U755 (N_755,In_2520,In_3193);
xnor U756 (N_756,In_4963,In_1982);
nand U757 (N_757,In_4748,In_4303);
xnor U758 (N_758,In_3418,In_2668);
xor U759 (N_759,In_1868,In_3284);
or U760 (N_760,In_3576,In_4759);
and U761 (N_761,In_959,In_1067);
nor U762 (N_762,In_2009,In_3106);
and U763 (N_763,In_1441,In_812);
nor U764 (N_764,In_2677,In_1060);
nor U765 (N_765,In_2786,In_201);
or U766 (N_766,In_797,In_4984);
nor U767 (N_767,In_3837,In_2909);
and U768 (N_768,In_2823,In_2188);
and U769 (N_769,In_479,In_3126);
xor U770 (N_770,In_0,In_3539);
nand U771 (N_771,In_814,In_3519);
or U772 (N_772,In_783,In_3156);
nand U773 (N_773,In_1350,In_4574);
nor U774 (N_774,In_2504,In_1698);
xnor U775 (N_775,In_3972,In_1955);
nand U776 (N_776,In_2113,In_3373);
xnor U777 (N_777,In_3077,In_4155);
and U778 (N_778,In_1482,In_4856);
nand U779 (N_779,In_1672,In_2442);
or U780 (N_780,In_3545,In_2565);
nand U781 (N_781,In_111,In_627);
and U782 (N_782,In_2492,In_2349);
nand U783 (N_783,In_1194,In_3761);
xor U784 (N_784,In_973,In_4570);
xor U785 (N_785,In_4044,In_1874);
and U786 (N_786,In_698,In_2976);
or U787 (N_787,In_2152,In_2469);
or U788 (N_788,In_4819,In_1880);
xor U789 (N_789,In_2769,In_82);
and U790 (N_790,In_4522,In_255);
nor U791 (N_791,In_1720,In_3167);
xnor U792 (N_792,In_839,In_2111);
or U793 (N_793,In_2079,In_4333);
or U794 (N_794,In_123,In_1113);
nand U795 (N_795,In_872,In_1826);
nor U796 (N_796,In_1376,In_1832);
and U797 (N_797,In_1799,In_1425);
and U798 (N_798,In_216,In_2959);
and U799 (N_799,In_3764,In_2811);
nor U800 (N_800,In_1809,In_1120);
nor U801 (N_801,In_1533,In_4260);
nor U802 (N_802,In_4343,In_836);
nor U803 (N_803,In_419,In_2534);
nand U804 (N_804,In_728,In_3532);
xor U805 (N_805,In_3204,In_3385);
or U806 (N_806,In_450,In_2641);
xor U807 (N_807,In_1064,In_366);
nor U808 (N_808,In_1985,In_3710);
xnor U809 (N_809,In_652,In_2843);
and U810 (N_810,In_2244,In_2150);
nand U811 (N_811,In_3927,In_428);
nand U812 (N_812,In_438,In_378);
xor U813 (N_813,In_1256,In_3146);
or U814 (N_814,In_4799,In_4681);
nand U815 (N_815,In_1946,In_4202);
nor U816 (N_816,In_2328,In_4489);
nand U817 (N_817,In_2703,In_4676);
xnor U818 (N_818,In_4817,In_1956);
or U819 (N_819,In_1319,In_2116);
and U820 (N_820,In_2949,In_1133);
nor U821 (N_821,In_3315,In_3036);
xnor U822 (N_822,In_4330,In_1182);
nand U823 (N_823,In_1301,In_3478);
or U824 (N_824,In_3416,In_1800);
nand U825 (N_825,In_3977,In_3820);
or U826 (N_826,In_4855,In_2421);
nand U827 (N_827,In_2899,In_3900);
nand U828 (N_828,In_4551,In_294);
nor U829 (N_829,In_682,In_458);
and U830 (N_830,In_4426,In_1234);
nand U831 (N_831,In_805,In_760);
xnor U832 (N_832,In_3505,In_858);
nand U833 (N_833,In_115,In_1474);
xnor U834 (N_834,In_3269,In_741);
and U835 (N_835,In_1161,In_925);
xnor U836 (N_836,In_2757,In_1933);
or U837 (N_837,In_3763,In_2859);
and U838 (N_838,In_1671,In_3827);
xnor U839 (N_839,In_844,In_2162);
and U840 (N_840,In_3758,In_1380);
nand U841 (N_841,In_3307,In_1850);
nand U842 (N_842,In_2006,In_2319);
nand U843 (N_843,In_1852,In_1302);
nand U844 (N_844,In_2841,In_2426);
or U845 (N_845,In_1841,In_2092);
xor U846 (N_846,In_1377,In_3509);
xor U847 (N_847,In_3869,In_2044);
nor U848 (N_848,In_615,In_309);
nor U849 (N_849,In_3819,In_512);
and U850 (N_850,In_4205,In_2687);
or U851 (N_851,In_3958,In_333);
nor U852 (N_852,In_3790,In_2471);
and U853 (N_853,In_2107,In_4012);
nor U854 (N_854,In_2924,In_2098);
or U855 (N_855,In_4796,In_506);
nand U856 (N_856,In_4492,In_2285);
nor U857 (N_857,In_417,In_972);
nor U858 (N_858,In_170,In_3933);
nor U859 (N_859,In_1966,In_4554);
nand U860 (N_860,In_4228,In_3465);
and U861 (N_861,In_3387,In_1109);
or U862 (N_862,In_1057,In_125);
and U863 (N_863,In_725,In_2064);
nor U864 (N_864,In_2511,In_1823);
nor U865 (N_865,In_2961,In_1184);
and U866 (N_866,In_763,In_2396);
nand U867 (N_867,In_1298,In_2913);
and U868 (N_868,In_2348,In_1447);
or U869 (N_869,In_1203,In_326);
or U870 (N_870,In_922,In_2289);
nor U871 (N_871,In_733,In_2059);
or U872 (N_872,In_1475,In_2754);
nand U873 (N_873,In_4329,In_4903);
nor U874 (N_874,In_2443,In_4200);
or U875 (N_875,In_3550,In_3651);
and U876 (N_876,In_1509,In_1662);
nor U877 (N_877,In_4277,In_470);
xnor U878 (N_878,In_1658,In_3817);
nor U879 (N_879,In_928,In_429);
or U880 (N_880,In_3637,In_4287);
nor U881 (N_881,In_1616,In_3946);
or U882 (N_882,In_4282,In_1151);
or U883 (N_883,In_2462,In_1965);
and U884 (N_884,In_2510,In_295);
xnor U885 (N_885,In_845,In_1661);
and U886 (N_886,In_3244,In_3639);
nand U887 (N_887,In_504,In_454);
or U888 (N_888,In_4892,In_1087);
or U889 (N_889,In_3806,In_2656);
xor U890 (N_890,In_2476,In_4781);
nor U891 (N_891,In_3929,In_1557);
nand U892 (N_892,In_4861,In_175);
and U893 (N_893,In_2545,In_2213);
nor U894 (N_894,In_4581,In_524);
nor U895 (N_895,In_3363,In_3775);
nand U896 (N_896,In_3934,In_2121);
and U897 (N_897,In_1999,In_4194);
or U898 (N_898,In_1743,In_1128);
nor U899 (N_899,In_2105,In_1633);
and U900 (N_900,In_2160,In_122);
nand U901 (N_901,In_683,In_81);
nand U902 (N_902,In_1042,In_3841);
nand U903 (N_903,In_610,In_2527);
or U904 (N_904,In_2625,In_4923);
or U905 (N_905,In_976,In_3955);
nand U906 (N_906,In_4514,In_1858);
and U907 (N_907,In_268,In_1074);
nor U908 (N_908,In_4377,In_2127);
nand U909 (N_909,In_4876,In_2479);
nor U910 (N_910,In_356,In_1638);
xor U911 (N_911,In_1519,In_569);
nor U912 (N_912,In_841,In_2286);
and U913 (N_913,In_1003,In_883);
or U914 (N_914,In_3514,In_1000);
or U915 (N_915,In_4062,In_4249);
xnor U916 (N_916,In_4324,In_2052);
nand U917 (N_917,In_647,In_1772);
and U918 (N_918,In_1465,In_307);
nor U919 (N_919,In_3480,In_293);
nand U920 (N_920,In_2973,In_1396);
or U921 (N_921,In_2362,In_3737);
xor U922 (N_922,In_2616,In_3814);
or U923 (N_923,In_943,In_3081);
or U924 (N_924,In_1384,In_3988);
xor U925 (N_925,In_573,In_4451);
or U926 (N_926,In_3671,In_1423);
and U927 (N_927,In_4569,In_3232);
nand U928 (N_928,In_2030,In_2377);
and U929 (N_929,In_172,In_869);
xor U930 (N_930,In_640,In_4909);
or U931 (N_931,In_4000,In_4125);
nand U932 (N_932,In_2050,In_4430);
nor U933 (N_933,In_3059,In_4870);
xnor U934 (N_934,In_1523,In_1712);
xnor U935 (N_935,In_3780,In_1364);
or U936 (N_936,In_2321,In_2548);
xnor U937 (N_937,In_3019,In_4592);
nand U938 (N_938,In_3910,In_1905);
xnor U939 (N_939,In_1945,In_4299);
nand U940 (N_940,In_1990,In_2132);
nand U941 (N_941,In_3504,In_3164);
nor U942 (N_942,In_126,In_2472);
nand U943 (N_943,In_449,In_1342);
nand U944 (N_944,In_2898,In_4416);
nor U945 (N_945,In_4729,In_2882);
xnor U946 (N_946,In_1269,In_2104);
nand U947 (N_947,In_1352,In_932);
nor U948 (N_948,In_3158,In_1328);
nor U949 (N_949,In_3866,In_749);
nor U950 (N_950,In_2224,In_489);
nand U951 (N_951,In_310,In_4160);
or U952 (N_952,In_1684,In_3727);
and U953 (N_953,In_3016,In_3720);
or U954 (N_954,In_4005,In_3132);
nor U955 (N_955,In_934,In_1230);
nor U956 (N_956,In_278,In_3413);
or U957 (N_957,In_2062,In_256);
or U958 (N_958,In_1180,In_617);
xnor U959 (N_959,In_2179,In_784);
or U960 (N_960,In_638,In_437);
nand U961 (N_961,In_141,In_3446);
and U962 (N_962,In_574,In_4686);
and U963 (N_963,In_1494,In_1752);
nand U964 (N_964,In_1134,In_4276);
nand U965 (N_965,In_3682,In_1449);
xor U966 (N_966,In_2489,In_395);
or U967 (N_967,In_4188,In_4041);
and U968 (N_968,In_3585,In_2047);
and U969 (N_969,In_4422,In_2669);
and U970 (N_970,In_2782,In_3008);
nand U971 (N_971,In_2855,In_601);
and U972 (N_972,In_901,In_1650);
nand U973 (N_973,In_2814,In_2562);
or U974 (N_974,In_752,In_22);
and U975 (N_975,In_2937,In_3461);
nor U976 (N_976,In_4864,In_4337);
and U977 (N_977,In_4264,In_1119);
xnor U978 (N_978,In_655,In_318);
nor U979 (N_979,In_4792,In_1939);
nand U980 (N_980,In_742,In_53);
nand U981 (N_981,In_4253,In_2288);
xnor U982 (N_982,In_1978,In_1843);
xor U983 (N_983,In_3510,In_1571);
xnor U984 (N_984,In_1784,In_3233);
nand U985 (N_985,In_3833,In_3256);
nand U986 (N_986,In_1077,In_2490);
nand U987 (N_987,In_1862,In_2826);
nor U988 (N_988,In_4382,In_1770);
xor U989 (N_989,In_11,In_3425);
or U990 (N_990,In_1726,In_2087);
nor U991 (N_991,In_3573,In_2835);
nand U992 (N_992,In_3441,In_1696);
nand U993 (N_993,In_1606,In_2474);
and U994 (N_994,In_3283,In_389);
or U995 (N_995,In_3966,In_625);
and U996 (N_996,In_1678,In_3791);
and U997 (N_997,In_4450,In_1366);
or U998 (N_998,In_1807,In_3445);
nor U999 (N_999,In_2849,In_1914);
nor U1000 (N_1000,In_4516,In_1864);
xnor U1001 (N_1001,In_3649,In_2296);
xor U1002 (N_1002,In_4719,In_3913);
or U1003 (N_1003,In_3850,In_3406);
nand U1004 (N_1004,In_3404,In_3225);
nor U1005 (N_1005,In_451,In_1627);
xnor U1006 (N_1006,In_3340,In_1338);
or U1007 (N_1007,In_1585,In_3612);
nor U1008 (N_1008,In_4994,In_4517);
xnor U1009 (N_1009,In_3311,In_3291);
and U1010 (N_1010,In_1595,In_3800);
and U1011 (N_1011,In_637,In_4743);
and U1012 (N_1012,In_962,In_244);
nor U1013 (N_1013,In_3116,In_744);
nor U1014 (N_1014,In_3450,In_2952);
nor U1015 (N_1015,In_2419,In_1443);
xor U1016 (N_1016,In_2923,In_2155);
xor U1017 (N_1017,In_4307,In_72);
and U1018 (N_1018,In_2464,In_708);
nand U1019 (N_1019,In_3530,In_4267);
nand U1020 (N_1020,In_3569,In_491);
nor U1021 (N_1021,In_1628,In_3316);
nand U1022 (N_1022,In_3578,In_1101);
or U1023 (N_1023,In_1818,In_1105);
nor U1024 (N_1024,In_1786,In_4136);
or U1025 (N_1025,In_1496,In_4709);
and U1026 (N_1026,In_390,In_3381);
xnor U1027 (N_1027,In_3675,In_308);
xor U1028 (N_1028,In_1198,In_3996);
xor U1029 (N_1029,In_1689,In_1205);
nand U1030 (N_1030,In_3751,In_1899);
nand U1031 (N_1031,In_1426,In_1322);
nand U1032 (N_1032,In_253,In_2339);
or U1033 (N_1033,In_4191,In_1259);
and U1034 (N_1034,In_3544,In_2276);
nor U1035 (N_1035,In_153,In_1630);
nand U1036 (N_1036,In_649,In_4017);
and U1037 (N_1037,In_824,In_1876);
xnor U1038 (N_1038,In_734,In_2273);
or U1039 (N_1039,In_3614,In_138);
or U1040 (N_1040,In_124,In_4493);
and U1041 (N_1041,In_981,In_598);
nor U1042 (N_1042,In_2798,In_3852);
or U1043 (N_1043,In_2448,In_1766);
nor U1044 (N_1044,In_139,In_4521);
and U1045 (N_1045,In_1129,In_1779);
xor U1046 (N_1046,In_4395,In_4240);
and U1047 (N_1047,In_2048,In_3502);
nand U1048 (N_1048,In_1392,In_1336);
xnor U1049 (N_1049,In_2458,In_2935);
xor U1050 (N_1050,In_4736,In_1845);
or U1051 (N_1051,In_2232,In_3899);
or U1052 (N_1052,In_1911,In_4090);
and U1053 (N_1053,In_3714,In_2372);
or U1054 (N_1054,In_715,In_3388);
or U1055 (N_1055,In_2146,In_1721);
xor U1056 (N_1056,In_3513,In_4498);
xnor U1057 (N_1057,In_63,In_2488);
nand U1058 (N_1058,In_1100,In_1135);
or U1059 (N_1059,In_1226,In_4721);
xor U1060 (N_1060,In_1791,In_339);
or U1061 (N_1061,In_4379,In_676);
xor U1062 (N_1062,In_1160,In_1176);
or U1063 (N_1063,In_1271,In_4671);
or U1064 (N_1064,In_411,In_1548);
or U1065 (N_1065,In_4279,In_2012);
nand U1066 (N_1066,In_2156,In_4407);
xor U1067 (N_1067,In_4210,In_456);
and U1068 (N_1068,In_4197,In_4401);
xnor U1069 (N_1069,In_1278,In_4757);
xor U1070 (N_1070,In_1817,In_660);
nor U1071 (N_1071,In_4111,In_1701);
and U1072 (N_1072,In_92,In_3367);
or U1073 (N_1073,In_2099,In_2537);
nand U1074 (N_1074,In_3305,In_964);
and U1075 (N_1075,In_1938,In_810);
or U1076 (N_1076,In_2991,In_4539);
nand U1077 (N_1077,In_3650,In_866);
xor U1078 (N_1078,In_2524,In_2233);
or U1079 (N_1079,In_4737,In_3759);
nand U1080 (N_1080,In_4960,In_4225);
nor U1081 (N_1081,In_1531,In_4765);
xnor U1082 (N_1082,In_2930,In_2078);
xor U1083 (N_1083,In_1275,In_3076);
xnor U1084 (N_1084,In_2070,In_4906);
nor U1085 (N_1085,In_4890,In_4564);
nor U1086 (N_1086,In_2205,In_4524);
xor U1087 (N_1087,In_1753,In_282);
nor U1088 (N_1088,In_1002,In_2893);
and U1089 (N_1089,In_2142,In_3072);
or U1090 (N_1090,In_4459,In_815);
nor U1091 (N_1091,In_3214,In_1767);
xor U1092 (N_1092,In_406,In_162);
or U1093 (N_1093,In_31,In_3410);
and U1094 (N_1094,In_3067,In_1405);
or U1095 (N_1095,In_3564,In_3503);
and U1096 (N_1096,In_2229,In_4768);
nor U1097 (N_1097,In_1574,In_1285);
xor U1098 (N_1098,In_88,In_2636);
xor U1099 (N_1099,In_3750,In_1520);
nand U1100 (N_1100,In_4758,In_488);
and U1101 (N_1101,In_4593,In_2173);
or U1102 (N_1102,In_1341,In_3318);
nor U1103 (N_1103,In_2688,In_3832);
and U1104 (N_1104,In_1524,In_185);
xor U1105 (N_1105,In_457,In_3571);
nor U1106 (N_1106,In_3224,In_13);
and U1107 (N_1107,In_4323,In_3186);
nand U1108 (N_1108,In_2020,In_4001);
or U1109 (N_1109,In_2388,In_2579);
nand U1110 (N_1110,In_2577,In_791);
and U1111 (N_1111,In_639,In_3255);
nand U1112 (N_1112,In_992,In_2507);
and U1113 (N_1113,In_21,In_1223);
and U1114 (N_1114,In_3341,In_4505);
nand U1115 (N_1115,In_2096,In_1645);
nand U1116 (N_1116,In_3264,In_4576);
nand U1117 (N_1117,In_2869,In_174);
xnor U1118 (N_1118,In_2570,In_3685);
or U1119 (N_1119,In_3702,In_1335);
xor U1120 (N_1120,In_1719,In_1699);
nor U1121 (N_1121,In_2832,In_4816);
nor U1122 (N_1122,In_1078,In_2872);
nand U1123 (N_1123,In_1206,In_4166);
and U1124 (N_1124,In_2324,In_3068);
xnor U1125 (N_1125,In_2227,In_4391);
and U1126 (N_1126,In_3281,In_548);
xnor U1127 (N_1127,In_2357,In_2796);
nand U1128 (N_1128,In_4212,In_3002);
nand U1129 (N_1129,In_3865,In_335);
or U1130 (N_1130,In_2355,In_2103);
and U1131 (N_1131,In_300,In_3698);
nand U1132 (N_1132,In_2222,In_2447);
or U1133 (N_1133,In_4951,In_2501);
xor U1134 (N_1134,In_4786,In_4885);
nor U1135 (N_1135,In_688,In_607);
nor U1136 (N_1136,In_4608,In_4255);
nor U1137 (N_1137,In_1056,In_949);
nand U1138 (N_1138,In_4654,In_1358);
nand U1139 (N_1139,In_2752,In_1458);
or U1140 (N_1140,In_550,In_195);
or U1141 (N_1141,In_1095,In_3240);
nor U1142 (N_1142,In_4708,In_4823);
nand U1143 (N_1143,In_1549,In_620);
nor U1144 (N_1144,In_1534,In_533);
xor U1145 (N_1145,In_1732,In_885);
nand U1146 (N_1146,In_363,In_2140);
and U1147 (N_1147,In_3752,In_2766);
xnor U1148 (N_1148,In_4268,In_2783);
and U1149 (N_1149,In_4263,In_2017);
nor U1150 (N_1150,In_2712,In_359);
and U1151 (N_1151,In_3010,In_767);
or U1152 (N_1152,In_2916,In_4306);
xnor U1153 (N_1153,In_930,In_3163);
and U1154 (N_1154,In_3642,In_2543);
and U1155 (N_1155,In_4693,In_362);
nor U1156 (N_1156,In_2395,In_4049);
nor U1157 (N_1157,In_4373,In_3496);
or U1158 (N_1158,In_399,In_4835);
xor U1159 (N_1159,In_209,In_642);
and U1160 (N_1160,In_758,In_4871);
nor U1161 (N_1161,In_4018,In_4463);
xnor U1162 (N_1162,In_3555,In_2902);
and U1163 (N_1163,In_3017,In_1889);
or U1164 (N_1164,In_103,In_64);
nand U1165 (N_1165,In_1483,In_4132);
nand U1166 (N_1166,In_3854,In_1934);
and U1167 (N_1167,In_4986,In_2049);
xnor U1168 (N_1168,In_381,In_675);
and U1169 (N_1169,In_4944,In_2279);
nand U1170 (N_1170,In_2678,In_3657);
nor U1171 (N_1171,In_2666,In_2483);
xnor U1172 (N_1172,In_3376,In_2327);
and U1173 (N_1173,In_1686,In_2879);
or U1174 (N_1174,In_2591,In_4336);
nand U1175 (N_1175,In_2165,In_3846);
nor U1176 (N_1176,In_1387,In_2637);
xnor U1177 (N_1177,In_3141,In_1063);
or U1178 (N_1178,In_2439,In_2951);
nor U1179 (N_1179,In_1124,In_3825);
and U1180 (N_1180,In_3200,In_3184);
nor U1181 (N_1181,In_1444,In_693);
or U1182 (N_1182,In_1932,In_2711);
or U1183 (N_1183,In_2981,In_4508);
nor U1184 (N_1184,In_1655,In_4033);
xnor U1185 (N_1185,In_2890,In_827);
and U1186 (N_1186,In_1884,In_4226);
nor U1187 (N_1187,In_2485,In_3999);
and U1188 (N_1188,In_1070,In_422);
and U1189 (N_1189,In_2002,In_4798);
nand U1190 (N_1190,In_3919,In_1061);
nor U1191 (N_1191,In_3920,In_1200);
or U1192 (N_1192,In_3082,In_3839);
nor U1193 (N_1193,In_4024,In_3595);
xor U1194 (N_1194,In_1090,In_24);
or U1195 (N_1195,In_583,In_2889);
xor U1196 (N_1196,In_1931,In_3128);
xor U1197 (N_1197,In_659,In_415);
xnor U1198 (N_1198,In_3982,In_4107);
or U1199 (N_1199,In_2310,In_2987);
or U1200 (N_1200,In_1915,In_1153);
nand U1201 (N_1201,In_2060,In_2779);
xor U1202 (N_1202,In_4772,In_3299);
and U1203 (N_1203,In_79,In_4192);
nand U1204 (N_1204,In_1033,In_1814);
and U1205 (N_1205,In_1013,In_2287);
or U1206 (N_1206,In_3079,In_1115);
nor U1207 (N_1207,In_2812,In_3906);
xor U1208 (N_1208,In_4553,In_1685);
xor U1209 (N_1209,In_4678,In_4648);
nor U1210 (N_1210,In_4429,In_2878);
and U1211 (N_1211,In_3362,In_4934);
xnor U1212 (N_1212,In_4004,In_3183);
or U1213 (N_1213,In_2822,In_1258);
or U1214 (N_1214,In_3891,In_1963);
nor U1215 (N_1215,In_3443,In_527);
nor U1216 (N_1216,In_2124,In_1609);
nor U1217 (N_1217,In_3334,In_2559);
nand U1218 (N_1218,In_1,In_4639);
nand U1219 (N_1219,In_2928,In_2029);
or U1220 (N_1220,In_4623,In_1500);
xnor U1221 (N_1221,In_4241,In_616);
and U1222 (N_1222,In_3176,In_3864);
nand U1223 (N_1223,In_1093,In_4820);
nand U1224 (N_1224,In_1091,In_193);
or U1225 (N_1225,In_1267,In_3471);
nor U1226 (N_1226,In_1502,In_3191);
or U1227 (N_1227,In_4585,In_1438);
or U1228 (N_1228,In_4374,In_107);
nor U1229 (N_1229,In_1881,In_1514);
or U1230 (N_1230,In_3093,In_3380);
and U1231 (N_1231,In_4297,In_802);
nand U1232 (N_1232,In_4785,In_4691);
or U1233 (N_1233,In_753,In_1973);
and U1234 (N_1234,In_3809,In_3483);
or U1235 (N_1235,In_4943,In_1019);
nand U1236 (N_1236,In_4827,In_58);
and U1237 (N_1237,In_1219,In_967);
or U1238 (N_1238,In_554,In_1015);
xor U1239 (N_1239,In_3207,In_4314);
and U1240 (N_1240,In_375,In_2042);
or U1241 (N_1241,In_1456,In_4669);
nand U1242 (N_1242,In_448,In_2386);
nor U1243 (N_1243,In_263,In_4233);
nor U1244 (N_1244,In_3230,In_4118);
and U1245 (N_1245,In_2546,In_3914);
nand U1246 (N_1246,In_3023,In_3795);
and U1247 (N_1247,In_4918,In_2236);
and U1248 (N_1248,In_2493,In_878);
nor U1249 (N_1249,In_2411,In_10);
or U1250 (N_1250,In_1044,In_2268);
nand U1251 (N_1251,In_3770,In_4751);
and U1252 (N_1252,In_2221,In_4734);
nand U1253 (N_1253,In_4766,In_980);
nand U1254 (N_1254,In_3411,In_202);
and U1255 (N_1255,In_3499,In_994);
xnor U1256 (N_1256,In_4696,In_4980);
or U1257 (N_1257,In_2158,In_4293);
and U1258 (N_1258,In_2228,In_2200);
and U1259 (N_1259,In_4006,In_4392);
nor U1260 (N_1260,In_1622,In_2218);
or U1261 (N_1261,In_3359,In_2563);
nor U1262 (N_1262,In_829,In_4597);
nand U1263 (N_1263,In_1986,In_1890);
xnor U1264 (N_1264,In_4126,In_4002);
xnor U1265 (N_1265,In_4425,In_382);
or U1266 (N_1266,In_4145,In_4712);
xor U1267 (N_1267,In_2821,In_2429);
or U1268 (N_1268,In_3454,In_3875);
or U1269 (N_1269,In_1516,In_3030);
nor U1270 (N_1270,In_2449,In_233);
and U1271 (N_1271,In_787,In_206);
nor U1272 (N_1272,In_2383,In_1190);
and U1273 (N_1273,In_471,In_1551);
xnor U1274 (N_1274,In_4052,In_2707);
nor U1275 (N_1275,In_969,In_1300);
xor U1276 (N_1276,In_1783,In_4060);
nand U1277 (N_1277,In_2732,In_2646);
and U1278 (N_1278,In_75,In_2572);
nor U1279 (N_1279,In_2966,In_4828);
and U1280 (N_1280,In_517,In_1450);
xor U1281 (N_1281,In_4795,In_2682);
xor U1282 (N_1282,In_1220,In_1122);
xnor U1283 (N_1283,In_3945,In_330);
or U1284 (N_1284,In_4367,In_3346);
nand U1285 (N_1285,In_1422,In_2080);
nor U1286 (N_1286,In_1560,In_4186);
and U1287 (N_1287,In_1081,In_3025);
nor U1288 (N_1288,In_3320,In_3261);
and U1289 (N_1289,In_2260,In_463);
nor U1290 (N_1290,In_1459,In_254);
xor U1291 (N_1291,In_2143,In_2943);
or U1292 (N_1292,In_2178,In_3683);
or U1293 (N_1293,In_48,In_4437);
or U1294 (N_1294,In_4058,In_2380);
and U1295 (N_1295,In_4797,In_3785);
nand U1296 (N_1296,In_4245,In_3366);
and U1297 (N_1297,In_4193,In_2011);
nor U1298 (N_1298,In_2550,In_350);
or U1299 (N_1299,In_614,In_1629);
nand U1300 (N_1300,In_2317,In_3994);
and U1301 (N_1301,In_570,In_4636);
xnor U1302 (N_1302,In_4902,In_148);
nor U1303 (N_1303,In_1086,In_1197);
and U1304 (N_1304,In_543,In_2963);
or U1305 (N_1305,In_1820,In_38);
xor U1306 (N_1306,In_2345,In_3324);
and U1307 (N_1307,In_813,In_2359);
nand U1308 (N_1308,In_4110,In_2329);
or U1309 (N_1309,In_353,In_251);
nor U1310 (N_1310,In_1210,In_2237);
and U1311 (N_1311,In_1409,In_1207);
nor U1312 (N_1312,In_4560,In_25);
and U1313 (N_1313,In_4703,In_4301);
nor U1314 (N_1314,In_4124,In_761);
or U1315 (N_1315,In_1434,In_1983);
or U1316 (N_1316,In_69,In_3928);
nand U1317 (N_1317,In_2201,In_3834);
nor U1318 (N_1318,In_4806,In_843);
nor U1319 (N_1319,In_1950,In_2451);
nor U1320 (N_1320,In_1903,In_210);
nand U1321 (N_1321,In_2884,In_1365);
xnor U1322 (N_1322,In_2671,In_4895);
or U1323 (N_1323,In_4275,In_1288);
or U1324 (N_1324,In_1654,In_3083);
or U1325 (N_1325,In_755,In_3656);
or U1326 (N_1326,In_4996,In_2717);
xor U1327 (N_1327,In_771,In_4084);
nor U1328 (N_1328,In_2532,In_2413);
nor U1329 (N_1329,In_3584,In_2438);
and U1330 (N_1330,In_4501,In_2558);
xnor U1331 (N_1331,In_4731,In_729);
xor U1332 (N_1332,In_823,In_1308);
xnor U1333 (N_1333,In_1611,In_1673);
xnor U1334 (N_1334,In_950,In_1553);
or U1335 (N_1335,In_914,In_899);
xor U1336 (N_1336,In_501,In_1397);
and U1337 (N_1337,In_4578,In_1695);
nand U1338 (N_1338,In_1224,In_3676);
xor U1339 (N_1339,In_631,In_4073);
and U1340 (N_1340,In_650,In_3681);
or U1341 (N_1341,In_2938,In_2840);
and U1342 (N_1342,In_1030,In_3647);
and U1343 (N_1343,In_3467,In_1104);
xnor U1344 (N_1344,In_1597,In_908);
and U1345 (N_1345,In_1831,In_2982);
or U1346 (N_1346,In_15,In_1541);
xnor U1347 (N_1347,In_646,In_2484);
xnor U1348 (N_1348,In_4151,In_2528);
xor U1349 (N_1349,In_1382,In_3040);
or U1350 (N_1350,In_2210,In_1588);
or U1351 (N_1351,In_4420,In_2068);
nand U1352 (N_1352,In_3562,In_1825);
or U1353 (N_1353,In_3674,In_3482);
nor U1354 (N_1354,In_1241,In_4752);
nand U1355 (N_1355,In_4689,In_4533);
and U1356 (N_1356,In_2647,In_4956);
nand U1357 (N_1357,In_485,In_867);
and U1358 (N_1358,In_1272,In_1360);
nand U1359 (N_1359,In_2692,In_4499);
or U1360 (N_1360,In_478,In_2015);
nor U1361 (N_1361,In_1290,In_4495);
and U1362 (N_1362,In_2306,In_2226);
xor U1363 (N_1363,In_2144,In_4350);
or U1364 (N_1364,In_3983,In_859);
xnor U1365 (N_1365,In_2214,In_3939);
and U1366 (N_1366,In_3386,In_3953);
nor U1367 (N_1367,In_2995,In_2632);
or U1368 (N_1368,In_1754,In_4515);
nor U1369 (N_1369,In_3655,In_1391);
or U1370 (N_1370,In_717,In_1920);
nor U1371 (N_1371,In_3709,In_1279);
nor U1372 (N_1372,In_4679,In_155);
nor U1373 (N_1373,In_588,In_712);
nor U1374 (N_1374,In_1233,In_776);
nor U1375 (N_1375,In_3857,In_2676);
xor U1376 (N_1376,In_1317,In_4484);
or U1377 (N_1377,In_1634,In_4730);
nor U1378 (N_1378,In_687,In_1195);
nand U1379 (N_1379,In_2016,In_1048);
nor U1380 (N_1380,In_1715,In_2644);
nor U1381 (N_1381,In_377,In_1949);
and U1382 (N_1382,In_3842,In_3589);
xor U1383 (N_1383,In_4531,In_2708);
and U1384 (N_1384,In_4384,In_2353);
nand U1385 (N_1385,In_1683,In_3154);
and U1386 (N_1386,In_4529,In_3950);
or U1387 (N_1387,In_3686,In_3234);
or U1388 (N_1388,In_147,In_3020);
nor U1389 (N_1389,In_1251,In_3099);
or U1390 (N_1390,In_4357,In_3730);
and U1391 (N_1391,In_4502,In_292);
and U1392 (N_1392,In_4853,In_4534);
xor U1393 (N_1393,In_151,In_3044);
nand U1394 (N_1394,In_1998,In_1873);
nand U1395 (N_1395,In_1020,In_55);
nand U1396 (N_1396,In_3252,In_4137);
and U1397 (N_1397,In_3056,In_987);
or U1398 (N_1398,In_2803,In_939);
and U1399 (N_1399,In_956,In_2385);
nor U1400 (N_1400,In_4602,In_1088);
xor U1401 (N_1401,In_4042,In_3660);
nand U1402 (N_1402,In_4698,In_2801);
and U1403 (N_1403,In_2263,In_847);
nand U1404 (N_1404,In_2560,In_496);
or U1405 (N_1405,In_3859,In_487);
nor U1406 (N_1406,In_2698,In_3524);
nor U1407 (N_1407,In_1345,In_3623);
and U1408 (N_1408,In_2084,In_1374);
and U1409 (N_1409,In_1941,In_1600);
nand U1410 (N_1410,In_3970,In_2301);
or U1411 (N_1411,In_4841,In_3776);
and U1412 (N_1412,In_4480,In_3312);
and U1413 (N_1413,In_135,In_595);
and U1414 (N_1414,In_1813,In_4859);
xnor U1415 (N_1415,In_4922,In_3405);
nand U1416 (N_1416,In_70,In_2135);
xor U1417 (N_1417,In_4632,In_403);
and U1418 (N_1418,In_2225,In_345);
nand U1419 (N_1419,In_2683,In_4294);
xnor U1420 (N_1420,In_778,In_3151);
nor U1421 (N_1421,In_157,In_1222);
and U1422 (N_1422,In_2942,In_4507);
and U1423 (N_1423,In_2257,In_564);
nand U1424 (N_1424,In_462,In_2095);
nand U1425 (N_1425,In_1010,In_1007);
or U1426 (N_1426,In_3332,In_2664);
nor U1427 (N_1427,In_35,In_3119);
nor U1428 (N_1428,In_2853,In_1667);
xnor U1429 (N_1429,In_4485,In_628);
or U1430 (N_1430,In_2022,In_2337);
or U1431 (N_1431,In_1156,In_275);
nand U1432 (N_1432,In_2340,In_158);
xor U1433 (N_1433,In_2764,In_4149);
nand U1434 (N_1434,In_1371,In_4328);
nand U1435 (N_1435,In_3917,In_4652);
xnor U1436 (N_1436,In_465,In_1024);
or U1437 (N_1437,In_4089,In_352);
and U1438 (N_1438,In_4500,In_1639);
and U1439 (N_1439,In_2373,In_738);
nand U1440 (N_1440,In_2581,In_4803);
or U1441 (N_1441,In_2897,In_2599);
nor U1442 (N_1442,In_4941,In_3608);
xnor U1443 (N_1443,In_4026,In_3098);
and U1444 (N_1444,In_1142,In_1536);
nor U1445 (N_1445,In_4793,In_941);
nand U1446 (N_1446,In_1640,In_2130);
xor U1447 (N_1447,In_1315,In_4948);
nor U1448 (N_1448,In_1907,In_4647);
nor U1449 (N_1449,In_4344,In_1957);
xnor U1450 (N_1450,In_2986,In_1346);
xnor U1451 (N_1451,In_4285,In_3235);
nand U1452 (N_1452,In_3802,In_3130);
and U1453 (N_1453,In_1406,In_2186);
and U1454 (N_1454,In_320,In_3989);
and U1455 (N_1455,In_4674,In_41);
xnor U1456 (N_1456,In_4256,In_4714);
and U1457 (N_1457,In_2726,In_97);
and U1458 (N_1458,In_1511,In_62);
and U1459 (N_1459,In_2223,In_1132);
nor U1460 (N_1460,In_3831,In_2309);
xnor U1461 (N_1461,In_3490,In_2748);
or U1462 (N_1462,In_1499,In_2547);
xnor U1463 (N_1463,In_4497,In_119);
nor U1464 (N_1464,In_3088,In_710);
and U1465 (N_1465,In_4831,In_3383);
or U1466 (N_1466,In_4889,In_4883);
and U1467 (N_1467,In_3560,In_1168);
and U1468 (N_1468,In_3783,In_4348);
nor U1469 (N_1469,In_2513,In_3961);
xnor U1470 (N_1470,In_4718,In_4064);
nor U1471 (N_1471,In_1260,In_2366);
or U1472 (N_1472,In_495,In_3355);
nor U1473 (N_1473,In_3326,In_711);
and U1474 (N_1474,In_393,In_3122);
or U1475 (N_1475,In_3475,In_4921);
or U1476 (N_1476,In_1051,In_1408);
nand U1477 (N_1477,In_4408,In_3394);
xnor U1478 (N_1478,In_319,In_826);
xor U1479 (N_1479,In_591,In_2730);
nand U1480 (N_1480,In_1103,In_3194);
xor U1481 (N_1481,In_68,In_4530);
or U1482 (N_1482,In_1707,In_3472);
or U1483 (N_1483,In_1218,In_3047);
and U1484 (N_1484,In_2264,In_4057);
nor U1485 (N_1485,In_1618,In_3173);
nand U1486 (N_1486,In_1043,In_1741);
nor U1487 (N_1487,In_4761,In_1668);
nor U1488 (N_1488,In_3638,In_4424);
nand U1489 (N_1489,In_159,In_846);
nor U1490 (N_1490,In_3517,In_3570);
and U1491 (N_1491,In_2746,In_4606);
and U1492 (N_1492,In_3338,In_1047);
xor U1493 (N_1493,In_4872,In_3024);
or U1494 (N_1494,In_4637,In_3556);
nor U1495 (N_1495,In_2905,In_1395);
nor U1496 (N_1496,In_750,In_1280);
and U1497 (N_1497,In_2885,In_2780);
nand U1498 (N_1498,In_2159,In_2789);
nor U1499 (N_1499,In_2368,In_1107);
nor U1500 (N_1500,In_3210,In_4099);
or U1501 (N_1501,In_3197,In_4048);
xor U1502 (N_1502,In_1355,In_536);
nor U1503 (N_1503,In_4582,In_929);
nor U1504 (N_1504,In_4846,In_181);
nor U1505 (N_1505,In_1214,In_3462);
and U1506 (N_1506,In_985,In_5);
or U1507 (N_1507,In_516,In_3070);
nor U1508 (N_1508,In_4929,In_1733);
xor U1509 (N_1509,In_864,In_4987);
nor U1510 (N_1510,In_3633,In_301);
nand U1511 (N_1511,In_3980,In_3382);
xor U1512 (N_1512,In_3202,In_4690);
nor U1513 (N_1513,In_4571,In_3468);
nor U1514 (N_1514,In_769,In_2813);
nor U1515 (N_1515,In_3140,In_1039);
and U1516 (N_1516,In_1517,In_2354);
or U1517 (N_1517,In_272,In_4972);
nor U1518 (N_1518,In_4715,In_3177);
and U1519 (N_1519,In_1424,In_2549);
and U1520 (N_1520,In_1058,In_3523);
and U1521 (N_1521,In_146,In_4035);
nand U1522 (N_1522,In_986,In_1008);
nor U1523 (N_1523,In_2638,In_1991);
nand U1524 (N_1524,In_4558,In_868);
nand U1525 (N_1525,In_2191,In_2238);
nor U1526 (N_1526,In_4308,In_2139);
and U1527 (N_1527,In_4694,In_3533);
xor U1528 (N_1528,In_1777,In_3845);
nor U1529 (N_1529,In_2956,In_1572);
and U1530 (N_1530,In_507,In_3402);
and U1531 (N_1531,In_1577,In_2410);
nand U1532 (N_1532,In_790,In_3690);
xor U1533 (N_1533,In_3740,In_32);
nand U1534 (N_1534,In_2206,In_1348);
xor U1535 (N_1535,In_3722,In_3275);
nand U1536 (N_1536,In_1072,In_4992);
or U1537 (N_1537,In_3372,In_3599);
or U1538 (N_1538,In_4542,In_4685);
and U1539 (N_1539,In_1923,In_3075);
nand U1540 (N_1540,In_4141,In_1829);
and U1541 (N_1541,In_3941,In_3263);
or U1542 (N_1542,In_388,In_1031);
nor U1543 (N_1543,In_4510,In_4465);
and U1544 (N_1544,In_3711,In_30);
nand U1545 (N_1545,In_1334,In_4942);
nor U1546 (N_1546,In_2172,In_3074);
nand U1547 (N_1547,In_1185,In_3166);
and U1548 (N_1548,In_2174,In_2774);
or U1549 (N_1549,In_3109,In_3984);
xnor U1550 (N_1550,In_1032,In_957);
or U1551 (N_1551,In_549,In_2945);
xor U1552 (N_1552,In_3617,In_2926);
and U1553 (N_1553,In_1242,In_184);
nand U1554 (N_1554,In_414,In_3492);
nand U1555 (N_1555,In_427,In_2391);
xnor U1556 (N_1556,In_480,In_3851);
or U1557 (N_1557,In_2583,In_2505);
or U1558 (N_1558,In_1700,In_3551);
or U1559 (N_1559,In_80,In_1759);
or U1560 (N_1560,In_800,In_4075);
and U1561 (N_1561,In_3793,In_4327);
or U1562 (N_1562,In_1693,In_4947);
xor U1563 (N_1563,In_4093,In_4862);
xnor U1564 (N_1564,In_3808,In_4496);
and U1565 (N_1565,In_3453,In_2631);
xnor U1566 (N_1566,In_1887,In_669);
nand U1567 (N_1567,In_3583,In_3774);
xnor U1568 (N_1568,In_3213,In_2145);
or U1569 (N_1569,In_4296,In_1626);
nor U1570 (N_1570,In_1675,In_1071);
and U1571 (N_1571,In_215,In_1281);
and U1572 (N_1572,In_4971,In_4342);
or U1573 (N_1573,In_4969,In_4388);
nand U1574 (N_1574,In_4866,In_1515);
nor U1575 (N_1575,In_1211,In_1875);
xnor U1576 (N_1576,In_618,In_2665);
or U1577 (N_1577,In_2737,In_2810);
nand U1578 (N_1578,In_3718,In_1138);
nand U1579 (N_1579,In_2864,In_551);
xor U1580 (N_1580,In_2046,In_2075);
nor U1581 (N_1581,In_1312,In_1900);
and U1582 (N_1582,In_7,In_2176);
and U1583 (N_1583,In_142,In_2603);
xnor U1584 (N_1584,In_4353,In_4204);
and U1585 (N_1585,In_870,In_94);
xnor U1586 (N_1586,In_492,In_1062);
nor U1587 (N_1587,In_17,In_3133);
and U1588 (N_1588,In_34,In_4071);
and U1589 (N_1589,In_3046,In_1697);
nor U1590 (N_1590,In_4009,In_4250);
nor U1591 (N_1591,In_2154,In_2602);
nor U1592 (N_1592,In_4998,In_4860);
or U1593 (N_1593,In_3424,In_2021);
or U1594 (N_1594,In_2300,In_3460);
or U1595 (N_1595,In_1566,In_4577);
xnor U1596 (N_1596,In_2597,In_1851);
xnor U1597 (N_1597,In_2181,In_1430);
nor U1598 (N_1598,In_3822,In_3629);
or U1599 (N_1599,In_2054,In_1961);
xor U1600 (N_1600,In_1367,In_1558);
xor U1601 (N_1601,In_1580,In_4254);
and U1602 (N_1602,In_2761,In_87);
and U1603 (N_1603,In_121,In_2045);
xnor U1604 (N_1604,In_2542,In_2992);
or U1605 (N_1605,In_1263,In_2661);
or U1606 (N_1606,In_825,In_1445);
xor U1607 (N_1607,In_3249,In_1592);
nor U1608 (N_1608,In_1466,In_3915);
or U1609 (N_1609,In_561,In_36);
and U1610 (N_1610,In_2061,In_1127);
or U1611 (N_1611,In_2787,In_4372);
nand U1612 (N_1612,In_919,In_1191);
and U1613 (N_1613,In_12,In_1046);
and U1614 (N_1614,In_1663,In_4019);
nor U1615 (N_1615,In_4927,In_2554);
nor U1616 (N_1616,In_938,In_265);
xnor U1617 (N_1617,In_3587,In_4635);
xnor U1618 (N_1618,In_1546,In_1356);
or U1619 (N_1619,In_3175,In_169);
nor U1620 (N_1620,In_2161,In_3491);
nor U1621 (N_1621,In_1725,In_1247);
nand U1622 (N_1622,In_1521,In_2404);
xor U1623 (N_1623,In_4779,In_2512);
nor U1624 (N_1624,In_3347,In_1929);
xor U1625 (N_1625,In_4310,In_3270);
nand U1626 (N_1626,In_2605,In_2133);
nor U1627 (N_1627,In_402,In_1463);
xor U1628 (N_1628,In_2856,In_990);
and U1629 (N_1629,In_911,In_2409);
and U1630 (N_1630,In_4605,In_4747);
xor U1631 (N_1631,In_173,In_3574);
or U1632 (N_1632,In_2686,In_370);
and U1633 (N_1633,In_1318,In_4538);
and U1634 (N_1634,In_2051,In_379);
and U1635 (N_1635,In_1554,In_447);
xnor U1636 (N_1636,In_2360,In_2364);
nand U1637 (N_1637,In_4396,In_4886);
and U1638 (N_1638,In_2929,In_4265);
or U1639 (N_1639,In_2250,In_1468);
or U1640 (N_1640,In_1178,In_579);
nor U1641 (N_1641,In_4899,In_916);
nand U1642 (N_1642,In_2523,In_54);
nand U1643 (N_1643,In_3206,In_2101);
nand U1644 (N_1644,In_1243,In_2627);
xor U1645 (N_1645,In_2953,In_3786);
and U1646 (N_1646,In_3379,In_298);
xnor U1647 (N_1647,In_189,In_4454);
and U1648 (N_1648,In_3951,In_3969);
nor U1649 (N_1649,In_3487,In_765);
nor U1650 (N_1650,In_2297,In_2654);
and U1651 (N_1651,In_4528,In_799);
or U1652 (N_1652,In_1872,In_1569);
nor U1653 (N_1653,In_730,In_3836);
or U1654 (N_1654,In_1857,In_3577);
xnor U1655 (N_1655,In_1183,In_1212);
and U1656 (N_1656,In_2566,In_2455);
nand U1657 (N_1657,In_3448,In_713);
nand U1658 (N_1658,In_2788,In_3767);
nand U1659 (N_1659,In_4471,In_2350);
nor U1660 (N_1660,In_2189,In_3626);
and U1661 (N_1661,In_3892,In_3248);
xor U1662 (N_1662,In_3691,In_3971);
or U1663 (N_1663,In_3918,In_2808);
nand U1664 (N_1664,In_4135,In_4290);
nand U1665 (N_1665,In_4447,In_1249);
nor U1666 (N_1666,In_3904,In_4272);
nor U1667 (N_1667,In_4096,In_759);
and U1668 (N_1668,In_2282,In_4665);
and U1669 (N_1669,In_4021,In_2858);
or U1670 (N_1670,In_2621,In_20);
nor U1671 (N_1671,In_2985,In_4658);
xor U1672 (N_1672,In_4316,In_1607);
or U1673 (N_1673,In_205,In_3139);
nor U1674 (N_1674,In_2983,In_3457);
or U1675 (N_1675,In_481,In_1068);
xnor U1676 (N_1676,In_937,In_4404);
or U1677 (N_1677,In_580,In_1819);
xnor U1678 (N_1678,In_3313,In_1478);
nor U1679 (N_1679,In_156,In_4695);
and U1680 (N_1680,In_1724,In_2433);
nand U1681 (N_1681,In_4352,In_2526);
nor U1682 (N_1682,In_746,In_4916);
or U1683 (N_1683,In_1262,In_191);
or U1684 (N_1684,In_3749,In_365);
xnor U1685 (N_1685,In_4520,In_3797);
and U1686 (N_1686,In_2875,In_2569);
nor U1687 (N_1687,In_4215,In_3888);
nand U1688 (N_1688,In_975,In_3351);
xnor U1689 (N_1689,In_4664,In_3136);
or U1690 (N_1690,In_2085,In_531);
xor U1691 (N_1691,In_498,In_2972);
and U1692 (N_1692,In_2939,In_3567);
nor U1693 (N_1693,In_91,In_1323);
and U1694 (N_1694,In_4881,In_323);
xnor U1695 (N_1695,In_4162,In_3322);
or U1696 (N_1696,In_3392,In_2498);
and U1697 (N_1697,In_245,In_834);
xor U1698 (N_1698,In_1369,In_2128);
and U1699 (N_1699,In_4518,In_4418);
nand U1700 (N_1700,In_4390,In_658);
nor U1701 (N_1701,In_613,In_2965);
nand U1702 (N_1702,In_2185,In_4050);
and U1703 (N_1703,In_3422,In_4154);
xor U1704 (N_1704,In_4475,In_51);
nor U1705 (N_1705,In_93,In_3364);
or U1706 (N_1706,In_3540,In_1018);
or U1707 (N_1707,In_3135,In_3719);
and U1708 (N_1708,In_1054,In_152);
and U1709 (N_1709,In_1736,In_4887);
nand U1710 (N_1710,In_3221,In_344);
or U1711 (N_1711,In_3239,In_4802);
xnor U1712 (N_1712,In_3703,In_3277);
nand U1713 (N_1713,In_2760,In_3160);
xnor U1714 (N_1714,In_4417,In_900);
xnor U1715 (N_1715,In_1381,In_2169);
or U1716 (N_1716,In_3536,In_983);
xnor U1717 (N_1717,In_2544,In_4003);
xnor U1718 (N_1718,In_3607,In_2342);
or U1719 (N_1719,In_1016,In_4195);
nor U1720 (N_1720,In_1565,In_2724);
nor U1721 (N_1721,In_4345,In_3201);
nor U1722 (N_1722,In_4631,In_3769);
xnor U1723 (N_1723,In_218,In_314);
or U1724 (N_1724,In_4016,In_4750);
nor U1725 (N_1725,In_4894,In_3265);
or U1726 (N_1726,In_4773,In_1471);
xor U1727 (N_1727,In_3725,In_2918);
or U1728 (N_1728,In_1025,In_1788);
and U1729 (N_1729,In_4175,In_1252);
or U1730 (N_1730,In_668,In_3561);
and U1731 (N_1731,In_4830,In_1888);
nand U1732 (N_1732,In_4911,In_3352);
or U1733 (N_1733,In_3558,In_2802);
or U1734 (N_1734,In_1274,In_1491);
and U1735 (N_1735,In_4315,In_4196);
and U1736 (N_1736,In_3203,In_1503);
or U1737 (N_1737,In_4979,In_166);
nor U1738 (N_1738,In_4624,In_4248);
or U1739 (N_1739,In_721,In_3741);
nand U1740 (N_1740,In_2824,In_1778);
and U1741 (N_1741,In_4121,In_1708);
nand U1742 (N_1742,In_3033,In_4700);
and U1743 (N_1743,In_2402,In_3303);
nor U1744 (N_1744,In_1581,In_3430);
nand U1745 (N_1745,In_4626,In_1231);
nor U1746 (N_1746,In_3771,In_3054);
nand U1747 (N_1747,In_2733,In_3868);
nand U1748 (N_1748,In_1594,In_1769);
or U1749 (N_1749,In_1370,In_4184);
or U1750 (N_1750,In_988,In_1758);
xnor U1751 (N_1751,In_23,In_1790);
or U1752 (N_1752,In_198,In_889);
and U1753 (N_1753,In_4153,In_2611);
nand U1754 (N_1754,In_2398,In_2148);
nand U1755 (N_1755,In_4945,In_65);
and U1756 (N_1756,In_129,In_132);
and U1757 (N_1757,In_2351,In_2950);
and U1758 (N_1758,In_226,In_3734);
xnor U1759 (N_1759,In_4398,In_970);
nand U1760 (N_1760,In_2258,In_207);
nor U1761 (N_1761,In_2618,In_552);
nand U1762 (N_1762,In_3182,In_895);
and U1763 (N_1763,In_3423,In_3262);
nor U1764 (N_1764,In_2598,In_1550);
nand U1765 (N_1765,In_762,In_1473);
nor U1766 (N_1766,In_266,In_584);
xor U1767 (N_1767,In_3048,In_3049);
nor U1768 (N_1768,In_811,In_3810);
nand U1769 (N_1769,In_3172,In_2347);
nand U1770 (N_1770,In_3065,In_3485);
or U1771 (N_1771,In_2785,In_2834);
or U1772 (N_1772,In_1265,In_4491);
xor U1773 (N_1773,In_4579,In_2609);
and U1774 (N_1774,In_2790,In_3658);
nor U1775 (N_1775,In_4659,In_117);
xor U1776 (N_1776,In_3354,In_4211);
xor U1777 (N_1777,In_2432,In_1610);
nand U1778 (N_1778,In_4724,In_3273);
nor U1779 (N_1779,In_3684,In_2343);
xnor U1780 (N_1780,In_3882,In_1827);
xor U1781 (N_1781,In_4305,In_1504);
and U1782 (N_1782,In_2530,In_2466);
xnor U1783 (N_1783,In_2108,In_188);
nand U1784 (N_1784,In_1599,In_1413);
xnor U1785 (N_1785,In_965,In_1165);
or U1786 (N_1786,In_902,In_1975);
and U1787 (N_1787,In_4335,In_105);
or U1788 (N_1788,In_3952,In_2809);
nor U1789 (N_1789,In_2596,In_3863);
nor U1790 (N_1790,In_1162,In_200);
and U1791 (N_1791,In_2580,In_2806);
xor U1792 (N_1792,In_4775,In_2470);
or U1793 (N_1793,In_4829,In_968);
or U1794 (N_1794,In_2323,In_674);
xor U1795 (N_1795,In_842,In_3439);
or U1796 (N_1796,In_525,In_1254);
nand U1797 (N_1797,In_1022,In_4010);
nor U1798 (N_1798,In_4882,In_4400);
nand U1799 (N_1799,In_3911,In_4900);
xnor U1800 (N_1800,In_594,In_4612);
nand U1801 (N_1801,In_1332,In_743);
nor U1802 (N_1802,In_795,In_2234);
nor U1803 (N_1803,In_4262,In_1177);
xnor U1804 (N_1804,In_3788,In_4512);
nand U1805 (N_1805,In_1665,In_466);
nor U1806 (N_1806,In_1692,In_3466);
nand U1807 (N_1807,In_4851,In_2412);
and U1808 (N_1808,In_1815,In_3195);
and U1809 (N_1809,In_459,In_562);
xnor U1810 (N_1810,In_586,In_1925);
xor U1811 (N_1811,In_3185,In_677);
or U1812 (N_1812,In_2873,In_3399);
or U1813 (N_1813,In_4869,In_2719);
nor U1814 (N_1814,In_4043,In_136);
nor U1815 (N_1815,In_1158,In_1904);
or U1816 (N_1816,In_442,In_2453);
nor U1817 (N_1817,In_3700,In_1579);
nor U1818 (N_1818,In_4919,In_2624);
nand U1819 (N_1819,In_3760,In_1131);
xor U1820 (N_1820,In_1540,In_3398);
nor U1821 (N_1821,In_1619,In_4232);
nand U1822 (N_1822,In_2568,In_2177);
or U1823 (N_1823,In_4251,In_966);
nand U1824 (N_1824,In_1228,In_4629);
or U1825 (N_1825,In_1506,In_3733);
or U1826 (N_1826,In_1221,In_4857);
and U1827 (N_1827,In_116,In_1489);
or U1828 (N_1828,In_1547,In_3500);
nand U1829 (N_1829,In_2635,In_4213);
or U1830 (N_1830,In_2502,In_2639);
nand U1831 (N_1831,In_3747,In_4847);
and U1832 (N_1832,In_1213,In_1389);
nand U1833 (N_1833,In_3665,In_3648);
xor U1834 (N_1834,In_3876,In_4130);
nand U1835 (N_1835,In_3250,In_1798);
xnor U1836 (N_1836,In_1149,In_3942);
and U1837 (N_1837,In_3645,In_490);
or U1838 (N_1838,In_3419,In_140);
and U1839 (N_1839,In_3464,In_50);
nor U1840 (N_1840,In_3429,In_4181);
nand U1841 (N_1841,In_192,In_3729);
xor U1842 (N_1842,In_3717,In_342);
xor U1843 (N_1843,In_1347,In_4375);
or U1844 (N_1844,In_2891,In_2248);
or U1845 (N_1845,In_2010,In_4458);
and U1846 (N_1846,In_3687,In_3944);
or U1847 (N_1847,In_2027,In_1623);
or U1848 (N_1848,In_2697,In_2648);
nor U1849 (N_1849,In_544,In_2584);
nor U1850 (N_1850,In_1485,In_1669);
xor U1851 (N_1851,In_2381,In_410);
xor U1852 (N_1852,In_1192,In_284);
nand U1853 (N_1853,In_952,In_1261);
nor U1854 (N_1854,In_383,In_440);
or U1855 (N_1855,In_4436,In_1421);
and U1856 (N_1856,In_2425,In_113);
and U1857 (N_1857,In_2482,In_703);
nand U1858 (N_1858,In_3115,In_1401);
or U1859 (N_1859,In_1052,In_3304);
and U1860 (N_1860,In_1775,In_178);
xnor U1861 (N_1861,In_2370,In_1582);
nor U1862 (N_1862,In_2014,In_777);
and U1863 (N_1863,In_2311,In_3605);
and U1864 (N_1864,In_2302,In_1761);
nor U1865 (N_1865,In_4386,In_2278);
or U1866 (N_1866,In_4177,In_3636);
xnor U1867 (N_1867,In_4575,In_804);
xor U1868 (N_1868,In_3481,In_2770);
nand U1869 (N_1869,In_285,In_1853);
xnor U1870 (N_1870,In_2000,In_3699);
and U1871 (N_1871,In_1487,In_1602);
xor U1872 (N_1872,In_2467,In_1861);
nor U1873 (N_1873,In_4403,In_699);
xnor U1874 (N_1874,In_186,In_2077);
nand U1875 (N_1875,In_4108,In_2525);
and U1876 (N_1876,In_3522,In_1357);
and U1877 (N_1877,In_4767,In_1994);
xnor U1878 (N_1878,In_3563,In_76);
xor U1879 (N_1879,In_299,In_1822);
or U1880 (N_1880,In_1208,In_3511);
xnor U1881 (N_1881,In_4954,In_1774);
or U1882 (N_1882,In_3241,In_360);
nand U1883 (N_1883,In_3976,In_4037);
xor U1884 (N_1884,In_112,In_4763);
and U1885 (N_1885,In_1705,In_3090);
nand U1886 (N_1886,In_2867,In_2674);
and U1887 (N_1887,In_3011,In_2619);
or U1888 (N_1888,In_2004,In_1293);
xor U1889 (N_1889,In_768,In_1393);
nor U1890 (N_1890,In_4549,In_609);
nand U1891 (N_1891,In_4536,In_1472);
and U1892 (N_1892,In_473,In_4974);
nor U1893 (N_1893,In_380,In_1614);
nand U1894 (N_1894,In_565,In_853);
xnor U1895 (N_1895,In_3028,In_2721);
xor U1896 (N_1896,In_2932,In_164);
or U1897 (N_1897,In_2685,In_871);
nand U1898 (N_1898,In_232,In_1084);
or U1899 (N_1899,In_3431,In_2756);
or U1900 (N_1900,In_4370,In_4309);
and U1901 (N_1901,In_1246,In_500);
nor U1902 (N_1902,In_662,In_1237);
xnor U1903 (N_1903,In_3114,In_4620);
nand U1904 (N_1904,In_446,In_2400);
and U1905 (N_1905,In_1045,In_2211);
and U1906 (N_1906,In_4788,In_705);
or U1907 (N_1907,In_4227,In_1617);
nor U1908 (N_1908,In_4997,In_697);
or U1909 (N_1909,In_4646,In_1776);
or U1910 (N_1910,In_4369,In_4159);
xor U1911 (N_1911,In_736,In_2758);
and U1912 (N_1912,In_4946,In_2622);
xnor U1913 (N_1913,In_2947,In_4878);
or U1914 (N_1914,In_2954,In_1919);
nor U1915 (N_1915,In_3548,In_1909);
nand U1916 (N_1916,In_3484,In_4445);
xor U1917 (N_1917,In_2720,In_1012);
xnor U1918 (N_1918,In_3936,In_2751);
nor U1919 (N_1919,In_46,In_225);
or U1920 (N_1920,In_3962,In_789);
xor U1921 (N_1921,In_2702,In_4523);
and U1922 (N_1922,In_2190,In_2971);
nand U1923 (N_1923,In_1028,In_2844);
and U1924 (N_1924,In_168,In_4397);
nand U1925 (N_1925,In_3527,In_891);
or U1926 (N_1926,In_3537,In_1897);
or U1927 (N_1927,In_3887,In_1250);
or U1928 (N_1928,In_4776,In_2089);
nor U1929 (N_1929,In_3816,In_1126);
and U1930 (N_1930,In_3995,In_3975);
nor U1931 (N_1931,In_3739,In_3328);
nor U1932 (N_1932,In_704,In_873);
xor U1933 (N_1933,In_271,In_441);
and U1934 (N_1934,In_737,In_3121);
and U1935 (N_1935,In_3652,In_1490);
nand U1936 (N_1936,In_2055,In_2634);
xor U1937 (N_1937,In_931,In_3493);
nor U1938 (N_1938,In_4616,In_1454);
nor U1939 (N_1939,In_3796,In_2778);
nor U1940 (N_1940,In_3860,In_3440);
or U1941 (N_1941,In_1642,In_903);
nor U1942 (N_1942,In_1898,In_3110);
nand U1943 (N_1943,In_1399,In_1646);
or U1944 (N_1944,In_3798,In_672);
xor U1945 (N_1945,In_4230,In_3602);
xor U1946 (N_1946,In_4999,In_1227);
nor U1947 (N_1947,In_3815,In_372);
nand U1948 (N_1948,In_4477,In_4402);
nand U1949 (N_1949,In_3300,In_4326);
or U1950 (N_1950,In_3694,In_1796);
nand U1951 (N_1951,In_2791,In_4645);
and U1952 (N_1952,In_4046,In_2850);
and U1953 (N_1953,In_2593,In_4600);
and U1954 (N_1954,In_1625,In_935);
xnor U1955 (N_1955,In_4452,In_3153);
xnor U1956 (N_1956,In_475,In_3022);
xor U1957 (N_1957,In_597,In_874);
xnor U1958 (N_1958,In_2679,In_1834);
nor U1959 (N_1959,In_4749,In_1431);
nand U1960 (N_1960,In_1836,In_604);
or U1961 (N_1961,In_2919,In_3276);
nor U1962 (N_1962,In_887,In_3922);
xor U1963 (N_1963,In_4321,In_1306);
xnor U1964 (N_1964,In_4266,In_1108);
or U1965 (N_1965,In_149,In_2270);
nand U1966 (N_1966,In_9,In_2363);
nand U1967 (N_1967,In_4221,In_4219);
nand U1968 (N_1968,In_1781,In_2259);
or U1969 (N_1969,In_4566,In_1289);
and U1970 (N_1970,In_3521,In_1816);
and U1971 (N_1971,In_4222,In_4556);
nor U1972 (N_1972,In_2700,In_3378);
or U1973 (N_1973,In_998,In_890);
or U1974 (N_1974,In_3391,In_3688);
and U1975 (N_1975,In_224,In_4483);
or U1976 (N_1976,In_4720,In_2076);
and U1977 (N_1977,In_1034,In_3073);
xor U1978 (N_1978,In_273,In_624);
and U1979 (N_1979,In_1528,In_4113);
nor U1980 (N_1980,In_2303,In_317);
or U1981 (N_1981,In_109,In_1981);
or U1982 (N_1982,In_2118,In_3565);
nor U1983 (N_1983,In_2299,In_3170);
and U1984 (N_1984,In_1330,In_3145);
or U1985 (N_1985,In_3178,In_2777);
and U1986 (N_1986,In_2290,In_4769);
or U1987 (N_1987,In_1187,In_26);
nand U1988 (N_1988,In_3909,In_4675);
xor U1989 (N_1989,In_1974,In_974);
or U1990 (N_1990,In_1833,In_636);
nor U1991 (N_1991,In_2538,In_3894);
or U1992 (N_1992,In_2736,In_511);
nand U1993 (N_1993,In_1927,In_3180);
nor U1994 (N_1994,In_641,In_2553);
or U1995 (N_1995,In_412,In_3327);
nor U1996 (N_1996,In_1481,In_3432);
nor U1997 (N_1997,In_3027,In_4609);
or U1998 (N_1998,In_4039,In_1202);
nand U1999 (N_1999,In_4317,In_49);
nor U2000 (N_2000,In_513,In_4158);
and U2001 (N_2001,In_4020,In_1780);
nand U2002 (N_2002,In_780,In_4076);
nor U2003 (N_2003,In_1709,In_3189);
nand U2004 (N_2004,In_2845,In_2607);
nor U2005 (N_2005,In_673,In_3659);
or U2006 (N_2006,In_3813,In_1964);
nand U2007 (N_2007,In_1189,In_1069);
and U2008 (N_2008,In_3938,In_71);
or U2009 (N_2009,In_423,In_1477);
nand U2010 (N_2010,In_1216,In_2192);
xor U2011 (N_2011,In_4144,In_2341);
and U2012 (N_2012,In_1404,In_3840);
xnor U2013 (N_2013,In_2040,In_3554);
and U2014 (N_2014,In_671,In_3279);
and U2015 (N_2015,In_313,In_4780);
or U2016 (N_2016,In_4668,In_1150);
xnor U2017 (N_2017,In_3974,In_3302);
nand U2018 (N_2018,In_2110,In_3297);
xor U2019 (N_2019,In_4543,In_4291);
nor U2020 (N_2020,In_1993,In_3168);
xnor U2021 (N_2021,In_3666,In_4661);
or U2022 (N_2022,In_4937,In_606);
or U2023 (N_2023,In_993,In_1414);
nor U2024 (N_2024,In_4457,In_180);
or U2025 (N_2025,In_881,In_2435);
and U2026 (N_2026,In_585,In_3259);
nor U2027 (N_2027,In_2587,In_2450);
xnor U2028 (N_2028,In_505,In_2245);
nand U2029 (N_2029,In_2870,In_4583);
or U2030 (N_2030,In_4705,In_4722);
and U2031 (N_2031,In_101,In_3954);
nand U2032 (N_2032,In_2667,In_1830);
or U2033 (N_2033,In_3331,In_236);
nand U2034 (N_2034,In_694,In_2960);
nand U2035 (N_2035,In_3287,In_819);
xnor U2036 (N_2036,In_444,In_3157);
xor U2037 (N_2037,In_2881,In_1953);
nor U2038 (N_2038,In_4100,In_4896);
nor U2039 (N_2039,In_4726,In_3507);
nor U2040 (N_2040,In_4811,In_2988);
nand U2041 (N_2041,In_2293,In_849);
or U2042 (N_2042,In_18,In_2487);
xnor U2043 (N_2043,In_431,In_2253);
xnor U2044 (N_2044,In_3267,In_2147);
and U2045 (N_2045,In_2759,In_696);
and U2046 (N_2046,In_3486,In_4613);
nor U2047 (N_2047,In_3884,In_3664);
nor U2048 (N_2048,In_2689,In_2086);
or U2049 (N_2049,In_3498,In_2216);
nand U2050 (N_2050,In_1691,In_2536);
xor U2051 (N_2051,In_4440,In_1238);
nor U2052 (N_2052,In_2863,In_190);
nand U2053 (N_2053,In_3329,In_494);
and U2054 (N_2054,In_4104,In_1593);
or U2055 (N_2055,In_3870,In_4702);
and U2056 (N_2056,In_3847,In_1229);
nand U2057 (N_2057,In_1273,In_1760);
nor U2058 (N_2058,In_1361,In_4982);
nand U2059 (N_2059,In_2437,In_3643);
nor U2060 (N_2060,In_1590,In_409);
or U2061 (N_2061,In_4774,In_4413);
and U2062 (N_2062,In_2358,In_3497);
nand U2063 (N_2063,In_223,In_2980);
nand U2064 (N_2064,In_691,In_3874);
xnor U2065 (N_2065,In_4511,In_623);
nor U2066 (N_2066,In_1204,In_311);
xor U2067 (N_2067,In_4237,In_2043);
and U2068 (N_2068,In_237,In_1075);
xnor U2069 (N_2069,In_951,In_2112);
and U2070 (N_2070,In_3290,In_4753);
or U2071 (N_2071,In_1329,In_1749);
and U2072 (N_2072,In_1631,In_2854);
nand U2073 (N_2073,In_2974,In_4078);
or U2074 (N_2074,In_3260,In_4940);
xnor U2075 (N_2075,In_1398,In_4800);
xor U2076 (N_2076,In_4339,In_3336);
and U2077 (N_2077,In_1976,In_2167);
nor U2078 (N_2078,In_850,In_695);
nor U2079 (N_2079,In_4462,In_3041);
and U2080 (N_2080,In_280,In_4782);
xor U2081 (N_2081,In_3009,In_1448);
or U2082 (N_2082,In_3534,In_2454);
xor U2083 (N_2083,In_3835,In_3535);
nand U2084 (N_2084,In_1756,In_78);
xor U2085 (N_2085,In_1545,In_2231);
nor U2086 (N_2086,In_1085,In_3625);
or U2087 (N_2087,In_3818,In_3125);
nor U2088 (N_2088,In_556,In_1321);
nand U2089 (N_2089,In_4066,In_3506);
or U2090 (N_2090,In_593,In_3743);
and U2091 (N_2091,In_4349,In_211);
or U2092 (N_2092,In_2367,In_2217);
xor U2093 (N_2093,In_3333,In_1562);
or U2094 (N_2094,In_508,In_3805);
nor U2095 (N_2095,In_3343,In_1615);
xor U2096 (N_2096,In_685,In_270);
nand U2097 (N_2097,In_4470,In_3005);
or U2098 (N_2098,In_2194,In_4347);
nand U2099 (N_2099,In_3732,In_3257);
xnor U2100 (N_2100,In_1586,In_297);
nor U2101 (N_2101,In_4053,In_96);
and U2102 (N_2102,In_83,In_1017);
or U2103 (N_2103,In_2921,In_2901);
xnor U2104 (N_2104,In_1001,In_2184);
nor U2105 (N_2105,In_3094,In_1428);
nor U2106 (N_2106,In_4877,In_2292);
or U2107 (N_2107,In_2887,In_3061);
xor U2108 (N_2108,In_3078,In_1505);
nand U2109 (N_2109,In_589,In_1704);
or U2110 (N_2110,In_1688,In_4628);
nor U2111 (N_2111,In_102,In_332);
or U2112 (N_2112,In_2610,In_4123);
nand U2113 (N_2113,In_2097,In_1041);
and U2114 (N_2114,In_1239,In_1785);
and U2115 (N_2115,In_2322,In_1437);
xnor U2116 (N_2116,In_4541,In_1944);
or U2117 (N_2117,In_3724,In_1922);
nor U2118 (N_2118,In_3227,In_4683);
nor U2119 (N_2119,In_2662,In_540);
or U2120 (N_2120,In_4591,In_2820);
nand U2121 (N_2121,In_3031,In_2235);
xnor U2122 (N_2122,In_3155,In_1648);
nand U2123 (N_2123,In_2946,In_1723);
or U2124 (N_2124,In_1573,In_2753);
or U2125 (N_2125,In_555,In_59);
nand U2126 (N_2126,In_3931,In_222);
nand U2127 (N_2127,In_635,In_2422);
nand U2128 (N_2128,In_612,In_3968);
and U2129 (N_2129,In_305,In_2734);
or U2130 (N_2130,In_4555,In_1139);
or U2131 (N_2131,In_848,In_413);
xnor U2132 (N_2132,In_3420,In_468);
xnor U2133 (N_2133,In_469,In_2540);
nor U2134 (N_2134,In_4366,In_4808);
nor U2135 (N_2135,In_4414,In_1196);
nand U2136 (N_2136,In_1735,In_1446);
xor U2137 (N_2137,In_316,In_1451);
xnor U2138 (N_2138,In_915,In_3923);
xor U2139 (N_2139,In_2681,In_2576);
nor U2140 (N_2140,In_2255,In_56);
xnor U2141 (N_2141,In_2880,In_145);
or U2142 (N_2142,In_1453,In_2716);
and U2143 (N_2143,In_3152,In_514);
nand U2144 (N_2144,In_3538,In_2325);
nand U2145 (N_2145,In_1412,In_1996);
or U2146 (N_2146,In_2312,In_1303);
and U2147 (N_2147,In_4596,In_242);
nor U2148 (N_2148,In_1006,In_1343);
or U2149 (N_2149,In_2750,In_2252);
or U2150 (N_2150,In_3943,In_809);
nand U2151 (N_2151,In_4873,In_4242);
nand U2152 (N_2152,In_1773,In_3830);
or U2153 (N_2153,In_3628,In_3319);
nand U2154 (N_2154,In_1728,In_3437);
and U2155 (N_2155,In_3212,In_2633);
xor U2156 (N_2156,In_1908,In_1497);
and U2157 (N_2157,In_45,In_374);
and U2158 (N_2158,In_2784,In_4169);
or U2159 (N_2159,In_700,In_3748);
and U2160 (N_2160,In_927,In_2163);
or U2161 (N_2161,In_3034,In_4025);
nor U2162 (N_2162,In_1745,In_2463);
nor U2163 (N_2163,In_3903,In_1793);
nor U2164 (N_2164,In_3898,In_28);
nand U2165 (N_2165,In_3755,In_3575);
or U2166 (N_2166,In_4990,In_3879);
xnor U2167 (N_2167,In_2093,In_6);
xor U2168 (N_2168,In_2414,In_510);
and U2169 (N_2169,In_1320,In_1576);
nor U2170 (N_2170,In_707,In_4701);
nand U2171 (N_2171,In_1608,In_2876);
xor U2172 (N_2172,In_4286,In_3358);
or U2173 (N_2173,In_3706,In_4133);
or U2174 (N_2174,In_4423,In_1680);
xnor U2175 (N_2175,In_150,In_2623);
xor U2176 (N_2176,In_4717,In_3893);
xnor U2177 (N_2177,In_4117,In_4904);
and U2178 (N_2178,In_3039,In_3807);
nand U2179 (N_2179,In_3455,In_1563);
nand U2180 (N_2180,In_3877,In_1632);
nor U2181 (N_2181,In_3624,In_1676);
nor U2182 (N_2182,In_2795,In_3080);
or U2183 (N_2183,In_529,In_4744);
and U2184 (N_2184,In_4148,In_3580);
nand U2185 (N_2185,In_3872,In_4914);
or U2186 (N_2186,In_2420,In_4444);
xor U2187 (N_2187,In_1863,In_4156);
nor U2188 (N_2188,In_4764,In_1706);
xnor U2189 (N_2189,In_2441,In_279);
nor U2190 (N_2190,In_945,In_1962);
nand U2191 (N_2191,In_2715,In_835);
nor U2192 (N_2192,In_1145,In_2100);
xor U2193 (N_2193,In_1488,In_4140);
nand U2194 (N_2194,In_1106,In_1123);
nand U2195 (N_2195,In_4446,In_1518);
nand U2196 (N_2196,In_4289,In_1859);
nand U2197 (N_2197,In_3661,In_252);
nand U2198 (N_2198,In_1942,In_4147);
or U2199 (N_2199,In_1418,In_1181);
or U2200 (N_2200,In_3045,In_2763);
nand U2201 (N_2201,In_2026,In_1539);
nand U2202 (N_2202,In_1532,In_3282);
or U2203 (N_2203,In_1559,In_2615);
xnor U2204 (N_2204,In_3435,In_267);
nor U2205 (N_2205,In_2745,In_1764);
nor U2206 (N_2206,In_2578,In_3627);
nor U2207 (N_2207,In_3417,In_4092);
nor U2208 (N_2208,In_3317,In_3965);
nand U2209 (N_2209,In_2460,In_4029);
and U2210 (N_2210,In_2330,In_2418);
nor U2211 (N_2211,In_130,In_3735);
or U2212 (N_2212,In_4187,In_854);
xor U2213 (N_2213,In_2126,In_2332);
nor U2214 (N_2214,In_4234,In_2706);
nand U2215 (N_2215,In_770,In_2166);
nor U2216 (N_2216,In_4273,In_4112);
and U2217 (N_2217,In_3120,In_3844);
xor U2218 (N_2218,In_4203,In_1682);
and U2219 (N_2219,In_806,In_3459);
or U2220 (N_2220,In_3451,In_689);
nor U2221 (N_2221,In_953,In_909);
or U2222 (N_2222,In_3867,In_4097);
and U2223 (N_2223,In_3963,In_4706);
or U2224 (N_2224,In_1694,In_4322);
nand U2225 (N_2225,In_4034,In_2335);
and U2226 (N_2226,In_128,In_4789);
or U2227 (N_2227,In_1835,In_684);
and U2228 (N_2228,In_2392,In_4559);
xor U2229 (N_2229,In_3369,In_1080);
or U2230 (N_2230,In_2131,In_4619);
nor U2231 (N_2231,In_1501,In_670);
xor U2232 (N_2232,In_3159,In_3268);
nor U2233 (N_2233,In_104,In_3781);
or U2234 (N_2234,In_2316,In_1578);
or U2235 (N_2235,In_4442,In_886);
and U2236 (N_2236,In_274,In_3142);
nand U2237 (N_2237,In_4760,In_3368);
and U2238 (N_2238,In_89,In_1294);
nand U2239 (N_2239,In_2436,In_1801);
nor U2240 (N_2240,In_1065,In_946);
nand U2241 (N_2241,In_3296,In_4732);
and U2242 (N_2242,In_4167,In_2399);
xor U2243 (N_2243,In_4754,In_2090);
xor U2244 (N_2244,In_1493,In_1349);
nor U2245 (N_2245,In_3123,In_1442);
nand U2246 (N_2246,In_241,In_1512);
or U2247 (N_2247,In_2393,In_1802);
nor U2248 (N_2248,In_4818,In_633);
or U2249 (N_2249,In_3930,In_4660);
xnor U2250 (N_2250,In_1561,In_4975);
and U2251 (N_2251,In_4119,In_1901);
and U2252 (N_2252,In_3298,In_1427);
nor U2253 (N_2253,In_467,In_4807);
xnor U2254 (N_2254,In_3271,In_1362);
xor U2255 (N_2255,In_4292,In_1283);
nand U2256 (N_2256,In_4854,In_3091);
nand U2257 (N_2257,In_1040,In_4082);
and U2258 (N_2258,In_3546,In_2136);
xor U2259 (N_2259,In_2557,In_2643);
xor U2260 (N_2260,In_4371,In_435);
and U2261 (N_2261,In_2,In_2762);
or U2262 (N_2262,In_1236,In_2741);
nand U2263 (N_2263,In_214,In_2157);
nor U2264 (N_2264,In_4584,In_445);
nand U2265 (N_2265,In_1118,In_3773);
or U2266 (N_2266,In_3878,In_133);
and U2267 (N_2267,In_1255,In_716);
nor U2268 (N_2268,In_1555,In_2911);
nand U2269 (N_2269,In_822,In_3188);
nor U2270 (N_2270,In_2407,In_4716);
nor U2271 (N_2271,In_2723,In_1711);
and U2272 (N_2272,In_2334,In_651);
nor U2273 (N_2273,In_1282,In_4655);
and U2274 (N_2274,In_3089,In_3231);
or U2275 (N_2275,In_4778,In_2573);
nand U2276 (N_2276,In_2109,In_2283);
xnor U2277 (N_2277,In_368,In_792);
xnor U2278 (N_2278,In_137,In_523);
nor U2279 (N_2279,In_521,In_2294);
xnor U2280 (N_2280,In_2705,In_4274);
xnor U2281 (N_2281,In_3198,In_114);
nand U2282 (N_2282,In_3606,In_727);
nand U2283 (N_2283,In_1416,In_2653);
and U2284 (N_2284,In_4086,In_4427);
xnor U2285 (N_2285,In_3218,In_2575);
xnor U2286 (N_2286,In_1894,In_4428);
and U2287 (N_2287,In_3337,In_1885);
or U2288 (N_2288,In_1121,In_2585);
nor U2289 (N_2289,In_4604,In_2308);
nand U2290 (N_2290,In_4627,In_1583);
or U2291 (N_2291,In_2180,In_1174);
nor U2292 (N_2292,In_2033,In_4680);
or U2293 (N_2293,In_4258,In_322);
nand U2294 (N_2294,In_2900,In_391);
nor U2295 (N_2295,In_1679,In_2491);
or U2296 (N_2296,In_2539,In_425);
nand U2297 (N_2297,In_3038,In_3529);
or U2298 (N_2298,In_2468,In_576);
nor U2299 (N_2299,In_1620,In_1806);
and U2300 (N_2300,In_4936,In_1167);
and U2301 (N_2301,In_4925,In_3754);
nor U2302 (N_2302,In_542,In_1038);
and U2303 (N_2303,In_4378,In_95);
nand U2304 (N_2304,In_4239,In_4022);
and U2305 (N_2305,In_2123,In_2315);
xnor U2306 (N_2306,In_3726,In_947);
xor U2307 (N_2307,In_2658,In_982);
nor U2308 (N_2308,In_1125,In_1882);
nand U2309 (N_2309,In_2970,In_398);
or U2310 (N_2310,In_2807,In_2212);
and U2311 (N_2311,In_385,In_1027);
or U2312 (N_2312,In_2833,In_3604);
xor U2313 (N_2313,In_4077,In_3147);
and U2314 (N_2314,In_3449,In_3205);
and U2315 (N_2315,In_2318,In_4567);
xor U2316 (N_2316,In_1589,In_4368);
nand U2317 (N_2317,In_1869,In_4537);
and U2318 (N_2318,In_4771,In_3559);
xor U2319 (N_2319,In_3285,In_2868);
xnor U2320 (N_2320,In_2125,In_2267);
xnor U2321 (N_2321,In_499,In_2767);
xor U2322 (N_2322,In_3216,In_4594);
xor U2323 (N_2323,In_3541,In_4393);
xor U2324 (N_2324,In_4056,In_2183);
and U2325 (N_2325,In_355,In_2830);
and U2326 (N_2326,In_1917,In_3708);
nor U2327 (N_2327,In_2057,In_4687);
and U2328 (N_2328,In_86,In_2013);
nand U2329 (N_2329,In_933,In_1670);
nor U2330 (N_2330,In_248,In_3508);
nor U2331 (N_2331,In_4684,In_2997);
xor U2332 (N_2332,In_3335,In_4603);
nor U2333 (N_2333,In_3342,In_163);
and U2334 (N_2334,In_1952,In_1386);
nor U2335 (N_2335,In_626,In_4745);
xnor U2336 (N_2336,In_3824,In_2896);
nor U2337 (N_2337,In_1656,In_4376);
xnor U2338 (N_2338,In_3843,In_3610);
and U2339 (N_2339,In_4481,In_4985);
xor U2340 (N_2340,In_855,In_404);
and U2341 (N_2341,In_2007,In_2415);
nand U2342 (N_2342,In_3715,In_4509);
or U2343 (N_2343,In_918,In_3470);
nand U2344 (N_2344,In_722,In_436);
nor U2345 (N_2345,In_1935,In_3723);
and U2346 (N_2346,In_528,In_1995);
or U2347 (N_2347,In_578,In_3543);
or U2348 (N_2348,In_329,In_4068);
nand U2349 (N_2349,In_257,In_4525);
xor U2350 (N_2350,In_1992,In_4088);
and U2351 (N_2351,In_3179,In_3174);
nand U2352 (N_2352,In_1538,In_1651);
or U2353 (N_2353,In_1879,In_2141);
nor U2354 (N_2354,In_1636,In_3289);
or U2355 (N_2355,In_2877,In_4666);
nand U2356 (N_2356,In_3105,In_4101);
xnor U2357 (N_2357,In_4884,In_3165);
xor U2358 (N_2358,In_4464,In_600);
nor U2359 (N_2359,In_4572,In_632);
nor U2360 (N_2360,In_3463,In_4932);
nor U2361 (N_2361,In_1402,In_1958);
or U2362 (N_2362,In_315,In_648);
nor U2363 (N_2363,In_2374,In_1797);
or U2364 (N_2364,In_66,In_3568);
xnor U2365 (N_2365,In_2427,In_1821);
xor U2366 (N_2366,In_3254,In_2710);
nand U2367 (N_2367,In_553,In_2445);
nand U2368 (N_2368,In_2742,In_401);
nand U2369 (N_2369,In_443,In_1163);
nand U2370 (N_2370,In_39,In_4098);
xor U2371 (N_2371,In_396,In_2262);
nand U2372 (N_2372,In_4809,In_90);
nand U2373 (N_2373,In_2804,In_3494);
xor U2374 (N_2374,In_334,In_4380);
or U2375 (N_2375,In_4434,In_4950);
nor U2376 (N_2376,In_1055,In_3566);
nor U2377 (N_2377,In_4412,In_2978);
nor U2378 (N_2378,In_2773,In_3981);
or U2379 (N_2379,In_3361,In_2999);
nand U2380 (N_2380,In_4325,In_3434);
nor U2381 (N_2381,In_369,In_4824);
nor U2382 (N_2382,In_2765,In_4051);
and U2383 (N_2383,In_4146,In_3053);
and U2384 (N_2384,In_3395,In_3266);
nor U2385 (N_2385,In_2094,In_4991);
xor U2386 (N_2386,In_2379,In_3641);
nor U2387 (N_2387,In_1522,In_4983);
nor U2388 (N_2388,In_2865,In_2704);
and U2389 (N_2389,In_331,In_4568);
xor U2390 (N_2390,In_1147,In_4804);
nand U2391 (N_2391,In_1918,In_1892);
and U2392 (N_2392,In_1311,In_537);
nand U2393 (N_2393,In_3594,In_4845);
or U2394 (N_2394,In_954,In_1789);
nor U2395 (N_2395,In_4300,In_3620);
or U2396 (N_2396,In_832,In_1440);
or U2397 (N_2397,In_955,In_645);
nor U2398 (N_2398,In_1635,In_1344);
and U2399 (N_2399,In_3330,In_3895);
or U2400 (N_2400,In_4079,In_2847);
nand U2401 (N_2401,In_3489,In_371);
and U2402 (N_2402,In_3621,In_2827);
and U2403 (N_2403,In_2910,In_522);
nand U2404 (N_2404,In_4080,In_786);
nor U2405 (N_2405,In_3243,In_3272);
nand U2406 (N_2406,In_4812,In_4540);
xnor U2407 (N_2407,In_2861,In_663);
xor U2408 (N_2408,In_433,In_430);
and U2409 (N_2409,In_3295,In_3055);
nor U2410 (N_2410,In_3593,In_1716);
nand U2411 (N_2411,In_1525,In_4850);
xor U2412 (N_2412,In_4338,In_3390);
and U2413 (N_2413,In_4879,In_4095);
nand U2414 (N_2414,In_4532,In_3986);
nor U2415 (N_2415,In_4131,In_4545);
and U2416 (N_2416,In_3144,In_4607);
or U2417 (N_2417,In_4411,In_779);
or U2418 (N_2418,In_1795,In_100);
or U2419 (N_2419,In_4271,In_3862);
and U2420 (N_2420,In_4735,In_2171);
nor U2421 (N_2421,In_2314,In_4468);
nand U2422 (N_2422,In_2320,In_3586);
or U2423 (N_2423,In_2376,In_4959);
nand U2424 (N_2424,In_1148,In_1363);
or U2425 (N_2425,In_127,In_1137);
nor U2426 (N_2426,In_3883,In_754);
xor U2427 (N_2427,In_3853,In_4939);
nor U2428 (N_2428,In_4688,In_351);
or U2429 (N_2429,In_785,In_3171);
nand U2430 (N_2430,In_3107,In_1073);
and U2431 (N_2431,In_1604,In_3644);
or U2432 (N_2432,In_4455,In_1415);
xnor U2433 (N_2433,In_2571,In_4931);
or U2434 (N_2434,In_3228,In_3219);
xnor U2435 (N_2435,In_801,In_3321);
or U2436 (N_2436,In_833,In_420);
xor U2437 (N_2437,In_1305,In_3374);
xnor U2438 (N_2438,In_3956,In_3557);
and U2439 (N_2439,In_1674,In_1895);
xnor U2440 (N_2440,In_3804,In_4028);
or U2441 (N_2441,In_3101,In_4015);
and U2442 (N_2442,In_3803,In_221);
or U2443 (N_2443,In_4662,In_4625);
or U2444 (N_2444,In_3469,In_4826);
or U2445 (N_2445,In_4913,In_1076);
and U2446 (N_2446,In_1284,In_1765);
or U2447 (N_2447,In_3310,In_2735);
or U2448 (N_2448,In_1209,In_3215);
nor U2449 (N_2449,In_2430,In_4216);
and U2450 (N_2450,In_2886,In_2423);
and U2451 (N_2451,In_281,In_4183);
and U2452 (N_2452,In_208,In_4723);
xnor U2453 (N_2453,In_1811,In_756);
or U2454 (N_2454,In_2405,In_43);
nor U2455 (N_2455,In_2564,In_1537);
nand U2456 (N_2456,In_3957,In_4116);
nand U2457 (N_2457,In_2478,In_4171);
and U2458 (N_2458,In_4087,In_349);
xor U2459 (N_2459,In_4298,In_1893);
or U2460 (N_2460,In_47,In_239);
nand U2461 (N_2461,In_1326,In_367);
xor U2462 (N_2462,In_4590,In_2397);
and U2463 (N_2463,In_2038,In_3447);
xor U2464 (N_2464,In_2106,In_2037);
nand U2465 (N_2465,In_472,In_453);
nor U2466 (N_2466,In_2298,In_340);
and U2467 (N_2467,In_3549,In_4214);
or U2468 (N_2468,In_3209,In_176);
and U2469 (N_2469,In_3821,In_2122);
or U2470 (N_2470,In_503,In_182);
or U2471 (N_2471,In_798,In_2696);
and U2472 (N_2472,In_1644,In_288);
xor U2473 (N_2473,In_2452,In_4122);
nand U2474 (N_2474,In_4790,In_1937);
nor U2475 (N_2475,In_3704,In_3855);
and U2476 (N_2476,In_4643,In_4506);
xor U2477 (N_2477,In_3192,In_3238);
nand U2478 (N_2478,In_4178,In_559);
nand U2479 (N_2479,In_2336,In_4201);
nor U2480 (N_2480,In_3501,In_1979);
xor U2481 (N_2481,In_1526,In_3979);
xor U2482 (N_2482,In_1702,In_1988);
nor U2483 (N_2483,In_547,In_464);
nand U2484 (N_2484,In_120,In_2866);
or U2485 (N_2485,In_2628,In_3547);
nor U2486 (N_2486,In_1383,In_4615);
and U2487 (N_2487,In_4926,In_818);
or U2488 (N_2488,In_566,In_2500);
xnor U2489 (N_2489,In_2815,In_2713);
and U2490 (N_2490,In_346,In_3015);
xnor U2491 (N_2491,In_817,In_2280);
or U2492 (N_2492,In_2219,In_2990);
xor U2493 (N_2493,In_167,In_2962);
or U2494 (N_2494,In_3779,In_3762);
or U2495 (N_2495,In_3433,In_2738);
and U2496 (N_2496,In_4677,In_2775);
nand U2497 (N_2497,In_757,In_3772);
and U2498 (N_2498,In_893,In_4739);
nor U2499 (N_2499,In_2408,In_958);
or U2500 (N_2500,In_4863,In_4032);
nand U2501 (N_2501,In_3764,In_3388);
or U2502 (N_2502,In_726,In_4449);
nor U2503 (N_2503,In_4438,In_4880);
xnor U2504 (N_2504,In_2324,In_2216);
or U2505 (N_2505,In_2557,In_3495);
nor U2506 (N_2506,In_1413,In_4397);
xnor U2507 (N_2507,In_4259,In_628);
nand U2508 (N_2508,In_3806,In_4415);
nor U2509 (N_2509,In_3523,In_1090);
nand U2510 (N_2510,In_1347,In_2688);
or U2511 (N_2511,In_1743,In_781);
nor U2512 (N_2512,In_402,In_3274);
nor U2513 (N_2513,In_2726,In_2332);
nor U2514 (N_2514,In_2463,In_3746);
nand U2515 (N_2515,In_4575,In_4205);
and U2516 (N_2516,In_2987,In_1482);
nand U2517 (N_2517,In_1129,In_637);
nor U2518 (N_2518,In_3740,In_4249);
or U2519 (N_2519,In_994,In_4866);
nand U2520 (N_2520,In_721,In_3902);
nand U2521 (N_2521,In_1995,In_4596);
xor U2522 (N_2522,In_2274,In_3100);
or U2523 (N_2523,In_3558,In_767);
and U2524 (N_2524,In_1217,In_1999);
nor U2525 (N_2525,In_3730,In_2172);
nand U2526 (N_2526,In_1984,In_1960);
nor U2527 (N_2527,In_508,In_3183);
nand U2528 (N_2528,In_4744,In_572);
nand U2529 (N_2529,In_1846,In_4769);
nor U2530 (N_2530,In_4334,In_3694);
and U2531 (N_2531,In_2706,In_4193);
xor U2532 (N_2532,In_1850,In_2647);
and U2533 (N_2533,In_2678,In_2932);
or U2534 (N_2534,In_3625,In_3650);
nand U2535 (N_2535,In_3518,In_2492);
nor U2536 (N_2536,In_1931,In_531);
nand U2537 (N_2537,In_547,In_1425);
xnor U2538 (N_2538,In_3105,In_1284);
or U2539 (N_2539,In_4552,In_4031);
nor U2540 (N_2540,In_1811,In_1568);
or U2541 (N_2541,In_3393,In_1027);
nand U2542 (N_2542,In_3328,In_4224);
nand U2543 (N_2543,In_3204,In_3599);
and U2544 (N_2544,In_2832,In_4016);
xor U2545 (N_2545,In_947,In_2120);
nor U2546 (N_2546,In_3618,In_1558);
nand U2547 (N_2547,In_4535,In_3410);
nand U2548 (N_2548,In_1371,In_1830);
xnor U2549 (N_2549,In_895,In_3384);
and U2550 (N_2550,In_176,In_3840);
or U2551 (N_2551,In_3422,In_4421);
and U2552 (N_2552,In_1900,In_898);
xnor U2553 (N_2553,In_4442,In_1085);
or U2554 (N_2554,In_1654,In_2294);
and U2555 (N_2555,In_4813,In_3960);
xor U2556 (N_2556,In_3646,In_896);
and U2557 (N_2557,In_4585,In_4393);
nor U2558 (N_2558,In_2695,In_533);
nand U2559 (N_2559,In_3086,In_1189);
or U2560 (N_2560,In_3528,In_4403);
xnor U2561 (N_2561,In_2253,In_2149);
xor U2562 (N_2562,In_3527,In_4682);
and U2563 (N_2563,In_4335,In_2694);
nand U2564 (N_2564,In_3866,In_3331);
or U2565 (N_2565,In_1521,In_4951);
nand U2566 (N_2566,In_4367,In_3007);
or U2567 (N_2567,In_2251,In_4830);
xnor U2568 (N_2568,In_4558,In_734);
nand U2569 (N_2569,In_447,In_1631);
nand U2570 (N_2570,In_4683,In_3961);
nand U2571 (N_2571,In_992,In_1498);
xnor U2572 (N_2572,In_2948,In_3824);
nor U2573 (N_2573,In_2783,In_1984);
nor U2574 (N_2574,In_3256,In_4899);
xnor U2575 (N_2575,In_4489,In_2178);
nor U2576 (N_2576,In_465,In_3825);
and U2577 (N_2577,In_2029,In_2051);
xnor U2578 (N_2578,In_4684,In_3843);
nor U2579 (N_2579,In_995,In_2392);
nor U2580 (N_2580,In_3647,In_2912);
or U2581 (N_2581,In_1684,In_2259);
or U2582 (N_2582,In_2242,In_4183);
nand U2583 (N_2583,In_4331,In_1188);
nor U2584 (N_2584,In_4934,In_1325);
nor U2585 (N_2585,In_4070,In_2738);
or U2586 (N_2586,In_2641,In_4975);
xnor U2587 (N_2587,In_2443,In_2486);
xnor U2588 (N_2588,In_4269,In_4273);
and U2589 (N_2589,In_1760,In_3263);
xnor U2590 (N_2590,In_4374,In_3155);
or U2591 (N_2591,In_4093,In_3901);
nor U2592 (N_2592,In_1326,In_3816);
and U2593 (N_2593,In_1185,In_1747);
or U2594 (N_2594,In_3616,In_4017);
nand U2595 (N_2595,In_4681,In_2049);
or U2596 (N_2596,In_4758,In_2986);
and U2597 (N_2597,In_3438,In_52);
or U2598 (N_2598,In_4307,In_3987);
nand U2599 (N_2599,In_4257,In_2054);
nand U2600 (N_2600,In_110,In_3740);
and U2601 (N_2601,In_3427,In_1566);
xor U2602 (N_2602,In_4655,In_2781);
nand U2603 (N_2603,In_1176,In_1314);
xor U2604 (N_2604,In_830,In_295);
or U2605 (N_2605,In_555,In_3405);
and U2606 (N_2606,In_901,In_4866);
nand U2607 (N_2607,In_232,In_934);
xnor U2608 (N_2608,In_2248,In_2915);
nand U2609 (N_2609,In_971,In_4385);
xnor U2610 (N_2610,In_1807,In_935);
nor U2611 (N_2611,In_2495,In_76);
nor U2612 (N_2612,In_3184,In_4952);
xor U2613 (N_2613,In_712,In_3835);
xor U2614 (N_2614,In_3637,In_3005);
or U2615 (N_2615,In_1901,In_3472);
and U2616 (N_2616,In_657,In_3668);
and U2617 (N_2617,In_1656,In_2808);
and U2618 (N_2618,In_1609,In_2035);
nor U2619 (N_2619,In_4863,In_545);
nand U2620 (N_2620,In_1093,In_741);
nand U2621 (N_2621,In_2321,In_2648);
nor U2622 (N_2622,In_1014,In_1356);
or U2623 (N_2623,In_1546,In_1230);
nor U2624 (N_2624,In_3220,In_6);
nor U2625 (N_2625,In_2378,In_2565);
or U2626 (N_2626,In_4348,In_4456);
xor U2627 (N_2627,In_3979,In_2595);
nand U2628 (N_2628,In_3711,In_4924);
xor U2629 (N_2629,In_2065,In_4332);
nand U2630 (N_2630,In_2474,In_3807);
or U2631 (N_2631,In_172,In_3981);
or U2632 (N_2632,In_2105,In_4624);
nand U2633 (N_2633,In_481,In_4134);
nor U2634 (N_2634,In_1721,In_3797);
nor U2635 (N_2635,In_1891,In_3945);
xor U2636 (N_2636,In_2879,In_2510);
nand U2637 (N_2637,In_4270,In_2237);
xnor U2638 (N_2638,In_4983,In_3520);
or U2639 (N_2639,In_3577,In_2623);
or U2640 (N_2640,In_49,In_4490);
nor U2641 (N_2641,In_2410,In_3941);
or U2642 (N_2642,In_1806,In_182);
nor U2643 (N_2643,In_2160,In_306);
or U2644 (N_2644,In_1889,In_1674);
or U2645 (N_2645,In_2045,In_3942);
or U2646 (N_2646,In_3074,In_4259);
or U2647 (N_2647,In_1405,In_3029);
or U2648 (N_2648,In_1201,In_1047);
nor U2649 (N_2649,In_3713,In_1069);
or U2650 (N_2650,In_2670,In_1973);
nor U2651 (N_2651,In_2623,In_1553);
nor U2652 (N_2652,In_1418,In_3899);
nor U2653 (N_2653,In_405,In_1941);
nor U2654 (N_2654,In_1663,In_3329);
nand U2655 (N_2655,In_1530,In_4531);
nor U2656 (N_2656,In_4972,In_1074);
xor U2657 (N_2657,In_2182,In_4036);
or U2658 (N_2658,In_4956,In_2749);
nor U2659 (N_2659,In_176,In_156);
xor U2660 (N_2660,In_451,In_790);
or U2661 (N_2661,In_943,In_4342);
nand U2662 (N_2662,In_1824,In_3929);
and U2663 (N_2663,In_2602,In_46);
nand U2664 (N_2664,In_3511,In_4158);
nor U2665 (N_2665,In_3956,In_3594);
or U2666 (N_2666,In_1766,In_3144);
nor U2667 (N_2667,In_4494,In_2528);
nand U2668 (N_2668,In_2059,In_4546);
xnor U2669 (N_2669,In_4530,In_2774);
xnor U2670 (N_2670,In_2113,In_4050);
or U2671 (N_2671,In_1747,In_2128);
and U2672 (N_2672,In_4887,In_1568);
xor U2673 (N_2673,In_3107,In_1770);
and U2674 (N_2674,In_3422,In_2753);
nor U2675 (N_2675,In_2836,In_4902);
and U2676 (N_2676,In_4015,In_274);
xor U2677 (N_2677,In_362,In_1021);
nand U2678 (N_2678,In_1188,In_4621);
nor U2679 (N_2679,In_4736,In_3260);
or U2680 (N_2680,In_2341,In_4644);
xnor U2681 (N_2681,In_2644,In_217);
nor U2682 (N_2682,In_4187,In_1733);
or U2683 (N_2683,In_4606,In_3780);
nand U2684 (N_2684,In_3168,In_468);
nand U2685 (N_2685,In_3587,In_186);
or U2686 (N_2686,In_4432,In_3762);
xnor U2687 (N_2687,In_4935,In_4066);
or U2688 (N_2688,In_44,In_728);
xor U2689 (N_2689,In_1244,In_2012);
or U2690 (N_2690,In_577,In_1588);
nand U2691 (N_2691,In_4551,In_3730);
or U2692 (N_2692,In_4188,In_3268);
nor U2693 (N_2693,In_4173,In_3642);
and U2694 (N_2694,In_2566,In_975);
nand U2695 (N_2695,In_101,In_4225);
xnor U2696 (N_2696,In_3142,In_1215);
and U2697 (N_2697,In_1380,In_3406);
or U2698 (N_2698,In_2924,In_1412);
nand U2699 (N_2699,In_293,In_569);
nand U2700 (N_2700,In_4152,In_4349);
nand U2701 (N_2701,In_2619,In_1593);
nor U2702 (N_2702,In_904,In_2784);
and U2703 (N_2703,In_717,In_3767);
xnor U2704 (N_2704,In_2740,In_4803);
and U2705 (N_2705,In_3737,In_763);
nor U2706 (N_2706,In_3812,In_1313);
and U2707 (N_2707,In_141,In_4925);
or U2708 (N_2708,In_297,In_3546);
nand U2709 (N_2709,In_3329,In_3991);
and U2710 (N_2710,In_3468,In_2296);
or U2711 (N_2711,In_1798,In_1888);
or U2712 (N_2712,In_1048,In_3507);
xnor U2713 (N_2713,In_99,In_2735);
and U2714 (N_2714,In_4298,In_1675);
and U2715 (N_2715,In_830,In_1094);
nand U2716 (N_2716,In_4561,In_4121);
or U2717 (N_2717,In_4956,In_2557);
nand U2718 (N_2718,In_3708,In_665);
and U2719 (N_2719,In_1925,In_3563);
xnor U2720 (N_2720,In_236,In_633);
xnor U2721 (N_2721,In_37,In_3073);
nor U2722 (N_2722,In_1069,In_1063);
nor U2723 (N_2723,In_703,In_1541);
xor U2724 (N_2724,In_2696,In_4325);
and U2725 (N_2725,In_3748,In_3362);
and U2726 (N_2726,In_992,In_1072);
nand U2727 (N_2727,In_3828,In_1848);
and U2728 (N_2728,In_4818,In_590);
or U2729 (N_2729,In_249,In_208);
nand U2730 (N_2730,In_571,In_4424);
xor U2731 (N_2731,In_1355,In_4114);
xnor U2732 (N_2732,In_2115,In_1007);
or U2733 (N_2733,In_318,In_3091);
nor U2734 (N_2734,In_523,In_4561);
nor U2735 (N_2735,In_1699,In_1807);
nor U2736 (N_2736,In_222,In_1667);
nand U2737 (N_2737,In_4573,In_1720);
or U2738 (N_2738,In_4859,In_148);
xnor U2739 (N_2739,In_1273,In_3975);
nor U2740 (N_2740,In_2282,In_323);
xnor U2741 (N_2741,In_1320,In_207);
and U2742 (N_2742,In_2810,In_1356);
xor U2743 (N_2743,In_2700,In_3389);
and U2744 (N_2744,In_3202,In_3565);
and U2745 (N_2745,In_582,In_684);
nand U2746 (N_2746,In_1974,In_4453);
xor U2747 (N_2747,In_3402,In_300);
or U2748 (N_2748,In_4836,In_3173);
xor U2749 (N_2749,In_1218,In_1973);
and U2750 (N_2750,In_2221,In_669);
nand U2751 (N_2751,In_517,In_3574);
xor U2752 (N_2752,In_2533,In_4903);
nor U2753 (N_2753,In_1821,In_3697);
or U2754 (N_2754,In_1049,In_438);
or U2755 (N_2755,In_2328,In_4665);
nor U2756 (N_2756,In_3435,In_915);
nor U2757 (N_2757,In_1410,In_1567);
and U2758 (N_2758,In_3294,In_1096);
nor U2759 (N_2759,In_3260,In_3731);
xnor U2760 (N_2760,In_3540,In_2515);
nand U2761 (N_2761,In_4243,In_1091);
xnor U2762 (N_2762,In_4471,In_3006);
and U2763 (N_2763,In_846,In_900);
or U2764 (N_2764,In_2579,In_4696);
or U2765 (N_2765,In_1527,In_4277);
nand U2766 (N_2766,In_4536,In_2353);
nor U2767 (N_2767,In_4729,In_3165);
or U2768 (N_2768,In_3581,In_174);
nand U2769 (N_2769,In_4884,In_3782);
and U2770 (N_2770,In_83,In_789);
or U2771 (N_2771,In_4921,In_1291);
nor U2772 (N_2772,In_643,In_305);
nand U2773 (N_2773,In_350,In_2042);
nand U2774 (N_2774,In_2858,In_4780);
and U2775 (N_2775,In_834,In_3670);
or U2776 (N_2776,In_2204,In_4837);
and U2777 (N_2777,In_3094,In_2085);
nand U2778 (N_2778,In_1007,In_3315);
and U2779 (N_2779,In_1682,In_2966);
or U2780 (N_2780,In_2776,In_2896);
nand U2781 (N_2781,In_2299,In_3386);
or U2782 (N_2782,In_3561,In_877);
nand U2783 (N_2783,In_3507,In_4742);
and U2784 (N_2784,In_3295,In_1997);
or U2785 (N_2785,In_4097,In_1302);
or U2786 (N_2786,In_722,In_2683);
or U2787 (N_2787,In_2095,In_469);
or U2788 (N_2788,In_37,In_3465);
nand U2789 (N_2789,In_4365,In_1436);
nand U2790 (N_2790,In_89,In_111);
nor U2791 (N_2791,In_676,In_3061);
or U2792 (N_2792,In_2701,In_2306);
nand U2793 (N_2793,In_2398,In_4263);
and U2794 (N_2794,In_4259,In_1804);
and U2795 (N_2795,In_3971,In_552);
or U2796 (N_2796,In_4816,In_684);
nor U2797 (N_2797,In_1419,In_210);
or U2798 (N_2798,In_4405,In_1699);
xnor U2799 (N_2799,In_1436,In_4572);
nor U2800 (N_2800,In_1941,In_4317);
or U2801 (N_2801,In_288,In_3206);
nor U2802 (N_2802,In_1790,In_4866);
xor U2803 (N_2803,In_4924,In_2245);
nand U2804 (N_2804,In_2129,In_3728);
and U2805 (N_2805,In_3534,In_3436);
and U2806 (N_2806,In_3899,In_842);
or U2807 (N_2807,In_2065,In_831);
nor U2808 (N_2808,In_2449,In_1789);
nand U2809 (N_2809,In_1807,In_361);
xnor U2810 (N_2810,In_4045,In_87);
nor U2811 (N_2811,In_4552,In_3592);
nand U2812 (N_2812,In_979,In_1458);
nand U2813 (N_2813,In_1473,In_54);
nand U2814 (N_2814,In_4158,In_345);
xor U2815 (N_2815,In_1696,In_2286);
xnor U2816 (N_2816,In_1411,In_4304);
nor U2817 (N_2817,In_2684,In_1451);
xor U2818 (N_2818,In_3100,In_1850);
nand U2819 (N_2819,In_3386,In_3590);
and U2820 (N_2820,In_2752,In_4093);
nand U2821 (N_2821,In_1735,In_437);
xnor U2822 (N_2822,In_4489,In_1301);
nor U2823 (N_2823,In_1367,In_163);
nand U2824 (N_2824,In_2294,In_2576);
and U2825 (N_2825,In_4615,In_3334);
xnor U2826 (N_2826,In_907,In_1399);
xnor U2827 (N_2827,In_2341,In_1488);
and U2828 (N_2828,In_2932,In_519);
nand U2829 (N_2829,In_2402,In_1760);
xor U2830 (N_2830,In_2334,In_1090);
nor U2831 (N_2831,In_2454,In_4411);
xnor U2832 (N_2832,In_509,In_1997);
nand U2833 (N_2833,In_4025,In_2785);
or U2834 (N_2834,In_2526,In_3144);
nand U2835 (N_2835,In_4609,In_2098);
nand U2836 (N_2836,In_3562,In_4740);
or U2837 (N_2837,In_1901,In_939);
xnor U2838 (N_2838,In_650,In_2033);
or U2839 (N_2839,In_4810,In_4114);
xnor U2840 (N_2840,In_4139,In_4785);
xor U2841 (N_2841,In_2758,In_1988);
nor U2842 (N_2842,In_523,In_4725);
nor U2843 (N_2843,In_1964,In_2417);
or U2844 (N_2844,In_3963,In_1616);
nor U2845 (N_2845,In_4543,In_3131);
nand U2846 (N_2846,In_4443,In_2407);
and U2847 (N_2847,In_1488,In_1720);
and U2848 (N_2848,In_1159,In_1728);
nor U2849 (N_2849,In_4171,In_1797);
or U2850 (N_2850,In_2555,In_1970);
or U2851 (N_2851,In_3119,In_908);
or U2852 (N_2852,In_1564,In_3307);
nand U2853 (N_2853,In_1040,In_102);
and U2854 (N_2854,In_201,In_3911);
xor U2855 (N_2855,In_2970,In_3541);
or U2856 (N_2856,In_3776,In_1323);
and U2857 (N_2857,In_3452,In_4753);
or U2858 (N_2858,In_1812,In_3556);
and U2859 (N_2859,In_263,In_4338);
or U2860 (N_2860,In_4040,In_222);
and U2861 (N_2861,In_2220,In_3691);
and U2862 (N_2862,In_1428,In_4855);
and U2863 (N_2863,In_2546,In_3372);
nand U2864 (N_2864,In_2025,In_4958);
nor U2865 (N_2865,In_4536,In_2373);
nand U2866 (N_2866,In_149,In_1225);
nor U2867 (N_2867,In_4710,In_3402);
or U2868 (N_2868,In_2570,In_3181);
or U2869 (N_2869,In_2355,In_1775);
or U2870 (N_2870,In_600,In_163);
and U2871 (N_2871,In_845,In_4984);
and U2872 (N_2872,In_136,In_694);
nand U2873 (N_2873,In_4264,In_1700);
or U2874 (N_2874,In_3784,In_4245);
nand U2875 (N_2875,In_507,In_1711);
and U2876 (N_2876,In_428,In_2057);
or U2877 (N_2877,In_4893,In_247);
nand U2878 (N_2878,In_4334,In_2632);
xnor U2879 (N_2879,In_301,In_3734);
nor U2880 (N_2880,In_3575,In_1517);
nand U2881 (N_2881,In_1483,In_4222);
and U2882 (N_2882,In_3771,In_217);
nor U2883 (N_2883,In_1139,In_1367);
and U2884 (N_2884,In_623,In_4714);
nand U2885 (N_2885,In_1555,In_3959);
or U2886 (N_2886,In_2237,In_4980);
nand U2887 (N_2887,In_4915,In_4282);
xnor U2888 (N_2888,In_3343,In_4050);
and U2889 (N_2889,In_3973,In_3265);
nor U2890 (N_2890,In_4477,In_1781);
nand U2891 (N_2891,In_2871,In_1350);
or U2892 (N_2892,In_2098,In_802);
nand U2893 (N_2893,In_3125,In_1912);
xnor U2894 (N_2894,In_2180,In_4060);
nand U2895 (N_2895,In_170,In_1829);
nand U2896 (N_2896,In_278,In_4897);
or U2897 (N_2897,In_1747,In_824);
or U2898 (N_2898,In_3767,In_3120);
and U2899 (N_2899,In_3410,In_1611);
xor U2900 (N_2900,In_4548,In_1409);
nor U2901 (N_2901,In_2394,In_943);
nor U2902 (N_2902,In_4636,In_1393);
xor U2903 (N_2903,In_3966,In_4336);
nand U2904 (N_2904,In_3827,In_1577);
or U2905 (N_2905,In_1507,In_1888);
nor U2906 (N_2906,In_3301,In_2208);
nand U2907 (N_2907,In_2670,In_3502);
nand U2908 (N_2908,In_1686,In_2292);
and U2909 (N_2909,In_3394,In_1349);
and U2910 (N_2910,In_4021,In_1481);
xor U2911 (N_2911,In_1675,In_279);
xor U2912 (N_2912,In_2412,In_320);
or U2913 (N_2913,In_4831,In_1561);
and U2914 (N_2914,In_4370,In_3690);
xnor U2915 (N_2915,In_2307,In_2969);
nor U2916 (N_2916,In_2508,In_4790);
or U2917 (N_2917,In_1236,In_4829);
nand U2918 (N_2918,In_2911,In_1703);
nand U2919 (N_2919,In_687,In_2734);
and U2920 (N_2920,In_988,In_1938);
or U2921 (N_2921,In_1792,In_520);
and U2922 (N_2922,In_2600,In_1798);
or U2923 (N_2923,In_1505,In_41);
nor U2924 (N_2924,In_2007,In_2981);
or U2925 (N_2925,In_10,In_3761);
and U2926 (N_2926,In_4605,In_2238);
nor U2927 (N_2927,In_1211,In_1819);
nor U2928 (N_2928,In_712,In_4160);
nand U2929 (N_2929,In_4566,In_1123);
nand U2930 (N_2930,In_3474,In_4129);
or U2931 (N_2931,In_673,In_2768);
and U2932 (N_2932,In_3032,In_4384);
xnor U2933 (N_2933,In_4130,In_625);
nand U2934 (N_2934,In_4041,In_3904);
nand U2935 (N_2935,In_358,In_1082);
nand U2936 (N_2936,In_3196,In_1781);
nor U2937 (N_2937,In_2661,In_592);
nor U2938 (N_2938,In_4515,In_728);
xnor U2939 (N_2939,In_3681,In_80);
xor U2940 (N_2940,In_4895,In_4627);
xor U2941 (N_2941,In_2952,In_3251);
or U2942 (N_2942,In_504,In_4569);
and U2943 (N_2943,In_3088,In_1402);
xor U2944 (N_2944,In_2448,In_4053);
nand U2945 (N_2945,In_4297,In_4589);
xor U2946 (N_2946,In_3886,In_1165);
and U2947 (N_2947,In_819,In_4939);
nor U2948 (N_2948,In_3074,In_4326);
or U2949 (N_2949,In_4257,In_1839);
or U2950 (N_2950,In_4163,In_3856);
xnor U2951 (N_2951,In_3939,In_1133);
and U2952 (N_2952,In_3206,In_3849);
nor U2953 (N_2953,In_4519,In_335);
and U2954 (N_2954,In_3961,In_1010);
nor U2955 (N_2955,In_3253,In_459);
or U2956 (N_2956,In_2862,In_2341);
nor U2957 (N_2957,In_4306,In_4030);
and U2958 (N_2958,In_3504,In_4548);
or U2959 (N_2959,In_4858,In_1470);
nand U2960 (N_2960,In_4552,In_3210);
nor U2961 (N_2961,In_3428,In_1632);
and U2962 (N_2962,In_2361,In_773);
or U2963 (N_2963,In_4898,In_77);
nor U2964 (N_2964,In_1072,In_1840);
nor U2965 (N_2965,In_4507,In_2054);
nand U2966 (N_2966,In_3182,In_4675);
and U2967 (N_2967,In_1568,In_4894);
and U2968 (N_2968,In_2909,In_2621);
or U2969 (N_2969,In_1120,In_1931);
or U2970 (N_2970,In_2950,In_897);
and U2971 (N_2971,In_1417,In_122);
nand U2972 (N_2972,In_938,In_4773);
nand U2973 (N_2973,In_1002,In_1582);
xor U2974 (N_2974,In_980,In_3546);
and U2975 (N_2975,In_1857,In_3515);
nand U2976 (N_2976,In_2617,In_3756);
nor U2977 (N_2977,In_78,In_289);
nand U2978 (N_2978,In_2622,In_1493);
or U2979 (N_2979,In_435,In_25);
nand U2980 (N_2980,In_1266,In_1114);
nor U2981 (N_2981,In_3223,In_3064);
xnor U2982 (N_2982,In_558,In_1997);
xnor U2983 (N_2983,In_2012,In_1213);
and U2984 (N_2984,In_56,In_3626);
nand U2985 (N_2985,In_1280,In_4316);
xnor U2986 (N_2986,In_1082,In_1541);
and U2987 (N_2987,In_1402,In_3020);
nand U2988 (N_2988,In_1756,In_1279);
xor U2989 (N_2989,In_1191,In_1115);
nand U2990 (N_2990,In_2978,In_565);
nand U2991 (N_2991,In_2005,In_4072);
and U2992 (N_2992,In_252,In_3009);
xnor U2993 (N_2993,In_3902,In_2281);
and U2994 (N_2994,In_541,In_4295);
or U2995 (N_2995,In_111,In_1075);
and U2996 (N_2996,In_4164,In_306);
nand U2997 (N_2997,In_4596,In_3540);
or U2998 (N_2998,In_111,In_2060);
nand U2999 (N_2999,In_2961,In_1997);
nor U3000 (N_3000,In_4693,In_2432);
nor U3001 (N_3001,In_1594,In_2122);
nor U3002 (N_3002,In_171,In_3713);
nor U3003 (N_3003,In_4109,In_680);
nand U3004 (N_3004,In_3231,In_312);
or U3005 (N_3005,In_780,In_2670);
xnor U3006 (N_3006,In_3335,In_910);
or U3007 (N_3007,In_4475,In_4421);
or U3008 (N_3008,In_1970,In_2620);
or U3009 (N_3009,In_4779,In_1932);
and U3010 (N_3010,In_856,In_2275);
xnor U3011 (N_3011,In_1700,In_2308);
or U3012 (N_3012,In_4760,In_3466);
xor U3013 (N_3013,In_996,In_4737);
xor U3014 (N_3014,In_4728,In_4198);
or U3015 (N_3015,In_3460,In_4482);
xnor U3016 (N_3016,In_3109,In_126);
nand U3017 (N_3017,In_2797,In_1098);
and U3018 (N_3018,In_4325,In_2755);
xor U3019 (N_3019,In_4017,In_4863);
nand U3020 (N_3020,In_3710,In_564);
or U3021 (N_3021,In_506,In_3300);
nor U3022 (N_3022,In_1258,In_2746);
nor U3023 (N_3023,In_3132,In_2212);
nor U3024 (N_3024,In_2808,In_1129);
xnor U3025 (N_3025,In_37,In_1186);
xnor U3026 (N_3026,In_3109,In_4707);
or U3027 (N_3027,In_3271,In_3944);
nor U3028 (N_3028,In_2672,In_1736);
xnor U3029 (N_3029,In_702,In_698);
nand U3030 (N_3030,In_1456,In_2999);
nor U3031 (N_3031,In_4084,In_595);
or U3032 (N_3032,In_3777,In_2275);
nor U3033 (N_3033,In_169,In_3203);
nor U3034 (N_3034,In_4445,In_4112);
xnor U3035 (N_3035,In_1,In_4375);
nor U3036 (N_3036,In_4356,In_3081);
and U3037 (N_3037,In_4591,In_2304);
or U3038 (N_3038,In_3481,In_1382);
and U3039 (N_3039,In_35,In_325);
or U3040 (N_3040,In_654,In_1666);
nor U3041 (N_3041,In_4125,In_875);
xnor U3042 (N_3042,In_1794,In_1774);
and U3043 (N_3043,In_4277,In_539);
nand U3044 (N_3044,In_4467,In_2616);
and U3045 (N_3045,In_4846,In_3271);
or U3046 (N_3046,In_659,In_365);
nor U3047 (N_3047,In_4151,In_879);
nor U3048 (N_3048,In_2982,In_4195);
nand U3049 (N_3049,In_2950,In_4523);
or U3050 (N_3050,In_3017,In_1046);
nor U3051 (N_3051,In_4514,In_2007);
and U3052 (N_3052,In_1220,In_931);
xor U3053 (N_3053,In_649,In_1962);
nand U3054 (N_3054,In_4892,In_4858);
or U3055 (N_3055,In_1079,In_156);
nand U3056 (N_3056,In_2130,In_3307);
nand U3057 (N_3057,In_2886,In_4161);
or U3058 (N_3058,In_3310,In_1075);
nand U3059 (N_3059,In_3342,In_1953);
or U3060 (N_3060,In_4860,In_1138);
nor U3061 (N_3061,In_3659,In_3646);
or U3062 (N_3062,In_2622,In_1990);
nor U3063 (N_3063,In_3597,In_3002);
nand U3064 (N_3064,In_2137,In_2422);
xnor U3065 (N_3065,In_1199,In_3286);
and U3066 (N_3066,In_4280,In_4572);
nor U3067 (N_3067,In_479,In_1288);
nand U3068 (N_3068,In_3624,In_1383);
or U3069 (N_3069,In_3375,In_2997);
nand U3070 (N_3070,In_1616,In_2994);
nor U3071 (N_3071,In_3428,In_1656);
nand U3072 (N_3072,In_1493,In_109);
nor U3073 (N_3073,In_3722,In_3091);
nand U3074 (N_3074,In_4016,In_4282);
and U3075 (N_3075,In_657,In_1601);
or U3076 (N_3076,In_2586,In_3662);
or U3077 (N_3077,In_3945,In_631);
and U3078 (N_3078,In_4556,In_1669);
xor U3079 (N_3079,In_49,In_442);
nor U3080 (N_3080,In_822,In_4603);
nor U3081 (N_3081,In_2045,In_4549);
or U3082 (N_3082,In_2322,In_3932);
xnor U3083 (N_3083,In_4436,In_3704);
or U3084 (N_3084,In_1931,In_73);
nor U3085 (N_3085,In_451,In_3976);
or U3086 (N_3086,In_2435,In_3267);
nor U3087 (N_3087,In_3406,In_2279);
or U3088 (N_3088,In_1628,In_1844);
xnor U3089 (N_3089,In_82,In_559);
nor U3090 (N_3090,In_4955,In_4427);
nor U3091 (N_3091,In_1443,In_1685);
or U3092 (N_3092,In_3048,In_306);
and U3093 (N_3093,In_2457,In_4989);
nand U3094 (N_3094,In_1863,In_857);
nor U3095 (N_3095,In_2253,In_1212);
or U3096 (N_3096,In_987,In_2862);
xor U3097 (N_3097,In_4344,In_1639);
and U3098 (N_3098,In_4864,In_4061);
or U3099 (N_3099,In_229,In_607);
and U3100 (N_3100,In_2550,In_3705);
nor U3101 (N_3101,In_2422,In_4951);
or U3102 (N_3102,In_2815,In_492);
nand U3103 (N_3103,In_1443,In_1297);
or U3104 (N_3104,In_477,In_305);
nor U3105 (N_3105,In_4433,In_3175);
and U3106 (N_3106,In_2918,In_3577);
nand U3107 (N_3107,In_2858,In_441);
or U3108 (N_3108,In_4465,In_4283);
nor U3109 (N_3109,In_1554,In_2568);
nand U3110 (N_3110,In_1625,In_4384);
and U3111 (N_3111,In_2868,In_4897);
and U3112 (N_3112,In_881,In_2576);
and U3113 (N_3113,In_121,In_3046);
nor U3114 (N_3114,In_3548,In_4796);
nand U3115 (N_3115,In_3331,In_4482);
nor U3116 (N_3116,In_740,In_2287);
and U3117 (N_3117,In_4795,In_2274);
and U3118 (N_3118,In_4227,In_2238);
or U3119 (N_3119,In_4838,In_1299);
or U3120 (N_3120,In_742,In_362);
nand U3121 (N_3121,In_2576,In_4548);
or U3122 (N_3122,In_3094,In_1242);
and U3123 (N_3123,In_2758,In_3374);
nand U3124 (N_3124,In_647,In_240);
and U3125 (N_3125,In_61,In_4452);
or U3126 (N_3126,In_3212,In_976);
xor U3127 (N_3127,In_3593,In_1654);
nor U3128 (N_3128,In_2025,In_175);
xor U3129 (N_3129,In_565,In_868);
nor U3130 (N_3130,In_4088,In_3190);
and U3131 (N_3131,In_168,In_54);
nand U3132 (N_3132,In_2779,In_3340);
and U3133 (N_3133,In_1004,In_3463);
and U3134 (N_3134,In_2220,In_3675);
and U3135 (N_3135,In_3607,In_3784);
and U3136 (N_3136,In_722,In_581);
nor U3137 (N_3137,In_1780,In_3964);
nor U3138 (N_3138,In_1783,In_2752);
nand U3139 (N_3139,In_4866,In_151);
xnor U3140 (N_3140,In_4570,In_4064);
nor U3141 (N_3141,In_3334,In_2226);
and U3142 (N_3142,In_4957,In_4342);
or U3143 (N_3143,In_256,In_3616);
or U3144 (N_3144,In_2138,In_4410);
nand U3145 (N_3145,In_1529,In_920);
nor U3146 (N_3146,In_3526,In_863);
or U3147 (N_3147,In_2361,In_1050);
nor U3148 (N_3148,In_3040,In_1828);
nand U3149 (N_3149,In_2870,In_1618);
xor U3150 (N_3150,In_2375,In_2092);
nor U3151 (N_3151,In_595,In_69);
or U3152 (N_3152,In_3996,In_4961);
and U3153 (N_3153,In_2318,In_3202);
or U3154 (N_3154,In_4453,In_3870);
and U3155 (N_3155,In_2140,In_2941);
and U3156 (N_3156,In_1701,In_169);
nor U3157 (N_3157,In_755,In_1038);
nand U3158 (N_3158,In_3838,In_845);
and U3159 (N_3159,In_8,In_1069);
or U3160 (N_3160,In_4727,In_910);
and U3161 (N_3161,In_1416,In_4586);
and U3162 (N_3162,In_1973,In_2445);
nand U3163 (N_3163,In_1546,In_151);
nand U3164 (N_3164,In_769,In_4348);
and U3165 (N_3165,In_2918,In_304);
xor U3166 (N_3166,In_3276,In_646);
and U3167 (N_3167,In_2927,In_4733);
and U3168 (N_3168,In_4969,In_2276);
nand U3169 (N_3169,In_4075,In_1238);
and U3170 (N_3170,In_1984,In_2386);
xnor U3171 (N_3171,In_2605,In_2777);
or U3172 (N_3172,In_4390,In_3113);
nand U3173 (N_3173,In_3951,In_2514);
nand U3174 (N_3174,In_2670,In_2634);
nor U3175 (N_3175,In_2599,In_4711);
or U3176 (N_3176,In_3726,In_973);
xnor U3177 (N_3177,In_586,In_4529);
nand U3178 (N_3178,In_3693,In_79);
or U3179 (N_3179,In_1614,In_4280);
nor U3180 (N_3180,In_2205,In_178);
xor U3181 (N_3181,In_4327,In_4686);
nand U3182 (N_3182,In_433,In_4981);
and U3183 (N_3183,In_2887,In_225);
nor U3184 (N_3184,In_3352,In_3758);
nand U3185 (N_3185,In_323,In_766);
nor U3186 (N_3186,In_3779,In_1803);
and U3187 (N_3187,In_417,In_1124);
xnor U3188 (N_3188,In_159,In_3674);
xnor U3189 (N_3189,In_2582,In_4727);
nand U3190 (N_3190,In_3963,In_3441);
or U3191 (N_3191,In_1397,In_2236);
nand U3192 (N_3192,In_1075,In_4981);
and U3193 (N_3193,In_3404,In_900);
and U3194 (N_3194,In_2243,In_230);
nor U3195 (N_3195,In_3256,In_2132);
nor U3196 (N_3196,In_3203,In_1367);
and U3197 (N_3197,In_1280,In_4944);
and U3198 (N_3198,In_2626,In_2970);
or U3199 (N_3199,In_2539,In_3636);
and U3200 (N_3200,In_1733,In_3441);
xnor U3201 (N_3201,In_4539,In_488);
nand U3202 (N_3202,In_1904,In_2349);
and U3203 (N_3203,In_4238,In_3574);
or U3204 (N_3204,In_4433,In_2088);
nand U3205 (N_3205,In_4245,In_3079);
or U3206 (N_3206,In_1695,In_4118);
and U3207 (N_3207,In_3862,In_2497);
nor U3208 (N_3208,In_952,In_415);
nand U3209 (N_3209,In_4320,In_2929);
nor U3210 (N_3210,In_3043,In_914);
and U3211 (N_3211,In_2326,In_4473);
nor U3212 (N_3212,In_1824,In_2729);
nor U3213 (N_3213,In_3444,In_785);
or U3214 (N_3214,In_4542,In_2714);
nor U3215 (N_3215,In_2995,In_3128);
nand U3216 (N_3216,In_4094,In_993);
and U3217 (N_3217,In_662,In_3862);
and U3218 (N_3218,In_3112,In_2984);
or U3219 (N_3219,In_2392,In_3929);
nor U3220 (N_3220,In_462,In_2477);
nor U3221 (N_3221,In_4295,In_3009);
xnor U3222 (N_3222,In_1199,In_4581);
nand U3223 (N_3223,In_2762,In_2219);
and U3224 (N_3224,In_124,In_740);
nor U3225 (N_3225,In_4453,In_4837);
xor U3226 (N_3226,In_901,In_1515);
xnor U3227 (N_3227,In_3477,In_4435);
or U3228 (N_3228,In_1559,In_4503);
nand U3229 (N_3229,In_1111,In_984);
nor U3230 (N_3230,In_1853,In_3940);
nor U3231 (N_3231,In_4484,In_117);
and U3232 (N_3232,In_4006,In_1826);
nand U3233 (N_3233,In_1704,In_2660);
nor U3234 (N_3234,In_81,In_1107);
nor U3235 (N_3235,In_2837,In_1708);
xor U3236 (N_3236,In_4955,In_3762);
nand U3237 (N_3237,In_2791,In_2191);
nand U3238 (N_3238,In_3715,In_1054);
nand U3239 (N_3239,In_2076,In_175);
xnor U3240 (N_3240,In_2324,In_1515);
and U3241 (N_3241,In_2398,In_1995);
xor U3242 (N_3242,In_2172,In_4356);
or U3243 (N_3243,In_3111,In_2519);
and U3244 (N_3244,In_3049,In_3666);
nor U3245 (N_3245,In_1223,In_1601);
nand U3246 (N_3246,In_4666,In_3876);
or U3247 (N_3247,In_3608,In_4456);
nand U3248 (N_3248,In_2383,In_4059);
and U3249 (N_3249,In_2681,In_645);
nor U3250 (N_3250,In_854,In_4432);
or U3251 (N_3251,In_767,In_3197);
and U3252 (N_3252,In_1124,In_1298);
or U3253 (N_3253,In_4011,In_372);
nand U3254 (N_3254,In_352,In_1756);
nand U3255 (N_3255,In_2381,In_2226);
nor U3256 (N_3256,In_4300,In_1065);
nand U3257 (N_3257,In_4865,In_1977);
nor U3258 (N_3258,In_1806,In_1969);
nor U3259 (N_3259,In_1238,In_565);
and U3260 (N_3260,In_1524,In_3753);
and U3261 (N_3261,In_185,In_3113);
nor U3262 (N_3262,In_1186,In_3096);
or U3263 (N_3263,In_1481,In_2909);
nor U3264 (N_3264,In_1453,In_809);
nand U3265 (N_3265,In_822,In_4772);
nand U3266 (N_3266,In_1468,In_68);
nor U3267 (N_3267,In_2265,In_654);
nand U3268 (N_3268,In_2269,In_1852);
nand U3269 (N_3269,In_1758,In_1322);
nand U3270 (N_3270,In_2734,In_2097);
nand U3271 (N_3271,In_1602,In_1799);
nor U3272 (N_3272,In_4227,In_1619);
and U3273 (N_3273,In_2786,In_2527);
or U3274 (N_3274,In_3706,In_985);
nor U3275 (N_3275,In_711,In_3225);
or U3276 (N_3276,In_3438,In_244);
or U3277 (N_3277,In_2909,In_2262);
xor U3278 (N_3278,In_465,In_1948);
and U3279 (N_3279,In_4912,In_3137);
nand U3280 (N_3280,In_4607,In_2185);
xor U3281 (N_3281,In_2977,In_44);
or U3282 (N_3282,In_1309,In_1808);
nor U3283 (N_3283,In_3771,In_1294);
xnor U3284 (N_3284,In_3325,In_3699);
nand U3285 (N_3285,In_4766,In_2226);
or U3286 (N_3286,In_1766,In_802);
or U3287 (N_3287,In_3835,In_2166);
xnor U3288 (N_3288,In_578,In_171);
nand U3289 (N_3289,In_4250,In_3215);
nand U3290 (N_3290,In_2122,In_476);
or U3291 (N_3291,In_112,In_4083);
nand U3292 (N_3292,In_2076,In_4432);
and U3293 (N_3293,In_3040,In_1745);
xor U3294 (N_3294,In_3694,In_492);
and U3295 (N_3295,In_2747,In_2708);
xor U3296 (N_3296,In_2869,In_4634);
nor U3297 (N_3297,In_166,In_3845);
or U3298 (N_3298,In_1270,In_1012);
nand U3299 (N_3299,In_2569,In_1780);
nand U3300 (N_3300,In_718,In_2522);
xnor U3301 (N_3301,In_3462,In_3694);
and U3302 (N_3302,In_864,In_4305);
xnor U3303 (N_3303,In_439,In_1555);
xnor U3304 (N_3304,In_4777,In_27);
or U3305 (N_3305,In_2017,In_4704);
xor U3306 (N_3306,In_4087,In_3469);
nand U3307 (N_3307,In_4836,In_4950);
xor U3308 (N_3308,In_1288,In_1727);
and U3309 (N_3309,In_3936,In_3587);
and U3310 (N_3310,In_2567,In_3736);
nand U3311 (N_3311,In_2071,In_3437);
xor U3312 (N_3312,In_94,In_3162);
nor U3313 (N_3313,In_4501,In_740);
or U3314 (N_3314,In_4039,In_3362);
xnor U3315 (N_3315,In_3910,In_1252);
and U3316 (N_3316,In_468,In_1840);
and U3317 (N_3317,In_2998,In_339);
and U3318 (N_3318,In_4337,In_696);
or U3319 (N_3319,In_4921,In_2546);
or U3320 (N_3320,In_3225,In_1329);
and U3321 (N_3321,In_1023,In_4831);
nand U3322 (N_3322,In_3418,In_4328);
and U3323 (N_3323,In_2108,In_1756);
nor U3324 (N_3324,In_4646,In_2815);
nand U3325 (N_3325,In_1615,In_71);
and U3326 (N_3326,In_3265,In_362);
nor U3327 (N_3327,In_627,In_709);
and U3328 (N_3328,In_2814,In_4859);
xor U3329 (N_3329,In_3933,In_2714);
and U3330 (N_3330,In_4019,In_2740);
nor U3331 (N_3331,In_4523,In_712);
xnor U3332 (N_3332,In_3557,In_696);
nand U3333 (N_3333,In_4854,In_2410);
or U3334 (N_3334,In_3442,In_4547);
or U3335 (N_3335,In_4169,In_3288);
nor U3336 (N_3336,In_2240,In_2879);
or U3337 (N_3337,In_322,In_2268);
or U3338 (N_3338,In_1640,In_2634);
xor U3339 (N_3339,In_2054,In_4907);
or U3340 (N_3340,In_957,In_2865);
or U3341 (N_3341,In_480,In_3891);
and U3342 (N_3342,In_4897,In_1180);
nor U3343 (N_3343,In_2901,In_788);
xor U3344 (N_3344,In_4780,In_2810);
or U3345 (N_3345,In_3106,In_4800);
and U3346 (N_3346,In_3077,In_3809);
or U3347 (N_3347,In_104,In_1833);
or U3348 (N_3348,In_2537,In_3067);
or U3349 (N_3349,In_3176,In_3783);
nand U3350 (N_3350,In_2709,In_4718);
and U3351 (N_3351,In_2879,In_864);
nand U3352 (N_3352,In_3690,In_486);
nor U3353 (N_3353,In_4454,In_502);
nor U3354 (N_3354,In_1086,In_3248);
and U3355 (N_3355,In_1788,In_3532);
or U3356 (N_3356,In_3768,In_4503);
or U3357 (N_3357,In_51,In_4168);
and U3358 (N_3358,In_4967,In_3967);
nor U3359 (N_3359,In_732,In_4611);
and U3360 (N_3360,In_1713,In_2056);
and U3361 (N_3361,In_2375,In_1416);
and U3362 (N_3362,In_749,In_3310);
and U3363 (N_3363,In_1610,In_2951);
or U3364 (N_3364,In_70,In_2484);
xor U3365 (N_3365,In_1392,In_4553);
and U3366 (N_3366,In_661,In_4082);
xnor U3367 (N_3367,In_4555,In_4578);
or U3368 (N_3368,In_3472,In_1845);
xor U3369 (N_3369,In_4096,In_1772);
nor U3370 (N_3370,In_4448,In_3730);
or U3371 (N_3371,In_21,In_889);
and U3372 (N_3372,In_1459,In_2327);
or U3373 (N_3373,In_1406,In_2667);
nor U3374 (N_3374,In_635,In_460);
and U3375 (N_3375,In_1607,In_3037);
and U3376 (N_3376,In_87,In_35);
xor U3377 (N_3377,In_3332,In_4976);
and U3378 (N_3378,In_4028,In_2576);
or U3379 (N_3379,In_2466,In_1196);
and U3380 (N_3380,In_4209,In_1630);
nand U3381 (N_3381,In_3213,In_3340);
or U3382 (N_3382,In_1249,In_4855);
nand U3383 (N_3383,In_3391,In_3539);
and U3384 (N_3384,In_2612,In_1361);
and U3385 (N_3385,In_3613,In_2568);
or U3386 (N_3386,In_4465,In_922);
nor U3387 (N_3387,In_4283,In_4282);
xor U3388 (N_3388,In_201,In_544);
and U3389 (N_3389,In_4353,In_3202);
and U3390 (N_3390,In_58,In_3322);
xnor U3391 (N_3391,In_2577,In_4079);
nand U3392 (N_3392,In_4530,In_4377);
and U3393 (N_3393,In_4210,In_1711);
nand U3394 (N_3394,In_3263,In_4491);
or U3395 (N_3395,In_2631,In_429);
nand U3396 (N_3396,In_2123,In_1615);
nand U3397 (N_3397,In_2913,In_4620);
xor U3398 (N_3398,In_1791,In_1664);
or U3399 (N_3399,In_444,In_2731);
nand U3400 (N_3400,In_967,In_901);
and U3401 (N_3401,In_2253,In_2136);
or U3402 (N_3402,In_2462,In_2668);
xor U3403 (N_3403,In_1816,In_3284);
xnor U3404 (N_3404,In_2668,In_326);
xor U3405 (N_3405,In_932,In_1889);
nand U3406 (N_3406,In_408,In_20);
nand U3407 (N_3407,In_4222,In_2830);
xnor U3408 (N_3408,In_3570,In_4191);
nor U3409 (N_3409,In_2178,In_1529);
nor U3410 (N_3410,In_247,In_3258);
and U3411 (N_3411,In_1660,In_2911);
or U3412 (N_3412,In_4172,In_2431);
and U3413 (N_3413,In_4148,In_3676);
nor U3414 (N_3414,In_635,In_3690);
nor U3415 (N_3415,In_4091,In_2983);
nor U3416 (N_3416,In_58,In_1719);
xnor U3417 (N_3417,In_457,In_2720);
xnor U3418 (N_3418,In_4078,In_1977);
nand U3419 (N_3419,In_4090,In_4156);
xor U3420 (N_3420,In_4220,In_4765);
and U3421 (N_3421,In_3668,In_3837);
nand U3422 (N_3422,In_4314,In_920);
nor U3423 (N_3423,In_4402,In_39);
xor U3424 (N_3424,In_4653,In_4919);
xnor U3425 (N_3425,In_3568,In_2152);
nand U3426 (N_3426,In_4115,In_4911);
nor U3427 (N_3427,In_1251,In_3539);
nor U3428 (N_3428,In_3326,In_4243);
nand U3429 (N_3429,In_2632,In_1278);
and U3430 (N_3430,In_2171,In_2738);
and U3431 (N_3431,In_2861,In_1862);
and U3432 (N_3432,In_3403,In_2229);
xor U3433 (N_3433,In_2382,In_2935);
nor U3434 (N_3434,In_4465,In_2487);
xnor U3435 (N_3435,In_1006,In_881);
and U3436 (N_3436,In_3304,In_2820);
nand U3437 (N_3437,In_1794,In_3843);
xor U3438 (N_3438,In_2833,In_4860);
nor U3439 (N_3439,In_4061,In_118);
nand U3440 (N_3440,In_4150,In_2759);
or U3441 (N_3441,In_72,In_4161);
nor U3442 (N_3442,In_3535,In_2146);
or U3443 (N_3443,In_2209,In_3586);
or U3444 (N_3444,In_2508,In_487);
xnor U3445 (N_3445,In_612,In_2807);
nand U3446 (N_3446,In_1418,In_189);
nand U3447 (N_3447,In_1996,In_2228);
nand U3448 (N_3448,In_1290,In_773);
nand U3449 (N_3449,In_4461,In_198);
nand U3450 (N_3450,In_1635,In_893);
or U3451 (N_3451,In_4821,In_1926);
or U3452 (N_3452,In_1924,In_3089);
or U3453 (N_3453,In_4490,In_3650);
and U3454 (N_3454,In_1211,In_1924);
xor U3455 (N_3455,In_2986,In_24);
and U3456 (N_3456,In_4566,In_1435);
nor U3457 (N_3457,In_2358,In_2388);
or U3458 (N_3458,In_1999,In_2123);
or U3459 (N_3459,In_2250,In_1536);
nor U3460 (N_3460,In_3220,In_1155);
or U3461 (N_3461,In_759,In_344);
xor U3462 (N_3462,In_888,In_2377);
and U3463 (N_3463,In_617,In_3182);
nand U3464 (N_3464,In_4244,In_558);
xor U3465 (N_3465,In_1743,In_2474);
nor U3466 (N_3466,In_3834,In_3489);
or U3467 (N_3467,In_774,In_2674);
and U3468 (N_3468,In_3412,In_2766);
or U3469 (N_3469,In_3174,In_3907);
nand U3470 (N_3470,In_1481,In_740);
or U3471 (N_3471,In_800,In_4728);
nor U3472 (N_3472,In_3821,In_2818);
and U3473 (N_3473,In_2871,In_606);
xor U3474 (N_3474,In_200,In_995);
xnor U3475 (N_3475,In_3873,In_3267);
and U3476 (N_3476,In_4432,In_4213);
nand U3477 (N_3477,In_3342,In_1159);
or U3478 (N_3478,In_922,In_3532);
xnor U3479 (N_3479,In_1023,In_4041);
or U3480 (N_3480,In_3542,In_2171);
and U3481 (N_3481,In_344,In_568);
nor U3482 (N_3482,In_1381,In_2249);
xnor U3483 (N_3483,In_2766,In_1870);
and U3484 (N_3484,In_2762,In_2650);
xnor U3485 (N_3485,In_870,In_4495);
nor U3486 (N_3486,In_233,In_4334);
nand U3487 (N_3487,In_1528,In_1511);
nor U3488 (N_3488,In_4269,In_3387);
nand U3489 (N_3489,In_4149,In_2912);
and U3490 (N_3490,In_23,In_3034);
or U3491 (N_3491,In_2614,In_4930);
xor U3492 (N_3492,In_3232,In_2923);
and U3493 (N_3493,In_199,In_1614);
nand U3494 (N_3494,In_2594,In_2627);
nand U3495 (N_3495,In_4191,In_1179);
nand U3496 (N_3496,In_1257,In_4763);
nand U3497 (N_3497,In_2229,In_202);
nand U3498 (N_3498,In_4924,In_1445);
xnor U3499 (N_3499,In_4975,In_3907);
and U3500 (N_3500,In_4081,In_4852);
nand U3501 (N_3501,In_4882,In_3352);
xnor U3502 (N_3502,In_2223,In_1010);
nor U3503 (N_3503,In_698,In_108);
nand U3504 (N_3504,In_412,In_1933);
and U3505 (N_3505,In_1098,In_1498);
xnor U3506 (N_3506,In_255,In_3009);
or U3507 (N_3507,In_4892,In_4543);
xor U3508 (N_3508,In_291,In_2732);
nor U3509 (N_3509,In_4851,In_2551);
nor U3510 (N_3510,In_3655,In_2123);
and U3511 (N_3511,In_4544,In_2999);
and U3512 (N_3512,In_988,In_981);
nand U3513 (N_3513,In_4725,In_1302);
nand U3514 (N_3514,In_960,In_1136);
xnor U3515 (N_3515,In_1096,In_3192);
nor U3516 (N_3516,In_2455,In_3091);
or U3517 (N_3517,In_4634,In_3258);
xor U3518 (N_3518,In_1733,In_3709);
xnor U3519 (N_3519,In_2066,In_26);
nor U3520 (N_3520,In_2093,In_2168);
or U3521 (N_3521,In_4608,In_2517);
and U3522 (N_3522,In_3790,In_3385);
nand U3523 (N_3523,In_4595,In_3458);
xnor U3524 (N_3524,In_3994,In_4031);
nand U3525 (N_3525,In_4632,In_4885);
nor U3526 (N_3526,In_2540,In_1537);
xor U3527 (N_3527,In_4236,In_4591);
nand U3528 (N_3528,In_3517,In_1028);
xor U3529 (N_3529,In_6,In_1674);
and U3530 (N_3530,In_2664,In_552);
nand U3531 (N_3531,In_4781,In_727);
xnor U3532 (N_3532,In_3683,In_4528);
nor U3533 (N_3533,In_2681,In_3895);
xor U3534 (N_3534,In_684,In_3029);
and U3535 (N_3535,In_3892,In_28);
or U3536 (N_3536,In_3802,In_4937);
xnor U3537 (N_3537,In_1386,In_1864);
and U3538 (N_3538,In_292,In_4041);
nand U3539 (N_3539,In_3189,In_2059);
xor U3540 (N_3540,In_1407,In_3952);
xnor U3541 (N_3541,In_2687,In_4153);
and U3542 (N_3542,In_1362,In_891);
or U3543 (N_3543,In_3552,In_3660);
xnor U3544 (N_3544,In_1413,In_888);
nor U3545 (N_3545,In_1414,In_3784);
nor U3546 (N_3546,In_3455,In_4813);
nand U3547 (N_3547,In_1832,In_4913);
xor U3548 (N_3548,In_730,In_3636);
and U3549 (N_3549,In_4549,In_1228);
xnor U3550 (N_3550,In_1662,In_724);
xnor U3551 (N_3551,In_4087,In_1108);
xnor U3552 (N_3552,In_2251,In_4821);
nand U3553 (N_3553,In_3465,In_4125);
xor U3554 (N_3554,In_2378,In_3096);
xor U3555 (N_3555,In_560,In_3);
nor U3556 (N_3556,In_4859,In_48);
xnor U3557 (N_3557,In_891,In_1927);
nor U3558 (N_3558,In_4586,In_4341);
and U3559 (N_3559,In_165,In_1328);
nor U3560 (N_3560,In_3835,In_2828);
nor U3561 (N_3561,In_403,In_443);
nor U3562 (N_3562,In_3354,In_3393);
or U3563 (N_3563,In_1545,In_2712);
xor U3564 (N_3564,In_4664,In_2066);
and U3565 (N_3565,In_2227,In_444);
xnor U3566 (N_3566,In_695,In_1233);
and U3567 (N_3567,In_3434,In_1212);
xor U3568 (N_3568,In_1094,In_922);
nand U3569 (N_3569,In_453,In_2128);
and U3570 (N_3570,In_4007,In_75);
nor U3571 (N_3571,In_2353,In_4505);
nand U3572 (N_3572,In_3736,In_1833);
nor U3573 (N_3573,In_1901,In_970);
nand U3574 (N_3574,In_4678,In_2714);
or U3575 (N_3575,In_3990,In_2525);
or U3576 (N_3576,In_4273,In_88);
nand U3577 (N_3577,In_1381,In_118);
nor U3578 (N_3578,In_4925,In_381);
xor U3579 (N_3579,In_1630,In_3412);
and U3580 (N_3580,In_945,In_1210);
or U3581 (N_3581,In_4659,In_4653);
and U3582 (N_3582,In_4476,In_1137);
or U3583 (N_3583,In_4684,In_831);
and U3584 (N_3584,In_560,In_3675);
xor U3585 (N_3585,In_943,In_3994);
xnor U3586 (N_3586,In_2791,In_3170);
or U3587 (N_3587,In_527,In_2472);
nand U3588 (N_3588,In_3926,In_4091);
or U3589 (N_3589,In_4777,In_2783);
or U3590 (N_3590,In_2677,In_4618);
nor U3591 (N_3591,In_4295,In_3253);
and U3592 (N_3592,In_4333,In_3193);
and U3593 (N_3593,In_4737,In_1037);
and U3594 (N_3594,In_1141,In_3472);
and U3595 (N_3595,In_3717,In_2645);
nor U3596 (N_3596,In_172,In_3835);
and U3597 (N_3597,In_4761,In_3127);
or U3598 (N_3598,In_2563,In_3318);
xnor U3599 (N_3599,In_3166,In_2895);
xor U3600 (N_3600,In_1096,In_2391);
nand U3601 (N_3601,In_3904,In_3453);
nor U3602 (N_3602,In_4493,In_3954);
or U3603 (N_3603,In_38,In_1997);
nand U3604 (N_3604,In_4732,In_3871);
and U3605 (N_3605,In_2145,In_1034);
nand U3606 (N_3606,In_174,In_2891);
xor U3607 (N_3607,In_3867,In_2427);
xnor U3608 (N_3608,In_2427,In_857);
nor U3609 (N_3609,In_4651,In_3005);
xnor U3610 (N_3610,In_4547,In_225);
nand U3611 (N_3611,In_1819,In_2425);
xor U3612 (N_3612,In_13,In_97);
or U3613 (N_3613,In_4406,In_2505);
nand U3614 (N_3614,In_3440,In_2898);
and U3615 (N_3615,In_2853,In_1304);
or U3616 (N_3616,In_2863,In_2552);
or U3617 (N_3617,In_1561,In_2420);
nor U3618 (N_3618,In_1674,In_439);
nor U3619 (N_3619,In_2570,In_2406);
nand U3620 (N_3620,In_1067,In_4772);
nor U3621 (N_3621,In_4782,In_1986);
and U3622 (N_3622,In_1850,In_886);
nor U3623 (N_3623,In_4491,In_3891);
or U3624 (N_3624,In_3854,In_3063);
xnor U3625 (N_3625,In_3825,In_4554);
nor U3626 (N_3626,In_585,In_450);
and U3627 (N_3627,In_4742,In_657);
or U3628 (N_3628,In_703,In_3567);
and U3629 (N_3629,In_3190,In_2157);
and U3630 (N_3630,In_301,In_3884);
nor U3631 (N_3631,In_3207,In_4227);
and U3632 (N_3632,In_1189,In_320);
xor U3633 (N_3633,In_4168,In_2744);
nor U3634 (N_3634,In_384,In_1613);
nor U3635 (N_3635,In_605,In_1779);
nand U3636 (N_3636,In_1404,In_1285);
nand U3637 (N_3637,In_1374,In_1747);
or U3638 (N_3638,In_4110,In_2080);
and U3639 (N_3639,In_809,In_2988);
nor U3640 (N_3640,In_3743,In_4917);
and U3641 (N_3641,In_2452,In_3846);
and U3642 (N_3642,In_2758,In_3036);
nor U3643 (N_3643,In_2511,In_3176);
xor U3644 (N_3644,In_3954,In_3323);
or U3645 (N_3645,In_866,In_3214);
or U3646 (N_3646,In_1618,In_1782);
nand U3647 (N_3647,In_3824,In_429);
nand U3648 (N_3648,In_4380,In_1212);
nand U3649 (N_3649,In_868,In_2377);
and U3650 (N_3650,In_1567,In_560);
nand U3651 (N_3651,In_4292,In_1445);
xnor U3652 (N_3652,In_3308,In_2626);
xnor U3653 (N_3653,In_2700,In_1616);
or U3654 (N_3654,In_4043,In_4897);
xnor U3655 (N_3655,In_4041,In_54);
nand U3656 (N_3656,In_4792,In_1042);
nor U3657 (N_3657,In_135,In_3283);
or U3658 (N_3658,In_381,In_1217);
nand U3659 (N_3659,In_3165,In_3916);
nor U3660 (N_3660,In_1001,In_2163);
nand U3661 (N_3661,In_3415,In_509);
or U3662 (N_3662,In_4408,In_3616);
or U3663 (N_3663,In_3533,In_1060);
or U3664 (N_3664,In_3057,In_517);
or U3665 (N_3665,In_1877,In_2553);
nor U3666 (N_3666,In_3816,In_2625);
nand U3667 (N_3667,In_2474,In_621);
xor U3668 (N_3668,In_4847,In_2213);
and U3669 (N_3669,In_563,In_1640);
nor U3670 (N_3670,In_4321,In_575);
or U3671 (N_3671,In_2497,In_1496);
xor U3672 (N_3672,In_2507,In_2889);
nor U3673 (N_3673,In_3271,In_4079);
nand U3674 (N_3674,In_3860,In_270);
nor U3675 (N_3675,In_3094,In_1141);
and U3676 (N_3676,In_3832,In_3397);
nand U3677 (N_3677,In_1779,In_529);
and U3678 (N_3678,In_3021,In_2495);
nand U3679 (N_3679,In_2793,In_3443);
xnor U3680 (N_3680,In_2551,In_4902);
nand U3681 (N_3681,In_396,In_2421);
or U3682 (N_3682,In_2282,In_4851);
nand U3683 (N_3683,In_2085,In_2020);
or U3684 (N_3684,In_3563,In_333);
or U3685 (N_3685,In_4904,In_3655);
nor U3686 (N_3686,In_4969,In_2338);
and U3687 (N_3687,In_1833,In_296);
nand U3688 (N_3688,In_3656,In_459);
xnor U3689 (N_3689,In_1388,In_1728);
nor U3690 (N_3690,In_2179,In_1110);
nor U3691 (N_3691,In_373,In_3112);
xor U3692 (N_3692,In_812,In_3901);
nor U3693 (N_3693,In_2800,In_540);
or U3694 (N_3694,In_2309,In_4147);
nand U3695 (N_3695,In_2671,In_757);
nor U3696 (N_3696,In_3809,In_456);
nor U3697 (N_3697,In_350,In_2936);
nor U3698 (N_3698,In_2277,In_3740);
nor U3699 (N_3699,In_1185,In_3371);
nor U3700 (N_3700,In_4272,In_2848);
nor U3701 (N_3701,In_2286,In_99);
and U3702 (N_3702,In_2955,In_2233);
nand U3703 (N_3703,In_1001,In_1354);
nand U3704 (N_3704,In_1300,In_272);
nand U3705 (N_3705,In_1718,In_3889);
or U3706 (N_3706,In_2410,In_2658);
or U3707 (N_3707,In_1881,In_3376);
nand U3708 (N_3708,In_713,In_3349);
xnor U3709 (N_3709,In_2123,In_1451);
xor U3710 (N_3710,In_2391,In_679);
or U3711 (N_3711,In_2308,In_1371);
nand U3712 (N_3712,In_2114,In_2484);
nor U3713 (N_3713,In_3930,In_4510);
nand U3714 (N_3714,In_988,In_783);
or U3715 (N_3715,In_3349,In_3148);
nand U3716 (N_3716,In_2406,In_2171);
nor U3717 (N_3717,In_319,In_97);
or U3718 (N_3718,In_2143,In_2772);
and U3719 (N_3719,In_3341,In_4625);
and U3720 (N_3720,In_1660,In_1093);
and U3721 (N_3721,In_4245,In_1403);
nor U3722 (N_3722,In_732,In_3207);
nand U3723 (N_3723,In_4018,In_3912);
nand U3724 (N_3724,In_3914,In_205);
nand U3725 (N_3725,In_2656,In_464);
or U3726 (N_3726,In_96,In_2070);
or U3727 (N_3727,In_798,In_4581);
xor U3728 (N_3728,In_3010,In_329);
nand U3729 (N_3729,In_3746,In_293);
nor U3730 (N_3730,In_3523,In_2232);
nand U3731 (N_3731,In_4936,In_1649);
xor U3732 (N_3732,In_3808,In_4359);
and U3733 (N_3733,In_1232,In_4660);
xor U3734 (N_3734,In_2880,In_3813);
xnor U3735 (N_3735,In_2213,In_3691);
xor U3736 (N_3736,In_4529,In_2162);
xnor U3737 (N_3737,In_4918,In_431);
nor U3738 (N_3738,In_1578,In_1230);
and U3739 (N_3739,In_3182,In_2547);
nor U3740 (N_3740,In_1242,In_1982);
and U3741 (N_3741,In_4209,In_1375);
nand U3742 (N_3742,In_2179,In_3573);
xnor U3743 (N_3743,In_3819,In_4403);
nand U3744 (N_3744,In_1521,In_4124);
nand U3745 (N_3745,In_1554,In_3058);
nor U3746 (N_3746,In_4079,In_2926);
and U3747 (N_3747,In_1662,In_992);
nand U3748 (N_3748,In_857,In_52);
and U3749 (N_3749,In_525,In_981);
or U3750 (N_3750,In_462,In_4249);
xor U3751 (N_3751,In_3836,In_915);
nor U3752 (N_3752,In_4181,In_3705);
or U3753 (N_3753,In_2078,In_2622);
and U3754 (N_3754,In_549,In_1805);
and U3755 (N_3755,In_2730,In_3498);
nand U3756 (N_3756,In_846,In_1478);
nor U3757 (N_3757,In_1716,In_4087);
nand U3758 (N_3758,In_2193,In_4501);
nand U3759 (N_3759,In_2689,In_2913);
nand U3760 (N_3760,In_243,In_4503);
nor U3761 (N_3761,In_2177,In_3773);
or U3762 (N_3762,In_845,In_169);
or U3763 (N_3763,In_2137,In_2622);
or U3764 (N_3764,In_265,In_2234);
and U3765 (N_3765,In_2928,In_2207);
or U3766 (N_3766,In_749,In_3015);
xnor U3767 (N_3767,In_1759,In_2140);
nand U3768 (N_3768,In_4473,In_708);
and U3769 (N_3769,In_1843,In_895);
or U3770 (N_3770,In_44,In_3303);
nand U3771 (N_3771,In_915,In_3217);
nand U3772 (N_3772,In_719,In_3461);
and U3773 (N_3773,In_469,In_1184);
or U3774 (N_3774,In_1461,In_1751);
nand U3775 (N_3775,In_3331,In_365);
or U3776 (N_3776,In_2046,In_4726);
and U3777 (N_3777,In_2986,In_1603);
nor U3778 (N_3778,In_2348,In_2650);
xor U3779 (N_3779,In_3748,In_1753);
nor U3780 (N_3780,In_3459,In_1615);
nor U3781 (N_3781,In_4435,In_4458);
and U3782 (N_3782,In_2575,In_3030);
xnor U3783 (N_3783,In_3857,In_272);
xnor U3784 (N_3784,In_1592,In_2098);
nor U3785 (N_3785,In_2829,In_1065);
or U3786 (N_3786,In_2864,In_3231);
nand U3787 (N_3787,In_1425,In_3421);
nor U3788 (N_3788,In_256,In_1434);
and U3789 (N_3789,In_4221,In_1157);
and U3790 (N_3790,In_2982,In_4493);
or U3791 (N_3791,In_3050,In_729);
nand U3792 (N_3792,In_1439,In_724);
xor U3793 (N_3793,In_1963,In_4617);
nand U3794 (N_3794,In_2577,In_1008);
or U3795 (N_3795,In_940,In_4417);
and U3796 (N_3796,In_1644,In_3322);
and U3797 (N_3797,In_3026,In_4965);
xor U3798 (N_3798,In_731,In_1284);
nand U3799 (N_3799,In_2206,In_1212);
or U3800 (N_3800,In_2792,In_1335);
nor U3801 (N_3801,In_695,In_207);
nand U3802 (N_3802,In_4647,In_1982);
and U3803 (N_3803,In_1377,In_3681);
and U3804 (N_3804,In_2450,In_1848);
nand U3805 (N_3805,In_4463,In_168);
nor U3806 (N_3806,In_4238,In_4351);
xor U3807 (N_3807,In_84,In_3898);
nor U3808 (N_3808,In_748,In_948);
xor U3809 (N_3809,In_3715,In_864);
nand U3810 (N_3810,In_1649,In_2039);
xnor U3811 (N_3811,In_3156,In_4155);
or U3812 (N_3812,In_2394,In_270);
nand U3813 (N_3813,In_2333,In_88);
or U3814 (N_3814,In_4182,In_1667);
nand U3815 (N_3815,In_348,In_2629);
nor U3816 (N_3816,In_2566,In_468);
nand U3817 (N_3817,In_4086,In_670);
nor U3818 (N_3818,In_3451,In_2209);
xnor U3819 (N_3819,In_823,In_4076);
and U3820 (N_3820,In_3599,In_2355);
nor U3821 (N_3821,In_770,In_3592);
nor U3822 (N_3822,In_1800,In_1865);
nor U3823 (N_3823,In_4946,In_576);
nand U3824 (N_3824,In_278,In_2029);
or U3825 (N_3825,In_4184,In_1952);
or U3826 (N_3826,In_133,In_2000);
nor U3827 (N_3827,In_4083,In_1673);
nor U3828 (N_3828,In_2952,In_4107);
xor U3829 (N_3829,In_1144,In_2913);
nor U3830 (N_3830,In_1976,In_3755);
xor U3831 (N_3831,In_246,In_3571);
nor U3832 (N_3832,In_1196,In_2066);
or U3833 (N_3833,In_2482,In_888);
or U3834 (N_3834,In_1299,In_2708);
nand U3835 (N_3835,In_2411,In_3474);
or U3836 (N_3836,In_3057,In_4283);
nor U3837 (N_3837,In_1971,In_1951);
and U3838 (N_3838,In_2930,In_2402);
and U3839 (N_3839,In_1395,In_400);
nor U3840 (N_3840,In_213,In_2169);
nand U3841 (N_3841,In_2950,In_4049);
or U3842 (N_3842,In_3645,In_3426);
or U3843 (N_3843,In_3491,In_4711);
nor U3844 (N_3844,In_1467,In_2639);
and U3845 (N_3845,In_4959,In_4675);
and U3846 (N_3846,In_2884,In_4797);
and U3847 (N_3847,In_994,In_2593);
nor U3848 (N_3848,In_4929,In_3606);
or U3849 (N_3849,In_392,In_1495);
xor U3850 (N_3850,In_728,In_569);
nand U3851 (N_3851,In_2413,In_3197);
nor U3852 (N_3852,In_334,In_3483);
nor U3853 (N_3853,In_3304,In_2150);
nor U3854 (N_3854,In_4480,In_4100);
nor U3855 (N_3855,In_1805,In_4099);
or U3856 (N_3856,In_4259,In_2384);
nor U3857 (N_3857,In_4124,In_723);
and U3858 (N_3858,In_3849,In_2101);
nand U3859 (N_3859,In_4672,In_3474);
nor U3860 (N_3860,In_629,In_2427);
nor U3861 (N_3861,In_2646,In_1845);
xnor U3862 (N_3862,In_1726,In_3217);
and U3863 (N_3863,In_3771,In_4684);
nand U3864 (N_3864,In_2802,In_4655);
nand U3865 (N_3865,In_2713,In_1747);
nand U3866 (N_3866,In_846,In_1226);
or U3867 (N_3867,In_3412,In_215);
or U3868 (N_3868,In_1613,In_547);
or U3869 (N_3869,In_1155,In_121);
and U3870 (N_3870,In_3721,In_3282);
and U3871 (N_3871,In_3855,In_953);
and U3872 (N_3872,In_3522,In_3763);
xor U3873 (N_3873,In_3260,In_3601);
and U3874 (N_3874,In_236,In_1053);
or U3875 (N_3875,In_1077,In_1624);
and U3876 (N_3876,In_422,In_4822);
and U3877 (N_3877,In_1158,In_1376);
and U3878 (N_3878,In_3474,In_3817);
nor U3879 (N_3879,In_3863,In_3720);
or U3880 (N_3880,In_313,In_4080);
nand U3881 (N_3881,In_266,In_4271);
xnor U3882 (N_3882,In_4035,In_4720);
and U3883 (N_3883,In_176,In_220);
and U3884 (N_3884,In_195,In_4241);
or U3885 (N_3885,In_4557,In_1648);
nor U3886 (N_3886,In_2766,In_3198);
and U3887 (N_3887,In_4428,In_492);
nor U3888 (N_3888,In_2751,In_931);
or U3889 (N_3889,In_3974,In_447);
xor U3890 (N_3890,In_720,In_946);
and U3891 (N_3891,In_480,In_3549);
and U3892 (N_3892,In_4340,In_3337);
xor U3893 (N_3893,In_1791,In_2823);
xor U3894 (N_3894,In_701,In_487);
nor U3895 (N_3895,In_2911,In_783);
nor U3896 (N_3896,In_3610,In_4386);
nand U3897 (N_3897,In_2185,In_4695);
or U3898 (N_3898,In_2879,In_452);
nand U3899 (N_3899,In_931,In_463);
or U3900 (N_3900,In_2740,In_2786);
or U3901 (N_3901,In_3658,In_2152);
and U3902 (N_3902,In_274,In_3432);
xnor U3903 (N_3903,In_3923,In_145);
or U3904 (N_3904,In_54,In_4625);
nor U3905 (N_3905,In_1783,In_1066);
and U3906 (N_3906,In_2861,In_4752);
and U3907 (N_3907,In_3428,In_257);
and U3908 (N_3908,In_4621,In_4769);
nor U3909 (N_3909,In_286,In_419);
and U3910 (N_3910,In_4341,In_3404);
and U3911 (N_3911,In_1212,In_2879);
nor U3912 (N_3912,In_3741,In_283);
nand U3913 (N_3913,In_2082,In_2058);
nand U3914 (N_3914,In_3893,In_4508);
or U3915 (N_3915,In_1574,In_1553);
or U3916 (N_3916,In_2606,In_3662);
nand U3917 (N_3917,In_3624,In_1434);
xor U3918 (N_3918,In_2115,In_785);
and U3919 (N_3919,In_1977,In_1855);
nor U3920 (N_3920,In_2255,In_2816);
xnor U3921 (N_3921,In_894,In_4978);
nor U3922 (N_3922,In_4036,In_937);
or U3923 (N_3923,In_2349,In_3802);
xor U3924 (N_3924,In_4329,In_4417);
nor U3925 (N_3925,In_2821,In_194);
or U3926 (N_3926,In_2750,In_3150);
nor U3927 (N_3927,In_2454,In_2193);
xnor U3928 (N_3928,In_1137,In_1300);
and U3929 (N_3929,In_3069,In_1257);
xnor U3930 (N_3930,In_1809,In_2458);
nand U3931 (N_3931,In_4476,In_208);
nor U3932 (N_3932,In_2796,In_1739);
xor U3933 (N_3933,In_231,In_1671);
or U3934 (N_3934,In_4164,In_2105);
nor U3935 (N_3935,In_2208,In_4673);
or U3936 (N_3936,In_4683,In_1488);
or U3937 (N_3937,In_169,In_4728);
nor U3938 (N_3938,In_1835,In_4429);
xor U3939 (N_3939,In_1855,In_2074);
nor U3940 (N_3940,In_4028,In_4921);
or U3941 (N_3941,In_1886,In_2362);
xor U3942 (N_3942,In_4610,In_2659);
or U3943 (N_3943,In_1975,In_3271);
xnor U3944 (N_3944,In_679,In_2420);
and U3945 (N_3945,In_3995,In_859);
xor U3946 (N_3946,In_2879,In_3873);
xnor U3947 (N_3947,In_4232,In_4857);
xnor U3948 (N_3948,In_3474,In_2804);
or U3949 (N_3949,In_4827,In_1543);
and U3950 (N_3950,In_4884,In_3177);
nor U3951 (N_3951,In_4312,In_3937);
and U3952 (N_3952,In_4643,In_3814);
nand U3953 (N_3953,In_1193,In_1951);
or U3954 (N_3954,In_599,In_1634);
xor U3955 (N_3955,In_3118,In_1514);
and U3956 (N_3956,In_420,In_2562);
nand U3957 (N_3957,In_170,In_4650);
nand U3958 (N_3958,In_3380,In_1225);
nor U3959 (N_3959,In_3022,In_3653);
xor U3960 (N_3960,In_1948,In_195);
or U3961 (N_3961,In_4319,In_2993);
xor U3962 (N_3962,In_4238,In_1962);
or U3963 (N_3963,In_1747,In_2830);
nor U3964 (N_3964,In_4689,In_4461);
or U3965 (N_3965,In_4467,In_3311);
nand U3966 (N_3966,In_3388,In_4228);
nand U3967 (N_3967,In_994,In_901);
and U3968 (N_3968,In_2647,In_652);
nor U3969 (N_3969,In_1241,In_108);
or U3970 (N_3970,In_1804,In_488);
xor U3971 (N_3971,In_929,In_4264);
and U3972 (N_3972,In_4331,In_4925);
xor U3973 (N_3973,In_3085,In_1521);
xnor U3974 (N_3974,In_2477,In_1067);
nor U3975 (N_3975,In_4296,In_428);
nor U3976 (N_3976,In_2253,In_802);
xor U3977 (N_3977,In_131,In_4982);
or U3978 (N_3978,In_2401,In_3332);
and U3979 (N_3979,In_4962,In_91);
nor U3980 (N_3980,In_2908,In_4591);
and U3981 (N_3981,In_2865,In_481);
nand U3982 (N_3982,In_1989,In_4158);
or U3983 (N_3983,In_321,In_1472);
or U3984 (N_3984,In_1606,In_535);
xor U3985 (N_3985,In_1501,In_4437);
nand U3986 (N_3986,In_4853,In_1265);
nor U3987 (N_3987,In_790,In_3238);
nand U3988 (N_3988,In_2975,In_1742);
or U3989 (N_3989,In_3789,In_883);
nor U3990 (N_3990,In_3620,In_934);
and U3991 (N_3991,In_1341,In_254);
xor U3992 (N_3992,In_2157,In_613);
or U3993 (N_3993,In_3676,In_1881);
or U3994 (N_3994,In_2407,In_3976);
and U3995 (N_3995,In_2163,In_542);
xnor U3996 (N_3996,In_4050,In_2296);
nand U3997 (N_3997,In_1260,In_4803);
and U3998 (N_3998,In_3886,In_3545);
or U3999 (N_3999,In_4429,In_4930);
nand U4000 (N_4000,In_2336,In_2681);
or U4001 (N_4001,In_2215,In_1983);
and U4002 (N_4002,In_1417,In_3917);
or U4003 (N_4003,In_2133,In_4321);
xnor U4004 (N_4004,In_4531,In_4543);
or U4005 (N_4005,In_3261,In_2063);
and U4006 (N_4006,In_4056,In_1382);
nand U4007 (N_4007,In_3356,In_1474);
nand U4008 (N_4008,In_3620,In_4900);
xnor U4009 (N_4009,In_2596,In_3326);
or U4010 (N_4010,In_630,In_3516);
xnor U4011 (N_4011,In_4006,In_130);
nand U4012 (N_4012,In_3262,In_1430);
nor U4013 (N_4013,In_870,In_3033);
and U4014 (N_4014,In_2478,In_3661);
nand U4015 (N_4015,In_560,In_716);
nor U4016 (N_4016,In_847,In_1555);
xnor U4017 (N_4017,In_4680,In_178);
nand U4018 (N_4018,In_4829,In_2233);
or U4019 (N_4019,In_4378,In_4975);
nor U4020 (N_4020,In_992,In_330);
xnor U4021 (N_4021,In_1017,In_1621);
or U4022 (N_4022,In_1429,In_195);
nand U4023 (N_4023,In_3086,In_4788);
nor U4024 (N_4024,In_3741,In_4564);
nor U4025 (N_4025,In_3025,In_2547);
nand U4026 (N_4026,In_3899,In_4903);
and U4027 (N_4027,In_490,In_898);
and U4028 (N_4028,In_2160,In_656);
or U4029 (N_4029,In_2033,In_4951);
nor U4030 (N_4030,In_1605,In_754);
and U4031 (N_4031,In_4190,In_726);
nand U4032 (N_4032,In_3185,In_2596);
nor U4033 (N_4033,In_2681,In_4638);
nand U4034 (N_4034,In_1897,In_1097);
nand U4035 (N_4035,In_3345,In_1164);
xnor U4036 (N_4036,In_3855,In_212);
or U4037 (N_4037,In_1863,In_72);
or U4038 (N_4038,In_3724,In_4950);
xnor U4039 (N_4039,In_4087,In_167);
and U4040 (N_4040,In_881,In_1514);
and U4041 (N_4041,In_2283,In_2369);
nor U4042 (N_4042,In_1900,In_1990);
xnor U4043 (N_4043,In_2062,In_1386);
xnor U4044 (N_4044,In_3539,In_4021);
or U4045 (N_4045,In_1616,In_554);
or U4046 (N_4046,In_1658,In_4767);
xnor U4047 (N_4047,In_307,In_2675);
and U4048 (N_4048,In_4565,In_2327);
and U4049 (N_4049,In_2356,In_2926);
nand U4050 (N_4050,In_968,In_174);
xor U4051 (N_4051,In_4428,In_4622);
xor U4052 (N_4052,In_455,In_4375);
and U4053 (N_4053,In_2150,In_2409);
and U4054 (N_4054,In_832,In_2671);
and U4055 (N_4055,In_1426,In_523);
xor U4056 (N_4056,In_441,In_4569);
nor U4057 (N_4057,In_2959,In_3469);
and U4058 (N_4058,In_2919,In_262);
nor U4059 (N_4059,In_3904,In_2356);
or U4060 (N_4060,In_2469,In_4802);
xnor U4061 (N_4061,In_2808,In_4377);
or U4062 (N_4062,In_3210,In_926);
nor U4063 (N_4063,In_1927,In_800);
xnor U4064 (N_4064,In_2560,In_3464);
nor U4065 (N_4065,In_1395,In_248);
xnor U4066 (N_4066,In_3152,In_4360);
xnor U4067 (N_4067,In_3764,In_2284);
and U4068 (N_4068,In_2017,In_1563);
xor U4069 (N_4069,In_537,In_99);
xnor U4070 (N_4070,In_2369,In_2169);
xor U4071 (N_4071,In_1939,In_2901);
and U4072 (N_4072,In_1084,In_3550);
nor U4073 (N_4073,In_1470,In_4986);
nor U4074 (N_4074,In_4975,In_2355);
or U4075 (N_4075,In_3069,In_2211);
or U4076 (N_4076,In_4184,In_131);
or U4077 (N_4077,In_3610,In_1190);
xor U4078 (N_4078,In_2718,In_276);
or U4079 (N_4079,In_4257,In_1223);
and U4080 (N_4080,In_3584,In_4841);
xnor U4081 (N_4081,In_3297,In_1936);
xor U4082 (N_4082,In_2516,In_1091);
and U4083 (N_4083,In_2676,In_1590);
nor U4084 (N_4084,In_2001,In_1926);
nor U4085 (N_4085,In_4142,In_143);
or U4086 (N_4086,In_2944,In_4055);
nand U4087 (N_4087,In_2980,In_2332);
nand U4088 (N_4088,In_360,In_2111);
xor U4089 (N_4089,In_4595,In_1312);
or U4090 (N_4090,In_1125,In_1049);
or U4091 (N_4091,In_3189,In_772);
or U4092 (N_4092,In_3453,In_2533);
nand U4093 (N_4093,In_1875,In_2220);
xnor U4094 (N_4094,In_2820,In_370);
and U4095 (N_4095,In_3945,In_1947);
and U4096 (N_4096,In_733,In_4835);
and U4097 (N_4097,In_2973,In_63);
nand U4098 (N_4098,In_2513,In_607);
or U4099 (N_4099,In_1651,In_1943);
xnor U4100 (N_4100,In_332,In_1360);
nor U4101 (N_4101,In_1487,In_3442);
and U4102 (N_4102,In_392,In_4947);
and U4103 (N_4103,In_4174,In_2359);
nand U4104 (N_4104,In_3876,In_4546);
and U4105 (N_4105,In_17,In_1769);
and U4106 (N_4106,In_3966,In_698);
or U4107 (N_4107,In_4586,In_2730);
nor U4108 (N_4108,In_4098,In_3544);
nand U4109 (N_4109,In_3765,In_3449);
or U4110 (N_4110,In_3116,In_3655);
or U4111 (N_4111,In_3458,In_1921);
and U4112 (N_4112,In_2135,In_528);
and U4113 (N_4113,In_3499,In_3785);
nand U4114 (N_4114,In_4586,In_3075);
nor U4115 (N_4115,In_368,In_697);
or U4116 (N_4116,In_3570,In_3052);
or U4117 (N_4117,In_4668,In_3647);
and U4118 (N_4118,In_4281,In_4598);
xor U4119 (N_4119,In_1521,In_53);
nand U4120 (N_4120,In_1871,In_2545);
nor U4121 (N_4121,In_503,In_1498);
or U4122 (N_4122,In_1704,In_3563);
nand U4123 (N_4123,In_2459,In_1867);
or U4124 (N_4124,In_2844,In_1057);
and U4125 (N_4125,In_1544,In_1547);
nor U4126 (N_4126,In_3974,In_2772);
nor U4127 (N_4127,In_2126,In_2497);
xor U4128 (N_4128,In_2350,In_4582);
or U4129 (N_4129,In_1776,In_1247);
nand U4130 (N_4130,In_1279,In_1202);
nand U4131 (N_4131,In_3689,In_2616);
nor U4132 (N_4132,In_4603,In_4602);
xnor U4133 (N_4133,In_470,In_2692);
or U4134 (N_4134,In_1973,In_3368);
or U4135 (N_4135,In_1621,In_2888);
xnor U4136 (N_4136,In_1125,In_1646);
nor U4137 (N_4137,In_3418,In_1592);
xnor U4138 (N_4138,In_1426,In_4344);
nor U4139 (N_4139,In_2428,In_3438);
and U4140 (N_4140,In_3239,In_3902);
nor U4141 (N_4141,In_4378,In_4683);
and U4142 (N_4142,In_4086,In_3704);
and U4143 (N_4143,In_975,In_897);
nand U4144 (N_4144,In_2347,In_3769);
or U4145 (N_4145,In_4037,In_14);
xnor U4146 (N_4146,In_1703,In_1181);
xnor U4147 (N_4147,In_2772,In_3937);
nor U4148 (N_4148,In_613,In_357);
nand U4149 (N_4149,In_1898,In_4177);
xor U4150 (N_4150,In_38,In_3795);
xor U4151 (N_4151,In_1590,In_3214);
nor U4152 (N_4152,In_4681,In_1284);
or U4153 (N_4153,In_2514,In_4962);
xnor U4154 (N_4154,In_3193,In_1652);
and U4155 (N_4155,In_4535,In_974);
and U4156 (N_4156,In_1525,In_4828);
xor U4157 (N_4157,In_3063,In_2380);
nor U4158 (N_4158,In_3634,In_2177);
or U4159 (N_4159,In_3689,In_3064);
nand U4160 (N_4160,In_3239,In_992);
nand U4161 (N_4161,In_805,In_274);
nor U4162 (N_4162,In_4979,In_1147);
nand U4163 (N_4163,In_3678,In_1180);
xnor U4164 (N_4164,In_4560,In_3414);
nand U4165 (N_4165,In_1132,In_395);
xnor U4166 (N_4166,In_669,In_388);
and U4167 (N_4167,In_4714,In_923);
nor U4168 (N_4168,In_759,In_1615);
nand U4169 (N_4169,In_1963,In_455);
and U4170 (N_4170,In_852,In_136);
nor U4171 (N_4171,In_4774,In_1607);
nand U4172 (N_4172,In_1844,In_1377);
and U4173 (N_4173,In_3335,In_2692);
xnor U4174 (N_4174,In_648,In_872);
and U4175 (N_4175,In_3980,In_1115);
xnor U4176 (N_4176,In_3517,In_1067);
and U4177 (N_4177,In_4040,In_1377);
xor U4178 (N_4178,In_1858,In_4060);
xor U4179 (N_4179,In_2401,In_1444);
and U4180 (N_4180,In_1711,In_3562);
nand U4181 (N_4181,In_4715,In_842);
and U4182 (N_4182,In_1285,In_1701);
and U4183 (N_4183,In_3107,In_1021);
nor U4184 (N_4184,In_4205,In_4617);
or U4185 (N_4185,In_2204,In_701);
and U4186 (N_4186,In_271,In_1375);
nor U4187 (N_4187,In_1725,In_4086);
nor U4188 (N_4188,In_2831,In_790);
and U4189 (N_4189,In_4026,In_4103);
nand U4190 (N_4190,In_3119,In_381);
and U4191 (N_4191,In_3359,In_4725);
and U4192 (N_4192,In_345,In_3747);
xnor U4193 (N_4193,In_3072,In_1599);
xnor U4194 (N_4194,In_1093,In_859);
xnor U4195 (N_4195,In_2336,In_537);
and U4196 (N_4196,In_296,In_2424);
xnor U4197 (N_4197,In_725,In_4159);
or U4198 (N_4198,In_4046,In_3179);
nor U4199 (N_4199,In_3202,In_2288);
nor U4200 (N_4200,In_517,In_4189);
nor U4201 (N_4201,In_3955,In_3712);
and U4202 (N_4202,In_4226,In_2974);
or U4203 (N_4203,In_3431,In_4082);
or U4204 (N_4204,In_1070,In_2177);
or U4205 (N_4205,In_3390,In_853);
xnor U4206 (N_4206,In_864,In_37);
nor U4207 (N_4207,In_4181,In_3813);
nand U4208 (N_4208,In_2096,In_1764);
or U4209 (N_4209,In_349,In_4103);
and U4210 (N_4210,In_1596,In_579);
nor U4211 (N_4211,In_1929,In_2319);
nand U4212 (N_4212,In_2433,In_3372);
xnor U4213 (N_4213,In_983,In_4637);
or U4214 (N_4214,In_280,In_3519);
xor U4215 (N_4215,In_1104,In_734);
or U4216 (N_4216,In_555,In_1137);
nand U4217 (N_4217,In_332,In_77);
nor U4218 (N_4218,In_2111,In_1841);
nand U4219 (N_4219,In_3944,In_4638);
xor U4220 (N_4220,In_2665,In_4514);
or U4221 (N_4221,In_2833,In_3141);
nand U4222 (N_4222,In_4222,In_121);
nor U4223 (N_4223,In_2121,In_3234);
and U4224 (N_4224,In_778,In_4460);
and U4225 (N_4225,In_2448,In_1336);
and U4226 (N_4226,In_300,In_1658);
and U4227 (N_4227,In_3295,In_635);
and U4228 (N_4228,In_1544,In_2859);
or U4229 (N_4229,In_2790,In_1626);
nor U4230 (N_4230,In_4049,In_4876);
or U4231 (N_4231,In_4753,In_3154);
nand U4232 (N_4232,In_582,In_4734);
and U4233 (N_4233,In_1663,In_84);
nand U4234 (N_4234,In_3722,In_2426);
xnor U4235 (N_4235,In_541,In_4335);
nor U4236 (N_4236,In_2554,In_2979);
xnor U4237 (N_4237,In_2653,In_4123);
nand U4238 (N_4238,In_3158,In_4727);
nor U4239 (N_4239,In_3768,In_4013);
nor U4240 (N_4240,In_752,In_3503);
nand U4241 (N_4241,In_2308,In_2942);
or U4242 (N_4242,In_162,In_4735);
nand U4243 (N_4243,In_42,In_4257);
xor U4244 (N_4244,In_1279,In_4909);
nand U4245 (N_4245,In_3566,In_1205);
nor U4246 (N_4246,In_1525,In_4357);
xor U4247 (N_4247,In_14,In_4333);
nand U4248 (N_4248,In_2580,In_2445);
or U4249 (N_4249,In_1914,In_1461);
or U4250 (N_4250,In_3931,In_3522);
nor U4251 (N_4251,In_1738,In_1647);
and U4252 (N_4252,In_1506,In_4093);
xor U4253 (N_4253,In_3734,In_477);
xnor U4254 (N_4254,In_1230,In_1726);
and U4255 (N_4255,In_1100,In_3760);
nor U4256 (N_4256,In_4869,In_3716);
and U4257 (N_4257,In_3672,In_2672);
nand U4258 (N_4258,In_3707,In_4554);
xnor U4259 (N_4259,In_929,In_464);
xnor U4260 (N_4260,In_4731,In_1591);
or U4261 (N_4261,In_2207,In_302);
nor U4262 (N_4262,In_976,In_4026);
xor U4263 (N_4263,In_2772,In_4431);
xor U4264 (N_4264,In_4401,In_4165);
nand U4265 (N_4265,In_868,In_2705);
nand U4266 (N_4266,In_2441,In_4153);
xnor U4267 (N_4267,In_1899,In_2885);
nor U4268 (N_4268,In_4023,In_1480);
xor U4269 (N_4269,In_2272,In_576);
xor U4270 (N_4270,In_1682,In_4892);
nand U4271 (N_4271,In_1490,In_50);
nor U4272 (N_4272,In_3768,In_722);
or U4273 (N_4273,In_156,In_4350);
nand U4274 (N_4274,In_4236,In_4465);
and U4275 (N_4275,In_585,In_2166);
xnor U4276 (N_4276,In_3682,In_2867);
nor U4277 (N_4277,In_400,In_2592);
or U4278 (N_4278,In_2096,In_3723);
and U4279 (N_4279,In_1524,In_4992);
nand U4280 (N_4280,In_4310,In_4844);
nor U4281 (N_4281,In_1036,In_2062);
nand U4282 (N_4282,In_1593,In_230);
xnor U4283 (N_4283,In_2899,In_4952);
nor U4284 (N_4284,In_1392,In_4373);
nand U4285 (N_4285,In_1115,In_4848);
xor U4286 (N_4286,In_2638,In_180);
xnor U4287 (N_4287,In_3295,In_2918);
xor U4288 (N_4288,In_2910,In_850);
and U4289 (N_4289,In_3774,In_1525);
and U4290 (N_4290,In_422,In_521);
nand U4291 (N_4291,In_3644,In_3871);
xnor U4292 (N_4292,In_1717,In_2079);
or U4293 (N_4293,In_160,In_4797);
nand U4294 (N_4294,In_2462,In_4954);
nor U4295 (N_4295,In_1693,In_2992);
nor U4296 (N_4296,In_3677,In_3419);
nand U4297 (N_4297,In_1916,In_815);
and U4298 (N_4298,In_3039,In_4748);
and U4299 (N_4299,In_81,In_3027);
and U4300 (N_4300,In_3862,In_1014);
and U4301 (N_4301,In_1527,In_4417);
nor U4302 (N_4302,In_3707,In_3702);
nand U4303 (N_4303,In_2109,In_3519);
or U4304 (N_4304,In_4564,In_674);
xor U4305 (N_4305,In_958,In_1237);
xnor U4306 (N_4306,In_2527,In_4226);
nand U4307 (N_4307,In_1279,In_2192);
nor U4308 (N_4308,In_2296,In_2177);
and U4309 (N_4309,In_2770,In_3729);
and U4310 (N_4310,In_2059,In_2193);
nor U4311 (N_4311,In_1655,In_4509);
nand U4312 (N_4312,In_4623,In_3465);
nand U4313 (N_4313,In_4064,In_4962);
nand U4314 (N_4314,In_319,In_1318);
nand U4315 (N_4315,In_4320,In_3097);
and U4316 (N_4316,In_4565,In_2970);
nand U4317 (N_4317,In_2487,In_1505);
or U4318 (N_4318,In_3850,In_2354);
and U4319 (N_4319,In_4149,In_860);
or U4320 (N_4320,In_985,In_3871);
xnor U4321 (N_4321,In_4224,In_3247);
or U4322 (N_4322,In_2735,In_1362);
xnor U4323 (N_4323,In_1928,In_2345);
nor U4324 (N_4324,In_4307,In_4205);
nand U4325 (N_4325,In_2165,In_4222);
nor U4326 (N_4326,In_2021,In_1147);
and U4327 (N_4327,In_3364,In_1528);
xnor U4328 (N_4328,In_3756,In_3081);
nor U4329 (N_4329,In_2976,In_2694);
nor U4330 (N_4330,In_754,In_4482);
nand U4331 (N_4331,In_10,In_3921);
and U4332 (N_4332,In_3210,In_4211);
or U4333 (N_4333,In_4658,In_3755);
xor U4334 (N_4334,In_2895,In_3430);
xnor U4335 (N_4335,In_2181,In_4477);
nor U4336 (N_4336,In_1368,In_4445);
nor U4337 (N_4337,In_3856,In_3909);
and U4338 (N_4338,In_2516,In_276);
xnor U4339 (N_4339,In_1286,In_1802);
and U4340 (N_4340,In_1589,In_2023);
xor U4341 (N_4341,In_2568,In_1684);
xor U4342 (N_4342,In_4863,In_4244);
nand U4343 (N_4343,In_4338,In_496);
nand U4344 (N_4344,In_2322,In_355);
xnor U4345 (N_4345,In_4347,In_368);
or U4346 (N_4346,In_2282,In_242);
or U4347 (N_4347,In_2729,In_4538);
and U4348 (N_4348,In_2942,In_2810);
and U4349 (N_4349,In_315,In_2196);
nor U4350 (N_4350,In_272,In_3881);
nor U4351 (N_4351,In_1682,In_3683);
xnor U4352 (N_4352,In_171,In_4283);
nor U4353 (N_4353,In_3574,In_4258);
nand U4354 (N_4354,In_2857,In_3381);
nand U4355 (N_4355,In_3632,In_4340);
and U4356 (N_4356,In_1066,In_4611);
xnor U4357 (N_4357,In_4761,In_797);
nor U4358 (N_4358,In_1720,In_1104);
nand U4359 (N_4359,In_4397,In_4014);
and U4360 (N_4360,In_3755,In_2249);
nor U4361 (N_4361,In_2931,In_1745);
nand U4362 (N_4362,In_779,In_4757);
nor U4363 (N_4363,In_4123,In_501);
nor U4364 (N_4364,In_2062,In_2303);
nor U4365 (N_4365,In_1175,In_2873);
nor U4366 (N_4366,In_2880,In_4856);
xnor U4367 (N_4367,In_4195,In_1258);
and U4368 (N_4368,In_3332,In_2908);
nor U4369 (N_4369,In_3618,In_2458);
xor U4370 (N_4370,In_3893,In_4664);
or U4371 (N_4371,In_4201,In_4174);
or U4372 (N_4372,In_3249,In_948);
nor U4373 (N_4373,In_2264,In_3940);
or U4374 (N_4374,In_2494,In_2967);
xor U4375 (N_4375,In_2998,In_3189);
or U4376 (N_4376,In_2918,In_3508);
or U4377 (N_4377,In_3767,In_3189);
and U4378 (N_4378,In_3161,In_316);
xnor U4379 (N_4379,In_2738,In_2308);
or U4380 (N_4380,In_1032,In_1442);
or U4381 (N_4381,In_4129,In_3065);
or U4382 (N_4382,In_55,In_674);
xnor U4383 (N_4383,In_3255,In_338);
or U4384 (N_4384,In_3205,In_2537);
and U4385 (N_4385,In_3015,In_1337);
and U4386 (N_4386,In_324,In_4680);
nor U4387 (N_4387,In_4835,In_1717);
nand U4388 (N_4388,In_125,In_3946);
nor U4389 (N_4389,In_3206,In_3449);
nor U4390 (N_4390,In_527,In_1655);
xor U4391 (N_4391,In_3932,In_3446);
nand U4392 (N_4392,In_2974,In_4114);
nand U4393 (N_4393,In_169,In_4504);
and U4394 (N_4394,In_3121,In_2958);
xnor U4395 (N_4395,In_315,In_2278);
nand U4396 (N_4396,In_762,In_3923);
nor U4397 (N_4397,In_3035,In_967);
or U4398 (N_4398,In_4731,In_3034);
xnor U4399 (N_4399,In_1775,In_4467);
or U4400 (N_4400,In_2126,In_4283);
and U4401 (N_4401,In_4904,In_3463);
nand U4402 (N_4402,In_2236,In_4453);
and U4403 (N_4403,In_1711,In_740);
nor U4404 (N_4404,In_1256,In_1707);
nor U4405 (N_4405,In_2815,In_3995);
or U4406 (N_4406,In_4734,In_3206);
or U4407 (N_4407,In_2040,In_2392);
and U4408 (N_4408,In_4756,In_124);
and U4409 (N_4409,In_2181,In_3829);
xor U4410 (N_4410,In_4354,In_4945);
or U4411 (N_4411,In_3196,In_2148);
nor U4412 (N_4412,In_669,In_4978);
nand U4413 (N_4413,In_4451,In_3445);
or U4414 (N_4414,In_3064,In_4380);
and U4415 (N_4415,In_970,In_1090);
nand U4416 (N_4416,In_1518,In_366);
nor U4417 (N_4417,In_2015,In_1178);
xnor U4418 (N_4418,In_4064,In_2525);
nor U4419 (N_4419,In_2352,In_814);
nor U4420 (N_4420,In_4273,In_1127);
or U4421 (N_4421,In_3506,In_3706);
xor U4422 (N_4422,In_3512,In_4888);
xor U4423 (N_4423,In_4292,In_1709);
xnor U4424 (N_4424,In_2442,In_4089);
xor U4425 (N_4425,In_3513,In_557);
nand U4426 (N_4426,In_4690,In_3508);
and U4427 (N_4427,In_4976,In_1764);
xor U4428 (N_4428,In_1161,In_3374);
nand U4429 (N_4429,In_4410,In_2989);
or U4430 (N_4430,In_2875,In_2308);
nand U4431 (N_4431,In_1098,In_1572);
or U4432 (N_4432,In_4100,In_1504);
or U4433 (N_4433,In_4768,In_3258);
and U4434 (N_4434,In_2089,In_2826);
and U4435 (N_4435,In_4450,In_46);
xor U4436 (N_4436,In_3016,In_1);
or U4437 (N_4437,In_2932,In_2083);
nor U4438 (N_4438,In_305,In_2243);
nor U4439 (N_4439,In_4950,In_2616);
nand U4440 (N_4440,In_2484,In_3561);
nor U4441 (N_4441,In_3593,In_2700);
and U4442 (N_4442,In_2362,In_3649);
xor U4443 (N_4443,In_39,In_4244);
and U4444 (N_4444,In_3208,In_3479);
nand U4445 (N_4445,In_2860,In_976);
nor U4446 (N_4446,In_2910,In_755);
and U4447 (N_4447,In_1193,In_1933);
nor U4448 (N_4448,In_4558,In_935);
xnor U4449 (N_4449,In_2087,In_4455);
nand U4450 (N_4450,In_3616,In_4044);
nand U4451 (N_4451,In_1284,In_2007);
xor U4452 (N_4452,In_876,In_1130);
nor U4453 (N_4453,In_2042,In_2180);
nand U4454 (N_4454,In_4798,In_3404);
nand U4455 (N_4455,In_391,In_3545);
or U4456 (N_4456,In_591,In_2330);
nor U4457 (N_4457,In_1021,In_3257);
xnor U4458 (N_4458,In_1481,In_1449);
or U4459 (N_4459,In_730,In_3785);
nand U4460 (N_4460,In_4876,In_784);
nand U4461 (N_4461,In_2886,In_4769);
and U4462 (N_4462,In_4770,In_1229);
xnor U4463 (N_4463,In_532,In_2866);
and U4464 (N_4464,In_485,In_4717);
xnor U4465 (N_4465,In_3338,In_4538);
xor U4466 (N_4466,In_4810,In_944);
nor U4467 (N_4467,In_526,In_4265);
nand U4468 (N_4468,In_361,In_4751);
and U4469 (N_4469,In_653,In_3087);
and U4470 (N_4470,In_4111,In_3013);
nor U4471 (N_4471,In_1986,In_496);
and U4472 (N_4472,In_549,In_3897);
or U4473 (N_4473,In_2681,In_2456);
xor U4474 (N_4474,In_1485,In_2043);
nor U4475 (N_4475,In_3702,In_3658);
or U4476 (N_4476,In_4937,In_3223);
nand U4477 (N_4477,In_3385,In_1201);
xor U4478 (N_4478,In_10,In_4988);
and U4479 (N_4479,In_4614,In_3780);
and U4480 (N_4480,In_1019,In_97);
or U4481 (N_4481,In_3657,In_893);
nand U4482 (N_4482,In_255,In_4468);
and U4483 (N_4483,In_1532,In_2221);
nand U4484 (N_4484,In_1290,In_3317);
xnor U4485 (N_4485,In_4678,In_1207);
nand U4486 (N_4486,In_741,In_4865);
nor U4487 (N_4487,In_2337,In_2691);
or U4488 (N_4488,In_4257,In_2495);
or U4489 (N_4489,In_2968,In_2406);
and U4490 (N_4490,In_344,In_4306);
xnor U4491 (N_4491,In_415,In_1063);
or U4492 (N_4492,In_1917,In_2730);
and U4493 (N_4493,In_1668,In_4899);
and U4494 (N_4494,In_1566,In_4574);
and U4495 (N_4495,In_4203,In_1746);
nand U4496 (N_4496,In_918,In_1878);
nor U4497 (N_4497,In_4771,In_1943);
xnor U4498 (N_4498,In_4150,In_3124);
or U4499 (N_4499,In_4782,In_372);
xnor U4500 (N_4500,In_2409,In_3985);
or U4501 (N_4501,In_3878,In_2822);
nor U4502 (N_4502,In_2291,In_1942);
or U4503 (N_4503,In_2012,In_3608);
nor U4504 (N_4504,In_414,In_789);
and U4505 (N_4505,In_4183,In_2887);
nor U4506 (N_4506,In_4106,In_902);
and U4507 (N_4507,In_1393,In_4559);
or U4508 (N_4508,In_4380,In_283);
xor U4509 (N_4509,In_1514,In_2696);
nand U4510 (N_4510,In_3705,In_2736);
nor U4511 (N_4511,In_4692,In_3820);
and U4512 (N_4512,In_819,In_2917);
or U4513 (N_4513,In_325,In_2973);
xnor U4514 (N_4514,In_4447,In_2139);
nor U4515 (N_4515,In_4801,In_3177);
xnor U4516 (N_4516,In_2502,In_2474);
or U4517 (N_4517,In_4155,In_3835);
and U4518 (N_4518,In_1310,In_3826);
or U4519 (N_4519,In_687,In_338);
xnor U4520 (N_4520,In_4708,In_1415);
xor U4521 (N_4521,In_1942,In_3397);
or U4522 (N_4522,In_2951,In_2267);
xnor U4523 (N_4523,In_4371,In_2191);
xnor U4524 (N_4524,In_702,In_4272);
nand U4525 (N_4525,In_937,In_4859);
xnor U4526 (N_4526,In_3767,In_3606);
nor U4527 (N_4527,In_2326,In_4767);
or U4528 (N_4528,In_3320,In_2776);
and U4529 (N_4529,In_102,In_682);
and U4530 (N_4530,In_4103,In_341);
xor U4531 (N_4531,In_341,In_3231);
xnor U4532 (N_4532,In_2034,In_2834);
xnor U4533 (N_4533,In_1822,In_3848);
or U4534 (N_4534,In_4497,In_1654);
xnor U4535 (N_4535,In_909,In_4863);
nor U4536 (N_4536,In_4378,In_2352);
xor U4537 (N_4537,In_1904,In_1853);
xnor U4538 (N_4538,In_4664,In_4133);
nand U4539 (N_4539,In_1650,In_3908);
nand U4540 (N_4540,In_4201,In_930);
nand U4541 (N_4541,In_3002,In_4443);
and U4542 (N_4542,In_1798,In_2086);
nand U4543 (N_4543,In_3859,In_2356);
nor U4544 (N_4544,In_2217,In_44);
xor U4545 (N_4545,In_2087,In_3306);
nor U4546 (N_4546,In_4887,In_292);
xor U4547 (N_4547,In_4987,In_1112);
or U4548 (N_4548,In_809,In_3185);
nand U4549 (N_4549,In_1283,In_2959);
or U4550 (N_4550,In_1129,In_3051);
xnor U4551 (N_4551,In_2146,In_2823);
nand U4552 (N_4552,In_1217,In_4370);
nor U4553 (N_4553,In_3791,In_2809);
nand U4554 (N_4554,In_971,In_2552);
or U4555 (N_4555,In_3447,In_144);
nor U4556 (N_4556,In_4496,In_2090);
nor U4557 (N_4557,In_4259,In_430);
or U4558 (N_4558,In_3434,In_2872);
xnor U4559 (N_4559,In_4092,In_2623);
xnor U4560 (N_4560,In_3341,In_2407);
nor U4561 (N_4561,In_4452,In_1406);
nor U4562 (N_4562,In_4594,In_3699);
or U4563 (N_4563,In_2447,In_911);
or U4564 (N_4564,In_1798,In_3173);
and U4565 (N_4565,In_4853,In_2813);
and U4566 (N_4566,In_1828,In_58);
and U4567 (N_4567,In_3446,In_4663);
xor U4568 (N_4568,In_4277,In_1298);
or U4569 (N_4569,In_2256,In_2277);
nor U4570 (N_4570,In_2605,In_2140);
nor U4571 (N_4571,In_4323,In_4394);
nor U4572 (N_4572,In_4724,In_1165);
and U4573 (N_4573,In_1344,In_4259);
and U4574 (N_4574,In_920,In_4519);
nor U4575 (N_4575,In_2299,In_4135);
or U4576 (N_4576,In_2064,In_2664);
xnor U4577 (N_4577,In_1130,In_2365);
nor U4578 (N_4578,In_3508,In_2084);
xor U4579 (N_4579,In_1212,In_994);
and U4580 (N_4580,In_849,In_2640);
nand U4581 (N_4581,In_307,In_245);
nand U4582 (N_4582,In_4074,In_2105);
nand U4583 (N_4583,In_1247,In_4556);
or U4584 (N_4584,In_4038,In_4935);
xor U4585 (N_4585,In_1007,In_672);
nand U4586 (N_4586,In_1963,In_4300);
xor U4587 (N_4587,In_2277,In_511);
nor U4588 (N_4588,In_4572,In_78);
xnor U4589 (N_4589,In_2810,In_4852);
nor U4590 (N_4590,In_428,In_3038);
nand U4591 (N_4591,In_152,In_1990);
and U4592 (N_4592,In_666,In_3582);
xnor U4593 (N_4593,In_2761,In_343);
nor U4594 (N_4594,In_1362,In_2911);
xnor U4595 (N_4595,In_1578,In_2822);
and U4596 (N_4596,In_1717,In_840);
or U4597 (N_4597,In_534,In_1773);
xnor U4598 (N_4598,In_1697,In_1619);
and U4599 (N_4599,In_1474,In_1378);
and U4600 (N_4600,In_548,In_1202);
and U4601 (N_4601,In_2967,In_2070);
or U4602 (N_4602,In_3100,In_888);
xor U4603 (N_4603,In_272,In_257);
and U4604 (N_4604,In_4521,In_3835);
nand U4605 (N_4605,In_281,In_4429);
nor U4606 (N_4606,In_1845,In_4791);
and U4607 (N_4607,In_523,In_3746);
xnor U4608 (N_4608,In_3822,In_4636);
xor U4609 (N_4609,In_339,In_2363);
and U4610 (N_4610,In_3367,In_3847);
nor U4611 (N_4611,In_278,In_684);
and U4612 (N_4612,In_1886,In_441);
or U4613 (N_4613,In_3522,In_21);
and U4614 (N_4614,In_1471,In_473);
and U4615 (N_4615,In_1502,In_4015);
nor U4616 (N_4616,In_1958,In_4306);
or U4617 (N_4617,In_4441,In_2882);
xor U4618 (N_4618,In_1129,In_3822);
and U4619 (N_4619,In_3521,In_3538);
nand U4620 (N_4620,In_4820,In_1529);
xnor U4621 (N_4621,In_171,In_4587);
nor U4622 (N_4622,In_2382,In_769);
and U4623 (N_4623,In_256,In_3824);
or U4624 (N_4624,In_2516,In_2781);
and U4625 (N_4625,In_4301,In_1437);
or U4626 (N_4626,In_4106,In_1677);
xnor U4627 (N_4627,In_4719,In_1944);
xnor U4628 (N_4628,In_2260,In_2566);
nor U4629 (N_4629,In_2213,In_1065);
nand U4630 (N_4630,In_1411,In_3544);
and U4631 (N_4631,In_1044,In_3220);
xnor U4632 (N_4632,In_3378,In_3117);
and U4633 (N_4633,In_4029,In_4561);
and U4634 (N_4634,In_2256,In_4524);
nor U4635 (N_4635,In_281,In_2562);
nand U4636 (N_4636,In_1262,In_3587);
and U4637 (N_4637,In_375,In_277);
nand U4638 (N_4638,In_3624,In_2779);
nand U4639 (N_4639,In_817,In_2680);
and U4640 (N_4640,In_3670,In_3924);
nor U4641 (N_4641,In_2306,In_4884);
nor U4642 (N_4642,In_4451,In_186);
and U4643 (N_4643,In_2117,In_3501);
nand U4644 (N_4644,In_2574,In_3434);
nand U4645 (N_4645,In_2262,In_4799);
or U4646 (N_4646,In_1748,In_1028);
and U4647 (N_4647,In_3422,In_2839);
and U4648 (N_4648,In_672,In_1474);
nand U4649 (N_4649,In_3267,In_3707);
nor U4650 (N_4650,In_3290,In_3950);
xnor U4651 (N_4651,In_1545,In_3161);
or U4652 (N_4652,In_971,In_1191);
or U4653 (N_4653,In_2534,In_2901);
nand U4654 (N_4654,In_2887,In_4635);
xnor U4655 (N_4655,In_875,In_2870);
nand U4656 (N_4656,In_3501,In_4137);
nand U4657 (N_4657,In_537,In_1923);
or U4658 (N_4658,In_1321,In_1263);
xor U4659 (N_4659,In_113,In_3452);
nor U4660 (N_4660,In_355,In_3657);
xnor U4661 (N_4661,In_3439,In_666);
and U4662 (N_4662,In_825,In_294);
nand U4663 (N_4663,In_651,In_4179);
and U4664 (N_4664,In_2726,In_4216);
or U4665 (N_4665,In_1320,In_1877);
and U4666 (N_4666,In_1650,In_3772);
nand U4667 (N_4667,In_1181,In_746);
or U4668 (N_4668,In_676,In_4116);
and U4669 (N_4669,In_4659,In_4026);
nor U4670 (N_4670,In_732,In_217);
nand U4671 (N_4671,In_4627,In_2430);
or U4672 (N_4672,In_1594,In_2675);
nor U4673 (N_4673,In_2208,In_1797);
nor U4674 (N_4674,In_3877,In_3091);
xnor U4675 (N_4675,In_3598,In_1306);
nand U4676 (N_4676,In_2365,In_2056);
or U4677 (N_4677,In_4314,In_3138);
and U4678 (N_4678,In_1594,In_1198);
nand U4679 (N_4679,In_3218,In_2174);
and U4680 (N_4680,In_1046,In_4788);
and U4681 (N_4681,In_4994,In_3578);
or U4682 (N_4682,In_3397,In_3615);
xnor U4683 (N_4683,In_4490,In_3991);
or U4684 (N_4684,In_2698,In_2061);
nand U4685 (N_4685,In_4993,In_2974);
xor U4686 (N_4686,In_3539,In_2259);
or U4687 (N_4687,In_1698,In_2363);
nand U4688 (N_4688,In_3377,In_3541);
and U4689 (N_4689,In_274,In_1276);
nand U4690 (N_4690,In_1635,In_4373);
and U4691 (N_4691,In_3939,In_123);
nand U4692 (N_4692,In_3917,In_2900);
and U4693 (N_4693,In_3290,In_2015);
xnor U4694 (N_4694,In_4146,In_3262);
nand U4695 (N_4695,In_634,In_2231);
nor U4696 (N_4696,In_2965,In_3014);
nor U4697 (N_4697,In_1101,In_34);
xor U4698 (N_4698,In_104,In_3467);
nand U4699 (N_4699,In_1386,In_2369);
and U4700 (N_4700,In_4836,In_2774);
nor U4701 (N_4701,In_3778,In_2649);
nor U4702 (N_4702,In_3127,In_4329);
nor U4703 (N_4703,In_4898,In_1797);
or U4704 (N_4704,In_4780,In_3656);
or U4705 (N_4705,In_3377,In_543);
nand U4706 (N_4706,In_1639,In_1955);
and U4707 (N_4707,In_24,In_4204);
or U4708 (N_4708,In_4481,In_4557);
and U4709 (N_4709,In_3640,In_2573);
xnor U4710 (N_4710,In_3200,In_49);
nand U4711 (N_4711,In_3265,In_3967);
nor U4712 (N_4712,In_2701,In_3858);
nor U4713 (N_4713,In_132,In_3543);
xnor U4714 (N_4714,In_152,In_3030);
and U4715 (N_4715,In_4792,In_3051);
xnor U4716 (N_4716,In_485,In_4901);
or U4717 (N_4717,In_3029,In_87);
nand U4718 (N_4718,In_14,In_2389);
nor U4719 (N_4719,In_4013,In_4028);
xnor U4720 (N_4720,In_4756,In_641);
and U4721 (N_4721,In_4496,In_3224);
nor U4722 (N_4722,In_1979,In_2897);
and U4723 (N_4723,In_4935,In_54);
nor U4724 (N_4724,In_603,In_4972);
xnor U4725 (N_4725,In_736,In_293);
nand U4726 (N_4726,In_3026,In_4024);
nand U4727 (N_4727,In_4390,In_1358);
xnor U4728 (N_4728,In_4544,In_2535);
or U4729 (N_4729,In_1063,In_2532);
nor U4730 (N_4730,In_1851,In_3025);
or U4731 (N_4731,In_4461,In_2510);
and U4732 (N_4732,In_234,In_217);
xor U4733 (N_4733,In_1152,In_1616);
xor U4734 (N_4734,In_4699,In_2912);
or U4735 (N_4735,In_4948,In_3015);
nor U4736 (N_4736,In_1129,In_3407);
nor U4737 (N_4737,In_4939,In_4832);
nor U4738 (N_4738,In_22,In_3433);
nor U4739 (N_4739,In_19,In_4153);
or U4740 (N_4740,In_1096,In_106);
xor U4741 (N_4741,In_2377,In_3918);
and U4742 (N_4742,In_1834,In_165);
nor U4743 (N_4743,In_1120,In_184);
xnor U4744 (N_4744,In_3468,In_612);
and U4745 (N_4745,In_1330,In_3367);
nand U4746 (N_4746,In_2995,In_1524);
and U4747 (N_4747,In_3328,In_640);
or U4748 (N_4748,In_4119,In_620);
nor U4749 (N_4749,In_4126,In_4012);
xnor U4750 (N_4750,In_4848,In_562);
xnor U4751 (N_4751,In_2379,In_4983);
nor U4752 (N_4752,In_3808,In_2678);
nand U4753 (N_4753,In_3085,In_66);
nand U4754 (N_4754,In_1437,In_2858);
xnor U4755 (N_4755,In_1100,In_4329);
xor U4756 (N_4756,In_43,In_3317);
or U4757 (N_4757,In_4076,In_1962);
and U4758 (N_4758,In_448,In_1525);
xnor U4759 (N_4759,In_4842,In_4771);
and U4760 (N_4760,In_471,In_3018);
and U4761 (N_4761,In_2335,In_2446);
or U4762 (N_4762,In_386,In_2394);
or U4763 (N_4763,In_814,In_2911);
or U4764 (N_4764,In_4327,In_3007);
xor U4765 (N_4765,In_4795,In_4964);
or U4766 (N_4766,In_3691,In_1047);
xnor U4767 (N_4767,In_3367,In_2916);
or U4768 (N_4768,In_2478,In_4324);
xor U4769 (N_4769,In_478,In_459);
nand U4770 (N_4770,In_45,In_745);
or U4771 (N_4771,In_1233,In_2684);
xor U4772 (N_4772,In_4094,In_4531);
or U4773 (N_4773,In_3141,In_847);
nor U4774 (N_4774,In_3087,In_4961);
nor U4775 (N_4775,In_4137,In_4651);
and U4776 (N_4776,In_1045,In_3934);
or U4777 (N_4777,In_1908,In_4670);
nor U4778 (N_4778,In_2203,In_4889);
or U4779 (N_4779,In_1457,In_1624);
xnor U4780 (N_4780,In_3072,In_1263);
nor U4781 (N_4781,In_3226,In_1287);
nand U4782 (N_4782,In_2922,In_3993);
or U4783 (N_4783,In_2415,In_2362);
and U4784 (N_4784,In_1741,In_4163);
or U4785 (N_4785,In_4263,In_3767);
or U4786 (N_4786,In_2949,In_1320);
and U4787 (N_4787,In_2070,In_2);
nor U4788 (N_4788,In_2945,In_2316);
and U4789 (N_4789,In_418,In_1938);
xnor U4790 (N_4790,In_4817,In_1306);
xnor U4791 (N_4791,In_4705,In_205);
nand U4792 (N_4792,In_1026,In_1982);
nand U4793 (N_4793,In_4726,In_3433);
nor U4794 (N_4794,In_4389,In_739);
and U4795 (N_4795,In_1707,In_4674);
and U4796 (N_4796,In_3827,In_4513);
or U4797 (N_4797,In_524,In_1941);
xnor U4798 (N_4798,In_1447,In_4730);
and U4799 (N_4799,In_2707,In_1588);
and U4800 (N_4800,In_1282,In_2963);
and U4801 (N_4801,In_1384,In_663);
xnor U4802 (N_4802,In_3847,In_3772);
or U4803 (N_4803,In_2441,In_2918);
nor U4804 (N_4804,In_4213,In_2520);
and U4805 (N_4805,In_4611,In_4366);
xor U4806 (N_4806,In_2071,In_4891);
nand U4807 (N_4807,In_2710,In_1317);
and U4808 (N_4808,In_808,In_2991);
or U4809 (N_4809,In_3694,In_2173);
nor U4810 (N_4810,In_2512,In_3026);
nand U4811 (N_4811,In_4461,In_1143);
and U4812 (N_4812,In_604,In_32);
and U4813 (N_4813,In_68,In_3359);
nor U4814 (N_4814,In_2310,In_2363);
nand U4815 (N_4815,In_4430,In_3176);
and U4816 (N_4816,In_4364,In_3106);
xor U4817 (N_4817,In_1979,In_2692);
and U4818 (N_4818,In_3003,In_2897);
nor U4819 (N_4819,In_837,In_1752);
nand U4820 (N_4820,In_2673,In_291);
xnor U4821 (N_4821,In_3427,In_2847);
nor U4822 (N_4822,In_3976,In_3917);
nor U4823 (N_4823,In_1400,In_3671);
and U4824 (N_4824,In_2263,In_807);
nand U4825 (N_4825,In_4248,In_525);
nor U4826 (N_4826,In_3087,In_1940);
nand U4827 (N_4827,In_4239,In_4038);
or U4828 (N_4828,In_2057,In_2027);
nand U4829 (N_4829,In_2294,In_3506);
nand U4830 (N_4830,In_1373,In_1608);
and U4831 (N_4831,In_930,In_3826);
nand U4832 (N_4832,In_4642,In_3007);
nand U4833 (N_4833,In_4662,In_4764);
nor U4834 (N_4834,In_4212,In_4762);
and U4835 (N_4835,In_1401,In_1989);
nor U4836 (N_4836,In_3364,In_4095);
and U4837 (N_4837,In_576,In_2279);
nand U4838 (N_4838,In_448,In_135);
nand U4839 (N_4839,In_551,In_2634);
xnor U4840 (N_4840,In_4301,In_1968);
xor U4841 (N_4841,In_1366,In_3908);
and U4842 (N_4842,In_3586,In_2349);
nand U4843 (N_4843,In_4351,In_154);
or U4844 (N_4844,In_601,In_3915);
xor U4845 (N_4845,In_3459,In_2375);
or U4846 (N_4846,In_1434,In_3799);
nor U4847 (N_4847,In_2897,In_3893);
xnor U4848 (N_4848,In_3780,In_1232);
and U4849 (N_4849,In_4504,In_3047);
xor U4850 (N_4850,In_2934,In_4749);
nor U4851 (N_4851,In_4063,In_3846);
or U4852 (N_4852,In_4288,In_1471);
xnor U4853 (N_4853,In_3830,In_1233);
and U4854 (N_4854,In_2040,In_4606);
or U4855 (N_4855,In_1032,In_2149);
nor U4856 (N_4856,In_3880,In_2809);
and U4857 (N_4857,In_4047,In_4958);
and U4858 (N_4858,In_4305,In_4845);
or U4859 (N_4859,In_3908,In_1034);
xnor U4860 (N_4860,In_1285,In_954);
nor U4861 (N_4861,In_676,In_2582);
nand U4862 (N_4862,In_1162,In_4051);
nor U4863 (N_4863,In_4609,In_1211);
xor U4864 (N_4864,In_1946,In_1178);
or U4865 (N_4865,In_169,In_2606);
nand U4866 (N_4866,In_1578,In_2006);
nor U4867 (N_4867,In_657,In_864);
or U4868 (N_4868,In_2745,In_299);
xnor U4869 (N_4869,In_2046,In_3531);
and U4870 (N_4870,In_479,In_784);
and U4871 (N_4871,In_3074,In_762);
xnor U4872 (N_4872,In_2919,In_1768);
and U4873 (N_4873,In_1234,In_4795);
and U4874 (N_4874,In_4837,In_4596);
or U4875 (N_4875,In_2531,In_2327);
nand U4876 (N_4876,In_4696,In_2525);
or U4877 (N_4877,In_1790,In_4792);
nand U4878 (N_4878,In_1420,In_4691);
xnor U4879 (N_4879,In_3764,In_9);
or U4880 (N_4880,In_187,In_3855);
nand U4881 (N_4881,In_2241,In_4048);
and U4882 (N_4882,In_3815,In_57);
nor U4883 (N_4883,In_4856,In_295);
nor U4884 (N_4884,In_806,In_4740);
and U4885 (N_4885,In_1854,In_4431);
nor U4886 (N_4886,In_4399,In_122);
nand U4887 (N_4887,In_4809,In_4056);
or U4888 (N_4888,In_1010,In_383);
nand U4889 (N_4889,In_2192,In_2803);
xor U4890 (N_4890,In_3005,In_2093);
or U4891 (N_4891,In_1026,In_2692);
xnor U4892 (N_4892,In_1845,In_2792);
nor U4893 (N_4893,In_2642,In_1850);
nor U4894 (N_4894,In_2303,In_2654);
and U4895 (N_4895,In_2208,In_92);
nor U4896 (N_4896,In_2567,In_3656);
nor U4897 (N_4897,In_523,In_2625);
nor U4898 (N_4898,In_3503,In_2691);
or U4899 (N_4899,In_14,In_3482);
xnor U4900 (N_4900,In_1538,In_654);
and U4901 (N_4901,In_656,In_1396);
and U4902 (N_4902,In_1173,In_3819);
or U4903 (N_4903,In_872,In_4031);
or U4904 (N_4904,In_3369,In_2832);
and U4905 (N_4905,In_2909,In_207);
xnor U4906 (N_4906,In_1391,In_2307);
and U4907 (N_4907,In_1526,In_874);
nor U4908 (N_4908,In_2514,In_3552);
xor U4909 (N_4909,In_657,In_252);
nor U4910 (N_4910,In_2683,In_4235);
nor U4911 (N_4911,In_4015,In_1372);
xor U4912 (N_4912,In_4691,In_91);
nand U4913 (N_4913,In_1045,In_3639);
nand U4914 (N_4914,In_967,In_2728);
and U4915 (N_4915,In_2444,In_2229);
or U4916 (N_4916,In_4965,In_3847);
and U4917 (N_4917,In_188,In_496);
nor U4918 (N_4918,In_4325,In_110);
or U4919 (N_4919,In_2072,In_1480);
xor U4920 (N_4920,In_4983,In_971);
or U4921 (N_4921,In_4037,In_180);
xor U4922 (N_4922,In_1938,In_3314);
nand U4923 (N_4923,In_4417,In_1036);
and U4924 (N_4924,In_2665,In_1189);
nor U4925 (N_4925,In_2636,In_2612);
xor U4926 (N_4926,In_1242,In_3833);
xnor U4927 (N_4927,In_4487,In_1541);
and U4928 (N_4928,In_1191,In_4894);
nor U4929 (N_4929,In_2202,In_2545);
xor U4930 (N_4930,In_771,In_4212);
and U4931 (N_4931,In_3128,In_1852);
xor U4932 (N_4932,In_731,In_649);
and U4933 (N_4933,In_2165,In_4783);
and U4934 (N_4934,In_1224,In_604);
nand U4935 (N_4935,In_3325,In_3519);
xor U4936 (N_4936,In_4748,In_822);
xor U4937 (N_4937,In_3162,In_2992);
or U4938 (N_4938,In_912,In_1528);
nand U4939 (N_4939,In_2729,In_589);
xnor U4940 (N_4940,In_1971,In_3304);
nand U4941 (N_4941,In_1447,In_236);
nor U4942 (N_4942,In_766,In_297);
nand U4943 (N_4943,In_3559,In_949);
xor U4944 (N_4944,In_1826,In_2125);
nand U4945 (N_4945,In_159,In_185);
nand U4946 (N_4946,In_2333,In_2784);
nor U4947 (N_4947,In_727,In_3043);
and U4948 (N_4948,In_3160,In_4611);
xor U4949 (N_4949,In_4229,In_3085);
and U4950 (N_4950,In_3884,In_1547);
or U4951 (N_4951,In_547,In_4741);
nand U4952 (N_4952,In_3254,In_1923);
xor U4953 (N_4953,In_2765,In_510);
xnor U4954 (N_4954,In_1086,In_2721);
and U4955 (N_4955,In_4694,In_2295);
and U4956 (N_4956,In_2918,In_3983);
and U4957 (N_4957,In_4057,In_684);
nand U4958 (N_4958,In_2604,In_3000);
or U4959 (N_4959,In_3084,In_352);
nand U4960 (N_4960,In_1117,In_4032);
nor U4961 (N_4961,In_1265,In_2686);
xor U4962 (N_4962,In_1695,In_3233);
nor U4963 (N_4963,In_2367,In_3621);
nor U4964 (N_4964,In_1419,In_4722);
nand U4965 (N_4965,In_182,In_1200);
and U4966 (N_4966,In_4981,In_2069);
nor U4967 (N_4967,In_397,In_3024);
xor U4968 (N_4968,In_2502,In_4547);
xor U4969 (N_4969,In_1088,In_4825);
or U4970 (N_4970,In_1767,In_3329);
xnor U4971 (N_4971,In_4993,In_48);
xor U4972 (N_4972,In_1986,In_4440);
and U4973 (N_4973,In_558,In_4608);
nor U4974 (N_4974,In_1941,In_2424);
xnor U4975 (N_4975,In_3941,In_1436);
nor U4976 (N_4976,In_3655,In_4844);
or U4977 (N_4977,In_4158,In_1095);
xor U4978 (N_4978,In_3315,In_1352);
or U4979 (N_4979,In_2775,In_4850);
nand U4980 (N_4980,In_4459,In_217);
nand U4981 (N_4981,In_3975,In_35);
xor U4982 (N_4982,In_909,In_829);
or U4983 (N_4983,In_624,In_264);
nor U4984 (N_4984,In_2931,In_1872);
or U4985 (N_4985,In_4812,In_476);
xor U4986 (N_4986,In_121,In_1783);
and U4987 (N_4987,In_1694,In_4078);
or U4988 (N_4988,In_2109,In_4968);
nor U4989 (N_4989,In_4086,In_2941);
nand U4990 (N_4990,In_4886,In_4129);
or U4991 (N_4991,In_4162,In_3647);
xnor U4992 (N_4992,In_2911,In_1748);
nand U4993 (N_4993,In_1186,In_1445);
nand U4994 (N_4994,In_1477,In_4474);
and U4995 (N_4995,In_2584,In_1658);
nor U4996 (N_4996,In_2865,In_1437);
and U4997 (N_4997,In_4295,In_2647);
nand U4998 (N_4998,In_1343,In_2458);
or U4999 (N_4999,In_910,In_2587);
xor U5000 (N_5000,N_1597,N_1433);
nor U5001 (N_5001,N_4058,N_379);
or U5002 (N_5002,N_1425,N_1338);
and U5003 (N_5003,N_1127,N_4380);
xnor U5004 (N_5004,N_1337,N_15);
xnor U5005 (N_5005,N_4055,N_905);
nor U5006 (N_5006,N_688,N_526);
and U5007 (N_5007,N_3709,N_2007);
and U5008 (N_5008,N_4390,N_88);
or U5009 (N_5009,N_4864,N_2789);
or U5010 (N_5010,N_1431,N_533);
or U5011 (N_5011,N_2676,N_3561);
and U5012 (N_5012,N_1032,N_4674);
or U5013 (N_5013,N_2513,N_1120);
or U5014 (N_5014,N_2812,N_833);
and U5015 (N_5015,N_876,N_4612);
and U5016 (N_5016,N_1605,N_2759);
nor U5017 (N_5017,N_3345,N_3245);
nor U5018 (N_5018,N_2981,N_2714);
xor U5019 (N_5019,N_476,N_4936);
and U5020 (N_5020,N_3381,N_1514);
and U5021 (N_5021,N_2288,N_1799);
nand U5022 (N_5022,N_2182,N_1414);
and U5023 (N_5023,N_2046,N_3021);
nand U5024 (N_5024,N_4983,N_2600);
xnor U5025 (N_5025,N_1716,N_3139);
nand U5026 (N_5026,N_1174,N_1457);
xor U5027 (N_5027,N_1576,N_696);
and U5028 (N_5028,N_4425,N_2788);
nand U5029 (N_5029,N_317,N_1460);
or U5030 (N_5030,N_1383,N_2341);
nor U5031 (N_5031,N_3630,N_2756);
xor U5032 (N_5032,N_377,N_3931);
xnor U5033 (N_5033,N_4335,N_626);
or U5034 (N_5034,N_76,N_4582);
nand U5035 (N_5035,N_669,N_316);
xnor U5036 (N_5036,N_1114,N_291);
xnor U5037 (N_5037,N_2819,N_2033);
nand U5038 (N_5038,N_2234,N_1620);
xnor U5039 (N_5039,N_3171,N_2066);
and U5040 (N_5040,N_2663,N_1082);
nor U5041 (N_5041,N_3358,N_2317);
xor U5042 (N_5042,N_881,N_415);
and U5043 (N_5043,N_1276,N_3273);
nor U5044 (N_5044,N_513,N_4362);
or U5045 (N_5045,N_3162,N_2994);
xnor U5046 (N_5046,N_2790,N_4053);
and U5047 (N_5047,N_1573,N_734);
and U5048 (N_5048,N_269,N_1051);
nand U5049 (N_5049,N_1874,N_497);
and U5050 (N_5050,N_4742,N_3946);
nand U5051 (N_5051,N_3847,N_4236);
or U5052 (N_5052,N_2154,N_4049);
nand U5053 (N_5053,N_3629,N_198);
and U5054 (N_5054,N_3572,N_2474);
and U5055 (N_5055,N_2476,N_3953);
and U5056 (N_5056,N_3750,N_3934);
nand U5057 (N_5057,N_1148,N_1316);
nor U5058 (N_5058,N_3564,N_1462);
nor U5059 (N_5059,N_3527,N_1057);
nand U5060 (N_5060,N_667,N_3004);
or U5061 (N_5061,N_4997,N_3743);
and U5062 (N_5062,N_3454,N_3996);
xor U5063 (N_5063,N_1357,N_1151);
xor U5064 (N_5064,N_3870,N_3951);
nor U5065 (N_5065,N_2316,N_4976);
xor U5066 (N_5066,N_4022,N_346);
nor U5067 (N_5067,N_2704,N_580);
nor U5068 (N_5068,N_1701,N_795);
xnor U5069 (N_5069,N_3145,N_1843);
and U5070 (N_5070,N_2520,N_93);
nand U5071 (N_5071,N_4109,N_3055);
xor U5072 (N_5072,N_2367,N_416);
xnor U5073 (N_5073,N_1271,N_1275);
xor U5074 (N_5074,N_81,N_808);
nor U5075 (N_5075,N_351,N_869);
nand U5076 (N_5076,N_2694,N_3195);
xor U5077 (N_5077,N_1633,N_2861);
xor U5078 (N_5078,N_1778,N_1961);
nand U5079 (N_5079,N_1652,N_678);
or U5080 (N_5080,N_2293,N_237);
xor U5081 (N_5081,N_4561,N_2507);
and U5082 (N_5082,N_2090,N_3801);
nand U5083 (N_5083,N_756,N_1606);
and U5084 (N_5084,N_4373,N_1073);
nand U5085 (N_5085,N_1291,N_559);
xnor U5086 (N_5086,N_370,N_1865);
nand U5087 (N_5087,N_4801,N_4006);
nand U5088 (N_5088,N_1679,N_4166);
and U5089 (N_5089,N_3637,N_214);
xor U5090 (N_5090,N_3278,N_3863);
nor U5091 (N_5091,N_331,N_2486);
and U5092 (N_5092,N_1964,N_4147);
nand U5093 (N_5093,N_1709,N_4164);
xnor U5094 (N_5094,N_3746,N_3272);
and U5095 (N_5095,N_1647,N_3445);
nand U5096 (N_5096,N_713,N_2282);
nand U5097 (N_5097,N_4887,N_298);
nor U5098 (N_5098,N_1988,N_1039);
xor U5099 (N_5099,N_1705,N_1583);
or U5100 (N_5100,N_1690,N_501);
xor U5101 (N_5101,N_483,N_3940);
nand U5102 (N_5102,N_4921,N_2947);
and U5103 (N_5103,N_4880,N_1826);
or U5104 (N_5104,N_822,N_3897);
xnor U5105 (N_5105,N_343,N_4126);
xor U5106 (N_5106,N_1128,N_3574);
and U5107 (N_5107,N_4306,N_1370);
and U5108 (N_5108,N_850,N_1984);
or U5109 (N_5109,N_4341,N_4506);
or U5110 (N_5110,N_1839,N_1250);
and U5111 (N_5111,N_2473,N_2678);
xnor U5112 (N_5112,N_4751,N_2987);
nor U5113 (N_5113,N_4077,N_3713);
xnor U5114 (N_5114,N_4688,N_1044);
nor U5115 (N_5115,N_1960,N_141);
xnor U5116 (N_5116,N_2924,N_2436);
or U5117 (N_5117,N_4500,N_4331);
nor U5118 (N_5118,N_1777,N_1156);
xnor U5119 (N_5119,N_4776,N_4803);
xor U5120 (N_5120,N_3677,N_2722);
xnor U5121 (N_5121,N_1225,N_2761);
nor U5122 (N_5122,N_2682,N_1036);
xnor U5123 (N_5123,N_2362,N_2307);
xnor U5124 (N_5124,N_3204,N_962);
xor U5125 (N_5125,N_3829,N_3288);
nand U5126 (N_5126,N_666,N_920);
and U5127 (N_5127,N_3938,N_3699);
or U5128 (N_5128,N_427,N_4549);
xnor U5129 (N_5129,N_2503,N_2271);
nor U5130 (N_5130,N_1065,N_985);
and U5131 (N_5131,N_2427,N_4656);
nand U5132 (N_5132,N_524,N_4903);
xor U5133 (N_5133,N_1177,N_1422);
xor U5134 (N_5134,N_1327,N_1890);
xor U5135 (N_5135,N_1458,N_4619);
nor U5136 (N_5136,N_692,N_2934);
or U5137 (N_5137,N_2057,N_2747);
xor U5138 (N_5138,N_4105,N_4133);
and U5139 (N_5139,N_3987,N_395);
and U5140 (N_5140,N_4945,N_310);
xor U5141 (N_5141,N_2811,N_1043);
xnor U5142 (N_5142,N_1509,N_138);
nor U5143 (N_5143,N_1665,N_208);
nor U5144 (N_5144,N_322,N_4322);
nor U5145 (N_5145,N_2283,N_2719);
nor U5146 (N_5146,N_4635,N_1328);
or U5147 (N_5147,N_870,N_3261);
xor U5148 (N_5148,N_2866,N_1171);
xor U5149 (N_5149,N_1915,N_4677);
and U5150 (N_5150,N_791,N_4289);
xnor U5151 (N_5151,N_3624,N_1943);
nor U5152 (N_5152,N_968,N_3899);
or U5153 (N_5153,N_4944,N_1612);
and U5154 (N_5154,N_1083,N_3366);
and U5155 (N_5155,N_1313,N_352);
or U5156 (N_5156,N_3134,N_4777);
nor U5157 (N_5157,N_4923,N_2772);
nor U5158 (N_5158,N_2312,N_4404);
xor U5159 (N_5159,N_970,N_407);
and U5160 (N_5160,N_54,N_3112);
nand U5161 (N_5161,N_3168,N_1902);
and U5162 (N_5162,N_193,N_2343);
xnor U5163 (N_5163,N_3242,N_4451);
xnor U5164 (N_5164,N_4138,N_1766);
nor U5165 (N_5165,N_3076,N_1437);
nor U5166 (N_5166,N_4483,N_1215);
xnor U5167 (N_5167,N_4630,N_4408);
nand U5168 (N_5168,N_3547,N_861);
xnor U5169 (N_5169,N_1207,N_838);
xor U5170 (N_5170,N_2272,N_374);
nor U5171 (N_5171,N_4488,N_3207);
xor U5172 (N_5172,N_897,N_503);
nand U5173 (N_5173,N_179,N_5);
nor U5174 (N_5174,N_934,N_4280);
and U5175 (N_5175,N_3529,N_4461);
xor U5176 (N_5176,N_649,N_1314);
xnor U5177 (N_5177,N_3775,N_1190);
and U5178 (N_5178,N_2675,N_2541);
and U5179 (N_5179,N_3176,N_3668);
nor U5180 (N_5180,N_3828,N_1521);
or U5181 (N_5181,N_4465,N_3675);
nor U5182 (N_5182,N_92,N_973);
and U5183 (N_5183,N_2415,N_2303);
nand U5184 (N_5184,N_2468,N_1382);
or U5185 (N_5185,N_3429,N_2273);
or U5186 (N_5186,N_4340,N_2519);
nand U5187 (N_5187,N_4848,N_4297);
nand U5188 (N_5188,N_187,N_4653);
and U5189 (N_5189,N_4965,N_2211);
or U5190 (N_5190,N_4876,N_3117);
nor U5191 (N_5191,N_247,N_4015);
nor U5192 (N_5192,N_3126,N_3715);
nor U5193 (N_5193,N_4261,N_3289);
xor U5194 (N_5194,N_2992,N_4134);
xnor U5195 (N_5195,N_4860,N_4243);
nand U5196 (N_5196,N_2280,N_1516);
and U5197 (N_5197,N_3632,N_2696);
nor U5198 (N_5198,N_770,N_3688);
nor U5199 (N_5199,N_1661,N_1793);
xnor U5200 (N_5200,N_4118,N_587);
xor U5201 (N_5201,N_1103,N_2948);
or U5202 (N_5202,N_2375,N_3905);
and U5203 (N_5203,N_455,N_4646);
nand U5204 (N_5204,N_1080,N_3158);
nor U5205 (N_5205,N_4173,N_1903);
or U5206 (N_5206,N_4512,N_708);
nand U5207 (N_5207,N_2188,N_1687);
nor U5208 (N_5208,N_4478,N_184);
xor U5209 (N_5209,N_2103,N_4087);
and U5210 (N_5210,N_4569,N_772);
and U5211 (N_5211,N_3724,N_1582);
or U5212 (N_5212,N_3900,N_436);
and U5213 (N_5213,N_2708,N_2326);
xor U5214 (N_5214,N_1400,N_385);
xnor U5215 (N_5215,N_4857,N_2522);
nor U5216 (N_5216,N_376,N_639);
xor U5217 (N_5217,N_1362,N_3385);
nand U5218 (N_5218,N_4604,N_3469);
or U5219 (N_5219,N_223,N_3177);
and U5220 (N_5220,N_202,N_2430);
and U5221 (N_5221,N_623,N_2502);
and U5222 (N_5222,N_3943,N_1512);
nor U5223 (N_5223,N_4479,N_1332);
nor U5224 (N_5224,N_279,N_2142);
nand U5225 (N_5225,N_2127,N_605);
xor U5226 (N_5226,N_4691,N_4245);
and U5227 (N_5227,N_26,N_2816);
nor U5228 (N_5228,N_4484,N_2223);
nand U5229 (N_5229,N_3571,N_4188);
or U5230 (N_5230,N_3045,N_2567);
nor U5231 (N_5231,N_1050,N_3369);
nand U5232 (N_5232,N_439,N_472);
nand U5233 (N_5233,N_4196,N_381);
nand U5234 (N_5234,N_236,N_2310);
nor U5235 (N_5235,N_1408,N_3078);
and U5236 (N_5236,N_793,N_3077);
or U5237 (N_5237,N_3325,N_2699);
nor U5238 (N_5238,N_2885,N_456);
xor U5239 (N_5239,N_4456,N_1415);
and U5240 (N_5240,N_723,N_3769);
nor U5241 (N_5241,N_835,N_646);
or U5242 (N_5242,N_681,N_2156);
nand U5243 (N_5243,N_3956,N_4050);
or U5244 (N_5244,N_1532,N_787);
nor U5245 (N_5245,N_2721,N_2642);
xor U5246 (N_5246,N_459,N_4292);
xor U5247 (N_5247,N_3155,N_1305);
nor U5248 (N_5248,N_947,N_312);
and U5249 (N_5249,N_309,N_4787);
or U5250 (N_5250,N_160,N_717);
nand U5251 (N_5251,N_2017,N_327);
nand U5252 (N_5252,N_2203,N_4939);
nor U5253 (N_5253,N_2966,N_4692);
nor U5254 (N_5254,N_3172,N_520);
nand U5255 (N_5255,N_4625,N_1161);
nor U5256 (N_5256,N_546,N_2441);
nand U5257 (N_5257,N_4013,N_1166);
nor U5258 (N_5258,N_1323,N_1420);
xor U5259 (N_5259,N_2974,N_661);
nand U5260 (N_5260,N_4667,N_1997);
nand U5261 (N_5261,N_819,N_468);
or U5262 (N_5262,N_3714,N_1554);
nand U5263 (N_5263,N_2794,N_4120);
or U5264 (N_5264,N_1478,N_4185);
xor U5265 (N_5265,N_2710,N_1900);
nand U5266 (N_5266,N_2650,N_2231);
xor U5267 (N_5267,N_4930,N_2775);
nand U5268 (N_5268,N_1140,N_2944);
and U5269 (N_5269,N_2392,N_1577);
or U5270 (N_5270,N_1263,N_1767);
xor U5271 (N_5271,N_2477,N_2830);
nor U5272 (N_5272,N_529,N_4905);
nor U5273 (N_5273,N_1945,N_2796);
xnor U5274 (N_5274,N_1117,N_2049);
nor U5275 (N_5275,N_711,N_3950);
xor U5276 (N_5276,N_3584,N_767);
and U5277 (N_5277,N_3635,N_2443);
nor U5278 (N_5278,N_1550,N_4293);
nor U5279 (N_5279,N_3865,N_3662);
nand U5280 (N_5280,N_4665,N_1026);
nor U5281 (N_5281,N_817,N_2099);
and U5282 (N_5282,N_1423,N_1999);
nor U5283 (N_5283,N_2933,N_3917);
nor U5284 (N_5284,N_1124,N_752);
nor U5285 (N_5285,N_3933,N_2281);
xnor U5286 (N_5286,N_7,N_3696);
or U5287 (N_5287,N_4181,N_3562);
xnor U5288 (N_5288,N_1153,N_3263);
and U5289 (N_5289,N_679,N_3538);
nand U5290 (N_5290,N_1780,N_63);
nand U5291 (N_5291,N_3188,N_4559);
nand U5292 (N_5292,N_442,N_2378);
nand U5293 (N_5293,N_273,N_647);
xnor U5294 (N_5294,N_1214,N_4144);
nor U5295 (N_5295,N_4774,N_1027);
and U5296 (N_5296,N_3658,N_4570);
nor U5297 (N_5297,N_2777,N_4186);
nand U5298 (N_5298,N_3720,N_2357);
or U5299 (N_5299,N_1293,N_4629);
nor U5300 (N_5300,N_2973,N_1424);
and U5301 (N_5301,N_41,N_4176);
or U5302 (N_5302,N_3974,N_1385);
or U5303 (N_5303,N_2639,N_2290);
and U5304 (N_5304,N_815,N_2657);
nor U5305 (N_5305,N_1591,N_1378);
nand U5306 (N_5306,N_1607,N_3485);
and U5307 (N_5307,N_2077,N_2327);
nand U5308 (N_5308,N_4648,N_3410);
nand U5309 (N_5309,N_2423,N_1618);
nand U5310 (N_5310,N_2347,N_4542);
or U5311 (N_5311,N_2419,N_3898);
and U5312 (N_5312,N_1930,N_726);
nand U5313 (N_5313,N_531,N_414);
and U5314 (N_5314,N_3767,N_3545);
nand U5315 (N_5315,N_3178,N_2198);
xor U5316 (N_5316,N_4645,N_3267);
or U5317 (N_5317,N_4723,N_360);
xor U5318 (N_5318,N_4869,N_3615);
or U5319 (N_5319,N_949,N_2259);
nor U5320 (N_5320,N_2172,N_776);
nor U5321 (N_5321,N_3731,N_4640);
nor U5322 (N_5322,N_3038,N_3067);
nand U5323 (N_5323,N_3739,N_378);
nor U5324 (N_5324,N_3339,N_2649);
and U5325 (N_5325,N_3248,N_4127);
xnor U5326 (N_5326,N_1038,N_2093);
or U5327 (N_5327,N_4088,N_4035);
nor U5328 (N_5328,N_3444,N_4423);
xor U5329 (N_5329,N_1531,N_446);
nor U5330 (N_5330,N_78,N_3842);
nor U5331 (N_5331,N_2314,N_577);
nor U5332 (N_5332,N_3302,N_673);
xnor U5333 (N_5333,N_1565,N_2533);
xnor U5334 (N_5334,N_4272,N_3378);
or U5335 (N_5335,N_3411,N_4762);
and U5336 (N_5336,N_3463,N_926);
xnor U5337 (N_5337,N_267,N_4003);
or U5338 (N_5338,N_1643,N_3832);
and U5339 (N_5339,N_1926,N_3484);
nor U5340 (N_5340,N_242,N_4269);
nand U5341 (N_5341,N_797,N_4826);
and U5342 (N_5342,N_140,N_1838);
xnor U5343 (N_5343,N_480,N_4583);
nand U5344 (N_5344,N_1998,N_2771);
or U5345 (N_5345,N_473,N_2634);
nor U5346 (N_5346,N_1367,N_2038);
nand U5347 (N_5347,N_1243,N_2518);
xor U5348 (N_5348,N_2815,N_4329);
nand U5349 (N_5349,N_412,N_2523);
and U5350 (N_5350,N_335,N_4866);
and U5351 (N_5351,N_4299,N_499);
or U5352 (N_5352,N_1788,N_386);
and U5353 (N_5353,N_3773,N_2920);
nand U5354 (N_5354,N_4573,N_4242);
or U5355 (N_5355,N_2020,N_115);
xnor U5356 (N_5356,N_1523,N_4831);
nand U5357 (N_5357,N_4952,N_2487);
and U5358 (N_5358,N_1613,N_345);
and U5359 (N_5359,N_1954,N_4135);
nor U5360 (N_5360,N_2851,N_2558);
or U5361 (N_5361,N_1211,N_2905);
xnor U5362 (N_5362,N_1791,N_1594);
or U5363 (N_5363,N_125,N_2045);
or U5364 (N_5364,N_397,N_2778);
xor U5365 (N_5365,N_1432,N_4676);
and U5366 (N_5366,N_3137,N_4989);
xnor U5367 (N_5367,N_2892,N_816);
nand U5368 (N_5368,N_1419,N_4810);
or U5369 (N_5369,N_3671,N_1031);
nor U5370 (N_5370,N_4900,N_891);
or U5371 (N_5371,N_1005,N_929);
nor U5372 (N_5372,N_2009,N_2592);
nor U5373 (N_5373,N_3111,N_2619);
or U5374 (N_5374,N_528,N_883);
xor U5375 (N_5375,N_4195,N_2988);
nor U5376 (N_5376,N_1773,N_4727);
nor U5377 (N_5377,N_301,N_4699);
and U5378 (N_5378,N_548,N_1800);
or U5379 (N_5379,N_4453,N_4139);
and U5380 (N_5380,N_1201,N_2850);
or U5381 (N_5381,N_3262,N_3200);
or U5382 (N_5382,N_257,N_4455);
xnor U5383 (N_5383,N_3152,N_2764);
nand U5384 (N_5384,N_2661,N_3970);
nand U5385 (N_5385,N_2845,N_544);
xnor U5386 (N_5386,N_4644,N_4529);
nand U5387 (N_5387,N_3011,N_4252);
nand U5388 (N_5388,N_3355,N_2927);
nand U5389 (N_5389,N_2346,N_550);
xor U5390 (N_5390,N_4370,N_4572);
nand U5391 (N_5391,N_4378,N_24);
nand U5392 (N_5392,N_2806,N_182);
and U5393 (N_5393,N_1446,N_1950);
nand U5394 (N_5394,N_59,N_2638);
and U5395 (N_5395,N_3238,N_4333);
nand U5396 (N_5396,N_2849,N_443);
and U5397 (N_5397,N_2904,N_2583);
nand U5398 (N_5398,N_4314,N_2589);
xor U5399 (N_5399,N_1410,N_2113);
or U5400 (N_5400,N_1831,N_1680);
xor U5401 (N_5401,N_2003,N_42);
nand U5402 (N_5402,N_0,N_3947);
or U5403 (N_5403,N_1341,N_831);
xnor U5404 (N_5404,N_3108,N_1588);
and U5405 (N_5405,N_2148,N_1299);
or U5406 (N_5406,N_3336,N_2799);
and U5407 (N_5407,N_2041,N_742);
and U5408 (N_5408,N_3215,N_625);
and U5409 (N_5409,N_1427,N_4621);
nand U5410 (N_5410,N_4096,N_1671);
nor U5411 (N_5411,N_1557,N_3493);
and U5412 (N_5412,N_2718,N_11);
or U5413 (N_5413,N_4060,N_2121);
or U5414 (N_5414,N_2688,N_3462);
nor U5415 (N_5415,N_1237,N_1209);
xor U5416 (N_5416,N_2820,N_4654);
nor U5417 (N_5417,N_1563,N_2683);
nand U5418 (N_5418,N_2371,N_1682);
xor U5419 (N_5419,N_3570,N_2488);
nor U5420 (N_5420,N_3114,N_1741);
nor U5421 (N_5421,N_2725,N_959);
nand U5422 (N_5422,N_1899,N_3118);
nand U5423 (N_5423,N_2137,N_2043);
and U5424 (N_5424,N_3846,N_2313);
xor U5425 (N_5425,N_4175,N_864);
xnor U5426 (N_5426,N_4706,N_545);
xnor U5427 (N_5427,N_2630,N_3164);
nor U5428 (N_5428,N_2695,N_4489);
or U5429 (N_5429,N_2229,N_4525);
or U5430 (N_5430,N_83,N_2318);
nor U5431 (N_5431,N_1466,N_2438);
nor U5432 (N_5432,N_2416,N_2984);
and U5433 (N_5433,N_203,N_2654);
and U5434 (N_5434,N_2405,N_2475);
nand U5435 (N_5435,N_305,N_200);
nand U5436 (N_5436,N_2387,N_3972);
and U5437 (N_5437,N_4216,N_159);
xor U5438 (N_5438,N_2680,N_3450);
and U5439 (N_5439,N_4639,N_1648);
nor U5440 (N_5440,N_2945,N_3525);
nor U5441 (N_5441,N_3908,N_164);
nor U5442 (N_5442,N_3659,N_1480);
nand U5443 (N_5443,N_1830,N_930);
and U5444 (N_5444,N_4950,N_515);
nand U5445 (N_5445,N_3580,N_2542);
nand U5446 (N_5446,N_296,N_3845);
nor U5447 (N_5447,N_3534,N_84);
or U5448 (N_5448,N_4701,N_1738);
and U5449 (N_5449,N_3729,N_856);
nor U5450 (N_5450,N_4286,N_4785);
nand U5451 (N_5451,N_810,N_4247);
nor U5452 (N_5452,N_2836,N_1189);
nor U5453 (N_5453,N_199,N_496);
nand U5454 (N_5454,N_4334,N_1872);
xnor U5455 (N_5455,N_2410,N_38);
or U5456 (N_5456,N_3969,N_1146);
xor U5457 (N_5457,N_4112,N_1624);
nand U5458 (N_5458,N_4204,N_2394);
xor U5459 (N_5459,N_3376,N_746);
and U5460 (N_5460,N_1137,N_3867);
xnor U5461 (N_5461,N_4814,N_1416);
and U5462 (N_5462,N_1343,N_4564);
nand U5463 (N_5463,N_2525,N_2136);
or U5464 (N_5464,N_3896,N_2301);
nor U5465 (N_5465,N_1506,N_85);
or U5466 (N_5466,N_4255,N_3935);
nor U5467 (N_5467,N_3284,N_1494);
xor U5468 (N_5468,N_2183,N_3024);
and U5469 (N_5469,N_4931,N_2989);
nor U5470 (N_5470,N_2300,N_2228);
nor U5471 (N_5471,N_1438,N_100);
or U5472 (N_5472,N_1349,N_3387);
and U5473 (N_5473,N_4424,N_3069);
xnor U5474 (N_5474,N_4100,N_3957);
nor U5475 (N_5475,N_1905,N_201);
nor U5476 (N_5476,N_4224,N_3730);
and U5477 (N_5477,N_4560,N_3554);
and U5478 (N_5478,N_4412,N_4153);
xor U5479 (N_5479,N_3085,N_2717);
nor U5480 (N_5480,N_1819,N_1059);
nand U5481 (N_5481,N_4310,N_3857);
and U5482 (N_5482,N_1195,N_2377);
nor U5483 (N_5483,N_4940,N_4494);
nor U5484 (N_5484,N_4799,N_3920);
xor U5485 (N_5485,N_1798,N_354);
xnor U5486 (N_5486,N_3567,N_4778);
xnor U5487 (N_5487,N_2773,N_4843);
and U5488 (N_5488,N_675,N_1035);
xor U5489 (N_5489,N_2685,N_4704);
nand U5490 (N_5490,N_4915,N_1786);
xor U5491 (N_5491,N_4215,N_4993);
nand U5492 (N_5492,N_2795,N_1789);
and U5493 (N_5493,N_798,N_4697);
and U5494 (N_5494,N_1084,N_4470);
or U5495 (N_5495,N_3211,N_4889);
nor U5496 (N_5496,N_2365,N_1732);
nor U5497 (N_5497,N_809,N_3408);
and U5498 (N_5498,N_1335,N_3367);
or U5499 (N_5499,N_1750,N_3487);
nor U5500 (N_5500,N_4082,N_1277);
xor U5501 (N_5501,N_4853,N_3505);
nand U5502 (N_5502,N_619,N_4394);
xnor U5503 (N_5503,N_2833,N_4368);
nand U5504 (N_5504,N_1049,N_329);
nand U5505 (N_5505,N_2027,N_500);
nor U5506 (N_5506,N_1692,N_4338);
nor U5507 (N_5507,N_4177,N_1574);
and U5508 (N_5508,N_844,N_3531);
and U5509 (N_5509,N_3048,N_1398);
or U5510 (N_5510,N_774,N_1745);
nand U5511 (N_5511,N_4917,N_1540);
xor U5512 (N_5512,N_3783,N_4482);
and U5513 (N_5513,N_3359,N_4967);
nand U5514 (N_5514,N_2181,N_1465);
nor U5515 (N_5515,N_2946,N_1555);
nand U5516 (N_5516,N_347,N_348);
and U5517 (N_5517,N_474,N_3116);
or U5518 (N_5518,N_802,N_2372);
nand U5519 (N_5519,N_943,N_4347);
or U5520 (N_5520,N_956,N_289);
or U5521 (N_5521,N_4441,N_4822);
nor U5522 (N_5522,N_4039,N_2186);
nand U5523 (N_5523,N_1658,N_1992);
xor U5524 (N_5524,N_91,N_2434);
xor U5525 (N_5525,N_3517,N_4416);
or U5526 (N_5526,N_2995,N_2728);
xor U5527 (N_5527,N_1763,N_1795);
or U5528 (N_5528,N_2595,N_2413);
xor U5529 (N_5529,N_4251,N_3756);
xor U5530 (N_5530,N_4136,N_3252);
or U5531 (N_5531,N_3184,N_2063);
nor U5532 (N_5532,N_336,N_3109);
nor U5533 (N_5533,N_4984,N_4471);
or U5534 (N_5534,N_2258,N_3961);
nand U5535 (N_5535,N_3704,N_2428);
and U5536 (N_5536,N_3903,N_1740);
nor U5537 (N_5537,N_4641,N_1487);
or U5538 (N_5538,N_2490,N_1562);
and U5539 (N_5539,N_4693,N_4695);
nand U5540 (N_5540,N_607,N_2384);
nor U5541 (N_5541,N_3174,N_1852);
or U5542 (N_5542,N_148,N_2999);
nor U5543 (N_5543,N_1862,N_4918);
xor U5544 (N_5544,N_4304,N_3804);
nand U5545 (N_5545,N_1363,N_849);
nand U5546 (N_5546,N_2494,N_2841);
or U5547 (N_5547,N_2990,N_4324);
or U5548 (N_5548,N_4047,N_1459);
nand U5549 (N_5549,N_3249,N_4393);
nand U5550 (N_5550,N_4437,N_4174);
and U5551 (N_5551,N_4910,N_3831);
or U5552 (N_5552,N_4791,N_2854);
xnor U5553 (N_5553,N_2874,N_635);
and U5554 (N_5554,N_3502,N_2321);
nand U5555 (N_5555,N_1063,N_2844);
and U5556 (N_5556,N_1150,N_1223);
or U5557 (N_5557,N_4107,N_4823);
nor U5558 (N_5558,N_3170,N_4157);
xor U5559 (N_5559,N_1447,N_3191);
or U5560 (N_5560,N_740,N_1079);
nand U5561 (N_5561,N_118,N_2814);
or U5562 (N_5562,N_137,N_4017);
xnor U5563 (N_5563,N_4197,N_3150);
xor U5564 (N_5564,N_227,N_1938);
and U5565 (N_5565,N_4526,N_693);
or U5566 (N_5566,N_652,N_239);
and U5567 (N_5567,N_364,N_3980);
xor U5568 (N_5568,N_506,N_2253);
nand U5569 (N_5569,N_685,N_3465);
and U5570 (N_5570,N_4379,N_3039);
nand U5571 (N_5571,N_4141,N_4627);
xor U5572 (N_5572,N_3955,N_1587);
xnor U5573 (N_5573,N_4231,N_4913);
xor U5574 (N_5574,N_1581,N_3028);
nor U5575 (N_5575,N_4395,N_25);
nand U5576 (N_5576,N_701,N_4769);
nor U5577 (N_5577,N_3861,N_2529);
xor U5578 (N_5578,N_3213,N_3327);
or U5579 (N_5579,N_2097,N_1381);
nor U5580 (N_5580,N_3723,N_2862);
nand U5581 (N_5581,N_3083,N_1106);
and U5582 (N_5582,N_2804,N_699);
nand U5583 (N_5583,N_828,N_3578);
and U5584 (N_5584,N_2540,N_3795);
or U5585 (N_5585,N_521,N_657);
xor U5586 (N_5586,N_1717,N_1451);
xnor U5587 (N_5587,N_2013,N_226);
or U5588 (N_5588,N_1895,N_3342);
nand U5589 (N_5589,N_4037,N_871);
nor U5590 (N_5590,N_3600,N_840);
nand U5591 (N_5591,N_705,N_2769);
and U5592 (N_5592,N_4859,N_4358);
xor U5593 (N_5593,N_358,N_4527);
nand U5594 (N_5594,N_1136,N_1813);
or U5595 (N_5595,N_709,N_2940);
nand U5596 (N_5596,N_3844,N_4397);
and U5597 (N_5597,N_2711,N_94);
and U5598 (N_5598,N_4613,N_447);
xor U5599 (N_5599,N_2262,N_2879);
xnor U5600 (N_5600,N_3937,N_2470);
xor U5601 (N_5601,N_3504,N_2393);
or U5602 (N_5602,N_1995,N_3653);
or U5603 (N_5603,N_1097,N_1175);
and U5604 (N_5604,N_1824,N_4374);
nand U5605 (N_5605,N_4406,N_4121);
xor U5606 (N_5606,N_4565,N_3921);
and U5607 (N_5607,N_2531,N_3399);
nand U5608 (N_5608,N_634,N_2957);
and U5609 (N_5609,N_211,N_3396);
xor U5610 (N_5610,N_4756,N_448);
and U5611 (N_5611,N_3990,N_1069);
nand U5612 (N_5612,N_800,N_4098);
nand U5613 (N_5613,N_1436,N_3901);
nand U5614 (N_5614,N_2409,N_4130);
xnor U5615 (N_5615,N_3051,N_1350);
xor U5616 (N_5616,N_3902,N_2035);
and U5617 (N_5617,N_3495,N_1751);
nand U5618 (N_5618,N_333,N_383);
nor U5619 (N_5619,N_2437,N_1855);
or U5620 (N_5620,N_4765,N_1391);
or U5621 (N_5621,N_1320,N_3672);
xor U5622 (N_5622,N_4896,N_4367);
nor U5623 (N_5623,N_4057,N_2004);
nor U5624 (N_5624,N_3265,N_4895);
nand U5625 (N_5625,N_3889,N_4167);
xor U5626 (N_5626,N_2528,N_2856);
and U5627 (N_5627,N_4080,N_2752);
and U5628 (N_5628,N_231,N_1145);
or U5629 (N_5629,N_1170,N_3218);
nand U5630 (N_5630,N_2237,N_1611);
nand U5631 (N_5631,N_2028,N_128);
or U5632 (N_5632,N_4432,N_4534);
xnor U5633 (N_5633,N_523,N_2376);
and U5634 (N_5634,N_2389,N_1808);
and U5635 (N_5635,N_1794,N_1066);
and U5636 (N_5636,N_482,N_4601);
xor U5637 (N_5637,N_884,N_1854);
nor U5638 (N_5638,N_2332,N_2664);
nand U5639 (N_5639,N_2478,N_4131);
nand U5640 (N_5640,N_169,N_1178);
nor U5641 (N_5641,N_4829,N_1444);
nand U5642 (N_5642,N_598,N_1675);
xnor U5643 (N_5643,N_3650,N_4541);
nand U5644 (N_5644,N_564,N_4804);
xor U5645 (N_5645,N_3402,N_1312);
nand U5646 (N_5646,N_2975,N_150);
and U5647 (N_5647,N_2545,N_1217);
xor U5648 (N_5648,N_747,N_2754);
nand U5649 (N_5649,N_2061,N_4746);
nor U5650 (N_5650,N_4218,N_2360);
nand U5651 (N_5651,N_3782,N_4933);
nand U5652 (N_5652,N_2245,N_4287);
and U5653 (N_5653,N_1033,N_1801);
nand U5654 (N_5654,N_1733,N_4624);
nand U5655 (N_5655,N_4249,N_2220);
xor U5656 (N_5656,N_609,N_2159);
nor U5657 (N_5657,N_3919,N_2252);
nor U5658 (N_5658,N_2500,N_4840);
nand U5659 (N_5659,N_4463,N_1649);
and U5660 (N_5660,N_4655,N_1617);
or U5661 (N_5661,N_1580,N_3924);
or U5662 (N_5662,N_3623,N_2461);
or U5663 (N_5663,N_4089,N_4142);
or U5664 (N_5664,N_2938,N_3065);
and U5665 (N_5665,N_3665,N_1534);
or U5666 (N_5666,N_3002,N_4413);
or U5667 (N_5667,N_3287,N_1922);
or U5668 (N_5668,N_2810,N_1859);
nor U5669 (N_5669,N_3983,N_4568);
and U5670 (N_5670,N_1289,N_2743);
and U5671 (N_5671,N_4159,N_4872);
and U5672 (N_5672,N_3886,N_4770);
and U5673 (N_5673,N_4070,N_834);
and U5674 (N_5674,N_105,N_1776);
nor U5675 (N_5675,N_818,N_3441);
xor U5676 (N_5676,N_3821,N_3703);
xor U5677 (N_5677,N_1202,N_4795);
nand U5678 (N_5678,N_2855,N_4363);
or U5679 (N_5679,N_1818,N_320);
nor U5680 (N_5680,N_645,N_3324);
nor U5681 (N_5681,N_4768,N_1390);
nor U5682 (N_5682,N_1775,N_1110);
nand U5683 (N_5683,N_3291,N_2514);
xor U5684 (N_5684,N_2269,N_892);
and U5685 (N_5685,N_158,N_3594);
xnor U5686 (N_5686,N_3,N_643);
and U5687 (N_5687,N_1657,N_3891);
xnor U5688 (N_5688,N_824,N_1702);
or U5689 (N_5689,N_1025,N_2881);
and U5690 (N_5690,N_4442,N_2878);
nor U5691 (N_5691,N_2263,N_3606);
xor U5692 (N_5692,N_2598,N_4719);
or U5693 (N_5693,N_1292,N_2958);
xor U5694 (N_5694,N_4323,N_4867);
nor U5695 (N_5695,N_759,N_1435);
or U5696 (N_5696,N_4018,N_3852);
nand U5697 (N_5697,N_3871,N_2919);
nor U5698 (N_5698,N_780,N_2129);
and U5699 (N_5699,N_1637,N_1014);
xnor U5700 (N_5700,N_2212,N_2098);
and U5701 (N_5701,N_868,N_1946);
xnor U5702 (N_5702,N_1845,N_2631);
nor U5703 (N_5703,N_2865,N_832);
and U5704 (N_5704,N_95,N_4538);
nor U5705 (N_5705,N_2031,N_4315);
nor U5706 (N_5706,N_3965,N_4576);
nand U5707 (N_5707,N_571,N_1236);
xnor U5708 (N_5708,N_3113,N_3244);
nor U5709 (N_5709,N_4873,N_3544);
xor U5710 (N_5710,N_2425,N_2823);
xor U5711 (N_5711,N_180,N_3740);
nor U5712 (N_5712,N_4366,N_72);
nand U5713 (N_5713,N_4326,N_3460);
and U5714 (N_5714,N_3185,N_1937);
xnor U5715 (N_5715,N_4283,N_434);
or U5716 (N_5716,N_3006,N_610);
nor U5717 (N_5717,N_1887,N_3885);
nor U5718 (N_5718,N_568,N_4021);
or U5719 (N_5719,N_2002,N_1956);
and U5720 (N_5720,N_4718,N_3115);
or U5721 (N_5721,N_2625,N_4508);
nand U5722 (N_5722,N_222,N_458);
nand U5723 (N_5723,N_1491,N_4354);
and U5724 (N_5724,N_4161,N_2298);
nor U5725 (N_5725,N_2898,N_3754);
xnor U5726 (N_5726,N_3464,N_4071);
nor U5727 (N_5727,N_1309,N_4816);
xnor U5728 (N_5728,N_4040,N_2614);
nand U5729 (N_5729,N_216,N_1696);
or U5730 (N_5730,N_1121,N_3467);
or U5731 (N_5731,N_2264,N_3555);
nor U5732 (N_5732,N_2082,N_1746);
nor U5733 (N_5733,N_1016,N_4496);
nor U5734 (N_5734,N_4433,N_4045);
and U5735 (N_5735,N_2167,N_1094);
or U5736 (N_5736,N_2119,N_3994);
nand U5737 (N_5737,N_4475,N_4078);
nor U5738 (N_5738,N_4745,N_4739);
nor U5739 (N_5739,N_18,N_2506);
and U5740 (N_5740,N_1850,N_2139);
or U5741 (N_5741,N_2388,N_3047);
and U5742 (N_5742,N_3827,N_4519);
or U5743 (N_5743,N_3190,N_220);
nand U5744 (N_5744,N_4793,N_2692);
or U5745 (N_5745,N_2080,N_1075);
and U5746 (N_5746,N_4369,N_1589);
xor U5747 (N_5747,N_676,N_2636);
xnor U5748 (N_5748,N_4230,N_1863);
or U5749 (N_5749,N_1708,N_2618);
nand U5750 (N_5750,N_4962,N_4248);
xor U5751 (N_5751,N_3823,N_4213);
nand U5752 (N_5752,N_4422,N_2732);
and U5753 (N_5753,N_4731,N_3121);
and U5754 (N_5754,N_2757,N_2010);
and U5755 (N_5755,N_636,N_2602);
or U5756 (N_5756,N_4845,N_3373);
and U5757 (N_5757,N_2408,N_452);
nand U5758 (N_5758,N_1912,N_3614);
or U5759 (N_5759,N_1520,N_1429);
nand U5760 (N_5760,N_4385,N_1041);
nand U5761 (N_5761,N_2278,N_603);
nand U5762 (N_5762,N_3397,N_151);
nand U5763 (N_5763,N_2496,N_3643);
xnor U5764 (N_5764,N_225,N_2706);
and U5765 (N_5765,N_1281,N_865);
xnor U5766 (N_5766,N_4513,N_44);
xnor U5767 (N_5767,N_2094,N_2042);
xnor U5768 (N_5768,N_1248,N_2135);
nand U5769 (N_5769,N_388,N_4546);
nand U5770 (N_5770,N_195,N_4955);
or U5771 (N_5771,N_4477,N_620);
xnor U5772 (N_5772,N_3770,N_4069);
nor U5773 (N_5773,N_245,N_4001);
nand U5774 (N_5774,N_3866,N_3346);
xnor U5775 (N_5775,N_2570,N_1870);
xnor U5776 (N_5776,N_660,N_651);
xnor U5777 (N_5777,N_1815,N_4389);
xor U5778 (N_5778,N_1958,N_1056);
xor U5779 (N_5779,N_1141,N_73);
or U5780 (N_5780,N_314,N_252);
nor U5781 (N_5781,N_411,N_573);
nor U5782 (N_5782,N_4146,N_3779);
xor U5783 (N_5783,N_2380,N_4717);
or U5784 (N_5784,N_2951,N_30);
xnor U5785 (N_5785,N_4462,N_1326);
nor U5786 (N_5786,N_3566,N_2238);
and U5787 (N_5787,N_716,N_467);
xnor U5788 (N_5788,N_2585,N_1021);
nand U5789 (N_5789,N_147,N_2344);
nor U5790 (N_5790,N_4636,N_27);
nand U5791 (N_5791,N_4327,N_2044);
nor U5792 (N_5792,N_2800,N_461);
and U5793 (N_5793,N_2446,N_4150);
xor U5794 (N_5794,N_1670,N_4260);
nand U5795 (N_5795,N_3010,N_3869);
nor U5796 (N_5796,N_3316,N_4171);
nand U5797 (N_5797,N_2712,N_432);
xor U5798 (N_5798,N_3061,N_4759);
nand U5799 (N_5799,N_2150,N_421);
nand U5800 (N_5800,N_988,N_853);
nand U5801 (N_5801,N_4290,N_3433);
xor U5802 (N_5802,N_1258,N_2289);
or U5803 (N_5803,N_3027,N_955);
nand U5804 (N_5804,N_1477,N_586);
nor U5805 (N_5805,N_2617,N_1663);
or U5806 (N_5806,N_486,N_28);
nor U5807 (N_5807,N_4579,N_3579);
xnor U5808 (N_5808,N_3319,N_481);
nor U5809 (N_5809,N_3438,N_1728);
and U5810 (N_5810,N_2493,N_4154);
nand U5811 (N_5811,N_256,N_2715);
or U5812 (N_5812,N_1218,N_4713);
and U5813 (N_5813,N_4600,N_2319);
nor U5814 (N_5814,N_4941,N_4850);
nor U5815 (N_5815,N_1973,N_2731);
nand U5816 (N_5816,N_2546,N_3377);
nand U5817 (N_5817,N_4295,N_2084);
xnor U5818 (N_5818,N_431,N_1274);
and U5819 (N_5819,N_3708,N_1388);
or U5820 (N_5820,N_4521,N_2770);
xor U5821 (N_5821,N_1976,N_4337);
xor U5822 (N_5822,N_938,N_1721);
nand U5823 (N_5823,N_4091,N_3224);
and U5824 (N_5824,N_1346,N_1226);
or U5825 (N_5825,N_1598,N_3585);
and U5826 (N_5826,N_3276,N_355);
or U5827 (N_5827,N_542,N_3744);
xor U5828 (N_5828,N_4439,N_4659);
and U5829 (N_5829,N_4246,N_2760);
or U5830 (N_5830,N_2242,N_1980);
or U5831 (N_5831,N_1067,N_4532);
or U5832 (N_5832,N_789,N_3835);
nand U5833 (N_5833,N_4874,N_4964);
nand U5834 (N_5834,N_463,N_2421);
or U5835 (N_5835,N_3966,N_1519);
nor U5836 (N_5836,N_3819,N_3275);
nand U5837 (N_5837,N_4844,N_3967);
and U5838 (N_5838,N_3026,N_1221);
nand U5839 (N_5839,N_1986,N_4978);
xnor U5840 (N_5840,N_4123,N_3664);
nor U5841 (N_5841,N_511,N_4398);
nand U5842 (N_5842,N_1584,N_1904);
xnor U5843 (N_5843,N_901,N_2239);
or U5844 (N_5844,N_3915,N_1430);
nor U5845 (N_5845,N_2550,N_3883);
or U5846 (N_5846,N_2199,N_1822);
or U5847 (N_5847,N_4657,N_3333);
nor U5848 (N_5848,N_4886,N_2315);
and U5849 (N_5849,N_1495,N_2606);
nand U5850 (N_5850,N_2091,N_2165);
and U5851 (N_5851,N_2381,N_2491);
nand U5852 (N_5852,N_4689,N_292);
or U5853 (N_5853,N_477,N_3808);
nor U5854 (N_5854,N_1913,N_4104);
nor U5855 (N_5855,N_2637,N_4675);
and U5856 (N_5856,N_1510,N_2641);
nor U5857 (N_5857,N_2564,N_3511);
and U5858 (N_5858,N_2218,N_4355);
or U5859 (N_5859,N_1304,N_1188);
nor U5860 (N_5860,N_4409,N_3776);
or U5861 (N_5861,N_1765,N_3149);
xnor U5862 (N_5862,N_1107,N_2768);
nor U5863 (N_5863,N_1650,N_3864);
nand U5864 (N_5864,N_3007,N_950);
or U5865 (N_5865,N_778,N_1488);
nand U5866 (N_5866,N_3044,N_644);
nor U5867 (N_5867,N_3549,N_3023);
nor U5868 (N_5868,N_794,N_3314);
or U5869 (N_5869,N_2083,N_775);
and U5870 (N_5870,N_2953,N_4906);
or U5871 (N_5871,N_1609,N_1499);
and U5872 (N_5872,N_2048,N_2669);
xor U5873 (N_5873,N_1882,N_4114);
and U5874 (N_5874,N_2730,N_3270);
nor U5875 (N_5875,N_1118,N_3144);
and U5876 (N_5876,N_1192,N_860);
xor U5877 (N_5877,N_1342,N_4786);
xor U5878 (N_5878,N_3586,N_562);
xor U5879 (N_5879,N_2166,N_1389);
nor U5880 (N_5880,N_1525,N_1394);
and U5881 (N_5881,N_4403,N_3560);
nor U5882 (N_5882,N_4779,N_1095);
nor U5883 (N_5883,N_2673,N_2569);
nor U5884 (N_5884,N_3559,N_4296);
nor U5885 (N_5885,N_2187,N_1099);
nand U5886 (N_5886,N_2560,N_4183);
and U5887 (N_5887,N_1939,N_3741);
xnor U5888 (N_5888,N_2467,N_3763);
or U5889 (N_5889,N_470,N_792);
or U5890 (N_5890,N_1553,N_718);
xor U5891 (N_5891,N_1713,N_730);
and U5892 (N_5892,N_2508,N_4074);
and U5893 (N_5893,N_3344,N_2824);
or U5894 (N_5894,N_404,N_3805);
or U5895 (N_5895,N_1678,N_977);
or U5896 (N_5896,N_2914,N_99);
and U5897 (N_5897,N_4454,N_1074);
or U5898 (N_5898,N_4628,N_3173);
nor U5899 (N_5899,N_2588,N_3893);
or U5900 (N_5900,N_196,N_1054);
xnor U5901 (N_5901,N_387,N_4837);
and U5902 (N_5902,N_3442,N_637);
nand U5903 (N_5903,N_4728,N_3417);
and U5904 (N_5904,N_1991,N_2527);
nor U5905 (N_5905,N_3131,N_3591);
or U5906 (N_5906,N_648,N_1603);
nor U5907 (N_5907,N_3160,N_1251);
or U5908 (N_5908,N_2869,N_932);
nand U5909 (N_5909,N_33,N_4651);
xor U5910 (N_5910,N_1560,N_3524);
nand U5911 (N_5911,N_4503,N_1779);
and U5912 (N_5912,N_1353,N_170);
and U5913 (N_5913,N_4191,N_2907);
xor U5914 (N_5914,N_558,N_4680);
or U5915 (N_5915,N_2813,N_3049);
or U5916 (N_5916,N_1853,N_449);
nor U5917 (N_5917,N_1931,N_1536);
or U5918 (N_5918,N_1115,N_4238);
nand U5919 (N_5919,N_3978,N_1135);
and U5920 (N_5920,N_3014,N_945);
and U5921 (N_5921,N_3616,N_2085);
xor U5922 (N_5922,N_2366,N_2783);
or U5923 (N_5923,N_4076,N_2345);
xor U5924 (N_5924,N_1694,N_3050);
and U5925 (N_5925,N_234,N_240);
or U5926 (N_5926,N_3601,N_75);
nor U5927 (N_5927,N_4712,N_1020);
nor U5928 (N_5928,N_3330,N_1635);
and U5929 (N_5929,N_3888,N_1152);
and U5930 (N_5930,N_1176,N_4509);
nand U5931 (N_5931,N_3691,N_4752);
xnor U5932 (N_5932,N_207,N_2249);
nand U5933 (N_5933,N_4396,N_2201);
xnor U5934 (N_5934,N_748,N_4187);
nand U5935 (N_5935,N_2023,N_244);
nor U5936 (N_5936,N_2196,N_3533);
nand U5937 (N_5937,N_1028,N_4097);
nand U5938 (N_5938,N_540,N_691);
nand U5939 (N_5939,N_3208,N_3040);
or U5940 (N_5940,N_2561,N_2276);
and U5941 (N_5941,N_190,N_680);
nor U5942 (N_5942,N_694,N_768);
nor U5943 (N_5943,N_2426,N_4929);
nand U5944 (N_5944,N_4266,N_4650);
or U5945 (N_5945,N_3879,N_1880);
nand U5946 (N_5946,N_4892,N_315);
nand U5947 (N_5947,N_3479,N_3165);
or U5948 (N_5948,N_554,N_278);
nand U5949 (N_5949,N_561,N_4158);
nor U5950 (N_5950,N_872,N_3459);
and U5951 (N_5951,N_1970,N_2665);
nor U5952 (N_5952,N_4391,N_253);
nor U5953 (N_5953,N_1241,N_4208);
and U5954 (N_5954,N_444,N_2162);
or U5955 (N_5955,N_1482,N_2857);
nor U5956 (N_5956,N_4501,N_3855);
or U5957 (N_5957,N_4830,N_3008);
nor U5958 (N_5958,N_3816,N_4922);
or U5959 (N_5959,N_440,N_1768);
xnor U5960 (N_5960,N_1674,N_2224);
xnor U5961 (N_5961,N_3942,N_553);
or U5962 (N_5962,N_4796,N_1091);
or U5963 (N_5963,N_3558,N_183);
nor U5964 (N_5964,N_3968,N_3930);
nand U5965 (N_5965,N_986,N_1898);
and U5966 (N_5966,N_64,N_4032);
or U5967 (N_5967,N_1232,N_3338);
nand U5968 (N_5968,N_3296,N_2177);
nand U5969 (N_5969,N_592,N_3473);
nor U5970 (N_5970,N_3153,N_1373);
nand U5971 (N_5971,N_4113,N_2116);
or U5972 (N_5972,N_2189,N_2955);
xor U5973 (N_5973,N_2922,N_1360);
xor U5974 (N_5974,N_2175,N_2628);
and U5975 (N_5975,N_283,N_2780);
xor U5976 (N_5976,N_4328,N_4530);
xor U5977 (N_5977,N_4652,N_1369);
nand U5978 (N_5978,N_2791,N_3592);
and U5979 (N_5979,N_4951,N_904);
or U5980 (N_5980,N_3132,N_4773);
nand U5981 (N_5981,N_3834,N_3995);
or U5982 (N_5982,N_2693,N_1406);
nor U5983 (N_5983,N_422,N_551);
nor U5984 (N_5984,N_3536,N_4902);
nor U5985 (N_5985,N_4059,N_640);
and U5986 (N_5986,N_4724,N_1355);
and U5987 (N_5987,N_4616,N_111);
or U5988 (N_5988,N_1985,N_1561);
nor U5989 (N_5989,N_4073,N_744);
xnor U5990 (N_5990,N_3693,N_282);
and U5991 (N_5991,N_1957,N_402);
and U5992 (N_5992,N_209,N_1655);
nand U5993 (N_5993,N_3764,N_286);
or U5994 (N_5994,N_3812,N_1947);
nor U5995 (N_5995,N_3128,N_1629);
xor U5996 (N_5996,N_3929,N_2215);
or U5997 (N_5997,N_3535,N_2566);
and U5998 (N_5998,N_1301,N_4233);
xor U5999 (N_5999,N_4959,N_2651);
nand U6000 (N_6000,N_1737,N_2822);
or U6001 (N_6001,N_4221,N_1393);
and U6002 (N_6002,N_471,N_2087);
and U6003 (N_6003,N_3985,N_1761);
xnor U6004 (N_6004,N_4291,N_82);
or U6005 (N_6005,N_3984,N_4865);
nand U6006 (N_6006,N_1273,N_4348);
xnor U6007 (N_6007,N_4459,N_4312);
or U6008 (N_6008,N_4298,N_1744);
or U6009 (N_6009,N_2723,N_1547);
and U6010 (N_6010,N_450,N_4700);
xor U6011 (N_6011,N_1315,N_3492);
xor U6012 (N_6012,N_274,N_4544);
nand U6013 (N_6013,N_2620,N_1288);
xor U6014 (N_6014,N_2716,N_246);
or U6015 (N_6015,N_1810,N_2640);
and U6016 (N_6016,N_2265,N_4392);
xnor U6017 (N_6017,N_4430,N_2134);
and U6018 (N_6018,N_3710,N_332);
nand U6019 (N_6019,N_265,N_4253);
nand U6020 (N_6020,N_4743,N_2100);
nand U6021 (N_6021,N_1322,N_935);
nor U6022 (N_6022,N_248,N_1356);
nor U6023 (N_6023,N_2018,N_2737);
nand U6024 (N_6024,N_547,N_594);
nor U6025 (N_6025,N_3507,N_4336);
and U6026 (N_6026,N_3159,N_4111);
nand U6027 (N_6027,N_371,N_851);
xor U6028 (N_6028,N_2328,N_403);
or U6029 (N_6029,N_4664,N_3542);
and U6030 (N_6030,N_1739,N_2998);
nand U6031 (N_6031,N_764,N_2672);
and U6032 (N_6032,N_1719,N_4316);
xnor U6033 (N_6033,N_627,N_2785);
and U6034 (N_6034,N_1962,N_1722);
nand U6035 (N_6035,N_2968,N_4294);
nor U6036 (N_6036,N_2051,N_3627);
nor U6037 (N_6037,N_4725,N_837);
and U6038 (N_6038,N_4472,N_719);
nor U6039 (N_6039,N_4309,N_3590);
xor U6040 (N_6040,N_3787,N_1407);
or U6041 (N_6041,N_229,N_485);
nor U6042 (N_6042,N_1187,N_2748);
and U6043 (N_6043,N_4273,N_4847);
and U6044 (N_6044,N_464,N_79);
xnor U6045 (N_6045,N_2005,N_3595);
nor U6046 (N_6046,N_2977,N_3250);
and U6047 (N_6047,N_3923,N_4709);
nand U6048 (N_6048,N_205,N_4168);
and U6049 (N_6049,N_1076,N_954);
xnor U6050 (N_6050,N_3013,N_1600);
nor U6051 (N_6051,N_4067,N_2451);
or U6052 (N_6052,N_108,N_2458);
nor U6053 (N_6053,N_4620,N_3406);
nand U6054 (N_6054,N_951,N_591);
or U6055 (N_6055,N_2864,N_3468);
or U6056 (N_6056,N_4415,N_3425);
nand U6057 (N_6057,N_3849,N_2548);
nand U6058 (N_6058,N_4575,N_3042);
nand U6059 (N_6059,N_3361,N_3521);
nor U6060 (N_6060,N_1421,N_3796);
or U6061 (N_6061,N_981,N_2629);
and U6062 (N_6062,N_4384,N_969);
nand U6063 (N_6063,N_4808,N_3954);
nor U6064 (N_6064,N_1216,N_2612);
or U6065 (N_6065,N_417,N_4418);
xor U6066 (N_6066,N_2551,N_3925);
nand U6067 (N_6067,N_4151,N_2985);
nor U6068 (N_6068,N_4661,N_2744);
nor U6069 (N_6069,N_4278,N_3759);
nand U6070 (N_6070,N_3235,N_1468);
nand U6071 (N_6071,N_618,N_2633);
nor U6072 (N_6072,N_2110,N_16);
and U6073 (N_6073,N_4030,N_684);
and U6074 (N_6074,N_2875,N_1527);
and U6075 (N_6075,N_2208,N_2960);
nor U6076 (N_6076,N_3851,N_863);
nand U6077 (N_6077,N_2935,N_3390);
and U6078 (N_6078,N_2054,N_3161);
nor U6079 (N_6079,N_410,N_1623);
or U6080 (N_6080,N_4132,N_3728);
nand U6081 (N_6081,N_3647,N_1464);
xor U6082 (N_6082,N_1848,N_641);
nand U6083 (N_6083,N_4178,N_1173);
and U6084 (N_6084,N_3053,N_537);
or U6085 (N_6085,N_154,N_2138);
nor U6086 (N_6086,N_2062,N_465);
or U6087 (N_6087,N_330,N_814);
or U6088 (N_6088,N_3059,N_4350);
xor U6089 (N_6089,N_3939,N_460);
nand U6090 (N_6090,N_2622,N_307);
xor U6091 (N_6091,N_4426,N_2308);
and U6092 (N_6092,N_3506,N_1070);
xnor U6093 (N_6093,N_720,N_2055);
nor U6094 (N_6094,N_2072,N_406);
and U6095 (N_6095,N_3607,N_887);
nand U6096 (N_6096,N_1714,N_880);
or U6097 (N_6097,N_3001,N_3998);
nand U6098 (N_6098,N_3230,N_976);
and U6099 (N_6099,N_3575,N_3070);
and U6100 (N_6100,N_2155,N_2608);
and U6101 (N_6101,N_2324,N_1987);
and U6102 (N_6102,N_4658,N_2733);
nand U6103 (N_6103,N_1029,N_3313);
xor U6104 (N_6104,N_2447,N_3229);
and U6105 (N_6105,N_655,N_1310);
nand U6106 (N_6106,N_784,N_3494);
nor U6107 (N_6107,N_129,N_4897);
nand U6108 (N_6108,N_4140,N_1982);
xnor U6109 (N_6109,N_662,N_3727);
nand U6110 (N_6110,N_2399,N_3694);
nor U6111 (N_6111,N_4714,N_3568);
nor U6112 (N_6112,N_1297,N_3872);
and U6113 (N_6113,N_913,N_555);
and U6114 (N_6114,N_1300,N_3784);
or U6115 (N_6115,N_3435,N_4214);
and U6116 (N_6116,N_3303,N_2338);
nand U6117 (N_6117,N_2610,N_4839);
xor U6118 (N_6118,N_4048,N_3906);
xor U6119 (N_6119,N_4748,N_3509);
nand U6120 (N_6120,N_1238,N_3129);
xnor U6121 (N_6121,N_773,N_4543);
and U6122 (N_6122,N_251,N_4075);
nor U6123 (N_6123,N_189,N_3353);
xor U6124 (N_6124,N_3557,N_2835);
xor U6125 (N_6125,N_4798,N_117);
or U6126 (N_6126,N_4875,N_3810);
and U6127 (N_6127,N_933,N_1640);
or U6128 (N_6128,N_2323,N_4924);
or U6129 (N_6129,N_1212,N_277);
and U6130 (N_6130,N_2070,N_2333);
and U6131 (N_6131,N_2086,N_4934);
or U6132 (N_6132,N_1673,N_2536);
nand U6133 (N_6133,N_682,N_1526);
nor U6134 (N_6134,N_516,N_113);
or U6135 (N_6135,N_2120,N_413);
and U6136 (N_6136,N_3712,N_1453);
or U6137 (N_6137,N_3133,N_3060);
and U6138 (N_6138,N_3666,N_3803);
or U6139 (N_6139,N_1286,N_3087);
xor U6140 (N_6140,N_1365,N_738);
and U6141 (N_6141,N_2784,N_1802);
xnor U6142 (N_6142,N_2232,N_3979);
and U6143 (N_6143,N_4,N_937);
or U6144 (N_6144,N_3110,N_4345);
nor U6145 (N_6145,N_1729,N_1823);
or U6146 (N_6146,N_43,N_2890);
and U6147 (N_6147,N_2834,N_1261);
nand U6148 (N_6148,N_204,N_2390);
and U6149 (N_6149,N_4265,N_4490);
nand U6150 (N_6150,N_260,N_611);
nor U6151 (N_6151,N_4707,N_2872);
or U6152 (N_6152,N_3046,N_4566);
and U6153 (N_6153,N_3948,N_4722);
nor U6154 (N_6154,N_3217,N_3932);
nand U6155 (N_6155,N_3752,N_4079);
and U6156 (N_6156,N_3401,N_1003);
nor U6157 (N_6157,N_4137,N_2901);
or U6158 (N_6158,N_1144,N_3209);
and U6159 (N_6159,N_4871,N_4852);
xnor U6160 (N_6160,N_712,N_596);
nor U6161 (N_6161,N_2831,N_2147);
and U6162 (N_6162,N_3030,N_4948);
nand U6163 (N_6163,N_3552,N_218);
and U6164 (N_6164,N_2782,N_4685);
and U6165 (N_6165,N_1700,N_3409);
or U6166 (N_6166,N_4448,N_4492);
xnor U6167 (N_6167,N_1022,N_462);
xor U6168 (N_6168,N_3532,N_882);
xor U6169 (N_6169,N_3977,N_4160);
xor U6170 (N_6170,N_535,N_4932);
nor U6171 (N_6171,N_2277,N_102);
nor U6172 (N_6172,N_3386,N_507);
and U6173 (N_6173,N_3621,N_1864);
xnor U6174 (N_6174,N_1180,N_536);
nand U6175 (N_6175,N_2686,N_4308);
or U6176 (N_6176,N_4026,N_4879);
nand U6177 (N_6177,N_3394,N_4754);
nand U6178 (N_6178,N_4102,N_3206);
nor U6179 (N_6179,N_4473,N_71);
or U6180 (N_6180,N_1048,N_4056);
or U6181 (N_6181,N_2144,N_2193);
and U6182 (N_6182,N_2429,N_4302);
or U6183 (N_6183,N_1296,N_912);
nand U6184 (N_6184,N_1833,N_2131);
nand U6185 (N_6185,N_3090,N_4163);
nand U6186 (N_6186,N_3404,N_3721);
xor U6187 (N_6187,N_3391,N_2891);
xnor U6188 (N_6188,N_3440,N_1347);
nand U6189 (N_6189,N_2296,N_766);
nand U6190 (N_6190,N_275,N_2452);
and U6191 (N_6191,N_4694,N_3095);
or U6192 (N_6192,N_1329,N_2396);
nand U6193 (N_6193,N_2304,N_3130);
nand U6194 (N_6194,N_3785,N_4957);
xor U6195 (N_6195,N_1470,N_2703);
and U6196 (N_6196,N_4244,N_1615);
nor U6197 (N_6197,N_2015,N_2884);
xnor U6198 (N_6198,N_4262,N_2504);
or U6199 (N_6199,N_3357,N_4584);
nand U6200 (N_6200,N_1760,N_2979);
and U6201 (N_6201,N_2219,N_4043);
or U6202 (N_6202,N_1846,N_4275);
or U6203 (N_6203,N_990,N_65);
nand U6204 (N_6204,N_2330,N_3873);
and U6205 (N_6205,N_3194,N_2039);
nand U6206 (N_6206,N_1645,N_4736);
nor U6207 (N_6207,N_2418,N_1290);
or U6208 (N_6208,N_114,N_478);
nor U6209 (N_6209,N_1448,N_2604);
xnor U6210 (N_6210,N_1011,N_2411);
nand U6211 (N_6211,N_4094,N_1037);
and U6212 (N_6212,N_4734,N_1279);
xor U6213 (N_6213,N_2656,N_3012);
or U6214 (N_6214,N_2965,N_1935);
or U6215 (N_6215,N_4344,N_1601);
and U6216 (N_6216,N_4708,N_3904);
and U6217 (N_6217,N_2929,N_670);
or U6218 (N_6218,N_4536,N_4916);
xnor U6219 (N_6219,N_2294,N_2071);
nor U6220 (N_6220,N_2256,N_1920);
or U6221 (N_6221,N_1807,N_2605);
xor U6222 (N_6222,N_1858,N_668);
xnor U6223 (N_6223,N_650,N_4912);
xor U6224 (N_6224,N_2509,N_1971);
xor U6225 (N_6225,N_87,N_2659);
nor U6226 (N_6226,N_4588,N_1889);
and U6227 (N_6227,N_1004,N_3148);
xnor U6228 (N_6228,N_994,N_2713);
or U6229 (N_6229,N_2361,N_2635);
xnor U6230 (N_6230,N_1959,N_3350);
nand U6231 (N_6231,N_284,N_3286);
nand U6232 (N_6232,N_3649,N_4349);
nand U6233 (N_6233,N_1654,N_2106);
and U6234 (N_6234,N_2817,N_281);
and U6235 (N_6235,N_398,N_3094);
or U6236 (N_6236,N_3135,N_1955);
nand U6237 (N_6237,N_3789,N_3892);
xnor U6238 (N_6238,N_1844,N_783);
nor U6239 (N_6239,N_2217,N_342);
or U6240 (N_6240,N_1503,N_1374);
nor U6241 (N_6241,N_4862,N_2267);
and U6242 (N_6242,N_4192,N_588);
nor U6243 (N_6243,N_3392,N_3372);
nand U6244 (N_6244,N_2724,N_3989);
and U6245 (N_6245,N_3477,N_4011);
xnor U6246 (N_6246,N_1253,N_2462);
or U6247 (N_6247,N_2750,N_2763);
nor U6248 (N_6248,N_4357,N_2928);
nand U6249 (N_6249,N_1230,N_4004);
nor U6250 (N_6250,N_29,N_356);
xnor U6251 (N_6251,N_1847,N_1283);
xor U6252 (N_6252,N_1689,N_212);
nor U6253 (N_6253,N_1927,N_3033);
xnor U6254 (N_6254,N_4673,N_2268);
nand U6255 (N_6255,N_758,N_390);
and U6256 (N_6256,N_1630,N_4617);
and U6257 (N_6257,N_2615,N_243);
nor U6258 (N_6258,N_2060,N_2373);
or U6259 (N_6259,N_2200,N_3836);
xnor U6260 (N_6260,N_585,N_451);
xor U6261 (N_6261,N_3105,N_1804);
nand U6262 (N_6262,N_3328,N_2257);
nor U6263 (N_6263,N_60,N_2079);
or U6264 (N_6264,N_2674,N_290);
nor U6265 (N_6265,N_1546,N_288);
nor U6266 (N_6266,N_110,N_2244);
xor U6267 (N_6267,N_4988,N_617);
or U6268 (N_6268,N_2971,N_4449);
nand U6269 (N_6269,N_745,N_2858);
nand U6270 (N_6270,N_3840,N_3352);
xnor U6271 (N_6271,N_2671,N_4784);
and U6272 (N_6272,N_3212,N_4596);
xnor U6273 (N_6273,N_14,N_1375);
nor U6274 (N_6274,N_1979,N_4775);
nor U6275 (N_6275,N_1693,N_3514);
and U6276 (N_6276,N_1163,N_372);
and U6277 (N_6277,N_1758,N_1399);
or U6278 (N_6278,N_3837,N_3582);
xor U6279 (N_6279,N_1496,N_4730);
xor U6280 (N_6280,N_3887,N_1242);
xor U6281 (N_6281,N_761,N_1198);
nand U6282 (N_6282,N_492,N_3519);
or U6283 (N_6283,N_3009,N_3254);
xor U6284 (N_6284,N_4716,N_1184);
and U6285 (N_6285,N_2284,N_62);
nor U6286 (N_6286,N_3518,N_2424);
xor U6287 (N_6287,N_4259,N_1836);
and U6288 (N_6288,N_3551,N_293);
nor U6289 (N_6289,N_68,N_1632);
nor U6290 (N_6290,N_3748,N_2074);
and U6291 (N_6291,N_4980,N_1264);
nor U6292 (N_6292,N_3510,N_4353);
and U6293 (N_6293,N_1456,N_2826);
xor U6294 (N_6294,N_1172,N_4824);
or U6295 (N_6295,N_965,N_653);
xnor U6296 (N_6296,N_1513,N_855);
nor U6297 (N_6297,N_894,N_1493);
or U6298 (N_6298,N_1803,N_4815);
xnor U6299 (N_6299,N_9,N_2433);
or U6300 (N_6300,N_706,N_3646);
or U6301 (N_6301,N_4356,N_153);
or U6302 (N_6302,N_391,N_777);
nand U6303 (N_6303,N_3733,N_3747);
or U6304 (N_6304,N_888,N_505);
and U6305 (N_6305,N_2355,N_3526);
nand U6306 (N_6306,N_4679,N_1017);
nor U6307 (N_6307,N_3707,N_3682);
nand U6308 (N_6308,N_921,N_2986);
or U6309 (N_6309,N_2143,N_4618);
nand U6310 (N_6310,N_4811,N_4431);
xnor U6311 (N_6311,N_157,N_3874);
nor U6312 (N_6312,N_181,N_3952);
or U6313 (N_6313,N_1975,N_3788);
nor U6314 (N_6314,N_4972,N_1249);
nor U6315 (N_6315,N_405,N_3447);
xor U6316 (N_6316,N_2151,N_4386);
xnor U6317 (N_6317,N_367,N_4505);
or U6318 (N_6318,N_1336,N_1412);
nand U6319 (N_6319,N_4172,N_1570);
nand U6320 (N_6320,N_1348,N_4992);
and U6321 (N_6321,N_2114,N_3856);
nor U6322 (N_6322,N_1875,N_606);
nor U6323 (N_6323,N_3512,N_4402);
and U6324 (N_6324,N_1442,N_152);
or U6325 (N_6325,N_3269,N_300);
nand U6326 (N_6326,N_2829,N_1529);
nor U6327 (N_6327,N_409,N_2913);
and U6328 (N_6328,N_3202,N_1196);
or U6329 (N_6329,N_4007,N_3732);
xnor U6330 (N_6330,N_3913,N_2184);
xnor U6331 (N_6331,N_1157,N_3660);
or U6332 (N_6332,N_3428,N_3500);
or U6333 (N_6333,N_1817,N_4780);
xor U6334 (N_6334,N_119,N_70);
and U6335 (N_6335,N_895,N_2956);
nand U6336 (N_6336,N_3684,N_847);
nor U6337 (N_6337,N_3488,N_1339);
xor U6338 (N_6338,N_1317,N_1552);
nor U6339 (N_6339,N_4686,N_1753);
xnor U6340 (N_6340,N_97,N_2505);
xor U6341 (N_6341,N_917,N_3294);
nor U6342 (N_6342,N_1047,N_4485);
or U6343 (N_6343,N_494,N_2180);
nand U6344 (N_6344,N_1785,N_2095);
xnor U6345 (N_6345,N_510,N_4637);
and U6346 (N_6346,N_228,N_3104);
nor U6347 (N_6347,N_4209,N_1948);
xor U6348 (N_6348,N_4868,N_3667);
or U6349 (N_6349,N_3449,N_4571);
nand U6350 (N_6350,N_3032,N_3895);
or U6351 (N_6351,N_1492,N_3916);
nand U6352 (N_6352,N_4190,N_2888);
and U6353 (N_6353,N_1666,N_3636);
nor U6354 (N_6354,N_3349,N_1024);
and U6355 (N_6355,N_1590,N_166);
and U6356 (N_6356,N_2305,N_2157);
or U6357 (N_6357,N_4210,N_530);
and U6358 (N_6358,N_3482,N_3986);
nor U6359 (N_6359,N_2221,N_4065);
nor U6360 (N_6360,N_4580,N_4551);
xnor U6361 (N_6361,N_1797,N_1450);
xnor U6362 (N_6362,N_1626,N_3093);
nor U6363 (N_6363,N_4548,N_2511);
and U6364 (N_6364,N_3448,N_4642);
nand U6365 (N_6365,N_4643,N_1402);
nand U6366 (N_6366,N_48,N_4914);
xnor U6367 (N_6367,N_2334,N_4365);
nor U6368 (N_6368,N_3800,N_2356);
and U6369 (N_6369,N_3179,N_2158);
nand U6370 (N_6370,N_624,N_1538);
nand U6371 (N_6371,N_1614,N_805);
and U6372 (N_6372,N_3656,N_4991);
or U6373 (N_6373,N_4460,N_1108);
xor U6374 (N_6374,N_4999,N_171);
nand U6375 (N_6375,N_4660,N_3768);
xor U6376 (N_6376,N_90,N_3089);
nand U6377 (N_6377,N_2498,N_1841);
nand U6378 (N_6378,N_674,N_375);
or U6379 (N_6379,N_4250,N_131);
nor U6380 (N_6380,N_3716,N_466);
and U6381 (N_6381,N_2190,N_4092);
and U6382 (N_6382,N_3322,N_2609);
nand U6383 (N_6383,N_2078,N_1078);
nand U6384 (N_6384,N_1088,N_4116);
nand U6385 (N_6385,N_3424,N_1387);
nor U6386 (N_6386,N_3237,N_155);
xnor U6387 (N_6387,N_517,N_2105);
nand U6388 (N_6388,N_1756,N_2206);
nor U6389 (N_6389,N_2065,N_4064);
nor U6390 (N_6390,N_295,N_2538);
or U6391 (N_6391,N_3122,N_3421);
nand U6392 (N_6392,N_2572,N_4662);
nor U6393 (N_6393,N_1475,N_4276);
and U6394 (N_6394,N_1994,N_1828);
nor U6395 (N_6395,N_144,N_3107);
nand U6396 (N_6396,N_1507,N_3271);
or U6397 (N_6397,N_17,N_3692);
and U6398 (N_6398,N_139,N_1125);
or U6399 (N_6399,N_593,N_2808);
and U6400 (N_6400,N_2895,N_1272);
and U6401 (N_6401,N_19,N_4450);
and U6402 (N_6402,N_1667,N_52);
nand U6403 (N_6403,N_3609,N_2480);
nand U6404 (N_6404,N_1101,N_2544);
nand U6405 (N_6405,N_2530,N_1757);
and U6406 (N_6406,N_3528,N_1851);
xor U6407 (N_6407,N_1386,N_2287);
or U6408 (N_6408,N_271,N_1749);
xnor U6409 (N_6409,N_3281,N_2069);
and U6410 (N_6410,N_2385,N_3661);
and U6411 (N_6411,N_1194,N_1138);
and U6412 (N_6412,N_2909,N_4603);
nand U6413 (N_6413,N_173,N_4920);
nand U6414 (N_6414,N_931,N_590);
nand U6415 (N_6415,N_4907,N_3734);
or U6416 (N_6416,N_4264,N_4771);
nand U6417 (N_6417,N_306,N_1774);
nor U6418 (N_6418,N_1119,N_4927);
and U6419 (N_6419,N_3140,N_4963);
nor U6420 (N_6420,N_2485,N_3848);
xor U6421 (N_6421,N_4545,N_2354);
xnor U6422 (N_6422,N_806,N_4202);
nand U6423 (N_6423,N_429,N_2204);
and U6424 (N_6424,N_2125,N_1941);
nand U6425 (N_6425,N_2404,N_4468);
and U6426 (N_6426,N_642,N_3431);
or U6427 (N_6427,N_1266,N_1476);
nor U6428 (N_6428,N_4761,N_1379);
or U6429 (N_6429,N_2937,N_1983);
nor U6430 (N_6430,N_2081,N_1792);
nor U6431 (N_6431,N_4825,N_4222);
and U6432 (N_6432,N_1318,N_4124);
nand U6433 (N_6433,N_4419,N_2102);
nor U6434 (N_6434,N_4533,N_3941);
and U6435 (N_6435,N_4330,N_4703);
nor U6436 (N_6436,N_3753,N_2152);
nand U6437 (N_6437,N_2801,N_4669);
nand U6438 (N_6438,N_4737,N_1578);
and U6439 (N_6439,N_4452,N_967);
nor U6440 (N_6440,N_334,N_3043);
xnor U6441 (N_6441,N_3626,N_3151);
xor U6442 (N_6442,N_2517,N_4744);
and U6443 (N_6443,N_4510,N_1285);
or U6444 (N_6444,N_2016,N_569);
or U6445 (N_6445,N_3960,N_2753);
xor U6446 (N_6446,N_2697,N_1060);
nor U6447 (N_6447,N_2207,N_3310);
nor U6448 (N_6448,N_3347,N_4376);
xnor U6449 (N_6449,N_4535,N_3405);
nor U6450 (N_6450,N_804,N_1012);
or U6451 (N_6451,N_1497,N_707);
nand U6452 (N_6452,N_2616,N_3169);
and U6453 (N_6453,N_710,N_4267);
xnor U6454 (N_6454,N_3427,N_532);
and U6455 (N_6455,N_1168,N_4194);
xor U6456 (N_6456,N_4985,N_1676);
nand U6457 (N_6457,N_1139,N_3341);
and U6458 (N_6458,N_4649,N_2185);
nor U6459 (N_6459,N_3628,N_534);
xnor U6460 (N_6460,N_3611,N_2403);
or U6461 (N_6461,N_1966,N_493);
and U6462 (N_6462,N_1164,N_4257);
or U6463 (N_6463,N_1413,N_1770);
nor U6464 (N_6464,N_1656,N_3771);
or U6465 (N_6465,N_2982,N_3301);
nor U6466 (N_6466,N_3260,N_1816);
xnor U6467 (N_6467,N_2161,N_1064);
or U6468 (N_6468,N_488,N_1743);
or U6469 (N_6469,N_3548,N_261);
nor U6470 (N_6470,N_2597,N_1636);
or U6471 (N_6471,N_1704,N_4025);
or U6472 (N_6472,N_3285,N_2482);
or U6473 (N_6473,N_3064,N_2320);
nor U6474 (N_6474,N_1918,N_3802);
nor U6475 (N_6475,N_4042,N_4467);
or U6476 (N_6476,N_297,N_2943);
nand U6477 (N_6477,N_3370,N_3279);
nand U6478 (N_6478,N_2983,N_911);
nor U6479 (N_6479,N_4125,N_1333);
nor U6480 (N_6480,N_2765,N_4117);
and U6481 (N_6481,N_4954,N_4428);
nand U6482 (N_6482,N_3498,N_4201);
nand U6483 (N_6483,N_86,N_839);
nand U6484 (N_6484,N_4861,N_2623);
nor U6485 (N_6485,N_2827,N_3516);
and U6486 (N_6486,N_2412,N_4550);
xor U6487 (N_6487,N_4036,N_178);
xor U6488 (N_6488,N_174,N_3774);
and U6489 (N_6489,N_3622,N_2194);
and U6490 (N_6490,N_1245,N_563);
xor U6491 (N_6491,N_3894,N_2101);
nor U6492 (N_6492,N_4589,N_2512);
nor U6493 (N_6493,N_2774,N_4738);
nand U6494 (N_6494,N_1344,N_663);
or U6495 (N_6495,N_1204,N_4687);
nor U6496 (N_6496,N_373,N_1358);
nand U6497 (N_6497,N_4346,N_4410);
and U6498 (N_6498,N_3205,N_3537);
or U6499 (N_6499,N_3725,N_1796);
nor U6500 (N_6500,N_1199,N_732);
nor U6501 (N_6501,N_3403,N_4320);
xnor U6502 (N_6502,N_2621,N_2853);
and U6503 (N_6503,N_3136,N_2906);
or U6504 (N_6504,N_2011,N_3539);
xor U6505 (N_6505,N_781,N_3019);
and U6506 (N_6506,N_4486,N_2793);
or U6507 (N_6507,N_980,N_1409);
or U6508 (N_6508,N_3850,N_2012);
nor U6509 (N_6509,N_2432,N_143);
nand U6510 (N_6510,N_1508,N_1392);
nand U6511 (N_6511,N_2912,N_3227);
nor U6512 (N_6512,N_632,N_3154);
nand U6513 (N_6513,N_4284,N_4256);
and U6514 (N_6514,N_2873,N_3097);
and U6515 (N_6515,N_3371,N_326);
nor U6516 (N_6516,N_1814,N_2897);
nand U6517 (N_6517,N_4182,N_3407);
or U6518 (N_6518,N_1149,N_2579);
nor U6519 (N_6519,N_3198,N_2575);
and U6520 (N_6520,N_3546,N_4061);
xor U6521 (N_6521,N_4375,N_4928);
and U6522 (N_6522,N_1669,N_3697);
and U6523 (N_6523,N_2939,N_3736);
and U6524 (N_6524,N_4968,N_4611);
nand U6525 (N_6525,N_539,N_384);
nor U6526 (N_6526,N_3652,N_1914);
xnor U6527 (N_6527,N_1710,N_4528);
or U6528 (N_6528,N_4223,N_2627);
nor U6529 (N_6529,N_638,N_3348);
or U6530 (N_6530,N_1441,N_4271);
nor U6531 (N_6531,N_1837,N_2336);
or U6532 (N_6532,N_4371,N_1868);
or U6533 (N_6533,N_3781,N_2250);
and U6534 (N_6534,N_4663,N_3452);
and U6535 (N_6535,N_725,N_3268);
xor U6536 (N_6536,N_3765,N_2014);
nor U6537 (N_6537,N_4343,N_946);
xnor U6538 (N_6538,N_2668,N_3414);
nor U6539 (N_6539,N_365,N_2030);
and U6540 (N_6540,N_2705,N_4388);
nand U6541 (N_6541,N_2450,N_3638);
nor U6542 (N_6542,N_3862,N_4720);
xnor U6543 (N_6543,N_285,N_2972);
or U6544 (N_6544,N_3326,N_4599);
nand U6545 (N_6545,N_369,N_4507);
xnor U6546 (N_6546,N_2749,N_1197);
or U6547 (N_6547,N_2883,N_3791);
and U6548 (N_6548,N_3503,N_2645);
xor U6549 (N_6549,N_4106,N_230);
xor U6550 (N_6550,N_3877,N_2171);
or U6551 (N_6551,N_3307,N_1869);
xnor U6552 (N_6552,N_2587,N_827);
nor U6553 (N_6553,N_3817,N_1604);
nand U6554 (N_6554,N_2241,N_2359);
nor U6555 (N_6555,N_1911,N_3700);
nand U6556 (N_6556,N_1155,N_1873);
nand U6557 (N_6557,N_3335,N_3216);
xor U6558 (N_6558,N_453,N_2701);
or U6559 (N_6559,N_4254,N_538);
xnor U6560 (N_6560,N_4009,N_4585);
and U6561 (N_6561,N_2174,N_3599);
and U6562 (N_6562,N_2591,N_4715);
and U6563 (N_6563,N_782,N_3124);
nand U6564 (N_6564,N_3422,N_3331);
xor U6565 (N_6565,N_2286,N_2440);
nand U6566 (N_6566,N_961,N_4956);
nor U6567 (N_6567,N_2896,N_4443);
xor U6568 (N_6568,N_3031,N_3321);
or U6569 (N_6569,N_1089,N_39);
nor U6570 (N_6570,N_1302,N_3982);
or U6571 (N_6571,N_2112,N_130);
xnor U6572 (N_6572,N_4180,N_194);
xnor U6573 (N_6573,N_1015,N_3416);
and U6574 (N_6574,N_728,N_4672);
nor U6575 (N_6575,N_2742,N_4884);
nor U6576 (N_6576,N_2818,N_1364);
xnor U6577 (N_6577,N_2209,N_1331);
or U6578 (N_6578,N_4446,N_2582);
nand U6579 (N_6579,N_621,N_1445);
xor U6580 (N_6580,N_1571,N_704);
xor U6581 (N_6581,N_4553,N_825);
xnor U6582 (N_6582,N_2908,N_2107);
xnor U6583 (N_6583,N_3880,N_2969);
nand U6584 (N_6584,N_3679,N_2526);
nor U6585 (N_6585,N_615,N_3318);
and U6586 (N_6586,N_1233,N_1784);
xor U6587 (N_6587,N_1295,N_4325);
nor U6588 (N_6588,N_906,N_2260);
and U6589 (N_6589,N_3437,N_2658);
and U6590 (N_6590,N_923,N_4750);
or U6591 (N_6591,N_509,N_4949);
nand U6592 (N_6592,N_2222,N_249);
nand U6593 (N_6593,N_3388,N_1754);
and U6594 (N_6594,N_3066,N_2092);
or U6595 (N_6595,N_4911,N_885);
nand U6596 (N_6596,N_3186,N_2923);
or U6597 (N_6597,N_1885,N_3717);
nand U6598 (N_6598,N_4898,N_4683);
nor U6599 (N_6599,N_3280,N_2662);
or U6600 (N_6600,N_4760,N_3221);
xnor U6601 (N_6601,N_843,N_3226);
xor U6602 (N_6602,N_4747,N_324);
and U6603 (N_6603,N_4893,N_597);
or U6604 (N_6604,N_518,N_3617);
and U6605 (N_6605,N_1222,N_3613);
and U6606 (N_6606,N_4766,N_2915);
and U6607 (N_6607,N_3825,N_3234);
and U6608 (N_6608,N_1686,N_2593);
nand U6609 (N_6609,N_1771,N_1371);
nand U6610 (N_6610,N_2295,N_3337);
and U6611 (N_6611,N_1967,N_2068);
and U6612 (N_6612,N_1505,N_974);
and U6613 (N_6613,N_1820,N_47);
xor U6614 (N_6614,N_4849,N_4878);
nor U6615 (N_6615,N_2590,N_2104);
and U6616 (N_6616,N_1894,N_2472);
xnor U6617 (N_6617,N_4038,N_900);
or U6618 (N_6618,N_1616,N_3706);
xnor U6619 (N_6619,N_3799,N_963);
nand U6620 (N_6620,N_2689,N_2766);
or U6621 (N_6621,N_1896,N_1989);
xor U6622 (N_6622,N_975,N_3486);
or U6623 (N_6623,N_323,N_4602);
nand U6624 (N_6624,N_3088,N_2247);
nand U6625 (N_6625,N_4733,N_4342);
xnor U6626 (N_6626,N_4735,N_4301);
and U6627 (N_6627,N_49,N_1712);
nor U6628 (N_6628,N_762,N_3563);
xor U6629 (N_6629,N_1112,N_3100);
nor U6630 (N_6630,N_3400,N_3598);
xnor U6631 (N_6631,N_3451,N_736);
or U6632 (N_6632,N_132,N_1280);
or U6633 (N_6633,N_1239,N_2179);
nand U6634 (N_6634,N_4598,N_4263);
nor U6635 (N_6635,N_1812,N_2809);
nor U6636 (N_6636,N_3156,N_2537);
nor U6637 (N_6637,N_3820,N_3423);
and U6638 (N_6638,N_2479,N_4199);
or U6639 (N_6639,N_2353,N_2145);
or U6640 (N_6640,N_4609,N_2767);
xor U6641 (N_6641,N_4832,N_32);
xor U6642 (N_6642,N_2379,N_3068);
nor U6643 (N_6643,N_1325,N_1718);
or U6644 (N_6644,N_53,N_2586);
nor U6645 (N_6645,N_1569,N_1129);
nand U6646 (N_6646,N_22,N_2798);
nand U6647 (N_6647,N_785,N_1879);
or U6648 (N_6648,N_2807,N_3814);
or U6649 (N_6649,N_3443,N_4152);
or U6650 (N_6650,N_3884,N_1449);
nor U6651 (N_6651,N_2096,N_1857);
nor U6652 (N_6652,N_2243,N_1220);
nand U6653 (N_6653,N_3792,N_2040);
nand U6654 (N_6654,N_4987,N_357);
xnor U6655 (N_6655,N_575,N_4794);
or U6656 (N_6656,N_2553,N_419);
nand U6657 (N_6657,N_3253,N_2173);
nand U6658 (N_6658,N_858,N_4979);
nand U6659 (N_6659,N_3749,N_671);
and U6660 (N_6660,N_3323,N_3476);
xor U6661 (N_6661,N_3520,N_790);
nor U6662 (N_6662,N_1473,N_3214);
or U6663 (N_6663,N_3418,N_254);
xnor U6664 (N_6664,N_3233,N_613);
nor U6665 (N_6665,N_3489,N_3103);
xor U6666 (N_6666,N_3199,N_4881);
xnor U6667 (N_6667,N_3918,N_936);
and U6668 (N_6668,N_3907,N_3243);
nor U6669 (N_6669,N_4682,N_133);
nor U6670 (N_6670,N_1081,N_1469);
nand U6671 (N_6671,N_3203,N_3383);
or U6672 (N_6672,N_3603,N_4033);
or U6673 (N_6673,N_4361,N_457);
xor U6674 (N_6674,N_3082,N_1321);
nor U6675 (N_6675,N_3295,N_4081);
xor U6676 (N_6676,N_2921,N_4995);
nor U6677 (N_6677,N_4434,N_3556);
or U6678 (N_6678,N_2274,N_2601);
and U6679 (N_6679,N_1210,N_1018);
and U6680 (N_6680,N_2170,N_2603);
and U6681 (N_6681,N_2444,N_2996);
or U6682 (N_6682,N_13,N_3604);
nand U6683 (N_6683,N_4054,N_2149);
or U6684 (N_6684,N_66,N_3593);
xor U6685 (N_6685,N_878,N_614);
nand U6686 (N_6686,N_3101,N_3685);
nand U6687 (N_6687,N_217,N_2275);
xor U6688 (N_6688,N_982,N_4539);
nor U6689 (N_6689,N_1631,N_2322);
and U6690 (N_6690,N_1105,N_4285);
nor U6691 (N_6691,N_1013,N_1085);
nand U6692 (N_6692,N_4014,N_268);
nand U6693 (N_6693,N_4023,N_4783);
xnor U6694 (N_6694,N_631,N_3639);
and U6695 (N_6695,N_3683,N_1165);
xor U6696 (N_6696,N_3726,N_845);
xnor U6697 (N_6697,N_3589,N_3673);
and U6698 (N_6698,N_4401,N_2903);
and U6699 (N_6699,N_1040,N_1764);
xnor U6700 (N_6700,N_1881,N_1042);
and U6701 (N_6701,N_3807,N_1916);
nor U6702 (N_6702,N_3798,N_4165);
xor U6703 (N_6703,N_4090,N_3738);
and U6704 (N_6704,N_2552,N_2925);
xnor U6705 (N_6705,N_2422,N_1755);
or U6706 (N_6706,N_250,N_2786);
nand U6707 (N_6707,N_1345,N_4767);
xnor U6708 (N_6708,N_1484,N_1596);
nor U6709 (N_6709,N_350,N_2489);
or U6710 (N_6710,N_4319,N_255);
xor U6711 (N_6711,N_484,N_127);
and U6712 (N_6712,N_4666,N_2887);
or U6713 (N_6713,N_3657,N_2846);
and U6714 (N_6714,N_4797,N_2417);
or U6715 (N_6715,N_1154,N_2291);
nor U6716 (N_6716,N_4110,N_2342);
nand U6717 (N_6717,N_656,N_4447);
nor U6718 (N_6718,N_3020,N_55);
and U6719 (N_6719,N_4445,N_1185);
nor U6720 (N_6720,N_749,N_441);
nor U6721 (N_6721,N_1783,N_924);
xor U6722 (N_6722,N_1706,N_1368);
nand U6723 (N_6723,N_1909,N_4821);
nor U6724 (N_6724,N_2910,N_4623);
and U6725 (N_6725,N_1883,N_971);
nor U6726 (N_6726,N_3826,N_1396);
xnor U6727 (N_6727,N_1832,N_2976);
xor U6728 (N_6728,N_3654,N_1093);
and U6729 (N_6729,N_1551,N_3530);
or U6730 (N_6730,N_908,N_4332);
nand U6731 (N_6731,N_3181,N_3815);
xnor U6732 (N_6732,N_2848,N_665);
nor U6733 (N_6733,N_2395,N_238);
xor U6734 (N_6734,N_3778,N_4998);
or U6735 (N_6735,N_4961,N_4994);
nand U6736 (N_6736,N_3742,N_2532);
or U6737 (N_6737,N_1734,N_3481);
xnor U6738 (N_6738,N_4515,N_2941);
nand U6739 (N_6739,N_3944,N_1542);
and U6740 (N_6740,N_3760,N_1000);
and U6741 (N_6741,N_185,N_4083);
xor U6742 (N_6742,N_1071,N_191);
and U6743 (N_6743,N_560,N_4894);
or U6744 (N_6744,N_3608,N_2460);
nand U6745 (N_6745,N_3074,N_4156);
nand U6746 (N_6746,N_123,N_4684);
or U6747 (N_6747,N_4626,N_3910);
and U6748 (N_6748,N_2058,N_3461);
nor U6749 (N_6749,N_1426,N_3651);
and U6750 (N_6750,N_823,N_1742);
and U6751 (N_6751,N_1878,N_541);
nand U6752 (N_6752,N_1259,N_1267);
and U6753 (N_6753,N_12,N_999);
xor U6754 (N_6754,N_4517,N_1483);
or U6755 (N_6755,N_4782,N_2926);
xor U6756 (N_6756,N_4690,N_3379);
or U6757 (N_6757,N_3822,N_2369);
nand U6758 (N_6758,N_2246,N_3436);
or U6759 (N_6759,N_3577,N_1471);
xor U6760 (N_6760,N_3258,N_522);
or U6761 (N_6761,N_4828,N_2581);
or U6762 (N_6762,N_2374,N_4634);
and U6763 (N_6763,N_1752,N_321);
xnor U6764 (N_6764,N_2931,N_703);
nand U6765 (N_6765,N_1096,N_3062);
and U6766 (N_6766,N_3550,N_830);
or U6767 (N_6767,N_4883,N_2740);
or U6768 (N_6768,N_1990,N_4444);
xnor U6769 (N_6769,N_2594,N_1372);
xnor U6770 (N_6770,N_1126,N_1627);
nand U6771 (N_6771,N_103,N_600);
nor U6772 (N_6772,N_4710,N_4842);
nand U6773 (N_6773,N_2599,N_1699);
or U6774 (N_6774,N_2133,N_3515);
or U6775 (N_6775,N_2383,N_2483);
and U6776 (N_6776,N_4807,N_836);
nand U6777 (N_6777,N_1621,N_1182);
or U6778 (N_6778,N_428,N_2573);
and U6779 (N_6779,N_1790,N_2306);
and U6780 (N_6780,N_3868,N_1486);
or U6781 (N_6781,N_1642,N_4790);
nand U6782 (N_6782,N_2524,N_3141);
or U6783 (N_6783,N_3838,N_4093);
nand U6784 (N_6784,N_2577,N_4698);
nor U6785 (N_6785,N_2191,N_2539);
nand U6786 (N_6786,N_4068,N_2666);
or U6787 (N_6787,N_1781,N_4457);
or U6788 (N_6788,N_2261,N_1504);
or U6789 (N_6789,N_3457,N_1397);
or U6790 (N_6790,N_1334,N_821);
nand U6791 (N_6791,N_2047,N_1684);
or U6792 (N_6792,N_4670,N_4086);
nor U6793 (N_6793,N_34,N_996);
nor U6794 (N_6794,N_1871,N_2632);
nand U6795 (N_6795,N_2459,N_4587);
nor U6796 (N_6796,N_61,N_1968);
or U6797 (N_6797,N_2670,N_4758);
and U6798 (N_6798,N_1167,N_4229);
nor U6799 (N_6799,N_659,N_3360);
or U6800 (N_6800,N_3035,N_1691);
xnor U6801 (N_6801,N_4567,N_328);
or U6802 (N_6802,N_796,N_1953);
nor U6803 (N_6803,N_4946,N_3458);
xnor U6804 (N_6804,N_3718,N_1949);
xor U6805 (N_6805,N_1951,N_4212);
nand U6806 (N_6806,N_2797,N_2781);
nand U6807 (N_6807,N_1772,N_683);
xor U6808 (N_6808,N_1908,N_1183);
xnor U6809 (N_6809,N_1730,N_1111);
nor U6810 (N_6810,N_2860,N_4975);
and U6811 (N_6811,N_2397,N_4311);
and U6812 (N_6812,N_4029,N_1463);
nor U6813 (N_6813,N_739,N_4085);
nor U6814 (N_6814,N_4429,N_727);
and U6815 (N_6815,N_697,N_2439);
or U6816 (N_6816,N_135,N_1213);
nand U6817 (N_6817,N_1703,N_1104);
xnor U6818 (N_6818,N_401,N_1892);
nor U6819 (N_6819,N_4318,N_57);
or U6820 (N_6820,N_3223,N_1502);
xnor U6821 (N_6821,N_4846,N_2534);
xor U6822 (N_6822,N_4942,N_156);
xor U6823 (N_6823,N_394,N_771);
xor U6824 (N_6824,N_3222,N_2029);
nor U6825 (N_6825,N_922,N_3225);
xnor U6826 (N_6826,N_1490,N_3175);
xor U6827 (N_6827,N_1685,N_4000);
and U6828 (N_6828,N_2868,N_2292);
xnor U6829 (N_6829,N_1664,N_4595);
nor U6830 (N_6830,N_1384,N_4919);
and U6831 (N_6831,N_820,N_1842);
nand U6832 (N_6832,N_3312,N_4977);
xor U6833 (N_6833,N_4417,N_50);
and U6834 (N_6834,N_1944,N_3446);
xor U6835 (N_6835,N_4597,N_1452);
xor U6836 (N_6836,N_2698,N_2197);
xnor U6837 (N_6837,N_1224,N_2613);
nor U6838 (N_6838,N_1924,N_801);
and U6839 (N_6839,N_1829,N_1361);
or U6840 (N_6840,N_4016,N_2596);
or U6841 (N_6841,N_1116,N_672);
nand U6842 (N_6842,N_3843,N_702);
xnor U6843 (N_6843,N_1906,N_3311);
and U6844 (N_6844,N_998,N_2644);
xor U6845 (N_6845,N_2556,N_4749);
and U6846 (N_6846,N_3187,N_3255);
or U6847 (N_6847,N_1287,N_2954);
or U6848 (N_6848,N_3277,N_4372);
xor U6849 (N_6849,N_2484,N_1575);
or U6850 (N_6850,N_3602,N_4207);
or U6851 (N_6851,N_4863,N_4877);
and U6852 (N_6852,N_4523,N_4547);
or U6853 (N_6853,N_4227,N_4578);
nand U6854 (N_6854,N_3183,N_4228);
or U6855 (N_6855,N_2132,N_3612);
or U6856 (N_6856,N_3655,N_4440);
nor U6857 (N_6857,N_3670,N_857);
xnor U6858 (N_6858,N_3964,N_2400);
xor U6859 (N_6859,N_3356,N_1876);
and U6860 (N_6860,N_1628,N_4502);
or U6861 (N_6861,N_1727,N_854);
nand U6862 (N_6862,N_4364,N_1524);
nor U6863 (N_6863,N_2510,N_1558);
or U6864 (N_6864,N_2840,N_966);
nand U6865 (N_6865,N_3413,N_2727);
xor U6866 (N_6866,N_2213,N_2420);
or U6867 (N_6867,N_1860,N_1092);
or U6868 (N_6868,N_1688,N_3389);
and U6869 (N_6869,N_4981,N_4466);
nand U6870 (N_6870,N_3633,N_866);
nor U6871 (N_6871,N_4203,N_3705);
xnor U6872 (N_6872,N_4753,N_1306);
nor U6873 (N_6873,N_608,N_2871);
nor U6874 (N_6874,N_4381,N_4010);
nor U6875 (N_6875,N_2734,N_1539);
and U6876 (N_6876,N_4066,N_36);
nand U6877 (N_6877,N_1825,N_4493);
or U6878 (N_6878,N_633,N_1567);
nor U6879 (N_6879,N_3219,N_4020);
xnor U6880 (N_6880,N_3430,N_1142);
and U6881 (N_6881,N_1782,N_2235);
nor U6882 (N_6882,N_3573,N_3737);
and U6883 (N_6883,N_3909,N_3981);
xnor U6884 (N_6884,N_2073,N_1179);
or U6885 (N_6885,N_3475,N_4495);
nand U6886 (N_6886,N_4300,N_2037);
and U6887 (N_6887,N_340,N_4237);
or U6888 (N_6888,N_311,N_1809);
nand U6889 (N_6889,N_3936,N_741);
or U6890 (N_6890,N_1644,N_604);
nand U6891 (N_6891,N_4072,N_2210);
nand U6892 (N_6892,N_3993,N_1933);
and U6893 (N_6893,N_3375,N_318);
nand U6894 (N_6894,N_848,N_197);
xor U6895 (N_6895,N_595,N_120);
nand U6896 (N_6896,N_4012,N_1090);
and U6897 (N_6897,N_2501,N_1359);
xor U6898 (N_6898,N_2351,N_1888);
nand U6899 (N_6899,N_2402,N_2584);
nand U6900 (N_6900,N_698,N_1932);
nor U6901 (N_6901,N_2543,N_3833);
nor U6902 (N_6902,N_399,N_3474);
and U6903 (N_6903,N_2463,N_1340);
or U6904 (N_6904,N_4947,N_2535);
or U6905 (N_6905,N_1923,N_3201);
nand U6906 (N_6906,N_602,N_2646);
or U6907 (N_6907,N_3147,N_2894);
nand U6908 (N_6908,N_3663,N_4899);
xnor U6909 (N_6909,N_4119,N_1);
nand U6910 (N_6910,N_4317,N_1058);
xor U6911 (N_6911,N_2707,N_3722);
and U6912 (N_6912,N_3999,N_3305);
or U6913 (N_6913,N_2251,N_2735);
and U6914 (N_6914,N_601,N_1485);
or U6915 (N_6915,N_489,N_4101);
and U6916 (N_6916,N_3640,N_1747);
and U6917 (N_6917,N_1929,N_4270);
or U6918 (N_6918,N_3466,N_2942);
or U6919 (N_6919,N_1046,N_3809);
and U6920 (N_6920,N_3317,N_1133);
or U6921 (N_6921,N_2702,N_2967);
or U6922 (N_6922,N_4834,N_525);
and U6923 (N_6923,N_565,N_2453);
nor U6924 (N_6924,N_4052,N_3292);
or U6925 (N_6925,N_958,N_2495);
nand U6926 (N_6926,N_842,N_690);
nor U6927 (N_6927,N_3309,N_3890);
nor U6928 (N_6928,N_3605,N_2930);
or U6929 (N_6929,N_1311,N_4407);
nor U6930 (N_6930,N_1849,N_4046);
xor U6931 (N_6931,N_4809,N_589);
and U6932 (N_6932,N_2471,N_3678);
nand U6933 (N_6933,N_3619,N_1113);
or U6934 (N_6934,N_3762,N_1549);
nor U6935 (N_6935,N_294,N_1886);
nor U6936 (N_6936,N_2741,N_3669);
xnor U6937 (N_6937,N_3127,N_3631);
nand U6938 (N_6938,N_3674,N_2164);
nand U6939 (N_6939,N_1403,N_1235);
xor U6940 (N_6940,N_2626,N_1723);
nor U6941 (N_6941,N_2435,N_3587);
or U6942 (N_6942,N_121,N_910);
nor U6943 (N_6943,N_1893,N_687);
nand U6944 (N_6944,N_4504,N_3264);
nand U6945 (N_6945,N_235,N_4882);
nor U6946 (N_6946,N_582,N_1324);
nor U6947 (N_6947,N_579,N_1759);
xnor U6948 (N_6948,N_4420,N_3508);
or U6949 (N_6949,N_1866,N_622);
and U6950 (N_6950,N_2036,N_2309);
xnor U6951 (N_6951,N_2364,N_1395);
and U6952 (N_6952,N_3343,N_1158);
nand U6953 (N_6953,N_3290,N_4986);
or U6954 (N_6954,N_1608,N_1545);
xnor U6955 (N_6955,N_4279,N_4615);
xnor U6956 (N_6956,N_628,N_2863);
nor U6957 (N_6957,N_508,N_2297);
or U6958 (N_6958,N_3232,N_2547);
xnor U6959 (N_6959,N_3299,N_1208);
nor U6960 (N_6960,N_266,N_3018);
xnor U6961 (N_6961,N_512,N_2034);
nand U6962 (N_6962,N_629,N_925);
nor U6963 (N_6963,N_2227,N_4339);
nor U6964 (N_6964,N_2088,N_3648);
nor U6965 (N_6965,N_1193,N_4149);
and U6966 (N_6966,N_2299,N_889);
and U6967 (N_6967,N_1972,N_3439);
and U6968 (N_6968,N_3420,N_3565);
or U6969 (N_6969,N_1219,N_344);
nor U6970 (N_6970,N_3480,N_175);
or U6971 (N_6971,N_2126,N_3236);
nand U6972 (N_6972,N_918,N_2414);
nor U6973 (N_6973,N_4524,N_3642);
or U6974 (N_6974,N_4591,N_3247);
nor U6975 (N_6975,N_2832,N_1897);
nor U6976 (N_6976,N_2576,N_567);
or U6977 (N_6977,N_1055,N_1572);
nor U6978 (N_6978,N_1282,N_2876);
nor U6979 (N_6979,N_4926,N_426);
and U6980 (N_6980,N_4870,N_3256);
nor U6981 (N_6981,N_1377,N_3625);
nand U6982 (N_6982,N_3138,N_3470);
and U6983 (N_6983,N_3041,N_4711);
nor U6984 (N_6984,N_896,N_3072);
nor U6985 (N_6985,N_1404,N_1585);
xor U6986 (N_6986,N_106,N_4051);
xnor U6987 (N_6987,N_3777,N_1610);
nor U6988 (N_6988,N_2611,N_4740);
nor U6989 (N_6989,N_3963,N_1726);
xnor U6990 (N_6990,N_1541,N_4812);
xor U6991 (N_6991,N_4696,N_948);
or U6992 (N_6992,N_829,N_873);
nor U6993 (N_6993,N_754,N_23);
nand U6994 (N_6994,N_3380,N_1981);
nor U6995 (N_6995,N_2192,N_1835);
and U6996 (N_6996,N_4170,N_4788);
xor U6997 (N_6997,N_654,N_2660);
nor U6998 (N_6998,N_1308,N_2932);
and U6999 (N_6999,N_2302,N_2052);
or U7000 (N_7000,N_3274,N_3300);
nand U7001 (N_7001,N_995,N_1228);
nand U7002 (N_7002,N_1535,N_10);
and U7003 (N_7003,N_695,N_2667);
nand U7004 (N_7004,N_2736,N_3073);
nand U7005 (N_7005,N_264,N_556);
xor U7006 (N_7006,N_3959,N_574);
xor U7007 (N_7007,N_760,N_4435);
nor U7008 (N_7008,N_341,N_2847);
nand U7009 (N_7009,N_1910,N_1861);
nor U7010 (N_7010,N_2442,N_3576);
or U7011 (N_7011,N_4458,N_4557);
or U7012 (N_7012,N_161,N_2574);
xnor U7013 (N_7013,N_4220,N_21);
or U7014 (N_7014,N_1009,N_1660);
or U7015 (N_7015,N_987,N_3818);
or U7016 (N_7016,N_2739,N_4781);
or U7017 (N_7017,N_3415,N_1278);
nor U7018 (N_7018,N_3681,N_1622);
xnor U7019 (N_7019,N_3102,N_1131);
and U7020 (N_7020,N_3540,N_4757);
nand U7021 (N_7021,N_4960,N_146);
nor U7022 (N_7022,N_4555,N_909);
nand U7023 (N_7023,N_3081,N_3490);
or U7024 (N_7024,N_4741,N_2349);
xor U7025 (N_7025,N_1925,N_4632);
xor U7026 (N_7026,N_2993,N_302);
xnor U7027 (N_7027,N_3497,N_280);
nand U7028 (N_7028,N_149,N_167);
and U7029 (N_7029,N_3228,N_490);
and U7030 (N_7030,N_3259,N_1489);
and U7031 (N_7031,N_2805,N_3084);
and U7032 (N_7032,N_2008,N_3231);
and U7033 (N_7033,N_3634,N_3962);
nor U7034 (N_7034,N_4108,N_914);
xor U7035 (N_7035,N_392,N_4531);
and U7036 (N_7036,N_2056,N_599);
and U7037 (N_7037,N_616,N_2911);
xnor U7038 (N_7038,N_1159,N_487);
nand U7039 (N_7039,N_2952,N_3719);
nand U7040 (N_7040,N_1677,N_1244);
and U7041 (N_7041,N_3096,N_304);
nor U7042 (N_7042,N_107,N_993);
or U7043 (N_7043,N_928,N_1061);
xnor U7044 (N_7044,N_3297,N_1077);
nand U7045 (N_7045,N_4103,N_2563);
nor U7046 (N_7046,N_3320,N_1940);
and U7047 (N_7047,N_983,N_1697);
xnor U7048 (N_7048,N_3120,N_37);
nor U7049 (N_7049,N_1053,N_3017);
and U7050 (N_7050,N_4891,N_4145);
nand U7051 (N_7051,N_4095,N_1936);
nor U7052 (N_7052,N_927,N_3841);
xor U7053 (N_7053,N_1625,N_2401);
xnor U7054 (N_7054,N_2178,N_4802);
xnor U7055 (N_7055,N_3772,N_2248);
nor U7056 (N_7056,N_3395,N_2325);
or U7057 (N_7057,N_1181,N_3351);
and U7058 (N_7058,N_4813,N_2991);
or U7059 (N_7059,N_2978,N_2270);
xor U7060 (N_7060,N_4274,N_3912);
and U7061 (N_7061,N_786,N_2936);
or U7062 (N_7062,N_3644,N_4966);
and U7063 (N_7063,N_1856,N_45);
nand U7064 (N_7064,N_4606,N_163);
or U7065 (N_7065,N_3016,N_433);
nor U7066 (N_7066,N_4115,N_270);
xor U7067 (N_7067,N_2828,N_2562);
or U7068 (N_7068,N_3034,N_2363);
nor U7069 (N_7069,N_3881,N_1566);
nor U7070 (N_7070,N_1206,N_2949);
xnor U7071 (N_7071,N_2279,N_3283);
nor U7072 (N_7072,N_907,N_3786);
xnor U7073 (N_7073,N_210,N_1901);
xnor U7074 (N_7074,N_1641,N_3240);
or U7075 (N_7075,N_1662,N_2653);
or U7076 (N_7076,N_984,N_2691);
xor U7077 (N_7077,N_2124,N_1002);
nand U7078 (N_7078,N_1229,N_4909);
and U7079 (N_7079,N_1651,N_1454);
xnor U7080 (N_7080,N_2448,N_2053);
xnor U7081 (N_7081,N_3455,N_4586);
or U7082 (N_7082,N_3686,N_420);
xnor U7083 (N_7083,N_4239,N_1007);
nand U7084 (N_7084,N_4885,N_735);
nand U7085 (N_7085,N_4974,N_1559);
xnor U7086 (N_7086,N_2624,N_2050);
and U7087 (N_7087,N_2492,N_2555);
nand U7088 (N_7088,N_1455,N_2466);
nand U7089 (N_7089,N_2214,N_2168);
or U7090 (N_7090,N_2019,N_3988);
and U7091 (N_7091,N_4851,N_3157);
xnor U7092 (N_7092,N_4537,N_495);
nand U7093 (N_7093,N_221,N_2340);
nor U7094 (N_7094,N_1695,N_4031);
xnor U7095 (N_7095,N_122,N_1500);
nand U7096 (N_7096,N_393,N_4480);
xor U7097 (N_7097,N_8,N_3755);
or U7098 (N_7098,N_978,N_1724);
xnor U7099 (N_7099,N_902,N_3790);
or U7100 (N_7100,N_3365,N_3824);
nor U7101 (N_7101,N_1806,N_2900);
xor U7102 (N_7102,N_4827,N_1548);
nand U7103 (N_7103,N_1068,N_3702);
nand U7104 (N_7104,N_3583,N_3143);
nor U7105 (N_7105,N_3854,N_3037);
xnor U7106 (N_7106,N_3163,N_1711);
or U7107 (N_7107,N_859,N_2406);
and U7108 (N_7108,N_104,N_1877);
nand U7109 (N_7109,N_134,N_366);
nor U7110 (N_7110,N_1498,N_4581);
or U7111 (N_7111,N_2647,N_4205);
and U7112 (N_7112,N_1537,N_368);
xnor U7113 (N_7113,N_2859,N_1417);
nor U7114 (N_7114,N_3029,N_1246);
and U7115 (N_7115,N_886,N_1303);
or U7116 (N_7116,N_2499,N_4817);
nand U7117 (N_7117,N_2837,N_2970);
or U7118 (N_7118,N_3063,N_4958);
nand U7119 (N_7119,N_3057,N_4481);
nor U7120 (N_7120,N_4198,N_4321);
xnor U7121 (N_7121,N_4148,N_3257);
nor U7122 (N_7122,N_1160,N_3971);
or U7123 (N_7123,N_1307,N_3491);
or U7124 (N_7124,N_112,N_1978);
nand U7125 (N_7125,N_3811,N_3975);
nand U7126 (N_7126,N_1257,N_4638);
nand U7127 (N_7127,N_4925,N_3364);
nor U7128 (N_7128,N_4062,N_2021);
nor U7129 (N_7129,N_1227,N_2745);
or U7130 (N_7130,N_1917,N_2700);
nand U7131 (N_7131,N_1977,N_349);
and U7132 (N_7132,N_3266,N_1518);
xnor U7133 (N_7133,N_58,N_4034);
nor U7134 (N_7134,N_3711,N_1517);
or U7135 (N_7135,N_2205,N_3676);
nand U7136 (N_7136,N_2838,N_2843);
and U7137 (N_7137,N_4514,N_1255);
and U7138 (N_7138,N_2792,N_4474);
nor U7139 (N_7139,N_584,N_658);
or U7140 (N_7140,N_3368,N_2655);
nor U7141 (N_7141,N_1461,N_4772);
xnor U7142 (N_7142,N_3005,N_3735);
nor U7143 (N_7143,N_2684,N_1528);
xor U7144 (N_7144,N_233,N_3182);
xnor U7145 (N_7145,N_1474,N_2025);
xor U7146 (N_7146,N_2578,N_3553);
and U7147 (N_7147,N_4678,N_2821);
or U7148 (N_7148,N_3354,N_2751);
and U7149 (N_7149,N_3098,N_903);
xnor U7150 (N_7150,N_423,N_2130);
nor U7151 (N_7151,N_1934,N_3690);
or U7152 (N_7152,N_101,N_1252);
nor U7153 (N_7153,N_2331,N_4019);
xnor U7154 (N_7154,N_1522,N_353);
nor U7155 (N_7155,N_1019,N_2445);
nor U7156 (N_7156,N_1952,N_3645);
and U7157 (N_7157,N_4605,N_4351);
or U7158 (N_7158,N_916,N_2000);
or U7159 (N_7159,N_2118,N_4671);
nor U7160 (N_7160,N_4383,N_2469);
or U7161 (N_7161,N_919,N_4562);
nor U7162 (N_7162,N_3813,N_1440);
xor U7163 (N_7163,N_3080,N_2726);
xnor U7164 (N_7164,N_4938,N_4732);
or U7165 (N_7165,N_4313,N_4200);
nor U7166 (N_7166,N_1376,N_2803);
or U7167 (N_7167,N_4705,N_3304);
xnor U7168 (N_7168,N_3958,N_4162);
or U7169 (N_7169,N_3251,N_3166);
xnor U7170 (N_7170,N_2076,N_2195);
xnor U7171 (N_7171,N_1401,N_1698);
or U7172 (N_7172,N_944,N_581);
or U7173 (N_7173,N_1707,N_2109);
nor U7174 (N_7174,N_4421,N_1472);
xnor U7175 (N_7175,N_89,N_1268);
and U7176 (N_7176,N_1006,N_811);
xnor U7177 (N_7177,N_3501,N_4518);
or U7178 (N_7178,N_3239,N_437);
nand U7179 (N_7179,N_1351,N_2738);
xnor U7180 (N_7180,N_890,N_3180);
xor U7181 (N_7181,N_425,N_262);
or U7182 (N_7182,N_1109,N_2709);
xnor U7183 (N_7183,N_31,N_1134);
and U7184 (N_7184,N_168,N_2877);
and U7185 (N_7185,N_4577,N_3398);
nand U7186 (N_7186,N_4128,N_3926);
and U7187 (N_7187,N_1735,N_2802);
or U7188 (N_7188,N_4608,N_4522);
nor U7189 (N_7189,N_3914,N_69);
xor U7190 (N_7190,N_1254,N_4498);
and U7191 (N_7191,N_2407,N_2163);
xnor U7192 (N_7192,N_2516,N_1186);
xor U7193 (N_7193,N_2226,N_3298);
nor U7194 (N_7194,N_2117,N_172);
and U7195 (N_7195,N_4005,N_4240);
or U7196 (N_7196,N_1653,N_4041);
and U7197 (N_7197,N_1034,N_751);
or U7198 (N_7198,N_1191,N_3196);
and U7199 (N_7199,N_3588,N_1122);
nor U7200 (N_7200,N_3569,N_4469);
xor U7201 (N_7201,N_4792,N_1147);
or U7202 (N_7202,N_1319,N_4206);
xor U7203 (N_7203,N_4399,N_700);
or U7204 (N_7204,N_2464,N_757);
and U7205 (N_7205,N_1736,N_3086);
xnor U7206 (N_7206,N_1270,N_3246);
nand U7207 (N_7207,N_2026,N_4833);
nor U7208 (N_7208,N_2255,N_3689);
nor U7209 (N_7209,N_1725,N_3382);
nand U7210 (N_7210,N_989,N_3499);
nor U7211 (N_7211,N_4219,N_1840);
and U7212 (N_7212,N_3698,N_4288);
nor U7213 (N_7213,N_572,N_964);
nand U7214 (N_7214,N_4789,N_3858);
xor U7215 (N_7215,N_1330,N_2779);
and U7216 (N_7216,N_3306,N_4217);
and U7217 (N_7217,N_2580,N_1586);
xnor U7218 (N_7218,N_576,N_3876);
or U7219 (N_7219,N_3412,N_3794);
xor U7220 (N_7220,N_1366,N_116);
or U7221 (N_7221,N_3945,N_308);
xor U7222 (N_7222,N_514,N_4556);
nand U7223 (N_7223,N_136,N_1001);
and U7224 (N_7224,N_2350,N_715);
nor U7225 (N_7225,N_940,N_1821);
nand U7226 (N_7226,N_2687,N_2755);
nand U7227 (N_7227,N_2240,N_3054);
or U7228 (N_7228,N_941,N_2962);
xnor U7229 (N_7229,N_4937,N_1921);
xnor U7230 (N_7230,N_287,N_1023);
and U7231 (N_7231,N_479,N_826);
nand U7232 (N_7232,N_2549,N_1996);
or U7233 (N_7233,N_689,N_731);
nor U7234 (N_7234,N_2329,N_1086);
and U7235 (N_7235,N_997,N_3022);
nand U7236 (N_7236,N_2348,N_4953);
xnor U7237 (N_7237,N_192,N_4702);
nand U7238 (N_7238,N_232,N_4226);
or U7239 (N_7239,N_4856,N_578);
nor U7240 (N_7240,N_4225,N_4970);
nand U7241 (N_7241,N_4084,N_4835);
or U7242 (N_7242,N_3797,N_3927);
nor U7243 (N_7243,N_1599,N_2456);
nand U7244 (N_7244,N_1579,N_1481);
and U7245 (N_7245,N_714,N_1102);
nand U7246 (N_7246,N_4099,N_3806);
or U7247 (N_7247,N_3220,N_4908);
and U7248 (N_7248,N_4427,N_4487);
and U7249 (N_7249,N_4024,N_1827);
nand U7250 (N_7250,N_1098,N_1052);
and U7251 (N_7251,N_3522,N_445);
and U7252 (N_7252,N_1132,N_3928);
nor U7253 (N_7253,N_1418,N_1247);
nand U7254 (N_7254,N_4277,N_2230);
or U7255 (N_7255,N_51,N_2515);
and U7256 (N_7256,N_1720,N_1439);
xnor U7257 (N_7257,N_729,N_2335);
or U7258 (N_7258,N_4973,N_867);
or U7259 (N_7259,N_2997,N_3830);
and U7260 (N_7260,N_3976,N_769);
xor U7261 (N_7261,N_2893,N_418);
nor U7262 (N_7262,N_1965,N_2557);
or U7263 (N_7263,N_527,N_4438);
nand U7264 (N_7264,N_1907,N_96);
or U7265 (N_7265,N_2202,N_362);
or U7266 (N_7266,N_812,N_813);
nand U7267 (N_7267,N_4476,N_1969);
nand U7268 (N_7268,N_3106,N_2128);
xnor U7269 (N_7269,N_2964,N_430);
nor U7270 (N_7270,N_1045,N_3991);
nand U7271 (N_7271,N_4235,N_1265);
nand U7272 (N_7272,N_1811,N_4819);
nor U7273 (N_7273,N_4841,N_4387);
or U7274 (N_7274,N_2059,N_3496);
or U7275 (N_7275,N_3092,N_1298);
or U7276 (N_7276,N_743,N_4721);
nand U7277 (N_7277,N_2169,N_3332);
xnor U7278 (N_7278,N_3192,N_3000);
or U7279 (N_7279,N_2902,N_4491);
nand U7280 (N_7280,N_3513,N_2358);
or U7281 (N_7281,N_3596,N_1672);
nand U7282 (N_7282,N_3071,N_1260);
nor U7283 (N_7283,N_1010,N_2889);
xor U7284 (N_7284,N_46,N_957);
nor U7285 (N_7285,N_1411,N_4303);
nand U7286 (N_7286,N_4268,N_3478);
and U7287 (N_7287,N_1762,N_299);
and U7288 (N_7288,N_2001,N_2568);
and U7289 (N_7289,N_1479,N_80);
xor U7290 (N_7290,N_2762,N_549);
or U7291 (N_7291,N_763,N_2565);
or U7292 (N_7292,N_4622,N_1668);
nor U7293 (N_7293,N_4633,N_4610);
and U7294 (N_7294,N_3241,N_4464);
or U7295 (N_7295,N_162,N_3471);
xor U7296 (N_7296,N_3079,N_1501);
nor U7297 (N_7297,N_1434,N_4607);
nand U7298 (N_7298,N_557,N_276);
xnor U7299 (N_7299,N_2882,N_1511);
nor U7300 (N_7300,N_2024,N_435);
and U7301 (N_7301,N_1919,N_4855);
and U7302 (N_7302,N_2787,N_145);
and U7303 (N_7303,N_952,N_566);
and U7304 (N_7304,N_2677,N_2216);
or U7305 (N_7305,N_424,N_4497);
and U7306 (N_7306,N_2337,N_77);
nor U7307 (N_7307,N_3610,N_3015);
or U7308 (N_7308,N_4281,N_359);
xnor U7309 (N_7309,N_4592,N_677);
or U7310 (N_7310,N_1405,N_1568);
nand U7311 (N_7311,N_3025,N_3766);
xnor U7312 (N_7312,N_2961,N_177);
nor U7313 (N_7313,N_3193,N_972);
nand U7314 (N_7314,N_2852,N_841);
xnor U7315 (N_7315,N_570,N_2398);
or U7316 (N_7316,N_737,N_724);
or U7317 (N_7317,N_2233,N_664);
nor U7318 (N_7318,N_4764,N_879);
and U7319 (N_7319,N_3757,N_1659);
and U7320 (N_7320,N_1352,N_2022);
or U7321 (N_7321,N_2980,N_2111);
xor U7322 (N_7322,N_4901,N_3793);
and U7323 (N_7323,N_3456,N_992);
nor U7324 (N_7324,N_502,N_1234);
nand U7325 (N_7325,N_313,N_2681);
or U7326 (N_7326,N_1284,N_2108);
or U7327 (N_7327,N_3618,N_915);
nand U7328 (N_7328,N_3056,N_1942);
xor U7329 (N_7329,N_1593,N_2916);
xnor U7330 (N_7330,N_2115,N_3911);
or U7331 (N_7331,N_2141,N_3597);
and U7332 (N_7332,N_3745,N_1638);
nand U7333 (N_7333,N_272,N_4969);
or U7334 (N_7334,N_2607,N_852);
xnor U7335 (N_7335,N_2370,N_4184);
nand U7336 (N_7336,N_1087,N_396);
or U7337 (N_7337,N_40,N_630);
nor U7338 (N_7338,N_4352,N_2455);
xor U7339 (N_7339,N_2867,N_389);
xnor U7340 (N_7340,N_438,N_3374);
and U7341 (N_7341,N_3997,N_1592);
and U7342 (N_7342,N_2746,N_2825);
and U7343 (N_7343,N_382,N_2554);
nand U7344 (N_7344,N_543,N_186);
and U7345 (N_7345,N_4726,N_3541);
and U7346 (N_7346,N_2679,N_3119);
nand U7347 (N_7347,N_899,N_862);
nor U7348 (N_7348,N_991,N_4996);
and U7349 (N_7349,N_4377,N_4631);
nand U7350 (N_7350,N_67,N_4552);
or U7351 (N_7351,N_552,N_1162);
xor U7352 (N_7352,N_2285,N_3293);
nor U7353 (N_7353,N_4858,N_498);
xnor U7354 (N_7354,N_188,N_1205);
and U7355 (N_7355,N_2842,N_2776);
nand U7356 (N_7356,N_4520,N_1891);
or U7357 (N_7357,N_176,N_219);
xnor U7358 (N_7358,N_4436,N_1805);
or U7359 (N_7359,N_1467,N_1008);
nand U7360 (N_7360,N_475,N_1169);
nand U7361 (N_7361,N_1530,N_4360);
xor U7362 (N_7362,N_74,N_109);
and U7363 (N_7363,N_1974,N_3123);
and U7364 (N_7364,N_4211,N_1543);
or U7365 (N_7365,N_4574,N_1203);
nor U7366 (N_7366,N_4189,N_1619);
or U7367 (N_7367,N_4593,N_3393);
xor U7368 (N_7368,N_4890,N_3384);
xnor U7369 (N_7369,N_2690,N_2352);
xnor U7370 (N_7370,N_4943,N_4820);
nand U7371 (N_7371,N_1834,N_4971);
nor U7372 (N_7372,N_2006,N_942);
or U7373 (N_7373,N_877,N_1030);
nand U7374 (N_7374,N_1928,N_612);
xor U7375 (N_7375,N_779,N_2497);
nor U7376 (N_7376,N_1428,N_3003);
or U7377 (N_7377,N_2075,N_3859);
nor U7378 (N_7378,N_1130,N_3761);
nor U7379 (N_7379,N_4729,N_126);
nand U7380 (N_7380,N_3780,N_3701);
xor U7381 (N_7381,N_4511,N_3058);
xnor U7382 (N_7382,N_2481,N_3210);
nor U7383 (N_7383,N_4647,N_380);
and U7384 (N_7384,N_3282,N_142);
or U7385 (N_7385,N_337,N_960);
or U7386 (N_7386,N_4002,N_4818);
nand U7387 (N_7387,N_4179,N_3146);
or U7388 (N_7388,N_4590,N_4806);
xor U7389 (N_7389,N_3853,N_213);
nand U7390 (N_7390,N_1515,N_803);
nor U7391 (N_7391,N_35,N_1354);
or U7392 (N_7392,N_1123,N_2839);
or U7393 (N_7393,N_1681,N_875);
and U7394 (N_7394,N_4305,N_2431);
nor U7395 (N_7395,N_3434,N_258);
xnor U7396 (N_7396,N_1269,N_4129);
xnor U7397 (N_7397,N_4888,N_1884);
nor U7398 (N_7398,N_2236,N_363);
and U7399 (N_7399,N_2391,N_206);
or U7400 (N_7400,N_2917,N_3197);
xor U7401 (N_7401,N_1602,N_2457);
and U7402 (N_7402,N_3973,N_2899);
nand U7403 (N_7403,N_4499,N_2648);
xor U7404 (N_7404,N_750,N_3543);
nand U7405 (N_7405,N_3680,N_2032);
or U7406 (N_7406,N_2339,N_2870);
xnor U7407 (N_7407,N_2153,N_4563);
xor U7408 (N_7408,N_3167,N_4282);
nor U7409 (N_7409,N_898,N_3363);
nand U7410 (N_7410,N_3362,N_4232);
and U7411 (N_7411,N_2950,N_3099);
xor U7412 (N_7412,N_583,N_3882);
xnor U7413 (N_7413,N_3687,N_4241);
xnor U7414 (N_7414,N_454,N_4307);
or U7415 (N_7415,N_3922,N_4540);
and U7416 (N_7416,N_4400,N_2454);
or U7417 (N_7417,N_2386,N_3878);
nand U7418 (N_7418,N_765,N_2886);
xnor U7419 (N_7419,N_504,N_686);
nor U7420 (N_7420,N_1556,N_3949);
and U7421 (N_7421,N_1100,N_4755);
or U7422 (N_7422,N_733,N_2652);
nor U7423 (N_7423,N_3189,N_1715);
nor U7424 (N_7424,N_1595,N_3839);
or U7425 (N_7425,N_799,N_4558);
and U7426 (N_7426,N_469,N_2729);
nor U7427 (N_7427,N_4594,N_2266);
nor U7428 (N_7428,N_1748,N_3472);
nand U7429 (N_7429,N_3860,N_1564);
and U7430 (N_7430,N_1683,N_3419);
nand U7431 (N_7431,N_2918,N_3483);
nor U7432 (N_7432,N_2176,N_4169);
nand U7433 (N_7433,N_6,N_4155);
xor U7434 (N_7434,N_4193,N_846);
xor U7435 (N_7435,N_2465,N_4763);
nand U7436 (N_7436,N_3142,N_1380);
nor U7437 (N_7437,N_4044,N_2720);
or U7438 (N_7438,N_2146,N_4838);
or U7439 (N_7439,N_4122,N_4028);
nor U7440 (N_7440,N_4516,N_1240);
xor U7441 (N_7441,N_2160,N_2758);
xnor U7442 (N_7442,N_4681,N_1639);
or U7443 (N_7443,N_303,N_2067);
or U7444 (N_7444,N_4854,N_3091);
nor U7445 (N_7445,N_165,N_3875);
or U7446 (N_7446,N_4027,N_408);
xnor U7447 (N_7447,N_338,N_491);
nand U7448 (N_7448,N_1646,N_400);
nand U7449 (N_7449,N_1062,N_4405);
xor U7450 (N_7450,N_4411,N_3758);
nor U7451 (N_7451,N_4982,N_3620);
nand U7452 (N_7452,N_2140,N_2880);
xor U7453 (N_7453,N_1867,N_339);
xnor U7454 (N_7454,N_361,N_2311);
or U7455 (N_7455,N_1072,N_2089);
nand U7456 (N_7456,N_3315,N_1634);
nor U7457 (N_7457,N_3453,N_874);
xor U7458 (N_7458,N_1262,N_2);
nand U7459 (N_7459,N_224,N_3581);
nor U7460 (N_7460,N_241,N_4904);
or U7461 (N_7461,N_4382,N_3308);
or U7462 (N_7462,N_20,N_4990);
or U7463 (N_7463,N_98,N_3432);
or U7464 (N_7464,N_979,N_2963);
or U7465 (N_7465,N_4554,N_2521);
nand U7466 (N_7466,N_2254,N_4063);
or U7467 (N_7467,N_1769,N_3426);
xor U7468 (N_7468,N_788,N_3036);
or U7469 (N_7469,N_1294,N_4143);
nand U7470 (N_7470,N_3329,N_215);
nand U7471 (N_7471,N_319,N_2382);
nor U7472 (N_7472,N_721,N_893);
nor U7473 (N_7473,N_124,N_3075);
nor U7474 (N_7474,N_3641,N_2122);
or U7475 (N_7475,N_4836,N_325);
and U7476 (N_7476,N_3523,N_3695);
nand U7477 (N_7477,N_1231,N_2959);
and U7478 (N_7478,N_4414,N_1200);
and U7479 (N_7479,N_1787,N_2064);
and U7480 (N_7480,N_2368,N_1256);
or U7481 (N_7481,N_1443,N_2449);
or U7482 (N_7482,N_1143,N_753);
and U7483 (N_7483,N_1533,N_1993);
nand U7484 (N_7484,N_3340,N_4258);
nor U7485 (N_7485,N_4614,N_722);
or U7486 (N_7486,N_939,N_2123);
or U7487 (N_7487,N_3125,N_4234);
and U7488 (N_7488,N_4805,N_1731);
nor U7489 (N_7489,N_1963,N_4008);
or U7490 (N_7490,N_263,N_2571);
nor U7491 (N_7491,N_56,N_4359);
xnor U7492 (N_7492,N_953,N_3052);
or U7493 (N_7493,N_2559,N_4935);
or U7494 (N_7494,N_3334,N_3751);
and U7495 (N_7495,N_2225,N_4668);
or U7496 (N_7496,N_2643,N_3992);
xnor U7497 (N_7497,N_807,N_519);
and U7498 (N_7498,N_1544,N_259);
nand U7499 (N_7499,N_4800,N_755);
or U7500 (N_7500,N_799,N_4162);
or U7501 (N_7501,N_2479,N_4442);
or U7502 (N_7502,N_4910,N_1321);
and U7503 (N_7503,N_3889,N_3938);
and U7504 (N_7504,N_3817,N_2342);
and U7505 (N_7505,N_1208,N_3064);
nand U7506 (N_7506,N_3519,N_704);
nor U7507 (N_7507,N_1406,N_3853);
or U7508 (N_7508,N_1585,N_628);
nand U7509 (N_7509,N_575,N_4579);
xor U7510 (N_7510,N_1791,N_294);
nand U7511 (N_7511,N_2335,N_2152);
and U7512 (N_7512,N_2072,N_2215);
nor U7513 (N_7513,N_2535,N_436);
and U7514 (N_7514,N_2000,N_3763);
xor U7515 (N_7515,N_4170,N_3701);
and U7516 (N_7516,N_3478,N_1050);
xor U7517 (N_7517,N_2017,N_4919);
and U7518 (N_7518,N_2574,N_4910);
nand U7519 (N_7519,N_237,N_4512);
nor U7520 (N_7520,N_4786,N_1226);
or U7521 (N_7521,N_1470,N_3634);
nand U7522 (N_7522,N_1896,N_1972);
or U7523 (N_7523,N_3526,N_3949);
nand U7524 (N_7524,N_2179,N_3671);
xnor U7525 (N_7525,N_764,N_4752);
xnor U7526 (N_7526,N_404,N_1607);
and U7527 (N_7527,N_195,N_547);
and U7528 (N_7528,N_2168,N_2011);
nand U7529 (N_7529,N_469,N_2797);
and U7530 (N_7530,N_4215,N_4533);
nand U7531 (N_7531,N_3788,N_1582);
nor U7532 (N_7532,N_649,N_4334);
nor U7533 (N_7533,N_254,N_2388);
xor U7534 (N_7534,N_3950,N_2947);
xnor U7535 (N_7535,N_4781,N_3246);
or U7536 (N_7536,N_2285,N_3657);
xnor U7537 (N_7537,N_2629,N_1850);
or U7538 (N_7538,N_1908,N_2437);
nand U7539 (N_7539,N_2693,N_4164);
xor U7540 (N_7540,N_1011,N_7);
nand U7541 (N_7541,N_3926,N_4075);
xor U7542 (N_7542,N_125,N_3164);
and U7543 (N_7543,N_1458,N_2770);
and U7544 (N_7544,N_4238,N_4321);
xor U7545 (N_7545,N_15,N_1575);
nand U7546 (N_7546,N_405,N_948);
nor U7547 (N_7547,N_4673,N_4608);
xnor U7548 (N_7548,N_3643,N_1359);
nor U7549 (N_7549,N_4877,N_2023);
or U7550 (N_7550,N_4959,N_4819);
and U7551 (N_7551,N_2197,N_892);
xor U7552 (N_7552,N_3591,N_387);
xnor U7553 (N_7553,N_249,N_1157);
nand U7554 (N_7554,N_3952,N_1099);
nand U7555 (N_7555,N_138,N_208);
nand U7556 (N_7556,N_1819,N_233);
or U7557 (N_7557,N_1182,N_3810);
and U7558 (N_7558,N_3649,N_3053);
nand U7559 (N_7559,N_4787,N_176);
xnor U7560 (N_7560,N_2160,N_3923);
nand U7561 (N_7561,N_1467,N_990);
xnor U7562 (N_7562,N_3378,N_4068);
and U7563 (N_7563,N_1004,N_3072);
nand U7564 (N_7564,N_3205,N_2380);
nand U7565 (N_7565,N_1603,N_2090);
or U7566 (N_7566,N_3814,N_827);
nand U7567 (N_7567,N_3594,N_1552);
nand U7568 (N_7568,N_2052,N_4794);
nand U7569 (N_7569,N_3647,N_3364);
or U7570 (N_7570,N_319,N_3259);
nand U7571 (N_7571,N_3125,N_2259);
nor U7572 (N_7572,N_3319,N_1277);
nand U7573 (N_7573,N_2781,N_2600);
nand U7574 (N_7574,N_3619,N_2705);
or U7575 (N_7575,N_2904,N_4837);
xor U7576 (N_7576,N_4725,N_1568);
nand U7577 (N_7577,N_469,N_3628);
nand U7578 (N_7578,N_1509,N_1148);
xnor U7579 (N_7579,N_619,N_783);
nand U7580 (N_7580,N_4149,N_173);
xnor U7581 (N_7581,N_389,N_1223);
or U7582 (N_7582,N_649,N_1706);
xor U7583 (N_7583,N_1941,N_3826);
xor U7584 (N_7584,N_3592,N_4489);
xor U7585 (N_7585,N_2700,N_4987);
xor U7586 (N_7586,N_121,N_3043);
xnor U7587 (N_7587,N_1851,N_3431);
nor U7588 (N_7588,N_4710,N_3919);
nand U7589 (N_7589,N_4380,N_4888);
nor U7590 (N_7590,N_321,N_2797);
and U7591 (N_7591,N_4772,N_2993);
nor U7592 (N_7592,N_4187,N_1928);
nand U7593 (N_7593,N_4487,N_4711);
xnor U7594 (N_7594,N_489,N_2157);
and U7595 (N_7595,N_1771,N_828);
or U7596 (N_7596,N_1405,N_4977);
nor U7597 (N_7597,N_2425,N_827);
nor U7598 (N_7598,N_2463,N_944);
nor U7599 (N_7599,N_4400,N_1334);
xor U7600 (N_7600,N_4180,N_3112);
and U7601 (N_7601,N_3236,N_9);
nor U7602 (N_7602,N_2563,N_1703);
nand U7603 (N_7603,N_2063,N_3678);
and U7604 (N_7604,N_3917,N_3171);
nor U7605 (N_7605,N_2346,N_311);
nor U7606 (N_7606,N_4785,N_3403);
nand U7607 (N_7607,N_4438,N_4666);
and U7608 (N_7608,N_4977,N_3746);
and U7609 (N_7609,N_4474,N_1374);
xnor U7610 (N_7610,N_4090,N_4446);
nor U7611 (N_7611,N_888,N_4747);
nand U7612 (N_7612,N_1743,N_3279);
or U7613 (N_7613,N_2456,N_746);
and U7614 (N_7614,N_4864,N_4549);
or U7615 (N_7615,N_195,N_1765);
xnor U7616 (N_7616,N_817,N_4111);
or U7617 (N_7617,N_314,N_3371);
or U7618 (N_7618,N_4328,N_3453);
nand U7619 (N_7619,N_130,N_4700);
xnor U7620 (N_7620,N_4764,N_1684);
nor U7621 (N_7621,N_3542,N_3751);
xnor U7622 (N_7622,N_2673,N_1223);
nor U7623 (N_7623,N_4117,N_925);
nor U7624 (N_7624,N_432,N_3013);
nand U7625 (N_7625,N_2525,N_4464);
xnor U7626 (N_7626,N_2496,N_4823);
nand U7627 (N_7627,N_4642,N_675);
nor U7628 (N_7628,N_1959,N_2325);
nor U7629 (N_7629,N_1983,N_1213);
or U7630 (N_7630,N_3142,N_3479);
nor U7631 (N_7631,N_1836,N_4841);
or U7632 (N_7632,N_255,N_2332);
or U7633 (N_7633,N_1450,N_2199);
nand U7634 (N_7634,N_4819,N_968);
xnor U7635 (N_7635,N_1611,N_4174);
nor U7636 (N_7636,N_2358,N_3216);
and U7637 (N_7637,N_2927,N_3383);
xnor U7638 (N_7638,N_1744,N_3855);
xor U7639 (N_7639,N_4517,N_448);
or U7640 (N_7640,N_1671,N_4759);
and U7641 (N_7641,N_3639,N_590);
nand U7642 (N_7642,N_3881,N_4387);
xor U7643 (N_7643,N_2162,N_3595);
or U7644 (N_7644,N_3647,N_1792);
xor U7645 (N_7645,N_4898,N_3612);
xnor U7646 (N_7646,N_35,N_909);
xnor U7647 (N_7647,N_2489,N_3388);
and U7648 (N_7648,N_124,N_3748);
xnor U7649 (N_7649,N_425,N_1273);
or U7650 (N_7650,N_1708,N_3615);
xor U7651 (N_7651,N_1527,N_4103);
xor U7652 (N_7652,N_4002,N_2871);
and U7653 (N_7653,N_3018,N_1961);
and U7654 (N_7654,N_3912,N_4500);
and U7655 (N_7655,N_1448,N_3161);
or U7656 (N_7656,N_74,N_4064);
or U7657 (N_7657,N_4839,N_1514);
xnor U7658 (N_7658,N_2583,N_4969);
or U7659 (N_7659,N_1588,N_2450);
xor U7660 (N_7660,N_3985,N_3824);
and U7661 (N_7661,N_1997,N_4703);
nor U7662 (N_7662,N_395,N_2155);
or U7663 (N_7663,N_2349,N_3729);
nor U7664 (N_7664,N_2706,N_3717);
nor U7665 (N_7665,N_2857,N_2507);
and U7666 (N_7666,N_2121,N_2629);
nand U7667 (N_7667,N_3952,N_3581);
nor U7668 (N_7668,N_1121,N_1475);
nand U7669 (N_7669,N_4162,N_1340);
and U7670 (N_7670,N_3503,N_1885);
and U7671 (N_7671,N_1687,N_3394);
and U7672 (N_7672,N_722,N_4865);
and U7673 (N_7673,N_125,N_139);
nor U7674 (N_7674,N_2001,N_4520);
and U7675 (N_7675,N_4099,N_3410);
xnor U7676 (N_7676,N_351,N_111);
nor U7677 (N_7677,N_4672,N_4712);
and U7678 (N_7678,N_4942,N_2894);
and U7679 (N_7679,N_4725,N_2163);
nor U7680 (N_7680,N_4512,N_1341);
nor U7681 (N_7681,N_1105,N_4089);
nand U7682 (N_7682,N_1539,N_1978);
or U7683 (N_7683,N_1857,N_4307);
nor U7684 (N_7684,N_3345,N_4182);
xnor U7685 (N_7685,N_570,N_2207);
xnor U7686 (N_7686,N_4921,N_3851);
and U7687 (N_7687,N_3616,N_4914);
or U7688 (N_7688,N_4736,N_512);
and U7689 (N_7689,N_4224,N_2553);
and U7690 (N_7690,N_1344,N_4467);
nor U7691 (N_7691,N_4527,N_4100);
nand U7692 (N_7692,N_3413,N_92);
nor U7693 (N_7693,N_416,N_3206);
nor U7694 (N_7694,N_4134,N_4926);
xnor U7695 (N_7695,N_776,N_2975);
or U7696 (N_7696,N_2124,N_860);
nand U7697 (N_7697,N_498,N_2851);
or U7698 (N_7698,N_1166,N_944);
nor U7699 (N_7699,N_1777,N_2445);
or U7700 (N_7700,N_2147,N_4398);
nor U7701 (N_7701,N_1119,N_3845);
or U7702 (N_7702,N_4031,N_3879);
and U7703 (N_7703,N_1571,N_3000);
nor U7704 (N_7704,N_2750,N_3335);
xor U7705 (N_7705,N_297,N_4376);
nor U7706 (N_7706,N_4979,N_370);
nor U7707 (N_7707,N_2876,N_3579);
and U7708 (N_7708,N_2894,N_789);
or U7709 (N_7709,N_1051,N_58);
or U7710 (N_7710,N_4702,N_3988);
nand U7711 (N_7711,N_4808,N_1755);
and U7712 (N_7712,N_1787,N_4950);
and U7713 (N_7713,N_3780,N_1426);
or U7714 (N_7714,N_3147,N_1409);
nand U7715 (N_7715,N_4790,N_1401);
nor U7716 (N_7716,N_2187,N_2296);
xor U7717 (N_7717,N_414,N_1770);
nor U7718 (N_7718,N_2737,N_609);
nand U7719 (N_7719,N_3504,N_2955);
and U7720 (N_7720,N_3253,N_2686);
nor U7721 (N_7721,N_4816,N_2159);
xor U7722 (N_7722,N_3729,N_4952);
and U7723 (N_7723,N_1746,N_3120);
and U7724 (N_7724,N_1640,N_2030);
or U7725 (N_7725,N_4253,N_4646);
xnor U7726 (N_7726,N_3542,N_4692);
nand U7727 (N_7727,N_3700,N_251);
and U7728 (N_7728,N_4108,N_2070);
xnor U7729 (N_7729,N_1685,N_4413);
and U7730 (N_7730,N_382,N_2168);
and U7731 (N_7731,N_1661,N_2949);
and U7732 (N_7732,N_2822,N_3570);
nand U7733 (N_7733,N_1380,N_2656);
nand U7734 (N_7734,N_1599,N_932);
nor U7735 (N_7735,N_785,N_2320);
and U7736 (N_7736,N_1743,N_3940);
or U7737 (N_7737,N_983,N_1049);
and U7738 (N_7738,N_4999,N_1082);
nand U7739 (N_7739,N_2602,N_4164);
nor U7740 (N_7740,N_4909,N_3388);
nand U7741 (N_7741,N_3087,N_453);
or U7742 (N_7742,N_272,N_2354);
and U7743 (N_7743,N_1809,N_3126);
nor U7744 (N_7744,N_2757,N_3968);
or U7745 (N_7745,N_2614,N_2956);
xnor U7746 (N_7746,N_1715,N_3354);
or U7747 (N_7747,N_4720,N_1452);
or U7748 (N_7748,N_1239,N_1070);
xor U7749 (N_7749,N_3610,N_675);
xnor U7750 (N_7750,N_4007,N_2731);
nand U7751 (N_7751,N_4105,N_4648);
xnor U7752 (N_7752,N_4061,N_3620);
nor U7753 (N_7753,N_4231,N_4324);
xnor U7754 (N_7754,N_4827,N_4440);
xnor U7755 (N_7755,N_3942,N_23);
xor U7756 (N_7756,N_823,N_2088);
and U7757 (N_7757,N_2134,N_4426);
nor U7758 (N_7758,N_3097,N_1554);
nand U7759 (N_7759,N_44,N_62);
and U7760 (N_7760,N_3687,N_4644);
xnor U7761 (N_7761,N_4512,N_3505);
nand U7762 (N_7762,N_4023,N_4634);
nor U7763 (N_7763,N_1621,N_1830);
xor U7764 (N_7764,N_4945,N_2052);
nor U7765 (N_7765,N_1687,N_1289);
xor U7766 (N_7766,N_1192,N_3004);
nand U7767 (N_7767,N_1972,N_146);
and U7768 (N_7768,N_2546,N_2137);
or U7769 (N_7769,N_2580,N_4658);
or U7770 (N_7770,N_93,N_3666);
nor U7771 (N_7771,N_1191,N_4034);
xor U7772 (N_7772,N_1977,N_2206);
or U7773 (N_7773,N_75,N_2735);
or U7774 (N_7774,N_2367,N_2596);
xor U7775 (N_7775,N_1156,N_352);
xor U7776 (N_7776,N_2975,N_589);
or U7777 (N_7777,N_1084,N_1479);
or U7778 (N_7778,N_1091,N_1981);
or U7779 (N_7779,N_4071,N_2162);
nor U7780 (N_7780,N_4569,N_3422);
and U7781 (N_7781,N_3491,N_1554);
nand U7782 (N_7782,N_2472,N_1572);
xnor U7783 (N_7783,N_2807,N_3742);
nand U7784 (N_7784,N_29,N_1775);
nor U7785 (N_7785,N_2481,N_1226);
xor U7786 (N_7786,N_1573,N_3765);
nand U7787 (N_7787,N_1025,N_4184);
nor U7788 (N_7788,N_1912,N_4932);
and U7789 (N_7789,N_4700,N_1587);
and U7790 (N_7790,N_2753,N_2425);
xor U7791 (N_7791,N_867,N_1667);
or U7792 (N_7792,N_652,N_2346);
or U7793 (N_7793,N_1153,N_1145);
or U7794 (N_7794,N_4093,N_2136);
nor U7795 (N_7795,N_625,N_4892);
nand U7796 (N_7796,N_3573,N_1526);
nand U7797 (N_7797,N_366,N_3481);
nor U7798 (N_7798,N_2786,N_4389);
xnor U7799 (N_7799,N_1142,N_4931);
xnor U7800 (N_7800,N_435,N_2315);
and U7801 (N_7801,N_2183,N_1157);
nor U7802 (N_7802,N_4196,N_1183);
xor U7803 (N_7803,N_2721,N_1483);
and U7804 (N_7804,N_639,N_4361);
and U7805 (N_7805,N_2121,N_3666);
nand U7806 (N_7806,N_4313,N_3447);
nor U7807 (N_7807,N_4803,N_4110);
xnor U7808 (N_7808,N_1771,N_4570);
and U7809 (N_7809,N_1943,N_739);
or U7810 (N_7810,N_4923,N_64);
or U7811 (N_7811,N_1158,N_121);
and U7812 (N_7812,N_1548,N_626);
and U7813 (N_7813,N_3076,N_1379);
nand U7814 (N_7814,N_1388,N_807);
xnor U7815 (N_7815,N_1412,N_1120);
nor U7816 (N_7816,N_1105,N_2205);
xor U7817 (N_7817,N_2498,N_4689);
nand U7818 (N_7818,N_1122,N_2615);
nor U7819 (N_7819,N_3919,N_3472);
nor U7820 (N_7820,N_3060,N_128);
xnor U7821 (N_7821,N_4548,N_2267);
or U7822 (N_7822,N_1634,N_1348);
and U7823 (N_7823,N_1154,N_3416);
xnor U7824 (N_7824,N_2388,N_1212);
or U7825 (N_7825,N_4429,N_1611);
nand U7826 (N_7826,N_3631,N_4005);
xnor U7827 (N_7827,N_4107,N_2066);
xnor U7828 (N_7828,N_3649,N_4238);
xnor U7829 (N_7829,N_3594,N_3804);
or U7830 (N_7830,N_3705,N_2488);
and U7831 (N_7831,N_932,N_1129);
or U7832 (N_7832,N_4231,N_1348);
nand U7833 (N_7833,N_103,N_372);
nand U7834 (N_7834,N_902,N_962);
nor U7835 (N_7835,N_785,N_2864);
xor U7836 (N_7836,N_2199,N_3170);
nand U7837 (N_7837,N_1023,N_1244);
nor U7838 (N_7838,N_2519,N_2940);
nand U7839 (N_7839,N_981,N_4401);
nand U7840 (N_7840,N_714,N_4254);
nand U7841 (N_7841,N_4180,N_2741);
and U7842 (N_7842,N_3228,N_4222);
xnor U7843 (N_7843,N_1155,N_2822);
or U7844 (N_7844,N_155,N_1886);
nand U7845 (N_7845,N_4718,N_2975);
xor U7846 (N_7846,N_1490,N_4776);
nor U7847 (N_7847,N_219,N_4470);
nor U7848 (N_7848,N_2756,N_521);
xnor U7849 (N_7849,N_1867,N_2575);
nor U7850 (N_7850,N_4753,N_1470);
or U7851 (N_7851,N_4981,N_2146);
or U7852 (N_7852,N_1979,N_1796);
or U7853 (N_7853,N_4048,N_4190);
xor U7854 (N_7854,N_1451,N_2835);
xnor U7855 (N_7855,N_1979,N_1582);
and U7856 (N_7856,N_698,N_3766);
nand U7857 (N_7857,N_2646,N_273);
nor U7858 (N_7858,N_170,N_3869);
or U7859 (N_7859,N_302,N_2769);
nor U7860 (N_7860,N_4414,N_3913);
nor U7861 (N_7861,N_55,N_4039);
or U7862 (N_7862,N_3292,N_3389);
xor U7863 (N_7863,N_2084,N_592);
nor U7864 (N_7864,N_4626,N_2504);
or U7865 (N_7865,N_4862,N_4039);
or U7866 (N_7866,N_1579,N_4058);
or U7867 (N_7867,N_16,N_1803);
and U7868 (N_7868,N_2516,N_3783);
nor U7869 (N_7869,N_1172,N_3848);
or U7870 (N_7870,N_1313,N_4786);
nand U7871 (N_7871,N_3328,N_2196);
nand U7872 (N_7872,N_2739,N_2118);
and U7873 (N_7873,N_2332,N_2203);
and U7874 (N_7874,N_3830,N_3421);
or U7875 (N_7875,N_4083,N_1749);
xor U7876 (N_7876,N_320,N_2308);
or U7877 (N_7877,N_2535,N_2326);
xor U7878 (N_7878,N_1667,N_1283);
and U7879 (N_7879,N_1437,N_3334);
nor U7880 (N_7880,N_2015,N_3974);
nand U7881 (N_7881,N_3311,N_977);
or U7882 (N_7882,N_190,N_4724);
and U7883 (N_7883,N_2266,N_680);
and U7884 (N_7884,N_3538,N_1711);
or U7885 (N_7885,N_557,N_209);
or U7886 (N_7886,N_3977,N_1636);
or U7887 (N_7887,N_2418,N_1566);
and U7888 (N_7888,N_2666,N_2665);
and U7889 (N_7889,N_3045,N_4845);
xnor U7890 (N_7890,N_3507,N_4645);
and U7891 (N_7891,N_4619,N_3426);
xnor U7892 (N_7892,N_4642,N_3057);
and U7893 (N_7893,N_273,N_3824);
xnor U7894 (N_7894,N_3677,N_1879);
and U7895 (N_7895,N_676,N_4265);
and U7896 (N_7896,N_830,N_3887);
xnor U7897 (N_7897,N_608,N_1272);
or U7898 (N_7898,N_2602,N_4733);
or U7899 (N_7899,N_1275,N_2132);
nand U7900 (N_7900,N_3822,N_2140);
nor U7901 (N_7901,N_2935,N_3980);
and U7902 (N_7902,N_4671,N_2986);
nor U7903 (N_7903,N_3247,N_3750);
or U7904 (N_7904,N_3362,N_2248);
and U7905 (N_7905,N_1428,N_4477);
and U7906 (N_7906,N_2419,N_548);
nand U7907 (N_7907,N_4441,N_3737);
nand U7908 (N_7908,N_1452,N_2078);
nor U7909 (N_7909,N_2356,N_2037);
xor U7910 (N_7910,N_1631,N_4732);
nor U7911 (N_7911,N_1096,N_2004);
or U7912 (N_7912,N_4917,N_4677);
xor U7913 (N_7913,N_2404,N_2205);
or U7914 (N_7914,N_1822,N_1638);
xnor U7915 (N_7915,N_4371,N_2194);
nor U7916 (N_7916,N_229,N_414);
or U7917 (N_7917,N_223,N_2997);
xor U7918 (N_7918,N_1694,N_233);
or U7919 (N_7919,N_658,N_50);
or U7920 (N_7920,N_1145,N_4152);
nand U7921 (N_7921,N_293,N_598);
xor U7922 (N_7922,N_4080,N_2544);
nor U7923 (N_7923,N_1781,N_2433);
or U7924 (N_7924,N_378,N_1160);
nand U7925 (N_7925,N_1682,N_521);
and U7926 (N_7926,N_1264,N_3514);
and U7927 (N_7927,N_1868,N_2977);
xnor U7928 (N_7928,N_3271,N_1040);
xnor U7929 (N_7929,N_4344,N_2667);
and U7930 (N_7930,N_3978,N_4195);
nand U7931 (N_7931,N_2174,N_220);
xor U7932 (N_7932,N_1337,N_3734);
nor U7933 (N_7933,N_1677,N_3031);
xnor U7934 (N_7934,N_562,N_57);
nand U7935 (N_7935,N_1014,N_3113);
nor U7936 (N_7936,N_3535,N_1045);
nor U7937 (N_7937,N_3382,N_3523);
nor U7938 (N_7938,N_1103,N_2050);
and U7939 (N_7939,N_3175,N_4368);
xnor U7940 (N_7940,N_4286,N_2068);
and U7941 (N_7941,N_3981,N_2886);
nor U7942 (N_7942,N_640,N_171);
nor U7943 (N_7943,N_780,N_1236);
nand U7944 (N_7944,N_272,N_4982);
xnor U7945 (N_7945,N_3411,N_238);
xnor U7946 (N_7946,N_3108,N_4197);
nand U7947 (N_7947,N_59,N_3613);
or U7948 (N_7948,N_944,N_3863);
or U7949 (N_7949,N_461,N_1319);
nand U7950 (N_7950,N_603,N_1942);
nor U7951 (N_7951,N_2271,N_254);
xor U7952 (N_7952,N_4561,N_71);
nand U7953 (N_7953,N_316,N_2626);
xnor U7954 (N_7954,N_1745,N_1228);
nand U7955 (N_7955,N_4347,N_4840);
and U7956 (N_7956,N_4255,N_511);
or U7957 (N_7957,N_2474,N_4289);
nor U7958 (N_7958,N_2295,N_1744);
nor U7959 (N_7959,N_481,N_3242);
and U7960 (N_7960,N_28,N_1055);
nor U7961 (N_7961,N_2276,N_2301);
nor U7962 (N_7962,N_944,N_4349);
or U7963 (N_7963,N_4986,N_2874);
nor U7964 (N_7964,N_1960,N_3556);
nor U7965 (N_7965,N_3708,N_285);
or U7966 (N_7966,N_2384,N_4043);
and U7967 (N_7967,N_298,N_1407);
and U7968 (N_7968,N_3996,N_364);
nand U7969 (N_7969,N_44,N_225);
nand U7970 (N_7970,N_3399,N_3701);
nor U7971 (N_7971,N_2867,N_1867);
xnor U7972 (N_7972,N_3919,N_3127);
nor U7973 (N_7973,N_1865,N_2707);
nor U7974 (N_7974,N_1372,N_2135);
nor U7975 (N_7975,N_1152,N_3546);
nor U7976 (N_7976,N_3252,N_1444);
or U7977 (N_7977,N_1382,N_450);
xnor U7978 (N_7978,N_3957,N_1255);
nor U7979 (N_7979,N_3487,N_3332);
or U7980 (N_7980,N_4871,N_3413);
or U7981 (N_7981,N_4670,N_2293);
xnor U7982 (N_7982,N_3380,N_1679);
xor U7983 (N_7983,N_3703,N_4849);
nand U7984 (N_7984,N_1976,N_3017);
nand U7985 (N_7985,N_1164,N_2730);
xnor U7986 (N_7986,N_3358,N_779);
xor U7987 (N_7987,N_4820,N_1746);
and U7988 (N_7988,N_1301,N_2867);
xnor U7989 (N_7989,N_1332,N_990);
and U7990 (N_7990,N_1417,N_2595);
nor U7991 (N_7991,N_3404,N_1152);
or U7992 (N_7992,N_4861,N_3185);
or U7993 (N_7993,N_2412,N_3765);
nor U7994 (N_7994,N_4691,N_2540);
and U7995 (N_7995,N_3110,N_2101);
and U7996 (N_7996,N_141,N_4604);
xnor U7997 (N_7997,N_368,N_4031);
and U7998 (N_7998,N_4282,N_2460);
nand U7999 (N_7999,N_3824,N_2229);
or U8000 (N_8000,N_504,N_2310);
and U8001 (N_8001,N_828,N_3861);
or U8002 (N_8002,N_4019,N_4674);
nor U8003 (N_8003,N_1367,N_2467);
nor U8004 (N_8004,N_4730,N_1736);
nand U8005 (N_8005,N_3844,N_481);
nand U8006 (N_8006,N_3274,N_3932);
nand U8007 (N_8007,N_2213,N_4574);
nor U8008 (N_8008,N_1386,N_1559);
and U8009 (N_8009,N_4885,N_2479);
nand U8010 (N_8010,N_3896,N_205);
nor U8011 (N_8011,N_2513,N_4734);
nand U8012 (N_8012,N_3865,N_135);
xnor U8013 (N_8013,N_1504,N_4249);
nor U8014 (N_8014,N_1306,N_4589);
or U8015 (N_8015,N_82,N_693);
xor U8016 (N_8016,N_3646,N_3409);
and U8017 (N_8017,N_3155,N_403);
nor U8018 (N_8018,N_637,N_4833);
and U8019 (N_8019,N_1288,N_4736);
nor U8020 (N_8020,N_503,N_1201);
nand U8021 (N_8021,N_3289,N_222);
or U8022 (N_8022,N_2860,N_721);
and U8023 (N_8023,N_1660,N_3668);
xnor U8024 (N_8024,N_2509,N_4392);
xor U8025 (N_8025,N_3207,N_214);
and U8026 (N_8026,N_4977,N_908);
nand U8027 (N_8027,N_4417,N_1044);
and U8028 (N_8028,N_573,N_1593);
and U8029 (N_8029,N_1251,N_1602);
and U8030 (N_8030,N_3231,N_2664);
or U8031 (N_8031,N_4567,N_1558);
nor U8032 (N_8032,N_2330,N_3577);
or U8033 (N_8033,N_4911,N_3460);
nand U8034 (N_8034,N_556,N_1688);
or U8035 (N_8035,N_3450,N_2087);
nand U8036 (N_8036,N_2471,N_46);
nand U8037 (N_8037,N_1703,N_1513);
or U8038 (N_8038,N_3932,N_2877);
nand U8039 (N_8039,N_2907,N_2030);
xnor U8040 (N_8040,N_497,N_283);
and U8041 (N_8041,N_9,N_829);
and U8042 (N_8042,N_2594,N_859);
nor U8043 (N_8043,N_1505,N_1782);
nor U8044 (N_8044,N_4979,N_3092);
nand U8045 (N_8045,N_3460,N_2413);
or U8046 (N_8046,N_666,N_2153);
nor U8047 (N_8047,N_2429,N_363);
nor U8048 (N_8048,N_1959,N_2136);
xnor U8049 (N_8049,N_4766,N_2953);
xnor U8050 (N_8050,N_1274,N_1609);
and U8051 (N_8051,N_1,N_4516);
nand U8052 (N_8052,N_4292,N_2543);
and U8053 (N_8053,N_1339,N_967);
or U8054 (N_8054,N_4490,N_3639);
nor U8055 (N_8055,N_3115,N_1183);
and U8056 (N_8056,N_4770,N_3901);
or U8057 (N_8057,N_4323,N_3199);
xnor U8058 (N_8058,N_1039,N_3848);
nor U8059 (N_8059,N_4558,N_2520);
nand U8060 (N_8060,N_252,N_872);
xor U8061 (N_8061,N_1195,N_3171);
nand U8062 (N_8062,N_1754,N_322);
xnor U8063 (N_8063,N_4623,N_748);
or U8064 (N_8064,N_2480,N_327);
xor U8065 (N_8065,N_2673,N_3645);
or U8066 (N_8066,N_1499,N_1013);
nor U8067 (N_8067,N_3677,N_2966);
nand U8068 (N_8068,N_2062,N_978);
xnor U8069 (N_8069,N_1260,N_4581);
xor U8070 (N_8070,N_929,N_3585);
nand U8071 (N_8071,N_1886,N_2543);
nor U8072 (N_8072,N_387,N_4714);
xor U8073 (N_8073,N_4137,N_2684);
and U8074 (N_8074,N_3593,N_2339);
nor U8075 (N_8075,N_2909,N_4392);
nand U8076 (N_8076,N_3706,N_1949);
and U8077 (N_8077,N_614,N_1326);
xnor U8078 (N_8078,N_4668,N_4311);
nor U8079 (N_8079,N_1221,N_1668);
xor U8080 (N_8080,N_711,N_4787);
and U8081 (N_8081,N_4632,N_3372);
or U8082 (N_8082,N_4544,N_81);
and U8083 (N_8083,N_1976,N_3416);
nor U8084 (N_8084,N_4666,N_36);
nor U8085 (N_8085,N_2605,N_3468);
and U8086 (N_8086,N_598,N_2187);
nor U8087 (N_8087,N_4339,N_1188);
xor U8088 (N_8088,N_1744,N_581);
and U8089 (N_8089,N_884,N_4893);
and U8090 (N_8090,N_4411,N_4505);
xor U8091 (N_8091,N_2261,N_2527);
xor U8092 (N_8092,N_3573,N_1862);
nand U8093 (N_8093,N_2505,N_2227);
nor U8094 (N_8094,N_4319,N_2475);
and U8095 (N_8095,N_4942,N_2554);
nand U8096 (N_8096,N_1206,N_1565);
nand U8097 (N_8097,N_3414,N_3946);
nand U8098 (N_8098,N_1389,N_3159);
and U8099 (N_8099,N_3657,N_1232);
nand U8100 (N_8100,N_2656,N_3862);
or U8101 (N_8101,N_2331,N_2054);
or U8102 (N_8102,N_1565,N_2480);
or U8103 (N_8103,N_1860,N_336);
xnor U8104 (N_8104,N_1337,N_1733);
and U8105 (N_8105,N_4750,N_4807);
nand U8106 (N_8106,N_389,N_4486);
and U8107 (N_8107,N_1559,N_1403);
xor U8108 (N_8108,N_1688,N_3363);
and U8109 (N_8109,N_916,N_4915);
xor U8110 (N_8110,N_3468,N_4701);
and U8111 (N_8111,N_250,N_645);
xnor U8112 (N_8112,N_2732,N_1772);
nand U8113 (N_8113,N_658,N_3668);
or U8114 (N_8114,N_697,N_1169);
and U8115 (N_8115,N_1015,N_584);
nand U8116 (N_8116,N_3569,N_3473);
nand U8117 (N_8117,N_4231,N_1144);
or U8118 (N_8118,N_3469,N_2932);
or U8119 (N_8119,N_2444,N_777);
and U8120 (N_8120,N_227,N_3200);
and U8121 (N_8121,N_4110,N_1729);
and U8122 (N_8122,N_1510,N_3319);
nand U8123 (N_8123,N_1006,N_3126);
and U8124 (N_8124,N_2736,N_2473);
nand U8125 (N_8125,N_2002,N_0);
nand U8126 (N_8126,N_3602,N_4205);
nand U8127 (N_8127,N_3600,N_24);
or U8128 (N_8128,N_4678,N_3324);
nand U8129 (N_8129,N_1237,N_1478);
xor U8130 (N_8130,N_1220,N_3526);
nand U8131 (N_8131,N_4318,N_194);
nor U8132 (N_8132,N_3544,N_98);
xnor U8133 (N_8133,N_1500,N_358);
nand U8134 (N_8134,N_2431,N_49);
nor U8135 (N_8135,N_3879,N_526);
and U8136 (N_8136,N_3330,N_4319);
or U8137 (N_8137,N_2864,N_444);
xnor U8138 (N_8138,N_3894,N_2705);
xnor U8139 (N_8139,N_4698,N_26);
xor U8140 (N_8140,N_2732,N_3716);
or U8141 (N_8141,N_3659,N_2854);
and U8142 (N_8142,N_1655,N_3579);
or U8143 (N_8143,N_1789,N_1465);
nand U8144 (N_8144,N_2323,N_470);
nor U8145 (N_8145,N_4343,N_4629);
nand U8146 (N_8146,N_4956,N_1366);
nand U8147 (N_8147,N_3944,N_3645);
and U8148 (N_8148,N_192,N_1366);
xnor U8149 (N_8149,N_1363,N_615);
or U8150 (N_8150,N_1847,N_3458);
xor U8151 (N_8151,N_469,N_842);
and U8152 (N_8152,N_1457,N_3489);
or U8153 (N_8153,N_2655,N_2996);
xnor U8154 (N_8154,N_3909,N_455);
xor U8155 (N_8155,N_1801,N_4101);
nand U8156 (N_8156,N_2408,N_227);
or U8157 (N_8157,N_3686,N_2625);
and U8158 (N_8158,N_286,N_3687);
or U8159 (N_8159,N_2576,N_882);
and U8160 (N_8160,N_3631,N_1344);
nand U8161 (N_8161,N_3316,N_4006);
nand U8162 (N_8162,N_1209,N_3808);
nand U8163 (N_8163,N_2663,N_2248);
or U8164 (N_8164,N_1146,N_2758);
and U8165 (N_8165,N_1998,N_3042);
xor U8166 (N_8166,N_146,N_3408);
xnor U8167 (N_8167,N_1687,N_1155);
nor U8168 (N_8168,N_1787,N_2065);
nand U8169 (N_8169,N_3200,N_217);
or U8170 (N_8170,N_954,N_2443);
and U8171 (N_8171,N_4291,N_2945);
nand U8172 (N_8172,N_3274,N_892);
or U8173 (N_8173,N_3918,N_4588);
nor U8174 (N_8174,N_764,N_4556);
or U8175 (N_8175,N_2565,N_2398);
xor U8176 (N_8176,N_2180,N_780);
or U8177 (N_8177,N_1054,N_3973);
or U8178 (N_8178,N_2556,N_4312);
xnor U8179 (N_8179,N_4666,N_3308);
nor U8180 (N_8180,N_2001,N_3194);
or U8181 (N_8181,N_2696,N_1425);
xor U8182 (N_8182,N_2212,N_3308);
nor U8183 (N_8183,N_3871,N_3518);
and U8184 (N_8184,N_3469,N_4192);
nor U8185 (N_8185,N_3930,N_3451);
nand U8186 (N_8186,N_1088,N_4147);
or U8187 (N_8187,N_901,N_326);
xnor U8188 (N_8188,N_4743,N_3268);
nand U8189 (N_8189,N_4995,N_1589);
xnor U8190 (N_8190,N_915,N_463);
and U8191 (N_8191,N_3408,N_27);
or U8192 (N_8192,N_642,N_4959);
or U8193 (N_8193,N_4504,N_4008);
and U8194 (N_8194,N_4077,N_842);
or U8195 (N_8195,N_281,N_1297);
nor U8196 (N_8196,N_518,N_3439);
xnor U8197 (N_8197,N_1865,N_844);
or U8198 (N_8198,N_1055,N_1850);
xor U8199 (N_8199,N_3209,N_3362);
and U8200 (N_8200,N_3148,N_3259);
or U8201 (N_8201,N_2203,N_2368);
xnor U8202 (N_8202,N_3034,N_3448);
or U8203 (N_8203,N_4712,N_4902);
xnor U8204 (N_8204,N_2059,N_4914);
nor U8205 (N_8205,N_3424,N_439);
or U8206 (N_8206,N_3443,N_1823);
or U8207 (N_8207,N_423,N_500);
nor U8208 (N_8208,N_3742,N_3037);
or U8209 (N_8209,N_4633,N_2501);
and U8210 (N_8210,N_1202,N_4654);
or U8211 (N_8211,N_1812,N_1229);
nor U8212 (N_8212,N_562,N_1240);
nor U8213 (N_8213,N_3952,N_2982);
xnor U8214 (N_8214,N_1025,N_444);
nand U8215 (N_8215,N_990,N_4418);
nor U8216 (N_8216,N_3594,N_4622);
or U8217 (N_8217,N_1358,N_2561);
nor U8218 (N_8218,N_330,N_4455);
nand U8219 (N_8219,N_2133,N_955);
and U8220 (N_8220,N_3005,N_2834);
or U8221 (N_8221,N_1492,N_3792);
xor U8222 (N_8222,N_4051,N_3176);
nor U8223 (N_8223,N_884,N_2324);
nand U8224 (N_8224,N_1023,N_2769);
or U8225 (N_8225,N_970,N_1669);
xor U8226 (N_8226,N_1924,N_658);
or U8227 (N_8227,N_50,N_443);
xnor U8228 (N_8228,N_3357,N_1895);
nor U8229 (N_8229,N_4257,N_614);
xnor U8230 (N_8230,N_2289,N_140);
or U8231 (N_8231,N_340,N_1292);
xor U8232 (N_8232,N_2396,N_166);
or U8233 (N_8233,N_2782,N_4035);
xor U8234 (N_8234,N_371,N_2715);
xor U8235 (N_8235,N_229,N_2866);
or U8236 (N_8236,N_4336,N_1188);
nand U8237 (N_8237,N_4191,N_1299);
nor U8238 (N_8238,N_524,N_1461);
or U8239 (N_8239,N_1643,N_2806);
and U8240 (N_8240,N_650,N_1685);
nand U8241 (N_8241,N_759,N_208);
nand U8242 (N_8242,N_2886,N_3670);
nand U8243 (N_8243,N_3972,N_4323);
or U8244 (N_8244,N_3811,N_1669);
nor U8245 (N_8245,N_2052,N_483);
nand U8246 (N_8246,N_962,N_4874);
nand U8247 (N_8247,N_486,N_1375);
or U8248 (N_8248,N_2746,N_3367);
xor U8249 (N_8249,N_1078,N_4637);
nor U8250 (N_8250,N_1355,N_4586);
nor U8251 (N_8251,N_231,N_2135);
nor U8252 (N_8252,N_2177,N_3468);
and U8253 (N_8253,N_4004,N_2647);
xor U8254 (N_8254,N_292,N_3782);
xor U8255 (N_8255,N_859,N_4989);
xnor U8256 (N_8256,N_2829,N_3689);
and U8257 (N_8257,N_16,N_1322);
nand U8258 (N_8258,N_3071,N_2434);
nand U8259 (N_8259,N_461,N_2536);
or U8260 (N_8260,N_627,N_137);
nand U8261 (N_8261,N_2417,N_2336);
xnor U8262 (N_8262,N_4788,N_1486);
xnor U8263 (N_8263,N_4995,N_1388);
nand U8264 (N_8264,N_4768,N_1589);
nor U8265 (N_8265,N_4086,N_4297);
and U8266 (N_8266,N_336,N_4965);
or U8267 (N_8267,N_2556,N_1468);
nand U8268 (N_8268,N_2680,N_171);
or U8269 (N_8269,N_1223,N_2637);
nand U8270 (N_8270,N_333,N_1531);
nand U8271 (N_8271,N_2633,N_2250);
nand U8272 (N_8272,N_4879,N_2597);
and U8273 (N_8273,N_4850,N_1290);
nor U8274 (N_8274,N_4122,N_3984);
nand U8275 (N_8275,N_4862,N_3397);
or U8276 (N_8276,N_1747,N_35);
and U8277 (N_8277,N_3058,N_626);
nand U8278 (N_8278,N_2992,N_3926);
xor U8279 (N_8279,N_1527,N_201);
xnor U8280 (N_8280,N_1653,N_1542);
nand U8281 (N_8281,N_3601,N_4190);
and U8282 (N_8282,N_36,N_3710);
nor U8283 (N_8283,N_4847,N_3901);
and U8284 (N_8284,N_1298,N_1809);
xnor U8285 (N_8285,N_4134,N_955);
and U8286 (N_8286,N_2848,N_4748);
nand U8287 (N_8287,N_2663,N_1799);
nor U8288 (N_8288,N_3745,N_3837);
and U8289 (N_8289,N_872,N_2458);
xor U8290 (N_8290,N_3862,N_4214);
xnor U8291 (N_8291,N_4647,N_2247);
nand U8292 (N_8292,N_190,N_3416);
xnor U8293 (N_8293,N_4482,N_3279);
nand U8294 (N_8294,N_2536,N_377);
xnor U8295 (N_8295,N_4166,N_3708);
or U8296 (N_8296,N_4614,N_3211);
or U8297 (N_8297,N_4910,N_4851);
or U8298 (N_8298,N_3167,N_355);
nor U8299 (N_8299,N_3868,N_2048);
and U8300 (N_8300,N_4236,N_968);
nor U8301 (N_8301,N_2809,N_1292);
xor U8302 (N_8302,N_111,N_73);
nand U8303 (N_8303,N_4397,N_848);
xor U8304 (N_8304,N_3554,N_4017);
and U8305 (N_8305,N_2639,N_3925);
nand U8306 (N_8306,N_4544,N_3471);
nand U8307 (N_8307,N_3588,N_417);
nand U8308 (N_8308,N_2428,N_1509);
nand U8309 (N_8309,N_3232,N_3362);
and U8310 (N_8310,N_2707,N_4486);
nand U8311 (N_8311,N_4581,N_3135);
or U8312 (N_8312,N_3452,N_158);
xnor U8313 (N_8313,N_4671,N_4867);
nor U8314 (N_8314,N_3391,N_4435);
xor U8315 (N_8315,N_1934,N_1509);
nor U8316 (N_8316,N_4933,N_3294);
xor U8317 (N_8317,N_3007,N_2425);
xnor U8318 (N_8318,N_2171,N_3158);
and U8319 (N_8319,N_2219,N_4874);
nor U8320 (N_8320,N_930,N_842);
nor U8321 (N_8321,N_3052,N_4715);
xor U8322 (N_8322,N_2720,N_4734);
nand U8323 (N_8323,N_3600,N_1807);
xor U8324 (N_8324,N_1313,N_1202);
or U8325 (N_8325,N_887,N_4975);
or U8326 (N_8326,N_3497,N_1665);
and U8327 (N_8327,N_3783,N_1773);
nand U8328 (N_8328,N_2177,N_1805);
or U8329 (N_8329,N_1292,N_1877);
xor U8330 (N_8330,N_243,N_1580);
or U8331 (N_8331,N_1915,N_2535);
nand U8332 (N_8332,N_618,N_1665);
and U8333 (N_8333,N_3309,N_4589);
and U8334 (N_8334,N_1286,N_1363);
nor U8335 (N_8335,N_129,N_1686);
nor U8336 (N_8336,N_3726,N_4781);
nand U8337 (N_8337,N_1331,N_2882);
nand U8338 (N_8338,N_1105,N_1500);
nor U8339 (N_8339,N_2512,N_4335);
xor U8340 (N_8340,N_1356,N_3131);
or U8341 (N_8341,N_138,N_820);
nand U8342 (N_8342,N_4012,N_3129);
nor U8343 (N_8343,N_3200,N_815);
nand U8344 (N_8344,N_4084,N_867);
or U8345 (N_8345,N_1103,N_3767);
xnor U8346 (N_8346,N_3546,N_3714);
or U8347 (N_8347,N_4012,N_900);
or U8348 (N_8348,N_3108,N_4898);
nor U8349 (N_8349,N_2910,N_1938);
nor U8350 (N_8350,N_1895,N_2238);
or U8351 (N_8351,N_773,N_435);
and U8352 (N_8352,N_3029,N_494);
and U8353 (N_8353,N_1678,N_4202);
nor U8354 (N_8354,N_4459,N_3853);
or U8355 (N_8355,N_4706,N_2392);
xor U8356 (N_8356,N_3396,N_529);
xnor U8357 (N_8357,N_2222,N_1908);
nand U8358 (N_8358,N_2359,N_1443);
or U8359 (N_8359,N_150,N_1962);
or U8360 (N_8360,N_1451,N_3494);
nor U8361 (N_8361,N_4207,N_87);
or U8362 (N_8362,N_2316,N_4250);
nand U8363 (N_8363,N_4804,N_3677);
nand U8364 (N_8364,N_2402,N_388);
xor U8365 (N_8365,N_2498,N_4118);
xor U8366 (N_8366,N_3715,N_970);
or U8367 (N_8367,N_4880,N_4638);
nor U8368 (N_8368,N_1372,N_4036);
xor U8369 (N_8369,N_3205,N_3812);
nor U8370 (N_8370,N_2771,N_2102);
nor U8371 (N_8371,N_2153,N_170);
nor U8372 (N_8372,N_3077,N_3517);
or U8373 (N_8373,N_2005,N_242);
nor U8374 (N_8374,N_4790,N_2763);
nand U8375 (N_8375,N_3222,N_4460);
and U8376 (N_8376,N_1872,N_232);
or U8377 (N_8377,N_4994,N_322);
and U8378 (N_8378,N_2234,N_2962);
or U8379 (N_8379,N_4714,N_2401);
or U8380 (N_8380,N_2184,N_2651);
or U8381 (N_8381,N_2957,N_3856);
xnor U8382 (N_8382,N_1638,N_2411);
nand U8383 (N_8383,N_2092,N_3451);
nor U8384 (N_8384,N_4542,N_133);
xnor U8385 (N_8385,N_941,N_426);
and U8386 (N_8386,N_3153,N_2949);
nand U8387 (N_8387,N_3444,N_418);
nor U8388 (N_8388,N_2821,N_2437);
or U8389 (N_8389,N_3201,N_4496);
and U8390 (N_8390,N_1545,N_1994);
and U8391 (N_8391,N_1330,N_1376);
nor U8392 (N_8392,N_1451,N_2019);
and U8393 (N_8393,N_69,N_2698);
and U8394 (N_8394,N_502,N_277);
xnor U8395 (N_8395,N_999,N_3595);
nand U8396 (N_8396,N_1821,N_1474);
and U8397 (N_8397,N_4226,N_838);
or U8398 (N_8398,N_1541,N_3683);
xnor U8399 (N_8399,N_2621,N_1780);
and U8400 (N_8400,N_2330,N_3283);
xnor U8401 (N_8401,N_2571,N_4037);
nor U8402 (N_8402,N_2716,N_720);
nand U8403 (N_8403,N_4248,N_241);
or U8404 (N_8404,N_1876,N_2976);
or U8405 (N_8405,N_3009,N_2741);
and U8406 (N_8406,N_4418,N_2115);
or U8407 (N_8407,N_4116,N_1391);
or U8408 (N_8408,N_882,N_3567);
xor U8409 (N_8409,N_3517,N_4021);
nand U8410 (N_8410,N_894,N_4095);
nand U8411 (N_8411,N_1973,N_1977);
or U8412 (N_8412,N_1638,N_2888);
or U8413 (N_8413,N_2012,N_2041);
xnor U8414 (N_8414,N_2733,N_4177);
nand U8415 (N_8415,N_1088,N_3548);
and U8416 (N_8416,N_2801,N_4661);
nand U8417 (N_8417,N_4776,N_3432);
nor U8418 (N_8418,N_348,N_1941);
xnor U8419 (N_8419,N_2169,N_4202);
xor U8420 (N_8420,N_433,N_4342);
nand U8421 (N_8421,N_3621,N_2349);
xor U8422 (N_8422,N_4537,N_2238);
or U8423 (N_8423,N_612,N_3407);
nand U8424 (N_8424,N_4443,N_4170);
nor U8425 (N_8425,N_3754,N_1145);
xnor U8426 (N_8426,N_1010,N_1963);
xnor U8427 (N_8427,N_3765,N_4824);
nor U8428 (N_8428,N_4751,N_4034);
xnor U8429 (N_8429,N_2573,N_1229);
or U8430 (N_8430,N_3159,N_4384);
and U8431 (N_8431,N_2476,N_3114);
nor U8432 (N_8432,N_1154,N_869);
xnor U8433 (N_8433,N_1891,N_3415);
xnor U8434 (N_8434,N_1914,N_3135);
nor U8435 (N_8435,N_2897,N_397);
xor U8436 (N_8436,N_4333,N_1142);
or U8437 (N_8437,N_402,N_915);
and U8438 (N_8438,N_1246,N_3243);
nand U8439 (N_8439,N_2432,N_3270);
and U8440 (N_8440,N_3268,N_1050);
xor U8441 (N_8441,N_773,N_376);
and U8442 (N_8442,N_86,N_1727);
nand U8443 (N_8443,N_4635,N_636);
xor U8444 (N_8444,N_1176,N_4188);
nor U8445 (N_8445,N_1230,N_3114);
or U8446 (N_8446,N_185,N_1445);
nand U8447 (N_8447,N_787,N_1405);
nor U8448 (N_8448,N_1649,N_2952);
xnor U8449 (N_8449,N_598,N_3876);
xor U8450 (N_8450,N_3134,N_2330);
or U8451 (N_8451,N_2359,N_4635);
nand U8452 (N_8452,N_2206,N_4649);
and U8453 (N_8453,N_64,N_3200);
nor U8454 (N_8454,N_1847,N_4391);
nand U8455 (N_8455,N_3041,N_3106);
xnor U8456 (N_8456,N_3972,N_2416);
nor U8457 (N_8457,N_2640,N_4422);
and U8458 (N_8458,N_1758,N_2324);
and U8459 (N_8459,N_1870,N_2333);
nor U8460 (N_8460,N_3861,N_1375);
and U8461 (N_8461,N_2587,N_4885);
nand U8462 (N_8462,N_4048,N_1801);
nor U8463 (N_8463,N_4405,N_1907);
xor U8464 (N_8464,N_1064,N_1111);
and U8465 (N_8465,N_3264,N_1902);
or U8466 (N_8466,N_2546,N_2610);
or U8467 (N_8467,N_2943,N_1033);
nor U8468 (N_8468,N_1734,N_1285);
or U8469 (N_8469,N_281,N_1068);
xnor U8470 (N_8470,N_986,N_2630);
xor U8471 (N_8471,N_653,N_4234);
xnor U8472 (N_8472,N_1393,N_62);
or U8473 (N_8473,N_1619,N_3065);
nand U8474 (N_8474,N_2443,N_730);
xnor U8475 (N_8475,N_4118,N_2399);
nand U8476 (N_8476,N_3143,N_42);
nor U8477 (N_8477,N_309,N_1238);
and U8478 (N_8478,N_2447,N_2601);
xnor U8479 (N_8479,N_3856,N_1159);
xor U8480 (N_8480,N_4411,N_4788);
nand U8481 (N_8481,N_2603,N_1446);
or U8482 (N_8482,N_3787,N_3211);
nand U8483 (N_8483,N_4104,N_3944);
or U8484 (N_8484,N_1932,N_4681);
nor U8485 (N_8485,N_3421,N_1940);
nor U8486 (N_8486,N_2467,N_3488);
or U8487 (N_8487,N_3508,N_2175);
and U8488 (N_8488,N_2834,N_2077);
or U8489 (N_8489,N_4666,N_682);
nand U8490 (N_8490,N_3689,N_4096);
and U8491 (N_8491,N_1051,N_2575);
and U8492 (N_8492,N_2848,N_2722);
nand U8493 (N_8493,N_3271,N_4482);
xnor U8494 (N_8494,N_3094,N_2879);
nand U8495 (N_8495,N_817,N_4937);
and U8496 (N_8496,N_4201,N_3319);
and U8497 (N_8497,N_1595,N_3049);
or U8498 (N_8498,N_1076,N_4419);
xnor U8499 (N_8499,N_46,N_4661);
nor U8500 (N_8500,N_4088,N_624);
or U8501 (N_8501,N_1182,N_4865);
or U8502 (N_8502,N_3,N_4396);
or U8503 (N_8503,N_4943,N_1590);
nor U8504 (N_8504,N_1052,N_693);
nor U8505 (N_8505,N_3178,N_2190);
nand U8506 (N_8506,N_3795,N_462);
and U8507 (N_8507,N_140,N_2278);
xnor U8508 (N_8508,N_1642,N_1270);
nand U8509 (N_8509,N_3798,N_3623);
xnor U8510 (N_8510,N_2109,N_4474);
or U8511 (N_8511,N_1835,N_1515);
nand U8512 (N_8512,N_4840,N_945);
xor U8513 (N_8513,N_580,N_3362);
and U8514 (N_8514,N_4106,N_2655);
or U8515 (N_8515,N_572,N_4548);
and U8516 (N_8516,N_1598,N_1877);
or U8517 (N_8517,N_425,N_387);
nand U8518 (N_8518,N_1560,N_2660);
xnor U8519 (N_8519,N_2925,N_2733);
or U8520 (N_8520,N_2129,N_830);
or U8521 (N_8521,N_457,N_1382);
nand U8522 (N_8522,N_1669,N_4787);
or U8523 (N_8523,N_4200,N_4420);
and U8524 (N_8524,N_3693,N_3537);
or U8525 (N_8525,N_4951,N_3245);
and U8526 (N_8526,N_4362,N_2415);
nand U8527 (N_8527,N_3277,N_3156);
nor U8528 (N_8528,N_4760,N_2051);
and U8529 (N_8529,N_3714,N_2800);
and U8530 (N_8530,N_4926,N_3080);
xnor U8531 (N_8531,N_2901,N_618);
and U8532 (N_8532,N_1895,N_1609);
nor U8533 (N_8533,N_955,N_504);
xor U8534 (N_8534,N_1268,N_2300);
nor U8535 (N_8535,N_4407,N_3139);
or U8536 (N_8536,N_3039,N_506);
nor U8537 (N_8537,N_2047,N_3930);
or U8538 (N_8538,N_709,N_3305);
or U8539 (N_8539,N_1308,N_3954);
or U8540 (N_8540,N_2913,N_3627);
or U8541 (N_8541,N_1687,N_2909);
or U8542 (N_8542,N_1794,N_4623);
nand U8543 (N_8543,N_1098,N_3096);
xor U8544 (N_8544,N_1036,N_4497);
or U8545 (N_8545,N_1084,N_2802);
nor U8546 (N_8546,N_2015,N_971);
or U8547 (N_8547,N_3444,N_767);
nor U8548 (N_8548,N_985,N_835);
or U8549 (N_8549,N_1612,N_4029);
nand U8550 (N_8550,N_2252,N_2498);
nor U8551 (N_8551,N_3503,N_1593);
or U8552 (N_8552,N_3895,N_3204);
xor U8553 (N_8553,N_4410,N_4289);
and U8554 (N_8554,N_96,N_433);
nand U8555 (N_8555,N_231,N_567);
nor U8556 (N_8556,N_4740,N_3168);
nor U8557 (N_8557,N_289,N_505);
nor U8558 (N_8558,N_1854,N_4918);
xnor U8559 (N_8559,N_1163,N_3733);
xnor U8560 (N_8560,N_2926,N_3718);
nand U8561 (N_8561,N_1529,N_1809);
nor U8562 (N_8562,N_2453,N_1748);
nand U8563 (N_8563,N_3377,N_3532);
nand U8564 (N_8564,N_4526,N_2824);
xor U8565 (N_8565,N_4544,N_4255);
nand U8566 (N_8566,N_535,N_3830);
nor U8567 (N_8567,N_1563,N_1727);
or U8568 (N_8568,N_4155,N_4352);
and U8569 (N_8569,N_3603,N_2722);
or U8570 (N_8570,N_343,N_3025);
and U8571 (N_8571,N_3581,N_3145);
nand U8572 (N_8572,N_4751,N_2762);
nand U8573 (N_8573,N_446,N_3983);
and U8574 (N_8574,N_449,N_4158);
or U8575 (N_8575,N_522,N_3436);
nand U8576 (N_8576,N_4005,N_1350);
nand U8577 (N_8577,N_3577,N_105);
nor U8578 (N_8578,N_1510,N_3071);
or U8579 (N_8579,N_2079,N_1348);
nor U8580 (N_8580,N_2408,N_2032);
and U8581 (N_8581,N_3784,N_42);
or U8582 (N_8582,N_1640,N_3044);
xor U8583 (N_8583,N_1286,N_207);
and U8584 (N_8584,N_3141,N_4644);
and U8585 (N_8585,N_1484,N_3781);
nand U8586 (N_8586,N_4487,N_4657);
or U8587 (N_8587,N_183,N_4984);
nand U8588 (N_8588,N_236,N_2785);
xnor U8589 (N_8589,N_3212,N_276);
and U8590 (N_8590,N_1387,N_74);
and U8591 (N_8591,N_1022,N_1241);
or U8592 (N_8592,N_2402,N_3655);
xnor U8593 (N_8593,N_2612,N_4405);
nand U8594 (N_8594,N_481,N_776);
and U8595 (N_8595,N_3224,N_3518);
and U8596 (N_8596,N_4893,N_216);
xor U8597 (N_8597,N_3648,N_3105);
or U8598 (N_8598,N_1429,N_219);
and U8599 (N_8599,N_2274,N_765);
or U8600 (N_8600,N_4920,N_3262);
xnor U8601 (N_8601,N_2711,N_2932);
and U8602 (N_8602,N_2416,N_3228);
and U8603 (N_8603,N_1884,N_2444);
nand U8604 (N_8604,N_4190,N_645);
xor U8605 (N_8605,N_3295,N_499);
or U8606 (N_8606,N_2671,N_3405);
nand U8607 (N_8607,N_725,N_817);
and U8608 (N_8608,N_360,N_1135);
nand U8609 (N_8609,N_3166,N_3980);
and U8610 (N_8610,N_800,N_1422);
or U8611 (N_8611,N_3622,N_1605);
or U8612 (N_8612,N_4833,N_3643);
xor U8613 (N_8613,N_3972,N_2531);
nand U8614 (N_8614,N_1196,N_2656);
nand U8615 (N_8615,N_3723,N_1225);
nor U8616 (N_8616,N_3602,N_3185);
and U8617 (N_8617,N_2487,N_4818);
nand U8618 (N_8618,N_4399,N_1742);
xor U8619 (N_8619,N_4841,N_4674);
nand U8620 (N_8620,N_4274,N_18);
nand U8621 (N_8621,N_4996,N_1866);
and U8622 (N_8622,N_2415,N_3287);
nand U8623 (N_8623,N_3962,N_893);
xor U8624 (N_8624,N_2448,N_845);
nand U8625 (N_8625,N_4076,N_381);
xor U8626 (N_8626,N_4978,N_3416);
or U8627 (N_8627,N_3296,N_1764);
or U8628 (N_8628,N_728,N_966);
nor U8629 (N_8629,N_3198,N_4649);
nand U8630 (N_8630,N_2666,N_4496);
nor U8631 (N_8631,N_1693,N_2520);
or U8632 (N_8632,N_3449,N_3725);
xor U8633 (N_8633,N_3096,N_3746);
xor U8634 (N_8634,N_1091,N_1067);
and U8635 (N_8635,N_2934,N_1974);
xnor U8636 (N_8636,N_4146,N_2262);
or U8637 (N_8637,N_4488,N_1813);
or U8638 (N_8638,N_110,N_463);
nand U8639 (N_8639,N_4920,N_1322);
nand U8640 (N_8640,N_114,N_2725);
nand U8641 (N_8641,N_1579,N_2943);
xor U8642 (N_8642,N_1962,N_4759);
nand U8643 (N_8643,N_4385,N_1019);
xnor U8644 (N_8644,N_732,N_719);
xnor U8645 (N_8645,N_4377,N_841);
and U8646 (N_8646,N_54,N_1079);
and U8647 (N_8647,N_3310,N_3269);
nor U8648 (N_8648,N_479,N_3567);
nand U8649 (N_8649,N_3610,N_11);
xnor U8650 (N_8650,N_1930,N_2646);
nor U8651 (N_8651,N_2236,N_67);
or U8652 (N_8652,N_362,N_4600);
nand U8653 (N_8653,N_1085,N_3623);
nand U8654 (N_8654,N_3151,N_79);
nor U8655 (N_8655,N_3009,N_3388);
nor U8656 (N_8656,N_4400,N_1387);
and U8657 (N_8657,N_2983,N_1544);
and U8658 (N_8658,N_4048,N_1032);
nand U8659 (N_8659,N_1984,N_3571);
or U8660 (N_8660,N_4935,N_1058);
nor U8661 (N_8661,N_3748,N_1464);
nor U8662 (N_8662,N_1031,N_280);
nand U8663 (N_8663,N_770,N_4683);
nand U8664 (N_8664,N_3960,N_2071);
or U8665 (N_8665,N_3156,N_2300);
nand U8666 (N_8666,N_1064,N_1740);
and U8667 (N_8667,N_2886,N_1998);
nand U8668 (N_8668,N_2965,N_1712);
nand U8669 (N_8669,N_4195,N_4264);
and U8670 (N_8670,N_3786,N_1933);
xnor U8671 (N_8671,N_3000,N_76);
or U8672 (N_8672,N_2776,N_645);
or U8673 (N_8673,N_4656,N_1679);
nand U8674 (N_8674,N_2437,N_4511);
xor U8675 (N_8675,N_4831,N_2758);
nor U8676 (N_8676,N_4021,N_4323);
nand U8677 (N_8677,N_3153,N_4122);
nand U8678 (N_8678,N_470,N_1218);
and U8679 (N_8679,N_3860,N_355);
nand U8680 (N_8680,N_4661,N_535);
nor U8681 (N_8681,N_4921,N_2556);
nand U8682 (N_8682,N_306,N_4752);
nor U8683 (N_8683,N_3883,N_4659);
nor U8684 (N_8684,N_3143,N_4990);
nor U8685 (N_8685,N_3255,N_4149);
xnor U8686 (N_8686,N_221,N_1143);
xor U8687 (N_8687,N_1464,N_3722);
xor U8688 (N_8688,N_1190,N_1709);
and U8689 (N_8689,N_3218,N_2873);
or U8690 (N_8690,N_3114,N_3141);
and U8691 (N_8691,N_3301,N_4113);
xor U8692 (N_8692,N_173,N_1197);
nor U8693 (N_8693,N_3880,N_3894);
nand U8694 (N_8694,N_820,N_2553);
or U8695 (N_8695,N_3440,N_773);
or U8696 (N_8696,N_1506,N_1961);
nor U8697 (N_8697,N_1980,N_2207);
nand U8698 (N_8698,N_4248,N_4754);
or U8699 (N_8699,N_4425,N_2743);
nor U8700 (N_8700,N_1708,N_883);
nand U8701 (N_8701,N_2669,N_1577);
and U8702 (N_8702,N_906,N_3411);
nand U8703 (N_8703,N_4040,N_1727);
nand U8704 (N_8704,N_4708,N_3143);
nand U8705 (N_8705,N_3192,N_3397);
xor U8706 (N_8706,N_3318,N_4637);
xor U8707 (N_8707,N_343,N_2821);
and U8708 (N_8708,N_2506,N_1460);
or U8709 (N_8709,N_2622,N_2279);
and U8710 (N_8710,N_4621,N_2747);
nand U8711 (N_8711,N_1821,N_2542);
nand U8712 (N_8712,N_1636,N_3076);
xnor U8713 (N_8713,N_2196,N_540);
xnor U8714 (N_8714,N_1749,N_2000);
nor U8715 (N_8715,N_2301,N_2906);
nand U8716 (N_8716,N_1205,N_535);
or U8717 (N_8717,N_2308,N_153);
and U8718 (N_8718,N_4083,N_4091);
xor U8719 (N_8719,N_2783,N_3725);
and U8720 (N_8720,N_3593,N_788);
nand U8721 (N_8721,N_1374,N_3691);
xnor U8722 (N_8722,N_3229,N_542);
xor U8723 (N_8723,N_3364,N_4003);
xor U8724 (N_8724,N_4320,N_3326);
xor U8725 (N_8725,N_534,N_2496);
xor U8726 (N_8726,N_2907,N_1270);
or U8727 (N_8727,N_3731,N_13);
nor U8728 (N_8728,N_3975,N_1660);
nor U8729 (N_8729,N_3410,N_828);
and U8730 (N_8730,N_1513,N_3876);
xnor U8731 (N_8731,N_4140,N_1165);
and U8732 (N_8732,N_4242,N_1409);
xnor U8733 (N_8733,N_2421,N_445);
and U8734 (N_8734,N_2899,N_3771);
nor U8735 (N_8735,N_3265,N_4079);
nor U8736 (N_8736,N_2425,N_211);
or U8737 (N_8737,N_3783,N_1766);
nand U8738 (N_8738,N_3746,N_3460);
nand U8739 (N_8739,N_3815,N_3319);
and U8740 (N_8740,N_662,N_2596);
xnor U8741 (N_8741,N_4246,N_4203);
xor U8742 (N_8742,N_3198,N_4433);
or U8743 (N_8743,N_3685,N_3341);
xnor U8744 (N_8744,N_1095,N_4983);
nor U8745 (N_8745,N_188,N_2837);
or U8746 (N_8746,N_4689,N_1754);
and U8747 (N_8747,N_4351,N_1412);
and U8748 (N_8748,N_2502,N_3877);
and U8749 (N_8749,N_783,N_525);
nor U8750 (N_8750,N_1575,N_4258);
nor U8751 (N_8751,N_3821,N_896);
nor U8752 (N_8752,N_827,N_1743);
nor U8753 (N_8753,N_449,N_1877);
or U8754 (N_8754,N_4948,N_801);
nor U8755 (N_8755,N_4981,N_4552);
or U8756 (N_8756,N_3259,N_864);
nor U8757 (N_8757,N_3951,N_1120);
nand U8758 (N_8758,N_4721,N_489);
nor U8759 (N_8759,N_2406,N_1260);
nor U8760 (N_8760,N_3889,N_2952);
xor U8761 (N_8761,N_3479,N_2379);
or U8762 (N_8762,N_1617,N_3541);
and U8763 (N_8763,N_1745,N_1570);
or U8764 (N_8764,N_1845,N_1032);
and U8765 (N_8765,N_4466,N_3944);
nor U8766 (N_8766,N_1655,N_1982);
xor U8767 (N_8767,N_1517,N_2361);
or U8768 (N_8768,N_1103,N_2342);
nand U8769 (N_8769,N_4464,N_503);
and U8770 (N_8770,N_4452,N_1194);
nor U8771 (N_8771,N_2537,N_911);
nor U8772 (N_8772,N_3048,N_1538);
or U8773 (N_8773,N_4664,N_2401);
nor U8774 (N_8774,N_3576,N_3032);
or U8775 (N_8775,N_692,N_3391);
nand U8776 (N_8776,N_1574,N_192);
nand U8777 (N_8777,N_340,N_538);
xor U8778 (N_8778,N_4668,N_121);
or U8779 (N_8779,N_2104,N_1023);
and U8780 (N_8780,N_4958,N_4620);
nor U8781 (N_8781,N_2671,N_3707);
and U8782 (N_8782,N_1978,N_2796);
or U8783 (N_8783,N_1252,N_3442);
xnor U8784 (N_8784,N_4588,N_4000);
or U8785 (N_8785,N_2593,N_4598);
xnor U8786 (N_8786,N_3308,N_4358);
xnor U8787 (N_8787,N_4747,N_2423);
nand U8788 (N_8788,N_1548,N_330);
nor U8789 (N_8789,N_1838,N_3065);
or U8790 (N_8790,N_3005,N_2258);
and U8791 (N_8791,N_2680,N_3570);
nor U8792 (N_8792,N_1117,N_1129);
nand U8793 (N_8793,N_3310,N_2142);
xor U8794 (N_8794,N_1561,N_3758);
and U8795 (N_8795,N_447,N_2852);
and U8796 (N_8796,N_400,N_304);
and U8797 (N_8797,N_2790,N_4373);
and U8798 (N_8798,N_2964,N_3327);
and U8799 (N_8799,N_1040,N_4548);
and U8800 (N_8800,N_3010,N_29);
nand U8801 (N_8801,N_2480,N_2291);
xor U8802 (N_8802,N_1628,N_26);
and U8803 (N_8803,N_2202,N_3315);
nand U8804 (N_8804,N_2509,N_2954);
xor U8805 (N_8805,N_2276,N_1491);
and U8806 (N_8806,N_1747,N_739);
xnor U8807 (N_8807,N_333,N_4129);
nor U8808 (N_8808,N_231,N_2303);
xor U8809 (N_8809,N_2378,N_1826);
nand U8810 (N_8810,N_2280,N_2423);
nand U8811 (N_8811,N_1507,N_3408);
or U8812 (N_8812,N_2159,N_2770);
or U8813 (N_8813,N_4454,N_1544);
nor U8814 (N_8814,N_4363,N_3305);
nand U8815 (N_8815,N_120,N_4476);
and U8816 (N_8816,N_1415,N_3572);
nand U8817 (N_8817,N_3449,N_4077);
and U8818 (N_8818,N_1104,N_1479);
and U8819 (N_8819,N_651,N_1405);
and U8820 (N_8820,N_4389,N_4511);
or U8821 (N_8821,N_2743,N_2104);
and U8822 (N_8822,N_3896,N_2810);
and U8823 (N_8823,N_1879,N_3765);
or U8824 (N_8824,N_1774,N_3394);
or U8825 (N_8825,N_2746,N_2450);
xnor U8826 (N_8826,N_1635,N_4676);
xnor U8827 (N_8827,N_1978,N_575);
or U8828 (N_8828,N_1654,N_2793);
nand U8829 (N_8829,N_3587,N_3804);
nor U8830 (N_8830,N_1275,N_2906);
or U8831 (N_8831,N_2231,N_2947);
and U8832 (N_8832,N_3028,N_2454);
nor U8833 (N_8833,N_718,N_3413);
xor U8834 (N_8834,N_2787,N_2487);
nor U8835 (N_8835,N_247,N_4429);
and U8836 (N_8836,N_444,N_4893);
or U8837 (N_8837,N_2473,N_4497);
nand U8838 (N_8838,N_3912,N_4511);
xnor U8839 (N_8839,N_2443,N_1938);
nand U8840 (N_8840,N_4897,N_1371);
and U8841 (N_8841,N_2915,N_3924);
nand U8842 (N_8842,N_4286,N_2675);
xnor U8843 (N_8843,N_2705,N_1940);
nor U8844 (N_8844,N_748,N_1500);
xor U8845 (N_8845,N_1689,N_17);
nand U8846 (N_8846,N_2445,N_1326);
or U8847 (N_8847,N_1922,N_4954);
nand U8848 (N_8848,N_4660,N_2547);
nor U8849 (N_8849,N_1987,N_2176);
and U8850 (N_8850,N_4412,N_2210);
nand U8851 (N_8851,N_3956,N_243);
nor U8852 (N_8852,N_3748,N_1403);
xnor U8853 (N_8853,N_1363,N_2570);
and U8854 (N_8854,N_1179,N_4414);
and U8855 (N_8855,N_1957,N_3433);
xnor U8856 (N_8856,N_3174,N_709);
xor U8857 (N_8857,N_2770,N_26);
nor U8858 (N_8858,N_3128,N_132);
nand U8859 (N_8859,N_99,N_4456);
xnor U8860 (N_8860,N_2020,N_4750);
or U8861 (N_8861,N_1673,N_679);
or U8862 (N_8862,N_4140,N_2053);
xor U8863 (N_8863,N_4954,N_937);
and U8864 (N_8864,N_3090,N_1701);
and U8865 (N_8865,N_1637,N_3467);
nor U8866 (N_8866,N_1196,N_766);
nand U8867 (N_8867,N_4643,N_3374);
and U8868 (N_8868,N_4340,N_3142);
nand U8869 (N_8869,N_4588,N_3902);
nor U8870 (N_8870,N_4487,N_2178);
and U8871 (N_8871,N_569,N_4752);
or U8872 (N_8872,N_1217,N_4638);
nor U8873 (N_8873,N_2187,N_1282);
or U8874 (N_8874,N_2004,N_3619);
nor U8875 (N_8875,N_4026,N_4318);
nand U8876 (N_8876,N_3584,N_2410);
or U8877 (N_8877,N_2647,N_2301);
and U8878 (N_8878,N_1725,N_1512);
nand U8879 (N_8879,N_1435,N_609);
nand U8880 (N_8880,N_2666,N_3765);
and U8881 (N_8881,N_527,N_347);
or U8882 (N_8882,N_2613,N_3939);
and U8883 (N_8883,N_1880,N_657);
and U8884 (N_8884,N_1015,N_2337);
or U8885 (N_8885,N_166,N_3997);
nand U8886 (N_8886,N_3108,N_619);
xnor U8887 (N_8887,N_220,N_1401);
or U8888 (N_8888,N_1966,N_585);
xor U8889 (N_8889,N_4348,N_4024);
nand U8890 (N_8890,N_2412,N_2739);
and U8891 (N_8891,N_94,N_4521);
and U8892 (N_8892,N_1700,N_3945);
nor U8893 (N_8893,N_2859,N_4283);
and U8894 (N_8894,N_2554,N_685);
nand U8895 (N_8895,N_109,N_3707);
nor U8896 (N_8896,N_2531,N_4744);
and U8897 (N_8897,N_4117,N_4979);
or U8898 (N_8898,N_564,N_3293);
xnor U8899 (N_8899,N_2194,N_1412);
and U8900 (N_8900,N_472,N_1222);
nor U8901 (N_8901,N_682,N_314);
nand U8902 (N_8902,N_2139,N_4524);
or U8903 (N_8903,N_603,N_737);
and U8904 (N_8904,N_35,N_4987);
or U8905 (N_8905,N_354,N_4729);
or U8906 (N_8906,N_2011,N_179);
xnor U8907 (N_8907,N_4872,N_4958);
or U8908 (N_8908,N_4617,N_2444);
nor U8909 (N_8909,N_391,N_3194);
and U8910 (N_8910,N_4230,N_3607);
or U8911 (N_8911,N_1122,N_1509);
and U8912 (N_8912,N_2147,N_925);
nand U8913 (N_8913,N_3169,N_326);
xnor U8914 (N_8914,N_2506,N_2890);
or U8915 (N_8915,N_630,N_1129);
nand U8916 (N_8916,N_3361,N_3006);
and U8917 (N_8917,N_2420,N_501);
nor U8918 (N_8918,N_4973,N_3113);
nand U8919 (N_8919,N_112,N_2702);
and U8920 (N_8920,N_4429,N_2251);
and U8921 (N_8921,N_4911,N_2969);
or U8922 (N_8922,N_184,N_1975);
or U8923 (N_8923,N_509,N_1831);
nand U8924 (N_8924,N_1322,N_112);
nand U8925 (N_8925,N_1307,N_373);
and U8926 (N_8926,N_3584,N_3424);
nor U8927 (N_8927,N_2866,N_589);
xnor U8928 (N_8928,N_659,N_2926);
and U8929 (N_8929,N_791,N_1785);
nand U8930 (N_8930,N_582,N_2355);
and U8931 (N_8931,N_302,N_2235);
xor U8932 (N_8932,N_976,N_2138);
nor U8933 (N_8933,N_778,N_2869);
xnor U8934 (N_8934,N_3937,N_3525);
or U8935 (N_8935,N_2424,N_2671);
or U8936 (N_8936,N_3954,N_3134);
and U8937 (N_8937,N_2004,N_339);
or U8938 (N_8938,N_694,N_3648);
or U8939 (N_8939,N_2096,N_3800);
and U8940 (N_8940,N_682,N_3758);
nor U8941 (N_8941,N_218,N_2598);
nand U8942 (N_8942,N_4943,N_4977);
nand U8943 (N_8943,N_656,N_2863);
nand U8944 (N_8944,N_1841,N_3639);
xor U8945 (N_8945,N_2881,N_2665);
xnor U8946 (N_8946,N_1407,N_1357);
or U8947 (N_8947,N_4699,N_2975);
and U8948 (N_8948,N_2778,N_2339);
xor U8949 (N_8949,N_1841,N_531);
and U8950 (N_8950,N_1769,N_3174);
nor U8951 (N_8951,N_1526,N_986);
xor U8952 (N_8952,N_4274,N_2941);
nand U8953 (N_8953,N_1716,N_4410);
xnor U8954 (N_8954,N_3584,N_2461);
and U8955 (N_8955,N_18,N_1689);
or U8956 (N_8956,N_1207,N_488);
and U8957 (N_8957,N_1610,N_1614);
and U8958 (N_8958,N_4612,N_694);
and U8959 (N_8959,N_4068,N_3701);
nand U8960 (N_8960,N_1053,N_376);
xnor U8961 (N_8961,N_1765,N_4164);
or U8962 (N_8962,N_249,N_1584);
or U8963 (N_8963,N_1296,N_2199);
or U8964 (N_8964,N_2612,N_2633);
nor U8965 (N_8965,N_2034,N_3327);
and U8966 (N_8966,N_1484,N_1430);
xnor U8967 (N_8967,N_3427,N_4053);
xor U8968 (N_8968,N_2739,N_4008);
or U8969 (N_8969,N_594,N_4953);
and U8970 (N_8970,N_470,N_2148);
and U8971 (N_8971,N_278,N_1372);
or U8972 (N_8972,N_2617,N_468);
nand U8973 (N_8973,N_1688,N_961);
nor U8974 (N_8974,N_1617,N_412);
nand U8975 (N_8975,N_839,N_4608);
xnor U8976 (N_8976,N_4459,N_1346);
and U8977 (N_8977,N_4949,N_3568);
nor U8978 (N_8978,N_2393,N_1913);
or U8979 (N_8979,N_598,N_4541);
xor U8980 (N_8980,N_656,N_3973);
and U8981 (N_8981,N_1876,N_4473);
xor U8982 (N_8982,N_677,N_1786);
nor U8983 (N_8983,N_3605,N_2431);
xor U8984 (N_8984,N_3763,N_2343);
or U8985 (N_8985,N_953,N_2110);
or U8986 (N_8986,N_2493,N_4444);
nand U8987 (N_8987,N_4372,N_2642);
nand U8988 (N_8988,N_3167,N_893);
or U8989 (N_8989,N_4814,N_2353);
nor U8990 (N_8990,N_4617,N_610);
and U8991 (N_8991,N_1453,N_495);
nand U8992 (N_8992,N_4027,N_2749);
nand U8993 (N_8993,N_1983,N_4711);
nor U8994 (N_8994,N_3726,N_4452);
xor U8995 (N_8995,N_1901,N_3320);
nand U8996 (N_8996,N_4160,N_535);
nor U8997 (N_8997,N_847,N_450);
xnor U8998 (N_8998,N_1642,N_250);
or U8999 (N_8999,N_4283,N_596);
nor U9000 (N_9000,N_2004,N_5);
xor U9001 (N_9001,N_4006,N_2261);
and U9002 (N_9002,N_2617,N_4246);
xnor U9003 (N_9003,N_4550,N_126);
and U9004 (N_9004,N_1820,N_1872);
xnor U9005 (N_9005,N_2463,N_1341);
or U9006 (N_9006,N_670,N_4220);
xnor U9007 (N_9007,N_2409,N_506);
nand U9008 (N_9008,N_1406,N_3302);
or U9009 (N_9009,N_2616,N_2300);
nor U9010 (N_9010,N_3422,N_380);
nor U9011 (N_9011,N_2375,N_4625);
and U9012 (N_9012,N_268,N_2263);
or U9013 (N_9013,N_1350,N_345);
or U9014 (N_9014,N_4353,N_1039);
xnor U9015 (N_9015,N_1398,N_4209);
or U9016 (N_9016,N_3207,N_4250);
and U9017 (N_9017,N_4275,N_4160);
and U9018 (N_9018,N_802,N_4360);
xnor U9019 (N_9019,N_1950,N_3995);
xor U9020 (N_9020,N_2775,N_3431);
nand U9021 (N_9021,N_4043,N_1563);
nor U9022 (N_9022,N_2019,N_4800);
and U9023 (N_9023,N_2893,N_3219);
and U9024 (N_9024,N_2232,N_3894);
nor U9025 (N_9025,N_3580,N_3248);
and U9026 (N_9026,N_659,N_3570);
and U9027 (N_9027,N_666,N_835);
nor U9028 (N_9028,N_1205,N_3152);
and U9029 (N_9029,N_37,N_1338);
or U9030 (N_9030,N_4511,N_4743);
nor U9031 (N_9031,N_1264,N_869);
xor U9032 (N_9032,N_796,N_316);
xor U9033 (N_9033,N_3656,N_1189);
nor U9034 (N_9034,N_488,N_2617);
or U9035 (N_9035,N_2371,N_4320);
xnor U9036 (N_9036,N_2007,N_3521);
nor U9037 (N_9037,N_2010,N_4564);
or U9038 (N_9038,N_4629,N_2093);
nand U9039 (N_9039,N_1168,N_4870);
or U9040 (N_9040,N_4675,N_2497);
nor U9041 (N_9041,N_758,N_1452);
nor U9042 (N_9042,N_3501,N_1871);
and U9043 (N_9043,N_3843,N_1319);
nand U9044 (N_9044,N_2070,N_283);
or U9045 (N_9045,N_3123,N_296);
nand U9046 (N_9046,N_1834,N_2326);
nand U9047 (N_9047,N_4552,N_3409);
nor U9048 (N_9048,N_3372,N_4723);
nand U9049 (N_9049,N_4793,N_4869);
and U9050 (N_9050,N_44,N_321);
nor U9051 (N_9051,N_707,N_1139);
nor U9052 (N_9052,N_3419,N_2938);
or U9053 (N_9053,N_3695,N_3814);
nor U9054 (N_9054,N_1776,N_4796);
xnor U9055 (N_9055,N_4862,N_184);
or U9056 (N_9056,N_378,N_1393);
nor U9057 (N_9057,N_3456,N_4168);
nor U9058 (N_9058,N_3814,N_1436);
xor U9059 (N_9059,N_4267,N_15);
and U9060 (N_9060,N_2176,N_1295);
xnor U9061 (N_9061,N_4114,N_2620);
and U9062 (N_9062,N_3541,N_732);
nor U9063 (N_9063,N_4662,N_3295);
nor U9064 (N_9064,N_2254,N_297);
xor U9065 (N_9065,N_4636,N_3079);
xor U9066 (N_9066,N_4022,N_454);
nor U9067 (N_9067,N_3349,N_1687);
xor U9068 (N_9068,N_1535,N_4044);
nor U9069 (N_9069,N_2106,N_4154);
nor U9070 (N_9070,N_4780,N_1706);
nand U9071 (N_9071,N_4770,N_1725);
and U9072 (N_9072,N_3207,N_3517);
nor U9073 (N_9073,N_2138,N_1918);
and U9074 (N_9074,N_766,N_1890);
nor U9075 (N_9075,N_3322,N_480);
and U9076 (N_9076,N_3916,N_4942);
nor U9077 (N_9077,N_2477,N_2293);
nor U9078 (N_9078,N_294,N_3746);
xor U9079 (N_9079,N_4995,N_3547);
nand U9080 (N_9080,N_3126,N_3040);
nand U9081 (N_9081,N_2029,N_3049);
and U9082 (N_9082,N_1499,N_1621);
or U9083 (N_9083,N_3684,N_2004);
nand U9084 (N_9084,N_3009,N_2298);
and U9085 (N_9085,N_1011,N_889);
or U9086 (N_9086,N_2106,N_4354);
nor U9087 (N_9087,N_784,N_1639);
or U9088 (N_9088,N_986,N_4266);
xor U9089 (N_9089,N_3274,N_3915);
and U9090 (N_9090,N_405,N_447);
and U9091 (N_9091,N_1955,N_606);
xnor U9092 (N_9092,N_743,N_333);
xor U9093 (N_9093,N_1003,N_2388);
or U9094 (N_9094,N_2940,N_2955);
xor U9095 (N_9095,N_1103,N_1695);
xor U9096 (N_9096,N_707,N_4246);
or U9097 (N_9097,N_836,N_2738);
nor U9098 (N_9098,N_1958,N_707);
nor U9099 (N_9099,N_1688,N_3885);
or U9100 (N_9100,N_3292,N_4128);
nor U9101 (N_9101,N_3330,N_4293);
nand U9102 (N_9102,N_2177,N_4777);
xor U9103 (N_9103,N_3991,N_1437);
nand U9104 (N_9104,N_3343,N_2414);
nand U9105 (N_9105,N_4848,N_1343);
nand U9106 (N_9106,N_888,N_203);
and U9107 (N_9107,N_2969,N_4050);
and U9108 (N_9108,N_87,N_3514);
or U9109 (N_9109,N_2691,N_90);
xor U9110 (N_9110,N_294,N_1019);
nor U9111 (N_9111,N_1296,N_2648);
nand U9112 (N_9112,N_1947,N_2784);
nor U9113 (N_9113,N_1542,N_2520);
or U9114 (N_9114,N_4717,N_2081);
nand U9115 (N_9115,N_4010,N_3647);
nor U9116 (N_9116,N_3437,N_4389);
and U9117 (N_9117,N_598,N_469);
xor U9118 (N_9118,N_1239,N_1742);
and U9119 (N_9119,N_2898,N_3239);
nor U9120 (N_9120,N_185,N_4907);
xnor U9121 (N_9121,N_4704,N_3719);
nand U9122 (N_9122,N_3598,N_2275);
xnor U9123 (N_9123,N_257,N_596);
xnor U9124 (N_9124,N_2809,N_4365);
nor U9125 (N_9125,N_1617,N_687);
and U9126 (N_9126,N_2337,N_342);
and U9127 (N_9127,N_4193,N_3930);
and U9128 (N_9128,N_4906,N_2709);
or U9129 (N_9129,N_4152,N_357);
xnor U9130 (N_9130,N_4549,N_3707);
nand U9131 (N_9131,N_2765,N_4579);
xnor U9132 (N_9132,N_3177,N_1475);
and U9133 (N_9133,N_1770,N_1076);
xor U9134 (N_9134,N_4265,N_665);
and U9135 (N_9135,N_918,N_3367);
xnor U9136 (N_9136,N_2099,N_3885);
and U9137 (N_9137,N_558,N_1388);
or U9138 (N_9138,N_4415,N_4205);
xor U9139 (N_9139,N_3715,N_3816);
and U9140 (N_9140,N_3236,N_1073);
or U9141 (N_9141,N_4705,N_752);
xor U9142 (N_9142,N_2695,N_3781);
nand U9143 (N_9143,N_697,N_3514);
xnor U9144 (N_9144,N_2391,N_3273);
nand U9145 (N_9145,N_2847,N_1551);
nand U9146 (N_9146,N_2472,N_3751);
or U9147 (N_9147,N_3892,N_3529);
or U9148 (N_9148,N_3163,N_1712);
and U9149 (N_9149,N_2037,N_3459);
nor U9150 (N_9150,N_1707,N_23);
nand U9151 (N_9151,N_4290,N_3659);
nor U9152 (N_9152,N_2926,N_3682);
nor U9153 (N_9153,N_1014,N_17);
xor U9154 (N_9154,N_4043,N_7);
nor U9155 (N_9155,N_2801,N_3689);
nor U9156 (N_9156,N_658,N_1067);
xnor U9157 (N_9157,N_1690,N_170);
nor U9158 (N_9158,N_1584,N_1317);
nand U9159 (N_9159,N_1636,N_789);
or U9160 (N_9160,N_1074,N_288);
and U9161 (N_9161,N_151,N_1041);
nor U9162 (N_9162,N_3875,N_651);
xnor U9163 (N_9163,N_4368,N_4000);
or U9164 (N_9164,N_1312,N_4110);
nand U9165 (N_9165,N_96,N_645);
xnor U9166 (N_9166,N_806,N_388);
nand U9167 (N_9167,N_4593,N_1945);
nor U9168 (N_9168,N_3226,N_2799);
or U9169 (N_9169,N_1941,N_4331);
nand U9170 (N_9170,N_4047,N_1462);
nor U9171 (N_9171,N_3730,N_4741);
xnor U9172 (N_9172,N_1587,N_307);
nand U9173 (N_9173,N_2945,N_3479);
nor U9174 (N_9174,N_2610,N_1555);
or U9175 (N_9175,N_808,N_1662);
xor U9176 (N_9176,N_4895,N_3899);
nor U9177 (N_9177,N_4530,N_409);
nor U9178 (N_9178,N_2994,N_3428);
nand U9179 (N_9179,N_3139,N_2538);
and U9180 (N_9180,N_2114,N_2477);
nand U9181 (N_9181,N_3289,N_3613);
xnor U9182 (N_9182,N_682,N_1055);
or U9183 (N_9183,N_3357,N_1772);
or U9184 (N_9184,N_218,N_4668);
nand U9185 (N_9185,N_2075,N_3940);
nand U9186 (N_9186,N_2364,N_1641);
nand U9187 (N_9187,N_3899,N_1638);
or U9188 (N_9188,N_3487,N_3316);
nor U9189 (N_9189,N_4371,N_1028);
xor U9190 (N_9190,N_2289,N_2055);
and U9191 (N_9191,N_4380,N_2009);
and U9192 (N_9192,N_2196,N_3346);
nor U9193 (N_9193,N_1970,N_2440);
or U9194 (N_9194,N_992,N_1721);
and U9195 (N_9195,N_4207,N_2097);
and U9196 (N_9196,N_1528,N_178);
nor U9197 (N_9197,N_4918,N_2192);
nand U9198 (N_9198,N_1228,N_2784);
xnor U9199 (N_9199,N_2624,N_469);
xor U9200 (N_9200,N_16,N_3876);
nor U9201 (N_9201,N_41,N_676);
nor U9202 (N_9202,N_2802,N_980);
xnor U9203 (N_9203,N_1417,N_2391);
nor U9204 (N_9204,N_3920,N_489);
and U9205 (N_9205,N_1243,N_2156);
xnor U9206 (N_9206,N_3513,N_3476);
nor U9207 (N_9207,N_2480,N_3211);
nand U9208 (N_9208,N_385,N_2714);
xor U9209 (N_9209,N_3083,N_307);
or U9210 (N_9210,N_3824,N_4337);
nor U9211 (N_9211,N_4081,N_4679);
nand U9212 (N_9212,N_4777,N_4470);
and U9213 (N_9213,N_1495,N_4406);
nand U9214 (N_9214,N_1866,N_973);
nand U9215 (N_9215,N_558,N_3961);
xor U9216 (N_9216,N_2222,N_3544);
and U9217 (N_9217,N_768,N_4502);
and U9218 (N_9218,N_2784,N_3677);
and U9219 (N_9219,N_18,N_482);
or U9220 (N_9220,N_3863,N_3855);
xnor U9221 (N_9221,N_549,N_605);
and U9222 (N_9222,N_3481,N_4096);
xor U9223 (N_9223,N_30,N_2611);
xor U9224 (N_9224,N_3174,N_367);
nand U9225 (N_9225,N_3025,N_3047);
nor U9226 (N_9226,N_3819,N_4220);
xnor U9227 (N_9227,N_1078,N_3101);
nor U9228 (N_9228,N_327,N_4522);
and U9229 (N_9229,N_4267,N_879);
nor U9230 (N_9230,N_3330,N_2397);
or U9231 (N_9231,N_1586,N_1684);
nand U9232 (N_9232,N_406,N_1665);
xnor U9233 (N_9233,N_4265,N_2128);
or U9234 (N_9234,N_2761,N_4682);
xor U9235 (N_9235,N_4261,N_43);
nor U9236 (N_9236,N_4679,N_453);
nor U9237 (N_9237,N_3738,N_2338);
or U9238 (N_9238,N_3267,N_1920);
nor U9239 (N_9239,N_2308,N_601);
nor U9240 (N_9240,N_1423,N_31);
xor U9241 (N_9241,N_1169,N_1367);
xnor U9242 (N_9242,N_2643,N_1430);
and U9243 (N_9243,N_533,N_3723);
nor U9244 (N_9244,N_1718,N_396);
or U9245 (N_9245,N_1306,N_481);
nor U9246 (N_9246,N_1015,N_2075);
nor U9247 (N_9247,N_3031,N_4519);
nand U9248 (N_9248,N_0,N_2480);
xnor U9249 (N_9249,N_2866,N_639);
or U9250 (N_9250,N_2463,N_179);
and U9251 (N_9251,N_419,N_3863);
or U9252 (N_9252,N_4382,N_2967);
nor U9253 (N_9253,N_1724,N_3562);
or U9254 (N_9254,N_2501,N_4628);
or U9255 (N_9255,N_2330,N_4219);
nand U9256 (N_9256,N_3568,N_726);
xnor U9257 (N_9257,N_2632,N_2545);
nor U9258 (N_9258,N_141,N_2813);
and U9259 (N_9259,N_1228,N_767);
xor U9260 (N_9260,N_3956,N_1657);
nor U9261 (N_9261,N_1065,N_3347);
or U9262 (N_9262,N_3824,N_1633);
or U9263 (N_9263,N_4737,N_2888);
and U9264 (N_9264,N_3249,N_2121);
and U9265 (N_9265,N_173,N_1851);
or U9266 (N_9266,N_4727,N_956);
nor U9267 (N_9267,N_4345,N_308);
nor U9268 (N_9268,N_1867,N_1947);
and U9269 (N_9269,N_207,N_1063);
and U9270 (N_9270,N_2971,N_1453);
nand U9271 (N_9271,N_22,N_2169);
nand U9272 (N_9272,N_2931,N_4058);
xnor U9273 (N_9273,N_949,N_1126);
nor U9274 (N_9274,N_119,N_1401);
xor U9275 (N_9275,N_242,N_1049);
and U9276 (N_9276,N_1928,N_84);
nor U9277 (N_9277,N_2925,N_1591);
nand U9278 (N_9278,N_4500,N_4045);
xnor U9279 (N_9279,N_520,N_4691);
and U9280 (N_9280,N_3272,N_3606);
or U9281 (N_9281,N_905,N_1229);
and U9282 (N_9282,N_1799,N_2650);
xor U9283 (N_9283,N_4424,N_2376);
nand U9284 (N_9284,N_2343,N_278);
or U9285 (N_9285,N_1938,N_4514);
nor U9286 (N_9286,N_977,N_1328);
nor U9287 (N_9287,N_3841,N_1711);
and U9288 (N_9288,N_266,N_4545);
nand U9289 (N_9289,N_146,N_4251);
xnor U9290 (N_9290,N_3284,N_885);
and U9291 (N_9291,N_963,N_4293);
and U9292 (N_9292,N_172,N_838);
and U9293 (N_9293,N_4066,N_4933);
or U9294 (N_9294,N_3699,N_4801);
xor U9295 (N_9295,N_1374,N_1977);
and U9296 (N_9296,N_4998,N_3356);
xor U9297 (N_9297,N_3272,N_4312);
nand U9298 (N_9298,N_3234,N_1511);
and U9299 (N_9299,N_965,N_3585);
nand U9300 (N_9300,N_4115,N_3468);
and U9301 (N_9301,N_2515,N_327);
nand U9302 (N_9302,N_1219,N_4758);
or U9303 (N_9303,N_41,N_1387);
and U9304 (N_9304,N_1428,N_578);
or U9305 (N_9305,N_730,N_4453);
and U9306 (N_9306,N_3443,N_2699);
nor U9307 (N_9307,N_416,N_3551);
and U9308 (N_9308,N_4056,N_3895);
nor U9309 (N_9309,N_1937,N_3190);
nor U9310 (N_9310,N_1732,N_3236);
nor U9311 (N_9311,N_4548,N_4227);
nand U9312 (N_9312,N_4541,N_3874);
nor U9313 (N_9313,N_4688,N_2610);
nor U9314 (N_9314,N_4236,N_393);
nor U9315 (N_9315,N_3715,N_3471);
nand U9316 (N_9316,N_1821,N_3420);
and U9317 (N_9317,N_2507,N_2989);
nand U9318 (N_9318,N_992,N_3466);
or U9319 (N_9319,N_1778,N_2733);
and U9320 (N_9320,N_1621,N_3789);
xor U9321 (N_9321,N_221,N_2007);
or U9322 (N_9322,N_4168,N_930);
or U9323 (N_9323,N_2805,N_3061);
xor U9324 (N_9324,N_2558,N_455);
nor U9325 (N_9325,N_2228,N_3981);
or U9326 (N_9326,N_4361,N_2899);
xnor U9327 (N_9327,N_4740,N_493);
and U9328 (N_9328,N_3495,N_2006);
or U9329 (N_9329,N_1449,N_2204);
and U9330 (N_9330,N_486,N_3018);
xor U9331 (N_9331,N_644,N_2879);
and U9332 (N_9332,N_3276,N_3388);
nand U9333 (N_9333,N_2421,N_4627);
or U9334 (N_9334,N_1695,N_829);
xnor U9335 (N_9335,N_3805,N_2003);
nor U9336 (N_9336,N_487,N_2255);
or U9337 (N_9337,N_4183,N_2308);
nor U9338 (N_9338,N_542,N_241);
and U9339 (N_9339,N_3654,N_2489);
xnor U9340 (N_9340,N_4991,N_4943);
or U9341 (N_9341,N_624,N_2755);
or U9342 (N_9342,N_4900,N_4176);
nor U9343 (N_9343,N_4602,N_4653);
nor U9344 (N_9344,N_3531,N_958);
nor U9345 (N_9345,N_3799,N_2195);
or U9346 (N_9346,N_29,N_4889);
or U9347 (N_9347,N_2643,N_2970);
nand U9348 (N_9348,N_3252,N_992);
and U9349 (N_9349,N_1512,N_2400);
nand U9350 (N_9350,N_3150,N_1147);
or U9351 (N_9351,N_4354,N_3526);
nor U9352 (N_9352,N_4030,N_1159);
nor U9353 (N_9353,N_559,N_178);
nand U9354 (N_9354,N_980,N_1752);
xnor U9355 (N_9355,N_2548,N_993);
nand U9356 (N_9356,N_1396,N_696);
xor U9357 (N_9357,N_4372,N_3077);
and U9358 (N_9358,N_1628,N_3136);
xnor U9359 (N_9359,N_2115,N_587);
and U9360 (N_9360,N_573,N_1767);
xnor U9361 (N_9361,N_1510,N_2351);
xor U9362 (N_9362,N_1829,N_3139);
or U9363 (N_9363,N_2107,N_2464);
nor U9364 (N_9364,N_3945,N_3982);
and U9365 (N_9365,N_774,N_318);
and U9366 (N_9366,N_2259,N_1041);
nor U9367 (N_9367,N_4374,N_1297);
and U9368 (N_9368,N_592,N_2902);
nand U9369 (N_9369,N_124,N_1666);
and U9370 (N_9370,N_4852,N_4797);
xor U9371 (N_9371,N_3408,N_2134);
or U9372 (N_9372,N_2731,N_2919);
and U9373 (N_9373,N_2297,N_4861);
nor U9374 (N_9374,N_4092,N_2049);
nand U9375 (N_9375,N_1535,N_3231);
nand U9376 (N_9376,N_3015,N_3004);
or U9377 (N_9377,N_4459,N_4319);
nand U9378 (N_9378,N_2390,N_2817);
nand U9379 (N_9379,N_2361,N_2163);
nor U9380 (N_9380,N_4956,N_1986);
nor U9381 (N_9381,N_3449,N_3752);
and U9382 (N_9382,N_486,N_1125);
nand U9383 (N_9383,N_4827,N_3186);
or U9384 (N_9384,N_4395,N_2228);
or U9385 (N_9385,N_909,N_2669);
and U9386 (N_9386,N_4404,N_141);
nand U9387 (N_9387,N_1728,N_2862);
nor U9388 (N_9388,N_3912,N_1826);
nand U9389 (N_9389,N_3329,N_4506);
or U9390 (N_9390,N_2414,N_4016);
nand U9391 (N_9391,N_1342,N_4880);
nand U9392 (N_9392,N_4017,N_4496);
xnor U9393 (N_9393,N_928,N_2672);
xor U9394 (N_9394,N_2312,N_2917);
xor U9395 (N_9395,N_2236,N_3010);
nand U9396 (N_9396,N_4622,N_4387);
or U9397 (N_9397,N_2955,N_2758);
nand U9398 (N_9398,N_2938,N_3352);
or U9399 (N_9399,N_3878,N_4582);
xor U9400 (N_9400,N_50,N_2037);
and U9401 (N_9401,N_2456,N_4081);
xor U9402 (N_9402,N_65,N_1160);
nor U9403 (N_9403,N_3597,N_2155);
nand U9404 (N_9404,N_1010,N_4012);
nand U9405 (N_9405,N_2000,N_3165);
nor U9406 (N_9406,N_4042,N_4419);
nand U9407 (N_9407,N_3574,N_958);
nand U9408 (N_9408,N_803,N_239);
and U9409 (N_9409,N_1902,N_3841);
nor U9410 (N_9410,N_2942,N_2790);
and U9411 (N_9411,N_1804,N_809);
and U9412 (N_9412,N_4807,N_2988);
xnor U9413 (N_9413,N_1563,N_336);
nor U9414 (N_9414,N_2661,N_2580);
nor U9415 (N_9415,N_544,N_3908);
xor U9416 (N_9416,N_1270,N_4607);
nor U9417 (N_9417,N_3875,N_222);
and U9418 (N_9418,N_855,N_3303);
or U9419 (N_9419,N_3987,N_3066);
xnor U9420 (N_9420,N_4296,N_4714);
nand U9421 (N_9421,N_3714,N_417);
and U9422 (N_9422,N_96,N_1670);
xnor U9423 (N_9423,N_1017,N_3167);
or U9424 (N_9424,N_2216,N_2885);
nand U9425 (N_9425,N_865,N_61);
xnor U9426 (N_9426,N_610,N_1658);
nand U9427 (N_9427,N_2194,N_4824);
and U9428 (N_9428,N_2211,N_4710);
nand U9429 (N_9429,N_4301,N_522);
nand U9430 (N_9430,N_2914,N_4637);
nand U9431 (N_9431,N_4538,N_2325);
nand U9432 (N_9432,N_1127,N_1093);
xnor U9433 (N_9433,N_2727,N_1406);
nand U9434 (N_9434,N_36,N_2886);
or U9435 (N_9435,N_4839,N_640);
xor U9436 (N_9436,N_324,N_1480);
xor U9437 (N_9437,N_654,N_4434);
nand U9438 (N_9438,N_889,N_2681);
or U9439 (N_9439,N_3307,N_1738);
nor U9440 (N_9440,N_2730,N_4870);
and U9441 (N_9441,N_2224,N_2871);
xnor U9442 (N_9442,N_4994,N_1032);
nor U9443 (N_9443,N_2627,N_4839);
nand U9444 (N_9444,N_1172,N_2021);
or U9445 (N_9445,N_943,N_391);
or U9446 (N_9446,N_4492,N_4951);
and U9447 (N_9447,N_3006,N_4751);
and U9448 (N_9448,N_1888,N_2115);
nor U9449 (N_9449,N_1135,N_4828);
or U9450 (N_9450,N_1504,N_3715);
nand U9451 (N_9451,N_2076,N_4906);
or U9452 (N_9452,N_2841,N_4582);
and U9453 (N_9453,N_1315,N_767);
nand U9454 (N_9454,N_1092,N_2155);
or U9455 (N_9455,N_1886,N_1258);
nand U9456 (N_9456,N_4853,N_4890);
and U9457 (N_9457,N_4209,N_3710);
nor U9458 (N_9458,N_4025,N_1110);
nand U9459 (N_9459,N_2065,N_3260);
or U9460 (N_9460,N_3227,N_1117);
nand U9461 (N_9461,N_4888,N_984);
and U9462 (N_9462,N_4447,N_3024);
nand U9463 (N_9463,N_732,N_1200);
and U9464 (N_9464,N_3943,N_1145);
or U9465 (N_9465,N_4874,N_4603);
xor U9466 (N_9466,N_4584,N_1054);
and U9467 (N_9467,N_1149,N_1375);
xor U9468 (N_9468,N_4779,N_4455);
or U9469 (N_9469,N_3977,N_2564);
xor U9470 (N_9470,N_911,N_1030);
xor U9471 (N_9471,N_159,N_2125);
nand U9472 (N_9472,N_1710,N_4608);
xor U9473 (N_9473,N_4432,N_4783);
and U9474 (N_9474,N_643,N_619);
and U9475 (N_9475,N_4391,N_2861);
xnor U9476 (N_9476,N_2535,N_1160);
and U9477 (N_9477,N_514,N_185);
xor U9478 (N_9478,N_4408,N_3664);
or U9479 (N_9479,N_24,N_2586);
nand U9480 (N_9480,N_314,N_4166);
and U9481 (N_9481,N_2517,N_4230);
nor U9482 (N_9482,N_2707,N_2157);
or U9483 (N_9483,N_3445,N_2364);
xnor U9484 (N_9484,N_4986,N_3564);
and U9485 (N_9485,N_3361,N_2735);
and U9486 (N_9486,N_3915,N_475);
nand U9487 (N_9487,N_3059,N_1989);
and U9488 (N_9488,N_3583,N_3961);
nor U9489 (N_9489,N_611,N_83);
and U9490 (N_9490,N_96,N_46);
nor U9491 (N_9491,N_3495,N_3464);
or U9492 (N_9492,N_3792,N_2125);
xnor U9493 (N_9493,N_489,N_1196);
xor U9494 (N_9494,N_1673,N_3171);
or U9495 (N_9495,N_4046,N_4002);
nand U9496 (N_9496,N_3908,N_781);
xnor U9497 (N_9497,N_1309,N_4587);
and U9498 (N_9498,N_3103,N_3737);
nand U9499 (N_9499,N_2114,N_1734);
xor U9500 (N_9500,N_3978,N_4745);
nand U9501 (N_9501,N_3506,N_4804);
nand U9502 (N_9502,N_2469,N_1622);
nor U9503 (N_9503,N_2247,N_2474);
xnor U9504 (N_9504,N_1486,N_703);
or U9505 (N_9505,N_3136,N_1959);
xor U9506 (N_9506,N_4629,N_1561);
xor U9507 (N_9507,N_2259,N_4821);
and U9508 (N_9508,N_4194,N_1370);
nand U9509 (N_9509,N_3917,N_3177);
or U9510 (N_9510,N_695,N_4247);
nand U9511 (N_9511,N_1174,N_3303);
and U9512 (N_9512,N_505,N_2736);
xor U9513 (N_9513,N_477,N_2950);
and U9514 (N_9514,N_1873,N_3151);
xnor U9515 (N_9515,N_3802,N_1720);
and U9516 (N_9516,N_2807,N_4235);
or U9517 (N_9517,N_417,N_297);
nand U9518 (N_9518,N_1825,N_1290);
or U9519 (N_9519,N_1907,N_1045);
and U9520 (N_9520,N_4257,N_4655);
nand U9521 (N_9521,N_3394,N_1459);
xor U9522 (N_9522,N_3202,N_1544);
xnor U9523 (N_9523,N_3920,N_1128);
xor U9524 (N_9524,N_1510,N_3686);
or U9525 (N_9525,N_3624,N_1890);
nand U9526 (N_9526,N_2327,N_1058);
nor U9527 (N_9527,N_3866,N_4812);
xor U9528 (N_9528,N_402,N_3842);
xnor U9529 (N_9529,N_4737,N_3897);
or U9530 (N_9530,N_836,N_2907);
xnor U9531 (N_9531,N_3936,N_1455);
nor U9532 (N_9532,N_123,N_444);
or U9533 (N_9533,N_4484,N_4074);
and U9534 (N_9534,N_2218,N_3247);
and U9535 (N_9535,N_3449,N_3733);
nand U9536 (N_9536,N_1629,N_3752);
nand U9537 (N_9537,N_4592,N_1088);
xor U9538 (N_9538,N_4487,N_2519);
or U9539 (N_9539,N_2011,N_4376);
nand U9540 (N_9540,N_3144,N_1615);
or U9541 (N_9541,N_1209,N_2011);
and U9542 (N_9542,N_4840,N_685);
and U9543 (N_9543,N_3580,N_3982);
and U9544 (N_9544,N_2253,N_1323);
or U9545 (N_9545,N_2870,N_182);
and U9546 (N_9546,N_1321,N_3431);
nor U9547 (N_9547,N_4722,N_4049);
and U9548 (N_9548,N_2780,N_2066);
and U9549 (N_9549,N_965,N_4160);
or U9550 (N_9550,N_1140,N_4784);
or U9551 (N_9551,N_1427,N_441);
xnor U9552 (N_9552,N_3241,N_4713);
or U9553 (N_9553,N_3886,N_1751);
nand U9554 (N_9554,N_3409,N_988);
or U9555 (N_9555,N_4489,N_2152);
or U9556 (N_9556,N_612,N_2042);
xnor U9557 (N_9557,N_1130,N_2219);
xnor U9558 (N_9558,N_4931,N_1820);
nand U9559 (N_9559,N_1149,N_1916);
or U9560 (N_9560,N_3557,N_854);
nand U9561 (N_9561,N_1371,N_3055);
or U9562 (N_9562,N_3369,N_3928);
nor U9563 (N_9563,N_4808,N_124);
xor U9564 (N_9564,N_2732,N_2001);
xnor U9565 (N_9565,N_1231,N_4350);
or U9566 (N_9566,N_1067,N_2101);
nand U9567 (N_9567,N_2246,N_3990);
and U9568 (N_9568,N_3661,N_721);
and U9569 (N_9569,N_1641,N_2550);
xor U9570 (N_9570,N_4356,N_2808);
or U9571 (N_9571,N_1349,N_4243);
and U9572 (N_9572,N_307,N_1420);
and U9573 (N_9573,N_720,N_3344);
and U9574 (N_9574,N_3203,N_2881);
or U9575 (N_9575,N_4862,N_3295);
xor U9576 (N_9576,N_3691,N_258);
xor U9577 (N_9577,N_708,N_1331);
nor U9578 (N_9578,N_628,N_774);
nor U9579 (N_9579,N_2450,N_1423);
and U9580 (N_9580,N_3608,N_2438);
or U9581 (N_9581,N_375,N_4335);
or U9582 (N_9582,N_2742,N_4102);
xnor U9583 (N_9583,N_4022,N_1941);
nor U9584 (N_9584,N_1248,N_1559);
nand U9585 (N_9585,N_825,N_1564);
nor U9586 (N_9586,N_1721,N_207);
nor U9587 (N_9587,N_2504,N_2815);
or U9588 (N_9588,N_1672,N_1996);
or U9589 (N_9589,N_1346,N_701);
xor U9590 (N_9590,N_2518,N_2579);
or U9591 (N_9591,N_1004,N_1545);
or U9592 (N_9592,N_4948,N_1964);
or U9593 (N_9593,N_2349,N_559);
and U9594 (N_9594,N_476,N_1610);
and U9595 (N_9595,N_2921,N_93);
or U9596 (N_9596,N_788,N_3426);
nand U9597 (N_9597,N_83,N_1997);
or U9598 (N_9598,N_4794,N_4693);
xnor U9599 (N_9599,N_1171,N_3056);
nand U9600 (N_9600,N_3741,N_1706);
nor U9601 (N_9601,N_3296,N_3644);
nor U9602 (N_9602,N_887,N_226);
and U9603 (N_9603,N_566,N_4110);
xor U9604 (N_9604,N_1621,N_4782);
and U9605 (N_9605,N_1157,N_185);
nor U9606 (N_9606,N_2323,N_2867);
nor U9607 (N_9607,N_1630,N_634);
xnor U9608 (N_9608,N_1482,N_1077);
xnor U9609 (N_9609,N_1285,N_825);
xor U9610 (N_9610,N_2737,N_673);
and U9611 (N_9611,N_4906,N_2584);
or U9612 (N_9612,N_4235,N_3225);
xnor U9613 (N_9613,N_3587,N_1206);
nand U9614 (N_9614,N_4675,N_4628);
and U9615 (N_9615,N_3421,N_1345);
nand U9616 (N_9616,N_1409,N_1113);
nand U9617 (N_9617,N_2654,N_4428);
or U9618 (N_9618,N_2643,N_1211);
and U9619 (N_9619,N_1921,N_3178);
nand U9620 (N_9620,N_781,N_4023);
nor U9621 (N_9621,N_705,N_3286);
or U9622 (N_9622,N_3078,N_2185);
xor U9623 (N_9623,N_2280,N_4136);
nor U9624 (N_9624,N_4575,N_4000);
and U9625 (N_9625,N_2715,N_2112);
or U9626 (N_9626,N_3163,N_2587);
nor U9627 (N_9627,N_4224,N_4411);
nor U9628 (N_9628,N_2813,N_1629);
or U9629 (N_9629,N_1102,N_619);
nor U9630 (N_9630,N_2320,N_2828);
nor U9631 (N_9631,N_3518,N_3019);
and U9632 (N_9632,N_4094,N_2712);
nor U9633 (N_9633,N_1780,N_3121);
nor U9634 (N_9634,N_3180,N_4776);
xnor U9635 (N_9635,N_2337,N_184);
and U9636 (N_9636,N_352,N_2319);
or U9637 (N_9637,N_3800,N_2950);
nor U9638 (N_9638,N_1627,N_1578);
nor U9639 (N_9639,N_922,N_4367);
nand U9640 (N_9640,N_923,N_4315);
nand U9641 (N_9641,N_1148,N_4354);
and U9642 (N_9642,N_1333,N_2276);
nor U9643 (N_9643,N_1734,N_4106);
nand U9644 (N_9644,N_4735,N_926);
or U9645 (N_9645,N_905,N_2106);
nand U9646 (N_9646,N_1580,N_3975);
and U9647 (N_9647,N_3884,N_3857);
and U9648 (N_9648,N_700,N_4219);
and U9649 (N_9649,N_3370,N_1069);
and U9650 (N_9650,N_2666,N_1014);
or U9651 (N_9651,N_3581,N_2759);
and U9652 (N_9652,N_1439,N_4913);
nor U9653 (N_9653,N_1089,N_450);
nor U9654 (N_9654,N_554,N_1643);
and U9655 (N_9655,N_775,N_4264);
and U9656 (N_9656,N_1247,N_628);
and U9657 (N_9657,N_2387,N_1328);
nor U9658 (N_9658,N_1780,N_402);
nor U9659 (N_9659,N_4470,N_1694);
nand U9660 (N_9660,N_2829,N_484);
nand U9661 (N_9661,N_4786,N_976);
xor U9662 (N_9662,N_3569,N_4850);
xor U9663 (N_9663,N_4568,N_1722);
nand U9664 (N_9664,N_70,N_3562);
nand U9665 (N_9665,N_1118,N_2967);
or U9666 (N_9666,N_1485,N_1957);
and U9667 (N_9667,N_1549,N_2397);
nor U9668 (N_9668,N_4620,N_1649);
xnor U9669 (N_9669,N_2060,N_1806);
xor U9670 (N_9670,N_3448,N_4811);
nand U9671 (N_9671,N_4870,N_1658);
or U9672 (N_9672,N_376,N_4490);
and U9673 (N_9673,N_4206,N_4092);
xnor U9674 (N_9674,N_947,N_3934);
and U9675 (N_9675,N_4736,N_2340);
nor U9676 (N_9676,N_985,N_3789);
nor U9677 (N_9677,N_783,N_2393);
nand U9678 (N_9678,N_2469,N_1111);
and U9679 (N_9679,N_2867,N_2106);
xnor U9680 (N_9680,N_4230,N_3802);
and U9681 (N_9681,N_2940,N_3444);
xnor U9682 (N_9682,N_1624,N_3430);
or U9683 (N_9683,N_2614,N_3936);
or U9684 (N_9684,N_780,N_2692);
nand U9685 (N_9685,N_433,N_228);
and U9686 (N_9686,N_3544,N_1062);
or U9687 (N_9687,N_3837,N_1633);
nor U9688 (N_9688,N_3106,N_4617);
or U9689 (N_9689,N_475,N_4960);
nor U9690 (N_9690,N_2719,N_4983);
and U9691 (N_9691,N_1482,N_3578);
xor U9692 (N_9692,N_574,N_4932);
and U9693 (N_9693,N_4773,N_1425);
nor U9694 (N_9694,N_4372,N_4586);
and U9695 (N_9695,N_366,N_4925);
and U9696 (N_9696,N_1709,N_4754);
nand U9697 (N_9697,N_3528,N_431);
xnor U9698 (N_9698,N_3102,N_2754);
nand U9699 (N_9699,N_3469,N_769);
nor U9700 (N_9700,N_1172,N_2681);
and U9701 (N_9701,N_2209,N_4847);
or U9702 (N_9702,N_4307,N_709);
nand U9703 (N_9703,N_73,N_842);
and U9704 (N_9704,N_3958,N_187);
xor U9705 (N_9705,N_2750,N_1789);
nor U9706 (N_9706,N_35,N_4082);
xnor U9707 (N_9707,N_3995,N_3004);
nand U9708 (N_9708,N_1384,N_4816);
or U9709 (N_9709,N_1872,N_519);
nand U9710 (N_9710,N_2760,N_3307);
xnor U9711 (N_9711,N_1281,N_2163);
nand U9712 (N_9712,N_3598,N_3232);
nand U9713 (N_9713,N_19,N_1290);
nor U9714 (N_9714,N_1510,N_437);
nand U9715 (N_9715,N_1824,N_4979);
nor U9716 (N_9716,N_3417,N_770);
nor U9717 (N_9717,N_3641,N_3331);
nand U9718 (N_9718,N_1296,N_2249);
and U9719 (N_9719,N_599,N_3752);
and U9720 (N_9720,N_2434,N_1415);
and U9721 (N_9721,N_1939,N_1584);
nand U9722 (N_9722,N_308,N_1388);
nor U9723 (N_9723,N_4487,N_483);
nand U9724 (N_9724,N_1519,N_902);
nor U9725 (N_9725,N_2579,N_1212);
or U9726 (N_9726,N_161,N_2054);
xnor U9727 (N_9727,N_3355,N_3419);
or U9728 (N_9728,N_3413,N_2666);
or U9729 (N_9729,N_4967,N_1794);
nand U9730 (N_9730,N_2506,N_3343);
nor U9731 (N_9731,N_1020,N_174);
and U9732 (N_9732,N_2665,N_1131);
or U9733 (N_9733,N_559,N_1068);
nor U9734 (N_9734,N_634,N_1432);
nor U9735 (N_9735,N_2536,N_3819);
nand U9736 (N_9736,N_1019,N_1231);
xor U9737 (N_9737,N_2765,N_1852);
or U9738 (N_9738,N_1419,N_582);
or U9739 (N_9739,N_2580,N_4133);
xnor U9740 (N_9740,N_2130,N_88);
nand U9741 (N_9741,N_1942,N_3707);
nor U9742 (N_9742,N_1290,N_3291);
xnor U9743 (N_9743,N_2296,N_661);
nand U9744 (N_9744,N_3867,N_868);
nand U9745 (N_9745,N_4407,N_1321);
xor U9746 (N_9746,N_4153,N_301);
and U9747 (N_9747,N_1806,N_4457);
nand U9748 (N_9748,N_2007,N_4709);
xor U9749 (N_9749,N_1751,N_171);
nand U9750 (N_9750,N_2795,N_3159);
nand U9751 (N_9751,N_2264,N_1856);
nor U9752 (N_9752,N_4818,N_1655);
nor U9753 (N_9753,N_1179,N_2004);
and U9754 (N_9754,N_2002,N_3633);
nand U9755 (N_9755,N_3406,N_4753);
xnor U9756 (N_9756,N_693,N_2196);
nor U9757 (N_9757,N_2678,N_2980);
xnor U9758 (N_9758,N_1125,N_4933);
or U9759 (N_9759,N_251,N_4821);
and U9760 (N_9760,N_1559,N_751);
nor U9761 (N_9761,N_2155,N_224);
or U9762 (N_9762,N_4965,N_1347);
and U9763 (N_9763,N_3583,N_3941);
nor U9764 (N_9764,N_3205,N_4657);
and U9765 (N_9765,N_2477,N_1254);
xor U9766 (N_9766,N_4162,N_840);
or U9767 (N_9767,N_2458,N_4834);
nor U9768 (N_9768,N_765,N_3588);
and U9769 (N_9769,N_4452,N_4257);
nor U9770 (N_9770,N_987,N_1158);
nor U9771 (N_9771,N_3306,N_3235);
and U9772 (N_9772,N_703,N_3797);
xor U9773 (N_9773,N_1484,N_556);
xnor U9774 (N_9774,N_1063,N_3262);
nor U9775 (N_9775,N_2844,N_1769);
and U9776 (N_9776,N_1633,N_485);
or U9777 (N_9777,N_1911,N_2929);
xnor U9778 (N_9778,N_2201,N_485);
or U9779 (N_9779,N_1415,N_1284);
nand U9780 (N_9780,N_4490,N_4293);
and U9781 (N_9781,N_2838,N_4394);
and U9782 (N_9782,N_1704,N_364);
nor U9783 (N_9783,N_1472,N_4142);
nor U9784 (N_9784,N_1375,N_2093);
xor U9785 (N_9785,N_1585,N_980);
nand U9786 (N_9786,N_4421,N_1646);
nor U9787 (N_9787,N_570,N_3521);
xnor U9788 (N_9788,N_4360,N_2402);
nand U9789 (N_9789,N_2375,N_1776);
or U9790 (N_9790,N_2841,N_679);
xor U9791 (N_9791,N_2627,N_2717);
and U9792 (N_9792,N_3074,N_424);
nand U9793 (N_9793,N_1241,N_870);
and U9794 (N_9794,N_3138,N_2552);
nand U9795 (N_9795,N_226,N_499);
or U9796 (N_9796,N_1904,N_2701);
nor U9797 (N_9797,N_3844,N_1320);
xnor U9798 (N_9798,N_2029,N_3503);
xor U9799 (N_9799,N_2973,N_1343);
xor U9800 (N_9800,N_3170,N_1462);
or U9801 (N_9801,N_1250,N_2510);
nand U9802 (N_9802,N_3592,N_2996);
xor U9803 (N_9803,N_3425,N_306);
or U9804 (N_9804,N_1469,N_973);
nor U9805 (N_9805,N_175,N_714);
nand U9806 (N_9806,N_4424,N_937);
and U9807 (N_9807,N_165,N_8);
or U9808 (N_9808,N_4961,N_4182);
or U9809 (N_9809,N_4343,N_1772);
xnor U9810 (N_9810,N_4905,N_1197);
nor U9811 (N_9811,N_2136,N_3555);
nand U9812 (N_9812,N_15,N_1882);
nand U9813 (N_9813,N_4472,N_2876);
nand U9814 (N_9814,N_3341,N_545);
xnor U9815 (N_9815,N_1087,N_4346);
or U9816 (N_9816,N_3028,N_952);
xnor U9817 (N_9817,N_4675,N_4414);
and U9818 (N_9818,N_2961,N_610);
xnor U9819 (N_9819,N_2947,N_3541);
nand U9820 (N_9820,N_1422,N_3330);
nor U9821 (N_9821,N_2465,N_4334);
xor U9822 (N_9822,N_1029,N_2866);
or U9823 (N_9823,N_1271,N_2397);
or U9824 (N_9824,N_3779,N_1807);
or U9825 (N_9825,N_4378,N_3888);
or U9826 (N_9826,N_2011,N_4262);
or U9827 (N_9827,N_2848,N_44);
nand U9828 (N_9828,N_3712,N_50);
nand U9829 (N_9829,N_2774,N_2576);
or U9830 (N_9830,N_1877,N_2914);
nor U9831 (N_9831,N_1656,N_2130);
nor U9832 (N_9832,N_3834,N_4633);
nor U9833 (N_9833,N_1822,N_4788);
and U9834 (N_9834,N_1038,N_532);
xnor U9835 (N_9835,N_2179,N_4628);
nor U9836 (N_9836,N_4254,N_4568);
and U9837 (N_9837,N_3689,N_34);
or U9838 (N_9838,N_3578,N_2459);
xnor U9839 (N_9839,N_1792,N_2675);
nor U9840 (N_9840,N_3480,N_637);
nand U9841 (N_9841,N_1185,N_4466);
or U9842 (N_9842,N_2645,N_3811);
and U9843 (N_9843,N_3102,N_3105);
nand U9844 (N_9844,N_2394,N_1244);
and U9845 (N_9845,N_1756,N_4379);
or U9846 (N_9846,N_3622,N_853);
or U9847 (N_9847,N_1232,N_4056);
xor U9848 (N_9848,N_1978,N_1808);
and U9849 (N_9849,N_389,N_149);
or U9850 (N_9850,N_3852,N_348);
or U9851 (N_9851,N_1145,N_4054);
or U9852 (N_9852,N_3790,N_3820);
or U9853 (N_9853,N_1884,N_3628);
xnor U9854 (N_9854,N_3807,N_2012);
nand U9855 (N_9855,N_1895,N_428);
or U9856 (N_9856,N_4486,N_847);
or U9857 (N_9857,N_3416,N_4015);
or U9858 (N_9858,N_2156,N_178);
or U9859 (N_9859,N_3309,N_1527);
and U9860 (N_9860,N_188,N_4168);
nand U9861 (N_9861,N_3349,N_3030);
and U9862 (N_9862,N_4238,N_1181);
xnor U9863 (N_9863,N_2703,N_3541);
xnor U9864 (N_9864,N_3742,N_2111);
or U9865 (N_9865,N_4033,N_504);
or U9866 (N_9866,N_3850,N_487);
or U9867 (N_9867,N_2181,N_2736);
nor U9868 (N_9868,N_2920,N_3276);
or U9869 (N_9869,N_4571,N_454);
and U9870 (N_9870,N_3447,N_4936);
nor U9871 (N_9871,N_778,N_2231);
and U9872 (N_9872,N_1455,N_1145);
nand U9873 (N_9873,N_3548,N_2093);
and U9874 (N_9874,N_4789,N_2252);
and U9875 (N_9875,N_1645,N_4478);
xnor U9876 (N_9876,N_964,N_433);
and U9877 (N_9877,N_2803,N_2681);
nand U9878 (N_9878,N_2056,N_482);
xor U9879 (N_9879,N_712,N_2500);
and U9880 (N_9880,N_1895,N_4935);
nor U9881 (N_9881,N_4593,N_1490);
and U9882 (N_9882,N_1640,N_4051);
xor U9883 (N_9883,N_2295,N_322);
nor U9884 (N_9884,N_4320,N_934);
and U9885 (N_9885,N_3773,N_4453);
xnor U9886 (N_9886,N_568,N_340);
xor U9887 (N_9887,N_2740,N_3941);
nor U9888 (N_9888,N_464,N_803);
xor U9889 (N_9889,N_3908,N_504);
nor U9890 (N_9890,N_3613,N_226);
nor U9891 (N_9891,N_3903,N_887);
or U9892 (N_9892,N_4285,N_4994);
nand U9893 (N_9893,N_553,N_2128);
nand U9894 (N_9894,N_1292,N_4384);
nand U9895 (N_9895,N_4516,N_4651);
nor U9896 (N_9896,N_4899,N_3302);
and U9897 (N_9897,N_2928,N_3368);
xnor U9898 (N_9898,N_3167,N_768);
nor U9899 (N_9899,N_3955,N_2278);
xnor U9900 (N_9900,N_3480,N_3363);
or U9901 (N_9901,N_1460,N_370);
xor U9902 (N_9902,N_4107,N_1023);
xnor U9903 (N_9903,N_3339,N_2583);
or U9904 (N_9904,N_4055,N_1147);
xnor U9905 (N_9905,N_2348,N_2473);
nand U9906 (N_9906,N_4885,N_2186);
nand U9907 (N_9907,N_2195,N_492);
xor U9908 (N_9908,N_2754,N_1803);
nor U9909 (N_9909,N_597,N_3444);
nor U9910 (N_9910,N_303,N_3083);
xor U9911 (N_9911,N_1042,N_2196);
nand U9912 (N_9912,N_2632,N_1452);
nor U9913 (N_9913,N_2208,N_589);
nor U9914 (N_9914,N_3350,N_3179);
or U9915 (N_9915,N_4042,N_2000);
nand U9916 (N_9916,N_2581,N_3332);
or U9917 (N_9917,N_420,N_4917);
or U9918 (N_9918,N_742,N_2940);
nor U9919 (N_9919,N_2508,N_2699);
and U9920 (N_9920,N_4500,N_4584);
and U9921 (N_9921,N_3685,N_1715);
nand U9922 (N_9922,N_4823,N_3752);
nor U9923 (N_9923,N_3156,N_2764);
nand U9924 (N_9924,N_2345,N_2138);
xnor U9925 (N_9925,N_3923,N_374);
nor U9926 (N_9926,N_1371,N_3240);
nor U9927 (N_9927,N_3828,N_403);
nand U9928 (N_9928,N_406,N_1210);
nor U9929 (N_9929,N_965,N_2794);
nor U9930 (N_9930,N_3546,N_48);
nand U9931 (N_9931,N_4184,N_1910);
and U9932 (N_9932,N_3507,N_1923);
and U9933 (N_9933,N_37,N_4497);
nor U9934 (N_9934,N_2317,N_2094);
xor U9935 (N_9935,N_2769,N_2278);
or U9936 (N_9936,N_2732,N_4883);
nor U9937 (N_9937,N_416,N_4363);
and U9938 (N_9938,N_1024,N_1243);
nand U9939 (N_9939,N_1599,N_1412);
nand U9940 (N_9940,N_1646,N_2568);
nor U9941 (N_9941,N_4709,N_4934);
xor U9942 (N_9942,N_1278,N_1489);
and U9943 (N_9943,N_822,N_3185);
or U9944 (N_9944,N_3576,N_3598);
nand U9945 (N_9945,N_201,N_1318);
xnor U9946 (N_9946,N_2179,N_4937);
and U9947 (N_9947,N_950,N_4969);
or U9948 (N_9948,N_4467,N_354);
xnor U9949 (N_9949,N_4390,N_4535);
and U9950 (N_9950,N_4459,N_3964);
nor U9951 (N_9951,N_4987,N_127);
or U9952 (N_9952,N_1142,N_3642);
nand U9953 (N_9953,N_110,N_3485);
nor U9954 (N_9954,N_2387,N_1498);
xor U9955 (N_9955,N_1852,N_4776);
xor U9956 (N_9956,N_2306,N_38);
xnor U9957 (N_9957,N_1449,N_2933);
nor U9958 (N_9958,N_3570,N_695);
nor U9959 (N_9959,N_2678,N_4420);
and U9960 (N_9960,N_54,N_4140);
nor U9961 (N_9961,N_148,N_2322);
nor U9962 (N_9962,N_203,N_4783);
or U9963 (N_9963,N_4819,N_775);
or U9964 (N_9964,N_3087,N_3668);
xnor U9965 (N_9965,N_1772,N_691);
or U9966 (N_9966,N_3089,N_4502);
xnor U9967 (N_9967,N_733,N_957);
nand U9968 (N_9968,N_1516,N_4292);
xor U9969 (N_9969,N_4346,N_1158);
or U9970 (N_9970,N_3529,N_2761);
or U9971 (N_9971,N_3397,N_2153);
nor U9972 (N_9972,N_11,N_3665);
nor U9973 (N_9973,N_4425,N_3152);
or U9974 (N_9974,N_276,N_1379);
and U9975 (N_9975,N_4651,N_3251);
xor U9976 (N_9976,N_4040,N_2551);
xnor U9977 (N_9977,N_2007,N_1475);
nor U9978 (N_9978,N_3559,N_3900);
and U9979 (N_9979,N_2328,N_2031);
nand U9980 (N_9980,N_2804,N_3700);
nor U9981 (N_9981,N_2822,N_4878);
nor U9982 (N_9982,N_26,N_273);
nand U9983 (N_9983,N_4446,N_4772);
nor U9984 (N_9984,N_714,N_3510);
and U9985 (N_9985,N_372,N_3770);
nor U9986 (N_9986,N_677,N_2596);
xor U9987 (N_9987,N_544,N_1191);
or U9988 (N_9988,N_3129,N_2982);
nor U9989 (N_9989,N_3871,N_2629);
and U9990 (N_9990,N_2907,N_1667);
xnor U9991 (N_9991,N_4937,N_4897);
or U9992 (N_9992,N_546,N_4460);
xor U9993 (N_9993,N_176,N_1882);
nor U9994 (N_9994,N_2051,N_4214);
nand U9995 (N_9995,N_1276,N_571);
or U9996 (N_9996,N_786,N_35);
nor U9997 (N_9997,N_3809,N_3149);
or U9998 (N_9998,N_385,N_200);
nand U9999 (N_9999,N_4301,N_1782);
and U10000 (N_10000,N_6990,N_9513);
or U10001 (N_10001,N_9972,N_5406);
nand U10002 (N_10002,N_6899,N_7187);
and U10003 (N_10003,N_9254,N_8662);
nand U10004 (N_10004,N_8910,N_9934);
nor U10005 (N_10005,N_8304,N_8594);
nand U10006 (N_10006,N_8463,N_7996);
or U10007 (N_10007,N_5950,N_8167);
nor U10008 (N_10008,N_6466,N_8113);
xnor U10009 (N_10009,N_6574,N_7451);
and U10010 (N_10010,N_7844,N_8558);
nand U10011 (N_10011,N_9383,N_6234);
xor U10012 (N_10012,N_6797,N_8582);
nand U10013 (N_10013,N_8494,N_5359);
and U10014 (N_10014,N_9275,N_6054);
nor U10015 (N_10015,N_8984,N_5333);
and U10016 (N_10016,N_8965,N_9241);
nand U10017 (N_10017,N_5530,N_5410);
nand U10018 (N_10018,N_7455,N_5450);
nand U10019 (N_10019,N_9425,N_9004);
nand U10020 (N_10020,N_5680,N_6471);
and U10021 (N_10021,N_6597,N_5768);
nand U10022 (N_10022,N_8520,N_9875);
xnor U10023 (N_10023,N_8367,N_8028);
xnor U10024 (N_10024,N_5673,N_8566);
nand U10025 (N_10025,N_8702,N_9252);
nor U10026 (N_10026,N_7832,N_5691);
xnor U10027 (N_10027,N_5546,N_6594);
nand U10028 (N_10028,N_9974,N_8243);
nor U10029 (N_10029,N_5755,N_9640);
and U10030 (N_10030,N_6892,N_7051);
nand U10031 (N_10031,N_5649,N_7034);
and U10032 (N_10032,N_5148,N_7108);
or U10033 (N_10033,N_7982,N_5064);
nand U10034 (N_10034,N_5591,N_6282);
nor U10035 (N_10035,N_7755,N_9825);
nand U10036 (N_10036,N_7714,N_5753);
nor U10037 (N_10037,N_7675,N_5794);
nand U10038 (N_10038,N_9551,N_9488);
or U10039 (N_10039,N_8715,N_8091);
or U10040 (N_10040,N_9466,N_9016);
nor U10041 (N_10041,N_8830,N_5675);
xnor U10042 (N_10042,N_5428,N_8901);
or U10043 (N_10043,N_7734,N_6329);
xnor U10044 (N_10044,N_6779,N_9651);
nor U10045 (N_10045,N_7517,N_6127);
xor U10046 (N_10046,N_6549,N_5026);
nor U10047 (N_10047,N_6739,N_8103);
and U10048 (N_10048,N_5809,N_6275);
nand U10049 (N_10049,N_8694,N_9322);
or U10050 (N_10050,N_8928,N_7364);
and U10051 (N_10051,N_7598,N_8477);
and U10052 (N_10052,N_6158,N_7251);
and U10053 (N_10053,N_8825,N_8992);
nand U10054 (N_10054,N_8302,N_9450);
nand U10055 (N_10055,N_8334,N_8378);
nand U10056 (N_10056,N_8711,N_5054);
and U10057 (N_10057,N_8400,N_7607);
xnor U10058 (N_10058,N_9007,N_8689);
or U10059 (N_10059,N_5391,N_6736);
xor U10060 (N_10060,N_6321,N_9802);
and U10061 (N_10061,N_6567,N_6408);
and U10062 (N_10062,N_5524,N_5004);
xnor U10063 (N_10063,N_7693,N_6979);
xnor U10064 (N_10064,N_7462,N_7708);
xor U10065 (N_10065,N_9618,N_5850);
nor U10066 (N_10066,N_9550,N_7204);
nor U10067 (N_10067,N_6188,N_9583);
xor U10068 (N_10068,N_5852,N_8050);
nor U10069 (N_10069,N_9721,N_7782);
xor U10070 (N_10070,N_7417,N_5412);
xnor U10071 (N_10071,N_5687,N_6871);
nor U10072 (N_10072,N_6418,N_8471);
xor U10073 (N_10073,N_9927,N_9514);
nor U10074 (N_10074,N_5408,N_7841);
and U10075 (N_10075,N_7669,N_6099);
or U10076 (N_10076,N_9088,N_8329);
nand U10077 (N_10077,N_7037,N_9922);
xnor U10078 (N_10078,N_6769,N_6897);
or U10079 (N_10079,N_5778,N_5287);
or U10080 (N_10080,N_5295,N_8282);
nand U10081 (N_10081,N_8426,N_7469);
and U10082 (N_10082,N_8253,N_8122);
nand U10083 (N_10083,N_6017,N_9462);
nand U10084 (N_10084,N_8062,N_8575);
xnor U10085 (N_10085,N_6117,N_8261);
nand U10086 (N_10086,N_7613,N_9365);
nor U10087 (N_10087,N_6236,N_9881);
nor U10088 (N_10088,N_5827,N_7423);
and U10089 (N_10089,N_7432,N_5678);
xor U10090 (N_10090,N_9108,N_9199);
xnor U10091 (N_10091,N_6636,N_5819);
nand U10092 (N_10092,N_9525,N_7765);
nor U10093 (N_10093,N_7837,N_5715);
and U10094 (N_10094,N_9384,N_8260);
xor U10095 (N_10095,N_5160,N_9848);
or U10096 (N_10096,N_6542,N_5919);
nand U10097 (N_10097,N_7622,N_5418);
nor U10098 (N_10098,N_8114,N_6124);
or U10099 (N_10099,N_9572,N_9696);
xor U10100 (N_10100,N_9484,N_5381);
nand U10101 (N_10101,N_5139,N_9459);
nor U10102 (N_10102,N_7929,N_8058);
nand U10103 (N_10103,N_7049,N_7788);
nor U10104 (N_10104,N_9478,N_5828);
and U10105 (N_10105,N_5003,N_7184);
nand U10106 (N_10106,N_8111,N_9768);
or U10107 (N_10107,N_5986,N_6679);
or U10108 (N_10108,N_6906,N_6625);
or U10109 (N_10109,N_7468,N_5149);
and U10110 (N_10110,N_5322,N_6762);
and U10111 (N_10111,N_6261,N_7316);
and U10112 (N_10112,N_6366,N_7602);
xor U10113 (N_10113,N_9142,N_9069);
nor U10114 (N_10114,N_8995,N_5871);
nor U10115 (N_10115,N_5757,N_6809);
nor U10116 (N_10116,N_5438,N_6505);
and U10117 (N_10117,N_5862,N_5093);
xnor U10118 (N_10118,N_9483,N_6307);
xor U10119 (N_10119,N_6123,N_7713);
or U10120 (N_10120,N_8423,N_5351);
nand U10121 (N_10121,N_5821,N_6239);
xnor U10122 (N_10122,N_6474,N_9127);
xor U10123 (N_10123,N_5383,N_5771);
nor U10124 (N_10124,N_5427,N_6498);
and U10125 (N_10125,N_5352,N_8456);
nand U10126 (N_10126,N_8262,N_6030);
nor U10127 (N_10127,N_7871,N_9853);
nor U10128 (N_10128,N_6641,N_7104);
xnor U10129 (N_10129,N_5329,N_6224);
nand U10130 (N_10130,N_8661,N_7609);
or U10131 (N_10131,N_9461,N_9884);
or U10132 (N_10132,N_9122,N_8972);
xnor U10133 (N_10133,N_5634,N_6079);
xor U10134 (N_10134,N_5196,N_9595);
nor U10135 (N_10135,N_6257,N_9697);
nand U10136 (N_10136,N_5700,N_6365);
nor U10137 (N_10137,N_5567,N_6805);
or U10138 (N_10138,N_9037,N_7939);
nand U10139 (N_10139,N_8223,N_5062);
or U10140 (N_10140,N_5595,N_5038);
or U10141 (N_10141,N_6345,N_9758);
nor U10142 (N_10142,N_6162,N_6431);
xor U10143 (N_10143,N_6951,N_7363);
xor U10144 (N_10144,N_6368,N_5811);
xnor U10145 (N_10145,N_8614,N_6263);
xor U10146 (N_10146,N_6849,N_5774);
nor U10147 (N_10147,N_7703,N_6080);
nor U10148 (N_10148,N_8770,N_8836);
and U10149 (N_10149,N_6798,N_5136);
nand U10150 (N_10150,N_5735,N_5937);
and U10151 (N_10151,N_5311,N_9346);
nor U10152 (N_10152,N_6443,N_6652);
or U10153 (N_10153,N_5244,N_6417);
nor U10154 (N_10154,N_5075,N_8299);
and U10155 (N_10155,N_5944,N_9440);
and U10156 (N_10156,N_9284,N_6037);
xor U10157 (N_10157,N_6572,N_6449);
nand U10158 (N_10158,N_5378,N_8930);
nor U10159 (N_10159,N_7698,N_5146);
nor U10160 (N_10160,N_6583,N_6435);
nand U10161 (N_10161,N_6294,N_8749);
or U10162 (N_10162,N_7560,N_6714);
nor U10163 (N_10163,N_5538,N_7088);
or U10164 (N_10164,N_7814,N_7087);
or U10165 (N_10165,N_8424,N_6580);
nand U10166 (N_10166,N_9617,N_9239);
nor U10167 (N_10167,N_6803,N_9098);
and U10168 (N_10168,N_7100,N_9059);
or U10169 (N_10169,N_5760,N_7071);
xnor U10170 (N_10170,N_8683,N_6202);
xor U10171 (N_10171,N_5155,N_6930);
and U10172 (N_10172,N_7769,N_7671);
xor U10173 (N_10173,N_8693,N_9585);
and U10174 (N_10174,N_5034,N_5293);
or U10175 (N_10175,N_7504,N_9285);
nand U10176 (N_10176,N_5888,N_8182);
xnor U10177 (N_10177,N_9702,N_7742);
nand U10178 (N_10178,N_9198,N_5480);
nand U10179 (N_10179,N_9442,N_6057);
nand U10180 (N_10180,N_5641,N_9055);
nor U10181 (N_10181,N_8977,N_7867);
or U10182 (N_10182,N_7717,N_6405);
nand U10183 (N_10183,N_5553,N_7011);
or U10184 (N_10184,N_5770,N_5371);
or U10185 (N_10185,N_8493,N_9282);
nor U10186 (N_10186,N_9887,N_6791);
xnor U10187 (N_10187,N_9081,N_6874);
or U10188 (N_10188,N_9178,N_5044);
nor U10189 (N_10189,N_9482,N_8840);
nand U10190 (N_10190,N_6947,N_6328);
and U10191 (N_10191,N_7330,N_5540);
or U10192 (N_10192,N_8917,N_8921);
xor U10193 (N_10193,N_7169,N_8875);
and U10194 (N_10194,N_8453,N_8331);
or U10195 (N_10195,N_9269,N_9872);
nand U10196 (N_10196,N_7284,N_5048);
nand U10197 (N_10197,N_9834,N_7321);
and U10198 (N_10198,N_8470,N_6869);
xnor U10199 (N_10199,N_9764,N_6469);
and U10200 (N_10200,N_6350,N_6961);
and U10201 (N_10201,N_8645,N_7311);
and U10202 (N_10202,N_5323,N_6976);
xor U10203 (N_10203,N_7440,N_9906);
xor U10204 (N_10204,N_7604,N_7747);
nor U10205 (N_10205,N_6831,N_7005);
nand U10206 (N_10206,N_8695,N_7259);
nand U10207 (N_10207,N_7157,N_9262);
xor U10208 (N_10208,N_5399,N_6393);
xor U10209 (N_10209,N_7375,N_7658);
nor U10210 (N_10210,N_9201,N_7620);
nor U10211 (N_10211,N_9729,N_9691);
and U10212 (N_10212,N_6318,N_6064);
nor U10213 (N_10213,N_7001,N_6219);
nor U10214 (N_10214,N_7345,N_7692);
xor U10215 (N_10215,N_9359,N_8443);
and U10216 (N_10216,N_9083,N_6663);
nand U10217 (N_10217,N_5379,N_9517);
nor U10218 (N_10218,N_9052,N_6260);
nor U10219 (N_10219,N_8742,N_7599);
or U10220 (N_10220,N_5242,N_5344);
nor U10221 (N_10221,N_8985,N_7524);
xor U10222 (N_10222,N_9772,N_7533);
nand U10223 (N_10223,N_5161,N_8462);
xnor U10224 (N_10224,N_6604,N_7502);
or U10225 (N_10225,N_8221,N_6903);
and U10226 (N_10226,N_6676,N_8069);
xnor U10227 (N_10227,N_8308,N_7979);
or U10228 (N_10228,N_6685,N_5968);
nand U10229 (N_10229,N_5125,N_9043);
nor U10230 (N_10230,N_8650,N_6948);
and U10231 (N_10231,N_9057,N_9784);
and U10232 (N_10232,N_5951,N_5665);
nor U10233 (N_10233,N_8633,N_6465);
and U10234 (N_10234,N_9920,N_9138);
xor U10235 (N_10235,N_5558,N_9975);
nor U10236 (N_10236,N_9472,N_7875);
nor U10237 (N_10237,N_8738,N_9362);
or U10238 (N_10238,N_6452,N_9711);
and U10239 (N_10239,N_7230,N_5599);
nor U10240 (N_10240,N_7722,N_7986);
or U10241 (N_10241,N_9349,N_7994);
or U10242 (N_10242,N_7276,N_7861);
and U10243 (N_10243,N_6927,N_7217);
nor U10244 (N_10244,N_9607,N_5957);
and U10245 (N_10245,N_5710,N_6729);
and U10246 (N_10246,N_8731,N_8599);
and U10247 (N_10247,N_7170,N_6422);
xor U10248 (N_10248,N_6727,N_9297);
or U10249 (N_10249,N_7195,N_7578);
and U10250 (N_10250,N_7799,N_6540);
nand U10251 (N_10251,N_8666,N_7803);
nor U10252 (N_10252,N_8580,N_9966);
xor U10253 (N_10253,N_6503,N_5049);
nor U10254 (N_10254,N_8796,N_8287);
nor U10255 (N_10255,N_6846,N_6657);
or U10256 (N_10256,N_5747,N_7800);
nand U10257 (N_10257,N_5101,N_8016);
or U10258 (N_10258,N_7020,N_9652);
xor U10259 (N_10259,N_8307,N_9712);
nor U10260 (N_10260,N_9996,N_8248);
or U10261 (N_10261,N_9794,N_6661);
nand U10262 (N_10262,N_8250,N_8532);
and U10263 (N_10263,N_8110,N_5928);
xor U10264 (N_10264,N_8318,N_5129);
and U10265 (N_10265,N_7296,N_8410);
xnor U10266 (N_10266,N_9842,N_7354);
nor U10267 (N_10267,N_6112,N_5625);
nor U10268 (N_10268,N_5086,N_7353);
or U10269 (N_10269,N_6154,N_6448);
or U10270 (N_10270,N_7357,N_8971);
xnor U10271 (N_10271,N_5415,N_7730);
nand U10272 (N_10272,N_7391,N_5973);
or U10273 (N_10273,N_7515,N_7780);
nand U10274 (N_10274,N_9333,N_7851);
xor U10275 (N_10275,N_5560,N_9502);
xor U10276 (N_10276,N_9412,N_5123);
nor U10277 (N_10277,N_5604,N_6886);
nor U10278 (N_10278,N_7485,N_5972);
xor U10279 (N_10279,N_6342,N_6140);
and U10280 (N_10280,N_6660,N_8912);
nand U10281 (N_10281,N_7074,N_8726);
xnor U10282 (N_10282,N_8322,N_5022);
and U10283 (N_10283,N_6792,N_6789);
xor U10284 (N_10284,N_5579,N_9646);
nand U10285 (N_10285,N_9181,N_7492);
nand U10286 (N_10286,N_6171,N_5395);
nor U10287 (N_10287,N_9791,N_7672);
or U10288 (N_10288,N_7829,N_9278);
or U10289 (N_10289,N_5452,N_9428);
nand U10290 (N_10290,N_6555,N_8806);
nor U10291 (N_10291,N_8822,N_5346);
xor U10292 (N_10292,N_9192,N_9167);
and U10293 (N_10293,N_9930,N_5298);
nor U10294 (N_10294,N_7210,N_6128);
xor U10295 (N_10295,N_5629,N_8154);
nor U10296 (N_10296,N_5615,N_7139);
xor U10297 (N_10297,N_5046,N_8397);
and U10298 (N_10298,N_7640,N_8120);
and U10299 (N_10299,N_8533,N_5009);
nand U10300 (N_10300,N_6967,N_6214);
xor U10301 (N_10301,N_5932,N_9800);
nor U10302 (N_10302,N_8979,N_9082);
or U10303 (N_10303,N_6599,N_5435);
nand U10304 (N_10304,N_5798,N_9866);
and U10305 (N_10305,N_5977,N_6168);
or U10306 (N_10306,N_8161,N_8712);
xnor U10307 (N_10307,N_9090,N_6426);
and U10308 (N_10308,N_7401,N_9206);
nor U10309 (N_10309,N_7807,N_5255);
nor U10310 (N_10310,N_9763,N_6339);
and U10311 (N_10311,N_6464,N_6493);
and U10312 (N_10312,N_7791,N_5921);
and U10313 (N_10313,N_9581,N_6069);
nor U10314 (N_10314,N_7854,N_5261);
xnor U10315 (N_10315,N_9248,N_7626);
nor U10316 (N_10316,N_7054,N_6222);
nor U10317 (N_10317,N_8510,N_6569);
xor U10318 (N_10318,N_9743,N_6723);
and U10319 (N_10319,N_7552,N_5721);
nor U10320 (N_10320,N_5580,N_8104);
or U10321 (N_10321,N_8046,N_6277);
xor U10322 (N_10322,N_7856,N_5555);
or U10323 (N_10323,N_6299,N_7924);
nor U10324 (N_10324,N_5947,N_6626);
nor U10325 (N_10325,N_8293,N_9695);
nand U10326 (N_10326,N_5441,N_7575);
xnor U10327 (N_10327,N_9542,N_8664);
nand U10328 (N_10328,N_5463,N_7315);
or U10329 (N_10329,N_5733,N_7762);
nor U10330 (N_10330,N_5751,N_8200);
or U10331 (N_10331,N_9809,N_5527);
or U10332 (N_10332,N_7431,N_7319);
xnor U10333 (N_10333,N_7294,N_8159);
nand U10334 (N_10334,N_9947,N_7787);
xor U10335 (N_10335,N_5117,N_7185);
nand U10336 (N_10336,N_8767,N_9154);
or U10337 (N_10337,N_8272,N_7885);
and U10338 (N_10338,N_9963,N_5204);
nor U10339 (N_10339,N_7751,N_8514);
or U10340 (N_10340,N_7110,N_9766);
nor U10341 (N_10341,N_5993,N_6244);
nand U10342 (N_10342,N_6889,N_9987);
nand U10343 (N_10343,N_7254,N_5754);
nor U10344 (N_10344,N_6119,N_7249);
nand U10345 (N_10345,N_7603,N_5095);
and U10346 (N_10346,N_7977,N_8136);
xnor U10347 (N_10347,N_9976,N_5313);
or U10348 (N_10348,N_7066,N_7082);
xor U10349 (N_10349,N_8679,N_5366);
and U10350 (N_10350,N_8829,N_8321);
nor U10351 (N_10351,N_5763,N_6519);
nand U10352 (N_10352,N_7715,N_5685);
or U10353 (N_10353,N_6494,N_8286);
nand U10354 (N_10354,N_8863,N_9399);
nor U10355 (N_10355,N_5787,N_9582);
xor U10356 (N_10356,N_8621,N_9878);
or U10357 (N_10357,N_8076,N_6880);
nor U10358 (N_10358,N_5780,N_6665);
nor U10359 (N_10359,N_6218,N_8482);
or U10360 (N_10360,N_9964,N_6781);
and U10361 (N_10361,N_7579,N_8503);
nor U10362 (N_10362,N_6609,N_5089);
and U10363 (N_10363,N_7749,N_9225);
nand U10364 (N_10364,N_7721,N_7687);
or U10365 (N_10365,N_6534,N_9431);
nor U10366 (N_10366,N_8399,N_8890);
and U10367 (N_10367,N_8506,N_8314);
or U10368 (N_10368,N_5534,N_7591);
xnor U10369 (N_10369,N_9505,N_5080);
nor U10370 (N_10370,N_7846,N_5069);
xor U10371 (N_10371,N_8049,N_6539);
xor U10372 (N_10372,N_9407,N_8414);
and U10373 (N_10373,N_8031,N_7916);
nand U10374 (N_10374,N_7244,N_7943);
xnor U10375 (N_10375,N_6851,N_9954);
or U10376 (N_10376,N_8512,N_6343);
or U10377 (N_10377,N_9161,N_6742);
nor U10378 (N_10378,N_6228,N_6308);
xor U10379 (N_10379,N_8359,N_8817);
xor U10380 (N_10380,N_9740,N_8475);
nor U10381 (N_10381,N_8156,N_8827);
xnor U10382 (N_10382,N_9056,N_7654);
xnor U10383 (N_10383,N_9329,N_8479);
or U10384 (N_10384,N_7189,N_5796);
nor U10385 (N_10385,N_5356,N_6738);
nand U10386 (N_10386,N_9408,N_5940);
or U10387 (N_10387,N_7221,N_8319);
or U10388 (N_10388,N_7477,N_9666);
xnor U10389 (N_10389,N_7080,N_8249);
or U10390 (N_10390,N_7618,N_9427);
nand U10391 (N_10391,N_5400,N_7739);
xor U10392 (N_10392,N_7368,N_9110);
and U10393 (N_10393,N_5677,N_5601);
and U10394 (N_10394,N_8570,N_7444);
xor U10395 (N_10395,N_6357,N_6490);
nor U10396 (N_10396,N_7608,N_6111);
nand U10397 (N_10397,N_5474,N_5752);
xnor U10398 (N_10398,N_8748,N_5788);
nand U10399 (N_10399,N_5559,N_6020);
xor U10400 (N_10400,N_8933,N_8908);
and U10401 (N_10401,N_6290,N_5725);
and U10402 (N_10402,N_7498,N_6845);
nor U10403 (N_10403,N_7014,N_6980);
nand U10404 (N_10404,N_8747,N_6866);
nor U10405 (N_10405,N_7981,N_9924);
and U10406 (N_10406,N_8017,N_9084);
and U10407 (N_10407,N_9435,N_7162);
nand U10408 (N_10408,N_5234,N_8184);
nor U10409 (N_10409,N_5726,N_6142);
nor U10410 (N_10410,N_7529,N_7968);
xor U10411 (N_10411,N_6115,N_8857);
nand U10412 (N_10412,N_7460,N_9971);
and U10413 (N_10413,N_5318,N_7834);
nand U10414 (N_10414,N_6481,N_7266);
and U10415 (N_10415,N_8531,N_9672);
and U10416 (N_10416,N_6701,N_9186);
nor U10417 (N_10417,N_5286,N_6761);
nor U10418 (N_10418,N_5238,N_5942);
or U10419 (N_10419,N_6454,N_5602);
nand U10420 (N_10420,N_8605,N_6457);
nor U10421 (N_10421,N_8343,N_7029);
xnor U10422 (N_10422,N_6850,N_5405);
or U10423 (N_10423,N_7526,N_9498);
nor U10424 (N_10424,N_6645,N_7932);
nor U10425 (N_10425,N_6149,N_9909);
xor U10426 (N_10426,N_9157,N_9632);
nor U10427 (N_10427,N_5609,N_9621);
nand U10428 (N_10428,N_7778,N_7246);
nand U10429 (N_10429,N_8981,N_5623);
xnor U10430 (N_10430,N_7313,N_7050);
nor U10431 (N_10431,N_6062,N_5392);
or U10432 (N_10432,N_9998,N_5698);
nand U10433 (N_10433,N_5954,N_9864);
nor U10434 (N_10434,N_7308,N_9242);
nor U10435 (N_10435,N_6658,N_9814);
and U10436 (N_10436,N_7196,N_5247);
and U10437 (N_10437,N_7150,N_6812);
or U10438 (N_10438,N_5390,N_8780);
nor U10439 (N_10439,N_9829,N_7232);
or U10440 (N_10440,N_7340,N_7253);
or U10441 (N_10441,N_6753,N_5817);
and U10442 (N_10442,N_9158,N_7137);
xor U10443 (N_10443,N_6700,N_9648);
or U10444 (N_10444,N_7828,N_5761);
or U10445 (N_10445,N_7325,N_8831);
xnor U10446 (N_10446,N_5734,N_5902);
and U10447 (N_10447,N_9737,N_6172);
or U10448 (N_10448,N_7773,N_5896);
nand U10449 (N_10449,N_7723,N_9641);
nand U10450 (N_10450,N_8276,N_8555);
nand U10451 (N_10451,N_5334,N_7464);
nor U10452 (N_10452,N_5657,N_7792);
nor U10453 (N_10453,N_6034,N_8360);
nor U10454 (N_10454,N_9313,N_8646);
xnor U10455 (N_10455,N_5158,N_9792);
nand U10456 (N_10456,N_8483,N_6501);
and U10457 (N_10457,N_8092,N_7306);
and U10458 (N_10458,N_7043,N_9446);
or U10459 (N_10459,N_5684,N_5923);
xor U10460 (N_10460,N_6447,N_6477);
nor U10461 (N_10461,N_5617,N_6994);
nand U10462 (N_10462,N_9576,N_9970);
and U10463 (N_10463,N_8931,N_7864);
xnor U10464 (N_10464,N_6790,N_8756);
nand U10465 (N_10465,N_7993,N_7877);
nand U10466 (N_10466,N_5007,N_5903);
nor U10467 (N_10467,N_5930,N_8192);
and U10468 (N_10468,N_8464,N_8497);
xor U10469 (N_10469,N_5099,N_7047);
nor U10470 (N_10470,N_6590,N_7384);
nand U10471 (N_10471,N_8821,N_6630);
nand U10472 (N_10472,N_5689,N_5631);
nor U10473 (N_10473,N_7655,N_8802);
or U10474 (N_10474,N_8824,N_9715);
nor U10475 (N_10475,N_7261,N_6024);
and U10476 (N_10476,N_9250,N_7868);
xnor U10477 (N_10477,N_8907,N_9174);
xnor U10478 (N_10478,N_9353,N_5036);
nor U10479 (N_10479,N_8498,N_8868);
nand U10480 (N_10480,N_9378,N_9799);
nand U10481 (N_10481,N_9591,N_7972);
and U10482 (N_10482,N_5504,N_8591);
xnor U10483 (N_10483,N_8030,N_7927);
nand U10484 (N_10484,N_7653,N_7203);
nor U10485 (N_10485,N_5398,N_9228);
or U10486 (N_10486,N_7165,N_5916);
nand U10487 (N_10487,N_6147,N_8925);
nand U10488 (N_10488,N_6153,N_6351);
nand U10489 (N_10489,N_8395,N_5597);
and U10490 (N_10490,N_6923,N_9544);
xor U10491 (N_10491,N_9166,N_9011);
xor U10492 (N_10492,N_8725,N_7328);
nand U10493 (N_10493,N_6944,N_7872);
or U10494 (N_10494,N_8081,N_9706);
nor U10495 (N_10495,N_6619,N_6073);
and U10496 (N_10496,N_7033,N_8187);
and U10497 (N_10497,N_8837,N_8980);
nor U10498 (N_10498,N_6843,N_6811);
nand U10499 (N_10499,N_6011,N_5370);
and U10500 (N_10500,N_6500,N_9893);
nand U10501 (N_10501,N_9936,N_6995);
nor U10502 (N_10502,N_5516,N_9050);
xnor U10503 (N_10503,N_8727,N_6386);
or U10504 (N_10504,N_5575,N_9149);
and U10505 (N_10505,N_5777,N_6303);
nor U10506 (N_10506,N_8189,N_6361);
nor U10507 (N_10507,N_9735,N_7124);
and U10508 (N_10508,N_8732,N_7397);
and U10509 (N_10509,N_9557,N_8766);
nor U10510 (N_10510,N_7081,N_7012);
xor U10511 (N_10511,N_5533,N_6433);
or U10512 (N_10512,N_7295,N_6411);
or U10513 (N_10513,N_6576,N_7659);
xor U10514 (N_10514,N_9000,N_6820);
nand U10515 (N_10515,N_6561,N_6400);
or U10516 (N_10516,N_8765,N_6352);
xnor U10517 (N_10517,N_8660,N_5728);
or U10518 (N_10518,N_8363,N_7003);
nor U10519 (N_10519,N_5468,N_6056);
or U10520 (N_10520,N_6830,N_9703);
nor U10521 (N_10521,N_8900,N_8613);
nand U10522 (N_10522,N_8958,N_7269);
and U10523 (N_10523,N_6362,N_6175);
nand U10524 (N_10524,N_5718,N_7992);
and U10525 (N_10525,N_5494,N_9840);
and U10526 (N_10526,N_7987,N_8859);
and U10527 (N_10527,N_5459,N_7534);
and U10528 (N_10528,N_5838,N_5193);
or U10529 (N_10529,N_7478,N_6806);
or U10530 (N_10530,N_6196,N_7369);
nor U10531 (N_10531,N_7912,N_6833);
nand U10532 (N_10532,N_7007,N_8415);
nand U10533 (N_10533,N_9801,N_7645);
or U10534 (N_10534,N_7951,N_6957);
and U10535 (N_10535,N_5076,N_6863);
nor U10536 (N_10536,N_9913,N_8590);
nand U10537 (N_10537,N_5090,N_9555);
or U10538 (N_10538,N_5249,N_5457);
or U10539 (N_10539,N_8568,N_8604);
nand U10540 (N_10540,N_5606,N_5207);
nand U10541 (N_10541,N_9476,N_5727);
xor U10542 (N_10542,N_9657,N_8133);
or U10543 (N_10543,N_9837,N_6637);
or U10544 (N_10544,N_5339,N_8425);
nand U10545 (N_10545,N_9810,N_8437);
and U10546 (N_10546,N_6415,N_8074);
nor U10547 (N_10547,N_7896,N_6682);
nor U10548 (N_10548,N_7733,N_9519);
or U10549 (N_10549,N_7663,N_8362);
nand U10550 (N_10550,N_5268,N_5327);
nor U10551 (N_10551,N_6675,N_7969);
and U10552 (N_10552,N_6712,N_9622);
and U10553 (N_10553,N_5825,N_5823);
and U10554 (N_10554,N_7078,N_9347);
nor U10555 (N_10555,N_9527,N_6004);
xnor U10556 (N_10556,N_9155,N_7129);
nand U10557 (N_10557,N_5859,N_8139);
and U10558 (N_10558,N_7719,N_7145);
nand U10559 (N_10559,N_9479,N_7320);
nor U10560 (N_10560,N_9079,N_7022);
nand U10561 (N_10561,N_8898,N_5302);
nand U10562 (N_10562,N_6243,N_8034);
nand U10563 (N_10563,N_7903,N_6216);
nand U10564 (N_10564,N_6799,N_6429);
xor U10565 (N_10565,N_6821,N_6287);
or U10566 (N_10566,N_5021,N_9653);
xnor U10567 (N_10567,N_8953,N_5775);
and U10568 (N_10568,N_9330,N_7274);
xnor U10569 (N_10569,N_5653,N_6265);
or U10570 (N_10570,N_5984,N_9833);
xnor U10571 (N_10571,N_8783,N_6536);
xnor U10572 (N_10572,N_8936,N_9164);
nand U10573 (N_10573,N_9245,N_5294);
nor U10574 (N_10574,N_8504,N_7167);
xor U10575 (N_10575,N_9116,N_5107);
xnor U10576 (N_10576,N_7105,N_5023);
xnor U10577 (N_10577,N_7745,N_7756);
and U10578 (N_10578,N_5372,N_8405);
xnor U10579 (N_10579,N_8145,N_8181);
nor U10580 (N_10580,N_7427,N_9309);
nand U10581 (N_10581,N_5460,N_7997);
nand U10582 (N_10582,N_5594,N_6817);
nand U10583 (N_10583,N_7116,N_8587);
xor U10584 (N_10584,N_7213,N_5834);
nand U10585 (N_10585,N_8768,N_8106);
xnor U10586 (N_10586,N_6130,N_8067);
or U10587 (N_10587,N_6673,N_9301);
or U10588 (N_10588,N_8722,N_8078);
nand U10589 (N_10589,N_6136,N_9403);
and U10590 (N_10590,N_7664,N_7786);
nand U10591 (N_10591,N_5522,N_9021);
nor U10592 (N_10592,N_5218,N_5425);
xnor U10593 (N_10593,N_6550,N_8881);
xor U10594 (N_10594,N_9229,N_7666);
nand U10595 (N_10595,N_7843,N_8450);
nand U10596 (N_10596,N_9685,N_6022);
and U10597 (N_10597,N_6562,N_6725);
and U10598 (N_10598,N_8801,N_6053);
nor U10599 (N_10599,N_8295,N_5472);
xor U10600 (N_10600,N_8847,N_5510);
nand U10601 (N_10601,N_7048,N_9549);
nand U10602 (N_10602,N_6211,N_5039);
xor U10603 (N_10603,N_8372,N_9759);
nor U10604 (N_10604,N_7257,N_8119);
nand U10605 (N_10605,N_5134,N_7839);
or U10606 (N_10606,N_9921,N_5866);
xnor U10607 (N_10607,N_9728,N_9426);
nor U10608 (N_10608,N_6006,N_9500);
nor U10609 (N_10609,N_6882,N_7271);
or U10610 (N_10610,N_9854,N_6522);
and U10611 (N_10611,N_8563,N_6425);
xor U10612 (N_10612,N_6483,N_5776);
nor U10613 (N_10613,N_9289,N_5731);
nor U10614 (N_10614,N_9841,N_9417);
or U10615 (N_10615,N_9633,N_5854);
and U10616 (N_10616,N_8220,N_6164);
nor U10617 (N_10617,N_7936,N_9969);
nand U10618 (N_10618,N_6424,N_7874);
or U10619 (N_10619,N_6659,N_7775);
or U10620 (N_10620,N_7949,N_8115);
or U10621 (N_10621,N_5439,N_9713);
nor U10622 (N_10622,N_7118,N_5240);
nand U10623 (N_10623,N_5458,N_7267);
xor U10624 (N_10624,N_5103,N_6063);
or U10625 (N_10625,N_9961,N_7920);
xor U10626 (N_10626,N_8354,N_8196);
nand U10627 (N_10627,N_9624,N_7428);
nor U10628 (N_10628,N_6516,N_8888);
and U10629 (N_10629,N_8976,N_9571);
and U10630 (N_10630,N_9175,N_8773);
nor U10631 (N_10631,N_6381,N_8126);
xnor U10632 (N_10632,N_9038,N_7009);
or U10633 (N_10633,N_8006,N_9942);
and U10634 (N_10634,N_5956,N_9400);
nor U10635 (N_10635,N_9001,N_9148);
nand U10636 (N_10636,N_5486,N_5363);
nor U10637 (N_10637,N_7387,N_7476);
and U10638 (N_10638,N_6807,N_5844);
xnor U10639 (N_10639,N_8518,N_9700);
or U10640 (N_10640,N_6841,N_9546);
or U10641 (N_10641,N_8403,N_7899);
xor U10642 (N_10642,N_9343,N_6414);
or U10643 (N_10643,N_5676,N_7774);
xnor U10644 (N_10644,N_5521,N_8446);
xor U10645 (N_10645,N_9773,N_5652);
nand U10646 (N_10646,N_8883,N_8609);
xor U10647 (N_10647,N_8713,N_7278);
and U10648 (N_10648,N_7676,N_6476);
and U10649 (N_10649,N_5264,N_6822);
or U10650 (N_10650,N_7435,N_5310);
nand U10651 (N_10651,N_7053,N_7439);
xnor U10652 (N_10652,N_6302,N_9770);
nor U10653 (N_10653,N_6598,N_5648);
xnor U10654 (N_10654,N_9890,N_8603);
xnor U10655 (N_10655,N_9986,N_6826);
nand U10656 (N_10656,N_8355,N_8164);
nor U10657 (N_10657,N_9778,N_8037);
nand U10658 (N_10658,N_9993,N_7231);
or U10659 (N_10659,N_9588,N_5904);
nor U10660 (N_10660,N_7283,N_5782);
nand U10661 (N_10661,N_5835,N_6853);
xnor U10662 (N_10662,N_7699,N_9797);
and U10663 (N_10663,N_8999,N_6012);
and U10664 (N_10664,N_5971,N_7390);
xor U10665 (N_10665,N_8779,N_5144);
xor U10666 (N_10666,N_5476,N_5960);
xor U10667 (N_10667,N_8778,N_9047);
xnor U10668 (N_10668,N_6942,N_6419);
nand U10669 (N_10669,N_5863,N_6316);
and U10670 (N_10670,N_5385,N_6177);
xnor U10671 (N_10671,N_7045,N_9009);
nor U10672 (N_10672,N_9029,N_5630);
nand U10673 (N_10673,N_8598,N_9465);
nand U10674 (N_10674,N_9689,N_8330);
or U10675 (N_10675,N_8368,N_9604);
nor U10676 (N_10676,N_9674,N_7706);
or U10677 (N_10677,N_5226,N_5679);
nor U10678 (N_10678,N_9506,N_6751);
or U10679 (N_10679,N_6108,N_7650);
and U10680 (N_10680,N_6907,N_8218);
xnor U10681 (N_10681,N_6910,N_7548);
or U10682 (N_10682,N_7612,N_9153);
nor U10683 (N_10683,N_6704,N_8897);
nand U10684 (N_10684,N_8624,N_6941);
nor U10685 (N_10685,N_8960,N_7120);
nor U10686 (N_10686,N_6992,N_7901);
or U10687 (N_10687,N_5925,N_5176);
nor U10688 (N_10688,N_8648,N_8775);
or U10689 (N_10689,N_8860,N_6377);
and U10690 (N_10690,N_7568,N_8927);
or U10691 (N_10691,N_5513,N_8002);
xnor U10692 (N_10692,N_8233,N_9813);
xnor U10693 (N_10693,N_6728,N_8672);
and U10694 (N_10694,N_8916,N_7940);
nor U10695 (N_10695,N_9644,N_7557);
and U10696 (N_10696,N_7701,N_9304);
and U10697 (N_10697,N_6526,N_9879);
nand U10698 (N_10698,N_7947,N_8585);
or U10699 (N_10699,N_9540,N_8361);
nor U10700 (N_10700,N_7509,N_9123);
nor U10701 (N_10701,N_9917,N_8391);
nor U10702 (N_10702,N_7662,N_8791);
or U10703 (N_10703,N_6122,N_9600);
and U10704 (N_10704,N_8215,N_9789);
xnor U10705 (N_10705,N_8404,N_5303);
xor U10706 (N_10706,N_9553,N_5868);
or U10707 (N_10707,N_9196,N_7093);
nor U10708 (N_10708,N_9914,N_6868);
xnor U10709 (N_10709,N_5804,N_9860);
nor U10710 (N_10710,N_7988,N_6199);
xor U10711 (N_10711,N_5490,N_8079);
and U10712 (N_10712,N_9738,N_9298);
or U10713 (N_10713,N_6566,N_5880);
xnor U10714 (N_10714,N_7911,N_5605);
xnor U10715 (N_10715,N_6283,N_8107);
nor U10716 (N_10716,N_6491,N_7378);
and U10717 (N_10717,N_8094,N_8014);
or U10718 (N_10718,N_5100,N_7490);
xor U10719 (N_10719,N_8753,N_5583);
xor U10720 (N_10720,N_5055,N_5669);
nor U10721 (N_10721,N_8990,N_5481);
and U10722 (N_10722,N_9410,N_9256);
and U10723 (N_10723,N_6655,N_8290);
nor U10724 (N_10724,N_6819,N_6146);
or U10725 (N_10725,N_6687,N_9070);
xnor U10726 (N_10726,N_6406,N_9965);
nor U10727 (N_10727,N_9005,N_9623);
and U10728 (N_10728,N_5495,N_7282);
or U10729 (N_10729,N_7121,N_8312);
nand U10730 (N_10730,N_8961,N_7349);
nand U10731 (N_10731,N_7408,N_9402);
or U10732 (N_10732,N_6060,N_5403);
or U10733 (N_10733,N_5169,N_6091);
or U10734 (N_10734,N_9786,N_6487);
nand U10735 (N_10735,N_7647,N_6949);
xor U10736 (N_10736,N_6775,N_6832);
nor U10737 (N_10737,N_6286,N_9288);
xor U10738 (N_10738,N_8441,N_7592);
and U10739 (N_10739,N_5404,N_9820);
or U10740 (N_10740,N_6925,N_8636);
xor U10741 (N_10741,N_9099,N_7026);
nor U10742 (N_10742,N_8593,N_6757);
or U10743 (N_10743,N_8724,N_9704);
nand U10744 (N_10744,N_6026,N_8994);
and U10745 (N_10745,N_7824,N_6148);
or U10746 (N_10746,N_8864,N_8365);
nand U10747 (N_10747,N_9337,N_5389);
nand U10748 (N_10748,N_6702,N_7342);
or U10749 (N_10749,N_6573,N_5536);
or U10750 (N_10750,N_8257,N_6276);
or U10751 (N_10751,N_8134,N_7225);
nand U10752 (N_10752,N_8627,N_8584);
nand U10753 (N_10753,N_9030,N_7380);
xnor U10754 (N_10754,N_6195,N_5975);
or U10755 (N_10755,N_8099,N_6186);
and U10756 (N_10756,N_6066,N_5939);
nand U10757 (N_10757,N_9128,N_5066);
and U10758 (N_10758,N_5257,N_5189);
nand U10759 (N_10759,N_8515,N_8112);
xor U10760 (N_10760,N_8799,N_7802);
nand U10761 (N_10761,N_9661,N_8377);
xnor U10762 (N_10762,N_7247,N_6489);
nor U10763 (N_10763,N_5229,N_5217);
nor U10764 (N_10764,N_5014,N_8600);
nor U10765 (N_10765,N_8655,N_5098);
xnor U10766 (N_10766,N_6297,N_9230);
or U10767 (N_10767,N_9223,N_9058);
or U10768 (N_10768,N_8042,N_7806);
and U10769 (N_10769,N_9326,N_5842);
nand U10770 (N_10770,N_6759,N_7711);
and U10771 (N_10771,N_5610,N_7057);
nand U10772 (N_10772,N_8059,N_7483);
and U10773 (N_10773,N_6268,N_8574);
nor U10774 (N_10774,N_7922,N_7928);
and U10775 (N_10775,N_5822,N_9422);
nor U10776 (N_10776,N_7860,N_5855);
nand U10777 (N_10777,N_6102,N_8970);
nand U10778 (N_10778,N_6755,N_8745);
or U10779 (N_10779,N_6315,N_5113);
and U10780 (N_10780,N_8708,N_8846);
xor U10781 (N_10781,N_7458,N_6964);
or U10782 (N_10782,N_6537,N_6392);
xor U10783 (N_10783,N_9503,N_8757);
or U10784 (N_10784,N_6086,N_5729);
or U10785 (N_10785,N_6628,N_8668);
nor U10786 (N_10786,N_9724,N_6732);
xnor U10787 (N_10787,N_9452,N_6279);
nand U10788 (N_10788,N_7630,N_8677);
and U10789 (N_10789,N_6467,N_7362);
nand U10790 (N_10790,N_6332,N_7373);
nor U10791 (N_10791,N_9932,N_6934);
nor U10792 (N_10792,N_8219,N_9949);
nor U10793 (N_10793,N_8744,N_9195);
xor U10794 (N_10794,N_7341,N_6028);
xnor U10795 (N_10795,N_5153,N_8044);
or U10796 (N_10796,N_5393,N_9547);
and U10797 (N_10797,N_8288,N_7983);
xnor U10798 (N_10798,N_7344,N_9017);
and U10799 (N_10799,N_6915,N_9526);
xor U10800 (N_10800,N_8168,N_8398);
or U10801 (N_10801,N_9036,N_7909);
nand U10802 (N_10802,N_5934,N_5265);
or U10803 (N_10803,N_6394,N_9566);
nand U10804 (N_10804,N_8567,N_6163);
or U10805 (N_10805,N_7409,N_5682);
xor U10806 (N_10806,N_8270,N_5712);
nor U10807 (N_10807,N_9790,N_7237);
nor U10808 (N_10808,N_7347,N_9573);
nor U10809 (N_10809,N_9575,N_8273);
nor U10810 (N_10810,N_9280,N_7097);
and U10811 (N_10811,N_9592,N_8394);
and U10812 (N_10812,N_9828,N_5965);
xor U10813 (N_10813,N_5998,N_5304);
or U10814 (N_10814,N_5328,N_5501);
nand U10815 (N_10815,N_5769,N_6450);
or U10816 (N_10816,N_6078,N_9111);
nand U10817 (N_10817,N_9504,N_5228);
or U10818 (N_10818,N_5477,N_8298);
xnor U10819 (N_10819,N_5614,N_7418);
nor U10820 (N_10820,N_5246,N_5664);
and U10821 (N_10821,N_7241,N_8969);
nand U10822 (N_10822,N_9628,N_8596);
nand U10823 (N_10823,N_8718,N_9350);
nand U10824 (N_10824,N_8628,N_5195);
xor U10825 (N_10825,N_5192,N_9855);
nand U10826 (N_10826,N_5814,N_8891);
xnor U10827 (N_10827,N_8607,N_5248);
and U10828 (N_10828,N_5805,N_7941);
xnor U10829 (N_10829,N_9586,N_8539);
or U10830 (N_10830,N_6227,N_9705);
or U10831 (N_10831,N_6437,N_6735);
and U10832 (N_10832,N_9281,N_7573);
or U10833 (N_10833,N_8246,N_5848);
xor U10834 (N_10834,N_5063,N_5430);
nor U10835 (N_10835,N_9769,N_5489);
xor U10836 (N_10836,N_8861,N_8686);
nor U10837 (N_10837,N_6106,N_6372);
nand U10838 (N_10838,N_8195,N_5083);
xor U10839 (N_10839,N_7683,N_6206);
nand U10840 (N_10840,N_6617,N_9665);
nor U10841 (N_10841,N_9742,N_9170);
nand U10842 (N_10842,N_6075,N_6093);
and U10843 (N_10843,N_5765,N_7503);
xnor U10844 (N_10844,N_5982,N_5622);
nor U10845 (N_10845,N_5523,N_7610);
or U10846 (N_10846,N_6475,N_5897);
and U10847 (N_10847,N_6565,N_9518);
and U10848 (N_10848,N_9593,N_9214);
nor U10849 (N_10849,N_7649,N_6747);
nand U10850 (N_10850,N_5453,N_8237);
nand U10851 (N_10851,N_6635,N_9977);
and U10852 (N_10852,N_5272,N_5988);
nand U10853 (N_10853,N_7790,N_5917);
nand U10854 (N_10854,N_5779,N_8935);
nor U10855 (N_10855,N_9392,N_5931);
or U10856 (N_10856,N_6204,N_6545);
nand U10857 (N_10857,N_7512,N_7226);
or U10858 (N_10858,N_9260,N_8294);
nor U10859 (N_10859,N_8040,N_8680);
and U10860 (N_10860,N_9815,N_9608);
and U10861 (N_10861,N_6622,N_9941);
or U10862 (N_10862,N_6051,N_8841);
xnor U10863 (N_10863,N_5618,N_5790);
or U10864 (N_10864,N_9699,N_8895);
or U10865 (N_10865,N_9257,N_7550);
nor U10866 (N_10866,N_5493,N_6159);
nor U10867 (N_10867,N_7808,N_5419);
xnor U10868 (N_10868,N_6407,N_8670);
xor U10869 (N_10869,N_5225,N_6932);
nor U10870 (N_10870,N_7168,N_6592);
xnor U10871 (N_10871,N_5588,N_5549);
nor U10872 (N_10872,N_5232,N_8205);
xor U10873 (N_10873,N_8162,N_5306);
or U10874 (N_10874,N_6748,N_5181);
xor U10875 (N_10875,N_5803,N_5396);
nor U10876 (N_10876,N_6320,N_5471);
xor U10877 (N_10877,N_8436,N_8941);
nor U10878 (N_10878,N_5291,N_8803);
or U10879 (N_10879,N_7190,N_7133);
or U10880 (N_10880,N_8467,N_9707);
and U10881 (N_10881,N_6325,N_8387);
nand U10882 (N_10882,N_8617,N_9434);
xnor U10883 (N_10883,N_7063,N_9308);
nor U10884 (N_10884,N_8269,N_9701);
or U10885 (N_10885,N_6298,N_8561);
nand U10886 (N_10886,N_5307,N_8056);
or U10887 (N_10887,N_8855,N_8835);
xor U10888 (N_10888,N_7297,N_8592);
and U10889 (N_10889,N_8379,N_9325);
and U10890 (N_10890,N_8902,N_8987);
nor U10891 (N_10891,N_6109,N_6480);
or U10892 (N_10892,N_8818,N_5152);
nor U10893 (N_10893,N_9804,N_9485);
and U10894 (N_10894,N_7119,N_7099);
or U10895 (N_10895,N_6848,N_5909);
nand U10896 (N_10896,N_7935,N_7265);
or U10897 (N_10897,N_9886,N_7700);
nand U10898 (N_10898,N_5767,N_6384);
nand U10899 (N_10899,N_8989,N_6269);
nand U10900 (N_10900,N_7955,N_7966);
xor U10901 (N_10901,N_6008,N_7900);
or U10902 (N_10902,N_5699,N_8486);
and U10903 (N_10903,N_5262,N_6065);
nor U10904 (N_10904,N_5537,N_6551);
and U10905 (N_10905,N_5147,N_8173);
xor U10906 (N_10906,N_8546,N_7600);
and U10907 (N_10907,N_6182,N_5651);
nand U10908 (N_10908,N_6602,N_7077);
nand U10909 (N_10909,N_5568,N_7198);
and U10910 (N_10910,N_5429,N_7978);
nand U10911 (N_10911,N_8588,N_5507);
or U10912 (N_10912,N_6289,N_9637);
xnor U10913 (N_10913,N_8022,N_9897);
and U10914 (N_10914,N_9568,N_7628);
xnor U10915 (N_10915,N_5282,N_9978);
nor U10916 (N_10916,N_7268,N_8944);
nand U10917 (N_10917,N_5661,N_6611);
and U10918 (N_10918,N_9190,N_5300);
or U10919 (N_10919,N_6281,N_9342);
or U10920 (N_10920,N_5843,N_9249);
and U10921 (N_10921,N_6674,N_9923);
and U10922 (N_10922,N_8513,N_5162);
and U10923 (N_10923,N_9183,N_6396);
and U10924 (N_10924,N_9356,N_9352);
xnor U10925 (N_10925,N_7377,N_6829);
and U10926 (N_10926,N_8306,N_7438);
xor U10927 (N_10927,N_9629,N_5343);
or U10928 (N_10928,N_9846,N_6586);
and U10929 (N_10929,N_7404,N_5110);
xnor U10930 (N_10930,N_7710,N_8488);
xor U10931 (N_10931,N_6690,N_6553);
or U10932 (N_10932,N_9765,N_8896);
nor U10933 (N_10933,N_5640,N_7566);
nor U10934 (N_10934,N_9220,N_9316);
nor U10935 (N_10935,N_9187,N_5382);
and U10936 (N_10936,N_7255,N_7690);
or U10937 (N_10937,N_8968,N_8597);
and U10938 (N_10938,N_5375,N_8833);
and U10939 (N_10939,N_7394,N_8808);
or U10940 (N_10940,N_6278,N_6232);
nor U10941 (N_10941,N_7753,N_8956);
or U10942 (N_10942,N_6300,N_5756);
xnor U10943 (N_10943,N_9670,N_5423);
or U10944 (N_10944,N_9447,N_5488);
or U10945 (N_10945,N_7386,N_9489);
or U10946 (N_10946,N_5883,N_5593);
nor U10947 (N_10947,N_5373,N_5266);
nand U10948 (N_10948,N_6970,N_9708);
xor U10949 (N_10949,N_9203,N_6322);
nand U10950 (N_10950,N_5933,N_9722);
nand U10951 (N_10951,N_8252,N_9634);
nor U10952 (N_10952,N_7164,N_7855);
xor U10953 (N_10953,N_6955,N_7897);
xnor U10954 (N_10954,N_8853,N_7359);
or U10955 (N_10955,N_6125,N_7836);
nand U10956 (N_10956,N_5898,N_8291);
and U10957 (N_10957,N_9638,N_5017);
or U10958 (N_10958,N_9339,N_6694);
nor U10959 (N_10959,N_7188,N_9045);
xnor U10960 (N_10960,N_7815,N_5467);
nor U10961 (N_10961,N_7131,N_7944);
nor U10962 (N_10962,N_5461,N_6556);
and U10963 (N_10963,N_9251,N_9344);
nor U10964 (N_10964,N_5227,N_7957);
or U10965 (N_10965,N_9687,N_5556);
or U10966 (N_10966,N_7095,N_6999);
nand U10967 (N_10967,N_8771,N_7991);
xor U10968 (N_10968,N_9276,N_9580);
or U10969 (N_10969,N_5209,N_9387);
nand U10970 (N_10970,N_9843,N_5672);
nand U10971 (N_10971,N_8224,N_5260);
or U10972 (N_10972,N_6003,N_6766);
and U10973 (N_10973,N_6780,N_7956);
or U10974 (N_10974,N_7889,N_8274);
xor U10975 (N_10975,N_7448,N_7665);
nand U10976 (N_10976,N_8812,N_7576);
or U10977 (N_10977,N_7400,N_5374);
nor U10978 (N_10978,N_7990,N_9404);
nand U10979 (N_10979,N_7332,N_7970);
and U10980 (N_10980,N_6035,N_9480);
or U10981 (N_10981,N_6528,N_8382);
and U10982 (N_10982,N_9374,N_8530);
or U10983 (N_10983,N_9601,N_6167);
or U10984 (N_10984,N_9681,N_6568);
or U10985 (N_10985,N_8721,N_7783);
nand U10986 (N_10986,N_5877,N_5040);
and U10987 (N_10987,N_8894,N_9130);
or U10988 (N_10988,N_9012,N_8750);
nor U10989 (N_10989,N_7399,N_9559);
xor U10990 (N_10990,N_6118,N_8186);
or U10991 (N_10991,N_9420,N_9124);
nand U10992 (N_10992,N_7835,N_8508);
and U10993 (N_10993,N_7472,N_8942);
and U10994 (N_10994,N_9054,N_9424);
or U10995 (N_10995,N_8373,N_6571);
or U10996 (N_10996,N_7547,N_5996);
xor U10997 (N_10997,N_6133,N_7302);
nand U10998 (N_10998,N_9443,N_6421);
xnor U10999 (N_10999,N_6001,N_5354);
and U11000 (N_11000,N_9380,N_5096);
nand U11001 (N_11001,N_5479,N_7553);
and U11002 (N_11002,N_5185,N_6643);
and U11003 (N_11003,N_6349,N_8844);
xor U11004 (N_11004,N_8032,N_5432);
nor U11005 (N_11005,N_7238,N_7372);
xor U11006 (N_11006,N_6143,N_6802);
nor U11007 (N_11007,N_8038,N_7823);
and U11008 (N_11008,N_8345,N_7805);
or U11009 (N_11009,N_5043,N_7263);
nand U11010 (N_11010,N_6559,N_7891);
xor U11011 (N_11011,N_9300,N_8647);
xor U11012 (N_11012,N_7967,N_5245);
nand U11013 (N_11013,N_9952,N_6391);
nand U11014 (N_11014,N_7256,N_6684);
nand U11015 (N_11015,N_8267,N_7046);
and U11016 (N_11016,N_9578,N_5860);
nor U11017 (N_11017,N_8213,N_5517);
or U11018 (N_11018,N_9097,N_9113);
or U11019 (N_11019,N_8946,N_8696);
or U11020 (N_11020,N_8129,N_9259);
xor U11021 (N_11021,N_9293,N_5231);
nor U11022 (N_11022,N_5578,N_5485);
nand U11023 (N_11023,N_8375,N_6782);
or U11024 (N_11024,N_7094,N_7309);
nor U11025 (N_11025,N_6633,N_5029);
and U11026 (N_11026,N_8913,N_9002);
nor U11027 (N_11027,N_6089,N_8551);
xnor U11028 (N_11028,N_8130,N_6885);
or U11029 (N_11029,N_6161,N_9224);
and U11030 (N_11030,N_5707,N_5317);
and U11031 (N_11031,N_7028,N_5345);
nor U11032 (N_11032,N_7729,N_5929);
nor U11033 (N_11033,N_8815,N_6914);
nand U11034 (N_11034,N_8204,N_5444);
and U11035 (N_11035,N_6249,N_5910);
and U11036 (N_11036,N_5639,N_8754);
nor U11037 (N_11037,N_6800,N_9822);
or U11038 (N_11038,N_5052,N_7716);
and U11039 (N_11039,N_5143,N_7661);
nor U11040 (N_11040,N_9667,N_7381);
nand U11041 (N_11041,N_6697,N_8141);
or U11042 (N_11042,N_7317,N_6061);
or U11043 (N_11043,N_8280,N_8320);
or U11044 (N_11044,N_9683,N_6412);
nand U11045 (N_11045,N_6962,N_8163);
or U11046 (N_11046,N_6824,N_6763);
nor U11047 (N_11047,N_7272,N_9014);
nand U11048 (N_11048,N_6401,N_5997);
nor U11049 (N_11049,N_6271,N_6966);
xor U11050 (N_11050,N_5283,N_5178);
nand U11051 (N_11051,N_8118,N_6554);
xor U11052 (N_11052,N_8255,N_8816);
nand U11053 (N_11053,N_6389,N_5926);
xnor U11054 (N_11054,N_5250,N_7127);
and U11055 (N_11055,N_5271,N_8199);
xnor U11056 (N_11056,N_9606,N_9244);
and U11057 (N_11057,N_5736,N_5171);
or U11058 (N_11058,N_7667,N_8612);
nor U11059 (N_11059,N_8877,N_8852);
nand U11060 (N_11060,N_8550,N_7627);
or U11061 (N_11061,N_6724,N_9415);
xor U11062 (N_11062,N_6884,N_8064);
xor U11063 (N_11063,N_9748,N_9419);
nand U11064 (N_11064,N_5908,N_5470);
or U11065 (N_11065,N_9753,N_7098);
nor U11066 (N_11066,N_9312,N_7822);
xnor U11067 (N_11067,N_9642,N_5469);
or U11068 (N_11068,N_6517,N_8073);
xnor U11069 (N_11069,N_8258,N_8547);
nor U11070 (N_11070,N_5424,N_9318);
nor U11071 (N_11071,N_5436,N_6786);
nand U11072 (N_11072,N_6973,N_9536);
nor U11073 (N_11073,N_5853,N_6027);
xnor U11074 (N_11074,N_7697,N_7010);
xor U11075 (N_11075,N_7580,N_5584);
nor U11076 (N_11076,N_9902,N_8704);
nand U11077 (N_11077,N_5890,N_7931);
nand U11078 (N_11078,N_5199,N_9093);
and U11079 (N_11079,N_9516,N_6496);
xor U11080 (N_11080,N_6672,N_6238);
nor U11081 (N_11081,N_9877,N_9876);
or U11082 (N_11082,N_8809,N_6521);
or U11083 (N_11083,N_9862,N_8552);
nand U11084 (N_11084,N_8554,N_7538);
nor U11085 (N_11085,N_9268,N_5886);
or U11086 (N_11086,N_5173,N_8328);
xnor U11087 (N_11087,N_6095,N_7030);
or U11088 (N_11088,N_9782,N_5577);
or U11089 (N_11089,N_7779,N_6306);
or U11090 (N_11090,N_6508,N_9752);
or U11091 (N_11091,N_5562,N_5270);
nor U11092 (N_11092,N_8843,N_6135);
xnor U11093 (N_11093,N_6603,N_7338);
nand U11094 (N_11094,N_5128,N_6312);
nor U11095 (N_11095,N_8915,N_7395);
nand U11096 (N_11096,N_9469,N_6067);
nand U11097 (N_11097,N_5208,N_6250);
nor U11098 (N_11098,N_9605,N_8740);
or U11099 (N_11099,N_7123,N_8481);
or U11100 (N_11100,N_5762,N_8461);
nor U11101 (N_11101,N_6353,N_8892);
xor U11102 (N_11102,N_9960,N_9105);
nor U11103 (N_11103,N_8878,N_6740);
and U11104 (N_11104,N_5607,N_7163);
xor U11105 (N_11105,N_8502,N_6883);
and U11106 (N_11106,N_6713,N_6670);
and U11107 (N_11107,N_6387,N_5223);
or U11108 (N_11108,N_8870,N_8828);
and U11109 (N_11109,N_7796,N_9775);
nand U11110 (N_11110,N_7572,N_8848);
or U11111 (N_11111,N_9287,N_7853);
nand U11112 (N_11112,N_5164,N_9912);
or U11113 (N_11113,N_6208,N_9078);
xor U11114 (N_11114,N_7677,N_8717);
xor U11115 (N_11115,N_8335,N_6327);
nor U11116 (N_11116,N_8451,N_8071);
nor U11117 (N_11117,N_5091,N_6081);
nor U11118 (N_11118,N_5188,N_9235);
nor U11119 (N_11119,N_5032,N_7136);
nor U11120 (N_11120,N_7199,N_7777);
and U11121 (N_11121,N_5550,N_9026);
nand U11122 (N_11122,N_5092,N_9125);
xor U11123 (N_11123,N_6646,N_5337);
nor U11124 (N_11124,N_6926,N_8658);
or U11125 (N_11125,N_5127,N_8940);
nand U11126 (N_11126,N_6169,N_9603);
nor U11127 (N_11127,N_9395,N_6499);
nor U11128 (N_11128,N_5620,N_7288);
or U11129 (N_11129,N_6292,N_6314);
or U11130 (N_11130,N_8336,N_8077);
nor U11131 (N_11131,N_5416,N_8346);
nor U11132 (N_11132,N_7724,N_9812);
or U11133 (N_11133,N_5024,N_6533);
xor U11134 (N_11134,N_7180,N_8667);
nand U11135 (N_11135,N_8408,N_9211);
or U11136 (N_11136,N_7801,N_8011);
xnor U11137 (N_11137,N_9218,N_6273);
and U11138 (N_11138,N_5420,N_8509);
nor U11139 (N_11139,N_9092,N_8549);
xnor U11140 (N_11140,N_9931,N_8311);
nand U11141 (N_11141,N_7292,N_5570);
nand U11142 (N_11142,N_8736,N_7567);
nor U11143 (N_11143,N_8341,N_9351);
nand U11144 (N_11144,N_7794,N_9615);
or U11145 (N_11145,N_5312,N_5554);
or U11146 (N_11146,N_7186,N_5349);
nor U11147 (N_11147,N_9838,N_5955);
nor U11148 (N_11148,N_5846,N_8013);
xnor U11149 (N_11149,N_9396,N_6705);
nor U11150 (N_11150,N_6986,N_8420);
xnor U11151 (N_11151,N_8865,N_9210);
and U11152 (N_11152,N_7726,N_9983);
and U11153 (N_11153,N_5511,N_5165);
nand U11154 (N_11154,N_7069,N_7334);
nor U11155 (N_11155,N_8385,N_5861);
nor U11156 (N_11156,N_8653,N_7999);
nor U11157 (N_11157,N_9627,N_6014);
xnor U11158 (N_11158,N_7816,N_7648);
nand U11159 (N_11159,N_7989,N_5781);
nand U11160 (N_11160,N_7243,N_9539);
xor U11161 (N_11161,N_7441,N_7343);
nand U11162 (N_11162,N_6103,N_7229);
or U11163 (N_11163,N_9747,N_7388);
nor U11164 (N_11164,N_7450,N_7463);
and U11165 (N_11165,N_7146,N_7245);
or U11166 (N_11166,N_9429,N_7507);
nor U11167 (N_11167,N_5276,N_7111);
nand U11168 (N_11168,N_7456,N_6319);
xnor U11169 (N_11169,N_6226,N_9331);
nor U11170 (N_11170,N_7605,N_8216);
or U11171 (N_11171,N_7277,N_5112);
or U11172 (N_11172,N_8885,N_8814);
nand U11173 (N_11173,N_6968,N_5845);
xnor U11174 (N_11174,N_5938,N_7374);
xor U11175 (N_11175,N_9205,N_5943);
xor U11176 (N_11176,N_5806,N_7784);
and U11177 (N_11177,N_5905,N_5981);
nand U11178 (N_11178,N_7952,N_8277);
nor U11179 (N_11179,N_9903,N_5350);
xnor U11180 (N_11180,N_9370,N_7679);
or U11181 (N_11181,N_6430,N_9077);
nand U11182 (N_11182,N_9231,N_7876);
or U11183 (N_11183,N_5839,N_7138);
and U11184 (N_11184,N_7273,N_7410);
or U11185 (N_11185,N_9796,N_9215);
or U11186 (N_11186,N_7651,N_8964);
nor U11187 (N_11187,N_8640,N_6180);
or U11188 (N_11188,N_6818,N_9354);
nor U11189 (N_11189,N_7153,N_7519);
xor U11190 (N_11190,N_7759,N_8642);
nand U11191 (N_11191,N_8782,N_9049);
or U11192 (N_11192,N_7696,N_7508);
nor U11193 (N_11193,N_6021,N_9611);
xnor U11194 (N_11194,N_8692,N_8084);
nand U11195 (N_11195,N_9911,N_8029);
nand U11196 (N_11196,N_6309,N_5239);
or U11197 (N_11197,N_8468,N_8759);
and U11198 (N_11198,N_6638,N_9957);
and U11199 (N_11199,N_7884,N_8789);
xnor U11200 (N_11200,N_7656,N_5157);
or U11201 (N_11201,N_9213,N_8432);
and U11202 (N_11202,N_7965,N_8348);
nor U11203 (N_11203,N_8967,N_9894);
nor U11204 (N_11204,N_5738,N_9531);
nand U11205 (N_11205,N_9861,N_5027);
or U11206 (N_11206,N_7379,N_8431);
or U11207 (N_11207,N_8544,N_8641);
or U11208 (N_11208,N_9369,N_9357);
nand U11209 (N_11209,N_7323,N_5279);
nor U11210 (N_11210,N_9491,N_5336);
xnor U11211 (N_11211,N_6141,N_6709);
nor U11212 (N_11212,N_6242,N_6872);
nand U11213 (N_11213,N_6246,N_5288);
xnor U11214 (N_11214,N_9184,N_6042);
nor U11215 (N_11215,N_9332,N_9982);
and U11216 (N_11216,N_6972,N_9345);
and U11217 (N_11217,N_9182,N_8795);
nor U11218 (N_11218,N_8409,N_8619);
xnor U11219 (N_11219,N_7910,N_5683);
nand U11220 (N_11220,N_7914,N_8871);
nand U11221 (N_11221,N_9662,N_8140);
nand U11222 (N_11222,N_6653,N_5499);
and U11223 (N_11223,N_8804,N_7818);
or U11224 (N_11224,N_6388,N_5131);
nor U11225 (N_11225,N_7718,N_6591);
nor U11226 (N_11226,N_8741,N_5596);
nand U11227 (N_11227,N_7632,N_9781);
xor U11228 (N_11228,N_5267,N_9880);
xnor U11229 (N_11229,N_7449,N_6960);
and U11230 (N_11230,N_6768,N_7545);
xor U11231 (N_11231,N_7385,N_7516);
nand U11232 (N_11232,N_7002,N_6774);
xor U11233 (N_11233,N_8241,N_8351);
nor U11234 (N_11234,N_9040,N_5870);
or U11235 (N_11235,N_7197,N_8606);
nor U11236 (N_11236,N_9507,N_6978);
nor U11237 (N_11237,N_5743,N_9534);
and U11238 (N_11238,N_9659,N_5137);
nand U11239 (N_11239,N_9754,N_6901);
or U11240 (N_11240,N_9680,N_7838);
xor U11241 (N_11241,N_7644,N_5627);
and U11242 (N_11242,N_8047,N_8838);
nand U11243 (N_11243,N_7421,N_7925);
and U11244 (N_11244,N_5115,N_7200);
nand U11245 (N_11245,N_8684,N_8430);
and U11246 (N_11246,N_7286,N_6823);
nand U11247 (N_11247,N_7122,N_6741);
nand U11248 (N_11248,N_6104,N_7581);
or U11249 (N_11249,N_8826,N_9398);
and U11250 (N_11250,N_5362,N_7532);
or U11251 (N_11251,N_5235,N_7072);
and U11252 (N_11252,N_5447,N_6010);
nand U11253 (N_11253,N_8781,N_9448);
xor U11254 (N_11254,N_5967,N_7454);
or U11255 (N_11255,N_5628,N_5674);
and U11256 (N_11256,N_8263,N_8500);
nand U11257 (N_11257,N_8411,N_6046);
and U11258 (N_11258,N_8637,N_8117);
and U11259 (N_11259,N_8849,N_9266);
nor U11260 (N_11260,N_7215,N_9314);
xnor U11261 (N_11261,N_6624,N_6201);
or U11262 (N_11262,N_6767,N_5475);
nand U11263 (N_11263,N_6876,N_7501);
or U11264 (N_11264,N_8873,N_5912);
xnor U11265 (N_11265,N_6511,N_9594);
xor U11266 (N_11266,N_8055,N_9112);
xnor U11267 (N_11267,N_8620,N_5791);
xor U11268 (N_11268,N_5658,N_8474);
and U11269 (N_11269,N_8611,N_9018);
and U11270 (N_11270,N_8762,N_6717);
or U11271 (N_11271,N_6255,N_8393);
and U11272 (N_11272,N_5316,N_6913);
nor U11273 (N_11273,N_7228,N_7337);
nand U11274 (N_11274,N_8185,N_8675);
or U11275 (N_11275,N_7549,N_6541);
and U11276 (N_11276,N_7985,N_6002);
or U11277 (N_11277,N_8635,N_9865);
nand U11278 (N_11278,N_9779,N_6369);
or U11279 (N_11279,N_7207,N_7242);
and U11280 (N_11280,N_5901,N_8786);
nor U11281 (N_11281,N_9538,N_8285);
or U11282 (N_11282,N_8438,N_9246);
xor U11283 (N_11283,N_9467,N_9523);
and U11284 (N_11284,N_5992,N_7625);
and U11285 (N_11285,N_8914,N_9327);
and U11286 (N_11286,N_7819,N_8934);
nand U11287 (N_11287,N_5251,N_6048);
nand U11288 (N_11288,N_9577,N_9216);
xnor U11289 (N_11289,N_5616,N_5646);
or U11290 (N_11290,N_9725,N_6203);
nor U11291 (N_11291,N_8095,N_8271);
nor U11292 (N_11292,N_5156,N_9944);
nand U11293 (N_11293,N_9335,N_5187);
nand U11294 (N_11294,N_5750,N_8823);
or U11295 (N_11295,N_7224,N_9719);
nor U11296 (N_11296,N_5686,N_7062);
xor U11297 (N_11297,N_8734,N_6495);
nand U11298 (N_11298,N_6212,N_9072);
nand U11299 (N_11299,N_5478,N_6423);
and U11300 (N_11300,N_8541,N_5011);
xor U11301 (N_11301,N_9454,N_7036);
or U11302 (N_11302,N_8242,N_9614);
and U11303 (N_11303,N_7820,N_7041);
xnor U11304 (N_11304,N_8595,N_6835);
xor U11305 (N_11305,N_8790,N_8540);
nand U11306 (N_11306,N_9371,N_8557);
and U11307 (N_11307,N_7938,N_9204);
xor U11308 (N_11308,N_8819,N_6059);
xor U11309 (N_11309,N_5719,N_5401);
xnor U11310 (N_11310,N_7959,N_8150);
nor U11311 (N_11311,N_6038,N_8376);
and U11312 (N_11312,N_7452,N_8303);
xor U11313 (N_11313,N_6808,N_5330);
or U11314 (N_11314,N_7056,N_7021);
and U11315 (N_11315,N_7420,N_5431);
nand U11316 (N_11316,N_9189,N_5057);
xnor U11317 (N_11317,N_8576,N_6529);
xor U11318 (N_11318,N_7426,N_9953);
nand U11319 (N_11319,N_5284,N_5966);
xnor U11320 (N_11320,N_5305,N_6587);
xor U11321 (N_11321,N_8492,N_6936);
nor U11322 (N_11322,N_8217,N_6094);
nor U11323 (N_11323,N_6058,N_8222);
xnor U11324 (N_11324,N_9915,N_6137);
xor U11325 (N_11325,N_5878,N_5571);
nand U11326 (N_11326,N_5613,N_8433);
or U11327 (N_11327,N_5301,N_5914);
or U11328 (N_11328,N_8703,N_8033);
or U11329 (N_11329,N_9598,N_6711);
or U11330 (N_11330,N_8615,N_6787);
nand U11331 (N_11331,N_5078,N_7830);
nor U11332 (N_11332,N_9867,N_7657);
and U11333 (N_11333,N_9140,N_5922);
nand U11334 (N_11334,N_6898,N_8374);
nor U11335 (N_11335,N_7013,N_5201);
nand U11336 (N_11336,N_7281,N_8206);
nand U11337 (N_11337,N_5849,N_7075);
nor U11338 (N_11338,N_6719,N_7770);
or U11339 (N_11339,N_7052,N_7845);
xnor U11340 (N_11340,N_5175,N_7058);
nand U11341 (N_11341,N_5409,N_8004);
or U11342 (N_11342,N_8457,N_8251);
nor U11343 (N_11343,N_6076,N_7106);
and U11344 (N_11344,N_5314,N_7586);
or U11345 (N_11345,N_8866,N_6492);
and U11346 (N_11346,N_8265,N_5918);
xor U11347 (N_11347,N_9221,N_5697);
nand U11348 (N_11348,N_7727,N_7304);
nand U11349 (N_11349,N_6049,N_7181);
or U11350 (N_11350,N_6221,N_6240);
nand U11351 (N_11351,N_9136,N_5873);
xnor U11352 (N_11352,N_9821,N_9366);
xnor U11353 (N_11353,N_9068,N_8279);
nand U11354 (N_11354,N_9874,N_5800);
or U11355 (N_11355,N_5473,N_7678);
nor U11356 (N_11356,N_7220,N_8296);
or U11357 (N_11357,N_5434,N_9761);
and U11358 (N_11358,N_8579,N_9172);
or U11359 (N_11359,N_5659,N_7360);
nor U11360 (N_11360,N_7101,N_6620);
nor U11361 (N_11361,N_7511,N_7746);
nor U11362 (N_11362,N_9073,N_7905);
or U11363 (N_11363,N_9202,N_6248);
and U11364 (N_11364,N_9323,N_6105);
and U11365 (N_11365,N_5668,N_9421);
or U11366 (N_11366,N_5884,N_7103);
xnor U11367 (N_11367,N_5881,N_5168);
nand U11368 (N_11368,N_5582,N_7291);
nand U11369 (N_11369,N_8190,N_7425);
xnor U11370 (N_11370,N_7280,N_7670);
or U11371 (N_11371,N_9334,N_8148);
nor U11372 (N_11372,N_8526,N_6678);
nor U11373 (N_11373,N_7500,N_6993);
and U11374 (N_11374,N_5927,N_8487);
or U11375 (N_11375,N_5421,N_6749);
xnor U11376 (N_11376,N_5455,N_9511);
and U11377 (N_11377,N_8324,N_5911);
nand U11378 (N_11378,N_5783,N_5241);
nand U11379 (N_11379,N_5109,N_8543);
xnor U11380 (N_11380,N_7083,N_8560);
nor U11381 (N_11381,N_9169,N_5047);
xor U11382 (N_11382,N_9449,N_9955);
nor U11383 (N_11383,N_6473,N_9609);
nor U11384 (N_11384,N_6756,N_5068);
and U11385 (N_11385,N_6828,N_7597);
nor U11386 (N_11386,N_9160,N_8203);
nand U11387 (N_11387,N_9264,N_6920);
and U11388 (N_11388,N_8009,N_8281);
nand U11389 (N_11389,N_6560,N_9321);
nor U11390 (N_11390,N_6547,N_5851);
xnor U11391 (N_11391,N_5042,N_8832);
and U11392 (N_11392,N_9967,N_8743);
nand U11393 (N_11393,N_6666,N_7327);
or U11394 (N_11394,N_7738,N_8674);
or U11395 (N_11395,N_7525,N_9959);
or U11396 (N_11396,N_5456,N_7857);
xor U11397 (N_11397,N_7488,N_9324);
xnor U11398 (N_11398,N_7998,N_5437);
and U11399 (N_11399,N_5633,N_6564);
nor U11400 (N_11400,N_6131,N_7530);
nor U11401 (N_11401,N_7582,N_9999);
xnor U11402 (N_11402,N_6929,N_5079);
nand U11403 (N_11403,N_9151,N_6814);
and U11404 (N_11404,N_6502,N_9562);
and U11405 (N_11405,N_8158,N_5941);
nand U11406 (N_11406,N_6341,N_8524);
nor U11407 (N_11407,N_6644,N_7827);
nor U11408 (N_11408,N_8292,N_8943);
xnor U11409 (N_11409,N_8700,N_8169);
nand U11410 (N_11410,N_9777,N_7660);
nand U11411 (N_11411,N_9095,N_9386);
or U11412 (N_11412,N_7833,N_6370);
xor U11413 (N_11413,N_7042,N_5151);
xor U11414 (N_11414,N_5041,N_6194);
nor U11415 (N_11415,N_7764,N_5621);
nand U11416 (N_11416,N_7125,N_9126);
or U11417 (N_11417,N_6839,N_7574);
nor U11418 (N_11418,N_8259,N_8651);
or U11419 (N_11419,N_5082,N_6771);
or U11420 (N_11420,N_5508,N_5174);
nand U11421 (N_11421,N_6378,N_9405);
nand U11422 (N_11422,N_5413,N_6259);
nor U11423 (N_11423,N_8959,N_9693);
or U11424 (N_11424,N_7352,N_6642);
nand U11425 (N_11425,N_6770,N_8511);
nand U11426 (N_11426,N_9745,N_6778);
and U11427 (N_11427,N_6760,N_6151);
or U11428 (N_11428,N_8983,N_8020);
or U11429 (N_11429,N_8349,N_6584);
nand U11430 (N_11430,N_9008,N_6904);
and U11431 (N_11431,N_6627,N_8063);
and U11432 (N_11432,N_9132,N_6862);
and U11433 (N_11433,N_9147,N_6340);
nand U11434 (N_11434,N_9232,N_9836);
nand U11435 (N_11435,N_7422,N_8876);
xnor U11436 (N_11436,N_8003,N_5565);
or U11437 (N_11437,N_5045,N_8157);
or U11438 (N_11438,N_6954,N_8323);
or U11439 (N_11439,N_6085,N_9945);
nor U11440 (N_11440,N_7482,N_6007);
and U11441 (N_11441,N_9537,N_8480);
or U11442 (N_11442,N_8236,N_6113);
and U11443 (N_11443,N_7351,N_8505);
xor U11444 (N_11444,N_8534,N_5206);
nor U11445 (N_11445,N_7637,N_6754);
nand U11446 (N_11446,N_6531,N_9682);
or U11447 (N_11447,N_5585,N_8101);
nor U11448 (N_11448,N_8991,N_6912);
nand U11449 (N_11449,N_9185,N_6173);
or U11450 (N_11450,N_5824,N_8998);
xnor U11451 (N_11451,N_8858,N_6453);
or U11452 (N_11452,N_6045,N_9520);
xnor U11453 (N_11453,N_7143,N_9973);
or U11454 (N_11454,N_6354,N_8097);
nor U11455 (N_11455,N_9451,N_5745);
nand U11456 (N_11456,N_8714,N_6854);
xor U11457 (N_11457,N_8144,N_9129);
nand U11458 (N_11458,N_8665,N_8854);
and U11459 (N_11459,N_8845,N_9564);
nor U11460 (N_11460,N_6185,N_7109);
xor U11461 (N_11461,N_8589,N_8525);
or U11462 (N_11462,N_7403,N_9492);
nor U11463 (N_11463,N_5820,N_6230);
xor U11464 (N_11464,N_7831,N_5644);
nand U11465 (N_11465,N_9569,N_6647);
nor U11466 (N_11466,N_7793,N_9937);
nand U11467 (N_11467,N_9100,N_5858);
xor U11468 (N_11468,N_7487,N_7016);
and U11469 (N_11469,N_7587,N_5840);
or U11470 (N_11470,N_9197,N_5913);
nor U11471 (N_11471,N_6997,N_9053);
or U11472 (N_11472,N_5978,N_5900);
nor U11473 (N_11473,N_7930,N_8562);
or U11474 (N_11474,N_5624,N_7405);
and U11475 (N_11475,N_6166,N_9490);
nor U11476 (N_11476,N_8673,N_7299);
nor U11477 (N_11477,N_8018,N_7092);
nand U11478 (N_11478,N_6677,N_5503);
xor U11479 (N_11479,N_9684,N_9328);
xor U11480 (N_11480,N_6088,N_5543);
xnor U11481 (N_11481,N_5670,N_5315);
or U11482 (N_11482,N_8706,N_7429);
and U11483 (N_11483,N_8485,N_8769);
xor U11484 (N_11484,N_8701,N_5072);
or U11485 (N_11485,N_8333,N_7642);
xnor U11486 (N_11486,N_5259,N_7883);
xnor U11487 (N_11487,N_6513,N_5230);
xor U11488 (N_11488,N_8639,N_8089);
or U11489 (N_11489,N_5028,N_7227);
and U11490 (N_11490,N_6070,N_5357);
and U11491 (N_11491,N_7740,N_5696);
nand U11492 (N_11492,N_7183,N_9716);
or U11493 (N_11493,N_8406,N_6486);
nand U11494 (N_11494,N_6585,N_5704);
nand U11495 (N_11495,N_8879,N_8950);
nand U11496 (N_11496,N_6348,N_9613);
nand U11497 (N_11497,N_8954,N_9234);
nand U11498 (N_11498,N_7518,N_6589);
and U11499 (N_11499,N_8625,N_5612);
nor U11500 (N_11500,N_9310,N_5407);
or U11501 (N_11501,N_7008,N_5205);
and U11502 (N_11502,N_5891,N_9677);
nor U11503 (N_11503,N_5526,N_5355);
nor U11504 (N_11504,N_9212,N_9438);
nand U11505 (N_11505,N_7735,N_5541);
xor U11506 (N_11506,N_9795,N_9686);
and U11507 (N_11507,N_7314,N_5764);
nor U11508 (N_11508,N_7239,N_9411);
and U11509 (N_11509,N_8000,N_8583);
nor U11510 (N_11510,N_7904,N_6145);
nand U11511 (N_11511,N_5116,N_7870);
and U11512 (N_11512,N_9720,N_7732);
xnor U11513 (N_11513,N_7817,N_5990);
or U11514 (N_11514,N_6293,N_5384);
nor U11515 (N_11515,N_9085,N_9731);
nand U11516 (N_11516,N_7826,N_9191);
and U11517 (N_11517,N_6258,N_8772);
nor U11518 (N_11518,N_8993,N_8152);
nand U11519 (N_11519,N_8962,N_7763);
or U11520 (N_11520,N_9746,N_5326);
nand U11521 (N_11521,N_7211,N_5915);
nand U11522 (N_11522,N_8339,N_9200);
or U11523 (N_11523,N_5140,N_9654);
xnor U11524 (N_11524,N_7117,N_8948);
nand U11525 (N_11525,N_8491,N_8325);
or U11526 (N_11526,N_6337,N_9545);
nor U11527 (N_11527,N_9240,N_6150);
nand U11528 (N_11528,N_9900,N_9401);
xor U11529 (N_11529,N_5708,N_5705);
or U11530 (N_11530,N_5183,N_9044);
or U11531 (N_11531,N_8342,N_5869);
or U11532 (N_11532,N_6785,N_5387);
and U11533 (N_11533,N_8978,N_6933);
xor U11534 (N_11534,N_8986,N_5320);
and U11535 (N_11535,N_6323,N_6864);
nand U11536 (N_11536,N_9830,N_5253);
xnor U11537 (N_11537,N_5269,N_9529);
nand U11538 (N_11538,N_9827,N_5104);
nor U11539 (N_11539,N_5342,N_8212);
nor U11540 (N_11540,N_5126,N_5974);
or U11541 (N_11541,N_5663,N_6442);
nand U11542 (N_11542,N_5018,N_5073);
nor U11543 (N_11543,N_7858,N_5812);
or U11544 (N_11544,N_5496,N_8039);
nand U11545 (N_11545,N_6247,N_5191);
and U11546 (N_11546,N_9475,N_5730);
nor U11547 (N_11547,N_6047,N_7067);
xnor U11548 (N_11548,N_9433,N_5275);
and U11549 (N_11549,N_5331,N_9658);
xnor U11550 (N_11550,N_5448,N_7402);
nor U11551 (N_11551,N_9859,N_5924);
xnor U11552 (N_11552,N_9663,N_8283);
xor U11553 (N_11553,N_7668,N_7555);
and U11554 (N_11554,N_8499,N_6656);
or U11555 (N_11555,N_9589,N_8146);
nor U11556 (N_11556,N_7065,N_5319);
nor U11557 (N_11557,N_9694,N_9512);
or U11558 (N_11558,N_8626,N_7760);
nand U11559 (N_11559,N_5525,N_7559);
or U11560 (N_11560,N_8155,N_7035);
or U11561 (N_11561,N_8904,N_9522);
or U11562 (N_11562,N_5019,N_7588);
xor U11563 (N_11563,N_8528,N_7382);
xnor U11564 (N_11564,N_8388,N_9709);
or U11565 (N_11565,N_9291,N_7863);
xnor U11566 (N_11566,N_7156,N_6364);
or U11567 (N_11567,N_7873,N_8787);
xor U11568 (N_11568,N_9080,N_6977);
xnor U11569 (N_11569,N_6688,N_8982);
or U11570 (N_11570,N_7584,N_9066);
nand U11571 (N_11571,N_8459,N_5722);
nand U11572 (N_11572,N_9750,N_9363);
and U11573 (N_11573,N_7300,N_5952);
xor U11574 (N_11574,N_5899,N_6708);
or U11575 (N_11575,N_5958,N_8015);
xnor U11576 (N_11576,N_9530,N_7771);
nor U11577 (N_11577,N_8472,N_8924);
nor U11578 (N_11578,N_5948,N_7570);
or U11579 (N_11579,N_8090,N_5120);
xnor U11580 (N_11580,N_9436,N_9109);
xor U11581 (N_11581,N_6827,N_8240);
nor U11582 (N_11582,N_6404,N_7497);
nand U11583 (N_11583,N_8764,N_6157);
xnor U11584 (N_11584,N_9430,N_7222);
xor U11585 (N_11585,N_8207,N_7556);
or U11586 (N_11586,N_5060,N_6891);
and U11587 (N_11587,N_7728,N_7652);
nor U11588 (N_11588,N_7443,N_6515);
or U11589 (N_11589,N_7091,N_5732);
xor U11590 (N_11590,N_9379,N_7144);
or U11591 (N_11591,N_8444,N_8428);
or U11592 (N_11592,N_7158,N_5882);
nor U11593 (N_11593,N_9710,N_7971);
or U11594 (N_11594,N_5216,N_8337);
nor U11595 (N_11595,N_8238,N_9296);
xnor U11596 (N_11596,N_6356,N_9916);
or U11597 (N_11597,N_7216,N_8997);
and U11598 (N_11598,N_8239,N_9762);
and U11599 (N_11599,N_7921,N_5987);
nor U11600 (N_11600,N_7480,N_6718);
xor U11601 (N_11601,N_6253,N_8402);
and U11602 (N_11602,N_8188,N_9532);
and U11603 (N_11603,N_5121,N_5364);
xor U11604 (N_11604,N_6859,N_8172);
nor U11605 (N_11605,N_5166,N_8228);
nand U11606 (N_11606,N_5273,N_5141);
nor U11607 (N_11607,N_7060,N_5563);
xor U11608 (N_11608,N_9741,N_9951);
xor U11609 (N_11609,N_6371,N_6908);
nand U11610 (N_11610,N_6497,N_8676);
xnor U11611 (N_11611,N_8065,N_5695);
nor U11612 (N_11612,N_7489,N_7505);
nor U11613 (N_11613,N_8193,N_6210);
nor U11614 (N_11614,N_9744,N_5365);
or U11615 (N_11615,N_7695,N_9493);
or U11616 (N_11616,N_5081,N_5889);
and U11617 (N_11617,N_8447,N_9882);
nand U11618 (N_11618,N_9515,N_9910);
nor U11619 (N_11619,N_8963,N_6579);
or U11620 (N_11620,N_6121,N_7061);
nor U11621 (N_11621,N_8973,N_9823);
or U11622 (N_11622,N_9338,N_8872);
nand U11623 (N_11623,N_9832,N_9788);
and U11624 (N_11624,N_9818,N_6975);
nor U11625 (N_11625,N_8147,N_5836);
and U11626 (N_11626,N_6654,N_7287);
and U11627 (N_11627,N_8538,N_7430);
or U11628 (N_11628,N_6945,N_7686);
nand U11629 (N_11629,N_6870,N_9432);
nor U11630 (N_11630,N_5529,N_5483);
nor U11631 (N_11631,N_7479,N_7707);
nor U11632 (N_11632,N_8465,N_9439);
or U11633 (N_11633,N_8974,N_5936);
and U11634 (N_11634,N_7177,N_9286);
xnor U11635 (N_11635,N_5243,N_8867);
or U11636 (N_11636,N_7895,N_8638);
xor U11637 (N_11637,N_6107,N_5368);
xnor U11638 (N_11638,N_5514,N_8682);
and U11639 (N_11639,N_6578,N_6825);
nand U11640 (N_11640,N_7038,N_8923);
nand U11641 (N_11641,N_7810,N_5020);
and U11642 (N_11642,N_9227,N_9025);
and U11643 (N_11643,N_9118,N_9381);
xnor U11644 (N_11644,N_5252,N_9258);
or U11645 (N_11645,N_5766,N_8102);
xnor U11646 (N_11646,N_6284,N_8171);
nor U11647 (N_11647,N_8842,N_8201);
nand U11648 (N_11648,N_6184,N_7289);
or U11649 (N_11649,N_9271,N_8390);
nand U11650 (N_11650,N_6374,N_9499);
or U11651 (N_11651,N_6613,N_7964);
xor U11652 (N_11652,N_9494,N_9565);
nor U11653 (N_11653,N_5949,N_6207);
or U11654 (N_11654,N_8527,N_7565);
and U11655 (N_11655,N_7161,N_7142);
or U11656 (N_11656,N_6110,N_5114);
nor U11657 (N_11657,N_9805,N_8903);
nand U11658 (N_11658,N_9134,N_9222);
xnor U11659 (N_11659,N_7862,N_7544);
and U11660 (N_11660,N_7235,N_8723);
nor U11661 (N_11661,N_9552,N_9933);
xnor U11662 (N_11662,N_5108,N_8517);
xnor U11663 (N_11663,N_5397,N_6847);
nand U11664 (N_11664,N_7219,N_8165);
nor U11665 (N_11665,N_9984,N_8383);
xnor U11666 (N_11666,N_9783,N_6860);
nor U11667 (N_11667,N_7486,N_7361);
nor U11668 (N_11668,N_7312,N_9377);
nor U11669 (N_11669,N_7209,N_6252);
xnor U11670 (N_11670,N_7290,N_7720);
or U11671 (N_11671,N_5236,N_8001);
xor U11672 (N_11672,N_8634,N_5502);
nor U11673 (N_11673,N_5792,N_6730);
and U11674 (N_11674,N_8366,N_7767);
or U11675 (N_11675,N_8108,N_5714);
xor U11676 (N_11676,N_6879,N_8911);
and U11677 (N_11677,N_6092,N_6295);
nor U11678 (N_11678,N_9535,N_7398);
xor U11679 (N_11679,N_8416,N_8211);
xnor U11680 (N_11680,N_9389,N_7346);
nor U11681 (N_11681,N_9306,N_9135);
and U11682 (N_11682,N_6581,N_6267);
nor U11683 (N_11683,N_7595,N_9528);
nand U11684 (N_11684,N_9760,N_6836);
and U11685 (N_11685,N_6877,N_5895);
nand U11686 (N_11686,N_9361,N_6538);
xor U11687 (N_11687,N_7906,N_5258);
nand U11688 (N_11688,N_5220,N_7089);
nand U11689 (N_11689,N_8266,N_7554);
nor U11690 (N_11690,N_8043,N_7453);
and U11691 (N_11691,N_7635,N_8776);
nor U11692 (N_11692,N_8553,N_6304);
nand U11693 (N_11693,N_8926,N_6535);
nand U11694 (N_11694,N_8618,N_5466);
and U11695 (N_11695,N_8788,N_7898);
nor U11696 (N_11696,N_7754,N_6187);
nor U11697 (N_11697,N_6570,N_7134);
nand U11698 (N_11698,N_6382,N_9042);
or U11699 (N_11699,N_9144,N_9367);
or U11700 (N_11700,N_9785,N_8685);
xnor U11701 (N_11701,N_7712,N_9487);
nor U11702 (N_11702,N_9751,N_7510);
nor U11703 (N_11703,N_9671,N_7888);
nor U11704 (N_11704,N_6527,N_9418);
or U11705 (N_11705,N_9883,N_7160);
or U11706 (N_11706,N_6225,N_7348);
and U11707 (N_11707,N_5667,N_9739);
and U11708 (N_11708,N_7437,N_8952);
nand U11709 (N_11709,N_5180,N_7059);
and U11710 (N_11710,N_6720,N_7850);
xnor U11711 (N_11711,N_9771,N_8194);
or U11712 (N_11712,N_7491,N_9032);
nand U11713 (N_11713,N_7339,N_7893);
and U11714 (N_11714,N_9888,N_5867);
nand U11715 (N_11715,N_6963,N_6596);
and U11716 (N_11716,N_7812,N_7915);
or U11717 (N_11717,N_7055,N_8777);
and U11718 (N_11718,N_7892,N_9277);
nor U11719 (N_11719,N_7471,N_7414);
xor U11720 (N_11720,N_6943,N_8586);
or U11721 (N_11721,N_5074,N_8025);
nand U11722 (N_11722,N_8202,N_7961);
and U11723 (N_11723,N_9341,N_7859);
or U11724 (N_11724,N_8792,N_5006);
or U11725 (N_11725,N_8235,N_7305);
xor U11726 (N_11726,N_8476,N_9819);
or U11727 (N_11727,N_7908,N_9690);
and U11728 (N_11728,N_7019,N_6922);
nand U11729 (N_11729,N_7621,N_7540);
and U11730 (N_11730,N_8834,N_8231);
xnor U11731 (N_11731,N_9020,N_5581);
nor U11732 (N_11732,N_9270,N_9639);
or U11733 (N_11733,N_5542,N_6441);
or U11734 (N_11734,N_9317,N_6152);
and U11735 (N_11735,N_5451,N_5388);
xnor U11736 (N_11736,N_7174,N_6928);
or U11737 (N_11737,N_8763,N_5071);
or U11738 (N_11738,N_6722,N_9087);
nor U11739 (N_11739,N_7590,N_6937);
and U11740 (N_11740,N_8501,N_8245);
and U11741 (N_11741,N_6601,N_7279);
and U11742 (N_11742,N_7942,N_6710);
nor U11743 (N_11743,N_8229,N_5010);
nor U11744 (N_11744,N_6706,N_6691);
and U11745 (N_11745,N_9265,N_5590);
nand U11746 (N_11746,N_9849,N_9950);
xor U11747 (N_11747,N_9048,N_6482);
xnor U11748 (N_11748,N_5816,N_5784);
xor U11749 (N_11749,N_9597,N_6272);
nor U11750 (N_11750,N_8690,N_8421);
xnor U11751 (N_11751,N_5841,N_9939);
and U11752 (N_11752,N_9273,N_6518);
and U11753 (N_11753,N_6470,N_9997);
nor U11754 (N_11754,N_9807,N_8739);
nand U11755 (N_11755,N_9217,N_6919);
nor U11756 (N_11756,N_7159,N_9899);
nor U11757 (N_11757,N_9806,N_7436);
nand U11758 (N_11758,N_9889,N_9107);
nor U11759 (N_11759,N_5449,N_5367);
nand U11760 (N_11760,N_7336,N_6514);
and U11761 (N_11761,N_5219,N_9464);
xnor U11762 (N_11762,N_8230,N_5801);
and U11763 (N_11763,N_5603,N_5280);
and U11764 (N_11764,N_9076,N_7457);
nand U11765 (N_11765,N_5662,N_9233);
nor U11766 (N_11766,N_7112,N_8209);
nor U11767 (N_11767,N_5094,N_9307);
xor U11768 (N_11768,N_5296,N_7205);
and U11769 (N_11769,N_7192,N_7980);
nor U11770 (N_11770,N_5737,N_6285);
xnor U11771 (N_11771,N_5492,N_8142);
or U11772 (N_11772,N_9019,N_9051);
nand U11773 (N_11773,N_7562,N_5031);
and U11774 (N_11774,N_7681,N_5688);
xor U11775 (N_11775,N_9590,N_9022);
nand U11776 (N_11776,N_7270,N_6331);
xor U11777 (N_11777,N_9460,N_9423);
nand U11778 (N_11778,N_5660,N_7393);
xor U11779 (N_11779,N_7615,N_8121);
or U11780 (N_11780,N_6071,N_7260);
nand U11781 (N_11781,N_9150,N_7171);
or U11782 (N_11782,N_5277,N_6631);
xor U11783 (N_11783,N_8197,N_6326);
nand U11784 (N_11784,N_6988,N_8256);
nor U11785 (N_11785,N_7673,N_9340);
xor U11786 (N_11786,N_8412,N_6623);
nor U11787 (N_11787,N_8315,N_5885);
xnor U11788 (N_11788,N_5445,N_7917);
nor U11789 (N_11789,N_6510,N_8309);
nand U11790 (N_11790,N_6120,N_5906);
nor U11791 (N_11791,N_8138,N_8310);
and U11792 (N_11792,N_5832,N_6446);
or U11793 (N_11793,N_8542,N_8137);
or U11794 (N_11794,N_5353,N_6616);
xnor U11795 (N_11795,N_9453,N_6023);
or U11796 (N_11796,N_9612,N_5059);
nor U11797 (N_11797,N_8737,N_6629);
or U11798 (N_11798,N_5587,N_6036);
and U11799 (N_11799,N_7593,N_7015);
or U11800 (N_11800,N_5186,N_8254);
and U11801 (N_11801,N_5723,N_7960);
nor U11802 (N_11802,N_8007,N_9858);
nand U11803 (N_11803,N_7954,N_8455);
nor U11804 (N_11804,N_9458,N_6181);
and U11805 (N_11805,N_7396,N_5772);
or U11806 (N_11806,N_7214,N_8807);
nor U11807 (N_11807,N_8716,N_9063);
or U11808 (N_11808,N_5053,N_5084);
nand U11809 (N_11809,N_5324,N_7772);
and U11810 (N_11810,N_9556,N_7705);
or U11811 (N_11811,N_7809,N_7149);
and U11812 (N_11812,N_6460,N_5773);
or U11813 (N_11813,N_9631,N_7212);
nand U11814 (N_11814,N_5532,N_7535);
and U11815 (N_11815,N_5465,N_7629);
and U11816 (N_11816,N_8301,N_9477);
and U11817 (N_11817,N_7933,N_8851);
nor U11818 (N_11818,N_5105,N_7191);
xor U11819 (N_11819,N_8988,N_5030);
xnor U11820 (N_11820,N_5215,N_6548);
nor U11821 (N_11821,N_7132,N_9988);
nor U11822 (N_11822,N_7293,N_7234);
or U11823 (N_11823,N_7811,N_6402);
nand U11824 (N_11824,N_9956,N_7018);
and U11825 (N_11825,N_5785,N_6179);
and U11826 (N_11826,N_9247,N_7882);
nand U11827 (N_11827,N_6745,N_9626);
nor U11828 (N_11828,N_9625,N_6176);
or U11829 (N_11829,N_9630,N_5237);
xor U11830 (N_11830,N_5874,N_5341);
or U11831 (N_11831,N_5491,N_9064);
xnor U11832 (N_11832,N_6543,N_6810);
and U11833 (N_11833,N_8371,N_7583);
xor U11834 (N_11834,N_8036,N_5589);
or U11835 (N_11835,N_7193,N_9119);
xnor U11836 (N_11836,N_7493,N_9146);
xor U11837 (N_11837,N_6618,N_8350);
nor U11838 (N_11838,N_5557,N_9413);
nor U11839 (N_11839,N_7750,N_8051);
xnor U11840 (N_11840,N_6347,N_6335);
nand U11841 (N_11841,N_5308,N_7358);
nor U11842 (N_11842,N_7333,N_8733);
xor U11843 (N_11843,N_9089,N_6733);
xor U11844 (N_11844,N_8573,N_6040);
nor U11845 (N_11845,N_6715,N_9871);
and U11846 (N_11846,N_8066,N_5626);
xor U11847 (N_11847,N_9115,N_7096);
xnor U11848 (N_11848,N_7520,N_7461);
nor U11849 (N_11849,N_8632,N_9533);
nor U11850 (N_11850,N_5711,N_6134);
or U11851 (N_11851,N_8906,N_9676);
xor U11852 (N_11852,N_7631,N_9141);
or U11853 (N_11853,N_8919,N_6544);
nand U11854 (N_11854,N_8024,N_8234);
xor U11855 (N_11855,N_7371,N_8082);
nand U11856 (N_11856,N_9567,N_6015);
or U11857 (N_11857,N_8338,N_6274);
and U11858 (N_11858,N_5656,N_5097);
and U11859 (N_11859,N_6612,N_5289);
or U11860 (N_11860,N_8671,N_7389);
nand U11861 (N_11861,N_6777,N_5000);
xnor U11862 (N_11862,N_5647,N_5213);
nand U11863 (N_11863,N_6981,N_8758);
and U11864 (N_11864,N_6264,N_8085);
nor U11865 (N_11865,N_9733,N_9620);
xor U11866 (N_11866,N_8384,N_9749);
nand U11867 (N_11867,N_6266,N_9817);
and U11868 (N_11868,N_7064,N_7537);
or U11869 (N_11869,N_7445,N_9734);
xor U11870 (N_11870,N_7684,N_6032);
nand U11871 (N_11871,N_9114,N_5377);
and U11872 (N_11872,N_5826,N_8179);
nand U11873 (N_11873,N_8075,N_7252);
nand U11874 (N_11874,N_8899,N_5837);
nand U11875 (N_11875,N_7467,N_5693);
xnor U11876 (N_11876,N_6280,N_8440);
nor U11877 (N_11877,N_7039,N_9776);
xnor U11878 (N_11878,N_9495,N_9904);
nor U11879 (N_11879,N_6198,N_5813);
nand U11880 (N_11880,N_9497,N_7913);
xnor U11881 (N_11881,N_5574,N_7704);
or U11882 (N_11882,N_7849,N_8644);
xnor U11883 (N_11883,N_5369,N_9844);
and U11884 (N_11884,N_6698,N_6334);
and U11885 (N_11885,N_7682,N_6896);
or U11886 (N_11886,N_9508,N_6895);
or U11887 (N_11887,N_7865,N_5632);
nand U11888 (N_11888,N_9756,N_8478);
nand U11889 (N_11889,N_9808,N_6917);
and U11890 (N_11890,N_8522,N_5203);
nor U11891 (N_11891,N_9803,N_6525);
and U11892 (N_11892,N_8932,N_5102);
or U11893 (N_11893,N_8996,N_5013);
nor U11894 (N_11894,N_9501,N_5016);
or U11895 (N_11895,N_7173,N_6772);
or U11896 (N_11896,N_8785,N_5070);
or U11897 (N_11897,N_8496,N_9856);
nor U11898 (N_11898,N_5744,N_7176);
nand U11899 (N_11899,N_5422,N_5394);
nand U11900 (N_11900,N_9787,N_7406);
or U11901 (N_11901,N_7166,N_7926);
or U11902 (N_11902,N_9034,N_6546);
or U11903 (N_11903,N_6484,N_6256);
or U11904 (N_11904,N_7495,N_6291);
nand U11905 (N_11905,N_7571,N_6251);
nand U11906 (N_11906,N_6838,N_6837);
or U11907 (N_11907,N_9929,N_9416);
or U11908 (N_11908,N_9091,N_6530);
nor U11909 (N_11909,N_6241,N_6126);
and U11910 (N_11910,N_5497,N_9868);
nor U11911 (N_11911,N_5999,N_5254);
nor U11912 (N_11912,N_5797,N_6005);
or U11913 (N_11913,N_5182,N_5694);
xor U11914 (N_11914,N_5212,N_5233);
nor U11915 (N_11915,N_5598,N_7307);
nand U11916 (N_11916,N_7506,N_6039);
nand U11917 (N_11917,N_9798,N_6649);
nand U11918 (N_11918,N_5552,N_6358);
nor U11919 (N_11919,N_9013,N_6082);
or U11920 (N_11920,N_9664,N_8125);
xnor U11921 (N_11921,N_6479,N_9156);
nor U11922 (N_11922,N_5720,N_6816);
or U11923 (N_11923,N_9723,N_9835);
or U11924 (N_11924,N_6614,N_5056);
nand U11925 (N_11925,N_6360,N_8364);
or U11926 (N_11926,N_6223,N_9315);
nand U11927 (N_11927,N_5935,N_8578);
nor U11928 (N_11928,N_5573,N_9376);
xor U11929 (N_11929,N_5907,N_7148);
nand U11930 (N_11930,N_8227,N_6375);
and U11931 (N_11931,N_7776,N_6716);
and U11932 (N_11932,N_9033,N_7084);
or U11933 (N_11933,N_6217,N_9311);
and U11934 (N_11934,N_7356,N_8813);
xnor U11935 (N_11935,N_5025,N_7310);
xor U11936 (N_11936,N_5348,N_6311);
or U11937 (N_11937,N_5528,N_9635);
or U11938 (N_11938,N_8947,N_6958);
nor U11939 (N_11939,N_7527,N_8214);
nand U11940 (N_11940,N_6788,N_9471);
xnor U11941 (N_11941,N_5833,N_6043);
xor U11942 (N_11942,N_9103,N_7689);
and U11943 (N_11943,N_8820,N_9901);
and U11944 (N_11944,N_8045,N_5177);
nor U11945 (N_11945,N_9675,N_6428);
or U11946 (N_11946,N_6750,N_5309);
nand U11947 (N_11947,N_9133,N_9726);
nand U11948 (N_11948,N_9041,N_9074);
or U11949 (N_11949,N_7958,N_8396);
nor U11950 (N_11950,N_5815,N_8811);
and U11951 (N_11951,N_9852,N_8048);
nor U11952 (N_11952,N_5872,N_8602);
xnor U11953 (N_11953,N_6939,N_9162);
nand U11954 (N_11954,N_5961,N_8123);
nand U11955 (N_11955,N_5969,N_7789);
or U11956 (N_11956,N_6074,N_5946);
and U11957 (N_11957,N_7523,N_6793);
and U11958 (N_11958,N_7178,N_7962);
xnor U11959 (N_11959,N_8569,N_5299);
and U11960 (N_11960,N_7350,N_8751);
or U11961 (N_11961,N_6615,N_5690);
and U11962 (N_11962,N_5894,N_7179);
nor U11963 (N_11963,N_6193,N_8143);
nand U11964 (N_11964,N_9946,N_5446);
or U11965 (N_11965,N_9457,N_9541);
and U11966 (N_11966,N_6984,N_9409);
xnor U11967 (N_11967,N_8945,N_9238);
xnor U11968 (N_11968,N_8052,N_8381);
or U11969 (N_11969,N_8023,N_6336);
nor U11970 (N_11970,N_5994,N_5572);
nor U11971 (N_11971,N_8418,N_6114);
nor U11972 (N_11972,N_5692,N_9958);
nand U11973 (N_11973,N_9015,N_8096);
xor U11974 (N_11974,N_6044,N_6921);
nor U11975 (N_11975,N_9563,N_7634);
nand U11976 (N_11976,N_8100,N_8244);
xor U11977 (N_11977,N_8545,N_9372);
xor U11978 (N_11978,N_8435,N_8669);
and U11979 (N_11979,N_8210,N_6758);
or U11980 (N_11980,N_9616,N_9104);
or U11981 (N_11981,N_5637,N_7744);
xor U11982 (N_11982,N_5482,N_7795);
or U11983 (N_11983,N_9320,N_8529);
and U11984 (N_11984,N_6504,N_6083);
and U11985 (N_11985,N_7869,N_6894);
nand U11986 (N_11986,N_9179,N_7076);
and U11987 (N_11987,N_5808,N_7233);
nor U11988 (N_11988,N_9139,N_6946);
xnor U11989 (N_11989,N_8072,N_8176);
nand U11990 (N_11990,N_6472,N_9851);
nand U11991 (N_11991,N_5576,N_6205);
and U11992 (N_11992,N_7258,N_7006);
nor U11993 (N_11993,N_6416,N_8905);
xor U11994 (N_11994,N_7522,N_9390);
xnor U11995 (N_11995,N_8810,N_5638);
and U11996 (N_11996,N_9714,N_6804);
or U11997 (N_11997,N_8784,N_8005);
nand U11998 (N_11998,N_7797,N_8389);
nor U11999 (N_11999,N_6577,N_9086);
nor U12000 (N_12000,N_7974,N_8709);
or U12001 (N_12001,N_7102,N_8093);
or U12002 (N_12002,N_9348,N_6639);
nand U12003 (N_12003,N_6873,N_8886);
xor U12004 (N_12004,N_6461,N_5703);
nor U12005 (N_12005,N_6427,N_5759);
xor U12006 (N_12006,N_5959,N_7031);
and U12007 (N_12007,N_9060,N_8175);
xor U12008 (N_12008,N_6911,N_7442);
nor U12009 (N_12009,N_8010,N_9236);
xnor U12010 (N_12010,N_5995,N_9650);
and U12011 (N_12011,N_7416,N_7680);
and U12012 (N_12012,N_8951,N_8663);
xnor U12013 (N_12013,N_5983,N_6438);
nor U12014 (N_12014,N_7934,N_8327);
xnor U12015 (N_12015,N_8893,N_5741);
and U12016 (N_12016,N_5642,N_5561);
or U12017 (N_12017,N_5487,N_5818);
or U12018 (N_12018,N_9645,N_6844);
nor U12019 (N_12019,N_8392,N_8429);
xnor U12020 (N_12020,N_8305,N_8469);
nand U12021 (N_12021,N_7736,N_5290);
or U12022 (N_12022,N_5037,N_6887);
or U12023 (N_12023,N_7821,N_9137);
nor U12024 (N_12024,N_5067,N_6379);
nor U12025 (N_12025,N_7025,N_5985);
and U12026 (N_12026,N_8313,N_7446);
xor U12027 (N_12027,N_8012,N_6355);
nor U12028 (N_12028,N_9643,N_5462);
and U12029 (N_12029,N_7685,N_7614);
xor U12030 (N_12030,N_6233,N_9774);
nand U12031 (N_12031,N_9145,N_8654);
or U12032 (N_12032,N_9496,N_6363);
nor U12033 (N_12033,N_6458,N_7781);
nor U12034 (N_12034,N_6144,N_7887);
nor U12035 (N_12035,N_7601,N_6783);
nor U12036 (N_12036,N_6403,N_6397);
nand U12037 (N_12037,N_7848,N_6296);
and U12038 (N_12038,N_8760,N_5654);
or U12039 (N_12039,N_9561,N_6132);
nor U12040 (N_12040,N_8019,N_5211);
xnor U12041 (N_12041,N_6582,N_9027);
or U12042 (N_12042,N_7264,N_8080);
nand U12043 (N_12043,N_6018,N_8105);
or U12044 (N_12044,N_6662,N_5749);
nand U12045 (N_12045,N_9010,N_7785);
and U12046 (N_12046,N_9811,N_8177);
nor U12047 (N_12047,N_9780,N_5876);
nand U12048 (N_12048,N_6965,N_5454);
and U12049 (N_12049,N_8225,N_5666);
nor U12050 (N_12050,N_9925,N_5857);
nand U12051 (N_12051,N_9062,N_9908);
xor U12052 (N_12052,N_9143,N_7617);
and U12053 (N_12053,N_5106,N_5058);
nand U12054 (N_12054,N_9474,N_8966);
and U12055 (N_12055,N_8326,N_5163);
nand U12056 (N_12056,N_7757,N_9692);
nand U12057 (N_12057,N_8728,N_7694);
nand U12058 (N_12058,N_7202,N_6488);
or U12059 (N_12059,N_6305,N_7419);
xnor U12060 (N_12060,N_6116,N_7902);
nand U12061 (N_12061,N_9319,N_6595);
xnor U12062 (N_12062,N_5278,N_7804);
xnor U12063 (N_12063,N_6608,N_8026);
and U12064 (N_12064,N_5865,N_8332);
nor U12065 (N_12065,N_8098,N_9061);
nand U12066 (N_12066,N_9470,N_9303);
nand U12067 (N_12067,N_8920,N_9290);
xnor U12068 (N_12068,N_7433,N_7329);
nor U12069 (N_12069,N_7950,N_7085);
and U12070 (N_12070,N_6410,N_9673);
or U12071 (N_12071,N_8616,N_6815);
nand U12072 (N_12072,N_5980,N_9368);
xnor U12073 (N_12073,N_8135,N_9163);
nor U12074 (N_12074,N_7248,N_6634);
or U12075 (N_12075,N_7521,N_6952);
xor U12076 (N_12076,N_8577,N_7798);
xnor U12077 (N_12077,N_8884,N_5340);
and U12078 (N_12078,N_9926,N_6668);
nor U12079 (N_12079,N_5989,N_8519);
and U12080 (N_12080,N_8705,N_8839);
and U12081 (N_12081,N_8054,N_8856);
nor U12082 (N_12082,N_7880,N_6439);
and U12083 (N_12083,N_9873,N_8649);
xnor U12084 (N_12084,N_8850,N_8178);
nor U12085 (N_12085,N_9816,N_8124);
and U12086 (N_12086,N_9101,N_9968);
xor U12087 (N_12087,N_6983,N_7528);
and U12088 (N_12088,N_5297,N_7128);
and U12089 (N_12089,N_8160,N_7481);
nor U12090 (N_12090,N_8289,N_7551);
nor U12091 (N_12091,N_6324,N_9391);
nand U12092 (N_12092,N_7585,N_9845);
nand U12093 (N_12093,N_8929,N_8340);
nor U12094 (N_12094,N_8735,N_7027);
or U12095 (N_12095,N_9003,N_8698);
xor U12096 (N_12096,N_5088,N_6013);
nand U12097 (N_12097,N_8659,N_5892);
and U12098 (N_12098,N_8083,N_6669);
nand U12099 (N_12099,N_5002,N_5256);
or U12100 (N_12100,N_9336,N_6888);
and U12101 (N_12101,N_5758,N_6632);
nor U12102 (N_12102,N_7589,N_8035);
or U12103 (N_12103,N_8053,N_7331);
nor U12104 (N_12104,N_6367,N_9120);
nor U12105 (N_12105,N_7017,N_8460);
nand U12106 (N_12106,N_5786,N_8088);
nor U12107 (N_12107,N_8937,N_9718);
nand U12108 (N_12108,N_5847,N_9028);
nand U12109 (N_12109,N_6857,N_5210);
nand U12110 (N_12110,N_5498,N_7285);
or U12111 (N_12111,N_9619,N_9891);
nor U12112 (N_12112,N_7130,N_6689);
or U12113 (N_12113,N_8128,N_6016);
and U12114 (N_12114,N_6096,N_5742);
xnor U12115 (N_12115,N_6288,N_9024);
nand U12116 (N_12116,N_7737,N_6395);
nor U12117 (N_12117,N_6890,N_7335);
xor U12118 (N_12118,N_7494,N_5138);
nand U12119 (N_12119,N_5065,N_6683);
nand U12120 (N_12120,N_5592,N_6693);
nor U12121 (N_12121,N_7126,N_6909);
and U12122 (N_12122,N_8352,N_8061);
or U12123 (N_12123,N_8523,N_6743);
nand U12124 (N_12124,N_5535,N_9669);
and U12125 (N_12125,N_7541,N_5746);
or U12126 (N_12126,N_8755,N_6746);
nand U12127 (N_12127,N_7024,N_7741);
or U12128 (N_12128,N_5611,N_8571);
and U12129 (N_12129,N_9895,N_6231);
xnor U12130 (N_12130,N_6765,N_6197);
and U12131 (N_12131,N_6100,N_9928);
or U12132 (N_12132,N_7324,N_9647);
and U12133 (N_12133,N_7702,N_5361);
xnor U12134 (N_12134,N_9267,N_7000);
and U12135 (N_12135,N_7842,N_5376);
nor U12136 (N_12136,N_8707,N_7322);
xnor U12137 (N_12137,N_6523,N_6507);
xor U12138 (N_12138,N_9437,N_5724);
xnor U12139 (N_12139,N_5325,N_8132);
nor U12140 (N_12140,N_9255,N_7141);
xnor U12141 (N_12141,N_8198,N_6680);
xnor U12142 (N_12142,N_9962,N_8889);
and U12143 (N_12143,N_7470,N_6440);
xor U12144 (N_12144,N_8060,N_9035);
nor U12145 (N_12145,N_9039,N_5433);
and U12146 (N_12146,N_8631,N_5172);
nand U12147 (N_12147,N_9299,N_8874);
and U12148 (N_12148,N_9979,N_9732);
or U12149 (N_12149,N_6621,N_5142);
xnor U12150 (N_12150,N_9406,N_5111);
or U12151 (N_12151,N_6436,N_5051);
xor U12152 (N_12152,N_6969,N_9468);
or U12153 (N_12153,N_7852,N_6160);
or U12154 (N_12154,N_5509,N_9919);
nand U12155 (N_12155,N_9948,N_5566);
xor U12156 (N_12156,N_8131,N_7937);
nor U12157 (N_12157,N_6861,N_6953);
nand U12158 (N_12158,N_5167,N_6524);
nand U12159 (N_12159,N_8957,N_9165);
nand U12160 (N_12160,N_6029,N_7152);
and U12161 (N_12161,N_7543,N_5671);
xor U12162 (N_12162,N_7275,N_6420);
or U12163 (N_12163,N_6734,N_7611);
or U12164 (N_12164,N_6019,N_6696);
xnor U12165 (N_12165,N_5008,N_6097);
nand U12166 (N_12166,N_5281,N_9393);
or U12167 (N_12167,N_9660,N_5118);
and U12168 (N_12168,N_6333,N_8344);
and U12169 (N_12169,N_9253,N_7383);
nand U12170 (N_12170,N_7688,N_6220);
xor U12171 (N_12171,N_6731,N_9981);
xor U12172 (N_12172,N_6924,N_7484);
and U12173 (N_12173,N_9587,N_8070);
nand U12174 (N_12174,N_8275,N_5202);
and U12175 (N_12175,N_7619,N_6852);
and U12176 (N_12176,N_6178,N_9106);
or U12177 (N_12177,N_6509,N_9863);
and U12178 (N_12178,N_8507,N_9896);
and U12179 (N_12179,N_7240,N_6918);
xor U12180 (N_12180,N_8681,N_7847);
xnor U12181 (N_12181,N_7564,N_9755);
nand U12182 (N_12182,N_5402,N_7473);
or U12183 (N_12183,N_5709,N_5856);
xor U12184 (N_12184,N_6900,N_5061);
nand U12185 (N_12185,N_8556,N_9131);
nand U12186 (N_12186,N_6129,N_5645);
nor U12187 (N_12187,N_5953,N_6588);
nor U12188 (N_12188,N_8449,N_6664);
xnor U12189 (N_12189,N_6940,N_9935);
xor U12190 (N_12190,N_6174,N_9943);
and U12191 (N_12191,N_9180,N_8434);
and U12192 (N_12192,N_6834,N_7691);
and U12193 (N_12193,N_8466,N_8356);
and U12194 (N_12194,N_5713,N_6344);
or U12195 (N_12195,N_7175,N_5464);
or U12196 (N_12196,N_8752,N_8882);
nor U12197 (N_12197,N_6801,N_5635);
and U12198 (N_12198,N_8422,N_5520);
and U12199 (N_12199,N_5506,N_6605);
and U12200 (N_12200,N_6192,N_9294);
and U12201 (N_12201,N_6671,N_6330);
or U12202 (N_12202,N_9414,N_6640);
and U12203 (N_12203,N_8407,N_5991);
or U12204 (N_12204,N_9209,N_7743);
nor U12205 (N_12205,N_6380,N_7318);
and U12206 (N_12206,N_8746,N_7115);
nand U12207 (N_12207,N_6842,N_6055);
xor U12208 (N_12208,N_6485,N_8057);
nand U12209 (N_12209,N_5440,N_6434);
nand U12210 (N_12210,N_5332,N_7813);
and U12211 (N_12211,N_6773,N_6681);
and U12212 (N_12212,N_9869,N_8975);
nand U12213 (N_12213,N_9046,N_7326);
and U12214 (N_12214,N_7596,N_5015);
nor U12215 (N_12215,N_6935,N_6699);
or U12216 (N_12216,N_6878,N_7866);
xnor U12217 (N_12217,N_8086,N_9584);
nor U12218 (N_12218,N_9261,N_9599);
and U12219 (N_12219,N_9394,N_6451);
xnor U12220 (N_12220,N_6000,N_5515);
nand U12221 (N_12221,N_7223,N_6359);
or U12222 (N_12222,N_7086,N_7044);
xnor U12223 (N_12223,N_9219,N_6237);
and U12224 (N_12224,N_5920,N_7392);
nor U12225 (N_12225,N_7370,N_9102);
nor U12226 (N_12226,N_8516,N_5132);
or U12227 (N_12227,N_7748,N_5197);
nor U12228 (N_12228,N_8572,N_8358);
or U12229 (N_12229,N_7975,N_5263);
or U12230 (N_12230,N_8232,N_5964);
xnor U12231 (N_12231,N_6101,N_5133);
xor U12232 (N_12232,N_7907,N_5539);
nand U12233 (N_12233,N_9292,N_8630);
nand U12234 (N_12234,N_9656,N_9305);
nand U12235 (N_12235,N_7536,N_7513);
nand U12236 (N_12236,N_5793,N_5519);
or U12237 (N_12237,N_9918,N_6189);
nand U12238 (N_12238,N_5360,N_7206);
nor U12239 (N_12239,N_7878,N_5124);
xnor U12240 (N_12240,N_9524,N_9176);
nand U12241 (N_12241,N_5979,N_5544);
or U12242 (N_12242,N_6744,N_8798);
xnor U12243 (N_12243,N_8629,N_5411);
nor U12244 (N_12244,N_5831,N_7447);
or U12245 (N_12245,N_7303,N_8284);
and U12246 (N_12246,N_6956,N_8938);
xor U12247 (N_12247,N_9171,N_9375);
xnor U12248 (N_12248,N_5716,N_5005);
nor U12249 (N_12249,N_7367,N_6444);
nor U12250 (N_12250,N_5221,N_7725);
xnor U12251 (N_12251,N_6050,N_8559);
xor U12252 (N_12252,N_6784,N_7068);
xnor U12253 (N_12253,N_8678,N_8300);
nor U12254 (N_12254,N_9892,N_7641);
nor U12255 (N_12255,N_6575,N_9636);
or U12256 (N_12256,N_9445,N_9717);
and U12257 (N_12257,N_7633,N_8370);
or U12258 (N_12258,N_6982,N_6893);
nand U12259 (N_12259,N_8880,N_8445);
xnor U12260 (N_12260,N_9444,N_5194);
nand U12261 (N_12261,N_6865,N_6707);
and U12262 (N_12262,N_8949,N_5119);
and U12263 (N_12263,N_9521,N_5179);
and U12264 (N_12264,N_5547,N_6752);
nor U12265 (N_12265,N_5001,N_5198);
nor U12266 (N_12266,N_7731,N_9193);
nand U12267 (N_12267,N_9907,N_8208);
nand U12268 (N_12268,N_8247,N_6385);
xor U12269 (N_12269,N_7201,N_5159);
and U12270 (N_12270,N_6902,N_9075);
and U12271 (N_12271,N_6413,N_8027);
nand U12272 (N_12272,N_8730,N_5170);
nand U12273 (N_12273,N_6721,N_6558);
or U12274 (N_12274,N_5531,N_6796);
nor U12275 (N_12275,N_6338,N_7995);
or U12276 (N_12276,N_8800,N_9655);
xor U12277 (N_12277,N_5214,N_5087);
nand U12278 (N_12278,N_9727,N_9885);
nor U12279 (N_12279,N_9898,N_6938);
and U12280 (N_12280,N_9543,N_8484);
nor U12281 (N_12281,N_7135,N_9006);
or U12282 (N_12282,N_6813,N_9857);
and U12283 (N_12283,N_5864,N_6478);
nand U12284 (N_12284,N_5414,N_5548);
or U12285 (N_12285,N_9826,N_6270);
or U12286 (N_12286,N_8278,N_5338);
nor U12287 (N_12287,N_9649,N_8797);
nor U12288 (N_12288,N_6432,N_6856);
nor U12289 (N_12289,N_6991,N_7155);
and U12290 (N_12290,N_5012,N_8317);
xnor U12291 (N_12291,N_9067,N_5702);
and U12292 (N_12292,N_8699,N_5976);
xnor U12293 (N_12293,N_5285,N_6998);
xor U12294 (N_12294,N_6190,N_7539);
xnor U12295 (N_12295,N_9096,N_7079);
nand U12296 (N_12296,N_9793,N_6794);
and U12297 (N_12297,N_9698,N_7407);
nand U12298 (N_12298,N_5830,N_5484);
nand U12299 (N_12299,N_5795,N_9274);
xor U12300 (N_12300,N_6041,N_9992);
nand U12301 (N_12301,N_9767,N_9560);
or U12302 (N_12302,N_7881,N_6459);
nor U12303 (N_12303,N_9441,N_8439);
nor U12304 (N_12304,N_5443,N_8922);
nand U12305 (N_12305,N_9456,N_9574);
or U12306 (N_12306,N_5292,N_7140);
nor U12307 (N_12307,N_6084,N_5799);
xor U12308 (N_12308,N_8869,N_7766);
nor U12309 (N_12309,N_7032,N_8116);
or U12310 (N_12310,N_9207,N_9994);
nand U12311 (N_12311,N_6156,N_7758);
and U12312 (N_12312,N_6398,N_9455);
and U12313 (N_12313,N_9463,N_9295);
and U12314 (N_12314,N_8452,N_8687);
xor U12315 (N_12315,N_9847,N_7638);
nand U12316 (N_12316,N_6245,N_6462);
or U12317 (N_12317,N_9023,N_5321);
xnor U12318 (N_12318,N_9302,N_7973);
and U12319 (N_12319,N_8623,N_5701);
xor U12320 (N_12320,N_8068,N_8697);
nor U12321 (N_12321,N_8008,N_6317);
nand U12322 (N_12322,N_6610,N_5150);
nand U12323 (N_12323,N_7639,N_9602);
xor U12324 (N_12324,N_8087,N_7107);
xnor U12325 (N_12325,N_9177,N_9579);
nor U12326 (N_12326,N_5077,N_6996);
nand U12327 (N_12327,N_8153,N_7194);
xor U12328 (N_12328,N_5500,N_8521);
or U12329 (N_12329,N_7976,N_9168);
and U12330 (N_12330,N_6512,N_6651);
xnor U12331 (N_12331,N_8417,N_7624);
or U12332 (N_12332,N_5586,N_8268);
xnor U12333 (N_12333,N_8688,N_5145);
xnor U12334 (N_12334,N_9850,N_7761);
nand U12335 (N_12335,N_5945,N_6881);
xnor U12336 (N_12336,N_9596,N_5358);
and U12337 (N_12337,N_8316,N_9991);
or U12338 (N_12338,N_9554,N_9558);
nor U12339 (N_12339,N_7945,N_6563);
nand U12340 (N_12340,N_8955,N_7923);
nand U12341 (N_12341,N_7236,N_5184);
nand U12342 (N_12342,N_6072,N_8719);
xor U12343 (N_12343,N_7172,N_8939);
xor U12344 (N_12344,N_7040,N_5748);
and U12345 (N_12345,N_7474,N_7073);
xnor U12346 (N_12346,N_5050,N_6916);
and U12347 (N_12347,N_6390,N_9824);
xnor U12348 (N_12348,N_7376,N_8774);
nand U12349 (N_12349,N_5608,N_7434);
and U12350 (N_12350,N_5085,N_6855);
nand U12351 (N_12351,N_6183,N_9194);
nor U12352 (N_12352,N_6031,N_7879);
nor U12353 (N_12353,N_8448,N_8127);
xnor U12354 (N_12354,N_8537,N_6170);
nand U12355 (N_12355,N_8041,N_7643);
nand U12356 (N_12356,N_6867,N_8183);
xnor U12357 (N_12357,N_7768,N_6695);
nor U12358 (N_12358,N_7218,N_6726);
nand U12359 (N_12359,N_7366,N_9839);
or U12360 (N_12360,N_7070,N_6737);
nor U12361 (N_12361,N_5810,N_7355);
nor U12362 (N_12362,N_7023,N_6764);
nand U12363 (N_12363,N_5512,N_7561);
and U12364 (N_12364,N_6200,N_6068);
nor U12365 (N_12365,N_5717,N_7558);
and U12366 (N_12366,N_6905,N_7424);
xnor U12367 (N_12367,N_7412,N_7886);
xnor U12368 (N_12368,N_6557,N_9152);
xnor U12369 (N_12369,N_5274,N_6593);
nor U12370 (N_12370,N_7594,N_9388);
or U12371 (N_12371,N_9989,N_7616);
and U12372 (N_12372,N_8581,N_6692);
nor U12373 (N_12373,N_5829,N_7953);
xnor U12374 (N_12374,N_6506,N_7646);
nand U12375 (N_12375,N_5035,N_9679);
xor U12376 (N_12376,N_5417,N_6959);
or U12377 (N_12377,N_7919,N_5190);
nand U12378 (N_12378,N_5875,N_6155);
xor U12379 (N_12379,N_7411,N_5681);
or U12380 (N_12380,N_7250,N_8174);
xor U12381 (N_12381,N_8353,N_7542);
xor U12382 (N_12382,N_7514,N_9208);
xor U12383 (N_12383,N_7825,N_7890);
nor U12384 (N_12384,N_8473,N_8887);
nand U12385 (N_12385,N_5386,N_6974);
and U12386 (N_12386,N_5879,N_8601);
or U12387 (N_12387,N_6703,N_6875);
nor U12388 (N_12388,N_6648,N_6795);
and U12389 (N_12389,N_7894,N_5545);
xnor U12390 (N_12390,N_9570,N_6532);
or U12391 (N_12391,N_5130,N_6985);
or U12392 (N_12392,N_5740,N_6229);
nand U12393 (N_12393,N_8793,N_6033);
nand U12394 (N_12394,N_7090,N_7475);
or U12395 (N_12395,N_6520,N_6971);
nand U12396 (N_12396,N_9071,N_5706);
and U12397 (N_12397,N_8442,N_5600);
or U12398 (N_12398,N_6165,N_5200);
and U12399 (N_12399,N_6235,N_6310);
and U12400 (N_12400,N_5569,N_6445);
nor U12401 (N_12401,N_6931,N_9031);
xor U12402 (N_12402,N_8357,N_9548);
xor U12403 (N_12403,N_9668,N_9980);
nand U12404 (N_12404,N_9985,N_6191);
nand U12405 (N_12405,N_8149,N_7113);
or U12406 (N_12406,N_6552,N_5963);
nor U12407 (N_12407,N_8264,N_8386);
nor U12408 (N_12408,N_6090,N_8454);
nor U12409 (N_12409,N_8495,N_5442);
and U12410 (N_12410,N_6455,N_6667);
xnor U12411 (N_12411,N_9486,N_6600);
and U12412 (N_12412,N_6776,N_8691);
nor U12413 (N_12413,N_8909,N_8369);
nor U12414 (N_12414,N_9678,N_7840);
and U12415 (N_12415,N_8761,N_6463);
xnor U12416 (N_12416,N_8180,N_5033);
nand U12417 (N_12417,N_5347,N_7301);
or U12418 (N_12418,N_9831,N_9610);
nand U12419 (N_12419,N_7577,N_9279);
nor U12420 (N_12420,N_8918,N_6468);
xor U12421 (N_12421,N_7948,N_5893);
and U12422 (N_12422,N_8151,N_7151);
xor U12423 (N_12423,N_9385,N_9173);
and U12424 (N_12424,N_7298,N_9757);
or U12425 (N_12425,N_5802,N_6009);
xnor U12426 (N_12426,N_6409,N_9990);
nand U12427 (N_12427,N_7459,N_6138);
xor U12428 (N_12428,N_9510,N_7674);
nand U12429 (N_12429,N_8489,N_5970);
and U12430 (N_12430,N_8720,N_7365);
xor U12431 (N_12431,N_6987,N_7606);
or U12432 (N_12432,N_5636,N_5122);
nor U12433 (N_12433,N_8191,N_7147);
xnor U12434 (N_12434,N_6254,N_9940);
xnor U12435 (N_12435,N_9355,N_6399);
nand U12436 (N_12436,N_8565,N_8610);
or U12437 (N_12437,N_9237,N_8643);
and U12438 (N_12438,N_6077,N_6606);
nor U12439 (N_12439,N_8729,N_7546);
xnor U12440 (N_12440,N_7004,N_9263);
and U12441 (N_12441,N_8413,N_7984);
nor U12442 (N_12442,N_9243,N_5619);
nor U12443 (N_12443,N_9283,N_7114);
xor U12444 (N_12444,N_9364,N_7531);
nand U12445 (N_12445,N_8419,N_6025);
or U12446 (N_12446,N_9995,N_7262);
xnor U12447 (N_12447,N_8535,N_7918);
nor U12448 (N_12448,N_6313,N_5222);
xor U12449 (N_12449,N_9373,N_7623);
and U12450 (N_12450,N_8427,N_6373);
or U12451 (N_12451,N_9730,N_9188);
or U12452 (N_12452,N_7154,N_8805);
nor U12453 (N_12453,N_8656,N_9121);
or U12454 (N_12454,N_9094,N_6383);
and U12455 (N_12455,N_8297,N_8458);
xor U12456 (N_12456,N_5518,N_7208);
or U12457 (N_12457,N_7946,N_8226);
and U12458 (N_12458,N_8166,N_9159);
nand U12459 (N_12459,N_9481,N_9360);
or U12460 (N_12460,N_8021,N_5962);
and U12461 (N_12461,N_6209,N_8109);
and U12462 (N_12462,N_5224,N_8548);
or U12463 (N_12463,N_6052,N_9938);
and U12464 (N_12464,N_9688,N_6301);
xor U12465 (N_12465,N_6858,N_5154);
or U12466 (N_12466,N_6686,N_6087);
nor U12467 (N_12467,N_7496,N_8380);
nand U12468 (N_12468,N_6376,N_6650);
nand U12469 (N_12469,N_5650,N_6840);
nor U12470 (N_12470,N_6950,N_9870);
xor U12471 (N_12471,N_9397,N_5739);
nand U12472 (N_12472,N_7415,N_8862);
xnor U12473 (N_12473,N_5426,N_6456);
xnor U12474 (N_12474,N_5887,N_7466);
xnor U12475 (N_12475,N_9226,N_7752);
and U12476 (N_12476,N_9736,N_7563);
and U12477 (N_12477,N_5807,N_9358);
and U12478 (N_12478,N_5335,N_6989);
xor U12479 (N_12479,N_7413,N_6607);
and U12480 (N_12480,N_5789,N_8794);
nand U12481 (N_12481,N_8652,N_5564);
xor U12482 (N_12482,N_6215,N_8657);
nand U12483 (N_12483,N_5643,N_5505);
or U12484 (N_12484,N_9382,N_5551);
or U12485 (N_12485,N_8347,N_8536);
or U12486 (N_12486,N_6098,N_9473);
or U12487 (N_12487,N_8490,N_8710);
nor U12488 (N_12488,N_6213,N_6139);
nand U12489 (N_12489,N_9117,N_6346);
nor U12490 (N_12490,N_8608,N_8622);
and U12491 (N_12491,N_5380,N_7465);
nor U12492 (N_12492,N_7499,N_8564);
and U12493 (N_12493,N_9272,N_7182);
xor U12494 (N_12494,N_7569,N_5135);
xor U12495 (N_12495,N_7963,N_9509);
nor U12496 (N_12496,N_9065,N_9905);
xnor U12497 (N_12497,N_8170,N_7709);
and U12498 (N_12498,N_5655,N_7636);
nor U12499 (N_12499,N_6262,N_8401);
nand U12500 (N_12500,N_5317,N_6125);
or U12501 (N_12501,N_5923,N_6788);
or U12502 (N_12502,N_8818,N_5291);
xor U12503 (N_12503,N_7983,N_7709);
nand U12504 (N_12504,N_8002,N_7236);
and U12505 (N_12505,N_8309,N_7518);
and U12506 (N_12506,N_7889,N_9314);
and U12507 (N_12507,N_7285,N_7904);
and U12508 (N_12508,N_6061,N_8113);
nand U12509 (N_12509,N_5401,N_9676);
and U12510 (N_12510,N_7492,N_7563);
and U12511 (N_12511,N_9068,N_6558);
and U12512 (N_12512,N_6513,N_7733);
nand U12513 (N_12513,N_8854,N_5387);
nor U12514 (N_12514,N_5697,N_5485);
xor U12515 (N_12515,N_9966,N_8199);
nand U12516 (N_12516,N_9557,N_8309);
or U12517 (N_12517,N_8342,N_5864);
nand U12518 (N_12518,N_9103,N_9289);
or U12519 (N_12519,N_9293,N_9577);
nor U12520 (N_12520,N_5612,N_8111);
xnor U12521 (N_12521,N_9245,N_7018);
nand U12522 (N_12522,N_6401,N_6521);
xnor U12523 (N_12523,N_6119,N_9993);
nand U12524 (N_12524,N_8616,N_5045);
and U12525 (N_12525,N_5985,N_6410);
or U12526 (N_12526,N_5862,N_5062);
xor U12527 (N_12527,N_9305,N_5527);
or U12528 (N_12528,N_5639,N_8055);
xnor U12529 (N_12529,N_8954,N_6642);
or U12530 (N_12530,N_7304,N_5363);
xor U12531 (N_12531,N_7872,N_8230);
or U12532 (N_12532,N_6316,N_8225);
nand U12533 (N_12533,N_5656,N_7394);
and U12534 (N_12534,N_8827,N_9744);
nand U12535 (N_12535,N_6351,N_5345);
nor U12536 (N_12536,N_6956,N_6671);
xnor U12537 (N_12537,N_9121,N_5317);
and U12538 (N_12538,N_9121,N_5617);
and U12539 (N_12539,N_6228,N_5425);
or U12540 (N_12540,N_6529,N_5647);
nor U12541 (N_12541,N_5990,N_5810);
and U12542 (N_12542,N_7780,N_9669);
and U12543 (N_12543,N_7609,N_5471);
and U12544 (N_12544,N_9115,N_6804);
or U12545 (N_12545,N_5163,N_5404);
and U12546 (N_12546,N_7796,N_5176);
nand U12547 (N_12547,N_6316,N_5707);
or U12548 (N_12548,N_6089,N_9734);
nor U12549 (N_12549,N_8745,N_6048);
nand U12550 (N_12550,N_7771,N_6673);
nand U12551 (N_12551,N_5442,N_6749);
and U12552 (N_12552,N_7614,N_7861);
and U12553 (N_12553,N_7172,N_9999);
and U12554 (N_12554,N_9270,N_8672);
nor U12555 (N_12555,N_5644,N_5093);
xnor U12556 (N_12556,N_9883,N_7997);
xor U12557 (N_12557,N_8820,N_6344);
and U12558 (N_12558,N_9380,N_6736);
nor U12559 (N_12559,N_8615,N_8278);
nand U12560 (N_12560,N_6610,N_6260);
and U12561 (N_12561,N_6310,N_9127);
nor U12562 (N_12562,N_6799,N_8023);
nand U12563 (N_12563,N_5971,N_6502);
xor U12564 (N_12564,N_6696,N_6790);
nand U12565 (N_12565,N_8334,N_7839);
or U12566 (N_12566,N_9408,N_6402);
or U12567 (N_12567,N_8136,N_9522);
and U12568 (N_12568,N_7364,N_9123);
nand U12569 (N_12569,N_9507,N_5856);
nor U12570 (N_12570,N_7464,N_7739);
nand U12571 (N_12571,N_9507,N_5212);
nor U12572 (N_12572,N_5329,N_9172);
xnor U12573 (N_12573,N_9333,N_6577);
nand U12574 (N_12574,N_8197,N_7030);
nor U12575 (N_12575,N_7910,N_9980);
nor U12576 (N_12576,N_5924,N_8823);
and U12577 (N_12577,N_8350,N_5178);
xor U12578 (N_12578,N_9747,N_9943);
nand U12579 (N_12579,N_9170,N_6948);
and U12580 (N_12580,N_6778,N_9193);
and U12581 (N_12581,N_6487,N_9776);
nand U12582 (N_12582,N_6998,N_7614);
nand U12583 (N_12583,N_7849,N_5888);
nand U12584 (N_12584,N_9303,N_8070);
nor U12585 (N_12585,N_6022,N_7537);
and U12586 (N_12586,N_5697,N_9694);
nor U12587 (N_12587,N_6329,N_5298);
nand U12588 (N_12588,N_7738,N_6774);
and U12589 (N_12589,N_6119,N_5129);
or U12590 (N_12590,N_9845,N_8383);
xnor U12591 (N_12591,N_5301,N_6635);
nor U12592 (N_12592,N_6248,N_5301);
and U12593 (N_12593,N_6739,N_8908);
nor U12594 (N_12594,N_6834,N_7833);
nand U12595 (N_12595,N_7251,N_9533);
xnor U12596 (N_12596,N_7299,N_6155);
nor U12597 (N_12597,N_8337,N_9706);
and U12598 (N_12598,N_7131,N_8851);
and U12599 (N_12599,N_5082,N_9104);
xnor U12600 (N_12600,N_7422,N_7068);
xor U12601 (N_12601,N_6823,N_8179);
and U12602 (N_12602,N_5682,N_5480);
nand U12603 (N_12603,N_6871,N_9248);
or U12604 (N_12604,N_6876,N_5063);
nor U12605 (N_12605,N_5144,N_5710);
and U12606 (N_12606,N_5757,N_9045);
and U12607 (N_12607,N_9137,N_7466);
or U12608 (N_12608,N_7649,N_6420);
or U12609 (N_12609,N_5865,N_8157);
xor U12610 (N_12610,N_7859,N_8120);
xor U12611 (N_12611,N_8781,N_9856);
or U12612 (N_12612,N_6475,N_5866);
xor U12613 (N_12613,N_8143,N_9274);
nor U12614 (N_12614,N_6733,N_9098);
nand U12615 (N_12615,N_8410,N_7626);
and U12616 (N_12616,N_5906,N_9005);
and U12617 (N_12617,N_8256,N_5438);
and U12618 (N_12618,N_9589,N_9627);
nand U12619 (N_12619,N_7126,N_9646);
nor U12620 (N_12620,N_8616,N_6261);
or U12621 (N_12621,N_8093,N_7299);
nor U12622 (N_12622,N_9392,N_6279);
nor U12623 (N_12623,N_9159,N_9516);
nor U12624 (N_12624,N_6581,N_5945);
xor U12625 (N_12625,N_8588,N_6987);
or U12626 (N_12626,N_5975,N_9493);
or U12627 (N_12627,N_6113,N_6551);
and U12628 (N_12628,N_7826,N_7840);
nor U12629 (N_12629,N_9650,N_8954);
or U12630 (N_12630,N_5400,N_5592);
or U12631 (N_12631,N_6067,N_5071);
xor U12632 (N_12632,N_7201,N_9121);
nand U12633 (N_12633,N_6262,N_9679);
nor U12634 (N_12634,N_8229,N_5509);
nand U12635 (N_12635,N_7812,N_6297);
xnor U12636 (N_12636,N_8842,N_7117);
nand U12637 (N_12637,N_6886,N_8908);
or U12638 (N_12638,N_5559,N_5211);
xor U12639 (N_12639,N_5872,N_7376);
and U12640 (N_12640,N_9806,N_8637);
nor U12641 (N_12641,N_9152,N_7639);
or U12642 (N_12642,N_6486,N_5244);
and U12643 (N_12643,N_9703,N_6693);
xnor U12644 (N_12644,N_6866,N_5282);
xor U12645 (N_12645,N_6089,N_8185);
xnor U12646 (N_12646,N_8032,N_7941);
or U12647 (N_12647,N_7481,N_9566);
nand U12648 (N_12648,N_6929,N_6141);
nor U12649 (N_12649,N_8453,N_6337);
nand U12650 (N_12650,N_9257,N_9271);
or U12651 (N_12651,N_9880,N_8206);
or U12652 (N_12652,N_8296,N_5237);
xor U12653 (N_12653,N_7554,N_6509);
and U12654 (N_12654,N_8387,N_9253);
xnor U12655 (N_12655,N_7081,N_9332);
or U12656 (N_12656,N_8568,N_6874);
xnor U12657 (N_12657,N_5273,N_7305);
or U12658 (N_12658,N_5564,N_5783);
or U12659 (N_12659,N_5623,N_6782);
xor U12660 (N_12660,N_6569,N_5274);
xnor U12661 (N_12661,N_5445,N_8762);
or U12662 (N_12662,N_6497,N_6948);
nand U12663 (N_12663,N_6822,N_6355);
nor U12664 (N_12664,N_8509,N_5903);
or U12665 (N_12665,N_7633,N_5627);
xnor U12666 (N_12666,N_8694,N_8997);
and U12667 (N_12667,N_9313,N_7706);
nor U12668 (N_12668,N_8269,N_7144);
nand U12669 (N_12669,N_9059,N_9981);
or U12670 (N_12670,N_9244,N_6611);
and U12671 (N_12671,N_9664,N_9799);
and U12672 (N_12672,N_5404,N_9241);
and U12673 (N_12673,N_9138,N_6130);
and U12674 (N_12674,N_9559,N_6574);
and U12675 (N_12675,N_6937,N_8704);
or U12676 (N_12676,N_5390,N_6546);
nand U12677 (N_12677,N_5791,N_5446);
nand U12678 (N_12678,N_9246,N_8503);
nand U12679 (N_12679,N_8929,N_5044);
and U12680 (N_12680,N_5889,N_7866);
nor U12681 (N_12681,N_9175,N_7242);
xor U12682 (N_12682,N_9742,N_7295);
xor U12683 (N_12683,N_8703,N_8658);
nor U12684 (N_12684,N_7152,N_5255);
and U12685 (N_12685,N_6995,N_5485);
nor U12686 (N_12686,N_5763,N_5184);
or U12687 (N_12687,N_5566,N_7373);
xnor U12688 (N_12688,N_6801,N_7538);
nand U12689 (N_12689,N_6890,N_6994);
and U12690 (N_12690,N_9570,N_9591);
and U12691 (N_12691,N_7006,N_7020);
nand U12692 (N_12692,N_9512,N_7339);
or U12693 (N_12693,N_6488,N_7290);
or U12694 (N_12694,N_7155,N_5196);
xor U12695 (N_12695,N_7946,N_8653);
and U12696 (N_12696,N_5151,N_9107);
nor U12697 (N_12697,N_7892,N_6058);
or U12698 (N_12698,N_9465,N_7016);
xnor U12699 (N_12699,N_8372,N_9471);
nand U12700 (N_12700,N_6803,N_5569);
nor U12701 (N_12701,N_9328,N_5707);
and U12702 (N_12702,N_8480,N_5742);
xor U12703 (N_12703,N_8598,N_6802);
nand U12704 (N_12704,N_6842,N_6988);
xor U12705 (N_12705,N_8160,N_8202);
nor U12706 (N_12706,N_8617,N_8543);
nand U12707 (N_12707,N_9392,N_6290);
nor U12708 (N_12708,N_9549,N_8502);
xor U12709 (N_12709,N_8606,N_6149);
nand U12710 (N_12710,N_6106,N_9590);
and U12711 (N_12711,N_6138,N_8188);
or U12712 (N_12712,N_9370,N_7387);
xor U12713 (N_12713,N_8552,N_7417);
nor U12714 (N_12714,N_5032,N_6714);
or U12715 (N_12715,N_7150,N_8289);
nor U12716 (N_12716,N_8086,N_9976);
and U12717 (N_12717,N_9070,N_5214);
and U12718 (N_12718,N_6190,N_6524);
xor U12719 (N_12719,N_9492,N_8622);
and U12720 (N_12720,N_5033,N_7062);
xor U12721 (N_12721,N_6264,N_9014);
or U12722 (N_12722,N_8228,N_6480);
xnor U12723 (N_12723,N_6324,N_8522);
xnor U12724 (N_12724,N_5187,N_6293);
xnor U12725 (N_12725,N_5818,N_8922);
nor U12726 (N_12726,N_9734,N_7576);
or U12727 (N_12727,N_7877,N_6265);
or U12728 (N_12728,N_8929,N_8607);
xor U12729 (N_12729,N_6786,N_9871);
nor U12730 (N_12730,N_6623,N_5097);
nor U12731 (N_12731,N_8269,N_7000);
or U12732 (N_12732,N_5242,N_6196);
nor U12733 (N_12733,N_7115,N_8667);
and U12734 (N_12734,N_5168,N_9214);
and U12735 (N_12735,N_6148,N_6530);
or U12736 (N_12736,N_7080,N_6080);
nor U12737 (N_12737,N_8357,N_8617);
nor U12738 (N_12738,N_6044,N_9580);
nand U12739 (N_12739,N_5301,N_6265);
nand U12740 (N_12740,N_5843,N_5353);
or U12741 (N_12741,N_5872,N_8346);
or U12742 (N_12742,N_7116,N_8078);
or U12743 (N_12743,N_6403,N_9579);
nor U12744 (N_12744,N_9302,N_5824);
or U12745 (N_12745,N_7705,N_9422);
or U12746 (N_12746,N_7309,N_5634);
or U12747 (N_12747,N_5071,N_7440);
nand U12748 (N_12748,N_5785,N_8318);
nand U12749 (N_12749,N_9218,N_5734);
xnor U12750 (N_12750,N_6309,N_8556);
and U12751 (N_12751,N_9509,N_8273);
nor U12752 (N_12752,N_9460,N_6831);
xnor U12753 (N_12753,N_9387,N_6708);
nand U12754 (N_12754,N_9951,N_9319);
and U12755 (N_12755,N_6570,N_6218);
nand U12756 (N_12756,N_9322,N_7172);
xnor U12757 (N_12757,N_9975,N_8245);
and U12758 (N_12758,N_9180,N_7708);
or U12759 (N_12759,N_9574,N_7390);
nand U12760 (N_12760,N_5021,N_9508);
nand U12761 (N_12761,N_9153,N_8210);
or U12762 (N_12762,N_8228,N_7565);
and U12763 (N_12763,N_7499,N_5945);
nand U12764 (N_12764,N_8799,N_5821);
or U12765 (N_12765,N_8454,N_8161);
xnor U12766 (N_12766,N_6476,N_8327);
nand U12767 (N_12767,N_6161,N_5716);
nor U12768 (N_12768,N_8799,N_8798);
nor U12769 (N_12769,N_6873,N_8520);
nand U12770 (N_12770,N_5826,N_7891);
and U12771 (N_12771,N_7480,N_8745);
xnor U12772 (N_12772,N_8030,N_9591);
xor U12773 (N_12773,N_6799,N_8908);
or U12774 (N_12774,N_8311,N_7144);
or U12775 (N_12775,N_8015,N_8617);
or U12776 (N_12776,N_5174,N_9359);
or U12777 (N_12777,N_8170,N_5822);
and U12778 (N_12778,N_9909,N_5534);
nand U12779 (N_12779,N_7591,N_8308);
and U12780 (N_12780,N_8831,N_5556);
nor U12781 (N_12781,N_5436,N_8798);
nand U12782 (N_12782,N_9549,N_5609);
or U12783 (N_12783,N_8185,N_7049);
nor U12784 (N_12784,N_7370,N_5828);
and U12785 (N_12785,N_6403,N_9722);
nand U12786 (N_12786,N_9199,N_7339);
nor U12787 (N_12787,N_7920,N_9426);
nand U12788 (N_12788,N_6590,N_8442);
and U12789 (N_12789,N_5143,N_5469);
xnor U12790 (N_12790,N_5648,N_7004);
nand U12791 (N_12791,N_7499,N_8953);
xnor U12792 (N_12792,N_7707,N_9058);
xor U12793 (N_12793,N_6763,N_9807);
xnor U12794 (N_12794,N_5097,N_8933);
nand U12795 (N_12795,N_9737,N_5529);
nor U12796 (N_12796,N_8709,N_6422);
nand U12797 (N_12797,N_9260,N_9997);
and U12798 (N_12798,N_8204,N_6202);
nor U12799 (N_12799,N_6812,N_5761);
xnor U12800 (N_12800,N_9506,N_9149);
nand U12801 (N_12801,N_6820,N_6565);
or U12802 (N_12802,N_7486,N_6848);
nor U12803 (N_12803,N_8825,N_9951);
nor U12804 (N_12804,N_6069,N_6738);
xor U12805 (N_12805,N_8595,N_7132);
nor U12806 (N_12806,N_8383,N_7354);
and U12807 (N_12807,N_5228,N_6953);
nor U12808 (N_12808,N_7784,N_9512);
xor U12809 (N_12809,N_9115,N_5595);
or U12810 (N_12810,N_8369,N_8109);
nor U12811 (N_12811,N_9802,N_7921);
xnor U12812 (N_12812,N_7753,N_7813);
nand U12813 (N_12813,N_8240,N_9335);
nand U12814 (N_12814,N_6446,N_8419);
xor U12815 (N_12815,N_7841,N_8994);
and U12816 (N_12816,N_5842,N_8869);
and U12817 (N_12817,N_7399,N_7610);
nor U12818 (N_12818,N_9532,N_9884);
and U12819 (N_12819,N_8161,N_9952);
xor U12820 (N_12820,N_8055,N_8811);
nor U12821 (N_12821,N_8988,N_9606);
or U12822 (N_12822,N_8924,N_8028);
or U12823 (N_12823,N_5057,N_6199);
nor U12824 (N_12824,N_9777,N_7282);
or U12825 (N_12825,N_9990,N_7430);
nand U12826 (N_12826,N_7890,N_7612);
and U12827 (N_12827,N_5273,N_6496);
or U12828 (N_12828,N_5131,N_7398);
nor U12829 (N_12829,N_5152,N_8840);
nand U12830 (N_12830,N_7596,N_6483);
nand U12831 (N_12831,N_9772,N_9547);
and U12832 (N_12832,N_8660,N_5907);
and U12833 (N_12833,N_8076,N_5478);
xor U12834 (N_12834,N_8388,N_9987);
nand U12835 (N_12835,N_6907,N_9135);
or U12836 (N_12836,N_8562,N_7983);
and U12837 (N_12837,N_5169,N_9016);
and U12838 (N_12838,N_8859,N_9302);
or U12839 (N_12839,N_5707,N_8602);
xor U12840 (N_12840,N_5696,N_6369);
and U12841 (N_12841,N_5807,N_8987);
xor U12842 (N_12842,N_9647,N_8629);
nand U12843 (N_12843,N_6575,N_8179);
xor U12844 (N_12844,N_8090,N_7596);
nand U12845 (N_12845,N_5099,N_5732);
and U12846 (N_12846,N_6945,N_5166);
nand U12847 (N_12847,N_6672,N_7829);
xnor U12848 (N_12848,N_9109,N_8855);
nand U12849 (N_12849,N_6905,N_6352);
nand U12850 (N_12850,N_6110,N_7755);
xor U12851 (N_12851,N_8300,N_5588);
nand U12852 (N_12852,N_7254,N_8599);
nor U12853 (N_12853,N_5659,N_9007);
nor U12854 (N_12854,N_9666,N_7131);
and U12855 (N_12855,N_7484,N_8915);
nor U12856 (N_12856,N_7026,N_7759);
xnor U12857 (N_12857,N_7416,N_6971);
nor U12858 (N_12858,N_9107,N_7749);
nor U12859 (N_12859,N_8790,N_6828);
xnor U12860 (N_12860,N_7821,N_5719);
and U12861 (N_12861,N_6441,N_5475);
and U12862 (N_12862,N_5340,N_9176);
nand U12863 (N_12863,N_7449,N_9845);
and U12864 (N_12864,N_8123,N_9494);
and U12865 (N_12865,N_6423,N_9758);
nand U12866 (N_12866,N_7239,N_9008);
and U12867 (N_12867,N_6637,N_7792);
xnor U12868 (N_12868,N_6773,N_6578);
xnor U12869 (N_12869,N_5926,N_5194);
nand U12870 (N_12870,N_5856,N_6586);
nor U12871 (N_12871,N_6349,N_8208);
or U12872 (N_12872,N_5465,N_7273);
and U12873 (N_12873,N_6785,N_7471);
and U12874 (N_12874,N_8091,N_6243);
nor U12875 (N_12875,N_8030,N_7699);
and U12876 (N_12876,N_5992,N_6634);
xnor U12877 (N_12877,N_7237,N_7279);
or U12878 (N_12878,N_7193,N_7756);
nor U12879 (N_12879,N_5482,N_8106);
or U12880 (N_12880,N_5800,N_9006);
and U12881 (N_12881,N_7337,N_5700);
or U12882 (N_12882,N_7768,N_7954);
and U12883 (N_12883,N_6857,N_5112);
xor U12884 (N_12884,N_8479,N_6864);
and U12885 (N_12885,N_7275,N_6608);
and U12886 (N_12886,N_6492,N_8376);
and U12887 (N_12887,N_8357,N_8147);
nand U12888 (N_12888,N_9801,N_6444);
nand U12889 (N_12889,N_9138,N_7568);
or U12890 (N_12890,N_7461,N_7921);
or U12891 (N_12891,N_6130,N_6753);
nor U12892 (N_12892,N_9880,N_5292);
and U12893 (N_12893,N_6282,N_8846);
xnor U12894 (N_12894,N_7307,N_7936);
or U12895 (N_12895,N_5699,N_5179);
or U12896 (N_12896,N_9507,N_6973);
and U12897 (N_12897,N_6894,N_6303);
nand U12898 (N_12898,N_6898,N_5249);
nor U12899 (N_12899,N_8634,N_7364);
nand U12900 (N_12900,N_8954,N_5663);
xor U12901 (N_12901,N_7548,N_5251);
or U12902 (N_12902,N_5901,N_6489);
nor U12903 (N_12903,N_6955,N_7315);
xnor U12904 (N_12904,N_5588,N_5246);
or U12905 (N_12905,N_6438,N_5554);
and U12906 (N_12906,N_6312,N_9835);
nand U12907 (N_12907,N_7698,N_6660);
nor U12908 (N_12908,N_9722,N_8209);
nor U12909 (N_12909,N_8293,N_9687);
nor U12910 (N_12910,N_5309,N_6964);
and U12911 (N_12911,N_7598,N_5484);
nor U12912 (N_12912,N_9928,N_8913);
nor U12913 (N_12913,N_6490,N_8034);
and U12914 (N_12914,N_8880,N_5184);
or U12915 (N_12915,N_9526,N_9755);
nor U12916 (N_12916,N_6553,N_7696);
and U12917 (N_12917,N_5410,N_7874);
xnor U12918 (N_12918,N_7885,N_6159);
and U12919 (N_12919,N_9375,N_5782);
and U12920 (N_12920,N_5184,N_9225);
nor U12921 (N_12921,N_9000,N_8355);
or U12922 (N_12922,N_8004,N_6634);
or U12923 (N_12923,N_9435,N_7558);
nor U12924 (N_12924,N_5301,N_5500);
nand U12925 (N_12925,N_6409,N_6146);
and U12926 (N_12926,N_9591,N_8042);
xnor U12927 (N_12927,N_5587,N_8235);
or U12928 (N_12928,N_8757,N_9059);
xnor U12929 (N_12929,N_8686,N_5412);
and U12930 (N_12930,N_9645,N_6883);
nand U12931 (N_12931,N_5028,N_6443);
nand U12932 (N_12932,N_7494,N_5933);
nand U12933 (N_12933,N_9124,N_9506);
xnor U12934 (N_12934,N_9933,N_5739);
xor U12935 (N_12935,N_8935,N_6812);
and U12936 (N_12936,N_5403,N_8468);
and U12937 (N_12937,N_8170,N_9254);
or U12938 (N_12938,N_9017,N_9739);
and U12939 (N_12939,N_7190,N_7468);
nor U12940 (N_12940,N_7605,N_9084);
or U12941 (N_12941,N_6974,N_8042);
xor U12942 (N_12942,N_5045,N_5960);
nand U12943 (N_12943,N_8481,N_5335);
nor U12944 (N_12944,N_5759,N_5498);
nor U12945 (N_12945,N_6492,N_5701);
and U12946 (N_12946,N_8124,N_8254);
nor U12947 (N_12947,N_5175,N_8100);
xor U12948 (N_12948,N_6930,N_9561);
and U12949 (N_12949,N_7865,N_9869);
nand U12950 (N_12950,N_8676,N_5438);
nor U12951 (N_12951,N_9244,N_6554);
xnor U12952 (N_12952,N_7207,N_8409);
xor U12953 (N_12953,N_7614,N_8085);
nand U12954 (N_12954,N_6036,N_6056);
and U12955 (N_12955,N_5794,N_5635);
xnor U12956 (N_12956,N_6972,N_7243);
xnor U12957 (N_12957,N_6785,N_8063);
nor U12958 (N_12958,N_8394,N_7169);
nor U12959 (N_12959,N_6725,N_8329);
nand U12960 (N_12960,N_9548,N_7345);
nand U12961 (N_12961,N_7092,N_8315);
and U12962 (N_12962,N_7280,N_8108);
and U12963 (N_12963,N_8261,N_7679);
nand U12964 (N_12964,N_8276,N_9936);
nand U12965 (N_12965,N_6118,N_7148);
and U12966 (N_12966,N_6174,N_9837);
nand U12967 (N_12967,N_9750,N_7790);
nor U12968 (N_12968,N_8407,N_9392);
nor U12969 (N_12969,N_8946,N_5216);
nand U12970 (N_12970,N_9752,N_8622);
or U12971 (N_12971,N_9971,N_6161);
and U12972 (N_12972,N_5697,N_9755);
nor U12973 (N_12973,N_8519,N_8706);
and U12974 (N_12974,N_7500,N_6954);
or U12975 (N_12975,N_6373,N_6082);
nor U12976 (N_12976,N_6653,N_8822);
nor U12977 (N_12977,N_5242,N_7751);
xnor U12978 (N_12978,N_7154,N_6197);
nand U12979 (N_12979,N_9628,N_6070);
nor U12980 (N_12980,N_7307,N_8984);
nand U12981 (N_12981,N_5331,N_6263);
nor U12982 (N_12982,N_8237,N_8843);
or U12983 (N_12983,N_6207,N_8850);
or U12984 (N_12984,N_8588,N_6955);
and U12985 (N_12985,N_8249,N_5778);
and U12986 (N_12986,N_6498,N_8209);
or U12987 (N_12987,N_8269,N_5933);
nand U12988 (N_12988,N_7245,N_9807);
xor U12989 (N_12989,N_9810,N_8525);
and U12990 (N_12990,N_6217,N_5514);
nor U12991 (N_12991,N_6430,N_9347);
and U12992 (N_12992,N_6181,N_5575);
or U12993 (N_12993,N_8375,N_7445);
nor U12994 (N_12994,N_5686,N_9895);
nand U12995 (N_12995,N_7065,N_5578);
xnor U12996 (N_12996,N_6260,N_9777);
and U12997 (N_12997,N_8991,N_6004);
nor U12998 (N_12998,N_8034,N_8953);
and U12999 (N_12999,N_6989,N_5799);
nor U13000 (N_13000,N_9219,N_9692);
nand U13001 (N_13001,N_9743,N_6038);
and U13002 (N_13002,N_8719,N_9741);
nor U13003 (N_13003,N_8101,N_5151);
and U13004 (N_13004,N_5037,N_9599);
nor U13005 (N_13005,N_7995,N_6273);
or U13006 (N_13006,N_8742,N_5490);
nor U13007 (N_13007,N_6045,N_5423);
nor U13008 (N_13008,N_8401,N_5140);
nand U13009 (N_13009,N_5733,N_7960);
nand U13010 (N_13010,N_9103,N_8976);
nor U13011 (N_13011,N_7813,N_6661);
and U13012 (N_13012,N_5094,N_5229);
or U13013 (N_13013,N_7340,N_7049);
xor U13014 (N_13014,N_7384,N_7013);
or U13015 (N_13015,N_9638,N_9174);
or U13016 (N_13016,N_7802,N_6444);
nand U13017 (N_13017,N_8619,N_6895);
xnor U13018 (N_13018,N_9016,N_5473);
or U13019 (N_13019,N_9118,N_7292);
nand U13020 (N_13020,N_9431,N_7278);
or U13021 (N_13021,N_7223,N_5491);
xnor U13022 (N_13022,N_9461,N_6285);
or U13023 (N_13023,N_6450,N_8651);
or U13024 (N_13024,N_7467,N_5412);
nor U13025 (N_13025,N_5205,N_5580);
and U13026 (N_13026,N_9669,N_6077);
nor U13027 (N_13027,N_8862,N_9653);
and U13028 (N_13028,N_7390,N_6695);
xor U13029 (N_13029,N_6809,N_9555);
nor U13030 (N_13030,N_9679,N_8188);
nor U13031 (N_13031,N_8862,N_5952);
and U13032 (N_13032,N_8756,N_9194);
nand U13033 (N_13033,N_8315,N_9482);
nand U13034 (N_13034,N_8862,N_8332);
and U13035 (N_13035,N_8847,N_9235);
and U13036 (N_13036,N_9176,N_5652);
nor U13037 (N_13037,N_8764,N_7649);
and U13038 (N_13038,N_5879,N_7954);
nor U13039 (N_13039,N_5506,N_6859);
xnor U13040 (N_13040,N_9463,N_9158);
nor U13041 (N_13041,N_8536,N_6990);
nor U13042 (N_13042,N_9337,N_6608);
nor U13043 (N_13043,N_7119,N_5490);
nor U13044 (N_13044,N_6916,N_7568);
nand U13045 (N_13045,N_6980,N_7627);
or U13046 (N_13046,N_9511,N_7514);
or U13047 (N_13047,N_9176,N_7297);
nand U13048 (N_13048,N_5256,N_6631);
xnor U13049 (N_13049,N_7150,N_6354);
nor U13050 (N_13050,N_5998,N_6638);
xor U13051 (N_13051,N_6985,N_7376);
nor U13052 (N_13052,N_8853,N_8398);
nand U13053 (N_13053,N_5691,N_6835);
nor U13054 (N_13054,N_9454,N_9289);
and U13055 (N_13055,N_8472,N_5848);
xor U13056 (N_13056,N_8876,N_8037);
and U13057 (N_13057,N_5307,N_7080);
nor U13058 (N_13058,N_5999,N_5781);
xor U13059 (N_13059,N_5252,N_7967);
or U13060 (N_13060,N_8062,N_9181);
or U13061 (N_13061,N_5544,N_5202);
xnor U13062 (N_13062,N_7004,N_5322);
nor U13063 (N_13063,N_8299,N_8354);
xnor U13064 (N_13064,N_8245,N_6259);
and U13065 (N_13065,N_5821,N_7343);
nor U13066 (N_13066,N_7107,N_6085);
nor U13067 (N_13067,N_5434,N_5401);
and U13068 (N_13068,N_8760,N_8565);
nand U13069 (N_13069,N_9171,N_5248);
nand U13070 (N_13070,N_9554,N_5238);
or U13071 (N_13071,N_8485,N_7917);
xor U13072 (N_13072,N_8553,N_6597);
nand U13073 (N_13073,N_6661,N_8172);
and U13074 (N_13074,N_5531,N_6012);
xor U13075 (N_13075,N_6354,N_6812);
or U13076 (N_13076,N_7677,N_8035);
nor U13077 (N_13077,N_8438,N_8979);
and U13078 (N_13078,N_6295,N_5246);
xor U13079 (N_13079,N_9502,N_9811);
nor U13080 (N_13080,N_7354,N_8965);
nand U13081 (N_13081,N_7827,N_9353);
xnor U13082 (N_13082,N_5197,N_7927);
and U13083 (N_13083,N_5310,N_8132);
and U13084 (N_13084,N_5838,N_5331);
nand U13085 (N_13085,N_5085,N_7237);
xor U13086 (N_13086,N_7647,N_5945);
or U13087 (N_13087,N_7593,N_6185);
or U13088 (N_13088,N_6228,N_8813);
nand U13089 (N_13089,N_5300,N_9036);
nor U13090 (N_13090,N_6141,N_7298);
nor U13091 (N_13091,N_9859,N_7868);
and U13092 (N_13092,N_9606,N_7241);
or U13093 (N_13093,N_6726,N_8746);
and U13094 (N_13094,N_9204,N_5617);
xor U13095 (N_13095,N_9605,N_8155);
xnor U13096 (N_13096,N_9956,N_8022);
and U13097 (N_13097,N_8301,N_5951);
xor U13098 (N_13098,N_7138,N_9966);
nand U13099 (N_13099,N_5741,N_9957);
nand U13100 (N_13100,N_8707,N_8962);
or U13101 (N_13101,N_9513,N_7160);
or U13102 (N_13102,N_5031,N_7361);
or U13103 (N_13103,N_6243,N_6963);
xor U13104 (N_13104,N_8759,N_8138);
xor U13105 (N_13105,N_5771,N_7041);
nor U13106 (N_13106,N_5822,N_5690);
or U13107 (N_13107,N_9279,N_6482);
nand U13108 (N_13108,N_6194,N_9562);
nand U13109 (N_13109,N_5853,N_8263);
or U13110 (N_13110,N_5506,N_5760);
nor U13111 (N_13111,N_6267,N_9231);
and U13112 (N_13112,N_9798,N_9405);
or U13113 (N_13113,N_7016,N_7770);
and U13114 (N_13114,N_8480,N_7328);
xor U13115 (N_13115,N_5007,N_5548);
and U13116 (N_13116,N_5392,N_9220);
xor U13117 (N_13117,N_5908,N_9575);
nor U13118 (N_13118,N_6530,N_8552);
nor U13119 (N_13119,N_9154,N_5999);
and U13120 (N_13120,N_5314,N_5384);
or U13121 (N_13121,N_8245,N_6629);
and U13122 (N_13122,N_6104,N_9745);
nand U13123 (N_13123,N_9585,N_5831);
nand U13124 (N_13124,N_8988,N_8962);
and U13125 (N_13125,N_7624,N_5300);
or U13126 (N_13126,N_5763,N_6403);
nor U13127 (N_13127,N_5626,N_8374);
xor U13128 (N_13128,N_9762,N_9593);
and U13129 (N_13129,N_6009,N_7814);
or U13130 (N_13130,N_8289,N_9838);
xnor U13131 (N_13131,N_5552,N_9159);
and U13132 (N_13132,N_6372,N_9359);
xnor U13133 (N_13133,N_7030,N_6808);
nor U13134 (N_13134,N_5972,N_5525);
nor U13135 (N_13135,N_8075,N_7422);
and U13136 (N_13136,N_8454,N_6224);
xor U13137 (N_13137,N_5065,N_6271);
or U13138 (N_13138,N_8933,N_7277);
and U13139 (N_13139,N_7421,N_5307);
and U13140 (N_13140,N_9924,N_7174);
xor U13141 (N_13141,N_6218,N_9096);
nand U13142 (N_13142,N_9328,N_7471);
xor U13143 (N_13143,N_6952,N_6528);
nor U13144 (N_13144,N_6549,N_6390);
and U13145 (N_13145,N_7234,N_5132);
xnor U13146 (N_13146,N_6296,N_5366);
nor U13147 (N_13147,N_8872,N_7565);
nor U13148 (N_13148,N_9783,N_8630);
and U13149 (N_13149,N_7454,N_8827);
xor U13150 (N_13150,N_8901,N_7828);
and U13151 (N_13151,N_9528,N_6173);
xor U13152 (N_13152,N_9411,N_9898);
xor U13153 (N_13153,N_5952,N_6269);
nand U13154 (N_13154,N_9304,N_8499);
xnor U13155 (N_13155,N_6642,N_5606);
nor U13156 (N_13156,N_8741,N_7432);
xor U13157 (N_13157,N_6718,N_9327);
or U13158 (N_13158,N_7137,N_8114);
and U13159 (N_13159,N_7367,N_5564);
nand U13160 (N_13160,N_6479,N_9039);
xnor U13161 (N_13161,N_8013,N_8157);
or U13162 (N_13162,N_7835,N_8006);
nand U13163 (N_13163,N_7584,N_7485);
xnor U13164 (N_13164,N_9856,N_6647);
nand U13165 (N_13165,N_8461,N_6531);
nor U13166 (N_13166,N_6567,N_9626);
xor U13167 (N_13167,N_9699,N_5577);
or U13168 (N_13168,N_9245,N_8039);
nand U13169 (N_13169,N_7414,N_7530);
nor U13170 (N_13170,N_6241,N_8414);
xnor U13171 (N_13171,N_9716,N_9593);
or U13172 (N_13172,N_8661,N_7719);
xor U13173 (N_13173,N_5493,N_5832);
nor U13174 (N_13174,N_8030,N_9047);
nand U13175 (N_13175,N_6983,N_6149);
nand U13176 (N_13176,N_7504,N_7028);
nor U13177 (N_13177,N_6420,N_6182);
and U13178 (N_13178,N_7296,N_7482);
and U13179 (N_13179,N_5908,N_8401);
nor U13180 (N_13180,N_6216,N_9526);
nor U13181 (N_13181,N_9646,N_7824);
xor U13182 (N_13182,N_8412,N_5220);
nand U13183 (N_13183,N_5227,N_7142);
and U13184 (N_13184,N_9036,N_8604);
or U13185 (N_13185,N_6648,N_5726);
nand U13186 (N_13186,N_9440,N_8270);
xnor U13187 (N_13187,N_5573,N_7965);
or U13188 (N_13188,N_7095,N_6411);
and U13189 (N_13189,N_5626,N_7444);
nor U13190 (N_13190,N_8335,N_6865);
xnor U13191 (N_13191,N_8779,N_7985);
and U13192 (N_13192,N_6761,N_8248);
nor U13193 (N_13193,N_6013,N_8409);
nor U13194 (N_13194,N_6738,N_5555);
and U13195 (N_13195,N_9014,N_5385);
nand U13196 (N_13196,N_6444,N_7554);
nor U13197 (N_13197,N_5366,N_8051);
nand U13198 (N_13198,N_5376,N_7011);
nor U13199 (N_13199,N_7850,N_7028);
nor U13200 (N_13200,N_6634,N_5752);
xor U13201 (N_13201,N_6993,N_6524);
or U13202 (N_13202,N_8977,N_8759);
nand U13203 (N_13203,N_7722,N_7350);
xnor U13204 (N_13204,N_8576,N_7172);
xor U13205 (N_13205,N_8342,N_7036);
and U13206 (N_13206,N_7290,N_8668);
nand U13207 (N_13207,N_5021,N_7418);
and U13208 (N_13208,N_6901,N_9875);
and U13209 (N_13209,N_6632,N_9542);
xnor U13210 (N_13210,N_5065,N_9657);
nor U13211 (N_13211,N_8419,N_7753);
nand U13212 (N_13212,N_8262,N_9941);
nand U13213 (N_13213,N_9507,N_5214);
nor U13214 (N_13214,N_5056,N_8164);
nor U13215 (N_13215,N_8450,N_5825);
and U13216 (N_13216,N_8583,N_7946);
nand U13217 (N_13217,N_5848,N_9746);
xor U13218 (N_13218,N_6171,N_5213);
and U13219 (N_13219,N_6291,N_6490);
nor U13220 (N_13220,N_6316,N_6138);
xnor U13221 (N_13221,N_5979,N_5724);
nor U13222 (N_13222,N_9069,N_5426);
nor U13223 (N_13223,N_7591,N_6595);
nor U13224 (N_13224,N_6646,N_8990);
or U13225 (N_13225,N_5710,N_8935);
and U13226 (N_13226,N_6226,N_7111);
xnor U13227 (N_13227,N_7683,N_9129);
nor U13228 (N_13228,N_9223,N_9951);
nor U13229 (N_13229,N_5349,N_7275);
nor U13230 (N_13230,N_5714,N_6634);
or U13231 (N_13231,N_6970,N_9104);
nand U13232 (N_13232,N_6650,N_5055);
nand U13233 (N_13233,N_9268,N_6046);
nand U13234 (N_13234,N_7783,N_9995);
nor U13235 (N_13235,N_6402,N_9937);
nor U13236 (N_13236,N_5476,N_7037);
nor U13237 (N_13237,N_6131,N_9888);
nor U13238 (N_13238,N_6577,N_7683);
nor U13239 (N_13239,N_7600,N_5082);
xnor U13240 (N_13240,N_9718,N_5612);
and U13241 (N_13241,N_6416,N_9836);
or U13242 (N_13242,N_9807,N_7287);
and U13243 (N_13243,N_7511,N_6714);
xor U13244 (N_13244,N_8105,N_6261);
and U13245 (N_13245,N_9233,N_7779);
nor U13246 (N_13246,N_8589,N_8475);
nand U13247 (N_13247,N_5982,N_9404);
and U13248 (N_13248,N_9101,N_5074);
nor U13249 (N_13249,N_8414,N_6550);
nor U13250 (N_13250,N_9488,N_7972);
nor U13251 (N_13251,N_9974,N_6749);
or U13252 (N_13252,N_5496,N_9745);
xor U13253 (N_13253,N_6139,N_9541);
nor U13254 (N_13254,N_5617,N_7350);
nand U13255 (N_13255,N_9548,N_5409);
xor U13256 (N_13256,N_5374,N_8325);
nor U13257 (N_13257,N_9112,N_8536);
and U13258 (N_13258,N_5088,N_5049);
xnor U13259 (N_13259,N_7038,N_6646);
nand U13260 (N_13260,N_8311,N_7254);
xnor U13261 (N_13261,N_7563,N_9381);
and U13262 (N_13262,N_9381,N_6456);
and U13263 (N_13263,N_8039,N_5918);
nor U13264 (N_13264,N_6657,N_8743);
and U13265 (N_13265,N_7651,N_9574);
or U13266 (N_13266,N_7636,N_9520);
or U13267 (N_13267,N_9417,N_8891);
xnor U13268 (N_13268,N_7334,N_5311);
or U13269 (N_13269,N_9775,N_6375);
nand U13270 (N_13270,N_5509,N_8013);
nor U13271 (N_13271,N_9004,N_7897);
nand U13272 (N_13272,N_5582,N_8883);
xor U13273 (N_13273,N_8110,N_5625);
nor U13274 (N_13274,N_5347,N_6534);
nor U13275 (N_13275,N_9155,N_9612);
and U13276 (N_13276,N_6890,N_5324);
xor U13277 (N_13277,N_7600,N_7298);
nor U13278 (N_13278,N_8687,N_6249);
xnor U13279 (N_13279,N_5036,N_8766);
xor U13280 (N_13280,N_6461,N_9818);
nor U13281 (N_13281,N_7186,N_9156);
and U13282 (N_13282,N_9763,N_5085);
xor U13283 (N_13283,N_5189,N_5752);
xnor U13284 (N_13284,N_8380,N_8164);
xnor U13285 (N_13285,N_6252,N_5410);
or U13286 (N_13286,N_5442,N_7853);
or U13287 (N_13287,N_7984,N_6145);
and U13288 (N_13288,N_6087,N_6515);
and U13289 (N_13289,N_6730,N_9464);
and U13290 (N_13290,N_6011,N_6211);
nor U13291 (N_13291,N_8508,N_7573);
nor U13292 (N_13292,N_9211,N_8696);
and U13293 (N_13293,N_7391,N_5258);
nor U13294 (N_13294,N_5178,N_6043);
or U13295 (N_13295,N_5815,N_7555);
nand U13296 (N_13296,N_5151,N_5103);
nand U13297 (N_13297,N_9466,N_9125);
and U13298 (N_13298,N_8579,N_9044);
xnor U13299 (N_13299,N_5621,N_6146);
nor U13300 (N_13300,N_6600,N_6447);
xnor U13301 (N_13301,N_8085,N_9079);
and U13302 (N_13302,N_9862,N_9026);
nor U13303 (N_13303,N_5038,N_8732);
and U13304 (N_13304,N_8436,N_8042);
nor U13305 (N_13305,N_9074,N_5200);
and U13306 (N_13306,N_5265,N_9176);
nor U13307 (N_13307,N_7487,N_7058);
or U13308 (N_13308,N_8992,N_9568);
nand U13309 (N_13309,N_7928,N_5435);
nor U13310 (N_13310,N_5531,N_6499);
xor U13311 (N_13311,N_9829,N_9254);
xnor U13312 (N_13312,N_5442,N_9842);
xor U13313 (N_13313,N_6665,N_5520);
nor U13314 (N_13314,N_7228,N_9892);
or U13315 (N_13315,N_6237,N_5180);
nand U13316 (N_13316,N_9205,N_5111);
and U13317 (N_13317,N_5645,N_8290);
nor U13318 (N_13318,N_5409,N_5475);
and U13319 (N_13319,N_7847,N_5899);
nor U13320 (N_13320,N_9505,N_8138);
nand U13321 (N_13321,N_7941,N_7335);
and U13322 (N_13322,N_9283,N_6701);
or U13323 (N_13323,N_7372,N_9333);
xnor U13324 (N_13324,N_5824,N_8502);
nor U13325 (N_13325,N_6879,N_9498);
xnor U13326 (N_13326,N_8802,N_8795);
nand U13327 (N_13327,N_6895,N_9791);
or U13328 (N_13328,N_9306,N_9177);
and U13329 (N_13329,N_6936,N_9607);
or U13330 (N_13330,N_8514,N_6965);
nor U13331 (N_13331,N_9531,N_5997);
and U13332 (N_13332,N_6565,N_5234);
nor U13333 (N_13333,N_8126,N_7434);
or U13334 (N_13334,N_8015,N_8152);
nand U13335 (N_13335,N_9800,N_8627);
and U13336 (N_13336,N_8669,N_8047);
and U13337 (N_13337,N_7242,N_5606);
xor U13338 (N_13338,N_6337,N_5665);
and U13339 (N_13339,N_9199,N_9787);
nand U13340 (N_13340,N_9742,N_5284);
or U13341 (N_13341,N_9459,N_5427);
xnor U13342 (N_13342,N_6922,N_9692);
xnor U13343 (N_13343,N_8942,N_5850);
xor U13344 (N_13344,N_9894,N_6628);
nand U13345 (N_13345,N_9063,N_5718);
and U13346 (N_13346,N_7758,N_5772);
nor U13347 (N_13347,N_6081,N_6984);
xnor U13348 (N_13348,N_6173,N_7227);
xnor U13349 (N_13349,N_6310,N_7673);
nor U13350 (N_13350,N_8242,N_6720);
or U13351 (N_13351,N_9843,N_8310);
nor U13352 (N_13352,N_6032,N_9066);
nand U13353 (N_13353,N_7989,N_6460);
nand U13354 (N_13354,N_6515,N_8930);
xnor U13355 (N_13355,N_5628,N_6617);
nand U13356 (N_13356,N_7125,N_7686);
and U13357 (N_13357,N_6392,N_9893);
nor U13358 (N_13358,N_6661,N_5495);
nor U13359 (N_13359,N_8678,N_8755);
xor U13360 (N_13360,N_8631,N_5273);
and U13361 (N_13361,N_8956,N_7797);
xor U13362 (N_13362,N_8507,N_7202);
and U13363 (N_13363,N_5708,N_8238);
nor U13364 (N_13364,N_7737,N_9472);
or U13365 (N_13365,N_8240,N_9665);
nand U13366 (N_13366,N_8698,N_7880);
and U13367 (N_13367,N_5757,N_8866);
xor U13368 (N_13368,N_5372,N_8955);
or U13369 (N_13369,N_8946,N_9255);
nor U13370 (N_13370,N_7957,N_8812);
xor U13371 (N_13371,N_5762,N_6924);
nor U13372 (N_13372,N_7277,N_7714);
nor U13373 (N_13373,N_5432,N_6202);
and U13374 (N_13374,N_5963,N_8498);
nor U13375 (N_13375,N_7888,N_5827);
and U13376 (N_13376,N_5778,N_9369);
and U13377 (N_13377,N_6602,N_7770);
and U13378 (N_13378,N_9810,N_9355);
or U13379 (N_13379,N_6085,N_6735);
nand U13380 (N_13380,N_8002,N_6176);
and U13381 (N_13381,N_8535,N_8531);
and U13382 (N_13382,N_9443,N_8878);
nand U13383 (N_13383,N_5416,N_6030);
or U13384 (N_13384,N_7304,N_7107);
nor U13385 (N_13385,N_7236,N_7303);
and U13386 (N_13386,N_6636,N_5759);
nor U13387 (N_13387,N_6568,N_5168);
and U13388 (N_13388,N_7247,N_9609);
and U13389 (N_13389,N_6256,N_6117);
nor U13390 (N_13390,N_7505,N_5586);
or U13391 (N_13391,N_8935,N_7577);
or U13392 (N_13392,N_9044,N_5753);
and U13393 (N_13393,N_9621,N_5484);
nand U13394 (N_13394,N_7747,N_9392);
and U13395 (N_13395,N_5272,N_5690);
nand U13396 (N_13396,N_9228,N_9116);
nand U13397 (N_13397,N_5953,N_9306);
xor U13398 (N_13398,N_6928,N_9363);
or U13399 (N_13399,N_9472,N_6711);
nand U13400 (N_13400,N_6513,N_5765);
nand U13401 (N_13401,N_9124,N_9983);
nand U13402 (N_13402,N_7580,N_8754);
xnor U13403 (N_13403,N_8546,N_7897);
xor U13404 (N_13404,N_5233,N_9438);
nand U13405 (N_13405,N_6079,N_6269);
or U13406 (N_13406,N_8377,N_5760);
nand U13407 (N_13407,N_6804,N_5285);
xnor U13408 (N_13408,N_6857,N_6220);
or U13409 (N_13409,N_5226,N_7257);
nand U13410 (N_13410,N_9742,N_6085);
or U13411 (N_13411,N_7384,N_5254);
xor U13412 (N_13412,N_8922,N_9983);
nand U13413 (N_13413,N_9636,N_5129);
nand U13414 (N_13414,N_9510,N_5460);
xnor U13415 (N_13415,N_8778,N_8432);
nand U13416 (N_13416,N_5836,N_6922);
nand U13417 (N_13417,N_8601,N_6961);
and U13418 (N_13418,N_9601,N_6460);
and U13419 (N_13419,N_8571,N_5736);
nor U13420 (N_13420,N_9945,N_7107);
and U13421 (N_13421,N_6004,N_9166);
nor U13422 (N_13422,N_6342,N_7507);
xor U13423 (N_13423,N_5284,N_5668);
nand U13424 (N_13424,N_8513,N_9287);
nand U13425 (N_13425,N_8521,N_9919);
or U13426 (N_13426,N_5239,N_7170);
xnor U13427 (N_13427,N_9261,N_8431);
nor U13428 (N_13428,N_5287,N_7988);
and U13429 (N_13429,N_9345,N_9316);
and U13430 (N_13430,N_9018,N_5949);
and U13431 (N_13431,N_9127,N_6145);
nand U13432 (N_13432,N_9547,N_8312);
nand U13433 (N_13433,N_5877,N_5171);
nor U13434 (N_13434,N_7248,N_5787);
xor U13435 (N_13435,N_8482,N_9634);
or U13436 (N_13436,N_9262,N_7726);
nor U13437 (N_13437,N_6642,N_9823);
and U13438 (N_13438,N_5916,N_8625);
xor U13439 (N_13439,N_6219,N_9073);
xor U13440 (N_13440,N_5797,N_5975);
xnor U13441 (N_13441,N_9355,N_9504);
xnor U13442 (N_13442,N_7635,N_7303);
xnor U13443 (N_13443,N_6221,N_5001);
nor U13444 (N_13444,N_9584,N_9914);
nor U13445 (N_13445,N_9262,N_8420);
and U13446 (N_13446,N_8913,N_7702);
or U13447 (N_13447,N_8140,N_7209);
nor U13448 (N_13448,N_7895,N_5399);
and U13449 (N_13449,N_8230,N_9164);
nand U13450 (N_13450,N_7779,N_6040);
and U13451 (N_13451,N_6531,N_7426);
or U13452 (N_13452,N_8886,N_8248);
and U13453 (N_13453,N_9429,N_9404);
nand U13454 (N_13454,N_8090,N_5612);
nand U13455 (N_13455,N_5856,N_9337);
nor U13456 (N_13456,N_7360,N_5722);
nand U13457 (N_13457,N_8005,N_6629);
nand U13458 (N_13458,N_6893,N_7306);
and U13459 (N_13459,N_9259,N_6588);
or U13460 (N_13460,N_9761,N_8437);
nand U13461 (N_13461,N_8294,N_6720);
nand U13462 (N_13462,N_9117,N_9163);
xnor U13463 (N_13463,N_6487,N_7159);
and U13464 (N_13464,N_5303,N_7738);
nor U13465 (N_13465,N_5262,N_5278);
or U13466 (N_13466,N_5992,N_7428);
and U13467 (N_13467,N_8871,N_6939);
or U13468 (N_13468,N_9905,N_6542);
xor U13469 (N_13469,N_6630,N_8758);
xnor U13470 (N_13470,N_6250,N_5729);
nand U13471 (N_13471,N_6490,N_9349);
xor U13472 (N_13472,N_8385,N_9857);
nand U13473 (N_13473,N_6238,N_5092);
xor U13474 (N_13474,N_5944,N_8940);
or U13475 (N_13475,N_5637,N_7254);
and U13476 (N_13476,N_8704,N_9243);
nor U13477 (N_13477,N_8711,N_6644);
and U13478 (N_13478,N_8524,N_8291);
nor U13479 (N_13479,N_6432,N_9348);
nor U13480 (N_13480,N_9893,N_9381);
or U13481 (N_13481,N_7680,N_7193);
nand U13482 (N_13482,N_9985,N_8763);
nor U13483 (N_13483,N_9933,N_5395);
xor U13484 (N_13484,N_6749,N_8784);
nand U13485 (N_13485,N_8294,N_5501);
nor U13486 (N_13486,N_8056,N_7993);
and U13487 (N_13487,N_9427,N_9207);
xnor U13488 (N_13488,N_9246,N_5061);
nor U13489 (N_13489,N_6140,N_8936);
nor U13490 (N_13490,N_7641,N_6092);
and U13491 (N_13491,N_8893,N_6017);
xnor U13492 (N_13492,N_7326,N_9833);
or U13493 (N_13493,N_5065,N_8554);
and U13494 (N_13494,N_7425,N_7482);
or U13495 (N_13495,N_7883,N_9014);
xor U13496 (N_13496,N_5650,N_6674);
or U13497 (N_13497,N_5880,N_5098);
nand U13498 (N_13498,N_9864,N_7329);
xnor U13499 (N_13499,N_8583,N_9520);
nand U13500 (N_13500,N_8959,N_7897);
nand U13501 (N_13501,N_5205,N_9396);
or U13502 (N_13502,N_6878,N_9708);
xnor U13503 (N_13503,N_8550,N_9190);
and U13504 (N_13504,N_7583,N_5683);
and U13505 (N_13505,N_6709,N_9328);
or U13506 (N_13506,N_8493,N_6391);
and U13507 (N_13507,N_8735,N_6174);
nor U13508 (N_13508,N_6331,N_6274);
nor U13509 (N_13509,N_8403,N_9962);
xnor U13510 (N_13510,N_7085,N_9361);
and U13511 (N_13511,N_6543,N_6251);
nor U13512 (N_13512,N_9947,N_7970);
xnor U13513 (N_13513,N_9053,N_8909);
xnor U13514 (N_13514,N_8773,N_7474);
and U13515 (N_13515,N_6740,N_6267);
xor U13516 (N_13516,N_8414,N_9277);
and U13517 (N_13517,N_7990,N_5407);
xor U13518 (N_13518,N_6059,N_8800);
nor U13519 (N_13519,N_5835,N_9104);
and U13520 (N_13520,N_9639,N_7666);
xnor U13521 (N_13521,N_7092,N_7746);
nor U13522 (N_13522,N_6228,N_8788);
xor U13523 (N_13523,N_7916,N_6185);
or U13524 (N_13524,N_8794,N_6893);
nand U13525 (N_13525,N_6987,N_8783);
nand U13526 (N_13526,N_8569,N_7657);
and U13527 (N_13527,N_8244,N_8582);
and U13528 (N_13528,N_5670,N_9957);
nor U13529 (N_13529,N_6744,N_9713);
nand U13530 (N_13530,N_6382,N_9530);
nand U13531 (N_13531,N_6010,N_7322);
xnor U13532 (N_13532,N_5359,N_6864);
xnor U13533 (N_13533,N_6139,N_8395);
nor U13534 (N_13534,N_8083,N_8248);
nor U13535 (N_13535,N_8716,N_9362);
nand U13536 (N_13536,N_5484,N_7192);
nor U13537 (N_13537,N_5465,N_5247);
or U13538 (N_13538,N_9559,N_7510);
and U13539 (N_13539,N_8556,N_8352);
nor U13540 (N_13540,N_9924,N_7183);
nor U13541 (N_13541,N_9557,N_5659);
and U13542 (N_13542,N_7270,N_7004);
xnor U13543 (N_13543,N_7591,N_7862);
xnor U13544 (N_13544,N_8610,N_8709);
xnor U13545 (N_13545,N_7598,N_7886);
nand U13546 (N_13546,N_6596,N_7602);
nand U13547 (N_13547,N_8474,N_9886);
xnor U13548 (N_13548,N_9306,N_9099);
nand U13549 (N_13549,N_6225,N_8340);
nor U13550 (N_13550,N_7154,N_6991);
and U13551 (N_13551,N_5156,N_6066);
xor U13552 (N_13552,N_5475,N_5299);
and U13553 (N_13553,N_5158,N_8239);
nor U13554 (N_13554,N_5834,N_8152);
or U13555 (N_13555,N_9774,N_5811);
and U13556 (N_13556,N_8911,N_8347);
or U13557 (N_13557,N_6051,N_8503);
and U13558 (N_13558,N_6174,N_5714);
xor U13559 (N_13559,N_6744,N_8612);
and U13560 (N_13560,N_7282,N_6337);
or U13561 (N_13561,N_9422,N_7554);
nor U13562 (N_13562,N_7668,N_7221);
and U13563 (N_13563,N_5946,N_6897);
nor U13564 (N_13564,N_5904,N_8007);
and U13565 (N_13565,N_5021,N_8068);
xor U13566 (N_13566,N_6784,N_9699);
xnor U13567 (N_13567,N_6127,N_8600);
nor U13568 (N_13568,N_8456,N_5255);
xnor U13569 (N_13569,N_6739,N_9013);
or U13570 (N_13570,N_8800,N_7985);
nor U13571 (N_13571,N_7610,N_6062);
nor U13572 (N_13572,N_8631,N_7489);
nor U13573 (N_13573,N_6505,N_6711);
or U13574 (N_13574,N_5706,N_5473);
or U13575 (N_13575,N_8746,N_5475);
xnor U13576 (N_13576,N_9964,N_7918);
nand U13577 (N_13577,N_5159,N_5385);
xor U13578 (N_13578,N_7949,N_9264);
or U13579 (N_13579,N_7388,N_8432);
nand U13580 (N_13580,N_9732,N_5231);
nand U13581 (N_13581,N_9292,N_7805);
nor U13582 (N_13582,N_6190,N_8900);
or U13583 (N_13583,N_5253,N_8695);
and U13584 (N_13584,N_6320,N_6564);
xor U13585 (N_13585,N_7806,N_5728);
xor U13586 (N_13586,N_7966,N_6799);
nand U13587 (N_13587,N_5384,N_6328);
nand U13588 (N_13588,N_6161,N_9456);
nand U13589 (N_13589,N_6480,N_6411);
xor U13590 (N_13590,N_5829,N_8541);
nand U13591 (N_13591,N_9622,N_8804);
nor U13592 (N_13592,N_7357,N_9103);
nand U13593 (N_13593,N_5414,N_6502);
nor U13594 (N_13594,N_8091,N_8793);
nand U13595 (N_13595,N_6021,N_5813);
or U13596 (N_13596,N_8981,N_7617);
xnor U13597 (N_13597,N_7357,N_8302);
and U13598 (N_13598,N_7748,N_9112);
nor U13599 (N_13599,N_7725,N_5333);
and U13600 (N_13600,N_9508,N_8900);
or U13601 (N_13601,N_8725,N_9435);
and U13602 (N_13602,N_6539,N_7317);
xnor U13603 (N_13603,N_8314,N_9787);
nand U13604 (N_13604,N_6130,N_5350);
nand U13605 (N_13605,N_7929,N_5021);
nand U13606 (N_13606,N_7060,N_8448);
nor U13607 (N_13607,N_9700,N_8543);
and U13608 (N_13608,N_5907,N_8686);
and U13609 (N_13609,N_9853,N_8139);
nor U13610 (N_13610,N_6770,N_6793);
nor U13611 (N_13611,N_8418,N_7067);
xnor U13612 (N_13612,N_8843,N_9532);
nor U13613 (N_13613,N_5370,N_8709);
nand U13614 (N_13614,N_5894,N_5118);
or U13615 (N_13615,N_8646,N_5216);
nand U13616 (N_13616,N_6606,N_6552);
or U13617 (N_13617,N_9242,N_5860);
and U13618 (N_13618,N_7534,N_5053);
or U13619 (N_13619,N_8106,N_8553);
nor U13620 (N_13620,N_6498,N_5691);
xor U13621 (N_13621,N_8817,N_7103);
nor U13622 (N_13622,N_8608,N_7655);
or U13623 (N_13623,N_5563,N_6964);
or U13624 (N_13624,N_6778,N_7344);
or U13625 (N_13625,N_5096,N_5416);
nand U13626 (N_13626,N_6218,N_8887);
and U13627 (N_13627,N_6273,N_6093);
xor U13628 (N_13628,N_6039,N_5663);
nand U13629 (N_13629,N_6749,N_7723);
nand U13630 (N_13630,N_7545,N_7750);
nor U13631 (N_13631,N_5269,N_9862);
and U13632 (N_13632,N_9347,N_5805);
nor U13633 (N_13633,N_9870,N_6933);
or U13634 (N_13634,N_5441,N_8374);
or U13635 (N_13635,N_9466,N_6099);
or U13636 (N_13636,N_8306,N_8021);
nor U13637 (N_13637,N_7483,N_9419);
and U13638 (N_13638,N_5858,N_6193);
xor U13639 (N_13639,N_5506,N_6675);
and U13640 (N_13640,N_7878,N_8395);
xor U13641 (N_13641,N_5872,N_7503);
xor U13642 (N_13642,N_8751,N_7605);
and U13643 (N_13643,N_9547,N_7234);
or U13644 (N_13644,N_7070,N_8742);
and U13645 (N_13645,N_8088,N_9197);
or U13646 (N_13646,N_6022,N_7211);
nand U13647 (N_13647,N_9653,N_7811);
or U13648 (N_13648,N_8966,N_5669);
nor U13649 (N_13649,N_6559,N_8409);
xor U13650 (N_13650,N_8707,N_9744);
or U13651 (N_13651,N_8476,N_8725);
or U13652 (N_13652,N_6402,N_5851);
nor U13653 (N_13653,N_5518,N_8499);
nand U13654 (N_13654,N_7362,N_6687);
nand U13655 (N_13655,N_5423,N_8292);
nor U13656 (N_13656,N_8360,N_8411);
nand U13657 (N_13657,N_9152,N_6549);
nand U13658 (N_13658,N_7884,N_6172);
or U13659 (N_13659,N_8614,N_9433);
and U13660 (N_13660,N_5167,N_7901);
and U13661 (N_13661,N_6196,N_8621);
or U13662 (N_13662,N_5439,N_7710);
and U13663 (N_13663,N_6013,N_9331);
nor U13664 (N_13664,N_8652,N_7537);
or U13665 (N_13665,N_9436,N_9730);
and U13666 (N_13666,N_8167,N_7318);
nand U13667 (N_13667,N_9907,N_8793);
or U13668 (N_13668,N_7890,N_7424);
or U13669 (N_13669,N_6704,N_7428);
xnor U13670 (N_13670,N_5503,N_8652);
nor U13671 (N_13671,N_9559,N_8317);
nand U13672 (N_13672,N_9364,N_6272);
or U13673 (N_13673,N_6021,N_7165);
and U13674 (N_13674,N_9847,N_5138);
xor U13675 (N_13675,N_6401,N_6026);
nor U13676 (N_13676,N_9449,N_8607);
xnor U13677 (N_13677,N_7872,N_9647);
and U13678 (N_13678,N_5236,N_6749);
nor U13679 (N_13679,N_9848,N_7025);
xnor U13680 (N_13680,N_5305,N_7891);
and U13681 (N_13681,N_8274,N_8837);
and U13682 (N_13682,N_7169,N_6311);
and U13683 (N_13683,N_6651,N_9106);
and U13684 (N_13684,N_8050,N_8341);
nor U13685 (N_13685,N_9893,N_7163);
nand U13686 (N_13686,N_6991,N_6660);
or U13687 (N_13687,N_9007,N_6236);
xnor U13688 (N_13688,N_8622,N_5896);
nor U13689 (N_13689,N_6449,N_5401);
nor U13690 (N_13690,N_7668,N_5120);
nand U13691 (N_13691,N_5687,N_7279);
nand U13692 (N_13692,N_8057,N_6170);
nor U13693 (N_13693,N_7992,N_7332);
nand U13694 (N_13694,N_5317,N_7204);
xor U13695 (N_13695,N_9925,N_9021);
nand U13696 (N_13696,N_9805,N_5844);
or U13697 (N_13697,N_6301,N_5626);
nor U13698 (N_13698,N_8420,N_9977);
or U13699 (N_13699,N_7886,N_8345);
or U13700 (N_13700,N_9562,N_6247);
and U13701 (N_13701,N_5303,N_8632);
and U13702 (N_13702,N_9357,N_9355);
xnor U13703 (N_13703,N_9019,N_7308);
nand U13704 (N_13704,N_6579,N_9046);
nor U13705 (N_13705,N_8317,N_5068);
or U13706 (N_13706,N_7554,N_7294);
nor U13707 (N_13707,N_6776,N_7597);
and U13708 (N_13708,N_5146,N_6184);
nand U13709 (N_13709,N_9261,N_5778);
xor U13710 (N_13710,N_6394,N_9063);
or U13711 (N_13711,N_8012,N_5893);
and U13712 (N_13712,N_6852,N_5516);
xnor U13713 (N_13713,N_9773,N_5348);
and U13714 (N_13714,N_5680,N_7790);
nor U13715 (N_13715,N_6349,N_5512);
xnor U13716 (N_13716,N_5077,N_9375);
nand U13717 (N_13717,N_8313,N_6025);
nand U13718 (N_13718,N_9551,N_6448);
nor U13719 (N_13719,N_5228,N_5825);
nor U13720 (N_13720,N_9579,N_5168);
nand U13721 (N_13721,N_8859,N_7056);
and U13722 (N_13722,N_7421,N_9616);
or U13723 (N_13723,N_9856,N_7077);
nor U13724 (N_13724,N_9434,N_8034);
or U13725 (N_13725,N_6331,N_9248);
nand U13726 (N_13726,N_6770,N_8948);
and U13727 (N_13727,N_8228,N_9940);
nand U13728 (N_13728,N_9485,N_9971);
nand U13729 (N_13729,N_6020,N_6395);
nand U13730 (N_13730,N_7874,N_9895);
nor U13731 (N_13731,N_6142,N_6538);
and U13732 (N_13732,N_9674,N_5606);
xor U13733 (N_13733,N_6041,N_7305);
or U13734 (N_13734,N_7219,N_9966);
or U13735 (N_13735,N_6450,N_9758);
and U13736 (N_13736,N_6557,N_8193);
or U13737 (N_13737,N_5231,N_8567);
nor U13738 (N_13738,N_9306,N_5990);
xor U13739 (N_13739,N_9439,N_7776);
or U13740 (N_13740,N_8152,N_7376);
nor U13741 (N_13741,N_9786,N_7454);
nand U13742 (N_13742,N_9277,N_8544);
nand U13743 (N_13743,N_5237,N_6639);
and U13744 (N_13744,N_9053,N_9057);
xnor U13745 (N_13745,N_8234,N_5933);
nand U13746 (N_13746,N_8114,N_9497);
or U13747 (N_13747,N_7982,N_9081);
nand U13748 (N_13748,N_6753,N_5246);
and U13749 (N_13749,N_8153,N_9678);
and U13750 (N_13750,N_6111,N_9313);
and U13751 (N_13751,N_7945,N_8336);
nor U13752 (N_13752,N_5373,N_6289);
xnor U13753 (N_13753,N_6716,N_9583);
nor U13754 (N_13754,N_5474,N_5301);
and U13755 (N_13755,N_6178,N_7852);
and U13756 (N_13756,N_7647,N_8843);
xor U13757 (N_13757,N_8650,N_5903);
nand U13758 (N_13758,N_7508,N_8899);
nor U13759 (N_13759,N_7927,N_5269);
nand U13760 (N_13760,N_8117,N_9707);
nor U13761 (N_13761,N_9054,N_7697);
nand U13762 (N_13762,N_9718,N_8178);
xor U13763 (N_13763,N_8731,N_7295);
nand U13764 (N_13764,N_7529,N_8468);
or U13765 (N_13765,N_5064,N_9184);
nand U13766 (N_13766,N_7646,N_8548);
and U13767 (N_13767,N_6134,N_5507);
nand U13768 (N_13768,N_7291,N_7106);
and U13769 (N_13769,N_7020,N_5480);
or U13770 (N_13770,N_8597,N_8611);
and U13771 (N_13771,N_7652,N_9173);
nor U13772 (N_13772,N_9078,N_8259);
and U13773 (N_13773,N_6914,N_8226);
xor U13774 (N_13774,N_7205,N_8129);
nor U13775 (N_13775,N_7419,N_7194);
nor U13776 (N_13776,N_6059,N_8443);
and U13777 (N_13777,N_5298,N_5260);
nor U13778 (N_13778,N_9505,N_7603);
xor U13779 (N_13779,N_7535,N_6940);
nor U13780 (N_13780,N_7558,N_5200);
or U13781 (N_13781,N_9425,N_5186);
nor U13782 (N_13782,N_8339,N_7300);
xor U13783 (N_13783,N_5800,N_8904);
or U13784 (N_13784,N_9317,N_5766);
nor U13785 (N_13785,N_7804,N_7816);
or U13786 (N_13786,N_5619,N_6507);
or U13787 (N_13787,N_5029,N_5124);
or U13788 (N_13788,N_7889,N_9271);
and U13789 (N_13789,N_6483,N_5321);
nand U13790 (N_13790,N_8779,N_5244);
or U13791 (N_13791,N_8338,N_7110);
nor U13792 (N_13792,N_7314,N_5046);
nor U13793 (N_13793,N_5029,N_5194);
or U13794 (N_13794,N_6380,N_8042);
xnor U13795 (N_13795,N_5053,N_8128);
nor U13796 (N_13796,N_9097,N_6694);
and U13797 (N_13797,N_7547,N_6064);
and U13798 (N_13798,N_8563,N_9042);
and U13799 (N_13799,N_6474,N_7545);
nand U13800 (N_13800,N_8986,N_5685);
xor U13801 (N_13801,N_9688,N_5876);
nand U13802 (N_13802,N_5054,N_6929);
or U13803 (N_13803,N_9176,N_6882);
or U13804 (N_13804,N_9135,N_6434);
xnor U13805 (N_13805,N_8053,N_5032);
nor U13806 (N_13806,N_5056,N_8004);
nand U13807 (N_13807,N_6448,N_6743);
xor U13808 (N_13808,N_9774,N_5060);
and U13809 (N_13809,N_8133,N_6201);
or U13810 (N_13810,N_7765,N_8117);
and U13811 (N_13811,N_8767,N_6070);
or U13812 (N_13812,N_5536,N_5676);
nor U13813 (N_13813,N_9003,N_5949);
xnor U13814 (N_13814,N_6071,N_8612);
and U13815 (N_13815,N_6910,N_7975);
and U13816 (N_13816,N_7300,N_9383);
nor U13817 (N_13817,N_9535,N_9284);
and U13818 (N_13818,N_6600,N_9158);
nand U13819 (N_13819,N_6572,N_6415);
nand U13820 (N_13820,N_9011,N_8985);
or U13821 (N_13821,N_8023,N_5575);
and U13822 (N_13822,N_8593,N_8869);
nand U13823 (N_13823,N_6868,N_6175);
nand U13824 (N_13824,N_7700,N_7200);
nand U13825 (N_13825,N_8732,N_8986);
or U13826 (N_13826,N_9680,N_6178);
nor U13827 (N_13827,N_8105,N_9937);
or U13828 (N_13828,N_6292,N_9931);
nor U13829 (N_13829,N_7068,N_5502);
and U13830 (N_13830,N_9023,N_9379);
or U13831 (N_13831,N_6898,N_5313);
nand U13832 (N_13832,N_6096,N_8299);
nand U13833 (N_13833,N_6217,N_6408);
nand U13834 (N_13834,N_9907,N_9386);
or U13835 (N_13835,N_9433,N_7598);
nor U13836 (N_13836,N_7577,N_6055);
nor U13837 (N_13837,N_6996,N_6932);
nand U13838 (N_13838,N_8350,N_8832);
xnor U13839 (N_13839,N_7088,N_9876);
nand U13840 (N_13840,N_9342,N_7804);
and U13841 (N_13841,N_7449,N_5640);
or U13842 (N_13842,N_7372,N_5854);
nor U13843 (N_13843,N_5567,N_6131);
or U13844 (N_13844,N_6010,N_5490);
and U13845 (N_13845,N_7730,N_5192);
or U13846 (N_13846,N_5685,N_7962);
nor U13847 (N_13847,N_7425,N_7692);
nor U13848 (N_13848,N_7290,N_7708);
or U13849 (N_13849,N_6153,N_9314);
xnor U13850 (N_13850,N_6310,N_9235);
or U13851 (N_13851,N_7988,N_5862);
nor U13852 (N_13852,N_8676,N_8096);
nor U13853 (N_13853,N_7381,N_5053);
xnor U13854 (N_13854,N_7634,N_6930);
xor U13855 (N_13855,N_6380,N_8870);
xnor U13856 (N_13856,N_8572,N_8355);
or U13857 (N_13857,N_5908,N_7497);
or U13858 (N_13858,N_8701,N_6264);
and U13859 (N_13859,N_5736,N_5812);
nand U13860 (N_13860,N_6248,N_5106);
and U13861 (N_13861,N_7345,N_8041);
and U13862 (N_13862,N_8606,N_8819);
xor U13863 (N_13863,N_6418,N_9691);
and U13864 (N_13864,N_6232,N_7140);
xor U13865 (N_13865,N_9261,N_6813);
or U13866 (N_13866,N_8940,N_8038);
and U13867 (N_13867,N_7470,N_6647);
and U13868 (N_13868,N_7602,N_8919);
and U13869 (N_13869,N_6206,N_5536);
nor U13870 (N_13870,N_7025,N_5780);
or U13871 (N_13871,N_5297,N_6901);
nand U13872 (N_13872,N_7823,N_5081);
or U13873 (N_13873,N_9111,N_5872);
and U13874 (N_13874,N_8861,N_8183);
and U13875 (N_13875,N_8940,N_9684);
and U13876 (N_13876,N_6699,N_8040);
nand U13877 (N_13877,N_7524,N_6587);
xor U13878 (N_13878,N_5749,N_6313);
xor U13879 (N_13879,N_7650,N_5591);
or U13880 (N_13880,N_5769,N_6697);
nor U13881 (N_13881,N_6566,N_9990);
and U13882 (N_13882,N_5757,N_6907);
xor U13883 (N_13883,N_5555,N_5353);
and U13884 (N_13884,N_6609,N_8457);
and U13885 (N_13885,N_6475,N_8699);
or U13886 (N_13886,N_6937,N_5970);
and U13887 (N_13887,N_6469,N_6613);
xor U13888 (N_13888,N_8197,N_8928);
and U13889 (N_13889,N_5736,N_6094);
xnor U13890 (N_13890,N_6200,N_6880);
nor U13891 (N_13891,N_6930,N_5761);
nand U13892 (N_13892,N_7455,N_5101);
nor U13893 (N_13893,N_5613,N_9860);
and U13894 (N_13894,N_5700,N_6799);
or U13895 (N_13895,N_5307,N_8907);
or U13896 (N_13896,N_9877,N_9557);
xor U13897 (N_13897,N_8013,N_9327);
nand U13898 (N_13898,N_5880,N_9679);
xor U13899 (N_13899,N_5299,N_9231);
and U13900 (N_13900,N_5044,N_6283);
and U13901 (N_13901,N_7991,N_5645);
xnor U13902 (N_13902,N_5391,N_8791);
nand U13903 (N_13903,N_7013,N_7515);
and U13904 (N_13904,N_5326,N_7054);
and U13905 (N_13905,N_6588,N_9013);
nand U13906 (N_13906,N_9325,N_7172);
and U13907 (N_13907,N_9193,N_8551);
xor U13908 (N_13908,N_6228,N_9858);
or U13909 (N_13909,N_6261,N_6054);
nor U13910 (N_13910,N_7586,N_8186);
nor U13911 (N_13911,N_6476,N_5183);
xnor U13912 (N_13912,N_8545,N_8159);
xor U13913 (N_13913,N_8538,N_8940);
and U13914 (N_13914,N_6970,N_8165);
nand U13915 (N_13915,N_7716,N_8202);
nor U13916 (N_13916,N_9124,N_7875);
nand U13917 (N_13917,N_5003,N_7166);
and U13918 (N_13918,N_5167,N_5123);
nor U13919 (N_13919,N_8473,N_8895);
xnor U13920 (N_13920,N_8270,N_9161);
nand U13921 (N_13921,N_7382,N_7746);
and U13922 (N_13922,N_9704,N_9030);
nor U13923 (N_13923,N_7927,N_7322);
nor U13924 (N_13924,N_5161,N_7869);
and U13925 (N_13925,N_8190,N_5748);
xor U13926 (N_13926,N_7967,N_9728);
nand U13927 (N_13927,N_9998,N_7950);
and U13928 (N_13928,N_5526,N_8250);
and U13929 (N_13929,N_6243,N_5320);
or U13930 (N_13930,N_7299,N_9330);
nor U13931 (N_13931,N_5440,N_9434);
and U13932 (N_13932,N_7808,N_9888);
xnor U13933 (N_13933,N_6293,N_6808);
and U13934 (N_13934,N_5689,N_6270);
nor U13935 (N_13935,N_9520,N_6526);
xor U13936 (N_13936,N_8225,N_8266);
or U13937 (N_13937,N_8499,N_9425);
or U13938 (N_13938,N_7285,N_6496);
xnor U13939 (N_13939,N_8537,N_8636);
and U13940 (N_13940,N_8888,N_6639);
and U13941 (N_13941,N_8649,N_5049);
or U13942 (N_13942,N_7548,N_9147);
xnor U13943 (N_13943,N_6555,N_7530);
xnor U13944 (N_13944,N_9616,N_6895);
nor U13945 (N_13945,N_5128,N_7919);
or U13946 (N_13946,N_5208,N_5839);
nor U13947 (N_13947,N_7527,N_5227);
and U13948 (N_13948,N_6342,N_5966);
and U13949 (N_13949,N_9036,N_5086);
nor U13950 (N_13950,N_9388,N_6574);
nor U13951 (N_13951,N_5657,N_8223);
nand U13952 (N_13952,N_5140,N_6891);
xor U13953 (N_13953,N_9436,N_5494);
xor U13954 (N_13954,N_8328,N_8780);
nor U13955 (N_13955,N_7580,N_6932);
nand U13956 (N_13956,N_7972,N_9462);
or U13957 (N_13957,N_8521,N_7207);
or U13958 (N_13958,N_6147,N_5971);
or U13959 (N_13959,N_8941,N_9545);
nand U13960 (N_13960,N_6245,N_8104);
xnor U13961 (N_13961,N_6061,N_6322);
xnor U13962 (N_13962,N_7657,N_9403);
xnor U13963 (N_13963,N_8467,N_7736);
nand U13964 (N_13964,N_8758,N_8849);
xor U13965 (N_13965,N_9785,N_7237);
and U13966 (N_13966,N_5911,N_7272);
xnor U13967 (N_13967,N_8770,N_6607);
and U13968 (N_13968,N_9608,N_7973);
xnor U13969 (N_13969,N_8990,N_8286);
and U13970 (N_13970,N_9527,N_7323);
or U13971 (N_13971,N_6909,N_7742);
nor U13972 (N_13972,N_7513,N_8456);
nand U13973 (N_13973,N_7156,N_6657);
nand U13974 (N_13974,N_5060,N_9326);
nor U13975 (N_13975,N_6232,N_5647);
nand U13976 (N_13976,N_7897,N_9287);
and U13977 (N_13977,N_6884,N_8815);
xor U13978 (N_13978,N_6816,N_5165);
or U13979 (N_13979,N_7022,N_5266);
xor U13980 (N_13980,N_9882,N_6816);
or U13981 (N_13981,N_5666,N_6412);
or U13982 (N_13982,N_7894,N_9686);
nand U13983 (N_13983,N_6296,N_9590);
nand U13984 (N_13984,N_5438,N_9498);
nor U13985 (N_13985,N_9705,N_6645);
or U13986 (N_13986,N_9143,N_8783);
xor U13987 (N_13987,N_8368,N_5782);
nand U13988 (N_13988,N_7087,N_8401);
and U13989 (N_13989,N_9461,N_9896);
xnor U13990 (N_13990,N_5738,N_9680);
nor U13991 (N_13991,N_9863,N_8528);
and U13992 (N_13992,N_6991,N_9579);
or U13993 (N_13993,N_7776,N_8342);
and U13994 (N_13994,N_7595,N_9236);
or U13995 (N_13995,N_8819,N_8799);
and U13996 (N_13996,N_6497,N_5664);
nand U13997 (N_13997,N_6309,N_7683);
and U13998 (N_13998,N_9087,N_9987);
and U13999 (N_13999,N_6801,N_5579);
xor U14000 (N_14000,N_8973,N_7590);
xor U14001 (N_14001,N_8284,N_7034);
and U14002 (N_14002,N_6997,N_8087);
or U14003 (N_14003,N_5993,N_8109);
or U14004 (N_14004,N_5956,N_9833);
nand U14005 (N_14005,N_8424,N_8505);
or U14006 (N_14006,N_5940,N_5428);
or U14007 (N_14007,N_6453,N_9999);
or U14008 (N_14008,N_5502,N_6581);
and U14009 (N_14009,N_7941,N_5247);
nand U14010 (N_14010,N_6961,N_6225);
xnor U14011 (N_14011,N_5175,N_6251);
nand U14012 (N_14012,N_7715,N_9360);
nor U14013 (N_14013,N_7489,N_6091);
xnor U14014 (N_14014,N_7148,N_6811);
or U14015 (N_14015,N_5281,N_6639);
xnor U14016 (N_14016,N_8531,N_5122);
xor U14017 (N_14017,N_6903,N_6005);
nor U14018 (N_14018,N_8470,N_9944);
nor U14019 (N_14019,N_9312,N_8833);
or U14020 (N_14020,N_7506,N_6204);
nand U14021 (N_14021,N_7929,N_7023);
nand U14022 (N_14022,N_8835,N_7191);
nand U14023 (N_14023,N_9728,N_7004);
xnor U14024 (N_14024,N_6696,N_9696);
and U14025 (N_14025,N_7044,N_9401);
or U14026 (N_14026,N_6060,N_7475);
nor U14027 (N_14027,N_6525,N_7806);
xnor U14028 (N_14028,N_7230,N_7432);
or U14029 (N_14029,N_6590,N_5392);
nor U14030 (N_14030,N_6637,N_6285);
xor U14031 (N_14031,N_5011,N_8136);
xor U14032 (N_14032,N_7897,N_8280);
nor U14033 (N_14033,N_6996,N_9869);
xnor U14034 (N_14034,N_8766,N_9876);
or U14035 (N_14035,N_9901,N_9194);
nor U14036 (N_14036,N_5052,N_5307);
nand U14037 (N_14037,N_8204,N_5935);
nand U14038 (N_14038,N_7635,N_8016);
nor U14039 (N_14039,N_8302,N_7363);
and U14040 (N_14040,N_5868,N_5980);
nor U14041 (N_14041,N_6822,N_6747);
nand U14042 (N_14042,N_9750,N_7055);
or U14043 (N_14043,N_8349,N_8341);
and U14044 (N_14044,N_5996,N_5191);
xor U14045 (N_14045,N_6251,N_8331);
nor U14046 (N_14046,N_6257,N_5622);
nand U14047 (N_14047,N_8251,N_6311);
nand U14048 (N_14048,N_8446,N_7044);
nand U14049 (N_14049,N_6980,N_8431);
or U14050 (N_14050,N_7049,N_6776);
nor U14051 (N_14051,N_8008,N_5491);
nand U14052 (N_14052,N_7397,N_9737);
nor U14053 (N_14053,N_9371,N_7664);
and U14054 (N_14054,N_6472,N_9549);
nand U14055 (N_14055,N_7782,N_6531);
xnor U14056 (N_14056,N_8578,N_9096);
or U14057 (N_14057,N_7983,N_7845);
nand U14058 (N_14058,N_6354,N_9532);
xnor U14059 (N_14059,N_8207,N_6049);
nand U14060 (N_14060,N_6989,N_6019);
and U14061 (N_14061,N_8470,N_7736);
or U14062 (N_14062,N_9738,N_5058);
and U14063 (N_14063,N_7173,N_7356);
or U14064 (N_14064,N_5085,N_7869);
nand U14065 (N_14065,N_7536,N_7984);
and U14066 (N_14066,N_5978,N_6413);
or U14067 (N_14067,N_9470,N_6995);
nand U14068 (N_14068,N_5273,N_5652);
and U14069 (N_14069,N_7701,N_5123);
xnor U14070 (N_14070,N_9240,N_9250);
xnor U14071 (N_14071,N_7908,N_6351);
and U14072 (N_14072,N_8676,N_6190);
and U14073 (N_14073,N_9338,N_9234);
nor U14074 (N_14074,N_8534,N_9184);
nor U14075 (N_14075,N_5267,N_7249);
nor U14076 (N_14076,N_7239,N_9247);
nand U14077 (N_14077,N_7088,N_7232);
or U14078 (N_14078,N_8405,N_5491);
nor U14079 (N_14079,N_5239,N_5669);
and U14080 (N_14080,N_6369,N_7349);
xor U14081 (N_14081,N_8578,N_5145);
and U14082 (N_14082,N_9857,N_9203);
nand U14083 (N_14083,N_5422,N_5595);
xor U14084 (N_14084,N_9165,N_8052);
and U14085 (N_14085,N_7639,N_7947);
or U14086 (N_14086,N_9057,N_8095);
or U14087 (N_14087,N_8060,N_5308);
or U14088 (N_14088,N_5982,N_8647);
and U14089 (N_14089,N_9509,N_6577);
xor U14090 (N_14090,N_5761,N_5927);
xnor U14091 (N_14091,N_8996,N_7758);
and U14092 (N_14092,N_9372,N_8239);
xnor U14093 (N_14093,N_9988,N_8233);
and U14094 (N_14094,N_5044,N_7555);
nor U14095 (N_14095,N_6101,N_8343);
and U14096 (N_14096,N_9346,N_7289);
or U14097 (N_14097,N_9324,N_6804);
or U14098 (N_14098,N_8677,N_8088);
nand U14099 (N_14099,N_9326,N_8079);
nand U14100 (N_14100,N_5956,N_7042);
nand U14101 (N_14101,N_7822,N_5079);
nor U14102 (N_14102,N_6286,N_6420);
and U14103 (N_14103,N_5068,N_7205);
nor U14104 (N_14104,N_9873,N_9963);
nor U14105 (N_14105,N_5240,N_9777);
or U14106 (N_14106,N_5034,N_7698);
and U14107 (N_14107,N_7578,N_9616);
and U14108 (N_14108,N_8219,N_8342);
nand U14109 (N_14109,N_8193,N_9726);
nor U14110 (N_14110,N_8436,N_9548);
xor U14111 (N_14111,N_5935,N_5270);
nand U14112 (N_14112,N_9286,N_6017);
or U14113 (N_14113,N_8680,N_5774);
nor U14114 (N_14114,N_7814,N_7405);
nor U14115 (N_14115,N_8233,N_9085);
xnor U14116 (N_14116,N_7258,N_5800);
nor U14117 (N_14117,N_7973,N_7125);
nand U14118 (N_14118,N_7325,N_5332);
xnor U14119 (N_14119,N_5563,N_9925);
and U14120 (N_14120,N_6973,N_7134);
xnor U14121 (N_14121,N_5479,N_7459);
or U14122 (N_14122,N_5549,N_8726);
nor U14123 (N_14123,N_5565,N_8900);
xor U14124 (N_14124,N_9753,N_7939);
and U14125 (N_14125,N_6270,N_6840);
xor U14126 (N_14126,N_7544,N_6983);
and U14127 (N_14127,N_6446,N_5212);
or U14128 (N_14128,N_8814,N_5313);
or U14129 (N_14129,N_7458,N_7514);
nand U14130 (N_14130,N_5226,N_8230);
xor U14131 (N_14131,N_9212,N_7306);
or U14132 (N_14132,N_7363,N_6120);
and U14133 (N_14133,N_5199,N_9642);
nand U14134 (N_14134,N_8115,N_7912);
xor U14135 (N_14135,N_9529,N_7670);
xor U14136 (N_14136,N_6339,N_6737);
nand U14137 (N_14137,N_5449,N_7151);
nand U14138 (N_14138,N_5926,N_8190);
or U14139 (N_14139,N_8700,N_5482);
and U14140 (N_14140,N_7452,N_8554);
nor U14141 (N_14141,N_7190,N_7626);
xnor U14142 (N_14142,N_5483,N_7366);
or U14143 (N_14143,N_8306,N_6336);
nand U14144 (N_14144,N_7931,N_8262);
and U14145 (N_14145,N_5237,N_8056);
xnor U14146 (N_14146,N_7396,N_7022);
nand U14147 (N_14147,N_8945,N_8427);
xor U14148 (N_14148,N_5261,N_8963);
or U14149 (N_14149,N_5722,N_8898);
and U14150 (N_14150,N_5878,N_9149);
xnor U14151 (N_14151,N_7473,N_5555);
xor U14152 (N_14152,N_8324,N_8210);
nor U14153 (N_14153,N_8124,N_9462);
nand U14154 (N_14154,N_7454,N_9103);
or U14155 (N_14155,N_5804,N_7460);
nor U14156 (N_14156,N_8373,N_9940);
and U14157 (N_14157,N_7371,N_8059);
xor U14158 (N_14158,N_5067,N_9724);
and U14159 (N_14159,N_9999,N_6254);
xor U14160 (N_14160,N_9311,N_5984);
or U14161 (N_14161,N_6163,N_5936);
nor U14162 (N_14162,N_5089,N_8643);
xor U14163 (N_14163,N_9154,N_9072);
xnor U14164 (N_14164,N_5327,N_6515);
xnor U14165 (N_14165,N_9021,N_7136);
nand U14166 (N_14166,N_6712,N_8267);
or U14167 (N_14167,N_6683,N_5084);
nand U14168 (N_14168,N_6844,N_8606);
or U14169 (N_14169,N_8806,N_9720);
nor U14170 (N_14170,N_8459,N_7197);
nand U14171 (N_14171,N_7571,N_5945);
or U14172 (N_14172,N_7104,N_9567);
nand U14173 (N_14173,N_5714,N_7728);
nand U14174 (N_14174,N_8175,N_7835);
nor U14175 (N_14175,N_8972,N_9027);
or U14176 (N_14176,N_7305,N_5894);
or U14177 (N_14177,N_8614,N_7866);
nor U14178 (N_14178,N_7743,N_6646);
and U14179 (N_14179,N_8489,N_9768);
and U14180 (N_14180,N_7597,N_9125);
xnor U14181 (N_14181,N_8749,N_6605);
or U14182 (N_14182,N_7078,N_6673);
and U14183 (N_14183,N_6986,N_5601);
nand U14184 (N_14184,N_5202,N_8885);
or U14185 (N_14185,N_6600,N_8843);
and U14186 (N_14186,N_5419,N_5925);
nor U14187 (N_14187,N_7966,N_5419);
xor U14188 (N_14188,N_8528,N_8402);
and U14189 (N_14189,N_5022,N_5161);
and U14190 (N_14190,N_5866,N_8143);
or U14191 (N_14191,N_6747,N_9265);
xnor U14192 (N_14192,N_6783,N_6754);
or U14193 (N_14193,N_7761,N_8329);
and U14194 (N_14194,N_8531,N_5422);
or U14195 (N_14195,N_6196,N_5694);
nor U14196 (N_14196,N_6452,N_6744);
nand U14197 (N_14197,N_9217,N_7018);
nor U14198 (N_14198,N_8498,N_7000);
and U14199 (N_14199,N_8707,N_6312);
nand U14200 (N_14200,N_9959,N_8833);
xor U14201 (N_14201,N_5567,N_8205);
nor U14202 (N_14202,N_7769,N_9275);
or U14203 (N_14203,N_6066,N_8880);
and U14204 (N_14204,N_6977,N_5164);
and U14205 (N_14205,N_5209,N_6593);
or U14206 (N_14206,N_7545,N_9457);
nand U14207 (N_14207,N_8942,N_5321);
or U14208 (N_14208,N_6638,N_6197);
and U14209 (N_14209,N_6184,N_6067);
or U14210 (N_14210,N_7302,N_5769);
nand U14211 (N_14211,N_9747,N_5261);
xor U14212 (N_14212,N_8538,N_5500);
xor U14213 (N_14213,N_9861,N_9394);
and U14214 (N_14214,N_7336,N_6699);
nor U14215 (N_14215,N_7595,N_5585);
and U14216 (N_14216,N_5866,N_7516);
and U14217 (N_14217,N_9295,N_5768);
nor U14218 (N_14218,N_8235,N_7104);
and U14219 (N_14219,N_5839,N_6974);
or U14220 (N_14220,N_5204,N_8698);
nand U14221 (N_14221,N_5520,N_5227);
or U14222 (N_14222,N_8683,N_8188);
and U14223 (N_14223,N_9640,N_7713);
nor U14224 (N_14224,N_5886,N_9095);
and U14225 (N_14225,N_7017,N_7684);
or U14226 (N_14226,N_9310,N_7227);
and U14227 (N_14227,N_8313,N_7215);
or U14228 (N_14228,N_9937,N_6920);
xor U14229 (N_14229,N_6945,N_5967);
and U14230 (N_14230,N_9654,N_8960);
nand U14231 (N_14231,N_5579,N_8913);
or U14232 (N_14232,N_7593,N_7383);
xor U14233 (N_14233,N_8476,N_6406);
nor U14234 (N_14234,N_6667,N_6625);
or U14235 (N_14235,N_7689,N_5603);
nand U14236 (N_14236,N_9673,N_5316);
or U14237 (N_14237,N_6241,N_9291);
nor U14238 (N_14238,N_8970,N_8815);
and U14239 (N_14239,N_7061,N_5085);
nor U14240 (N_14240,N_6607,N_7087);
xnor U14241 (N_14241,N_6182,N_9093);
or U14242 (N_14242,N_9795,N_9770);
or U14243 (N_14243,N_5757,N_6146);
or U14244 (N_14244,N_6564,N_9277);
or U14245 (N_14245,N_7493,N_5000);
xnor U14246 (N_14246,N_5552,N_8040);
nand U14247 (N_14247,N_8155,N_8305);
nand U14248 (N_14248,N_9507,N_8012);
and U14249 (N_14249,N_5559,N_6256);
and U14250 (N_14250,N_6225,N_9605);
xnor U14251 (N_14251,N_8376,N_9042);
or U14252 (N_14252,N_9110,N_6768);
xor U14253 (N_14253,N_9256,N_9105);
nor U14254 (N_14254,N_9401,N_7692);
or U14255 (N_14255,N_5094,N_6336);
nand U14256 (N_14256,N_6712,N_9607);
nand U14257 (N_14257,N_8154,N_8800);
xnor U14258 (N_14258,N_9824,N_7476);
nand U14259 (N_14259,N_7026,N_8334);
nand U14260 (N_14260,N_8471,N_6747);
nand U14261 (N_14261,N_7754,N_7953);
or U14262 (N_14262,N_5224,N_8154);
and U14263 (N_14263,N_6723,N_7876);
nand U14264 (N_14264,N_6729,N_9772);
xnor U14265 (N_14265,N_9173,N_6278);
nand U14266 (N_14266,N_8507,N_7593);
nand U14267 (N_14267,N_5149,N_8563);
nor U14268 (N_14268,N_7285,N_7303);
nor U14269 (N_14269,N_6005,N_5188);
or U14270 (N_14270,N_8773,N_7662);
and U14271 (N_14271,N_8885,N_7799);
and U14272 (N_14272,N_5157,N_8902);
nand U14273 (N_14273,N_7933,N_7257);
xnor U14274 (N_14274,N_9924,N_6073);
nor U14275 (N_14275,N_6317,N_5569);
xor U14276 (N_14276,N_5371,N_8786);
and U14277 (N_14277,N_7024,N_8524);
or U14278 (N_14278,N_7491,N_7314);
or U14279 (N_14279,N_6834,N_9121);
and U14280 (N_14280,N_9858,N_9735);
nand U14281 (N_14281,N_9257,N_8363);
nor U14282 (N_14282,N_9369,N_8131);
xnor U14283 (N_14283,N_5822,N_8459);
nor U14284 (N_14284,N_7958,N_6280);
nor U14285 (N_14285,N_8518,N_6850);
nor U14286 (N_14286,N_7589,N_7203);
nand U14287 (N_14287,N_6012,N_5465);
nand U14288 (N_14288,N_9327,N_9168);
and U14289 (N_14289,N_8094,N_9647);
nor U14290 (N_14290,N_7231,N_5866);
xor U14291 (N_14291,N_6124,N_9484);
or U14292 (N_14292,N_9421,N_6514);
nand U14293 (N_14293,N_5882,N_9296);
nor U14294 (N_14294,N_7571,N_8329);
xor U14295 (N_14295,N_8176,N_7763);
xor U14296 (N_14296,N_8751,N_5365);
nor U14297 (N_14297,N_6563,N_9694);
or U14298 (N_14298,N_6885,N_8827);
and U14299 (N_14299,N_7363,N_8819);
nor U14300 (N_14300,N_5201,N_7364);
xnor U14301 (N_14301,N_7982,N_6509);
nand U14302 (N_14302,N_9068,N_8460);
nor U14303 (N_14303,N_7959,N_8849);
nor U14304 (N_14304,N_6075,N_6956);
nand U14305 (N_14305,N_7537,N_8227);
nand U14306 (N_14306,N_8888,N_5626);
nor U14307 (N_14307,N_8813,N_6575);
xor U14308 (N_14308,N_7007,N_9990);
or U14309 (N_14309,N_6319,N_9490);
or U14310 (N_14310,N_6661,N_5263);
nand U14311 (N_14311,N_6583,N_9419);
xnor U14312 (N_14312,N_5710,N_9014);
xor U14313 (N_14313,N_9197,N_7213);
or U14314 (N_14314,N_7053,N_7433);
and U14315 (N_14315,N_8909,N_8996);
xnor U14316 (N_14316,N_7216,N_5447);
nor U14317 (N_14317,N_9588,N_9048);
nand U14318 (N_14318,N_7179,N_9254);
xnor U14319 (N_14319,N_9002,N_8525);
and U14320 (N_14320,N_8143,N_7246);
and U14321 (N_14321,N_6086,N_6913);
nand U14322 (N_14322,N_8793,N_7714);
nor U14323 (N_14323,N_6097,N_5201);
and U14324 (N_14324,N_9350,N_5570);
nand U14325 (N_14325,N_8282,N_9295);
nor U14326 (N_14326,N_9843,N_9510);
nor U14327 (N_14327,N_9935,N_9113);
nor U14328 (N_14328,N_8619,N_5230);
xnor U14329 (N_14329,N_9574,N_6478);
nand U14330 (N_14330,N_8981,N_7922);
xor U14331 (N_14331,N_6671,N_5066);
xor U14332 (N_14332,N_8490,N_6987);
nor U14333 (N_14333,N_6384,N_5474);
and U14334 (N_14334,N_8372,N_8989);
nor U14335 (N_14335,N_7964,N_6304);
nor U14336 (N_14336,N_5120,N_5062);
xor U14337 (N_14337,N_6495,N_9744);
nand U14338 (N_14338,N_5138,N_8002);
nand U14339 (N_14339,N_5116,N_9875);
nand U14340 (N_14340,N_7288,N_7473);
and U14341 (N_14341,N_9331,N_5377);
and U14342 (N_14342,N_7416,N_7368);
nand U14343 (N_14343,N_7304,N_9692);
nor U14344 (N_14344,N_5010,N_7486);
xor U14345 (N_14345,N_7553,N_7292);
xor U14346 (N_14346,N_8713,N_5239);
nor U14347 (N_14347,N_9413,N_6887);
nor U14348 (N_14348,N_8635,N_9293);
nor U14349 (N_14349,N_7000,N_6512);
xor U14350 (N_14350,N_8120,N_5854);
and U14351 (N_14351,N_7761,N_6086);
xor U14352 (N_14352,N_7969,N_7015);
and U14353 (N_14353,N_5297,N_8561);
xor U14354 (N_14354,N_9310,N_6896);
xor U14355 (N_14355,N_6181,N_5331);
xnor U14356 (N_14356,N_6865,N_5420);
or U14357 (N_14357,N_8355,N_5124);
xnor U14358 (N_14358,N_8156,N_6850);
or U14359 (N_14359,N_7081,N_9240);
and U14360 (N_14360,N_9040,N_5516);
and U14361 (N_14361,N_8730,N_9093);
or U14362 (N_14362,N_8380,N_8776);
and U14363 (N_14363,N_9639,N_6283);
nor U14364 (N_14364,N_5684,N_8044);
or U14365 (N_14365,N_6343,N_5457);
and U14366 (N_14366,N_9584,N_5241);
or U14367 (N_14367,N_9580,N_6980);
and U14368 (N_14368,N_9184,N_8570);
nand U14369 (N_14369,N_8755,N_5805);
nor U14370 (N_14370,N_9977,N_6436);
nor U14371 (N_14371,N_9222,N_8685);
nand U14372 (N_14372,N_8102,N_6497);
xnor U14373 (N_14373,N_7593,N_8997);
xor U14374 (N_14374,N_6387,N_6784);
nor U14375 (N_14375,N_7220,N_8788);
or U14376 (N_14376,N_6941,N_5922);
and U14377 (N_14377,N_7181,N_7911);
or U14378 (N_14378,N_7650,N_7252);
xor U14379 (N_14379,N_8160,N_7066);
or U14380 (N_14380,N_6703,N_7901);
nor U14381 (N_14381,N_9275,N_6024);
nor U14382 (N_14382,N_9019,N_7529);
nor U14383 (N_14383,N_6744,N_8886);
xor U14384 (N_14384,N_7965,N_9456);
xor U14385 (N_14385,N_6544,N_6215);
nand U14386 (N_14386,N_7121,N_8857);
xor U14387 (N_14387,N_5056,N_6623);
nand U14388 (N_14388,N_8505,N_8995);
nand U14389 (N_14389,N_9266,N_7497);
and U14390 (N_14390,N_9424,N_8632);
nor U14391 (N_14391,N_5454,N_9045);
and U14392 (N_14392,N_6377,N_5318);
or U14393 (N_14393,N_7662,N_9108);
nand U14394 (N_14394,N_9435,N_7416);
nor U14395 (N_14395,N_8737,N_9692);
nor U14396 (N_14396,N_5859,N_5037);
or U14397 (N_14397,N_7283,N_5215);
and U14398 (N_14398,N_8849,N_6614);
nor U14399 (N_14399,N_8999,N_6878);
nand U14400 (N_14400,N_8576,N_8702);
nor U14401 (N_14401,N_8493,N_9305);
or U14402 (N_14402,N_9919,N_6786);
nor U14403 (N_14403,N_7888,N_8669);
nor U14404 (N_14404,N_5230,N_7588);
nand U14405 (N_14405,N_9621,N_9326);
xor U14406 (N_14406,N_9041,N_9165);
xor U14407 (N_14407,N_8812,N_9512);
xor U14408 (N_14408,N_7178,N_8213);
nand U14409 (N_14409,N_8953,N_7256);
xnor U14410 (N_14410,N_7656,N_5540);
nand U14411 (N_14411,N_8835,N_9949);
and U14412 (N_14412,N_6430,N_9332);
xnor U14413 (N_14413,N_5024,N_7027);
xnor U14414 (N_14414,N_7659,N_6156);
nand U14415 (N_14415,N_7387,N_9082);
or U14416 (N_14416,N_5640,N_7172);
xor U14417 (N_14417,N_6314,N_5994);
nand U14418 (N_14418,N_9768,N_8717);
xor U14419 (N_14419,N_9584,N_6505);
nor U14420 (N_14420,N_9601,N_6879);
and U14421 (N_14421,N_5087,N_6027);
nor U14422 (N_14422,N_6791,N_6199);
or U14423 (N_14423,N_7256,N_7410);
nand U14424 (N_14424,N_7639,N_5337);
nand U14425 (N_14425,N_8314,N_8622);
nand U14426 (N_14426,N_8373,N_6586);
and U14427 (N_14427,N_5114,N_8042);
nand U14428 (N_14428,N_5360,N_7213);
nor U14429 (N_14429,N_8800,N_7991);
nand U14430 (N_14430,N_9276,N_5748);
and U14431 (N_14431,N_6609,N_9716);
xnor U14432 (N_14432,N_8955,N_5007);
or U14433 (N_14433,N_6875,N_7178);
nand U14434 (N_14434,N_7788,N_9647);
or U14435 (N_14435,N_7335,N_7926);
nor U14436 (N_14436,N_5601,N_6008);
or U14437 (N_14437,N_5480,N_7422);
nand U14438 (N_14438,N_5405,N_6784);
nor U14439 (N_14439,N_8333,N_8569);
xor U14440 (N_14440,N_5591,N_6200);
xor U14441 (N_14441,N_9069,N_5805);
and U14442 (N_14442,N_5292,N_5865);
and U14443 (N_14443,N_7359,N_5966);
and U14444 (N_14444,N_5424,N_9554);
or U14445 (N_14445,N_6276,N_5152);
nor U14446 (N_14446,N_8304,N_5460);
or U14447 (N_14447,N_7970,N_9627);
or U14448 (N_14448,N_8361,N_6910);
xor U14449 (N_14449,N_5030,N_6374);
nor U14450 (N_14450,N_8574,N_7771);
and U14451 (N_14451,N_7920,N_9239);
nand U14452 (N_14452,N_5116,N_8800);
nand U14453 (N_14453,N_8314,N_8362);
nor U14454 (N_14454,N_5899,N_9760);
and U14455 (N_14455,N_7783,N_7726);
nand U14456 (N_14456,N_6818,N_5717);
and U14457 (N_14457,N_6045,N_8667);
xnor U14458 (N_14458,N_5038,N_5530);
xor U14459 (N_14459,N_9610,N_8009);
xnor U14460 (N_14460,N_8600,N_5449);
nor U14461 (N_14461,N_8703,N_8424);
nor U14462 (N_14462,N_6702,N_7933);
nand U14463 (N_14463,N_5813,N_5357);
nor U14464 (N_14464,N_9482,N_7407);
nand U14465 (N_14465,N_7125,N_7810);
nor U14466 (N_14466,N_8708,N_6298);
nor U14467 (N_14467,N_9315,N_6588);
and U14468 (N_14468,N_5437,N_9723);
nor U14469 (N_14469,N_8900,N_9941);
nand U14470 (N_14470,N_9450,N_8429);
and U14471 (N_14471,N_6891,N_6204);
or U14472 (N_14472,N_8667,N_5561);
and U14473 (N_14473,N_7320,N_8029);
or U14474 (N_14474,N_7777,N_5136);
or U14475 (N_14475,N_9013,N_9164);
xnor U14476 (N_14476,N_6578,N_9680);
or U14477 (N_14477,N_5592,N_5887);
xnor U14478 (N_14478,N_6397,N_6788);
xnor U14479 (N_14479,N_8258,N_5617);
nand U14480 (N_14480,N_9486,N_8472);
nand U14481 (N_14481,N_5574,N_7582);
nor U14482 (N_14482,N_9185,N_8014);
and U14483 (N_14483,N_6169,N_9368);
nor U14484 (N_14484,N_6652,N_5944);
nand U14485 (N_14485,N_6028,N_9071);
and U14486 (N_14486,N_9372,N_9707);
and U14487 (N_14487,N_7995,N_8079);
nor U14488 (N_14488,N_9696,N_6800);
xor U14489 (N_14489,N_8109,N_8525);
or U14490 (N_14490,N_8447,N_7611);
nor U14491 (N_14491,N_7642,N_9819);
and U14492 (N_14492,N_5063,N_9066);
xnor U14493 (N_14493,N_7269,N_8567);
xnor U14494 (N_14494,N_5083,N_8316);
or U14495 (N_14495,N_9037,N_9267);
nand U14496 (N_14496,N_6940,N_6058);
nand U14497 (N_14497,N_6023,N_7939);
nand U14498 (N_14498,N_7152,N_6859);
nor U14499 (N_14499,N_8348,N_7799);
nand U14500 (N_14500,N_7874,N_7772);
or U14501 (N_14501,N_7172,N_6613);
and U14502 (N_14502,N_6221,N_9495);
xnor U14503 (N_14503,N_9292,N_6188);
nor U14504 (N_14504,N_9100,N_8265);
nand U14505 (N_14505,N_7387,N_7291);
nand U14506 (N_14506,N_6675,N_6771);
and U14507 (N_14507,N_8100,N_6315);
nand U14508 (N_14508,N_6497,N_8538);
and U14509 (N_14509,N_5754,N_6856);
or U14510 (N_14510,N_6130,N_9203);
xnor U14511 (N_14511,N_5875,N_8196);
nor U14512 (N_14512,N_7975,N_9794);
nand U14513 (N_14513,N_6911,N_7641);
xnor U14514 (N_14514,N_7413,N_9899);
nor U14515 (N_14515,N_9204,N_5267);
xnor U14516 (N_14516,N_9104,N_9010);
or U14517 (N_14517,N_6152,N_9258);
or U14518 (N_14518,N_8761,N_6163);
and U14519 (N_14519,N_6312,N_5748);
and U14520 (N_14520,N_6528,N_8081);
nand U14521 (N_14521,N_7749,N_7369);
nor U14522 (N_14522,N_8825,N_8841);
or U14523 (N_14523,N_5836,N_9228);
and U14524 (N_14524,N_7063,N_6836);
or U14525 (N_14525,N_7084,N_8354);
nand U14526 (N_14526,N_9278,N_5292);
xor U14527 (N_14527,N_7854,N_7186);
or U14528 (N_14528,N_7741,N_8762);
xor U14529 (N_14529,N_7727,N_8653);
or U14530 (N_14530,N_6711,N_7636);
nand U14531 (N_14531,N_9117,N_5199);
or U14532 (N_14532,N_8360,N_8846);
nor U14533 (N_14533,N_5010,N_8251);
nand U14534 (N_14534,N_8252,N_7423);
nor U14535 (N_14535,N_5503,N_8604);
nand U14536 (N_14536,N_9586,N_7269);
xor U14537 (N_14537,N_9721,N_8941);
and U14538 (N_14538,N_5572,N_6192);
nand U14539 (N_14539,N_9326,N_5852);
or U14540 (N_14540,N_7561,N_9826);
and U14541 (N_14541,N_9880,N_6594);
xor U14542 (N_14542,N_6051,N_5123);
and U14543 (N_14543,N_8692,N_9643);
or U14544 (N_14544,N_7391,N_5099);
nor U14545 (N_14545,N_6816,N_5288);
nor U14546 (N_14546,N_7071,N_7694);
nand U14547 (N_14547,N_8332,N_6759);
and U14548 (N_14548,N_5481,N_9652);
and U14549 (N_14549,N_5404,N_5558);
or U14550 (N_14550,N_8129,N_7643);
and U14551 (N_14551,N_6705,N_7862);
nor U14552 (N_14552,N_7461,N_9385);
xor U14553 (N_14553,N_5148,N_9877);
and U14554 (N_14554,N_7085,N_5199);
or U14555 (N_14555,N_8147,N_7362);
nand U14556 (N_14556,N_5829,N_9987);
or U14557 (N_14557,N_8118,N_7022);
and U14558 (N_14558,N_9784,N_6160);
and U14559 (N_14559,N_5979,N_6945);
and U14560 (N_14560,N_7841,N_5937);
xor U14561 (N_14561,N_5126,N_8451);
nand U14562 (N_14562,N_5128,N_6663);
or U14563 (N_14563,N_9048,N_9304);
nand U14564 (N_14564,N_7577,N_6309);
nor U14565 (N_14565,N_7431,N_6213);
and U14566 (N_14566,N_9717,N_8151);
and U14567 (N_14567,N_6385,N_6046);
nor U14568 (N_14568,N_9866,N_5711);
nor U14569 (N_14569,N_5991,N_5535);
or U14570 (N_14570,N_6689,N_5185);
xnor U14571 (N_14571,N_8002,N_9406);
and U14572 (N_14572,N_9572,N_5663);
and U14573 (N_14573,N_8657,N_6262);
and U14574 (N_14574,N_6445,N_8311);
xnor U14575 (N_14575,N_7709,N_9239);
xnor U14576 (N_14576,N_9361,N_7452);
xnor U14577 (N_14577,N_9242,N_7872);
and U14578 (N_14578,N_8165,N_9093);
and U14579 (N_14579,N_8867,N_7412);
and U14580 (N_14580,N_8402,N_7383);
or U14581 (N_14581,N_9786,N_9887);
and U14582 (N_14582,N_5162,N_7616);
xor U14583 (N_14583,N_5522,N_8726);
nand U14584 (N_14584,N_8922,N_6121);
nor U14585 (N_14585,N_8879,N_6239);
nand U14586 (N_14586,N_9039,N_6162);
or U14587 (N_14587,N_8681,N_9199);
nor U14588 (N_14588,N_8333,N_9235);
nor U14589 (N_14589,N_8530,N_5536);
and U14590 (N_14590,N_6650,N_8870);
xnor U14591 (N_14591,N_5260,N_8071);
nor U14592 (N_14592,N_9304,N_5153);
xor U14593 (N_14593,N_6569,N_8962);
xnor U14594 (N_14594,N_8695,N_6932);
nor U14595 (N_14595,N_7309,N_6203);
nor U14596 (N_14596,N_8048,N_9239);
xor U14597 (N_14597,N_8453,N_8387);
xnor U14598 (N_14598,N_7419,N_5198);
or U14599 (N_14599,N_7349,N_7626);
or U14600 (N_14600,N_9335,N_5473);
and U14601 (N_14601,N_9032,N_8928);
xnor U14602 (N_14602,N_7529,N_6062);
nand U14603 (N_14603,N_6590,N_7618);
nand U14604 (N_14604,N_8270,N_9683);
or U14605 (N_14605,N_9589,N_7550);
xor U14606 (N_14606,N_8462,N_9296);
nor U14607 (N_14607,N_7729,N_7837);
or U14608 (N_14608,N_6117,N_5839);
nand U14609 (N_14609,N_8905,N_6102);
or U14610 (N_14610,N_7422,N_6252);
nand U14611 (N_14611,N_5964,N_6703);
and U14612 (N_14612,N_5171,N_6502);
xor U14613 (N_14613,N_9953,N_7327);
xnor U14614 (N_14614,N_6073,N_8094);
xor U14615 (N_14615,N_8265,N_6614);
nor U14616 (N_14616,N_6256,N_7939);
or U14617 (N_14617,N_7725,N_5757);
nor U14618 (N_14618,N_6557,N_8742);
xnor U14619 (N_14619,N_5899,N_9128);
nor U14620 (N_14620,N_9051,N_8770);
nor U14621 (N_14621,N_8002,N_7768);
and U14622 (N_14622,N_7155,N_5855);
and U14623 (N_14623,N_6283,N_6137);
nor U14624 (N_14624,N_9658,N_5136);
xor U14625 (N_14625,N_6163,N_6340);
xor U14626 (N_14626,N_9859,N_9109);
or U14627 (N_14627,N_7351,N_7151);
xnor U14628 (N_14628,N_6622,N_8326);
or U14629 (N_14629,N_8181,N_8286);
nand U14630 (N_14630,N_6120,N_5491);
or U14631 (N_14631,N_8971,N_5470);
and U14632 (N_14632,N_9580,N_5650);
nand U14633 (N_14633,N_5624,N_7764);
and U14634 (N_14634,N_8526,N_7093);
and U14635 (N_14635,N_8304,N_8241);
or U14636 (N_14636,N_9407,N_8408);
xor U14637 (N_14637,N_5415,N_8910);
nor U14638 (N_14638,N_7283,N_7795);
nand U14639 (N_14639,N_9568,N_5430);
nand U14640 (N_14640,N_5049,N_5679);
and U14641 (N_14641,N_7923,N_9412);
or U14642 (N_14642,N_6827,N_8909);
and U14643 (N_14643,N_5867,N_9670);
nand U14644 (N_14644,N_8467,N_7488);
xor U14645 (N_14645,N_5802,N_8542);
xor U14646 (N_14646,N_5512,N_6208);
xor U14647 (N_14647,N_6259,N_5752);
xnor U14648 (N_14648,N_8114,N_8911);
or U14649 (N_14649,N_9385,N_7480);
and U14650 (N_14650,N_9132,N_5416);
and U14651 (N_14651,N_5303,N_8666);
or U14652 (N_14652,N_5319,N_5026);
xor U14653 (N_14653,N_9125,N_5188);
nor U14654 (N_14654,N_5168,N_9888);
nor U14655 (N_14655,N_5424,N_7415);
xnor U14656 (N_14656,N_7632,N_7016);
nor U14657 (N_14657,N_6719,N_8113);
and U14658 (N_14658,N_6884,N_9848);
or U14659 (N_14659,N_9340,N_5569);
nand U14660 (N_14660,N_7896,N_6297);
nor U14661 (N_14661,N_9416,N_8468);
or U14662 (N_14662,N_7194,N_8527);
nand U14663 (N_14663,N_8018,N_7207);
and U14664 (N_14664,N_9764,N_6131);
or U14665 (N_14665,N_8378,N_6446);
and U14666 (N_14666,N_7358,N_6234);
nor U14667 (N_14667,N_6389,N_7068);
nor U14668 (N_14668,N_8228,N_7917);
nand U14669 (N_14669,N_7559,N_6175);
nor U14670 (N_14670,N_7054,N_9711);
xnor U14671 (N_14671,N_6831,N_9113);
nor U14672 (N_14672,N_5566,N_6320);
or U14673 (N_14673,N_8539,N_8713);
nor U14674 (N_14674,N_8058,N_8344);
or U14675 (N_14675,N_6075,N_8169);
xnor U14676 (N_14676,N_5066,N_8814);
or U14677 (N_14677,N_9940,N_8494);
nand U14678 (N_14678,N_9601,N_5578);
and U14679 (N_14679,N_6359,N_8453);
nor U14680 (N_14680,N_5737,N_6731);
or U14681 (N_14681,N_9649,N_9906);
xor U14682 (N_14682,N_9133,N_5504);
xor U14683 (N_14683,N_9510,N_8426);
nand U14684 (N_14684,N_9491,N_8750);
nor U14685 (N_14685,N_8437,N_8271);
or U14686 (N_14686,N_5729,N_8985);
nand U14687 (N_14687,N_5689,N_9552);
xor U14688 (N_14688,N_6076,N_8478);
nand U14689 (N_14689,N_6582,N_5580);
nor U14690 (N_14690,N_9163,N_8304);
and U14691 (N_14691,N_6374,N_7675);
nor U14692 (N_14692,N_5505,N_9091);
nand U14693 (N_14693,N_8380,N_6614);
nor U14694 (N_14694,N_8349,N_8901);
or U14695 (N_14695,N_6224,N_9130);
or U14696 (N_14696,N_5566,N_5761);
and U14697 (N_14697,N_6695,N_6031);
or U14698 (N_14698,N_9045,N_8038);
nor U14699 (N_14699,N_9116,N_7978);
nor U14700 (N_14700,N_5881,N_6463);
nor U14701 (N_14701,N_8027,N_6486);
and U14702 (N_14702,N_9038,N_5027);
xor U14703 (N_14703,N_6488,N_6159);
or U14704 (N_14704,N_5584,N_6314);
nand U14705 (N_14705,N_6396,N_9704);
nand U14706 (N_14706,N_8636,N_9332);
or U14707 (N_14707,N_8106,N_5018);
nor U14708 (N_14708,N_7477,N_9346);
xnor U14709 (N_14709,N_5222,N_8949);
or U14710 (N_14710,N_9652,N_7250);
nand U14711 (N_14711,N_5458,N_5478);
and U14712 (N_14712,N_6515,N_7007);
nand U14713 (N_14713,N_9767,N_7051);
xnor U14714 (N_14714,N_5551,N_8790);
xnor U14715 (N_14715,N_5914,N_9655);
and U14716 (N_14716,N_9802,N_7350);
nand U14717 (N_14717,N_9164,N_6354);
nor U14718 (N_14718,N_9294,N_7845);
nor U14719 (N_14719,N_7746,N_6812);
xor U14720 (N_14720,N_6797,N_8845);
nor U14721 (N_14721,N_8026,N_6730);
or U14722 (N_14722,N_7849,N_8532);
xnor U14723 (N_14723,N_6622,N_9137);
nand U14724 (N_14724,N_8386,N_8960);
and U14725 (N_14725,N_9332,N_6421);
xnor U14726 (N_14726,N_7004,N_5450);
and U14727 (N_14727,N_6808,N_6500);
nand U14728 (N_14728,N_7752,N_6999);
nand U14729 (N_14729,N_7409,N_7050);
nand U14730 (N_14730,N_7957,N_5878);
xor U14731 (N_14731,N_7002,N_6050);
and U14732 (N_14732,N_7631,N_5468);
xor U14733 (N_14733,N_5102,N_8903);
xor U14734 (N_14734,N_7283,N_5283);
nor U14735 (N_14735,N_9319,N_6795);
or U14736 (N_14736,N_9944,N_5371);
nand U14737 (N_14737,N_7656,N_6337);
or U14738 (N_14738,N_8967,N_5544);
xnor U14739 (N_14739,N_9233,N_5757);
or U14740 (N_14740,N_7591,N_9253);
nor U14741 (N_14741,N_8388,N_6132);
nor U14742 (N_14742,N_8515,N_9690);
or U14743 (N_14743,N_9468,N_6429);
xor U14744 (N_14744,N_9064,N_7328);
xor U14745 (N_14745,N_7333,N_5525);
nor U14746 (N_14746,N_6452,N_5406);
or U14747 (N_14747,N_7044,N_5915);
and U14748 (N_14748,N_6656,N_6358);
nand U14749 (N_14749,N_8400,N_7258);
and U14750 (N_14750,N_8345,N_9137);
or U14751 (N_14751,N_5075,N_5020);
nor U14752 (N_14752,N_7539,N_8201);
xor U14753 (N_14753,N_8962,N_5779);
and U14754 (N_14754,N_8698,N_8707);
xor U14755 (N_14755,N_8747,N_5594);
and U14756 (N_14756,N_7428,N_7148);
or U14757 (N_14757,N_8063,N_9515);
nand U14758 (N_14758,N_8172,N_9694);
nor U14759 (N_14759,N_7495,N_5373);
nor U14760 (N_14760,N_6051,N_7340);
or U14761 (N_14761,N_8640,N_8857);
and U14762 (N_14762,N_8428,N_7197);
and U14763 (N_14763,N_8699,N_8175);
nand U14764 (N_14764,N_7328,N_5718);
or U14765 (N_14765,N_6160,N_5289);
nor U14766 (N_14766,N_9884,N_8670);
and U14767 (N_14767,N_5021,N_9766);
nand U14768 (N_14768,N_5730,N_5495);
nand U14769 (N_14769,N_5442,N_6532);
and U14770 (N_14770,N_9440,N_6129);
nor U14771 (N_14771,N_6509,N_7157);
or U14772 (N_14772,N_5467,N_5097);
and U14773 (N_14773,N_8661,N_5197);
xnor U14774 (N_14774,N_7307,N_7373);
xnor U14775 (N_14775,N_7868,N_9965);
nand U14776 (N_14776,N_8624,N_5411);
nor U14777 (N_14777,N_5062,N_7284);
nor U14778 (N_14778,N_7129,N_5632);
xor U14779 (N_14779,N_5738,N_8598);
nand U14780 (N_14780,N_8841,N_6716);
and U14781 (N_14781,N_7470,N_5758);
and U14782 (N_14782,N_5837,N_6686);
and U14783 (N_14783,N_5031,N_8171);
xnor U14784 (N_14784,N_5783,N_7975);
nand U14785 (N_14785,N_8532,N_9926);
and U14786 (N_14786,N_7900,N_5901);
or U14787 (N_14787,N_6227,N_8271);
and U14788 (N_14788,N_7834,N_8578);
and U14789 (N_14789,N_8492,N_6333);
nor U14790 (N_14790,N_9435,N_9322);
or U14791 (N_14791,N_6009,N_9292);
nand U14792 (N_14792,N_8934,N_5975);
or U14793 (N_14793,N_5069,N_7222);
nand U14794 (N_14794,N_9184,N_7460);
or U14795 (N_14795,N_6769,N_6684);
nor U14796 (N_14796,N_7798,N_9510);
nand U14797 (N_14797,N_7982,N_9428);
or U14798 (N_14798,N_6456,N_9375);
xor U14799 (N_14799,N_9730,N_6706);
or U14800 (N_14800,N_6384,N_6284);
or U14801 (N_14801,N_9132,N_6271);
xnor U14802 (N_14802,N_8301,N_9303);
xnor U14803 (N_14803,N_7572,N_9249);
and U14804 (N_14804,N_8900,N_7493);
nor U14805 (N_14805,N_7140,N_6170);
and U14806 (N_14806,N_9646,N_9100);
nand U14807 (N_14807,N_9269,N_8731);
nor U14808 (N_14808,N_9327,N_5522);
nand U14809 (N_14809,N_7331,N_5303);
nand U14810 (N_14810,N_6986,N_7020);
and U14811 (N_14811,N_5947,N_8258);
and U14812 (N_14812,N_5280,N_6551);
and U14813 (N_14813,N_9489,N_6741);
or U14814 (N_14814,N_8745,N_8500);
or U14815 (N_14815,N_5510,N_5836);
or U14816 (N_14816,N_5227,N_7385);
nor U14817 (N_14817,N_7124,N_6702);
and U14818 (N_14818,N_6530,N_7287);
xnor U14819 (N_14819,N_9494,N_6242);
or U14820 (N_14820,N_7594,N_6814);
or U14821 (N_14821,N_9277,N_5898);
xor U14822 (N_14822,N_7896,N_6767);
nand U14823 (N_14823,N_7662,N_7546);
nor U14824 (N_14824,N_6347,N_8122);
and U14825 (N_14825,N_9930,N_5581);
nor U14826 (N_14826,N_6492,N_9959);
and U14827 (N_14827,N_9846,N_7045);
and U14828 (N_14828,N_6141,N_7605);
xnor U14829 (N_14829,N_8942,N_5344);
nor U14830 (N_14830,N_9543,N_7151);
or U14831 (N_14831,N_8607,N_9718);
and U14832 (N_14832,N_7548,N_9720);
and U14833 (N_14833,N_5514,N_6352);
nand U14834 (N_14834,N_5783,N_8457);
xnor U14835 (N_14835,N_7364,N_9565);
nand U14836 (N_14836,N_9040,N_8772);
or U14837 (N_14837,N_6898,N_7567);
or U14838 (N_14838,N_8223,N_7920);
xnor U14839 (N_14839,N_5068,N_8114);
nand U14840 (N_14840,N_6336,N_6129);
xnor U14841 (N_14841,N_8530,N_5369);
and U14842 (N_14842,N_8051,N_5247);
nor U14843 (N_14843,N_9414,N_8047);
xnor U14844 (N_14844,N_9362,N_6970);
xor U14845 (N_14845,N_5178,N_9936);
nor U14846 (N_14846,N_9155,N_8636);
nor U14847 (N_14847,N_6066,N_8297);
and U14848 (N_14848,N_8452,N_8740);
nand U14849 (N_14849,N_9814,N_5939);
nand U14850 (N_14850,N_8136,N_7641);
nand U14851 (N_14851,N_9033,N_7221);
or U14852 (N_14852,N_7204,N_8044);
xor U14853 (N_14853,N_7307,N_6934);
and U14854 (N_14854,N_8907,N_5470);
xor U14855 (N_14855,N_7215,N_9459);
and U14856 (N_14856,N_5411,N_6634);
and U14857 (N_14857,N_9533,N_9970);
or U14858 (N_14858,N_5874,N_6478);
nand U14859 (N_14859,N_8076,N_6369);
and U14860 (N_14860,N_8424,N_5418);
and U14861 (N_14861,N_5783,N_5548);
xnor U14862 (N_14862,N_9412,N_8918);
nor U14863 (N_14863,N_5024,N_8261);
nand U14864 (N_14864,N_9695,N_9859);
and U14865 (N_14865,N_7724,N_7463);
nand U14866 (N_14866,N_6443,N_9638);
xor U14867 (N_14867,N_7652,N_6746);
nor U14868 (N_14868,N_7476,N_9951);
and U14869 (N_14869,N_9570,N_9883);
or U14870 (N_14870,N_5539,N_9348);
nand U14871 (N_14871,N_7934,N_8330);
xnor U14872 (N_14872,N_7662,N_7531);
nor U14873 (N_14873,N_8934,N_9048);
or U14874 (N_14874,N_8094,N_5242);
nor U14875 (N_14875,N_7183,N_7405);
xor U14876 (N_14876,N_9216,N_9918);
or U14877 (N_14877,N_9371,N_5120);
xnor U14878 (N_14878,N_9355,N_6536);
nor U14879 (N_14879,N_7248,N_7643);
and U14880 (N_14880,N_9040,N_8597);
xnor U14881 (N_14881,N_9528,N_8414);
nand U14882 (N_14882,N_9065,N_5991);
nand U14883 (N_14883,N_9774,N_9919);
nand U14884 (N_14884,N_5601,N_6646);
or U14885 (N_14885,N_6379,N_9852);
xnor U14886 (N_14886,N_9157,N_6220);
nand U14887 (N_14887,N_8743,N_9444);
or U14888 (N_14888,N_5125,N_5321);
and U14889 (N_14889,N_8541,N_7609);
nand U14890 (N_14890,N_5954,N_8764);
nor U14891 (N_14891,N_6229,N_9679);
and U14892 (N_14892,N_8631,N_5184);
nor U14893 (N_14893,N_6872,N_9285);
nor U14894 (N_14894,N_9812,N_7669);
and U14895 (N_14895,N_5624,N_6365);
nand U14896 (N_14896,N_6643,N_7387);
nand U14897 (N_14897,N_5521,N_9375);
and U14898 (N_14898,N_6169,N_6749);
nor U14899 (N_14899,N_8440,N_7525);
and U14900 (N_14900,N_5414,N_7756);
xnor U14901 (N_14901,N_9560,N_6753);
xnor U14902 (N_14902,N_9942,N_5004);
or U14903 (N_14903,N_9288,N_6777);
nand U14904 (N_14904,N_9171,N_8758);
or U14905 (N_14905,N_7797,N_6197);
nor U14906 (N_14906,N_6151,N_5596);
or U14907 (N_14907,N_9268,N_6595);
and U14908 (N_14908,N_7462,N_6605);
nor U14909 (N_14909,N_5557,N_9770);
xnor U14910 (N_14910,N_9236,N_5406);
nand U14911 (N_14911,N_8509,N_6938);
nor U14912 (N_14912,N_9732,N_6293);
xnor U14913 (N_14913,N_6168,N_5554);
or U14914 (N_14914,N_5367,N_8071);
nor U14915 (N_14915,N_9226,N_7672);
or U14916 (N_14916,N_6844,N_7876);
nand U14917 (N_14917,N_7453,N_9104);
nand U14918 (N_14918,N_5409,N_5187);
xnor U14919 (N_14919,N_8929,N_6912);
nor U14920 (N_14920,N_5126,N_8333);
and U14921 (N_14921,N_8270,N_6640);
xor U14922 (N_14922,N_6788,N_6350);
or U14923 (N_14923,N_7824,N_8929);
nor U14924 (N_14924,N_5021,N_5363);
nand U14925 (N_14925,N_9296,N_7735);
and U14926 (N_14926,N_5133,N_7060);
and U14927 (N_14927,N_5590,N_8273);
or U14928 (N_14928,N_6276,N_7878);
nor U14929 (N_14929,N_7768,N_8381);
or U14930 (N_14930,N_9436,N_9153);
and U14931 (N_14931,N_9581,N_5846);
nor U14932 (N_14932,N_5669,N_8424);
nand U14933 (N_14933,N_8862,N_7346);
and U14934 (N_14934,N_8177,N_7066);
nor U14935 (N_14935,N_7787,N_6331);
and U14936 (N_14936,N_6965,N_8944);
nor U14937 (N_14937,N_8897,N_7008);
nor U14938 (N_14938,N_8395,N_5575);
xor U14939 (N_14939,N_9744,N_6576);
nand U14940 (N_14940,N_8934,N_7411);
and U14941 (N_14941,N_7786,N_7043);
xnor U14942 (N_14942,N_9839,N_7239);
xnor U14943 (N_14943,N_9722,N_8767);
nand U14944 (N_14944,N_8225,N_6408);
nor U14945 (N_14945,N_6241,N_5739);
and U14946 (N_14946,N_7279,N_9870);
nor U14947 (N_14947,N_8927,N_6009);
or U14948 (N_14948,N_8738,N_7689);
nand U14949 (N_14949,N_7365,N_5889);
nor U14950 (N_14950,N_8005,N_5124);
nand U14951 (N_14951,N_9838,N_6501);
or U14952 (N_14952,N_9039,N_7358);
and U14953 (N_14953,N_8874,N_5124);
xnor U14954 (N_14954,N_5366,N_6139);
nand U14955 (N_14955,N_9352,N_7629);
nor U14956 (N_14956,N_6382,N_9629);
or U14957 (N_14957,N_5924,N_5003);
nand U14958 (N_14958,N_5920,N_5896);
xnor U14959 (N_14959,N_7829,N_8899);
nand U14960 (N_14960,N_9205,N_9180);
nand U14961 (N_14961,N_5096,N_5068);
nand U14962 (N_14962,N_9620,N_6369);
xnor U14963 (N_14963,N_8880,N_8180);
nand U14964 (N_14964,N_8233,N_7538);
nor U14965 (N_14965,N_6928,N_9675);
and U14966 (N_14966,N_6891,N_5005);
nand U14967 (N_14967,N_5043,N_9586);
and U14968 (N_14968,N_9009,N_7515);
and U14969 (N_14969,N_5360,N_5328);
nor U14970 (N_14970,N_6174,N_7187);
nand U14971 (N_14971,N_8903,N_9551);
nor U14972 (N_14972,N_5689,N_5718);
nor U14973 (N_14973,N_5490,N_8895);
xnor U14974 (N_14974,N_9855,N_7906);
nor U14975 (N_14975,N_5210,N_6627);
nand U14976 (N_14976,N_8471,N_5960);
nand U14977 (N_14977,N_8989,N_9171);
xnor U14978 (N_14978,N_8545,N_6221);
nor U14979 (N_14979,N_9638,N_9097);
or U14980 (N_14980,N_6258,N_9340);
nand U14981 (N_14981,N_7354,N_5248);
and U14982 (N_14982,N_5105,N_7974);
nor U14983 (N_14983,N_6068,N_9907);
xor U14984 (N_14984,N_8561,N_8720);
and U14985 (N_14985,N_6944,N_9074);
and U14986 (N_14986,N_7054,N_9954);
and U14987 (N_14987,N_6110,N_8820);
nor U14988 (N_14988,N_7145,N_8447);
and U14989 (N_14989,N_9559,N_7371);
nor U14990 (N_14990,N_5081,N_9891);
nor U14991 (N_14991,N_8995,N_9790);
nand U14992 (N_14992,N_5684,N_9436);
and U14993 (N_14993,N_9194,N_5538);
and U14994 (N_14994,N_7780,N_7564);
and U14995 (N_14995,N_8406,N_9506);
or U14996 (N_14996,N_5017,N_6301);
nand U14997 (N_14997,N_6809,N_5880);
nand U14998 (N_14998,N_9989,N_9752);
xor U14999 (N_14999,N_6932,N_7587);
and U15000 (N_15000,N_14178,N_14799);
xnor U15001 (N_15001,N_13751,N_13307);
or U15002 (N_15002,N_12450,N_13743);
nand U15003 (N_15003,N_12723,N_13150);
nor U15004 (N_15004,N_13355,N_14617);
or U15005 (N_15005,N_10384,N_14082);
nand U15006 (N_15006,N_10918,N_10887);
nor U15007 (N_15007,N_13034,N_11146);
xnor U15008 (N_15008,N_10343,N_14759);
or U15009 (N_15009,N_14935,N_12800);
nor U15010 (N_15010,N_10685,N_14129);
nand U15011 (N_15011,N_10341,N_12710);
nand U15012 (N_15012,N_13461,N_12234);
nand U15013 (N_15013,N_12199,N_11319);
nor U15014 (N_15014,N_14830,N_11625);
xor U15015 (N_15015,N_14398,N_12842);
or U15016 (N_15016,N_12062,N_11426);
nor U15017 (N_15017,N_10060,N_11102);
nor U15018 (N_15018,N_10693,N_10418);
nor U15019 (N_15019,N_13117,N_10789);
or U15020 (N_15020,N_12014,N_13046);
or U15021 (N_15021,N_13844,N_10428);
or U15022 (N_15022,N_13599,N_12791);
nand U15023 (N_15023,N_11691,N_11989);
and U15024 (N_15024,N_12275,N_12492);
xnor U15025 (N_15025,N_10199,N_10217);
nor U15026 (N_15026,N_12099,N_11866);
xnor U15027 (N_15027,N_14580,N_10210);
or U15028 (N_15028,N_13540,N_12498);
nand U15029 (N_15029,N_13947,N_11499);
nand U15030 (N_15030,N_10301,N_12342);
xnor U15031 (N_15031,N_11757,N_10406);
or U15032 (N_15032,N_12712,N_14939);
or U15033 (N_15033,N_14681,N_14371);
xor U15034 (N_15034,N_10815,N_14290);
and U15035 (N_15035,N_12551,N_12088);
xnor U15036 (N_15036,N_10013,N_14737);
or U15037 (N_15037,N_13526,N_13183);
nor U15038 (N_15038,N_12749,N_14523);
nand U15039 (N_15039,N_14447,N_14784);
xor U15040 (N_15040,N_13240,N_10886);
nand U15041 (N_15041,N_13496,N_14825);
nand U15042 (N_15042,N_12726,N_14189);
or U15043 (N_15043,N_12966,N_13655);
nand U15044 (N_15044,N_12894,N_11111);
xnor U15045 (N_15045,N_12489,N_13939);
nor U15046 (N_15046,N_11799,N_14876);
nand U15047 (N_15047,N_14802,N_10419);
nand U15048 (N_15048,N_14285,N_14567);
nand U15049 (N_15049,N_14906,N_13032);
or U15050 (N_15050,N_12796,N_10345);
and U15051 (N_15051,N_11658,N_13741);
nand U15052 (N_15052,N_11399,N_11155);
nor U15053 (N_15053,N_12029,N_11020);
nand U15054 (N_15054,N_10166,N_12269);
nor U15055 (N_15055,N_12801,N_14659);
or U15056 (N_15056,N_13777,N_13267);
or U15057 (N_15057,N_14730,N_12019);
nor U15058 (N_15058,N_12636,N_11208);
nand U15059 (N_15059,N_14303,N_13852);
nand U15060 (N_15060,N_11404,N_11141);
or U15061 (N_15061,N_12613,N_14384);
nor U15062 (N_15062,N_11693,N_11096);
or U15063 (N_15063,N_14302,N_11117);
and U15064 (N_15064,N_11311,N_12627);
nor U15065 (N_15065,N_12882,N_11440);
xnor U15066 (N_15066,N_13624,N_10644);
nand U15067 (N_15067,N_13796,N_10973);
and U15068 (N_15068,N_13625,N_12438);
xor U15069 (N_15069,N_12428,N_12987);
nand U15070 (N_15070,N_10032,N_12709);
nor U15071 (N_15071,N_11082,N_10501);
xnor U15072 (N_15072,N_14305,N_10005);
xor U15073 (N_15073,N_13289,N_12421);
nand U15074 (N_15074,N_14150,N_13265);
nor U15075 (N_15075,N_12962,N_13611);
nor U15076 (N_15076,N_10881,N_12872);
and U15077 (N_15077,N_10022,N_13467);
nor U15078 (N_15078,N_14750,N_13366);
nand U15079 (N_15079,N_10938,N_12748);
xor U15080 (N_15080,N_10972,N_14902);
xnor U15081 (N_15081,N_10940,N_14268);
or U15082 (N_15082,N_13560,N_10328);
xor U15083 (N_15083,N_14550,N_12182);
xor U15084 (N_15084,N_10641,N_14708);
or U15085 (N_15085,N_11559,N_14872);
nand U15086 (N_15086,N_10425,N_11543);
nor U15087 (N_15087,N_14201,N_10643);
nand U15088 (N_15088,N_12189,N_12706);
nand U15089 (N_15089,N_10868,N_11685);
xor U15090 (N_15090,N_11118,N_10719);
or U15091 (N_15091,N_12971,N_12540);
and U15092 (N_15092,N_11126,N_12990);
xor U15093 (N_15093,N_13692,N_11151);
or U15094 (N_15094,N_10703,N_11002);
xnor U15095 (N_15095,N_12494,N_14787);
or U15096 (N_15096,N_13895,N_12402);
xnor U15097 (N_15097,N_14612,N_14110);
or U15098 (N_15098,N_11500,N_14814);
xor U15099 (N_15099,N_13563,N_13356);
nor U15100 (N_15100,N_10159,N_12389);
xnor U15101 (N_15101,N_13039,N_10064);
and U15102 (N_15102,N_13010,N_10389);
nand U15103 (N_15103,N_11986,N_13119);
nand U15104 (N_15104,N_14454,N_10051);
xnor U15105 (N_15105,N_13425,N_11938);
nor U15106 (N_15106,N_11527,N_11755);
nor U15107 (N_15107,N_11479,N_11392);
nand U15108 (N_15108,N_10556,N_12208);
nand U15109 (N_15109,N_13394,N_11664);
or U15110 (N_15110,N_11354,N_14630);
nand U15111 (N_15111,N_12352,N_12977);
and U15112 (N_15112,N_14130,N_11814);
nand U15113 (N_15113,N_11488,N_13343);
nand U15114 (N_15114,N_14450,N_11598);
nand U15115 (N_15115,N_12720,N_10714);
or U15116 (N_15116,N_11867,N_10490);
or U15117 (N_15117,N_11886,N_10848);
or U15118 (N_15118,N_13206,N_13063);
or U15119 (N_15119,N_13633,N_14918);
nand U15120 (N_15120,N_10371,N_12906);
nor U15121 (N_15121,N_12102,N_14931);
xnor U15122 (N_15122,N_11717,N_14419);
or U15123 (N_15123,N_12912,N_10000);
nand U15124 (N_15124,N_14278,N_11695);
nand U15125 (N_15125,N_10098,N_12171);
nand U15126 (N_15126,N_13249,N_11150);
xor U15127 (N_15127,N_14966,N_11475);
nand U15128 (N_15128,N_11184,N_14469);
or U15129 (N_15129,N_10441,N_11909);
nand U15130 (N_15130,N_11191,N_12694);
or U15131 (N_15131,N_14196,N_14696);
or U15132 (N_15132,N_13442,N_11337);
nor U15133 (N_15133,N_10144,N_10087);
nand U15134 (N_15134,N_12301,N_11729);
nor U15135 (N_15135,N_14312,N_11406);
and U15136 (N_15136,N_10566,N_10409);
and U15137 (N_15137,N_12158,N_14175);
or U15138 (N_15138,N_13301,N_14381);
xor U15139 (N_15139,N_11099,N_13190);
nand U15140 (N_15140,N_10110,N_12325);
nand U15141 (N_15141,N_14553,N_14838);
nor U15142 (N_15142,N_11130,N_13713);
and U15143 (N_15143,N_10924,N_11393);
or U15144 (N_15144,N_14800,N_10543);
xnor U15145 (N_15145,N_11144,N_14903);
nor U15146 (N_15146,N_12671,N_14829);
and U15147 (N_15147,N_14832,N_13836);
nor U15148 (N_15148,N_11346,N_13718);
or U15149 (N_15149,N_14275,N_13996);
and U15150 (N_15150,N_12594,N_12004);
xor U15151 (N_15151,N_14085,N_14555);
nand U15152 (N_15152,N_10382,N_10509);
xnor U15153 (N_15153,N_13326,N_11632);
or U15154 (N_15154,N_10932,N_13497);
nor U15155 (N_15155,N_14353,N_13932);
and U15156 (N_15156,N_10113,N_13234);
or U15157 (N_15157,N_14232,N_12861);
or U15158 (N_15158,N_14765,N_13327);
xor U15159 (N_15159,N_14342,N_11350);
xnor U15160 (N_15160,N_13440,N_11995);
nand U15161 (N_15161,N_14560,N_14531);
and U15162 (N_15162,N_14456,N_12967);
nor U15163 (N_15163,N_14247,N_13924);
and U15164 (N_15164,N_13035,N_10776);
xnor U15165 (N_15165,N_13538,N_14017);
or U15166 (N_15166,N_11927,N_10361);
nand U15167 (N_15167,N_12224,N_11171);
nor U15168 (N_15168,N_10598,N_14326);
and U15169 (N_15169,N_11396,N_12360);
or U15170 (N_15170,N_11865,N_11473);
nor U15171 (N_15171,N_10132,N_10127);
nor U15172 (N_15172,N_10024,N_10473);
and U15173 (N_15173,N_11302,N_10505);
or U15174 (N_15174,N_13084,N_10744);
and U15175 (N_15175,N_11548,N_13421);
or U15176 (N_15176,N_13480,N_11743);
and U15177 (N_15177,N_11216,N_12873);
or U15178 (N_15178,N_10901,N_12931);
nand U15179 (N_15179,N_12302,N_11160);
or U15180 (N_15180,N_13826,N_13772);
nand U15181 (N_15181,N_14936,N_12607);
nand U15182 (N_15182,N_14658,N_12898);
nor U15183 (N_15183,N_11149,N_12405);
nand U15184 (N_15184,N_12953,N_14265);
xor U15185 (N_15185,N_13458,N_11248);
and U15186 (N_15186,N_13885,N_11858);
xor U15187 (N_15187,N_11330,N_10727);
and U15188 (N_15188,N_14297,N_13170);
nand U15189 (N_15189,N_12160,N_12368);
nand U15190 (N_15190,N_10621,N_12771);
and U15191 (N_15191,N_10810,N_14923);
or U15192 (N_15192,N_14778,N_10062);
and U15193 (N_15193,N_10268,N_10679);
xor U15194 (N_15194,N_13709,N_10721);
xnor U15195 (N_15195,N_10966,N_11601);
nor U15196 (N_15196,N_12543,N_12164);
xor U15197 (N_15197,N_14788,N_11110);
or U15198 (N_15198,N_10209,N_10831);
and U15199 (N_15199,N_10321,N_13926);
or U15200 (N_15200,N_14688,N_13830);
xnor U15201 (N_15201,N_12612,N_10580);
nand U15202 (N_15202,N_14368,N_11095);
nor U15203 (N_15203,N_10423,N_13057);
or U15204 (N_15204,N_12338,N_11622);
and U15205 (N_15205,N_12683,N_13004);
or U15206 (N_15206,N_12697,N_14524);
nand U15207 (N_15207,N_13755,N_13522);
or U15208 (N_15208,N_11273,N_14393);
nand U15209 (N_15209,N_14960,N_11803);
xor U15210 (N_15210,N_11247,N_12386);
nor U15211 (N_15211,N_13521,N_11575);
or U15212 (N_15212,N_11620,N_10800);
or U15213 (N_15213,N_10451,N_11097);
nor U15214 (N_15214,N_11763,N_10385);
nand U15215 (N_15215,N_10174,N_10877);
and U15216 (N_15216,N_13834,N_13971);
nor U15217 (N_15217,N_14723,N_14719);
and U15218 (N_15218,N_11566,N_13665);
or U15219 (N_15219,N_12241,N_12954);
nor U15220 (N_15220,N_10525,N_11778);
nand U15221 (N_15221,N_12985,N_13260);
and U15222 (N_15222,N_13101,N_11198);
nor U15223 (N_15223,N_14164,N_12226);
nor U15224 (N_15224,N_10760,N_10250);
or U15225 (N_15225,N_10965,N_13431);
nand U15226 (N_15226,N_12702,N_10284);
xor U15227 (N_15227,N_11568,N_12657);
and U15228 (N_15228,N_10526,N_13349);
nor U15229 (N_15229,N_14241,N_13871);
xor U15230 (N_15230,N_13629,N_12351);
xnor U15231 (N_15231,N_14508,N_14894);
and U15232 (N_15232,N_12391,N_10373);
and U15233 (N_15233,N_13095,N_10033);
or U15234 (N_15234,N_13827,N_13818);
xor U15235 (N_15235,N_14539,N_10656);
xnor U15236 (N_15236,N_10185,N_11914);
nor U15237 (N_15237,N_14764,N_13545);
nor U15238 (N_15238,N_10813,N_14392);
nor U15239 (N_15239,N_12643,N_13085);
nor U15240 (N_15240,N_14103,N_14760);
nand U15241 (N_15241,N_14233,N_12205);
xor U15242 (N_15242,N_11035,N_12409);
nand U15243 (N_15243,N_13438,N_12526);
xnor U15244 (N_15244,N_10456,N_10858);
or U15245 (N_15245,N_13104,N_10657);
and U15246 (N_15246,N_10704,N_14027);
xor U15247 (N_15247,N_11700,N_12291);
xor U15248 (N_15248,N_14137,N_11573);
xor U15249 (N_15249,N_12908,N_12343);
and U15250 (N_15250,N_11895,N_14350);
nand U15251 (N_15251,N_12120,N_14237);
nor U15252 (N_15252,N_11551,N_10592);
and U15253 (N_15253,N_12106,N_10133);
xor U15254 (N_15254,N_12186,N_13570);
nand U15255 (N_15255,N_11599,N_13965);
and U15256 (N_15256,N_12948,N_10500);
and U15257 (N_15257,N_12737,N_12765);
nor U15258 (N_15258,N_12986,N_14004);
and U15259 (N_15259,N_13378,N_10890);
nor U15260 (N_15260,N_10928,N_12168);
nand U15261 (N_15261,N_10583,N_10529);
nor U15262 (N_15262,N_11048,N_12693);
xnor U15263 (N_15263,N_10307,N_12395);
nor U15264 (N_15264,N_10767,N_10817);
xnor U15265 (N_15265,N_10731,N_14645);
xnor U15266 (N_15266,N_11892,N_10909);
nand U15267 (N_15267,N_13679,N_12200);
nand U15268 (N_15268,N_13177,N_11434);
or U15269 (N_15269,N_12745,N_11720);
xor U15270 (N_15270,N_11244,N_13581);
nor U15271 (N_15271,N_10988,N_12022);
nand U15272 (N_15272,N_14308,N_10460);
and U15273 (N_15273,N_14083,N_10053);
or U15274 (N_15274,N_14074,N_14286);
or U15275 (N_15275,N_11969,N_10978);
nand U15276 (N_15276,N_12432,N_10646);
and U15277 (N_15277,N_11315,N_11194);
nor U15278 (N_15278,N_14924,N_11574);
and U15279 (N_15279,N_11080,N_14208);
nand U15280 (N_15280,N_12115,N_11924);
and U15281 (N_15281,N_10093,N_11061);
xor U15282 (N_15282,N_12258,N_10686);
or U15283 (N_15283,N_11467,N_14486);
and U15284 (N_15284,N_12760,N_10180);
nand U15285 (N_15285,N_12167,N_11761);
and U15286 (N_15286,N_12778,N_10593);
and U15287 (N_15287,N_14458,N_12490);
xnor U15288 (N_15288,N_12777,N_11973);
nand U15289 (N_15289,N_13166,N_11493);
xnor U15290 (N_15290,N_14881,N_12349);
nor U15291 (N_15291,N_11432,N_10778);
nand U15292 (N_15292,N_11943,N_12978);
or U15293 (N_15293,N_10129,N_11231);
and U15294 (N_15294,N_14430,N_11207);
nand U15295 (N_15295,N_12895,N_13649);
and U15296 (N_15296,N_10177,N_14457);
or U15297 (N_15297,N_13091,N_14711);
xnor U15298 (N_15298,N_12844,N_13300);
xnor U15299 (N_15299,N_12910,N_14360);
xnor U15300 (N_15300,N_14597,N_13200);
and U15301 (N_15301,N_14141,N_10066);
nand U15302 (N_15302,N_14335,N_11565);
and U15303 (N_15303,N_11830,N_12864);
or U15304 (N_15304,N_13319,N_12111);
nand U15305 (N_15305,N_12462,N_13102);
and U15306 (N_15306,N_13475,N_13168);
xnor U15307 (N_15307,N_14172,N_11848);
or U15308 (N_15308,N_11526,N_12121);
nor U15309 (N_15309,N_14819,N_12052);
nor U15310 (N_15310,N_12630,N_11400);
nand U15311 (N_15311,N_10452,N_13710);
xor U15312 (N_15312,N_11712,N_12030);
or U15313 (N_15313,N_14061,N_13353);
or U15314 (N_15314,N_10926,N_12118);
xor U15315 (N_15315,N_12312,N_13833);
nand U15316 (N_15316,N_14926,N_10216);
or U15317 (N_15317,N_12843,N_12220);
nor U15318 (N_15318,N_10707,N_10619);
nor U15319 (N_15319,N_14258,N_11544);
xnor U15320 (N_15320,N_10194,N_14151);
xor U15321 (N_15321,N_12590,N_12027);
nand U15322 (N_15322,N_10483,N_14938);
or U15323 (N_15323,N_11039,N_12708);
xor U15324 (N_15324,N_14420,N_11287);
and U15325 (N_15325,N_10981,N_13262);
xnor U15326 (N_15326,N_13857,N_14041);
or U15327 (N_15327,N_11368,N_13550);
and U15328 (N_15328,N_14763,N_14562);
xor U15329 (N_15329,N_14476,N_11863);
xnor U15330 (N_15330,N_13116,N_14768);
nor U15331 (N_15331,N_11293,N_10557);
and U15332 (N_15332,N_14714,N_10884);
nor U15333 (N_15333,N_11576,N_10453);
and U15334 (N_15334,N_11379,N_10709);
or U15335 (N_15335,N_14490,N_11294);
nand U15336 (N_15336,N_14994,N_14383);
nor U15337 (N_15337,N_11724,N_11905);
and U15338 (N_15338,N_11193,N_11896);
or U15339 (N_15339,N_13987,N_12707);
or U15340 (N_15340,N_11859,N_12501);
xnor U15341 (N_15341,N_13683,N_10058);
nand U15342 (N_15342,N_12431,N_13992);
and U15343 (N_15343,N_11425,N_10647);
nand U15344 (N_15344,N_10521,N_10499);
nor U15345 (N_15345,N_11525,N_12806);
xnor U15346 (N_15346,N_10450,N_11617);
nand U15347 (N_15347,N_12392,N_12236);
nand U15348 (N_15348,N_13731,N_14274);
xor U15349 (N_15349,N_13769,N_12812);
nor U15350 (N_15350,N_13452,N_10038);
or U15351 (N_15351,N_10235,N_10045);
nand U15352 (N_15352,N_11329,N_14394);
and U15353 (N_15353,N_10663,N_10690);
xnor U15354 (N_15354,N_14611,N_13093);
or U15355 (N_15355,N_13955,N_12877);
and U15356 (N_15356,N_10176,N_11104);
xor U15357 (N_15357,N_12684,N_10394);
nand U15358 (N_15358,N_12065,N_11148);
nand U15359 (N_15359,N_11898,N_10114);
nor U15360 (N_15360,N_11648,N_10444);
nor U15361 (N_15361,N_14843,N_14549);
or U15362 (N_15362,N_12348,N_14943);
and U15363 (N_15363,N_14299,N_12834);
and U15364 (N_15364,N_14281,N_11623);
xnor U15365 (N_15365,N_14889,N_13215);
or U15366 (N_15366,N_11832,N_11063);
xnor U15367 (N_15367,N_12824,N_13055);
and U15368 (N_15368,N_14435,N_12646);
xnor U15369 (N_15369,N_14417,N_13621);
xor U15370 (N_15370,N_10358,N_13041);
xor U15371 (N_15371,N_13840,N_11305);
or U15372 (N_15372,N_11619,N_12488);
nand U15373 (N_15373,N_10290,N_10173);
and U15374 (N_15374,N_14228,N_10870);
nor U15375 (N_15375,N_14815,N_11255);
nor U15376 (N_15376,N_10838,N_10678);
and U15377 (N_15377,N_11779,N_13925);
xnor U15378 (N_15378,N_10157,N_13586);
and U15379 (N_15379,N_13388,N_14331);
and U15380 (N_15380,N_14410,N_12570);
and U15381 (N_15381,N_12394,N_13567);
xnor U15382 (N_15382,N_13359,N_13362);
nor U15383 (N_15383,N_11621,N_13537);
nand U15384 (N_15384,N_10183,N_13943);
nor U15385 (N_15385,N_11139,N_10262);
and U15386 (N_15386,N_12609,N_12309);
nand U15387 (N_15387,N_10796,N_14259);
nor U15388 (N_15388,N_14856,N_10211);
xor U15389 (N_15389,N_12519,N_11897);
or U15390 (N_15390,N_10604,N_14239);
and U15391 (N_15391,N_13436,N_10003);
nor U15392 (N_15392,N_10849,N_12610);
and U15393 (N_15393,N_14969,N_10416);
or U15394 (N_15394,N_13798,N_13509);
xor U15395 (N_15395,N_11366,N_13174);
nand U15396 (N_15396,N_12107,N_12276);
and U15397 (N_15397,N_10458,N_14808);
nand U15398 (N_15398,N_10930,N_14927);
and U15399 (N_15399,N_10370,N_12562);
xnor U15400 (N_15400,N_14615,N_12383);
and U15401 (N_15401,N_10238,N_11046);
nor U15402 (N_15402,N_12981,N_12614);
or U15403 (N_15403,N_13324,N_14874);
nand U15404 (N_15404,N_12449,N_13974);
nand U15405 (N_15405,N_10794,N_12900);
nor U15406 (N_15406,N_12686,N_13697);
nor U15407 (N_15407,N_13429,N_12297);
nor U15408 (N_15408,N_11558,N_12204);
and U15409 (N_15409,N_14098,N_11744);
nor U15410 (N_15410,N_10811,N_12142);
and U15411 (N_15411,N_11569,N_13179);
or U15412 (N_15412,N_10336,N_10737);
nand U15413 (N_15413,N_14461,N_13428);
nor U15414 (N_15414,N_11522,N_10626);
nand U15415 (N_15415,N_12346,N_11441);
and U15416 (N_15416,N_14003,N_14442);
or U15417 (N_15417,N_13400,N_10883);
nor U15418 (N_15418,N_14485,N_10056);
nor U15419 (N_15419,N_12157,N_11667);
nor U15420 (N_15420,N_14244,N_13571);
or U15421 (N_15421,N_12850,N_10705);
xnor U15422 (N_15422,N_13828,N_11663);
nor U15423 (N_15423,N_13899,N_10182);
and U15424 (N_15424,N_10306,N_13450);
nand U15425 (N_15425,N_13862,N_11815);
xor U15426 (N_15426,N_14160,N_11480);
nand U15427 (N_15427,N_10606,N_11413);
nand U15428 (N_15428,N_12270,N_14627);
or U15429 (N_15429,N_14373,N_12165);
xor U15430 (N_15430,N_11917,N_12375);
xor U15431 (N_15431,N_11060,N_10152);
nand U15432 (N_15432,N_12382,N_11183);
nor U15433 (N_15433,N_10624,N_10079);
or U15434 (N_15434,N_14761,N_13244);
nor U15435 (N_15435,N_12403,N_10750);
xor U15436 (N_15436,N_13700,N_10960);
xor U15437 (N_15437,N_10330,N_14691);
and U15438 (N_15438,N_14411,N_14873);
and U15439 (N_15439,N_10272,N_13719);
and U15440 (N_15440,N_11173,N_14010);
and U15441 (N_15441,N_14229,N_14097);
and U15442 (N_15442,N_14434,N_10929);
and U15443 (N_15443,N_13884,N_12530);
and U15444 (N_15444,N_12175,N_10314);
nor U15445 (N_15445,N_14493,N_13776);
nand U15446 (N_15446,N_12510,N_11359);
nand U15447 (N_15447,N_14128,N_13444);
or U15448 (N_15448,N_11062,N_10354);
xnor U15449 (N_15449,N_14727,N_12716);
and U15450 (N_15450,N_12776,N_12251);
and U15451 (N_15451,N_13077,N_13515);
nand U15452 (N_15452,N_14124,N_14610);
xnor U15453 (N_15453,N_10855,N_14365);
and U15454 (N_15454,N_13261,N_11230);
and U15455 (N_15455,N_13859,N_12629);
or U15456 (N_15456,N_10324,N_12670);
xor U15457 (N_15457,N_13280,N_11659);
nor U15458 (N_15458,N_14415,N_11510);
nand U15459 (N_15459,N_13835,N_13744);
and U15460 (N_15460,N_10491,N_11971);
nand U15461 (N_15461,N_11785,N_13361);
xor U15462 (N_15462,N_12642,N_13125);
xnor U15463 (N_15463,N_13654,N_13439);
xor U15464 (N_15464,N_14257,N_12534);
or U15465 (N_15465,N_14868,N_13533);
xnor U15466 (N_15466,N_14197,N_13294);
and U15467 (N_15467,N_10313,N_13671);
xnor U15468 (N_15468,N_14766,N_13456);
nor U15469 (N_15469,N_13381,N_12597);
nor U15470 (N_15470,N_10323,N_14826);
nand U15471 (N_15471,N_14385,N_10964);
nor U15472 (N_15472,N_14670,N_12997);
and U15473 (N_15473,N_14706,N_13008);
nand U15474 (N_15474,N_13787,N_11105);
or U15475 (N_15475,N_13462,N_14589);
and U15476 (N_15476,N_13304,N_14882);
and U15477 (N_15477,N_12867,N_10148);
or U15478 (N_15478,N_12905,N_13573);
and U15479 (N_15479,N_10091,N_12180);
nor U15480 (N_15480,N_10522,N_12412);
and U15481 (N_15481,N_10432,N_13345);
or U15482 (N_15482,N_11236,N_10193);
nor U15483 (N_15483,N_11388,N_13688);
xnor U15484 (N_15484,N_12439,N_10048);
or U15485 (N_15485,N_14336,N_14852);
and U15486 (N_15486,N_11052,N_12538);
or U15487 (N_15487,N_10535,N_11857);
or U15488 (N_15488,N_11324,N_14520);
nor U15489 (N_15489,N_10618,N_11474);
nand U15490 (N_15490,N_14254,N_10864);
and U15491 (N_15491,N_11835,N_13645);
and U15492 (N_15492,N_10463,N_11214);
nand U15493 (N_15493,N_12440,N_12659);
nor U15494 (N_15494,N_10899,N_14724);
nor U15495 (N_15495,N_14579,N_11394);
nor U15496 (N_15496,N_14685,N_11817);
and U15497 (N_15497,N_12685,N_11999);
nor U15498 (N_15498,N_12416,N_14592);
and U15499 (N_15499,N_11732,N_13404);
xnor U15500 (N_15500,N_14263,N_13569);
nor U15501 (N_15501,N_11899,N_14609);
xnor U15502 (N_15502,N_11307,N_10962);
and U15503 (N_15503,N_14112,N_12921);
and U15504 (N_15504,N_11931,N_14642);
nor U15505 (N_15505,N_14492,N_14619);
xor U15506 (N_15506,N_13157,N_13724);
nand U15507 (N_15507,N_13220,N_11353);
xor U15508 (N_15508,N_14015,N_13016);
xnor U15509 (N_15509,N_14644,N_12715);
and U15510 (N_15510,N_13303,N_11810);
or U15511 (N_15511,N_14180,N_13099);
and U15512 (N_15512,N_10508,N_11395);
xnor U15513 (N_15513,N_10387,N_12444);
xnor U15514 (N_15514,N_12536,N_10061);
nor U15515 (N_15515,N_10562,N_11026);
xor U15516 (N_15516,N_14726,N_11683);
or U15517 (N_15517,N_10923,N_12766);
xor U15518 (N_15518,N_14292,N_12056);
nand U15519 (N_15519,N_12193,N_10523);
nand U15520 (N_15520,N_14715,N_11627);
and U15521 (N_15521,N_10627,N_12914);
or U15522 (N_15522,N_11541,N_13075);
or U15523 (N_15523,N_10191,N_14947);
nor U15524 (N_15524,N_14222,N_10026);
xnor U15525 (N_15525,N_12188,N_14816);
or U15526 (N_15526,N_13952,N_11812);
nor U15527 (N_15527,N_10950,N_12314);
nor U15528 (N_15528,N_13295,N_10758);
or U15529 (N_15529,N_10167,N_14162);
or U15530 (N_15530,N_12733,N_14684);
or U15531 (N_15531,N_14352,N_13288);
or U15532 (N_15532,N_14198,N_13580);
nand U15533 (N_15533,N_10459,N_10747);
nand U15534 (N_15534,N_12470,N_11801);
nor U15535 (N_15535,N_13805,N_12257);
and U15536 (N_15536,N_11920,N_10919);
nand U15537 (N_15537,N_13318,N_14806);
nand U15538 (N_15538,N_14482,N_11014);
nand U15539 (N_15539,N_12072,N_13370);
or U15540 (N_15540,N_10516,N_12696);
nand U15541 (N_15541,N_13194,N_13914);
and U15542 (N_15542,N_12384,N_11553);
nand U15543 (N_15543,N_10320,N_13508);
nor U15544 (N_15544,N_14131,N_14203);
xor U15545 (N_15545,N_10340,N_12362);
xor U15546 (N_15546,N_12289,N_13453);
nor U15547 (N_15547,N_13790,N_10741);
nand U15548 (N_15548,N_13457,N_12545);
or U15549 (N_15549,N_14176,N_13178);
xnor U15550 (N_15550,N_12340,N_11825);
xor U15551 (N_15551,N_13419,N_13962);
or U15552 (N_15552,N_11735,N_11768);
nor U15553 (N_15553,N_11361,N_11420);
nand U15554 (N_15554,N_13948,N_11703);
or U15555 (N_15555,N_13762,N_14672);
and U15556 (N_15556,N_11719,N_13158);
or U15557 (N_15557,N_14051,N_12768);
and U15558 (N_15558,N_12074,N_10445);
or U15559 (N_15559,N_14246,N_10305);
or U15560 (N_15560,N_12013,N_11570);
nand U15561 (N_15561,N_14917,N_14181);
nand U15562 (N_15562,N_14603,N_13893);
and U15563 (N_15563,N_11089,N_14713);
nand U15564 (N_15564,N_14340,N_14296);
nor U15565 (N_15565,N_11129,N_12154);
or U15566 (N_15566,N_10970,N_14171);
nor U15567 (N_15567,N_13412,N_11027);
or U15568 (N_15568,N_12947,N_12425);
xnor U15569 (N_15569,N_12119,N_14845);
nand U15570 (N_15570,N_14102,N_14961);
nand U15571 (N_15571,N_11053,N_12316);
and U15572 (N_15572,N_11265,N_14138);
xor U15573 (N_15573,N_12836,N_11745);
or U15574 (N_15574,N_10958,N_13137);
nand U15575 (N_15575,N_14123,N_13367);
or U15576 (N_15576,N_12145,N_12255);
nand U15577 (N_15577,N_13314,N_10489);
nand U15578 (N_15578,N_12937,N_12732);
nor U15579 (N_15579,N_10772,N_14797);
or U15580 (N_15580,N_13883,N_12831);
nor U15581 (N_15581,N_12284,N_12079);
or U15582 (N_15582,N_14270,N_12058);
and U15583 (N_15583,N_10878,N_10135);
and U15584 (N_15584,N_12991,N_14416);
xnor U15585 (N_15585,N_11088,N_14401);
or U15586 (N_15586,N_10186,N_14252);
nand U15587 (N_15587,N_10150,N_14387);
nor U15588 (N_15588,N_12741,N_14341);
nand U15589 (N_15589,N_12077,N_11472);
nand U15590 (N_15590,N_10649,N_14170);
xor U15591 (N_15591,N_10485,N_11654);
nand U15592 (N_15592,N_10540,N_13636);
xor U15593 (N_15593,N_12277,N_13141);
and U15594 (N_15594,N_11131,N_10588);
nand U15595 (N_15595,N_12047,N_13618);
nand U15596 (N_15596,N_14835,N_12653);
nand U15597 (N_15597,N_13347,N_11636);
xnor U15598 (N_15598,N_13905,N_13706);
and U15599 (N_15599,N_11878,N_12288);
nand U15600 (N_15600,N_12303,N_11980);
nor U15601 (N_15601,N_14443,N_11463);
nor U15602 (N_15602,N_11269,N_13309);
and U15603 (N_15603,N_13729,N_14020);
xnor U15604 (N_15604,N_12995,N_13210);
xor U15605 (N_15605,N_13596,N_12020);
or U15606 (N_15606,N_12336,N_13484);
and U15607 (N_15607,N_12666,N_14746);
nor U15608 (N_15608,N_11747,N_12372);
and U15609 (N_15609,N_11197,N_13385);
nor U15610 (N_15610,N_10407,N_10348);
nand U15611 (N_15611,N_11579,N_14223);
nor U15612 (N_15612,N_13896,N_10533);
nand U15613 (N_15613,N_12976,N_12883);
nor U15614 (N_15614,N_14216,N_12717);
nand U15615 (N_15615,N_13072,N_10298);
nor U15616 (N_15616,N_10882,N_11618);
nand U15617 (N_15617,N_10271,N_13045);
xnor U15618 (N_15618,N_11107,N_12135);
nand U15619 (N_15619,N_11070,N_11701);
nor U15620 (N_15620,N_12243,N_10146);
or U15621 (N_15621,N_13615,N_11612);
and U15622 (N_15622,N_10814,N_12734);
and U15623 (N_15623,N_14586,N_10997);
xor U15624 (N_15624,N_13292,N_12485);
nor U15625 (N_15625,N_13493,N_11811);
and U15626 (N_15626,N_14565,N_13513);
or U15627 (N_15627,N_14516,N_11733);
xnor U15628 (N_15628,N_11725,N_13911);
nand U15629 (N_15629,N_12794,N_12411);
xor U15630 (N_15630,N_14188,N_11127);
or U15631 (N_15631,N_10665,N_12690);
or U15632 (N_15632,N_13670,N_13504);
xor U15633 (N_15633,N_10659,N_13471);
or U15634 (N_15634,N_11809,N_12730);
nand U15635 (N_15635,N_12133,N_14052);
or U15636 (N_15636,N_11588,N_13708);
xnor U15637 (N_15637,N_14261,N_13323);
and U15638 (N_15638,N_11501,N_11823);
nand U15639 (N_15639,N_14899,N_12127);
nor U15640 (N_15640,N_14515,N_12637);
or U15641 (N_15641,N_13845,N_12153);
nand U15642 (N_15642,N_12083,N_13232);
or U15643 (N_15643,N_13891,N_14517);
and U15644 (N_15644,N_10820,N_14320);
and U15645 (N_15645,N_10718,N_11028);
xnor U15646 (N_15646,N_10948,N_14911);
nand U15647 (N_15647,N_11790,N_11535);
and U15648 (N_15648,N_10987,N_10078);
nand U15649 (N_15649,N_13953,N_12472);
nor U15650 (N_15650,N_11954,N_12820);
and U15651 (N_15651,N_13842,N_12600);
nor U15652 (N_15652,N_13799,N_11478);
xor U15653 (N_15653,N_14949,N_14530);
and U15654 (N_15654,N_14841,N_13779);
or U15655 (N_15655,N_11912,N_13960);
nor U15656 (N_15656,N_13752,N_11949);
or U15657 (N_15657,N_14654,N_13238);
nor U15658 (N_15658,N_10706,N_10573);
and U15659 (N_15659,N_12330,N_13111);
nand U15660 (N_15660,N_12930,N_13082);
and U15661 (N_15661,N_13674,N_13809);
nor U15662 (N_15662,N_10668,N_14289);
nand U15663 (N_15663,N_10004,N_12839);
nand U15664 (N_15664,N_10118,N_14480);
xor U15665 (N_15665,N_12926,N_10270);
xor U15666 (N_15666,N_12274,N_11585);
xor U15667 (N_15667,N_14590,N_14844);
or U15668 (N_15668,N_11290,N_12869);
xor U15669 (N_15669,N_12248,N_11939);
nor U15670 (N_15670,N_11534,N_10147);
or U15671 (N_15671,N_12758,N_13640);
xnor U15672 (N_15672,N_11401,N_14412);
and U15673 (N_15673,N_11524,N_13464);
xnor U15674 (N_15674,N_14921,N_12959);
and U15675 (N_15675,N_11891,N_11765);
nand U15676 (N_15676,N_12875,N_11270);
nand U15677 (N_15677,N_10755,N_12576);
nor U15678 (N_15678,N_14731,N_10339);
and U15679 (N_15679,N_12786,N_13191);
nor U15680 (N_15680,N_13276,N_10140);
nand U15681 (N_15681,N_14090,N_10565);
and U15682 (N_15682,N_11655,N_14739);
xor U15683 (N_15683,N_12890,N_10792);
and U15684 (N_15684,N_10857,N_12306);
and U15685 (N_15685,N_10998,N_11457);
and U15686 (N_15686,N_11291,N_11443);
nand U15687 (N_15687,N_10429,N_14984);
xor U15688 (N_15688,N_12051,N_12093);
xnor U15689 (N_15689,N_13219,N_13189);
and U15690 (N_15690,N_11257,N_10843);
or U15691 (N_15691,N_13216,N_12772);
nor U15692 (N_15692,N_10720,N_11232);
or U15693 (N_15693,N_10130,N_12729);
nand U15694 (N_15694,N_14937,N_11748);
xor U15695 (N_15695,N_12569,N_10795);
or U15696 (N_15696,N_11157,N_10481);
and U15697 (N_15697,N_11731,N_11992);
xnor U15698 (N_15698,N_11687,N_11981);
nand U15699 (N_15699,N_12999,N_14380);
and U15700 (N_15700,N_13589,N_14756);
and U15701 (N_15701,N_12790,N_14184);
nand U15702 (N_15702,N_10232,N_11607);
nor U15703 (N_15703,N_11182,N_10829);
and U15704 (N_15704,N_12747,N_14907);
nand U15705 (N_15705,N_13934,N_12752);
and U15706 (N_15706,N_11122,N_10654);
or U15707 (N_15707,N_14646,N_10824);
or U15708 (N_15708,N_13118,N_11958);
nand U15709 (N_15709,N_11398,N_14348);
or U15710 (N_15710,N_13676,N_13770);
xnor U15711 (N_15711,N_11128,N_10391);
or U15712 (N_15712,N_13663,N_14640);
nand U15713 (N_15713,N_10070,N_11482);
nor U15714 (N_15714,N_13163,N_12884);
or U15715 (N_15715,N_13208,N_14230);
or U15716 (N_15716,N_13864,N_12584);
or U15717 (N_15717,N_12893,N_13585);
nor U15718 (N_15718,N_12994,N_10833);
or U15719 (N_15719,N_10297,N_13005);
xor U15720 (N_15720,N_13678,N_13623);
xnor U15721 (N_15721,N_14429,N_10691);
nand U15722 (N_15722,N_10124,N_11429);
and U15723 (N_15723,N_14242,N_12499);
nand U15724 (N_15724,N_11323,N_14709);
or U15725 (N_15725,N_14818,N_13494);
and U15726 (N_15726,N_14432,N_11657);
nor U15727 (N_15727,N_12979,N_10922);
nor U15728 (N_15728,N_13126,N_12032);
or U15729 (N_15729,N_13921,N_14745);
and U15730 (N_15730,N_13320,N_13352);
or U15731 (N_15731,N_12662,N_10438);
nor U15732 (N_15732,N_12502,N_14140);
and U15733 (N_15733,N_12265,N_11133);
nand U15734 (N_15734,N_11040,N_10196);
xnor U15735 (N_15735,N_10123,N_11932);
nand U15736 (N_15736,N_14699,N_11494);
nor U15737 (N_15737,N_11364,N_14992);
nand U15738 (N_15738,N_11961,N_13002);
nand U15739 (N_15739,N_10688,N_12982);
or U15740 (N_15740,N_10101,N_14925);
and U15741 (N_15741,N_12143,N_12380);
and U15742 (N_15742,N_12009,N_13881);
or U15743 (N_15743,N_13546,N_14993);
nand U15744 (N_15744,N_12059,N_10967);
or U15745 (N_15745,N_14616,N_11517);
nand U15746 (N_15746,N_14050,N_12669);
xor U15747 (N_15747,N_12652,N_10037);
nand U15748 (N_15748,N_14667,N_13967);
and U15749 (N_15749,N_12326,N_11454);
nor U15750 (N_15750,N_10326,N_14668);
and U15751 (N_15751,N_13721,N_13114);
nor U15752 (N_15752,N_12374,N_14031);
or U15753 (N_15753,N_12533,N_10819);
xor U15754 (N_15754,N_13747,N_12549);
nor U15755 (N_15755,N_13340,N_13549);
or U15756 (N_15756,N_10850,N_10049);
and U15757 (N_15757,N_14692,N_10251);
nand U15758 (N_15758,N_10198,N_11951);
xnor U15759 (N_15759,N_13527,N_12112);
and U15760 (N_15760,N_11885,N_13865);
nor U15761 (N_15761,N_11728,N_10860);
and U15762 (N_15762,N_13363,N_13284);
nand U15763 (N_15763,N_12779,N_13848);
xnor U15764 (N_15764,N_13311,N_12984);
xor U15765 (N_15765,N_11772,N_14733);
nor U15766 (N_15766,N_12632,N_13368);
and U15767 (N_15767,N_13651,N_13048);
xor U15768 (N_15768,N_11556,N_13602);
nand U15769 (N_15769,N_12735,N_10233);
nand U15770 (N_15770,N_10559,N_13644);
nor U15771 (N_15771,N_13698,N_11583);
and U15772 (N_15772,N_13524,N_13474);
or U15773 (N_15773,N_11421,N_13933);
or U15774 (N_15774,N_10564,N_10903);
xnor U15775 (N_15775,N_12212,N_10954);
nand U15776 (N_15776,N_14325,N_13737);
and U15777 (N_15777,N_10230,N_13006);
and U15778 (N_15778,N_10835,N_14721);
and U15779 (N_15779,N_12082,N_13794);
xnor U15780 (N_15780,N_13874,N_10697);
or U15781 (N_15781,N_12604,N_10818);
nor U15782 (N_15782,N_11030,N_12816);
or U15783 (N_15783,N_12808,N_13561);
and U15784 (N_15784,N_12860,N_14067);
nor U15785 (N_15785,N_13374,N_13096);
and U15786 (N_15786,N_12687,N_14626);
xnor U15787 (N_15787,N_11037,N_13941);
nand U15788 (N_15788,N_10969,N_12680);
and U15789 (N_15789,N_11455,N_12809);
nand U15790 (N_15790,N_11310,N_12479);
xor U15791 (N_15791,N_11328,N_10599);
and U15792 (N_15792,N_11162,N_13140);
xor U15793 (N_15793,N_11827,N_10372);
nor U15794 (N_15794,N_11024,N_10617);
nor U15795 (N_15795,N_10920,N_10280);
xor U15796 (N_15796,N_13892,N_12968);
xnor U15797 (N_15797,N_10069,N_13511);
or U15798 (N_15798,N_10812,N_11956);
nor U15799 (N_15799,N_14828,N_14673);
xor U15800 (N_15800,N_10545,N_10935);
or U15801 (N_15801,N_14045,N_14475);
or U15802 (N_15802,N_12192,N_12092);
nor U15803 (N_15803,N_11285,N_13069);
and U15804 (N_15804,N_11202,N_14770);
nand U15805 (N_15805,N_11665,N_12067);
or U15806 (N_15806,N_10682,N_11722);
or U15807 (N_15807,N_13564,N_10154);
or U15808 (N_15808,N_12711,N_13218);
or U15809 (N_15809,N_11590,N_12582);
nor U15810 (N_15810,N_12434,N_11038);
nor U15811 (N_15811,N_11447,N_13333);
nor U15812 (N_15812,N_12952,N_14272);
nand U15813 (N_15813,N_13078,N_12464);
or U15814 (N_15814,N_12596,N_13603);
and U15815 (N_15815,N_13423,N_10637);
nand U15816 (N_15816,N_11300,N_12003);
nor U15817 (N_15817,N_12246,N_13418);
nand U15818 (N_15818,N_12520,N_13824);
and U15819 (N_15819,N_14125,N_14134);
nand U15820 (N_15820,N_11240,N_10075);
and U15821 (N_15821,N_10761,N_12922);
nand U15822 (N_15822,N_14219,N_14587);
nor U15823 (N_15823,N_11370,N_14117);
nor U15824 (N_15824,N_14948,N_10579);
nor U15825 (N_15825,N_13383,N_10457);
nand U15826 (N_15826,N_12042,N_12282);
and U15827 (N_15827,N_14682,N_14069);
nor U15828 (N_15828,N_13716,N_14426);
xnor U15829 (N_15829,N_10660,N_12070);
xor U15830 (N_15830,N_10266,N_11491);
nor U15831 (N_15831,N_12958,N_14571);
xnor U15832 (N_15832,N_10145,N_10239);
xnor U15833 (N_15833,N_12463,N_12951);
or U15834 (N_15834,N_11888,N_11022);
nor U15835 (N_15835,N_12678,N_14912);
nand U15836 (N_15836,N_10187,N_12795);
xor U15837 (N_15837,N_12674,N_10254);
nand U15838 (N_15838,N_11634,N_13507);
nor U15839 (N_15839,N_12344,N_14751);
nand U15840 (N_15840,N_11074,N_10661);
xnor U15841 (N_15841,N_13247,N_14701);
and U15842 (N_15842,N_12341,N_13846);
or U15843 (N_15843,N_11605,N_11955);
or U15844 (N_15844,N_11045,N_13728);
xnor U15845 (N_15845,N_11266,N_14624);
xnor U15846 (N_15846,N_12803,N_12049);
or U15847 (N_15847,N_14909,N_14028);
or U15848 (N_15848,N_11386,N_11545);
nand U15849 (N_15849,N_11782,N_11837);
or U15850 (N_15850,N_12089,N_12211);
xor U15851 (N_15851,N_14855,N_13013);
and U15852 (N_15852,N_11477,N_13315);
nor U15853 (N_15853,N_14343,N_12481);
xor U15854 (N_15854,N_14149,N_14786);
nor U15855 (N_15855,N_11204,N_12024);
xor U15856 (N_15856,N_11295,N_12938);
or U15857 (N_15857,N_13608,N_10278);
or U15858 (N_15858,N_12996,N_10733);
xor U15859 (N_15859,N_12940,N_10554);
and U15860 (N_15860,N_11807,N_10042);
or U15861 (N_15861,N_10638,N_12602);
nor U15862 (N_15862,N_10227,N_13975);
nand U15863 (N_15863,N_11383,N_10467);
nand U15864 (N_15864,N_10830,N_13969);
xor U15865 (N_15865,N_12466,N_14206);
nand U15866 (N_15866,N_11246,N_13898);
xor U15867 (N_15867,N_13377,N_14310);
and U15868 (N_15868,N_13160,N_13154);
and U15869 (N_15869,N_10653,N_11412);
and U15870 (N_15870,N_13328,N_10139);
nand U15871 (N_15871,N_11378,N_13090);
xor U15872 (N_15872,N_10240,N_11326);
and U15873 (N_15873,N_14794,N_13588);
or U15874 (N_15874,N_11461,N_13299);
nor U15875 (N_15875,N_11280,N_12535);
xnor U15876 (N_15876,N_13532,N_10745);
nor U15877 (N_15877,N_12705,N_14200);
nor U15878 (N_15878,N_10979,N_11180);
or U15879 (N_15879,N_13587,N_14671);
nand U15880 (N_15880,N_11103,N_11726);
xor U15881 (N_15881,N_10837,N_10862);
and U15882 (N_15882,N_10602,N_14000);
or U15883 (N_15883,N_11221,N_12010);
and U15884 (N_15884,N_12845,N_10510);
nand U15885 (N_15885,N_13460,N_14204);
nor U15886 (N_15886,N_10780,N_13814);
xor U15887 (N_15887,N_13341,N_14888);
and U15888 (N_15888,N_13410,N_13638);
and U15889 (N_15889,N_13228,N_10375);
nor U15890 (N_15890,N_12719,N_11019);
nor U15891 (N_15891,N_13142,N_12060);
nand U15892 (N_15892,N_13791,N_12868);
and U15893 (N_15893,N_12223,N_10625);
and U15894 (N_15894,N_11530,N_11978);
and U15895 (N_15895,N_12537,N_11222);
xor U15896 (N_15896,N_13534,N_12046);
nand U15897 (N_15897,N_11481,N_13134);
or U15898 (N_15898,N_13958,N_14118);
and U15899 (N_15899,N_10507,N_14922);
nand U15900 (N_15900,N_14332,N_11490);
or U15901 (N_15901,N_14998,N_12353);
nor U15902 (N_15902,N_13468,N_12599);
or U15903 (N_15903,N_13693,N_12369);
or U15904 (N_15904,N_12580,N_10414);
nor U15905 (N_15905,N_13876,N_12458);
xor U15906 (N_15906,N_12913,N_12187);
and U15907 (N_15907,N_14389,N_14322);
nor U15908 (N_15908,N_12521,N_12792);
and U15909 (N_15909,N_11085,N_10933);
and U15910 (N_15910,N_11669,N_12357);
nor U15911 (N_15911,N_13127,N_14282);
xnor U15912 (N_15912,N_11997,N_10590);
and U15913 (N_15913,N_14405,N_12113);
nor U15914 (N_15914,N_14781,N_10895);
or U15915 (N_15915,N_14820,N_13397);
xor U15916 (N_15916,N_10379,N_10454);
nand U15917 (N_15917,N_12401,N_14892);
and U15918 (N_15918,N_12963,N_14053);
nand U15919 (N_15919,N_14040,N_12150);
or U15920 (N_15920,N_13109,N_11879);
nand U15921 (N_15921,N_11120,N_12992);
xor U15922 (N_15922,N_13466,N_14091);
or U15923 (N_15923,N_14316,N_10942);
nor U15924 (N_15924,N_13643,N_12159);
and U15925 (N_15925,N_13011,N_13322);
nor U15926 (N_15926,N_11065,N_12442);
nand U15927 (N_15927,N_10009,N_13495);
and U15928 (N_15928,N_12804,N_13089);
nand U15929 (N_15929,N_14900,N_13073);
or U15930 (N_15930,N_12849,N_11391);
nand U15931 (N_15931,N_12057,N_12713);
nor U15932 (N_15932,N_11119,N_13186);
nand U15933 (N_15933,N_13364,N_12764);
or U15934 (N_15934,N_12506,N_13448);
xor U15935 (N_15935,N_11581,N_12879);
xnor U15936 (N_15936,N_14725,N_14573);
or U15937 (N_15937,N_10393,N_11941);
nor U15938 (N_15938,N_13227,N_13765);
nand U15939 (N_15939,N_10252,N_12218);
nor U15940 (N_15940,N_10738,N_10121);
nor U15941 (N_15941,N_11357,N_10670);
or U15942 (N_15942,N_10867,N_10898);
xor U15943 (N_15943,N_13302,N_14056);
nor U15944 (N_15944,N_11718,N_12084);
and U15945 (N_15945,N_13822,N_11179);
or U15946 (N_15946,N_12400,N_13018);
and U15947 (N_15947,N_12589,N_12285);
nor U15948 (N_15948,N_12718,N_13756);
nand U15949 (N_15949,N_11935,N_14534);
nand U15950 (N_15950,N_12855,N_13817);
nor U15951 (N_15951,N_13552,N_13935);
nor U15952 (N_15952,N_10427,N_10991);
and U15953 (N_15953,N_10547,N_13202);
nand U15954 (N_15954,N_13235,N_13786);
and U15955 (N_15955,N_12663,N_13435);
and U15956 (N_15956,N_13110,N_13882);
xor U15957 (N_15957,N_13802,N_13612);
nor U15958 (N_15958,N_10401,N_10447);
nand U15959 (N_15959,N_14104,N_14100);
or U15960 (N_15960,N_10612,N_11615);
nand U15961 (N_15961,N_13887,N_10012);
nand U15962 (N_15962,N_12313,N_10584);
or U15963 (N_15963,N_10392,N_14940);
or U15964 (N_15964,N_12202,N_12542);
nor U15965 (N_15965,N_10465,N_10897);
xor U15966 (N_15966,N_13607,N_10403);
nor U15967 (N_15967,N_12078,N_10353);
or U15968 (N_15968,N_14470,N_10615);
nand U15969 (N_15969,N_11872,N_11994);
nand U15970 (N_15970,N_13487,N_10212);
nor U15971 (N_15971,N_11875,N_10190);
xnor U15972 (N_15972,N_13040,N_10982);
or U15973 (N_15973,N_11979,N_14980);
nand U15974 (N_15974,N_14029,N_14337);
nor U15975 (N_15975,N_10006,N_13812);
nor U15976 (N_15976,N_12497,N_14220);
nor U15977 (N_15977,N_13181,N_13691);
nand U15978 (N_15978,N_14545,N_12891);
or U15979 (N_15979,N_10043,N_11419);
xor U15980 (N_15980,N_12622,N_13384);
nor U15981 (N_15981,N_13022,N_12961);
nor U15982 (N_15982,N_12935,N_14535);
nand U15983 (N_15983,N_11660,N_11578);
and U15984 (N_15984,N_12138,N_10357);
nand U15985 (N_15985,N_13193,N_11335);
xnor U15986 (N_15986,N_10466,N_10264);
and U15987 (N_15987,N_10904,N_11972);
or U15988 (N_15988,N_12332,N_12650);
nand U15989 (N_15989,N_13003,N_12974);
or U15990 (N_15990,N_11200,N_13454);
and U15991 (N_15991,N_13336,N_12483);
xnor U15992 (N_15992,N_14779,N_14541);
or U15993 (N_15993,N_11254,N_12404);
or U15994 (N_15994,N_14113,N_13804);
or U15995 (N_15995,N_12742,N_13838);
and U15996 (N_15996,N_10841,N_14215);
or U15997 (N_15997,N_14146,N_10220);
or U15998 (N_15998,N_12242,N_14607);
or U15999 (N_15999,N_13994,N_12943);
xnor U16000 (N_16000,N_14554,N_13201);
or U16001 (N_16001,N_13767,N_11224);
xnor U16002 (N_16002,N_11528,N_10256);
nand U16003 (N_16003,N_11697,N_10316);
xnor U16004 (N_16004,N_12245,N_11167);
xnor U16005 (N_16005,N_13479,N_11212);
xnor U16006 (N_16006,N_10386,N_14810);
xor U16007 (N_16007,N_12151,N_10086);
and U16008 (N_16008,N_13019,N_12162);
and U16009 (N_16009,N_12292,N_12555);
nand U16010 (N_16010,N_10560,N_12335);
nor U16011 (N_16011,N_12287,N_10687);
or U16012 (N_16012,N_14408,N_10536);
nor U16013 (N_16013,N_12448,N_12950);
xor U16014 (N_16014,N_13847,N_13136);
nor U16015 (N_16015,N_13088,N_11762);
and U16016 (N_16016,N_13357,N_14762);
or U16017 (N_16017,N_13634,N_14851);
or U16018 (N_16018,N_12559,N_13486);
or U16019 (N_16019,N_12105,N_10757);
nand U16020 (N_16020,N_13473,N_14717);
and U16021 (N_16021,N_12759,N_10219);
nand U16022 (N_16022,N_10952,N_14614);
xor U16023 (N_16023,N_11029,N_11673);
and U16024 (N_16024,N_13647,N_10846);
or U16025 (N_16025,N_13810,N_13929);
nand U16026 (N_16026,N_13030,N_13829);
nand U16027 (N_16027,N_13963,N_11563);
and U16028 (N_16028,N_11540,N_14057);
xor U16029 (N_16029,N_12354,N_13736);
or U16030 (N_16030,N_11893,N_13176);
nor U16031 (N_16031,N_10265,N_12574);
xor U16032 (N_16032,N_13470,N_10681);
xnor U16033 (N_16033,N_11584,N_13233);
and U16034 (N_16034,N_12975,N_13528);
nor U16035 (N_16035,N_14240,N_11864);
xor U16036 (N_16036,N_11967,N_13730);
or U16037 (N_16037,N_13979,N_13880);
nor U16038 (N_16038,N_11520,N_14996);
or U16039 (N_16039,N_14989,N_11233);
or U16040 (N_16040,N_11225,N_14011);
nor U16041 (N_16041,N_10763,N_11641);
or U16042 (N_16042,N_13007,N_10613);
xnor U16043 (N_16043,N_10683,N_14008);
and U16044 (N_16044,N_13863,N_10570);
and U16045 (N_16045,N_14372,N_12528);
xor U16046 (N_16046,N_11076,N_10031);
nand U16047 (N_16047,N_14502,N_12881);
nand U16048 (N_16048,N_11808,N_13646);
nor U16049 (N_16049,N_10677,N_14648);
and U16050 (N_16050,N_11555,N_14634);
xor U16051 (N_16051,N_11562,N_13519);
nor U16052 (N_16052,N_10633,N_14093);
xnor U16053 (N_16053,N_11968,N_10434);
nand U16054 (N_16054,N_11509,N_12681);
xor U16055 (N_16055,N_11983,N_10474);
nand U16056 (N_16056,N_10623,N_10143);
nand U16057 (N_16057,N_13139,N_14221);
and U16058 (N_16058,N_12553,N_11736);
and U16059 (N_16059,N_14211,N_14755);
nor U16060 (N_16060,N_10575,N_13920);
nand U16061 (N_16061,N_12237,N_11805);
and U16062 (N_16062,N_11199,N_14928);
and U16063 (N_16063,N_11016,N_12214);
xor U16064 (N_16064,N_14101,N_14604);
nand U16065 (N_16065,N_10934,N_12424);
nand U16066 (N_16066,N_13478,N_11769);
nor U16067 (N_16067,N_10480,N_12104);
nor U16068 (N_16068,N_10050,N_11154);
nand U16069 (N_16069,N_14865,N_14946);
or U16070 (N_16070,N_12152,N_14537);
and U16071 (N_16071,N_10134,N_10845);
nor U16072 (N_16072,N_14697,N_11775);
or U16073 (N_16073,N_13051,N_14016);
nor U16074 (N_16074,N_13601,N_11114);
or U16075 (N_16075,N_14328,N_10764);
nor U16076 (N_16076,N_11650,N_10636);
nand U16077 (N_16077,N_11159,N_10640);
nand U16078 (N_16078,N_12144,N_14661);
nand U16079 (N_16079,N_12100,N_11834);
xnor U16080 (N_16080,N_13658,N_11681);
or U16081 (N_16081,N_10616,N_12561);
nor U16082 (N_16082,N_12293,N_14879);
or U16083 (N_16083,N_10762,N_14955);
and U16084 (N_16084,N_14861,N_12927);
or U16085 (N_16085,N_11902,N_12061);
nand U16086 (N_16086,N_12731,N_12048);
xor U16087 (N_16087,N_12254,N_11181);
nor U16088 (N_16088,N_12407,N_10996);
nor U16089 (N_16089,N_13025,N_10989);
xor U16090 (N_16090,N_14279,N_10255);
nor U16091 (N_16091,N_10364,N_12756);
nand U16092 (N_16092,N_13707,N_13877);
nor U16093 (N_16093,N_11288,N_14910);
or U16094 (N_16094,N_10742,N_13434);
nand U16095 (N_16095,N_10010,N_11064);
or U16096 (N_16096,N_10277,N_14652);
xnor U16097 (N_16097,N_10947,N_10350);
xnor U16098 (N_16098,N_14606,N_11770);
xor U16099 (N_16099,N_10077,N_11844);
nor U16100 (N_16100,N_12454,N_12945);
or U16101 (N_16101,N_11797,N_13594);
and U16102 (N_16102,N_12227,N_14094);
and U16103 (N_16103,N_11868,N_14789);
nor U16104 (N_16104,N_12469,N_13242);
nand U16105 (N_16105,N_11318,N_10600);
nor U16106 (N_16106,N_10360,N_11018);
nand U16107 (N_16107,N_10367,N_10497);
nor U16108 (N_16108,N_14618,N_10317);
nor U16109 (N_16109,N_12916,N_12660);
or U16110 (N_16110,N_14977,N_10083);
nor U16111 (N_16111,N_10702,N_11017);
xor U16112 (N_16112,N_13583,N_13321);
nor U16113 (N_16113,N_14559,N_10245);
and U16114 (N_16114,N_14990,N_11852);
and U16115 (N_16115,N_14033,N_14202);
nor U16116 (N_16116,N_12754,N_14886);
and U16117 (N_16117,N_11908,N_11228);
and U16118 (N_16118,N_14631,N_14473);
or U16119 (N_16119,N_11564,N_11213);
xnor U16120 (N_16120,N_13087,N_12426);
and U16121 (N_16121,N_14474,N_11433);
xor U16122 (N_16122,N_11734,N_10249);
nor U16123 (N_16123,N_14803,N_10319);
and U16124 (N_16124,N_13773,N_13086);
nor U16125 (N_16125,N_14860,N_14152);
or U16126 (N_16126,N_12098,N_14712);
nand U16127 (N_16127,N_12437,N_12957);
or U16128 (N_16128,N_10611,N_13889);
nand U16129 (N_16129,N_14747,N_12846);
and U16130 (N_16130,N_14813,N_14950);
xnor U16131 (N_16131,N_10908,N_11241);
nor U16132 (N_16132,N_12620,N_11245);
nor U16133 (N_16133,N_13557,N_14976);
xnor U16134 (N_16134,N_11186,N_10470);
nand U16135 (N_16135,N_11838,N_11296);
nand U16136 (N_16136,N_12173,N_11629);
nor U16137 (N_16137,N_14647,N_10034);
xor U16138 (N_16138,N_10594,N_10851);
and U16139 (N_16139,N_10234,N_14623);
nor U16140 (N_16140,N_10482,N_14452);
nor U16141 (N_16141,N_14507,N_13626);
or U16142 (N_16142,N_13806,N_11613);
and U16143 (N_16143,N_14116,N_13266);
nor U16144 (N_16144,N_12436,N_13530);
or U16145 (N_16145,N_13554,N_12822);
or U16146 (N_16146,N_10936,N_14155);
nor U16147 (N_16147,N_11143,N_11505);
nor U16148 (N_16148,N_11603,N_10549);
or U16149 (N_16149,N_11702,N_11819);
nand U16150 (N_16150,N_11643,N_14111);
nand U16151 (N_16151,N_14758,N_10426);
nor U16152 (N_16152,N_13758,N_14388);
or U16153 (N_16153,N_14783,N_13605);
xor U16154 (N_16154,N_12767,N_14504);
or U16155 (N_16155,N_13338,N_11846);
xor U16156 (N_16156,N_14987,N_13900);
nand U16157 (N_16157,N_11511,N_14468);
or U16158 (N_16158,N_10542,N_14014);
and U16159 (N_16159,N_10722,N_13399);
nand U16160 (N_16160,N_10442,N_12263);
and U16161 (N_16161,N_13147,N_11740);
nor U16162 (N_16162,N_10957,N_13619);
or U16163 (N_16163,N_14752,N_10131);
nor U16164 (N_16164,N_11970,N_10179);
xnor U16165 (N_16165,N_14638,N_11164);
or U16166 (N_16166,N_14449,N_11793);
nor U16167 (N_16167,N_12329,N_10404);
xor U16168 (N_16168,N_11373,N_11073);
nor U16169 (N_16169,N_13339,N_10362);
nand U16170 (N_16170,N_10369,N_11067);
and U16171 (N_16171,N_10844,N_12591);
and U16172 (N_16172,N_12423,N_12692);
nand U16173 (N_16173,N_11798,N_10164);
nor U16174 (N_16174,N_13684,N_11507);
or U16175 (N_16175,N_10876,N_10603);
nand U16176 (N_16176,N_10551,N_11430);
and U16177 (N_16177,N_11498,N_10968);
or U16178 (N_16178,N_10866,N_14249);
xnor U16179 (N_16179,N_10951,N_14660);
and U16180 (N_16180,N_14722,N_12396);
nand U16181 (N_16181,N_10842,N_12886);
nand U16182 (N_16182,N_11656,N_14743);
nand U16183 (N_16183,N_13774,N_10701);
xnor U16184 (N_16184,N_11614,N_13196);
nand U16185 (N_16185,N_11948,N_11678);
xor U16186 (N_16186,N_10052,N_11903);
nor U16187 (N_16187,N_12478,N_12575);
xor U16188 (N_16188,N_12179,N_11690);
or U16189 (N_16189,N_10992,N_13401);
xor U16190 (N_16190,N_12307,N_14536);
and U16191 (N_16191,N_12008,N_14451);
or U16192 (N_16192,N_10413,N_14514);
xor U16193 (N_16193,N_10243,N_10487);
and U16194 (N_16194,N_11646,N_13659);
xnor U16195 (N_16195,N_10840,N_13282);
and U16196 (N_16196,N_14018,N_13763);
nor U16197 (N_16197,N_14769,N_11226);
or U16198 (N_16198,N_14306,N_11238);
and U16199 (N_16199,N_11806,N_11833);
nor U16200 (N_16200,N_10854,N_14441);
or U16201 (N_16201,N_12471,N_10089);
nor U16202 (N_16202,N_11289,N_13922);
xnor U16203 (N_16203,N_12197,N_10823);
nand U16204 (N_16204,N_14600,N_12320);
or U16205 (N_16205,N_14330,N_13672);
nor U16206 (N_16206,N_12587,N_13562);
nand U16207 (N_16207,N_13066,N_11533);
or U16208 (N_16208,N_14941,N_11313);
and U16209 (N_16209,N_11651,N_13989);
nor U16210 (N_16210,N_11253,N_14678);
nor U16211 (N_16211,N_14498,N_13516);
or U16212 (N_16212,N_13907,N_12840);
or U16213 (N_16213,N_13038,N_11784);
and U16214 (N_16214,N_14403,N_12229);
and U16215 (N_16215,N_14518,N_10285);
nor U16216 (N_16216,N_12023,N_12252);
and U16217 (N_16217,N_14037,N_12964);
xnor U16218 (N_16218,N_11572,N_13422);
nor U16219 (N_16219,N_11708,N_14561);
nor U16220 (N_16220,N_11464,N_14656);
xor U16221 (N_16221,N_14157,N_10402);
and U16222 (N_16222,N_10253,N_10826);
or U16223 (N_16223,N_10717,N_13703);
xnor U16224 (N_16224,N_12821,N_11407);
and U16225 (N_16225,N_12983,N_14166);
and U16226 (N_16226,N_13335,N_14177);
nor U16227 (N_16227,N_11707,N_11004);
and U16228 (N_16228,N_11055,N_13740);
or U16229 (N_16229,N_14538,N_10631);
or U16230 (N_16230,N_12253,N_12149);
nand U16231 (N_16231,N_11645,N_12413);
xor U16232 (N_16232,N_12631,N_13582);
or U16233 (N_16233,N_12233,N_12960);
and U16234 (N_16234,N_13476,N_12249);
or U16235 (N_16235,N_11134,N_11855);
and U16236 (N_16236,N_13180,N_13330);
nand U16237 (N_16237,N_12177,N_14311);
or U16238 (N_16238,N_10237,N_12826);
nor U16239 (N_16239,N_13031,N_12308);
xnor U16240 (N_16240,N_13165,N_14471);
nand U16241 (N_16241,N_12639,N_12398);
nor U16242 (N_16242,N_12568,N_13940);
nor U16243 (N_16243,N_13591,N_12969);
xnor U16244 (N_16244,N_11560,N_14602);
nand U16245 (N_16245,N_11521,N_13662);
nor U16246 (N_16246,N_10917,N_11072);
or U16247 (N_16247,N_12130,N_10335);
nor U16248 (N_16248,N_12863,N_11013);
or U16249 (N_16249,N_11489,N_14877);
or U16250 (N_16250,N_10806,N_12928);
nor U16251 (N_16251,N_13151,N_11005);
nor U16252 (N_16252,N_12294,N_13867);
nand U16253 (N_16253,N_12358,N_12811);
or U16254 (N_16254,N_14641,N_13565);
or U16255 (N_16255,N_13717,N_11001);
xor U16256 (N_16256,N_13433,N_14414);
xor U16257 (N_16257,N_12017,N_14757);
nand U16258 (N_16258,N_11504,N_12503);
nand U16259 (N_16259,N_13923,N_13424);
and U16260 (N_16260,N_13430,N_10257);
nor U16261 (N_16261,N_14558,N_11075);
or U16262 (N_16262,N_13972,N_12445);
xnor U16263 (N_16263,N_11780,N_14837);
and U16264 (N_16264,N_12451,N_12475);
nor U16265 (N_16265,N_10074,N_11642);
or U16266 (N_16266,N_10975,N_14519);
or U16267 (N_16267,N_10338,N_10896);
nor U16268 (N_16268,N_13198,N_11767);
nand U16269 (N_16269,N_11688,N_10498);
or U16270 (N_16270,N_11900,N_11953);
or U16271 (N_16271,N_14022,N_12798);
nor U16272 (N_16272,N_10949,N_14382);
nand U16273 (N_16273,N_11069,N_11284);
nor U16274 (N_16274,N_10411,N_11881);
and U16275 (N_16275,N_10153,N_14186);
nand U16276 (N_16276,N_13575,N_13574);
and U16277 (N_16277,N_11604,N_13108);
or U16278 (N_16278,N_12068,N_13396);
or U16279 (N_16279,N_11608,N_10366);
nor U16280 (N_16280,N_11086,N_12161);
nand U16281 (N_16281,N_11428,N_12324);
and U16282 (N_16282,N_14071,N_11422);
xor U16283 (N_16283,N_10365,N_14893);
nand U16284 (N_16284,N_10735,N_14804);
nand U16285 (N_16285,N_13351,N_11156);
xnor U16286 (N_16286,N_11539,N_13797);
and U16287 (N_16287,N_13949,N_14771);
xnor U16288 (N_16288,N_13978,N_14639);
or U16289 (N_16289,N_12655,N_11963);
and U16290 (N_16290,N_11851,N_10974);
and U16291 (N_16291,N_12848,N_10808);
nand U16292 (N_16292,N_13182,N_12477);
and U16293 (N_16293,N_14608,N_12552);
nand U16294 (N_16294,N_11756,N_13221);
nor U16295 (N_16295,N_13568,N_10782);
nand U16296 (N_16296,N_13403,N_10809);
or U16297 (N_16297,N_12304,N_10517);
xnor U16298 (N_16298,N_14404,N_14801);
xor U16299 (N_16299,N_10383,N_14588);
and U16300 (N_16300,N_10018,N_14657);
or U16301 (N_16301,N_12487,N_13152);
nor U16302 (N_16302,N_12876,N_14821);
or U16303 (N_16303,N_11438,N_10927);
nor U16304 (N_16304,N_13749,N_14792);
nand U16305 (N_16305,N_11317,N_11008);
and U16306 (N_16306,N_12955,N_14793);
xor U16307 (N_16307,N_14570,N_13886);
and U16308 (N_16308,N_11223,N_11137);
nor U16309 (N_16309,N_12170,N_10943);
and U16310 (N_16310,N_10739,N_12508);
or U16311 (N_16311,N_12704,N_10218);
nor U16312 (N_16312,N_14897,N_13723);
xnor U16313 (N_16313,N_10801,N_13653);
and U16314 (N_16314,N_10099,N_11000);
xor U16315 (N_16315,N_10672,N_13712);
nor U16316 (N_16316,N_13873,N_12865);
or U16317 (N_16317,N_12989,N_13445);
or U16318 (N_16318,N_13946,N_10568);
xnor U16319 (N_16319,N_12544,N_10477);
or U16320 (N_16320,N_14651,N_11068);
xor U16321 (N_16321,N_12904,N_13705);
nand U16322 (N_16322,N_13332,N_10561);
nor U16323 (N_16323,N_14144,N_12770);
and U16324 (N_16324,N_11675,N_10775);
and U16325 (N_16325,N_10258,N_13373);
or U16326 (N_16326,N_10119,N_13714);
nor U16327 (N_16327,N_10475,N_14076);
xor U16328 (N_16328,N_11431,N_10017);
nand U16329 (N_16329,N_13103,N_10713);
xnor U16330 (N_16330,N_10861,N_11286);
or U16331 (N_16331,N_12347,N_12427);
xor U16332 (N_16332,N_11922,N_10675);
and U16333 (N_16333,N_12213,N_14245);
xor U16334 (N_16334,N_13677,N_14875);
or U16335 (N_16335,N_12385,N_10296);
or U16336 (N_16336,N_14260,N_10359);
and U16337 (N_16337,N_11940,N_11884);
or U16338 (N_16338,N_12207,N_11056);
and U16339 (N_16339,N_13988,N_11828);
or U16340 (N_16340,N_10327,N_11347);
and U16341 (N_16341,N_14109,N_12751);
nor U16342 (N_16342,N_11976,N_12280);
or U16343 (N_16343,N_14944,N_10246);
xor U16344 (N_16344,N_13595,N_13058);
nand U16345 (N_16345,N_11332,N_10650);
nor U16346 (N_16346,N_10629,N_14662);
xor U16347 (N_16347,N_13037,N_12897);
nand U16348 (N_16348,N_12588,N_13252);
and U16349 (N_16349,N_12117,N_11339);
or U16350 (N_16350,N_11057,N_14323);
and U16351 (N_16351,N_13185,N_10388);
nor U16352 (N_16352,N_12278,N_14226);
nor U16353 (N_16353,N_13609,N_14397);
and U16354 (N_16354,N_10891,N_12031);
nand U16355 (N_16355,N_14622,N_10597);
or U16356 (N_16356,N_14095,N_10054);
nor U16357 (N_16357,N_12787,N_14464);
nor U16358 (N_16358,N_12738,N_14235);
nand U16359 (N_16359,N_10368,N_14965);
nor U16360 (N_16360,N_12217,N_13360);
or U16361 (N_16361,N_11003,N_10015);
and U16362 (N_16362,N_11042,N_10743);
and U16363 (N_16363,N_10710,N_10214);
xnor U16364 (N_16364,N_11175,N_12775);
and U16365 (N_16365,N_13246,N_11910);
xor U16366 (N_16366,N_13138,N_12493);
and U16367 (N_16367,N_12601,N_11355);
and U16368 (N_16368,N_10269,N_13021);
or U16369 (N_16369,N_11738,N_10546);
nor U16370 (N_16370,N_10449,N_10244);
nor U16371 (N_16371,N_12473,N_10601);
xnor U16372 (N_16372,N_11369,N_13673);
xnor U16373 (N_16373,N_12410,N_10971);
and U16374 (N_16374,N_12452,N_13656);
xnor U16375 (N_16375,N_14842,N_13124);
and U16376 (N_16376,N_14455,N_13257);
nor U16377 (N_16377,N_14702,N_10937);
or U16378 (N_16378,N_12239,N_13539);
and U16379 (N_16379,N_12210,N_10380);
nor U16380 (N_16380,N_11870,N_10342);
and U16381 (N_16381,N_14741,N_10911);
or U16382 (N_16382,N_13337,N_10905);
and U16383 (N_16383,N_10847,N_14025);
nand U16384 (N_16384,N_10609,N_13982);
or U16385 (N_16385,N_12260,N_10700);
or U16386 (N_16386,N_12797,N_13113);
or U16387 (N_16387,N_12295,N_14463);
and U16388 (N_16388,N_12364,N_11100);
xnor U16389 (N_16389,N_10825,N_11135);
nor U16390 (N_16390,N_14728,N_14951);
xnor U16391 (N_16391,N_10756,N_11263);
nor U16392 (N_16392,N_14072,N_13811);
and U16393 (N_16393,N_14114,N_12203);
or U16394 (N_16394,N_14744,N_13820);
or U16395 (N_16395,N_13054,N_14012);
and U16396 (N_16396,N_14002,N_13680);
xnor U16397 (N_16397,N_12571,N_13803);
nor U16398 (N_16398,N_14001,N_14669);
or U16399 (N_16399,N_14459,N_11831);
or U16400 (N_16400,N_10071,N_12956);
xnor U16401 (N_16401,N_10759,N_11470);
nor U16402 (N_16402,N_12755,N_13100);
or U16403 (N_16403,N_10222,N_13406);
or U16404 (N_16404,N_12000,N_11930);
or U16405 (N_16405,N_14248,N_14674);
nand U16406 (N_16406,N_14477,N_12505);
nor U16407 (N_16407,N_13780,N_12101);
and U16408 (N_16408,N_12221,N_10726);
or U16409 (N_16409,N_10963,N_14716);
xnor U16410 (N_16410,N_10063,N_14834);
nand U16411 (N_16411,N_10544,N_12854);
and U16412 (N_16412,N_14934,N_14878);
xnor U16413 (N_16413,N_12238,N_11338);
nor U16414 (N_16414,N_10541,N_11795);
xor U16415 (N_16415,N_14437,N_12414);
or U16416 (N_16416,N_12036,N_12039);
nor U16417 (N_16417,N_10798,N_14481);
xor U16418 (N_16418,N_10163,N_11639);
or U16419 (N_16419,N_11007,N_10524);
nor U16420 (N_16420,N_10945,N_14655);
xor U16421 (N_16421,N_10344,N_14431);
nand U16422 (N_16422,N_12656,N_14968);
nand U16423 (N_16423,N_12939,N_11532);
nand U16424 (N_16424,N_14864,N_14732);
xor U16425 (N_16425,N_10128,N_12172);
nor U16426 (N_16426,N_13382,N_10725);
and U16427 (N_16427,N_10651,N_14190);
xnor U16428 (N_16428,N_13839,N_14528);
nor U16429 (N_16429,N_14313,N_14169);
xnor U16430 (N_16430,N_14007,N_14307);
nand U16431 (N_16431,N_14108,N_14009);
xor U16432 (N_16432,N_14991,N_12500);
nand U16433 (N_16433,N_13052,N_13411);
xor U16434 (N_16434,N_14145,N_12240);
xor U16435 (N_16435,N_11638,N_13043);
and U16436 (N_16436,N_10576,N_14139);
and U16437 (N_16437,N_14777,N_11506);
and U16438 (N_16438,N_11083,N_13657);
xor U16439 (N_16439,N_12525,N_12871);
nor U16440 (N_16440,N_13250,N_10448);
xor U16441 (N_16441,N_13746,N_13079);
nor U16442 (N_16442,N_11081,N_14255);
nor U16443 (N_16443,N_13970,N_12698);
xnor U16444 (N_16444,N_12832,N_14891);
and U16445 (N_16445,N_12736,N_14243);
and U16446 (N_16446,N_13931,N_11229);
nor U16447 (N_16447,N_13888,N_11794);
and U16448 (N_16448,N_13286,N_11699);
xor U16449 (N_16449,N_11672,N_14857);
xor U16450 (N_16450,N_12484,N_14084);
nor U16451 (N_16451,N_11826,N_10875);
nor U16452 (N_16452,N_10639,N_12675);
or U16453 (N_16453,N_11554,N_12833);
and U16454 (N_16454,N_10192,N_14236);
or U16455 (N_16455,N_10980,N_11242);
xor U16456 (N_16456,N_10939,N_13501);
or U16457 (N_16457,N_13727,N_14689);
or U16458 (N_16458,N_10170,N_10420);
and U16459 (N_16459,N_13945,N_13869);
or U16460 (N_16460,N_10439,N_11250);
nor U16461 (N_16461,N_14147,N_12350);
and U16462 (N_16462,N_13990,N_12901);
nor U16463 (N_16463,N_11676,N_14453);
nor U16464 (N_16464,N_13281,N_13285);
xnor U16465 (N_16465,N_13766,N_12370);
and U16466 (N_16466,N_12496,N_14707);
xor U16467 (N_16467,N_11196,N_12373);
xnor U16468 (N_16468,N_10421,N_10605);
and U16469 (N_16469,N_10076,N_10440);
or U16470 (N_16470,N_14444,N_12746);
and U16471 (N_16471,N_11933,N_13667);
xor U16472 (N_16472,N_11552,N_13823);
xnor U16473 (N_16473,N_10944,N_13036);
nor U16474 (N_16474,N_13855,N_14321);
nand U16475 (N_16475,N_12474,N_14238);
nor U16476 (N_16476,N_10953,N_11786);
and U16477 (N_16477,N_11450,N_11169);
nor U16478 (N_16478,N_13369,N_10446);
xor U16479 (N_16479,N_14277,N_11345);
and U16480 (N_16480,N_10724,N_10430);
and U16481 (N_16481,N_13023,N_13379);
nand U16482 (N_16482,N_12903,N_11258);
or U16483 (N_16483,N_14904,N_10097);
xnor U16484 (N_16484,N_10081,N_14062);
and U16485 (N_16485,N_14970,N_10698);
or U16486 (N_16486,N_12907,N_10674);
and U16487 (N_16487,N_12156,N_12819);
nand U16488 (N_16488,N_13854,N_12603);
and U16489 (N_16489,N_13556,N_13199);
or U16490 (N_16490,N_11304,N_10607);
xnor U16491 (N_16491,N_12852,N_11640);
nand U16492 (N_16492,N_12605,N_10312);
nand U16493 (N_16493,N_11561,N_11616);
or U16494 (N_16494,N_11546,N_13542);
xnor U16495 (N_16495,N_10553,N_11974);
nand U16496 (N_16496,N_14121,N_12094);
nand U16497 (N_16497,N_10816,N_14483);
nand U16498 (N_16498,N_14585,N_14135);
or U16499 (N_16499,N_14665,N_12682);
and U16500 (N_16500,N_11390,N_11166);
nor U16501 (N_16501,N_11626,N_13271);
xnor U16502 (N_16502,N_10476,N_10468);
xnor U16503 (N_16503,N_14213,N_14210);
or U16504 (N_16504,N_10025,N_10080);
xnor U16505 (N_16505,N_10634,N_10223);
xor U16506 (N_16506,N_14402,N_14795);
or U16507 (N_16507,N_14314,N_11356);
nor U16508 (N_16508,N_12244,N_14295);
and U16509 (N_16509,N_13491,N_14327);
nand U16510 (N_16510,N_10749,N_13906);
xor U16511 (N_16511,N_12321,N_13131);
or U16512 (N_16512,N_11298,N_13661);
xnor U16513 (N_16513,N_13754,N_11754);
nor U16514 (N_16514,N_12933,N_13393);
nand U16515 (N_16515,N_10068,N_11108);
nand U16516 (N_16516,N_10260,N_12103);
and U16517 (N_16517,N_14952,N_11742);
nor U16518 (N_16518,N_14315,N_12050);
nand U16519 (N_16519,N_12946,N_14883);
xnor U16520 (N_16520,N_10802,N_12870);
nor U16521 (N_16521,N_11101,N_11381);
nor U16522 (N_16522,N_14354,N_13631);
or U16523 (N_16523,N_10513,N_11649);
nor U16524 (N_16524,N_10105,N_14694);
nor U16525 (N_16525,N_11975,N_13843);
nand U16526 (N_16526,N_10108,N_12665);
or U16527 (N_16527,N_11365,N_13229);
or U16528 (N_16528,N_13951,N_14869);
nor U16529 (N_16529,N_11316,N_11542);
nor U16530 (N_16530,N_14693,N_12327);
and U16531 (N_16531,N_14548,N_12673);
nor U16532 (N_16532,N_12310,N_10241);
and U16533 (N_16533,N_12847,N_13968);
and U16534 (N_16534,N_14522,N_11523);
nand U16535 (N_16535,N_12345,N_14427);
nand U16536 (N_16536,N_13482,N_10236);
xnor U16537 (N_16537,N_13112,N_10865);
and U16538 (N_16538,N_13203,N_13704);
xor U16539 (N_16539,N_11348,N_12633);
and U16540 (N_16540,N_11887,N_13648);
and U16541 (N_16541,N_12606,N_13915);
and U16542 (N_16542,N_13441,N_11387);
nor U16543 (N_16543,N_13816,N_10374);
nor U16544 (N_16544,N_13291,N_12818);
nand U16545 (N_16545,N_13296,N_11760);
xnor U16546 (N_16546,N_14827,N_11567);
xnor U16547 (N_16547,N_11417,N_10055);
or U16548 (N_16548,N_11904,N_12085);
nand U16549 (N_16549,N_14338,N_10931);
nand U16550 (N_16550,N_13627,N_13146);
nor U16551 (N_16551,N_13759,N_13536);
or U16552 (N_16552,N_10503,N_11256);
and U16553 (N_16553,N_13372,N_12267);
or U16554 (N_16554,N_11059,N_12045);
or U16555 (N_16555,N_10184,N_10995);
nor U16556 (N_16556,N_11268,N_14319);
and U16557 (N_16557,N_10117,N_13417);
nor U16558 (N_16558,N_12279,N_12190);
or U16559 (N_16559,N_14870,N_14088);
or U16560 (N_16560,N_14796,N_11299);
nor U16561 (N_16561,N_13067,N_12654);
and U16562 (N_16562,N_11448,N_12359);
and U16563 (N_16563,N_10019,N_14748);
xnor U16564 (N_16564,N_13047,N_12198);
xor U16565 (N_16565,N_14817,N_10915);
or U16566 (N_16566,N_13760,N_14848);
or U16567 (N_16567,N_14425,N_12334);
xor U16568 (N_16568,N_11098,N_12815);
nand U16569 (N_16569,N_11906,N_10016);
xnor U16570 (N_16570,N_13604,N_13049);
nor U16571 (N_16571,N_11459,N_11937);
or U16572 (N_16572,N_13502,N_10494);
nor U16573 (N_16573,N_13297,N_12021);
or U16574 (N_16574,N_12942,N_11984);
and U16575 (N_16575,N_13492,N_14046);
nor U16576 (N_16576,N_12667,N_13669);
xnor U16577 (N_16577,N_14532,N_12300);
and U16578 (N_16578,N_13334,N_14933);
or U16579 (N_16579,N_10395,N_10730);
and U16580 (N_16580,N_11384,N_14039);
or U16581 (N_16581,N_11624,N_11281);
or U16582 (N_16582,N_14407,N_13750);
nand U16583 (N_16583,N_13715,N_14153);
or U16584 (N_16584,N_13387,N_12323);
and U16585 (N_16585,N_13789,N_14546);
nor U16586 (N_16586,N_14831,N_13074);
nand U16587 (N_16587,N_11877,N_12523);
nor U16588 (N_16588,N_13632,N_11531);
nand U16589 (N_16589,N_10351,N_12443);
nand U16590 (N_16590,N_12857,N_10188);
nor U16591 (N_16591,N_14916,N_14298);
and U16592 (N_16592,N_12677,N_13878);
xor U16593 (N_16593,N_11446,N_13098);
xnor U16594 (N_16594,N_13944,N_11818);
nor U16595 (N_16595,N_11411,N_11344);
or U16596 (N_16596,N_14264,N_14997);
or U16597 (N_16597,N_13026,N_12703);
xor U16598 (N_16598,N_12290,N_13489);
and U16599 (N_16599,N_13917,N_13559);
or U16600 (N_16600,N_11633,N_14698);
nand U16601 (N_16601,N_11445,N_13020);
nand U16602 (N_16602,N_12040,N_12615);
nand U16603 (N_16603,N_11277,N_12096);
or U16604 (N_16604,N_10999,N_13875);
xor U16605 (N_16605,N_12780,N_14569);
or U16606 (N_16606,N_11630,N_10581);
xnor U16607 (N_16607,N_12856,N_10781);
and U16608 (N_16608,N_12644,N_10786);
or U16609 (N_16609,N_10471,N_11508);
xor U16610 (N_16610,N_13070,N_12114);
nor U16611 (N_16611,N_14999,N_12874);
nor U16612 (N_16612,N_13443,N_11170);
nor U16613 (N_16613,N_10515,N_12219);
nor U16614 (N_16614,N_10748,N_10552);
or U16615 (N_16615,N_10346,N_11275);
and U16616 (N_16616,N_10785,N_12467);
xor U16617 (N_16617,N_14495,N_11033);
and U16618 (N_16618,N_10793,N_12033);
nor U16619 (N_16619,N_10106,N_13000);
or U16620 (N_16620,N_10478,N_10784);
nor U16621 (N_16621,N_10035,N_12934);
and U16622 (N_16622,N_13094,N_13957);
nand U16623 (N_16623,N_14491,N_14742);
nand U16624 (N_16624,N_13254,N_14087);
nand U16625 (N_16625,N_11451,N_13105);
xnor U16626 (N_16626,N_11449,N_14217);
nand U16627 (N_16627,N_11839,N_11174);
and U16628 (N_16628,N_12390,N_14120);
nor U16629 (N_16629,N_14421,N_10329);
and U16630 (N_16630,N_11380,N_14822);
xor U16631 (N_16631,N_12924,N_12206);
and U16632 (N_16632,N_12649,N_14006);
or U16633 (N_16633,N_12919,N_13413);
nor U16634 (N_16634,N_11787,N_13483);
or U16635 (N_16635,N_13995,N_14143);
nor U16636 (N_16636,N_13579,N_11435);
or U16637 (N_16637,N_12195,N_14059);
or U16638 (N_16638,N_13897,N_12539);
nor U16639 (N_16639,N_13938,N_14055);
or U16640 (N_16640,N_13159,N_10586);
xnor U16641 (N_16641,N_11796,N_10863);
xnor U16642 (N_16642,N_13427,N_13872);
or U16643 (N_16643,N_10961,N_11670);
nor U16644 (N_16644,N_14399,N_12418);
or U16645 (N_16645,N_10856,N_11880);
nor U16646 (N_16646,N_13666,N_10275);
xnor U16647 (N_16647,N_10648,N_14366);
xor U16648 (N_16648,N_13860,N_14356);
or U16649 (N_16649,N_11483,N_12887);
nor U16650 (N_16650,N_13735,N_10088);
xnor U16651 (N_16651,N_13437,N_11721);
nand U16652 (N_16652,N_11327,N_11926);
and U16653 (N_16653,N_12829,N_14344);
or U16654 (N_16654,N_14205,N_12936);
or U16655 (N_16655,N_13517,N_13053);
and U16656 (N_16656,N_13668,N_12725);
nand U16657 (N_16657,N_14445,N_13908);
nand U16658 (N_16658,N_13172,N_14048);
or U16659 (N_16659,N_12456,N_11360);
nor U16660 (N_16660,N_12037,N_14979);
or U16661 (N_16661,N_12567,N_13273);
nand U16662 (N_16662,N_13702,N_13447);
nor U16663 (N_16663,N_14317,N_13785);
and U16664 (N_16664,N_10065,N_14710);
and U16665 (N_16665,N_11850,N_12566);
xnor U16666 (N_16666,N_14064,N_12640);
nand U16667 (N_16667,N_10261,N_11918);
or U16668 (N_16668,N_14582,N_13606);
xor U16669 (N_16669,N_11771,N_12813);
and U16670 (N_16670,N_13788,N_12124);
xnor U16671 (N_16671,N_12459,N_11966);
nor U16672 (N_16672,N_14159,N_11495);
or U16673 (N_16673,N_11349,N_13997);
xnor U16674 (N_16674,N_10287,N_12750);
xor U16675 (N_16675,N_14465,N_12581);
nor U16676 (N_16676,N_12136,N_12169);
xnor U16677 (N_16677,N_13130,N_10363);
nand U16678 (N_16678,N_10712,N_11550);
nor U16679 (N_16679,N_10376,N_11829);
and U16680 (N_16680,N_14107,N_12899);
xnor U16681 (N_16681,N_12073,N_11883);
nor U16682 (N_16682,N_11090,N_13950);
or U16683 (N_16683,N_12572,N_10914);
and U16684 (N_16684,N_11010,N_11753);
xnor U16685 (N_16685,N_11925,N_13122);
nand U16686 (N_16686,N_10149,N_11206);
nor U16687 (N_16687,N_13510,N_11093);
xnor U16688 (N_16688,N_12944,N_13316);
and U16689 (N_16689,N_10412,N_11668);
or U16690 (N_16690,N_14158,N_14905);
nand U16691 (N_16691,N_10959,N_11312);
or U16692 (N_16692,N_12980,N_10303);
xor U16693 (N_16693,N_14487,N_10225);
nand U16694 (N_16694,N_12638,N_11071);
or U16695 (N_16695,N_12744,N_13918);
and U16696 (N_16696,N_11025,N_14635);
or U16697 (N_16697,N_13690,N_13106);
or U16698 (N_16698,N_11462,N_11168);
xnor U16699 (N_16699,N_13783,N_13916);
nand U16700 (N_16700,N_14472,N_14840);
and U16701 (N_16701,N_14406,N_12256);
nand U16702 (N_16702,N_10247,N_13722);
xor U16703 (N_16703,N_13071,N_12441);
nand U16704 (N_16704,N_11402,N_12785);
and U16705 (N_16705,N_10283,N_10912);
xnor U16706 (N_16706,N_13966,N_12457);
or U16707 (N_16707,N_13465,N_12166);
nor U16708 (N_16708,N_12002,N_12222);
nand U16709 (N_16709,N_10462,N_14224);
and U16710 (N_16710,N_12805,N_11047);
nor U16711 (N_16711,N_14058,N_11647);
or U16712 (N_16712,N_12110,N_13558);
nand U16713 (N_16713,N_12618,N_12837);
or U16714 (N_16714,N_13274,N_13488);
and U16715 (N_16715,N_10662,N_13781);
xor U16716 (N_16716,N_13409,N_10788);
nand U16717 (N_16717,N_14167,N_11113);
and U16718 (N_16718,N_13551,N_14484);
nor U16719 (N_16719,N_12137,N_13490);
and U16720 (N_16720,N_14738,N_12337);
nor U16721 (N_16721,N_12608,N_14266);
xnor U16722 (N_16722,N_14898,N_10591);
nand U16723 (N_16723,N_12550,N_14705);
or U16724 (N_16724,N_13277,N_13027);
and U16725 (N_16725,N_14460,N_14785);
or U16726 (N_16726,N_10008,N_10669);
xor U16727 (N_16727,N_13162,N_12825);
nor U16728 (N_16728,N_14859,N_13983);
nor U16729 (N_16729,N_10502,N_14526);
or U16730 (N_16730,N_10044,N_14494);
nor U16731 (N_16731,N_14218,N_12435);
xor U16732 (N_16732,N_12807,N_13213);
and U16733 (N_16733,N_13572,N_11813);
or U16734 (N_16734,N_11730,N_12087);
and U16735 (N_16735,N_10585,N_12356);
nand U16736 (N_16736,N_11934,N_13485);
or U16737 (N_16737,N_14467,N_11203);
and U16738 (N_16738,N_11916,N_13725);
nor U16739 (N_16739,N_11737,N_11822);
nand U16740 (N_16740,N_14035,N_12230);
or U16741 (N_16741,N_13059,N_11847);
xor U16742 (N_16742,N_12132,N_11458);
or U16743 (N_16743,N_12006,N_11592);
nand U16744 (N_16744,N_14563,N_14957);
or U16745 (N_16745,N_14972,N_14358);
xnor U16746 (N_16746,N_12688,N_14649);
xor U16747 (N_16747,N_11054,N_11178);
nand U16748 (N_16748,N_14521,N_14079);
nand U16749 (N_16749,N_13308,N_14772);
nand U16750 (N_16750,N_11716,N_12701);
and U16751 (N_16751,N_13205,N_10090);
and U16752 (N_16752,N_12086,N_10047);
and U16753 (N_16753,N_12311,N_13123);
nand U16754 (N_16754,N_14182,N_11791);
xor U16755 (N_16755,N_13358,N_10206);
nor U16756 (N_16756,N_14664,N_11176);
nand U16757 (N_16757,N_11189,N_10822);
or U16758 (N_16758,N_11705,N_11145);
nor U16759 (N_16759,N_10484,N_11112);
or U16760 (N_16760,N_11423,N_14988);
or U16761 (N_16761,N_12973,N_11964);
xnor U16762 (N_16762,N_13757,N_10492);
nand U16763 (N_16763,N_10295,N_13514);
xnor U16764 (N_16764,N_11582,N_11427);
or U16765 (N_16765,N_13459,N_10504);
xnor U16766 (N_16766,N_11911,N_13009);
and U16767 (N_16767,N_14049,N_10417);
nor U16768 (N_16768,N_13782,N_10804);
nor U16769 (N_16769,N_11367,N_12728);
nand U16770 (N_16770,N_10300,N_10666);
nand U16771 (N_16771,N_13998,N_10699);
and U16772 (N_16772,N_11840,N_13169);
and U16773 (N_16773,N_14839,N_12793);
xnor U16774 (N_16774,N_14598,N_11777);
nor U16775 (N_16775,N_12076,N_14488);
or U16776 (N_16776,N_12322,N_11587);
and U16777 (N_16777,N_12272,N_12689);
nor U16778 (N_16778,N_14423,N_13144);
and U16779 (N_16779,N_11036,N_11308);
xor U16780 (N_16780,N_10112,N_13451);
nand U16781 (N_16781,N_12298,N_14301);
xnor U16782 (N_16782,N_11571,N_10680);
and U16783 (N_16783,N_14964,N_14858);
nor U16784 (N_16784,N_13391,N_12554);
or U16785 (N_16785,N_13566,N_10910);
nand U16786 (N_16786,N_13506,N_13263);
xor U16787 (N_16787,N_12531,N_13617);
nand U16788 (N_16788,N_12482,N_14345);
and U16789 (N_16789,N_10534,N_14309);
nand U16790 (N_16790,N_13738,N_13808);
xor U16791 (N_16791,N_12556,N_10519);
or U16792 (N_16792,N_13976,N_10073);
xor U16793 (N_16793,N_12565,N_10518);
or U16794 (N_16794,N_11783,N_11928);
nor U16795 (N_16795,N_10408,N_11414);
nor U16796 (N_16796,N_14179,N_10213);
or U16797 (N_16797,N_11363,N_14503);
and U16798 (N_16798,N_14995,N_12139);
nand U16799 (N_16799,N_10095,N_14823);
nand U16800 (N_16800,N_12524,N_11437);
xor U16801 (N_16801,N_13890,N_13065);
nand U16802 (N_16802,N_12491,N_13512);
nand U16803 (N_16803,N_11078,N_10736);
or U16804 (N_16804,N_10839,N_12194);
and U16805 (N_16805,N_11234,N_10595);
nor U16806 (N_16806,N_13544,N_14168);
xnor U16807 (N_16807,N_12043,N_10337);
xor U16808 (N_16808,N_14227,N_10925);
nor U16809 (N_16809,N_13980,N_10874);
or U16810 (N_16810,N_10976,N_14363);
or U16811 (N_16811,N_11416,N_11595);
xor U16812 (N_16812,N_11136,N_13675);
or U16813 (N_16813,N_14269,N_10902);
nor U16814 (N_16814,N_12617,N_12406);
xnor U16815 (N_16815,N_13187,N_10488);
xor U16816 (N_16816,N_11410,N_14283);
and U16817 (N_16817,N_14192,N_12228);
or U16818 (N_16818,N_11710,N_10165);
xnor U16819 (N_16819,N_10085,N_11988);
nor U16820 (N_16820,N_14812,N_11606);
nand U16821 (N_16821,N_12557,N_10832);
xnor U16822 (N_16822,N_14038,N_14849);
nor U16823 (N_16823,N_11704,N_12181);
xnor U16824 (N_16824,N_13903,N_13342);
or U16825 (N_16825,N_11637,N_12034);
or U16826 (N_16826,N_14212,N_10628);
nand U16827 (N_16827,N_14954,N_11066);
nand U16828 (N_16828,N_10732,N_11192);
nor U16829 (N_16829,N_11631,N_14776);
xor U16830 (N_16830,N_14945,N_13686);
and U16831 (N_16831,N_10990,N_12379);
xnor U16832 (N_16832,N_12232,N_11371);
and U16833 (N_16833,N_14863,N_12830);
or U16834 (N_16834,N_13064,N_11376);
or U16835 (N_16835,N_12858,N_11486);
nor U16836 (N_16836,N_11965,N_11342);
and U16837 (N_16837,N_14060,N_11031);
nor U16838 (N_16838,N_12911,N_14479);
xor U16839 (N_16839,N_14880,N_14054);
or U16840 (N_16840,N_10752,N_13584);
and U16841 (N_16841,N_14193,N_13305);
nor U16842 (N_16842,N_14629,N_13687);
nor U16843 (N_16843,N_10563,N_11962);
xnor U16844 (N_16844,N_10853,N_11274);
or U16845 (N_16845,N_13350,N_13518);
nor U16846 (N_16846,N_14633,N_12783);
nor U16847 (N_16847,N_11276,N_10151);
xnor U16848 (N_16848,N_13851,N_14621);
xor U16849 (N_16849,N_10267,N_14024);
or U16850 (N_16850,N_12041,N_11766);
or U16851 (N_16851,N_12724,N_14351);
nor U16852 (N_16852,N_12264,N_13505);
or U16853 (N_16853,N_10215,N_11739);
nand U16854 (N_16854,N_13598,N_10436);
xor U16855 (N_16855,N_14374,N_11820);
or U16856 (N_16856,N_13239,N_13405);
xor U16857 (N_16857,N_11351,N_12641);
and U16858 (N_16858,N_10102,N_12387);
nand U16859 (N_16859,N_14510,N_14370);
or U16860 (N_16860,N_10096,N_13390);
nor U16861 (N_16861,N_13936,N_13616);
nand U16862 (N_16862,N_13902,N_11746);
xnor U16863 (N_16863,N_11205,N_13209);
xnor U16864 (N_16864,N_11252,N_12699);
or U16865 (N_16865,N_12063,N_13901);
nand U16866 (N_16866,N_12949,N_11802);
nor U16867 (N_16867,N_10228,N_11023);
nand U16868 (N_16868,N_11677,N_11325);
nand U16869 (N_16869,N_12664,N_14042);
or U16870 (N_16870,N_11547,N_12422);
nand U16871 (N_16871,N_11985,N_11512);
nand U16872 (N_16872,N_12647,N_11549);
and U16873 (N_16873,N_14276,N_10569);
or U16874 (N_16874,N_11362,N_14556);
or U16875 (N_16875,N_13290,N_14552);
nand U16876 (N_16876,N_11187,N_14867);
xor U16877 (N_16877,N_10859,N_13699);
xor U16878 (N_16878,N_11950,N_14718);
nor U16879 (N_16879,N_14809,N_14963);
nor U16880 (N_16880,N_12095,N_12513);
or U16881 (N_16881,N_13107,N_11600);
and U16882 (N_16882,N_10495,N_10405);
or U16883 (N_16883,N_14214,N_12080);
or U16884 (N_16884,N_12007,N_11519);
nor U16885 (N_16885,N_12972,N_11343);
and U16886 (N_16886,N_12183,N_13628);
nor U16887 (N_16887,N_10349,N_13800);
nor U16888 (N_16888,N_12810,N_13061);
nand U16889 (N_16889,N_13275,N_14636);
xnor U16890 (N_16890,N_13256,N_10531);
and U16891 (N_16891,N_10994,N_14981);
or U16892 (N_16892,N_11698,N_14637);
xnor U16893 (N_16893,N_14749,N_11352);
xor U16894 (N_16894,N_13248,N_10729);
xnor U16895 (N_16895,N_13858,N_12361);
and U16896 (N_16896,N_11444,N_13879);
nand U16897 (N_16897,N_12012,N_11536);
or U16898 (N_16898,N_11609,N_12885);
and U16899 (N_16899,N_14807,N_10836);
xor U16900 (N_16900,N_13211,N_12122);
nor U16901 (N_16901,N_12672,N_10472);
xnor U16902 (N_16902,N_10292,N_12923);
nand U16903 (N_16903,N_10007,N_11377);
or U16904 (N_16904,N_10224,N_11682);
nand U16905 (N_16905,N_10906,N_13272);
nor U16906 (N_16906,N_11484,N_12201);
xnor U16907 (N_16907,N_10111,N_11251);
nand U16908 (N_16908,N_13420,N_13801);
nor U16909 (N_16909,N_14174,N_13115);
nor U16910 (N_16910,N_11529,N_12743);
nand U16911 (N_16911,N_14740,N_10538);
nand U16912 (N_16912,N_10103,N_12296);
or U16913 (N_16913,N_12920,N_14754);
nor U16914 (N_16914,N_14584,N_10582);
or U16915 (N_16915,N_13230,N_11043);
or U16916 (N_16916,N_14080,N_10205);
nand U16917 (N_16917,N_12420,N_14026);
nand U16918 (N_16918,N_10302,N_13145);
and U16919 (N_16919,N_11741,N_14887);
nor U16920 (N_16920,N_11596,N_11201);
nand U16921 (N_16921,N_10263,N_13650);
xor U16922 (N_16922,N_12573,N_10567);
and U16923 (N_16923,N_12507,N_12376);
or U16924 (N_16924,N_10550,N_14915);
and U16925 (N_16925,N_13614,N_11436);
nand U16926 (N_16926,N_14884,N_11372);
nor U16927 (N_16927,N_13819,N_12447);
nor U16928 (N_16928,N_11789,N_12998);
nor U16929 (N_16929,N_10807,N_11282);
xor U16930 (N_16930,N_14574,N_12658);
nand U16931 (N_16931,N_13348,N_12146);
nand U16932 (N_16932,N_13312,N_13402);
xor U16933 (N_16933,N_11152,N_14890);
or U16934 (N_16934,N_12761,N_10390);
nand U16935 (N_16935,N_11172,N_12147);
or U16936 (N_16936,N_10399,N_13831);
and U16937 (N_16937,N_10779,N_12547);
and U16938 (N_16938,N_11409,N_10021);
xor U16939 (N_16939,N_13832,N_13778);
or U16940 (N_16940,N_14929,N_11259);
nor U16941 (N_16941,N_12461,N_13068);
nand U16942 (N_16942,N_14154,N_11901);
or U16943 (N_16943,N_13028,N_11092);
and U16944 (N_16944,N_10512,N_12054);
or U16945 (N_16945,N_11696,N_11723);
nor U16946 (N_16946,N_14824,N_13578);
nand U16947 (N_16947,N_10352,N_12261);
xnor U16948 (N_16948,N_14161,N_10514);
and U16949 (N_16949,N_12828,N_13207);
nor U16950 (N_16950,N_10125,N_14291);
xnor U16951 (N_16951,N_12266,N_10548);
nor U16952 (N_16952,N_14920,N_13555);
and U16953 (N_16953,N_11890,N_11759);
xor U16954 (N_16954,N_12773,N_13371);
xnor U16955 (N_16955,N_14677,N_10889);
xor U16956 (N_16956,N_10115,N_12044);
and U16957 (N_16957,N_10791,N_11389);
nor U16958 (N_16958,N_10746,N_14078);
or U16959 (N_16959,N_12378,N_11267);
nand U16960 (N_16960,N_12429,N_12769);
nand U16961 (N_16961,N_11021,N_10281);
or U16962 (N_16962,N_10985,N_13236);
or U16963 (N_16963,N_10608,N_14540);
nand U16964 (N_16964,N_11116,N_13195);
or U16965 (N_16965,N_11058,N_10695);
and U16966 (N_16966,N_10415,N_11692);
xnor U16967 (N_16967,N_12176,N_10723);
or U16968 (N_16968,N_12367,N_13012);
xnor U16969 (N_16969,N_14036,N_13081);
or U16970 (N_16970,N_11262,N_14962);
and U16971 (N_16971,N_14376,N_14632);
or U16972 (N_16972,N_14720,N_12585);
and U16973 (N_16973,N_14594,N_14361);
and U16974 (N_16974,N_10162,N_12739);
xnor U16975 (N_16975,N_10658,N_11322);
xor U16976 (N_16976,N_13593,N_13660);
or U16977 (N_16977,N_14287,N_14439);
nand U16978 (N_16978,N_10916,N_11944);
or U16979 (N_16979,N_13613,N_12069);
nand U16980 (N_16980,N_10001,N_12299);
or U16981 (N_16981,N_12802,N_13748);
or U16982 (N_16982,N_11752,N_14034);
or U16983 (N_16983,N_10011,N_13711);
nor U16984 (N_16984,N_11334,N_14942);
and U16985 (N_16985,N_14187,N_12915);
nor U16986 (N_16986,N_13164,N_14019);
nor U16987 (N_16987,N_13553,N_12271);
and U16988 (N_16988,N_10571,N_11301);
and U16989 (N_16989,N_13167,N_10986);
nand U16990 (N_16990,N_14375,N_14329);
nand U16991 (N_16991,N_12578,N_13173);
nand U16992 (N_16992,N_14413,N_13535);
nor U16993 (N_16993,N_14529,N_11439);
nor U16994 (N_16994,N_11044,N_13237);
nand U16995 (N_16995,N_11856,N_14231);
or U16996 (N_16996,N_14967,N_13761);
xor U16997 (N_16997,N_13928,N_14908);
xnor U16998 (N_16998,N_10871,N_14982);
nand U16999 (N_16999,N_12993,N_11188);
nor U17000 (N_17000,N_10667,N_12225);
nand U17001 (N_17001,N_10201,N_10771);
nor U17002 (N_17002,N_10109,N_13376);
and U17003 (N_17003,N_13171,N_11219);
and U17004 (N_17004,N_14043,N_11689);
nor U17005 (N_17005,N_11591,N_13354);
or U17006 (N_17006,N_10355,N_13807);
nor U17007 (N_17007,N_11190,N_13042);
or U17008 (N_17008,N_12835,N_14106);
nand U17009 (N_17009,N_11195,N_14021);
or U17010 (N_17010,N_13764,N_10464);
and U17011 (N_17011,N_14390,N_14628);
xor U17012 (N_17012,N_14958,N_10799);
and U17013 (N_17013,N_10907,N_13639);
nand U17014 (N_17014,N_12611,N_12583);
nor U17015 (N_17015,N_12648,N_12714);
xnor U17016 (N_17016,N_12892,N_13664);
nand U17017 (N_17017,N_12859,N_13733);
and U17018 (N_17018,N_11006,N_10171);
xnor U17019 (N_17019,N_14680,N_14132);
xnor U17020 (N_17020,N_11513,N_12862);
nand U17021 (N_17021,N_12377,N_12328);
or U17022 (N_17022,N_13734,N_11749);
xnor U17023 (N_17023,N_11260,N_13837);
xnor U17024 (N_17024,N_11153,N_13592);
nand U17025 (N_17025,N_11496,N_12016);
and U17026 (N_17026,N_12397,N_14293);
nor U17027 (N_17027,N_13942,N_12616);
nor U17028 (N_17028,N_10431,N_11694);
nand U17029 (N_17029,N_14096,N_10983);
nor U17030 (N_17030,N_13620,N_11518);
and U17031 (N_17031,N_13821,N_13695);
or U17032 (N_17032,N_10161,N_13344);
nand U17033 (N_17033,N_13132,N_10893);
or U17034 (N_17034,N_10589,N_13050);
or U17035 (N_17035,N_10433,N_11341);
nor U17036 (N_17036,N_14596,N_12774);
nor U17037 (N_17037,N_14081,N_13365);
and U17038 (N_17038,N_10197,N_10652);
or U17039 (N_17039,N_10318,N_14133);
and U17040 (N_17040,N_10311,N_14183);
or U17041 (N_17041,N_10289,N_14780);
and U17042 (N_17042,N_11469,N_11594);
or U17043 (N_17043,N_10486,N_13768);
nand U17044 (N_17044,N_12038,N_11041);
xnor U17045 (N_17045,N_10325,N_14424);
and U17046 (N_17046,N_14509,N_14613);
xnor U17047 (N_17047,N_12399,N_11261);
nand U17048 (N_17048,N_12419,N_11009);
or U17049 (N_17049,N_12305,N_11644);
or U17050 (N_17050,N_14377,N_14971);
nand U17051 (N_17051,N_11235,N_12753);
xnor U17052 (N_17052,N_13696,N_14650);
nor U17053 (N_17053,N_10104,N_11666);
xnor U17054 (N_17054,N_11593,N_11249);
or U17055 (N_17055,N_11680,N_12005);
nor U17056 (N_17056,N_14267,N_14347);
nor U17057 (N_17057,N_14505,N_12126);
or U17058 (N_17058,N_12516,N_14126);
or U17059 (N_17059,N_13062,N_14914);
and U17060 (N_17060,N_13076,N_12880);
or U17061 (N_17061,N_10158,N_10684);
nor U17062 (N_17062,N_14686,N_14846);
nor U17063 (N_17063,N_14605,N_11485);
xor U17064 (N_17064,N_12514,N_12486);
xnor U17065 (N_17065,N_10558,N_12838);
or U17066 (N_17066,N_11849,N_10803);
and U17067 (N_17067,N_10852,N_12721);
and U17068 (N_17068,N_13477,N_14833);
xnor U17069 (N_17069,N_12415,N_14378);
nor U17070 (N_17070,N_10332,N_14666);
or U17071 (N_17071,N_14533,N_13472);
nand U17072 (N_17072,N_14591,N_10946);
and U17073 (N_17073,N_14433,N_10322);
nand U17074 (N_17074,N_10740,N_10610);
xnor U17075 (N_17075,N_11776,N_10027);
or U17076 (N_17076,N_14030,N_14367);
or U17077 (N_17077,N_13792,N_13414);
or U17078 (N_17078,N_10635,N_11957);
nor U17079 (N_17079,N_10291,N_11788);
nand U17080 (N_17080,N_14032,N_13525);
and U17081 (N_17081,N_14466,N_14364);
xor U17082 (N_17082,N_13909,N_11358);
or U17083 (N_17083,N_12624,N_10181);
or U17084 (N_17084,N_13446,N_10766);
nor U17085 (N_17085,N_13287,N_11147);
or U17086 (N_17086,N_11279,N_11862);
nand U17087 (N_17087,N_11860,N_11869);
and U17088 (N_17088,N_11424,N_10286);
and U17089 (N_17089,N_14359,N_14790);
xnor U17090 (N_17090,N_14324,N_14396);
nand U17091 (N_17091,N_13682,N_13637);
nand U17092 (N_17092,N_10769,N_14142);
nor U17093 (N_17093,N_13217,N_14983);
and U17094 (N_17094,N_12518,N_12148);
nand U17095 (N_17095,N_13283,N_14199);
nor U17096 (N_17096,N_14687,N_11706);
xor U17097 (N_17097,N_12527,N_14499);
or U17098 (N_17098,N_11271,N_10377);
and U17099 (N_17099,N_10422,N_13977);
xor U17100 (N_17100,N_13313,N_13904);
nor U17101 (N_17101,N_11303,N_13044);
nand U17102 (N_17102,N_13685,N_13298);
or U17103 (N_17103,N_10400,N_13241);
or U17104 (N_17104,N_13255,N_13739);
xnor U17105 (N_17105,N_14862,N_10310);
nor U17106 (N_17106,N_10347,N_13407);
or U17107 (N_17107,N_12909,N_12371);
or U17108 (N_17108,N_12799,N_11715);
and U17109 (N_17109,N_12318,N_10437);
or U17110 (N_17110,N_14191,N_12782);
xor U17111 (N_17111,N_12317,N_13188);
nor U17112 (N_17112,N_12035,N_13128);
or U17113 (N_17113,N_11514,N_11996);
nand U17114 (N_17114,N_10790,N_11051);
xnor U17115 (N_17115,N_14734,N_13959);
xnor U17116 (N_17116,N_13529,N_14930);
and U17117 (N_17117,N_10126,N_14478);
xnor U17118 (N_17118,N_12365,N_11418);
nor U17119 (N_17119,N_13999,N_12141);
xnor U17120 (N_17120,N_11468,N_13024);
nand U17121 (N_17121,N_11471,N_12446);
xnor U17122 (N_17122,N_14047,N_14194);
and U17123 (N_17123,N_13395,N_12433);
nand U17124 (N_17124,N_10304,N_13630);
or U17125 (N_17125,N_12453,N_12651);
xor U17126 (N_17126,N_10783,N_12888);
nor U17127 (N_17127,N_13329,N_10040);
xnor U17128 (N_17128,N_11709,N_14975);
nand U17129 (N_17129,N_11397,N_13815);
nor U17130 (N_17130,N_11503,N_10202);
and U17131 (N_17131,N_10398,N_11243);
or U17132 (N_17132,N_13463,N_14422);
nand U17133 (N_17133,N_11034,N_12286);
and U17134 (N_17134,N_11597,N_13408);
and U17135 (N_17135,N_11611,N_14513);
and U17136 (N_17136,N_14092,N_11977);
or U17137 (N_17137,N_10777,N_13270);
and U17138 (N_17138,N_11538,N_12247);
or U17139 (N_17139,N_12676,N_12740);
and U17140 (N_17140,N_10880,N_11106);
and U17141 (N_17141,N_10172,N_13973);
or U17142 (N_17142,N_11889,N_12131);
xnor U17143 (N_17143,N_10116,N_11011);
and U17144 (N_17144,N_10160,N_12064);
or U17145 (N_17145,N_13415,N_10461);
nand U17146 (N_17146,N_11610,N_12517);
xnor U17147 (N_17147,N_11653,N_13015);
nand U17148 (N_17148,N_13642,N_10259);
xor U17149 (N_17149,N_13641,N_10136);
xnor U17150 (N_17150,N_11375,N_10092);
and U17151 (N_17151,N_11218,N_11084);
nand U17152 (N_17152,N_13753,N_12827);
and U17153 (N_17153,N_13689,N_13161);
and U17154 (N_17154,N_11998,N_11589);
nor U17155 (N_17155,N_14127,N_13726);
nor U17156 (N_17156,N_14318,N_12592);
or U17157 (N_17157,N_14497,N_12216);
or U17158 (N_17158,N_14653,N_11292);
nand U17159 (N_17159,N_11845,N_12841);
nand U17160 (N_17160,N_10273,N_12918);
nand U17161 (N_17161,N_13930,N_13870);
nand U17162 (N_17162,N_10555,N_13056);
and U17163 (N_17163,N_11165,N_12896);
nand U17164 (N_17164,N_13622,N_12388);
xor U17165 (N_17165,N_13120,N_14119);
or U17166 (N_17166,N_12215,N_11161);
nor U17167 (N_17167,N_14273,N_11264);
nor U17168 (N_17168,N_10689,N_10288);
xnor U17169 (N_17169,N_12355,N_11115);
xnor U17170 (N_17170,N_13259,N_13426);
and U17171 (N_17171,N_11824,N_11537);
and U17172 (N_17172,N_14400,N_10028);
or U17173 (N_17173,N_10734,N_13325);
nor U17174 (N_17174,N_13269,N_13499);
and U17175 (N_17175,N_13017,N_12853);
or U17176 (N_17176,N_11050,N_13793);
nand U17177 (N_17177,N_12558,N_10279);
nor U17178 (N_17178,N_14959,N_13825);
or U17179 (N_17179,N_14073,N_14956);
nand U17180 (N_17180,N_11138,N_12259);
or U17181 (N_17181,N_13225,N_14583);
nand U17182 (N_17182,N_12586,N_14568);
or U17183 (N_17183,N_10122,N_10014);
nand U17184 (N_17184,N_12125,N_14973);
nand U17185 (N_17185,N_14543,N_12250);
nand U17186 (N_17186,N_13204,N_12116);
nor U17187 (N_17187,N_14885,N_14595);
xor U17188 (N_17188,N_10036,N_13910);
xor U17189 (N_17189,N_10692,N_12851);
nand U17190 (N_17190,N_12522,N_14256);
and U17191 (N_17191,N_13243,N_14207);
or U17192 (N_17192,N_13694,N_12546);
and U17193 (N_17193,N_14284,N_14163);
and U17194 (N_17194,N_14063,N_13033);
xor U17195 (N_17195,N_10204,N_13380);
and U17196 (N_17196,N_11382,N_11960);
and U17197 (N_17197,N_13498,N_13251);
or U17198 (N_17198,N_13224,N_11185);
nor U17199 (N_17199,N_14288,N_13813);
nand U17200 (N_17200,N_11211,N_11764);
and U17201 (N_17201,N_10537,N_11309);
or U17202 (N_17202,N_12480,N_10041);
nand U17203 (N_17203,N_11460,N_12053);
or U17204 (N_17204,N_12430,N_11340);
xnor U17205 (N_17205,N_11946,N_10169);
xnor U17206 (N_17206,N_10315,N_11320);
nand U17207 (N_17207,N_10207,N_11577);
xnor U17208 (N_17208,N_10002,N_12134);
and U17209 (N_17209,N_11142,N_11466);
or U17210 (N_17210,N_10142,N_12495);
and U17211 (N_17211,N_11861,N_13264);
nand U17212 (N_17212,N_14501,N_13523);
nor U17213 (N_17213,N_10921,N_13701);
nand U17214 (N_17214,N_10655,N_14105);
and U17215 (N_17215,N_14643,N_14729);
and U17216 (N_17216,N_14919,N_11272);
nand U17217 (N_17217,N_11821,N_14871);
or U17218 (N_17218,N_11686,N_13503);
nand U17219 (N_17219,N_11853,N_14985);
or U17220 (N_17220,N_11239,N_14593);
nand U17221 (N_17221,N_12988,N_10424);
or U17222 (N_17222,N_14225,N_13652);
nor U17223 (N_17223,N_10900,N_14446);
xor U17224 (N_17224,N_11278,N_11217);
and U17225 (N_17225,N_12965,N_10708);
xnor U17226 (N_17226,N_10879,N_10137);
nand U17227 (N_17227,N_12108,N_10774);
xor U17228 (N_17228,N_10039,N_13092);
and U17229 (N_17229,N_11711,N_12679);
xnor U17230 (N_17230,N_10869,N_11321);
nand U17231 (N_17231,N_12515,N_13083);
and U17232 (N_17232,N_13184,N_14448);
xor U17233 (N_17233,N_10941,N_10469);
and U17234 (N_17234,N_12789,N_10334);
nand U17235 (N_17235,N_10694,N_11442);
nand U17236 (N_17236,N_12668,N_12129);
nor U17237 (N_17237,N_14625,N_10195);
xor U17238 (N_17238,N_12917,N_13937);
nand U17239 (N_17239,N_10331,N_13919);
nor U17240 (N_17240,N_13258,N_12028);
and U17241 (N_17241,N_10532,N_14854);
and U17242 (N_17242,N_11854,N_12817);
or U17243 (N_17243,N_14089,N_10084);
xnor U17244 (N_17244,N_14599,N_10396);
nand U17245 (N_17245,N_12235,N_13278);
and U17246 (N_17246,N_13720,N_14527);
nand U17247 (N_17247,N_12598,N_12381);
or U17248 (N_17248,N_10527,N_13346);
xor U17249 (N_17249,N_12511,N_10506);
nor U17250 (N_17250,N_14773,N_10231);
nand U17251 (N_17251,N_13775,N_10754);
or U17252 (N_17252,N_10834,N_14572);
nor U17253 (N_17253,N_12763,N_14409);
xnor U17254 (N_17254,N_10539,N_11792);
nand U17255 (N_17255,N_11515,N_14836);
xor U17256 (N_17256,N_13306,N_13153);
or U17257 (N_17257,N_11751,N_11959);
nor U17258 (N_17258,N_12529,N_14676);
nand U17259 (N_17259,N_12196,N_10208);
xor U17260 (N_17260,N_11628,N_14675);
nand U17261 (N_17261,N_12018,N_13961);
nor U17262 (N_17262,N_12184,N_12283);
xor U17263 (N_17263,N_14294,N_13192);
xnor U17264 (N_17264,N_10082,N_13226);
and U17265 (N_17265,N_11453,N_11297);
nand U17266 (N_17266,N_12071,N_10156);
and U17267 (N_17267,N_13392,N_12626);
or U17268 (N_17268,N_12925,N_12625);
and U17269 (N_17269,N_10728,N_11929);
and U17270 (N_17270,N_14791,N_11586);
and U17271 (N_17271,N_10676,N_10356);
nand U17272 (N_17272,N_13317,N_14357);
xor U17273 (N_17273,N_14165,N_11662);
or U17274 (N_17274,N_14346,N_14542);
nand U17275 (N_17275,N_12621,N_13742);
xor U17276 (N_17276,N_10030,N_11091);
or U17277 (N_17277,N_11121,N_10057);
nand U17278 (N_17278,N_12066,N_11773);
xor U17279 (N_17279,N_10673,N_14023);
xor U17280 (N_17280,N_10630,N_10885);
or U17281 (N_17281,N_12268,N_10787);
xnor U17282 (N_17282,N_14339,N_11635);
xor U17283 (N_17283,N_11227,N_14300);
xor U17284 (N_17284,N_11894,N_13175);
or U17285 (N_17285,N_12140,N_10984);
or U17286 (N_17286,N_13993,N_12097);
and U17287 (N_17287,N_14271,N_12468);
xor U17288 (N_17288,N_10046,N_12408);
xor U17289 (N_17289,N_11921,N_12560);
and U17290 (N_17290,N_10029,N_14978);
nor U17291 (N_17291,N_11987,N_12026);
and U17292 (N_17292,N_10200,N_13732);
and U17293 (N_17293,N_12011,N_13469);
and U17294 (N_17294,N_11331,N_14068);
xor U17295 (N_17295,N_12634,N_14185);
xor U17296 (N_17296,N_12532,N_10956);
nor U17297 (N_17297,N_14506,N_10308);
xor U17298 (N_17298,N_12970,N_14362);
and U17299 (N_17299,N_10120,N_10620);
nor U17300 (N_17300,N_12333,N_14395);
or U17301 (N_17301,N_13745,N_11314);
nand U17302 (N_17302,N_12262,N_10293);
nor U17303 (N_17303,N_10242,N_14895);
and U17304 (N_17304,N_11125,N_14044);
and U17305 (N_17305,N_11283,N_12932);
xnor U17306 (N_17306,N_10203,N_12081);
xnor U17307 (N_17307,N_11750,N_13080);
nor U17308 (N_17308,N_10309,N_10511);
nand U17309 (N_17309,N_11012,N_11209);
xnor U17310 (N_17310,N_14913,N_13155);
nand U17311 (N_17311,N_11403,N_10023);
or U17312 (N_17312,N_10530,N_13398);
nor U17313 (N_17313,N_12331,N_13135);
nand U17314 (N_17314,N_13268,N_11936);
or U17315 (N_17315,N_11456,N_13389);
nor U17316 (N_17316,N_11385,N_11993);
nand U17317 (N_17317,N_11671,N_10155);
and U17318 (N_17318,N_13964,N_14386);
or U17319 (N_17319,N_10805,N_12628);
or U17320 (N_17320,N_14005,N_14438);
nor U17321 (N_17321,N_11991,N_13577);
xnor U17322 (N_17322,N_13597,N_11158);
and U17323 (N_17323,N_10765,N_11915);
xor U17324 (N_17324,N_10797,N_14209);
nor U17325 (N_17325,N_10828,N_10020);
nor U17326 (N_17326,N_13386,N_14086);
xnor U17327 (N_17327,N_12339,N_11220);
and U17328 (N_17328,N_10977,N_12619);
nand U17329 (N_17329,N_14663,N_13449);
nand U17330 (N_17330,N_13853,N_13956);
and U17331 (N_17331,N_13156,N_13531);
nand U17332 (N_17332,N_10596,N_11982);
nor U17333 (N_17333,N_11163,N_12281);
nand U17334 (N_17334,N_14703,N_14334);
and U17335 (N_17335,N_10894,N_14496);
or U17336 (N_17336,N_11842,N_14566);
or U17337 (N_17337,N_10664,N_14253);
nor U17338 (N_17338,N_11336,N_11032);
and U17339 (N_17339,N_14156,N_13245);
and U17340 (N_17340,N_13784,N_10913);
nor U17341 (N_17341,N_14953,N_10715);
and U17342 (N_17342,N_14753,N_11942);
nand U17343 (N_17343,N_13541,N_11952);
and U17344 (N_17344,N_14075,N_14853);
nor U17345 (N_17345,N_10577,N_12273);
xnor U17346 (N_17346,N_10282,N_13293);
and U17347 (N_17347,N_13850,N_14575);
or U17348 (N_17348,N_13455,N_13841);
and U17349 (N_17349,N_13121,N_14066);
or U17350 (N_17350,N_11333,N_11452);
and U17351 (N_17351,N_13861,N_11405);
xnor U17352 (N_17352,N_10888,N_14704);
nand U17353 (N_17353,N_13635,N_12579);
and U17354 (N_17354,N_11502,N_11557);
and U17355 (N_17355,N_12757,N_14251);
and U17356 (N_17356,N_12548,N_13143);
nand U17357 (N_17357,N_14355,N_10168);
or U17358 (N_17358,N_11049,N_13500);
nor U17359 (N_17359,N_14173,N_12185);
nand U17360 (N_17360,N_12784,N_12090);
nand U17361 (N_17361,N_11679,N_14847);
and U17362 (N_17362,N_11781,N_10274);
nor U17363 (N_17363,N_11876,N_11816);
nor U17364 (N_17364,N_11882,N_12178);
and U17365 (N_17365,N_11836,N_10381);
nand U17366 (N_17366,N_14136,N_12788);
nand U17367 (N_17367,N_10248,N_12191);
xnor U17368 (N_17368,N_14581,N_14805);
and U17369 (N_17369,N_14333,N_11109);
xor U17370 (N_17370,N_10528,N_11077);
xor U17371 (N_17371,N_10221,N_13148);
nand U17372 (N_17372,N_13375,N_10059);
nand U17373 (N_17373,N_12001,N_11923);
nand U17374 (N_17374,N_11408,N_14262);
and U17375 (N_17375,N_11079,N_10751);
or U17376 (N_17376,N_14349,N_14065);
xnor U17377 (N_17377,N_10175,N_11094);
nand U17378 (N_17378,N_14418,N_10671);
nand U17379 (N_17379,N_14428,N_14115);
nor U17380 (N_17380,N_13432,N_10410);
nor U17381 (N_17381,N_13014,N_10378);
nor U17382 (N_17382,N_13795,N_12695);
or U17383 (N_17383,N_10574,N_11210);
xnor U17384 (N_17384,N_14700,N_10773);
nand U17385 (N_17385,N_13543,N_14280);
nand U17386 (N_17386,N_10578,N_14195);
or U17387 (N_17387,N_13149,N_14601);
nand U17388 (N_17388,N_14932,N_14774);
and U17389 (N_17389,N_14489,N_14974);
xnor U17390 (N_17390,N_12814,N_11497);
nor U17391 (N_17391,N_13954,N_14436);
nand U17392 (N_17392,N_11580,N_12075);
nand U17393 (N_17393,N_13481,N_12902);
xnor U17394 (N_17394,N_14866,N_11947);
and U17395 (N_17395,N_11727,N_12163);
and U17396 (N_17396,N_11913,N_14070);
nor U17397 (N_17397,N_13913,N_14547);
nand U17398 (N_17398,N_12635,N_11945);
and U17399 (N_17399,N_10873,N_13771);
or U17400 (N_17400,N_14379,N_11919);
nor U17401 (N_17401,N_13986,N_11758);
nor U17402 (N_17402,N_12781,N_12123);
and U17403 (N_17403,N_13231,N_12315);
and U17404 (N_17404,N_10753,N_12563);
and U17405 (N_17405,N_12762,N_12319);
nor U17406 (N_17406,N_14013,N_13547);
xnor U17407 (N_17407,N_11674,N_12393);
nor U17408 (N_17408,N_10294,N_13029);
xnor U17409 (N_17409,N_10768,N_11465);
nand U17410 (N_17410,N_10493,N_14736);
or U17411 (N_17411,N_10226,N_11684);
nand U17412 (N_17412,N_10067,N_11774);
nand U17413 (N_17413,N_14798,N_11652);
nor U17414 (N_17414,N_10141,N_14896);
nand U17415 (N_17415,N_14122,N_12417);
and U17416 (N_17416,N_13279,N_10189);
or U17417 (N_17417,N_14564,N_12509);
nand U17418 (N_17418,N_14462,N_14148);
xnor U17419 (N_17419,N_10716,N_11140);
nand U17420 (N_17420,N_14511,N_12564);
xnor U17421 (N_17421,N_12595,N_13097);
and U17422 (N_17422,N_11804,N_10645);
nand U17423 (N_17423,N_11123,N_14304);
nand U17424 (N_17424,N_14775,N_10587);
or U17425 (N_17425,N_11841,N_12866);
nand U17426 (N_17426,N_13214,N_14735);
and U17427 (N_17427,N_11871,N_12623);
or U17428 (N_17428,N_14811,N_11602);
or U17429 (N_17429,N_11714,N_10632);
or U17430 (N_17430,N_13253,N_10622);
nor U17431 (N_17431,N_10711,N_13548);
or U17432 (N_17432,N_12015,N_12645);
and U17433 (N_17433,N_12823,N_13212);
nor U17434 (N_17434,N_14690,N_14440);
nand U17435 (N_17435,N_10333,N_11907);
nand U17436 (N_17436,N_10094,N_14250);
nor U17437 (N_17437,N_12109,N_12155);
nand U17438 (N_17438,N_10276,N_13849);
xor U17439 (N_17439,N_13223,N_10770);
or U17440 (N_17440,N_14369,N_11990);
or U17441 (N_17441,N_13133,N_11476);
or U17442 (N_17442,N_12504,N_13197);
and U17443 (N_17443,N_14683,N_13866);
nand U17444 (N_17444,N_11713,N_14551);
or U17445 (N_17445,N_10138,N_10572);
nor U17446 (N_17446,N_12055,N_13060);
nor U17447 (N_17447,N_13129,N_10614);
nand U17448 (N_17448,N_10229,N_13001);
or U17449 (N_17449,N_11843,N_10993);
xor U17450 (N_17450,N_11087,N_12661);
xor U17451 (N_17451,N_14391,N_11306);
or U17452 (N_17452,N_14850,N_12593);
nand U17453 (N_17453,N_10520,N_14500);
nand U17454 (N_17454,N_14901,N_12455);
nor U17455 (N_17455,N_14525,N_10642);
xor U17456 (N_17456,N_11492,N_12722);
and U17457 (N_17457,N_12929,N_14099);
and U17458 (N_17458,N_12025,N_14077);
nor U17459 (N_17459,N_13590,N_14578);
or U17460 (N_17460,N_13984,N_14544);
and U17461 (N_17461,N_13600,N_10178);
nand U17462 (N_17462,N_10107,N_11124);
xor U17463 (N_17463,N_14679,N_13927);
nand U17464 (N_17464,N_12460,N_12091);
xor U17465 (N_17465,N_10435,N_12174);
xor U17466 (N_17466,N_12691,N_12363);
xnor U17467 (N_17467,N_11132,N_13681);
xor U17468 (N_17468,N_12878,N_12889);
xor U17469 (N_17469,N_12512,N_13981);
and U17470 (N_17470,N_13991,N_12366);
xnor U17471 (N_17471,N_10299,N_10397);
nor U17472 (N_17472,N_11661,N_10955);
or U17473 (N_17473,N_10072,N_10872);
or U17474 (N_17474,N_11215,N_12476);
and U17475 (N_17475,N_12941,N_14557);
nor U17476 (N_17476,N_14695,N_11516);
nor U17477 (N_17477,N_11237,N_10100);
nor U17478 (N_17478,N_11487,N_11015);
nand U17479 (N_17479,N_13222,N_10479);
or U17480 (N_17480,N_12700,N_10455);
xor U17481 (N_17481,N_11374,N_10821);
and U17482 (N_17482,N_14234,N_12465);
nor U17483 (N_17483,N_13894,N_10827);
and U17484 (N_17484,N_11873,N_12727);
and U17485 (N_17485,N_13520,N_10496);
or U17486 (N_17486,N_11415,N_13868);
nand U17487 (N_17487,N_13610,N_12209);
or U17488 (N_17488,N_11800,N_12231);
nor U17489 (N_17489,N_14986,N_13576);
or U17490 (N_17490,N_12577,N_14577);
nand U17491 (N_17491,N_13310,N_11177);
or U17492 (N_17492,N_13416,N_12541);
xor U17493 (N_17493,N_14512,N_13912);
or U17494 (N_17494,N_13856,N_10696);
or U17495 (N_17495,N_14782,N_13985);
and U17496 (N_17496,N_13331,N_12128);
nor U17497 (N_17497,N_14576,N_11874);
or U17498 (N_17498,N_10443,N_14620);
xor U17499 (N_17499,N_10892,N_14767);
nor U17500 (N_17500,N_13752,N_14799);
nor U17501 (N_17501,N_13148,N_14474);
and U17502 (N_17502,N_12809,N_12887);
and U17503 (N_17503,N_11916,N_14376);
and U17504 (N_17504,N_11221,N_11372);
xnor U17505 (N_17505,N_14729,N_14332);
or U17506 (N_17506,N_11277,N_14364);
nor U17507 (N_17507,N_10871,N_14169);
xnor U17508 (N_17508,N_13611,N_10198);
or U17509 (N_17509,N_14020,N_10348);
xnor U17510 (N_17510,N_11575,N_11486);
nand U17511 (N_17511,N_10987,N_13246);
nand U17512 (N_17512,N_14849,N_10864);
xnor U17513 (N_17513,N_13266,N_11452);
xor U17514 (N_17514,N_12607,N_14466);
and U17515 (N_17515,N_11130,N_13002);
or U17516 (N_17516,N_12295,N_14736);
nand U17517 (N_17517,N_13833,N_11887);
xor U17518 (N_17518,N_11646,N_10223);
nand U17519 (N_17519,N_14425,N_12529);
xnor U17520 (N_17520,N_13611,N_12640);
nand U17521 (N_17521,N_11610,N_11811);
or U17522 (N_17522,N_12857,N_14144);
or U17523 (N_17523,N_12735,N_10426);
or U17524 (N_17524,N_10663,N_12812);
nand U17525 (N_17525,N_13668,N_13972);
xnor U17526 (N_17526,N_13691,N_12284);
and U17527 (N_17527,N_12338,N_10637);
and U17528 (N_17528,N_11867,N_10639);
and U17529 (N_17529,N_11335,N_12524);
nand U17530 (N_17530,N_13056,N_11230);
nor U17531 (N_17531,N_13784,N_14967);
and U17532 (N_17532,N_13839,N_14103);
or U17533 (N_17533,N_12811,N_13374);
xor U17534 (N_17534,N_14004,N_11637);
nand U17535 (N_17535,N_12315,N_14484);
nor U17536 (N_17536,N_11298,N_13801);
or U17537 (N_17537,N_11290,N_11750);
xor U17538 (N_17538,N_11377,N_12324);
nor U17539 (N_17539,N_12912,N_12216);
nor U17540 (N_17540,N_11458,N_12608);
and U17541 (N_17541,N_14493,N_11009);
and U17542 (N_17542,N_11209,N_12788);
nand U17543 (N_17543,N_10061,N_10795);
nand U17544 (N_17544,N_12229,N_11675);
and U17545 (N_17545,N_12276,N_11032);
nor U17546 (N_17546,N_10785,N_13847);
xnor U17547 (N_17547,N_10202,N_10948);
nor U17548 (N_17548,N_11884,N_12884);
or U17549 (N_17549,N_13120,N_14069);
or U17550 (N_17550,N_11656,N_14317);
and U17551 (N_17551,N_13058,N_11216);
nand U17552 (N_17552,N_13521,N_13995);
or U17553 (N_17553,N_11888,N_14937);
xnor U17554 (N_17554,N_14454,N_10870);
nand U17555 (N_17555,N_13020,N_10855);
nor U17556 (N_17556,N_10922,N_12969);
and U17557 (N_17557,N_14555,N_14835);
nand U17558 (N_17558,N_11409,N_10827);
xnor U17559 (N_17559,N_10149,N_13736);
nand U17560 (N_17560,N_11573,N_13526);
and U17561 (N_17561,N_11870,N_10823);
nand U17562 (N_17562,N_11229,N_12278);
or U17563 (N_17563,N_12397,N_10693);
and U17564 (N_17564,N_14550,N_12354);
xor U17565 (N_17565,N_11861,N_11402);
nor U17566 (N_17566,N_10211,N_13662);
nor U17567 (N_17567,N_13582,N_12542);
xor U17568 (N_17568,N_12456,N_10224);
xor U17569 (N_17569,N_11998,N_10119);
or U17570 (N_17570,N_11269,N_10782);
or U17571 (N_17571,N_10372,N_10167);
xnor U17572 (N_17572,N_14022,N_11752);
or U17573 (N_17573,N_14789,N_14942);
xnor U17574 (N_17574,N_11353,N_10861);
xnor U17575 (N_17575,N_12463,N_10610);
nand U17576 (N_17576,N_13197,N_10876);
nand U17577 (N_17577,N_10029,N_14195);
nand U17578 (N_17578,N_13672,N_14689);
xnor U17579 (N_17579,N_11823,N_13780);
or U17580 (N_17580,N_14079,N_10506);
xor U17581 (N_17581,N_12464,N_11229);
or U17582 (N_17582,N_13053,N_14893);
or U17583 (N_17583,N_13114,N_13926);
xor U17584 (N_17584,N_10302,N_12401);
nor U17585 (N_17585,N_12927,N_14606);
or U17586 (N_17586,N_12554,N_10028);
xor U17587 (N_17587,N_13711,N_14856);
xnor U17588 (N_17588,N_14497,N_14526);
nor U17589 (N_17589,N_11839,N_12163);
and U17590 (N_17590,N_13679,N_14218);
and U17591 (N_17591,N_14312,N_11197);
nand U17592 (N_17592,N_11391,N_13232);
nor U17593 (N_17593,N_11447,N_10400);
and U17594 (N_17594,N_11428,N_11104);
and U17595 (N_17595,N_11106,N_12327);
and U17596 (N_17596,N_14323,N_10431);
nor U17597 (N_17597,N_13446,N_14092);
nor U17598 (N_17598,N_13709,N_13710);
nor U17599 (N_17599,N_14403,N_12367);
xor U17600 (N_17600,N_12687,N_11925);
and U17601 (N_17601,N_11998,N_14313);
nand U17602 (N_17602,N_10965,N_14397);
or U17603 (N_17603,N_13380,N_11441);
nor U17604 (N_17604,N_14397,N_11174);
and U17605 (N_17605,N_11168,N_10556);
nand U17606 (N_17606,N_13170,N_10843);
and U17607 (N_17607,N_14339,N_14376);
nand U17608 (N_17608,N_13199,N_14172);
or U17609 (N_17609,N_14013,N_14433);
nor U17610 (N_17610,N_11605,N_11544);
nand U17611 (N_17611,N_13841,N_10035);
and U17612 (N_17612,N_11789,N_11766);
or U17613 (N_17613,N_14664,N_11639);
nor U17614 (N_17614,N_12576,N_12893);
and U17615 (N_17615,N_14269,N_10118);
nand U17616 (N_17616,N_11340,N_10306);
or U17617 (N_17617,N_12916,N_14311);
nor U17618 (N_17618,N_13072,N_12998);
nor U17619 (N_17619,N_11509,N_12487);
xor U17620 (N_17620,N_13427,N_10890);
nand U17621 (N_17621,N_12605,N_10411);
and U17622 (N_17622,N_11527,N_13783);
and U17623 (N_17623,N_11767,N_14246);
nand U17624 (N_17624,N_12489,N_14079);
nor U17625 (N_17625,N_12562,N_11335);
or U17626 (N_17626,N_14709,N_12057);
xor U17627 (N_17627,N_10321,N_14213);
xor U17628 (N_17628,N_10969,N_13975);
xnor U17629 (N_17629,N_10243,N_10278);
xnor U17630 (N_17630,N_14480,N_10256);
xnor U17631 (N_17631,N_10622,N_14543);
xor U17632 (N_17632,N_11301,N_14459);
xor U17633 (N_17633,N_11522,N_12981);
and U17634 (N_17634,N_10853,N_12739);
or U17635 (N_17635,N_11041,N_11738);
nor U17636 (N_17636,N_13866,N_10352);
nand U17637 (N_17637,N_11670,N_11829);
and U17638 (N_17638,N_10010,N_10622);
xnor U17639 (N_17639,N_14866,N_13421);
and U17640 (N_17640,N_13363,N_12923);
and U17641 (N_17641,N_12778,N_10246);
or U17642 (N_17642,N_12924,N_10181);
and U17643 (N_17643,N_14523,N_12012);
and U17644 (N_17644,N_14027,N_14596);
nand U17645 (N_17645,N_10763,N_10103);
nor U17646 (N_17646,N_10466,N_14658);
nor U17647 (N_17647,N_10222,N_12026);
xor U17648 (N_17648,N_10242,N_10117);
nand U17649 (N_17649,N_10503,N_11215);
xnor U17650 (N_17650,N_12111,N_11156);
or U17651 (N_17651,N_10653,N_13567);
or U17652 (N_17652,N_10735,N_13445);
and U17653 (N_17653,N_12311,N_13608);
xnor U17654 (N_17654,N_12324,N_14285);
nor U17655 (N_17655,N_10634,N_12189);
nand U17656 (N_17656,N_11613,N_12424);
nor U17657 (N_17657,N_12890,N_11469);
and U17658 (N_17658,N_14691,N_14404);
xnor U17659 (N_17659,N_13951,N_12477);
nand U17660 (N_17660,N_11105,N_14887);
nand U17661 (N_17661,N_13994,N_12909);
and U17662 (N_17662,N_13068,N_12293);
nor U17663 (N_17663,N_12724,N_11205);
nor U17664 (N_17664,N_11584,N_14656);
nand U17665 (N_17665,N_13162,N_12872);
and U17666 (N_17666,N_14207,N_13757);
xnor U17667 (N_17667,N_11424,N_13042);
nand U17668 (N_17668,N_12068,N_10446);
nand U17669 (N_17669,N_13383,N_12461);
nor U17670 (N_17670,N_12462,N_11915);
xnor U17671 (N_17671,N_14639,N_11812);
nand U17672 (N_17672,N_13816,N_10421);
xnor U17673 (N_17673,N_13441,N_14073);
nor U17674 (N_17674,N_11479,N_14149);
xnor U17675 (N_17675,N_13105,N_13127);
or U17676 (N_17676,N_11716,N_12245);
and U17677 (N_17677,N_14614,N_13550);
and U17678 (N_17678,N_10930,N_13566);
xor U17679 (N_17679,N_10937,N_11522);
or U17680 (N_17680,N_11709,N_13554);
or U17681 (N_17681,N_12266,N_12987);
and U17682 (N_17682,N_13366,N_13481);
nor U17683 (N_17683,N_11917,N_13998);
nand U17684 (N_17684,N_13786,N_11329);
xor U17685 (N_17685,N_14371,N_12616);
and U17686 (N_17686,N_13144,N_13835);
or U17687 (N_17687,N_14072,N_10502);
and U17688 (N_17688,N_11740,N_13630);
or U17689 (N_17689,N_10450,N_11780);
nor U17690 (N_17690,N_12173,N_13970);
and U17691 (N_17691,N_11536,N_11825);
nand U17692 (N_17692,N_13845,N_10498);
xnor U17693 (N_17693,N_10555,N_12679);
or U17694 (N_17694,N_14959,N_12633);
nand U17695 (N_17695,N_11417,N_10141);
or U17696 (N_17696,N_12330,N_10975);
nor U17697 (N_17697,N_11599,N_12464);
or U17698 (N_17698,N_13738,N_11329);
and U17699 (N_17699,N_12703,N_11820);
or U17700 (N_17700,N_13365,N_13515);
and U17701 (N_17701,N_14145,N_10098);
nand U17702 (N_17702,N_14747,N_12731);
nand U17703 (N_17703,N_11172,N_12505);
or U17704 (N_17704,N_11443,N_12826);
xnor U17705 (N_17705,N_14797,N_12212);
nand U17706 (N_17706,N_14795,N_14382);
nor U17707 (N_17707,N_14724,N_12402);
and U17708 (N_17708,N_14812,N_12555);
xor U17709 (N_17709,N_12369,N_14772);
or U17710 (N_17710,N_11395,N_12913);
xor U17711 (N_17711,N_11315,N_11152);
and U17712 (N_17712,N_13315,N_12725);
nor U17713 (N_17713,N_11969,N_10586);
or U17714 (N_17714,N_10019,N_10468);
nand U17715 (N_17715,N_11907,N_14451);
or U17716 (N_17716,N_14600,N_12166);
xnor U17717 (N_17717,N_11876,N_11450);
or U17718 (N_17718,N_14810,N_12496);
nor U17719 (N_17719,N_11280,N_11746);
nand U17720 (N_17720,N_12667,N_13022);
nor U17721 (N_17721,N_10084,N_12996);
or U17722 (N_17722,N_14011,N_12662);
nor U17723 (N_17723,N_12474,N_12731);
or U17724 (N_17724,N_14215,N_10420);
nor U17725 (N_17725,N_12426,N_12138);
xnor U17726 (N_17726,N_12351,N_14481);
xnor U17727 (N_17727,N_14401,N_11413);
or U17728 (N_17728,N_10127,N_13145);
and U17729 (N_17729,N_13373,N_12155);
or U17730 (N_17730,N_13885,N_14485);
xnor U17731 (N_17731,N_11342,N_12396);
nor U17732 (N_17732,N_14129,N_14197);
nor U17733 (N_17733,N_12856,N_13480);
xor U17734 (N_17734,N_12602,N_12671);
nor U17735 (N_17735,N_13164,N_14912);
nand U17736 (N_17736,N_13354,N_11108);
nand U17737 (N_17737,N_14522,N_14374);
nand U17738 (N_17738,N_11078,N_13748);
xor U17739 (N_17739,N_13340,N_10874);
nand U17740 (N_17740,N_10065,N_12793);
or U17741 (N_17741,N_13141,N_12090);
or U17742 (N_17742,N_10470,N_14916);
nand U17743 (N_17743,N_10285,N_14432);
and U17744 (N_17744,N_12049,N_13846);
nor U17745 (N_17745,N_11183,N_10117);
or U17746 (N_17746,N_14110,N_14947);
xnor U17747 (N_17747,N_13548,N_12244);
nor U17748 (N_17748,N_14884,N_14565);
nand U17749 (N_17749,N_13838,N_14200);
nand U17750 (N_17750,N_12698,N_13536);
xor U17751 (N_17751,N_10774,N_13102);
nand U17752 (N_17752,N_10892,N_14091);
nor U17753 (N_17753,N_13847,N_11287);
nor U17754 (N_17754,N_11416,N_11946);
nor U17755 (N_17755,N_10388,N_10242);
and U17756 (N_17756,N_13886,N_11453);
and U17757 (N_17757,N_14517,N_14598);
and U17758 (N_17758,N_10885,N_10479);
or U17759 (N_17759,N_13706,N_12635);
nor U17760 (N_17760,N_14884,N_12409);
and U17761 (N_17761,N_12774,N_11685);
xnor U17762 (N_17762,N_12347,N_11676);
nor U17763 (N_17763,N_11781,N_13687);
xnor U17764 (N_17764,N_14206,N_12743);
xnor U17765 (N_17765,N_11826,N_13787);
nand U17766 (N_17766,N_11553,N_14331);
xnor U17767 (N_17767,N_11701,N_10034);
xor U17768 (N_17768,N_12922,N_12377);
or U17769 (N_17769,N_11760,N_13263);
and U17770 (N_17770,N_14672,N_14544);
xor U17771 (N_17771,N_10640,N_10230);
or U17772 (N_17772,N_14181,N_12797);
nand U17773 (N_17773,N_10713,N_12391);
or U17774 (N_17774,N_13436,N_11592);
nand U17775 (N_17775,N_10147,N_10855);
or U17776 (N_17776,N_10739,N_11695);
nand U17777 (N_17777,N_14130,N_13230);
nor U17778 (N_17778,N_14305,N_13161);
nand U17779 (N_17779,N_10192,N_14184);
or U17780 (N_17780,N_13758,N_10909);
xnor U17781 (N_17781,N_12489,N_12134);
nand U17782 (N_17782,N_11177,N_12747);
and U17783 (N_17783,N_14135,N_10846);
nor U17784 (N_17784,N_10546,N_14531);
xnor U17785 (N_17785,N_14066,N_12006);
xor U17786 (N_17786,N_10556,N_12473);
or U17787 (N_17787,N_10142,N_10441);
and U17788 (N_17788,N_12313,N_13956);
or U17789 (N_17789,N_11455,N_12291);
and U17790 (N_17790,N_13226,N_14483);
xnor U17791 (N_17791,N_13073,N_11097);
nor U17792 (N_17792,N_11385,N_11174);
and U17793 (N_17793,N_10577,N_11414);
nand U17794 (N_17794,N_10779,N_14243);
or U17795 (N_17795,N_13650,N_11029);
nor U17796 (N_17796,N_12536,N_11884);
nand U17797 (N_17797,N_11850,N_14046);
and U17798 (N_17798,N_14371,N_12437);
nor U17799 (N_17799,N_13603,N_13975);
nand U17800 (N_17800,N_10966,N_12671);
and U17801 (N_17801,N_14625,N_10793);
xor U17802 (N_17802,N_11922,N_11578);
nand U17803 (N_17803,N_13974,N_10648);
and U17804 (N_17804,N_13436,N_12912);
xnor U17805 (N_17805,N_12312,N_10748);
nor U17806 (N_17806,N_12455,N_13471);
nand U17807 (N_17807,N_12800,N_13053);
and U17808 (N_17808,N_10701,N_11818);
nand U17809 (N_17809,N_12852,N_13704);
or U17810 (N_17810,N_10948,N_13648);
and U17811 (N_17811,N_11558,N_11581);
and U17812 (N_17812,N_14083,N_13312);
nor U17813 (N_17813,N_14678,N_14698);
nor U17814 (N_17814,N_10977,N_14257);
nand U17815 (N_17815,N_13832,N_11180);
or U17816 (N_17816,N_10880,N_12844);
or U17817 (N_17817,N_10822,N_10223);
or U17818 (N_17818,N_11317,N_13496);
nand U17819 (N_17819,N_12654,N_10520);
or U17820 (N_17820,N_11898,N_12551);
nor U17821 (N_17821,N_14587,N_10984);
nand U17822 (N_17822,N_12626,N_10596);
and U17823 (N_17823,N_12202,N_10446);
nor U17824 (N_17824,N_13812,N_10262);
nand U17825 (N_17825,N_11816,N_10079);
nor U17826 (N_17826,N_14121,N_12600);
nor U17827 (N_17827,N_12713,N_13278);
or U17828 (N_17828,N_14168,N_13560);
nor U17829 (N_17829,N_14595,N_13177);
xor U17830 (N_17830,N_14973,N_10618);
nand U17831 (N_17831,N_11411,N_14355);
and U17832 (N_17832,N_11867,N_10364);
nand U17833 (N_17833,N_11596,N_14296);
xnor U17834 (N_17834,N_11060,N_13894);
nand U17835 (N_17835,N_14963,N_13365);
or U17836 (N_17836,N_10312,N_14828);
xnor U17837 (N_17837,N_14710,N_13178);
or U17838 (N_17838,N_11505,N_13483);
and U17839 (N_17839,N_14454,N_12767);
or U17840 (N_17840,N_11816,N_11288);
nand U17841 (N_17841,N_11166,N_12765);
xnor U17842 (N_17842,N_14103,N_14439);
nor U17843 (N_17843,N_10004,N_13997);
nand U17844 (N_17844,N_13053,N_11887);
nand U17845 (N_17845,N_12518,N_10851);
nor U17846 (N_17846,N_14084,N_14351);
nor U17847 (N_17847,N_14763,N_10815);
xnor U17848 (N_17848,N_11108,N_14982);
or U17849 (N_17849,N_12633,N_11923);
and U17850 (N_17850,N_12105,N_13600);
or U17851 (N_17851,N_14436,N_13640);
xnor U17852 (N_17852,N_14276,N_10324);
nand U17853 (N_17853,N_14839,N_13128);
or U17854 (N_17854,N_10508,N_13890);
nor U17855 (N_17855,N_10620,N_13468);
nand U17856 (N_17856,N_10267,N_13511);
xor U17857 (N_17857,N_12485,N_11339);
nor U17858 (N_17858,N_12043,N_14512);
or U17859 (N_17859,N_11276,N_13750);
xnor U17860 (N_17860,N_13939,N_10239);
nor U17861 (N_17861,N_12460,N_12816);
xnor U17862 (N_17862,N_10398,N_11246);
nor U17863 (N_17863,N_12157,N_10487);
nand U17864 (N_17864,N_13012,N_14902);
nor U17865 (N_17865,N_14583,N_11197);
or U17866 (N_17866,N_14489,N_11329);
or U17867 (N_17867,N_11148,N_13854);
xor U17868 (N_17868,N_13811,N_10490);
xor U17869 (N_17869,N_12655,N_13576);
xor U17870 (N_17870,N_12377,N_14499);
xor U17871 (N_17871,N_14515,N_10565);
xnor U17872 (N_17872,N_12277,N_11979);
nand U17873 (N_17873,N_13424,N_13413);
xor U17874 (N_17874,N_13396,N_12295);
xnor U17875 (N_17875,N_12719,N_10891);
nand U17876 (N_17876,N_14461,N_11449);
xor U17877 (N_17877,N_10162,N_12501);
nor U17878 (N_17878,N_13189,N_13484);
xor U17879 (N_17879,N_11948,N_11404);
or U17880 (N_17880,N_13502,N_10883);
xor U17881 (N_17881,N_13367,N_10206);
nor U17882 (N_17882,N_10849,N_11000);
nor U17883 (N_17883,N_12697,N_14338);
xnor U17884 (N_17884,N_14488,N_11110);
nand U17885 (N_17885,N_12751,N_10857);
xnor U17886 (N_17886,N_12631,N_11650);
and U17887 (N_17887,N_10538,N_11506);
xor U17888 (N_17888,N_11032,N_13068);
or U17889 (N_17889,N_12548,N_11764);
nand U17890 (N_17890,N_14432,N_14772);
nor U17891 (N_17891,N_14626,N_13448);
and U17892 (N_17892,N_10183,N_13759);
or U17893 (N_17893,N_11976,N_12570);
nand U17894 (N_17894,N_11464,N_10769);
xnor U17895 (N_17895,N_13001,N_10297);
xor U17896 (N_17896,N_11410,N_12754);
nand U17897 (N_17897,N_13561,N_13528);
nor U17898 (N_17898,N_12065,N_10835);
nor U17899 (N_17899,N_11331,N_10150);
nand U17900 (N_17900,N_14461,N_13345);
nand U17901 (N_17901,N_12959,N_13872);
and U17902 (N_17902,N_11864,N_12309);
xnor U17903 (N_17903,N_13123,N_13228);
xnor U17904 (N_17904,N_14704,N_12902);
xnor U17905 (N_17905,N_13305,N_11442);
nand U17906 (N_17906,N_14079,N_12520);
xnor U17907 (N_17907,N_12011,N_14567);
and U17908 (N_17908,N_14989,N_12428);
nand U17909 (N_17909,N_10052,N_12733);
and U17910 (N_17910,N_12353,N_13334);
xor U17911 (N_17911,N_14703,N_10189);
and U17912 (N_17912,N_14507,N_10872);
or U17913 (N_17913,N_13736,N_11757);
or U17914 (N_17914,N_12500,N_11956);
and U17915 (N_17915,N_14571,N_14333);
or U17916 (N_17916,N_13558,N_13279);
xnor U17917 (N_17917,N_13566,N_11703);
xor U17918 (N_17918,N_11782,N_12967);
nor U17919 (N_17919,N_13440,N_14624);
nand U17920 (N_17920,N_12796,N_13022);
or U17921 (N_17921,N_10520,N_14673);
nand U17922 (N_17922,N_10145,N_14054);
nand U17923 (N_17923,N_13111,N_11339);
nor U17924 (N_17924,N_14537,N_11542);
nor U17925 (N_17925,N_14742,N_11408);
and U17926 (N_17926,N_11997,N_13537);
nor U17927 (N_17927,N_14095,N_14967);
or U17928 (N_17928,N_12445,N_13733);
nor U17929 (N_17929,N_12665,N_13845);
and U17930 (N_17930,N_14025,N_10379);
and U17931 (N_17931,N_10825,N_14937);
or U17932 (N_17932,N_13648,N_13307);
nand U17933 (N_17933,N_12194,N_14521);
or U17934 (N_17934,N_10464,N_10699);
or U17935 (N_17935,N_10647,N_10723);
nor U17936 (N_17936,N_11891,N_11454);
nor U17937 (N_17937,N_10819,N_12886);
nand U17938 (N_17938,N_11688,N_11904);
nor U17939 (N_17939,N_13217,N_13985);
nand U17940 (N_17940,N_11766,N_10496);
nand U17941 (N_17941,N_13276,N_14107);
or U17942 (N_17942,N_12597,N_12552);
and U17943 (N_17943,N_12120,N_12785);
nor U17944 (N_17944,N_13829,N_11070);
nand U17945 (N_17945,N_14973,N_10896);
nand U17946 (N_17946,N_11629,N_14918);
or U17947 (N_17947,N_14139,N_13345);
xnor U17948 (N_17948,N_10240,N_10802);
xor U17949 (N_17949,N_11740,N_12898);
nor U17950 (N_17950,N_11543,N_10631);
and U17951 (N_17951,N_13527,N_14070);
nand U17952 (N_17952,N_14265,N_11098);
or U17953 (N_17953,N_11020,N_12218);
and U17954 (N_17954,N_14570,N_11698);
xnor U17955 (N_17955,N_10389,N_14396);
nand U17956 (N_17956,N_11743,N_11772);
or U17957 (N_17957,N_10619,N_10630);
and U17958 (N_17958,N_10395,N_13822);
xnor U17959 (N_17959,N_11765,N_12325);
nor U17960 (N_17960,N_14071,N_14648);
xor U17961 (N_17961,N_10657,N_13944);
nor U17962 (N_17962,N_11991,N_14220);
or U17963 (N_17963,N_11178,N_14625);
nor U17964 (N_17964,N_10636,N_14347);
nand U17965 (N_17965,N_12181,N_14729);
nor U17966 (N_17966,N_11149,N_13079);
xor U17967 (N_17967,N_14814,N_13490);
nor U17968 (N_17968,N_11702,N_13785);
and U17969 (N_17969,N_13220,N_12822);
xnor U17970 (N_17970,N_13066,N_12635);
and U17971 (N_17971,N_10275,N_11719);
nand U17972 (N_17972,N_13517,N_12653);
xnor U17973 (N_17973,N_13329,N_12288);
nor U17974 (N_17974,N_14611,N_13034);
nand U17975 (N_17975,N_14163,N_13797);
and U17976 (N_17976,N_10963,N_11989);
and U17977 (N_17977,N_12811,N_10867);
and U17978 (N_17978,N_14404,N_13570);
and U17979 (N_17979,N_11074,N_14566);
and U17980 (N_17980,N_12506,N_14896);
xor U17981 (N_17981,N_13538,N_11337);
nand U17982 (N_17982,N_10871,N_13901);
xor U17983 (N_17983,N_11293,N_14552);
nor U17984 (N_17984,N_13097,N_14790);
and U17985 (N_17985,N_14029,N_11034);
xnor U17986 (N_17986,N_13726,N_12646);
xnor U17987 (N_17987,N_14211,N_14447);
and U17988 (N_17988,N_10201,N_10990);
or U17989 (N_17989,N_11520,N_10600);
or U17990 (N_17990,N_12287,N_14434);
xnor U17991 (N_17991,N_14618,N_10946);
or U17992 (N_17992,N_13430,N_13456);
and U17993 (N_17993,N_10475,N_14423);
or U17994 (N_17994,N_10969,N_10290);
nor U17995 (N_17995,N_10213,N_10977);
and U17996 (N_17996,N_10067,N_13836);
nor U17997 (N_17997,N_14812,N_13482);
and U17998 (N_17998,N_13802,N_11215);
nand U17999 (N_17999,N_14538,N_11858);
and U18000 (N_18000,N_11277,N_13998);
or U18001 (N_18001,N_12963,N_14702);
nand U18002 (N_18002,N_12416,N_10440);
xor U18003 (N_18003,N_10312,N_12395);
or U18004 (N_18004,N_11868,N_11441);
xor U18005 (N_18005,N_14924,N_13562);
nand U18006 (N_18006,N_14788,N_13711);
nor U18007 (N_18007,N_11822,N_10755);
or U18008 (N_18008,N_13549,N_10313);
and U18009 (N_18009,N_12625,N_12614);
or U18010 (N_18010,N_13645,N_11984);
nand U18011 (N_18011,N_11260,N_13483);
or U18012 (N_18012,N_13462,N_12775);
and U18013 (N_18013,N_12323,N_13716);
xnor U18014 (N_18014,N_13877,N_14925);
or U18015 (N_18015,N_12871,N_10647);
nand U18016 (N_18016,N_12104,N_12822);
or U18017 (N_18017,N_11152,N_13891);
and U18018 (N_18018,N_11617,N_14874);
nor U18019 (N_18019,N_13542,N_12286);
nand U18020 (N_18020,N_13732,N_13267);
xnor U18021 (N_18021,N_13650,N_12903);
nor U18022 (N_18022,N_10551,N_13298);
nand U18023 (N_18023,N_10330,N_13136);
xnor U18024 (N_18024,N_12522,N_14160);
or U18025 (N_18025,N_10679,N_14731);
nand U18026 (N_18026,N_13345,N_11840);
and U18027 (N_18027,N_10441,N_10082);
and U18028 (N_18028,N_11754,N_14400);
nand U18029 (N_18029,N_11581,N_11674);
or U18030 (N_18030,N_10791,N_10710);
nor U18031 (N_18031,N_14210,N_12590);
nand U18032 (N_18032,N_10848,N_13924);
nand U18033 (N_18033,N_10467,N_12748);
and U18034 (N_18034,N_13500,N_12637);
or U18035 (N_18035,N_13817,N_11419);
xor U18036 (N_18036,N_12571,N_11916);
nor U18037 (N_18037,N_12092,N_13544);
and U18038 (N_18038,N_10799,N_12739);
or U18039 (N_18039,N_11552,N_14910);
xnor U18040 (N_18040,N_10000,N_14609);
xnor U18041 (N_18041,N_14964,N_12292);
and U18042 (N_18042,N_10263,N_11761);
and U18043 (N_18043,N_10423,N_14223);
or U18044 (N_18044,N_14015,N_11225);
nor U18045 (N_18045,N_14620,N_14743);
nand U18046 (N_18046,N_12502,N_12935);
nor U18047 (N_18047,N_11273,N_10760);
or U18048 (N_18048,N_10278,N_10862);
xnor U18049 (N_18049,N_13986,N_12064);
nand U18050 (N_18050,N_12983,N_12495);
nor U18051 (N_18051,N_10097,N_14973);
nor U18052 (N_18052,N_10214,N_12480);
and U18053 (N_18053,N_11476,N_12913);
nand U18054 (N_18054,N_11849,N_13293);
nand U18055 (N_18055,N_14497,N_13345);
xnor U18056 (N_18056,N_13921,N_11037);
and U18057 (N_18057,N_10008,N_14254);
or U18058 (N_18058,N_12062,N_14105);
xnor U18059 (N_18059,N_11520,N_12666);
and U18060 (N_18060,N_12201,N_12640);
xor U18061 (N_18061,N_10213,N_10003);
or U18062 (N_18062,N_14597,N_14053);
or U18063 (N_18063,N_10887,N_10919);
nand U18064 (N_18064,N_10208,N_12387);
or U18065 (N_18065,N_14797,N_14907);
or U18066 (N_18066,N_12323,N_14585);
nor U18067 (N_18067,N_12144,N_14076);
nor U18068 (N_18068,N_13448,N_14351);
xor U18069 (N_18069,N_13683,N_12234);
xor U18070 (N_18070,N_12603,N_14358);
nand U18071 (N_18071,N_13147,N_11339);
and U18072 (N_18072,N_14635,N_10710);
nand U18073 (N_18073,N_11951,N_11997);
or U18074 (N_18074,N_13920,N_13075);
xor U18075 (N_18075,N_11654,N_14969);
xor U18076 (N_18076,N_11781,N_14470);
xnor U18077 (N_18077,N_14027,N_11708);
nand U18078 (N_18078,N_10381,N_10962);
xnor U18079 (N_18079,N_12957,N_10553);
nor U18080 (N_18080,N_14197,N_10458);
or U18081 (N_18081,N_14108,N_14770);
nor U18082 (N_18082,N_12969,N_13142);
xnor U18083 (N_18083,N_11819,N_12085);
xor U18084 (N_18084,N_10274,N_11421);
and U18085 (N_18085,N_11958,N_14288);
nor U18086 (N_18086,N_10024,N_11345);
xor U18087 (N_18087,N_12425,N_10229);
xnor U18088 (N_18088,N_11394,N_11045);
or U18089 (N_18089,N_11256,N_14408);
or U18090 (N_18090,N_11592,N_11902);
and U18091 (N_18091,N_13394,N_10171);
xor U18092 (N_18092,N_13557,N_14341);
nor U18093 (N_18093,N_14880,N_12016);
nand U18094 (N_18094,N_13746,N_13552);
nor U18095 (N_18095,N_14147,N_13563);
xnor U18096 (N_18096,N_11686,N_12589);
nand U18097 (N_18097,N_11344,N_13279);
and U18098 (N_18098,N_12480,N_10289);
nor U18099 (N_18099,N_13175,N_12903);
xor U18100 (N_18100,N_14603,N_13283);
nand U18101 (N_18101,N_10151,N_13213);
xnor U18102 (N_18102,N_10938,N_12726);
nand U18103 (N_18103,N_13587,N_14341);
nor U18104 (N_18104,N_11715,N_13976);
and U18105 (N_18105,N_13399,N_11621);
and U18106 (N_18106,N_12381,N_10884);
and U18107 (N_18107,N_13633,N_14863);
xnor U18108 (N_18108,N_14082,N_10779);
nor U18109 (N_18109,N_10535,N_12481);
xnor U18110 (N_18110,N_12120,N_14299);
nor U18111 (N_18111,N_13157,N_10325);
nand U18112 (N_18112,N_13206,N_13216);
nand U18113 (N_18113,N_11820,N_13059);
xnor U18114 (N_18114,N_14180,N_11319);
or U18115 (N_18115,N_10328,N_14504);
xnor U18116 (N_18116,N_12770,N_14608);
or U18117 (N_18117,N_13358,N_13431);
or U18118 (N_18118,N_13296,N_10772);
nor U18119 (N_18119,N_13188,N_11428);
and U18120 (N_18120,N_10234,N_14575);
nand U18121 (N_18121,N_11643,N_11857);
nor U18122 (N_18122,N_14792,N_12667);
nand U18123 (N_18123,N_12715,N_13214);
nor U18124 (N_18124,N_12450,N_14358);
and U18125 (N_18125,N_13170,N_11589);
nand U18126 (N_18126,N_14836,N_13463);
and U18127 (N_18127,N_12140,N_12914);
nor U18128 (N_18128,N_10013,N_12481);
xnor U18129 (N_18129,N_10418,N_12223);
nand U18130 (N_18130,N_13954,N_10473);
or U18131 (N_18131,N_13624,N_10957);
nor U18132 (N_18132,N_10120,N_12640);
or U18133 (N_18133,N_10858,N_11532);
and U18134 (N_18134,N_10728,N_14697);
nand U18135 (N_18135,N_13009,N_14170);
nor U18136 (N_18136,N_11886,N_13201);
nand U18137 (N_18137,N_14341,N_11815);
nor U18138 (N_18138,N_10361,N_14729);
and U18139 (N_18139,N_14014,N_11145);
nand U18140 (N_18140,N_11075,N_14960);
or U18141 (N_18141,N_12962,N_11507);
xor U18142 (N_18142,N_12288,N_12958);
or U18143 (N_18143,N_12629,N_11012);
nand U18144 (N_18144,N_11659,N_13487);
or U18145 (N_18145,N_14923,N_13911);
xor U18146 (N_18146,N_10485,N_12571);
nor U18147 (N_18147,N_10978,N_11094);
nor U18148 (N_18148,N_12333,N_14921);
nor U18149 (N_18149,N_11012,N_12685);
xor U18150 (N_18150,N_13650,N_11002);
and U18151 (N_18151,N_13243,N_12279);
nor U18152 (N_18152,N_13085,N_14619);
nor U18153 (N_18153,N_12743,N_13560);
nand U18154 (N_18154,N_11306,N_10251);
and U18155 (N_18155,N_13504,N_13380);
xor U18156 (N_18156,N_12831,N_13500);
nor U18157 (N_18157,N_14851,N_14643);
or U18158 (N_18158,N_13964,N_10236);
and U18159 (N_18159,N_11021,N_11775);
or U18160 (N_18160,N_13714,N_13857);
or U18161 (N_18161,N_12307,N_11132);
xor U18162 (N_18162,N_13937,N_10131);
nor U18163 (N_18163,N_12022,N_13805);
xor U18164 (N_18164,N_12213,N_13985);
and U18165 (N_18165,N_10706,N_13523);
nand U18166 (N_18166,N_11368,N_10359);
nand U18167 (N_18167,N_12516,N_14537);
or U18168 (N_18168,N_13693,N_11457);
nor U18169 (N_18169,N_10202,N_12167);
and U18170 (N_18170,N_10398,N_12950);
nand U18171 (N_18171,N_13750,N_10701);
and U18172 (N_18172,N_10251,N_10188);
and U18173 (N_18173,N_13609,N_12323);
or U18174 (N_18174,N_10281,N_14409);
and U18175 (N_18175,N_10892,N_12279);
xnor U18176 (N_18176,N_10118,N_13001);
nand U18177 (N_18177,N_11473,N_11781);
or U18178 (N_18178,N_10913,N_14648);
nor U18179 (N_18179,N_14978,N_13553);
xnor U18180 (N_18180,N_11231,N_14403);
and U18181 (N_18181,N_12049,N_11790);
nor U18182 (N_18182,N_10358,N_10534);
and U18183 (N_18183,N_13785,N_11959);
nand U18184 (N_18184,N_10899,N_13244);
or U18185 (N_18185,N_13513,N_12492);
nor U18186 (N_18186,N_12297,N_10794);
nor U18187 (N_18187,N_13087,N_13182);
and U18188 (N_18188,N_14170,N_11278);
nand U18189 (N_18189,N_14835,N_14533);
nand U18190 (N_18190,N_12243,N_10223);
nand U18191 (N_18191,N_11194,N_13974);
and U18192 (N_18192,N_11910,N_14164);
and U18193 (N_18193,N_12886,N_11819);
nand U18194 (N_18194,N_10144,N_14603);
and U18195 (N_18195,N_10047,N_10064);
and U18196 (N_18196,N_13862,N_11056);
or U18197 (N_18197,N_13882,N_10928);
nand U18198 (N_18198,N_11053,N_13228);
and U18199 (N_18199,N_13644,N_13019);
nand U18200 (N_18200,N_14996,N_12469);
or U18201 (N_18201,N_13921,N_14334);
nand U18202 (N_18202,N_11111,N_10267);
or U18203 (N_18203,N_12916,N_12319);
nand U18204 (N_18204,N_14914,N_14306);
and U18205 (N_18205,N_13869,N_10986);
nor U18206 (N_18206,N_10504,N_14623);
nand U18207 (N_18207,N_14313,N_12118);
nor U18208 (N_18208,N_14296,N_13490);
xor U18209 (N_18209,N_12540,N_12593);
xnor U18210 (N_18210,N_11658,N_11293);
and U18211 (N_18211,N_14024,N_10691);
nand U18212 (N_18212,N_14912,N_12293);
xnor U18213 (N_18213,N_12760,N_14795);
nor U18214 (N_18214,N_14849,N_11052);
nor U18215 (N_18215,N_11083,N_11574);
xor U18216 (N_18216,N_11277,N_14093);
or U18217 (N_18217,N_14425,N_11834);
xor U18218 (N_18218,N_12033,N_13104);
nor U18219 (N_18219,N_11596,N_11735);
xnor U18220 (N_18220,N_14860,N_12235);
nor U18221 (N_18221,N_10293,N_10566);
nand U18222 (N_18222,N_12124,N_14473);
nand U18223 (N_18223,N_12671,N_14868);
and U18224 (N_18224,N_11505,N_11695);
nand U18225 (N_18225,N_10524,N_10875);
nor U18226 (N_18226,N_14008,N_12981);
xor U18227 (N_18227,N_10581,N_14001);
and U18228 (N_18228,N_10548,N_11355);
or U18229 (N_18229,N_14282,N_13361);
nand U18230 (N_18230,N_12374,N_13938);
or U18231 (N_18231,N_11807,N_10782);
nand U18232 (N_18232,N_14856,N_12298);
nor U18233 (N_18233,N_14505,N_13248);
nand U18234 (N_18234,N_14452,N_11901);
xor U18235 (N_18235,N_14432,N_14871);
nor U18236 (N_18236,N_14645,N_11066);
or U18237 (N_18237,N_12764,N_11981);
or U18238 (N_18238,N_13520,N_10104);
xnor U18239 (N_18239,N_14657,N_12841);
nor U18240 (N_18240,N_13238,N_14898);
xnor U18241 (N_18241,N_10426,N_13333);
nor U18242 (N_18242,N_12386,N_14169);
and U18243 (N_18243,N_14110,N_12867);
and U18244 (N_18244,N_13862,N_13821);
xor U18245 (N_18245,N_14457,N_13285);
nand U18246 (N_18246,N_10906,N_12235);
nand U18247 (N_18247,N_10205,N_12043);
or U18248 (N_18248,N_13712,N_12981);
nor U18249 (N_18249,N_12317,N_12427);
nand U18250 (N_18250,N_13337,N_13998);
nor U18251 (N_18251,N_12093,N_10949);
xor U18252 (N_18252,N_10141,N_12910);
xnor U18253 (N_18253,N_11492,N_13706);
nand U18254 (N_18254,N_11783,N_13566);
nand U18255 (N_18255,N_11319,N_13068);
and U18256 (N_18256,N_13646,N_12035);
nand U18257 (N_18257,N_14572,N_10711);
or U18258 (N_18258,N_10046,N_14272);
nand U18259 (N_18259,N_12499,N_10115);
and U18260 (N_18260,N_12194,N_14411);
nor U18261 (N_18261,N_10138,N_12363);
or U18262 (N_18262,N_14685,N_14688);
nor U18263 (N_18263,N_12990,N_12478);
xor U18264 (N_18264,N_14227,N_12421);
nand U18265 (N_18265,N_12204,N_10395);
or U18266 (N_18266,N_14971,N_13789);
xnor U18267 (N_18267,N_14074,N_11956);
or U18268 (N_18268,N_11032,N_13605);
or U18269 (N_18269,N_12661,N_12884);
nor U18270 (N_18270,N_10505,N_11088);
nand U18271 (N_18271,N_11391,N_10998);
or U18272 (N_18272,N_14878,N_11612);
and U18273 (N_18273,N_11591,N_14841);
nand U18274 (N_18274,N_10085,N_12427);
or U18275 (N_18275,N_10278,N_12211);
and U18276 (N_18276,N_12529,N_12029);
nor U18277 (N_18277,N_11579,N_11458);
or U18278 (N_18278,N_10882,N_14757);
xor U18279 (N_18279,N_14433,N_11038);
nor U18280 (N_18280,N_10890,N_10619);
xnor U18281 (N_18281,N_10981,N_11306);
and U18282 (N_18282,N_10678,N_11686);
nor U18283 (N_18283,N_14870,N_12282);
xnor U18284 (N_18284,N_14385,N_10849);
or U18285 (N_18285,N_10374,N_10525);
nor U18286 (N_18286,N_10780,N_12065);
nand U18287 (N_18287,N_12944,N_10105);
and U18288 (N_18288,N_14988,N_14044);
nor U18289 (N_18289,N_11311,N_10399);
nand U18290 (N_18290,N_12596,N_14657);
xor U18291 (N_18291,N_14528,N_10731);
nor U18292 (N_18292,N_14135,N_10246);
nand U18293 (N_18293,N_12525,N_10071);
or U18294 (N_18294,N_13118,N_10718);
nor U18295 (N_18295,N_11784,N_13679);
nor U18296 (N_18296,N_14385,N_14979);
or U18297 (N_18297,N_11812,N_12120);
and U18298 (N_18298,N_14533,N_12290);
or U18299 (N_18299,N_12658,N_12586);
and U18300 (N_18300,N_11373,N_11385);
xnor U18301 (N_18301,N_14723,N_12216);
nor U18302 (N_18302,N_12077,N_14715);
or U18303 (N_18303,N_13181,N_13944);
and U18304 (N_18304,N_13618,N_11780);
nand U18305 (N_18305,N_10834,N_13398);
xnor U18306 (N_18306,N_10036,N_14382);
and U18307 (N_18307,N_10241,N_10211);
and U18308 (N_18308,N_10452,N_13105);
nand U18309 (N_18309,N_11647,N_11719);
or U18310 (N_18310,N_13703,N_10608);
and U18311 (N_18311,N_14002,N_10910);
xor U18312 (N_18312,N_12990,N_12663);
or U18313 (N_18313,N_12410,N_14975);
and U18314 (N_18314,N_13344,N_13909);
xnor U18315 (N_18315,N_11643,N_12841);
and U18316 (N_18316,N_12748,N_13306);
and U18317 (N_18317,N_10724,N_13192);
or U18318 (N_18318,N_10021,N_13411);
nand U18319 (N_18319,N_12516,N_12831);
xnor U18320 (N_18320,N_10549,N_12222);
xor U18321 (N_18321,N_11955,N_10450);
nand U18322 (N_18322,N_10361,N_11218);
or U18323 (N_18323,N_11273,N_11038);
and U18324 (N_18324,N_12449,N_13694);
nor U18325 (N_18325,N_14103,N_12638);
nor U18326 (N_18326,N_11990,N_10332);
nor U18327 (N_18327,N_11509,N_11336);
nor U18328 (N_18328,N_14482,N_11575);
nor U18329 (N_18329,N_12793,N_10957);
and U18330 (N_18330,N_13082,N_12125);
nor U18331 (N_18331,N_10571,N_12582);
nor U18332 (N_18332,N_13827,N_11801);
or U18333 (N_18333,N_13826,N_10605);
or U18334 (N_18334,N_14950,N_13620);
and U18335 (N_18335,N_11013,N_12412);
xnor U18336 (N_18336,N_13474,N_10214);
nor U18337 (N_18337,N_12835,N_14748);
nand U18338 (N_18338,N_11672,N_13119);
and U18339 (N_18339,N_13040,N_12523);
and U18340 (N_18340,N_12908,N_12473);
nor U18341 (N_18341,N_10990,N_11652);
nor U18342 (N_18342,N_13411,N_14450);
and U18343 (N_18343,N_13705,N_12288);
or U18344 (N_18344,N_13805,N_10542);
nor U18345 (N_18345,N_12105,N_10333);
xnor U18346 (N_18346,N_11166,N_14379);
xor U18347 (N_18347,N_14384,N_13413);
xor U18348 (N_18348,N_13571,N_12102);
nor U18349 (N_18349,N_13848,N_10840);
xnor U18350 (N_18350,N_11707,N_11005);
nor U18351 (N_18351,N_10398,N_14705);
nand U18352 (N_18352,N_13061,N_12968);
xor U18353 (N_18353,N_11025,N_10505);
nand U18354 (N_18354,N_11512,N_14643);
nor U18355 (N_18355,N_11024,N_12022);
and U18356 (N_18356,N_13555,N_13469);
nor U18357 (N_18357,N_11955,N_11800);
xnor U18358 (N_18358,N_13484,N_10808);
and U18359 (N_18359,N_13670,N_12483);
nor U18360 (N_18360,N_10999,N_12771);
or U18361 (N_18361,N_14424,N_12052);
and U18362 (N_18362,N_12603,N_12753);
nand U18363 (N_18363,N_13838,N_13320);
or U18364 (N_18364,N_11708,N_11648);
and U18365 (N_18365,N_13865,N_10367);
xor U18366 (N_18366,N_14878,N_13663);
or U18367 (N_18367,N_12820,N_11031);
xnor U18368 (N_18368,N_11852,N_11670);
nor U18369 (N_18369,N_13654,N_14102);
and U18370 (N_18370,N_10199,N_13012);
or U18371 (N_18371,N_10455,N_10338);
and U18372 (N_18372,N_11469,N_13572);
nand U18373 (N_18373,N_10619,N_12630);
and U18374 (N_18374,N_14211,N_12174);
or U18375 (N_18375,N_12792,N_10951);
or U18376 (N_18376,N_10852,N_12115);
and U18377 (N_18377,N_14564,N_10286);
nor U18378 (N_18378,N_14444,N_11999);
and U18379 (N_18379,N_14842,N_11234);
xnor U18380 (N_18380,N_12042,N_12045);
nor U18381 (N_18381,N_14069,N_10794);
nand U18382 (N_18382,N_11342,N_13688);
or U18383 (N_18383,N_13603,N_14322);
and U18384 (N_18384,N_12657,N_14992);
nor U18385 (N_18385,N_12429,N_13866);
nand U18386 (N_18386,N_13457,N_11186);
xnor U18387 (N_18387,N_14896,N_13489);
xnor U18388 (N_18388,N_11537,N_12724);
nor U18389 (N_18389,N_14394,N_13478);
and U18390 (N_18390,N_13791,N_11784);
xor U18391 (N_18391,N_11901,N_13159);
nor U18392 (N_18392,N_12650,N_10761);
or U18393 (N_18393,N_12766,N_11854);
and U18394 (N_18394,N_11814,N_12549);
nand U18395 (N_18395,N_11209,N_10173);
or U18396 (N_18396,N_10324,N_14099);
or U18397 (N_18397,N_14818,N_14809);
nor U18398 (N_18398,N_13854,N_11105);
and U18399 (N_18399,N_11504,N_12565);
nor U18400 (N_18400,N_12832,N_14215);
nor U18401 (N_18401,N_14958,N_11324);
xor U18402 (N_18402,N_12347,N_12836);
xnor U18403 (N_18403,N_11691,N_14422);
xor U18404 (N_18404,N_14980,N_13759);
nor U18405 (N_18405,N_14223,N_14597);
and U18406 (N_18406,N_11556,N_13997);
xor U18407 (N_18407,N_14629,N_11262);
nand U18408 (N_18408,N_14444,N_12796);
nand U18409 (N_18409,N_11301,N_12279);
and U18410 (N_18410,N_12295,N_13970);
nor U18411 (N_18411,N_11930,N_14996);
and U18412 (N_18412,N_10237,N_12062);
nor U18413 (N_18413,N_10162,N_11205);
xor U18414 (N_18414,N_12215,N_14330);
nand U18415 (N_18415,N_11492,N_12640);
nand U18416 (N_18416,N_14989,N_14979);
nand U18417 (N_18417,N_10533,N_10549);
nor U18418 (N_18418,N_12978,N_13018);
or U18419 (N_18419,N_12020,N_11137);
and U18420 (N_18420,N_13256,N_12972);
or U18421 (N_18421,N_11763,N_13117);
and U18422 (N_18422,N_10277,N_14347);
nor U18423 (N_18423,N_14302,N_11605);
or U18424 (N_18424,N_13567,N_13685);
or U18425 (N_18425,N_13115,N_12740);
xor U18426 (N_18426,N_10308,N_13389);
and U18427 (N_18427,N_13744,N_11860);
nand U18428 (N_18428,N_12809,N_11938);
xor U18429 (N_18429,N_13341,N_10417);
xnor U18430 (N_18430,N_14919,N_11082);
nand U18431 (N_18431,N_12640,N_14388);
xor U18432 (N_18432,N_13753,N_12697);
or U18433 (N_18433,N_12971,N_14634);
nand U18434 (N_18434,N_12057,N_11510);
and U18435 (N_18435,N_11657,N_14714);
or U18436 (N_18436,N_12751,N_14865);
xor U18437 (N_18437,N_14255,N_11973);
nor U18438 (N_18438,N_14535,N_10759);
or U18439 (N_18439,N_13089,N_13186);
nor U18440 (N_18440,N_13062,N_14659);
or U18441 (N_18441,N_11058,N_13882);
and U18442 (N_18442,N_14121,N_10129);
and U18443 (N_18443,N_12735,N_12812);
nand U18444 (N_18444,N_11519,N_13156);
or U18445 (N_18445,N_10436,N_14439);
nand U18446 (N_18446,N_11477,N_12462);
and U18447 (N_18447,N_13080,N_10382);
nand U18448 (N_18448,N_13402,N_14219);
and U18449 (N_18449,N_10048,N_13762);
xnor U18450 (N_18450,N_10793,N_11517);
xnor U18451 (N_18451,N_10538,N_10580);
nor U18452 (N_18452,N_14922,N_13400);
nor U18453 (N_18453,N_14831,N_10478);
and U18454 (N_18454,N_14066,N_14283);
xor U18455 (N_18455,N_13009,N_13958);
or U18456 (N_18456,N_14425,N_10170);
or U18457 (N_18457,N_14722,N_10075);
or U18458 (N_18458,N_10503,N_12797);
xnor U18459 (N_18459,N_13214,N_14011);
nand U18460 (N_18460,N_11643,N_11380);
or U18461 (N_18461,N_10992,N_11417);
nand U18462 (N_18462,N_11835,N_14447);
nand U18463 (N_18463,N_12042,N_10034);
or U18464 (N_18464,N_14871,N_11239);
nor U18465 (N_18465,N_11957,N_14205);
nor U18466 (N_18466,N_14184,N_13802);
xor U18467 (N_18467,N_11251,N_10330);
and U18468 (N_18468,N_12032,N_13186);
xor U18469 (N_18469,N_14984,N_11638);
nand U18470 (N_18470,N_12279,N_13193);
xor U18471 (N_18471,N_12954,N_10593);
nor U18472 (N_18472,N_13645,N_13077);
nand U18473 (N_18473,N_10703,N_14052);
and U18474 (N_18474,N_12257,N_12495);
xnor U18475 (N_18475,N_13445,N_11150);
or U18476 (N_18476,N_14700,N_10174);
or U18477 (N_18477,N_12593,N_10818);
nor U18478 (N_18478,N_12893,N_14431);
nor U18479 (N_18479,N_12196,N_13223);
nor U18480 (N_18480,N_11762,N_14955);
xnor U18481 (N_18481,N_13180,N_13913);
and U18482 (N_18482,N_12101,N_11348);
and U18483 (N_18483,N_12701,N_11755);
nor U18484 (N_18484,N_11156,N_11804);
or U18485 (N_18485,N_12825,N_13350);
nand U18486 (N_18486,N_10131,N_12417);
or U18487 (N_18487,N_11538,N_12838);
xor U18488 (N_18488,N_14637,N_11394);
xnor U18489 (N_18489,N_13270,N_10577);
or U18490 (N_18490,N_10627,N_14910);
nand U18491 (N_18491,N_13261,N_14763);
and U18492 (N_18492,N_13203,N_10637);
nand U18493 (N_18493,N_12901,N_10456);
xor U18494 (N_18494,N_13412,N_11753);
xnor U18495 (N_18495,N_11559,N_10823);
and U18496 (N_18496,N_14959,N_12244);
or U18497 (N_18497,N_13304,N_12501);
or U18498 (N_18498,N_11632,N_13945);
nor U18499 (N_18499,N_10048,N_11721);
nor U18500 (N_18500,N_14140,N_13470);
nand U18501 (N_18501,N_14861,N_14469);
and U18502 (N_18502,N_11322,N_14770);
nand U18503 (N_18503,N_14944,N_14118);
xnor U18504 (N_18504,N_11619,N_11227);
xnor U18505 (N_18505,N_10356,N_13318);
and U18506 (N_18506,N_12098,N_14600);
nor U18507 (N_18507,N_11259,N_10333);
or U18508 (N_18508,N_11411,N_12063);
nand U18509 (N_18509,N_13199,N_13147);
nor U18510 (N_18510,N_12065,N_10165);
nand U18511 (N_18511,N_12229,N_10769);
nand U18512 (N_18512,N_12242,N_13059);
xnor U18513 (N_18513,N_14954,N_14966);
xnor U18514 (N_18514,N_11074,N_14985);
xor U18515 (N_18515,N_10120,N_10873);
or U18516 (N_18516,N_10845,N_14027);
and U18517 (N_18517,N_11628,N_10234);
nor U18518 (N_18518,N_12156,N_13988);
nand U18519 (N_18519,N_12923,N_12569);
or U18520 (N_18520,N_12187,N_13335);
nor U18521 (N_18521,N_12407,N_12188);
or U18522 (N_18522,N_12257,N_11074);
nor U18523 (N_18523,N_13230,N_10283);
nand U18524 (N_18524,N_11859,N_10884);
and U18525 (N_18525,N_10995,N_11915);
and U18526 (N_18526,N_12030,N_14204);
xor U18527 (N_18527,N_14515,N_11625);
nor U18528 (N_18528,N_14743,N_12740);
or U18529 (N_18529,N_11311,N_14172);
or U18530 (N_18530,N_10275,N_14061);
and U18531 (N_18531,N_14544,N_13006);
xnor U18532 (N_18532,N_12335,N_13880);
or U18533 (N_18533,N_13062,N_13584);
xnor U18534 (N_18534,N_11896,N_14637);
xnor U18535 (N_18535,N_10954,N_11079);
xor U18536 (N_18536,N_12525,N_11715);
nand U18537 (N_18537,N_10151,N_10958);
and U18538 (N_18538,N_13987,N_11586);
nor U18539 (N_18539,N_13967,N_12330);
xnor U18540 (N_18540,N_10121,N_13472);
or U18541 (N_18541,N_10132,N_14270);
or U18542 (N_18542,N_10365,N_14118);
and U18543 (N_18543,N_11454,N_11332);
nand U18544 (N_18544,N_14661,N_14965);
nand U18545 (N_18545,N_14714,N_10643);
nor U18546 (N_18546,N_12696,N_14677);
nand U18547 (N_18547,N_12165,N_11386);
nand U18548 (N_18548,N_11814,N_10983);
or U18549 (N_18549,N_14671,N_11020);
xnor U18550 (N_18550,N_10824,N_11700);
xor U18551 (N_18551,N_13774,N_13094);
nand U18552 (N_18552,N_14627,N_11421);
nor U18553 (N_18553,N_14548,N_11537);
xnor U18554 (N_18554,N_12424,N_10596);
xnor U18555 (N_18555,N_13676,N_10097);
and U18556 (N_18556,N_14320,N_11948);
nor U18557 (N_18557,N_10904,N_12493);
or U18558 (N_18558,N_14184,N_11027);
nor U18559 (N_18559,N_12674,N_13489);
and U18560 (N_18560,N_14674,N_13081);
or U18561 (N_18561,N_10384,N_14151);
xor U18562 (N_18562,N_13748,N_12961);
nand U18563 (N_18563,N_11300,N_13597);
and U18564 (N_18564,N_14957,N_13368);
nand U18565 (N_18565,N_14542,N_12589);
nor U18566 (N_18566,N_11836,N_12757);
nor U18567 (N_18567,N_13444,N_10257);
nor U18568 (N_18568,N_13267,N_10176);
xnor U18569 (N_18569,N_12527,N_11263);
or U18570 (N_18570,N_13943,N_11894);
and U18571 (N_18571,N_13771,N_10066);
and U18572 (N_18572,N_10077,N_12668);
nand U18573 (N_18573,N_12235,N_10375);
xor U18574 (N_18574,N_13275,N_12218);
nor U18575 (N_18575,N_12231,N_14234);
and U18576 (N_18576,N_12918,N_10036);
and U18577 (N_18577,N_12753,N_14740);
and U18578 (N_18578,N_11095,N_12385);
and U18579 (N_18579,N_11317,N_13137);
xnor U18580 (N_18580,N_11926,N_11025);
nand U18581 (N_18581,N_13184,N_13092);
and U18582 (N_18582,N_11719,N_11001);
and U18583 (N_18583,N_14607,N_11299);
nor U18584 (N_18584,N_11501,N_13465);
xnor U18585 (N_18585,N_13437,N_12965);
nor U18586 (N_18586,N_10176,N_11203);
xnor U18587 (N_18587,N_13242,N_12796);
or U18588 (N_18588,N_10325,N_12923);
nor U18589 (N_18589,N_14508,N_11699);
xor U18590 (N_18590,N_13589,N_13212);
xnor U18591 (N_18591,N_12212,N_10319);
xor U18592 (N_18592,N_13172,N_11048);
nor U18593 (N_18593,N_13773,N_13265);
and U18594 (N_18594,N_11156,N_10882);
and U18595 (N_18595,N_14619,N_14275);
xnor U18596 (N_18596,N_13608,N_14604);
and U18597 (N_18597,N_14417,N_12374);
xor U18598 (N_18598,N_12156,N_14537);
or U18599 (N_18599,N_14702,N_12503);
nor U18600 (N_18600,N_12114,N_11600);
nand U18601 (N_18601,N_12905,N_14509);
nor U18602 (N_18602,N_10222,N_14044);
xnor U18603 (N_18603,N_10348,N_11321);
and U18604 (N_18604,N_14442,N_12923);
nor U18605 (N_18605,N_11192,N_12837);
nor U18606 (N_18606,N_12513,N_13230);
nand U18607 (N_18607,N_10186,N_14747);
nor U18608 (N_18608,N_14308,N_13104);
and U18609 (N_18609,N_11604,N_13218);
xor U18610 (N_18610,N_11775,N_14211);
and U18611 (N_18611,N_13433,N_12798);
and U18612 (N_18612,N_13725,N_14744);
xnor U18613 (N_18613,N_11333,N_10588);
or U18614 (N_18614,N_11888,N_12520);
or U18615 (N_18615,N_12325,N_12040);
or U18616 (N_18616,N_10268,N_10624);
nor U18617 (N_18617,N_10946,N_11810);
xor U18618 (N_18618,N_10857,N_12510);
nor U18619 (N_18619,N_10175,N_10003);
xor U18620 (N_18620,N_12435,N_11222);
or U18621 (N_18621,N_12353,N_14707);
nor U18622 (N_18622,N_10276,N_13421);
xor U18623 (N_18623,N_10992,N_14461);
nand U18624 (N_18624,N_14059,N_12885);
nor U18625 (N_18625,N_13674,N_13305);
nor U18626 (N_18626,N_14292,N_14343);
xor U18627 (N_18627,N_10871,N_14620);
nand U18628 (N_18628,N_12768,N_11381);
nor U18629 (N_18629,N_11403,N_14831);
or U18630 (N_18630,N_12947,N_14201);
and U18631 (N_18631,N_10543,N_12821);
xnor U18632 (N_18632,N_14489,N_12897);
or U18633 (N_18633,N_11780,N_13685);
and U18634 (N_18634,N_13988,N_14590);
and U18635 (N_18635,N_11748,N_10940);
or U18636 (N_18636,N_13505,N_12184);
nor U18637 (N_18637,N_11428,N_10156);
nor U18638 (N_18638,N_13996,N_14518);
or U18639 (N_18639,N_12299,N_10544);
and U18640 (N_18640,N_10427,N_13179);
nor U18641 (N_18641,N_11497,N_10878);
nor U18642 (N_18642,N_11555,N_13044);
xnor U18643 (N_18643,N_11096,N_13344);
or U18644 (N_18644,N_11213,N_12951);
or U18645 (N_18645,N_12582,N_11548);
or U18646 (N_18646,N_14608,N_12452);
nor U18647 (N_18647,N_11431,N_11562);
nand U18648 (N_18648,N_14876,N_13063);
and U18649 (N_18649,N_10336,N_14352);
xor U18650 (N_18650,N_10286,N_14850);
or U18651 (N_18651,N_14451,N_12448);
nor U18652 (N_18652,N_10915,N_13304);
xor U18653 (N_18653,N_10984,N_12398);
nor U18654 (N_18654,N_14725,N_14789);
or U18655 (N_18655,N_10427,N_12468);
nand U18656 (N_18656,N_10083,N_14949);
or U18657 (N_18657,N_12437,N_12169);
xor U18658 (N_18658,N_10564,N_11521);
and U18659 (N_18659,N_13952,N_13914);
and U18660 (N_18660,N_14907,N_14516);
nand U18661 (N_18661,N_12970,N_12257);
nand U18662 (N_18662,N_13173,N_14737);
nor U18663 (N_18663,N_10353,N_13744);
and U18664 (N_18664,N_13701,N_12673);
nor U18665 (N_18665,N_12333,N_12304);
nor U18666 (N_18666,N_13749,N_11089);
nor U18667 (N_18667,N_12439,N_11471);
and U18668 (N_18668,N_11028,N_12410);
xor U18669 (N_18669,N_13327,N_12698);
and U18670 (N_18670,N_11390,N_11811);
and U18671 (N_18671,N_10829,N_10583);
nand U18672 (N_18672,N_13403,N_10075);
nor U18673 (N_18673,N_10603,N_14327);
nor U18674 (N_18674,N_12274,N_11498);
or U18675 (N_18675,N_11492,N_12816);
and U18676 (N_18676,N_14504,N_11981);
or U18677 (N_18677,N_10719,N_11332);
nor U18678 (N_18678,N_13301,N_14939);
and U18679 (N_18679,N_14906,N_13084);
nor U18680 (N_18680,N_11109,N_11631);
or U18681 (N_18681,N_12802,N_14299);
or U18682 (N_18682,N_10680,N_14759);
nand U18683 (N_18683,N_12670,N_13621);
and U18684 (N_18684,N_11003,N_13905);
nor U18685 (N_18685,N_13995,N_10080);
and U18686 (N_18686,N_10670,N_12877);
and U18687 (N_18687,N_11577,N_11970);
nor U18688 (N_18688,N_14509,N_11079);
and U18689 (N_18689,N_13235,N_11981);
and U18690 (N_18690,N_13913,N_13662);
nand U18691 (N_18691,N_10827,N_12060);
and U18692 (N_18692,N_11585,N_11937);
and U18693 (N_18693,N_14183,N_11365);
xor U18694 (N_18694,N_10721,N_10589);
nand U18695 (N_18695,N_13939,N_10988);
nand U18696 (N_18696,N_13633,N_14490);
or U18697 (N_18697,N_11270,N_10822);
xor U18698 (N_18698,N_12073,N_11501);
xnor U18699 (N_18699,N_14330,N_12650);
or U18700 (N_18700,N_10925,N_12369);
nor U18701 (N_18701,N_14029,N_14858);
nor U18702 (N_18702,N_14257,N_11362);
or U18703 (N_18703,N_14548,N_11346);
and U18704 (N_18704,N_12261,N_13902);
xor U18705 (N_18705,N_13134,N_11706);
and U18706 (N_18706,N_11914,N_11850);
nand U18707 (N_18707,N_10159,N_14492);
and U18708 (N_18708,N_12477,N_13178);
and U18709 (N_18709,N_12116,N_11617);
nand U18710 (N_18710,N_10059,N_14567);
nor U18711 (N_18711,N_13691,N_14614);
xor U18712 (N_18712,N_14681,N_10806);
and U18713 (N_18713,N_11948,N_13983);
and U18714 (N_18714,N_10035,N_12957);
or U18715 (N_18715,N_10171,N_12372);
nor U18716 (N_18716,N_13934,N_11823);
nand U18717 (N_18717,N_11541,N_11600);
xor U18718 (N_18718,N_14954,N_13982);
xor U18719 (N_18719,N_12930,N_10974);
xor U18720 (N_18720,N_10706,N_10412);
nor U18721 (N_18721,N_13842,N_14661);
xnor U18722 (N_18722,N_13518,N_14406);
and U18723 (N_18723,N_12249,N_10694);
nand U18724 (N_18724,N_10304,N_13916);
and U18725 (N_18725,N_11040,N_11578);
nand U18726 (N_18726,N_12478,N_13225);
nand U18727 (N_18727,N_12920,N_14298);
nor U18728 (N_18728,N_10171,N_13183);
nor U18729 (N_18729,N_12382,N_10342);
and U18730 (N_18730,N_13172,N_12029);
nor U18731 (N_18731,N_11445,N_13282);
xnor U18732 (N_18732,N_10119,N_10678);
xor U18733 (N_18733,N_12797,N_13168);
nand U18734 (N_18734,N_14342,N_10862);
nand U18735 (N_18735,N_10181,N_12747);
xnor U18736 (N_18736,N_13813,N_11920);
xnor U18737 (N_18737,N_13518,N_12762);
or U18738 (N_18738,N_13469,N_11532);
nand U18739 (N_18739,N_11159,N_13593);
or U18740 (N_18740,N_11456,N_13371);
nand U18741 (N_18741,N_12976,N_10063);
xnor U18742 (N_18742,N_13407,N_10677);
nor U18743 (N_18743,N_11832,N_12600);
nand U18744 (N_18744,N_11157,N_13095);
or U18745 (N_18745,N_14990,N_11134);
nor U18746 (N_18746,N_13711,N_14536);
nand U18747 (N_18747,N_13344,N_12653);
xnor U18748 (N_18748,N_10989,N_14568);
and U18749 (N_18749,N_10438,N_10900);
nand U18750 (N_18750,N_14464,N_11888);
nand U18751 (N_18751,N_12593,N_12761);
or U18752 (N_18752,N_10948,N_11080);
xnor U18753 (N_18753,N_14213,N_10064);
nand U18754 (N_18754,N_14362,N_10334);
nor U18755 (N_18755,N_11464,N_12328);
nand U18756 (N_18756,N_10832,N_12958);
nor U18757 (N_18757,N_10461,N_12790);
and U18758 (N_18758,N_14389,N_13594);
nor U18759 (N_18759,N_12014,N_11374);
xnor U18760 (N_18760,N_12697,N_10968);
and U18761 (N_18761,N_10991,N_13727);
or U18762 (N_18762,N_11439,N_11503);
nor U18763 (N_18763,N_13109,N_13070);
or U18764 (N_18764,N_10237,N_11925);
nor U18765 (N_18765,N_11790,N_10964);
nand U18766 (N_18766,N_11361,N_14894);
and U18767 (N_18767,N_12322,N_13440);
nor U18768 (N_18768,N_13859,N_12053);
or U18769 (N_18769,N_14324,N_14068);
xor U18770 (N_18770,N_13837,N_14577);
and U18771 (N_18771,N_12760,N_12892);
nand U18772 (N_18772,N_12562,N_14752);
nor U18773 (N_18773,N_14821,N_12626);
xnor U18774 (N_18774,N_10574,N_12819);
xnor U18775 (N_18775,N_10289,N_11469);
xnor U18776 (N_18776,N_10539,N_11527);
or U18777 (N_18777,N_13736,N_12214);
nand U18778 (N_18778,N_11189,N_12213);
nand U18779 (N_18779,N_11586,N_13800);
and U18780 (N_18780,N_12331,N_12477);
or U18781 (N_18781,N_14817,N_14713);
nor U18782 (N_18782,N_13744,N_10703);
nand U18783 (N_18783,N_10444,N_10035);
and U18784 (N_18784,N_12799,N_10450);
nand U18785 (N_18785,N_13892,N_11709);
xor U18786 (N_18786,N_12978,N_10056);
xnor U18787 (N_18787,N_14919,N_11909);
or U18788 (N_18788,N_12057,N_13617);
nor U18789 (N_18789,N_13199,N_14715);
nand U18790 (N_18790,N_11602,N_11844);
or U18791 (N_18791,N_11971,N_12131);
and U18792 (N_18792,N_14118,N_13886);
nor U18793 (N_18793,N_10133,N_11057);
nor U18794 (N_18794,N_14588,N_11389);
nand U18795 (N_18795,N_14998,N_11418);
nor U18796 (N_18796,N_11498,N_13518);
or U18797 (N_18797,N_12277,N_11474);
and U18798 (N_18798,N_13174,N_11554);
xor U18799 (N_18799,N_14464,N_11388);
xnor U18800 (N_18800,N_13511,N_10075);
or U18801 (N_18801,N_12057,N_13857);
nand U18802 (N_18802,N_13512,N_10978);
nor U18803 (N_18803,N_14928,N_12611);
nor U18804 (N_18804,N_10660,N_10187);
nand U18805 (N_18805,N_14593,N_14351);
and U18806 (N_18806,N_13743,N_10276);
xor U18807 (N_18807,N_13197,N_12311);
xnor U18808 (N_18808,N_11850,N_12786);
xor U18809 (N_18809,N_14985,N_12764);
nand U18810 (N_18810,N_14382,N_11734);
or U18811 (N_18811,N_10545,N_12971);
nand U18812 (N_18812,N_10553,N_14515);
or U18813 (N_18813,N_12561,N_10460);
nor U18814 (N_18814,N_11969,N_10865);
xor U18815 (N_18815,N_11646,N_11559);
xnor U18816 (N_18816,N_10700,N_11495);
or U18817 (N_18817,N_11844,N_14844);
nor U18818 (N_18818,N_12577,N_14880);
or U18819 (N_18819,N_11995,N_12802);
nor U18820 (N_18820,N_10141,N_11432);
and U18821 (N_18821,N_10702,N_14718);
and U18822 (N_18822,N_12435,N_10184);
nand U18823 (N_18823,N_10451,N_10745);
xnor U18824 (N_18824,N_12800,N_13511);
nor U18825 (N_18825,N_10357,N_10513);
and U18826 (N_18826,N_12999,N_12683);
nand U18827 (N_18827,N_10618,N_14763);
xor U18828 (N_18828,N_13381,N_11595);
or U18829 (N_18829,N_14529,N_14680);
or U18830 (N_18830,N_10828,N_14728);
and U18831 (N_18831,N_13413,N_11172);
xor U18832 (N_18832,N_12804,N_11209);
and U18833 (N_18833,N_11238,N_10186);
nand U18834 (N_18834,N_13013,N_13907);
and U18835 (N_18835,N_11918,N_11764);
xor U18836 (N_18836,N_14779,N_11842);
nand U18837 (N_18837,N_11859,N_11305);
and U18838 (N_18838,N_13642,N_13551);
nor U18839 (N_18839,N_13060,N_11235);
nor U18840 (N_18840,N_11047,N_12872);
xnor U18841 (N_18841,N_13109,N_12806);
nor U18842 (N_18842,N_13451,N_14310);
nand U18843 (N_18843,N_10342,N_13476);
xnor U18844 (N_18844,N_11544,N_13288);
nor U18845 (N_18845,N_11620,N_14559);
nand U18846 (N_18846,N_11815,N_12878);
nor U18847 (N_18847,N_13252,N_14377);
nand U18848 (N_18848,N_11258,N_10093);
nor U18849 (N_18849,N_11782,N_12939);
nor U18850 (N_18850,N_11954,N_13353);
and U18851 (N_18851,N_12810,N_14742);
xor U18852 (N_18852,N_12267,N_14660);
nand U18853 (N_18853,N_11925,N_12371);
nor U18854 (N_18854,N_14984,N_14287);
nand U18855 (N_18855,N_12498,N_13893);
and U18856 (N_18856,N_12713,N_10806);
or U18857 (N_18857,N_13510,N_10076);
and U18858 (N_18858,N_10951,N_11298);
and U18859 (N_18859,N_10501,N_10072);
or U18860 (N_18860,N_13196,N_11897);
nor U18861 (N_18861,N_14833,N_11022);
nand U18862 (N_18862,N_12663,N_14698);
xor U18863 (N_18863,N_12121,N_14226);
xnor U18864 (N_18864,N_12402,N_14693);
or U18865 (N_18865,N_12525,N_14056);
or U18866 (N_18866,N_11792,N_13448);
and U18867 (N_18867,N_14269,N_12043);
nand U18868 (N_18868,N_12232,N_11324);
nand U18869 (N_18869,N_13533,N_10346);
or U18870 (N_18870,N_13648,N_11745);
nor U18871 (N_18871,N_14541,N_11894);
nand U18872 (N_18872,N_14405,N_14157);
nor U18873 (N_18873,N_14689,N_12231);
xnor U18874 (N_18874,N_13900,N_13825);
or U18875 (N_18875,N_10867,N_12132);
xor U18876 (N_18876,N_10278,N_14869);
nand U18877 (N_18877,N_10752,N_14194);
nor U18878 (N_18878,N_12907,N_11464);
xor U18879 (N_18879,N_10998,N_11176);
nand U18880 (N_18880,N_13427,N_11818);
xor U18881 (N_18881,N_14087,N_11465);
xor U18882 (N_18882,N_13668,N_12858);
nand U18883 (N_18883,N_10167,N_13856);
nor U18884 (N_18884,N_10292,N_12805);
and U18885 (N_18885,N_11009,N_13600);
nor U18886 (N_18886,N_10887,N_11201);
xor U18887 (N_18887,N_10106,N_13740);
nor U18888 (N_18888,N_10190,N_14400);
or U18889 (N_18889,N_10446,N_10403);
xnor U18890 (N_18890,N_13413,N_11833);
or U18891 (N_18891,N_10594,N_10649);
nor U18892 (N_18892,N_12839,N_14564);
nand U18893 (N_18893,N_14084,N_11617);
and U18894 (N_18894,N_11425,N_11315);
or U18895 (N_18895,N_11763,N_10994);
or U18896 (N_18896,N_11361,N_12159);
and U18897 (N_18897,N_13968,N_13732);
nor U18898 (N_18898,N_11743,N_12689);
nor U18899 (N_18899,N_13722,N_10319);
nor U18900 (N_18900,N_13079,N_12133);
or U18901 (N_18901,N_10710,N_14678);
and U18902 (N_18902,N_10756,N_10956);
nor U18903 (N_18903,N_14991,N_12934);
or U18904 (N_18904,N_11398,N_10484);
and U18905 (N_18905,N_11764,N_10285);
or U18906 (N_18906,N_13491,N_14872);
or U18907 (N_18907,N_11336,N_11330);
nand U18908 (N_18908,N_11540,N_12235);
and U18909 (N_18909,N_13310,N_10305);
and U18910 (N_18910,N_10920,N_10195);
nor U18911 (N_18911,N_14187,N_14273);
nand U18912 (N_18912,N_14121,N_12950);
nand U18913 (N_18913,N_13257,N_13376);
and U18914 (N_18914,N_10488,N_14951);
or U18915 (N_18915,N_11717,N_13557);
nor U18916 (N_18916,N_11524,N_10264);
xor U18917 (N_18917,N_14534,N_11912);
nor U18918 (N_18918,N_13916,N_13574);
nor U18919 (N_18919,N_13988,N_13612);
xor U18920 (N_18920,N_13856,N_10930);
nor U18921 (N_18921,N_11378,N_13901);
nor U18922 (N_18922,N_12189,N_12748);
and U18923 (N_18923,N_13470,N_12439);
nand U18924 (N_18924,N_12444,N_13562);
nor U18925 (N_18925,N_12551,N_11315);
and U18926 (N_18926,N_14583,N_10004);
and U18927 (N_18927,N_10508,N_12803);
and U18928 (N_18928,N_10871,N_12134);
xnor U18929 (N_18929,N_11089,N_12750);
xnor U18930 (N_18930,N_11377,N_13680);
xnor U18931 (N_18931,N_14651,N_10434);
and U18932 (N_18932,N_12017,N_11615);
and U18933 (N_18933,N_11715,N_12753);
or U18934 (N_18934,N_10948,N_13932);
nor U18935 (N_18935,N_10518,N_12167);
and U18936 (N_18936,N_13606,N_10838);
or U18937 (N_18937,N_13590,N_12970);
or U18938 (N_18938,N_13901,N_10267);
xnor U18939 (N_18939,N_14005,N_11733);
and U18940 (N_18940,N_10134,N_11202);
and U18941 (N_18941,N_14655,N_14014);
nor U18942 (N_18942,N_14725,N_14378);
and U18943 (N_18943,N_14383,N_11539);
nand U18944 (N_18944,N_14639,N_13813);
or U18945 (N_18945,N_11978,N_13039);
or U18946 (N_18946,N_10283,N_12534);
nand U18947 (N_18947,N_13908,N_10143);
and U18948 (N_18948,N_10347,N_14546);
nor U18949 (N_18949,N_14977,N_14380);
and U18950 (N_18950,N_10576,N_11000);
or U18951 (N_18951,N_13460,N_14063);
and U18952 (N_18952,N_10524,N_12939);
and U18953 (N_18953,N_11746,N_10615);
nor U18954 (N_18954,N_14505,N_12335);
and U18955 (N_18955,N_11404,N_14967);
nand U18956 (N_18956,N_12955,N_10346);
or U18957 (N_18957,N_10603,N_14806);
nor U18958 (N_18958,N_12045,N_11467);
nor U18959 (N_18959,N_12030,N_11603);
or U18960 (N_18960,N_13500,N_11597);
and U18961 (N_18961,N_14690,N_12839);
nand U18962 (N_18962,N_10421,N_10962);
xor U18963 (N_18963,N_14342,N_10695);
or U18964 (N_18964,N_13948,N_12150);
nor U18965 (N_18965,N_12173,N_12584);
nor U18966 (N_18966,N_14351,N_11586);
and U18967 (N_18967,N_11278,N_10953);
nor U18968 (N_18968,N_12925,N_12428);
or U18969 (N_18969,N_13012,N_11631);
or U18970 (N_18970,N_13318,N_13593);
nand U18971 (N_18971,N_11412,N_14283);
and U18972 (N_18972,N_14581,N_11386);
nand U18973 (N_18973,N_11907,N_12198);
and U18974 (N_18974,N_13790,N_12909);
nor U18975 (N_18975,N_10304,N_14204);
nor U18976 (N_18976,N_10279,N_10150);
nand U18977 (N_18977,N_12572,N_10957);
and U18978 (N_18978,N_10430,N_10934);
and U18979 (N_18979,N_12255,N_12512);
xnor U18980 (N_18980,N_12302,N_13216);
xnor U18981 (N_18981,N_12202,N_11686);
nand U18982 (N_18982,N_11426,N_14146);
xor U18983 (N_18983,N_10030,N_14164);
nand U18984 (N_18984,N_14540,N_14390);
and U18985 (N_18985,N_14260,N_10824);
xnor U18986 (N_18986,N_11797,N_14683);
and U18987 (N_18987,N_12250,N_14322);
xor U18988 (N_18988,N_13514,N_13225);
and U18989 (N_18989,N_10250,N_12659);
or U18990 (N_18990,N_14855,N_12380);
xnor U18991 (N_18991,N_11845,N_12600);
and U18992 (N_18992,N_10909,N_14733);
and U18993 (N_18993,N_12258,N_14565);
xnor U18994 (N_18994,N_11688,N_12908);
nand U18995 (N_18995,N_13366,N_11281);
or U18996 (N_18996,N_14905,N_14899);
xnor U18997 (N_18997,N_13797,N_13751);
nor U18998 (N_18998,N_12720,N_11868);
or U18999 (N_18999,N_12422,N_11445);
xnor U19000 (N_19000,N_12238,N_11442);
nor U19001 (N_19001,N_14955,N_13505);
xnor U19002 (N_19002,N_14175,N_11816);
nand U19003 (N_19003,N_12158,N_11993);
and U19004 (N_19004,N_11463,N_14016);
nand U19005 (N_19005,N_10777,N_11731);
nor U19006 (N_19006,N_12184,N_11526);
or U19007 (N_19007,N_11549,N_10258);
or U19008 (N_19008,N_12237,N_10763);
xnor U19009 (N_19009,N_13081,N_11335);
nor U19010 (N_19010,N_10251,N_12179);
xor U19011 (N_19011,N_11911,N_13520);
nand U19012 (N_19012,N_11790,N_14567);
or U19013 (N_19013,N_14446,N_13518);
or U19014 (N_19014,N_11105,N_10075);
nand U19015 (N_19015,N_10830,N_14695);
nand U19016 (N_19016,N_11721,N_13260);
nor U19017 (N_19017,N_10914,N_10885);
or U19018 (N_19018,N_11520,N_13582);
xnor U19019 (N_19019,N_14405,N_11342);
or U19020 (N_19020,N_11426,N_11849);
xnor U19021 (N_19021,N_10051,N_12479);
or U19022 (N_19022,N_14884,N_10061);
xnor U19023 (N_19023,N_14156,N_12013);
xor U19024 (N_19024,N_13615,N_13712);
and U19025 (N_19025,N_12794,N_11449);
nor U19026 (N_19026,N_10365,N_11083);
nor U19027 (N_19027,N_14609,N_10784);
xor U19028 (N_19028,N_13626,N_13297);
nor U19029 (N_19029,N_12385,N_11988);
and U19030 (N_19030,N_13062,N_11446);
nand U19031 (N_19031,N_14426,N_13889);
xnor U19032 (N_19032,N_11717,N_11255);
or U19033 (N_19033,N_11260,N_13677);
xor U19034 (N_19034,N_12701,N_13509);
nor U19035 (N_19035,N_10844,N_14812);
and U19036 (N_19036,N_10496,N_12519);
xnor U19037 (N_19037,N_11330,N_10581);
nand U19038 (N_19038,N_13832,N_10463);
and U19039 (N_19039,N_11185,N_12353);
and U19040 (N_19040,N_10092,N_11968);
xnor U19041 (N_19041,N_12635,N_14955);
and U19042 (N_19042,N_14420,N_13376);
or U19043 (N_19043,N_12428,N_11138);
nor U19044 (N_19044,N_10825,N_14559);
or U19045 (N_19045,N_13215,N_13655);
nor U19046 (N_19046,N_13104,N_11591);
nand U19047 (N_19047,N_12803,N_12984);
nor U19048 (N_19048,N_14097,N_11764);
nor U19049 (N_19049,N_14229,N_10413);
nor U19050 (N_19050,N_10097,N_11631);
xor U19051 (N_19051,N_12913,N_12135);
xor U19052 (N_19052,N_11368,N_12474);
and U19053 (N_19053,N_14070,N_11133);
xnor U19054 (N_19054,N_12811,N_11378);
nand U19055 (N_19055,N_10927,N_10697);
nand U19056 (N_19056,N_10951,N_11081);
nand U19057 (N_19057,N_11213,N_10809);
or U19058 (N_19058,N_11028,N_11293);
nand U19059 (N_19059,N_11236,N_14133);
or U19060 (N_19060,N_11387,N_11526);
nand U19061 (N_19061,N_12987,N_10403);
or U19062 (N_19062,N_11653,N_14389);
or U19063 (N_19063,N_10374,N_10969);
nand U19064 (N_19064,N_13327,N_10624);
nand U19065 (N_19065,N_10449,N_11256);
nor U19066 (N_19066,N_13273,N_13601);
or U19067 (N_19067,N_10434,N_10999);
nand U19068 (N_19068,N_11454,N_11175);
or U19069 (N_19069,N_14219,N_13562);
xor U19070 (N_19070,N_12936,N_11987);
nand U19071 (N_19071,N_12871,N_13491);
nand U19072 (N_19072,N_14985,N_12646);
nor U19073 (N_19073,N_13140,N_10657);
xnor U19074 (N_19074,N_13311,N_12318);
nor U19075 (N_19075,N_14379,N_10351);
xnor U19076 (N_19076,N_14459,N_10353);
nand U19077 (N_19077,N_14391,N_13662);
or U19078 (N_19078,N_14838,N_11165);
xnor U19079 (N_19079,N_14715,N_13313);
and U19080 (N_19080,N_13211,N_14919);
nor U19081 (N_19081,N_13095,N_14712);
nor U19082 (N_19082,N_11449,N_10159);
and U19083 (N_19083,N_12419,N_11354);
and U19084 (N_19084,N_12072,N_12540);
nand U19085 (N_19085,N_14885,N_12507);
xor U19086 (N_19086,N_12292,N_14125);
and U19087 (N_19087,N_13306,N_10921);
and U19088 (N_19088,N_11482,N_14446);
xnor U19089 (N_19089,N_14252,N_11468);
or U19090 (N_19090,N_13226,N_13184);
nand U19091 (N_19091,N_12850,N_11382);
or U19092 (N_19092,N_11567,N_10828);
nor U19093 (N_19093,N_11895,N_12864);
or U19094 (N_19094,N_11196,N_12410);
nand U19095 (N_19095,N_11243,N_14605);
nor U19096 (N_19096,N_11657,N_13567);
or U19097 (N_19097,N_10667,N_13904);
or U19098 (N_19098,N_10651,N_10081);
nor U19099 (N_19099,N_14264,N_13831);
or U19100 (N_19100,N_13788,N_10641);
and U19101 (N_19101,N_13424,N_11760);
xor U19102 (N_19102,N_13959,N_13518);
and U19103 (N_19103,N_11705,N_13088);
or U19104 (N_19104,N_11090,N_10916);
nor U19105 (N_19105,N_14526,N_11576);
nor U19106 (N_19106,N_13321,N_14048);
and U19107 (N_19107,N_14123,N_14513);
nor U19108 (N_19108,N_10143,N_13395);
xor U19109 (N_19109,N_14311,N_12477);
and U19110 (N_19110,N_14740,N_14618);
nor U19111 (N_19111,N_11635,N_14545);
and U19112 (N_19112,N_11701,N_14097);
and U19113 (N_19113,N_10198,N_12546);
nand U19114 (N_19114,N_12821,N_12872);
nor U19115 (N_19115,N_14366,N_11137);
and U19116 (N_19116,N_14510,N_11896);
nor U19117 (N_19117,N_13140,N_11035);
and U19118 (N_19118,N_14601,N_11198);
nor U19119 (N_19119,N_13768,N_11482);
nand U19120 (N_19120,N_12389,N_14617);
nor U19121 (N_19121,N_10918,N_10510);
nand U19122 (N_19122,N_14606,N_13404);
nor U19123 (N_19123,N_11124,N_11043);
nor U19124 (N_19124,N_11531,N_11272);
xor U19125 (N_19125,N_13548,N_12468);
nor U19126 (N_19126,N_11801,N_11947);
nor U19127 (N_19127,N_13246,N_10435);
or U19128 (N_19128,N_14518,N_13000);
and U19129 (N_19129,N_11682,N_11347);
xnor U19130 (N_19130,N_10427,N_12765);
nand U19131 (N_19131,N_11099,N_12860);
or U19132 (N_19132,N_11645,N_13469);
or U19133 (N_19133,N_13275,N_13416);
or U19134 (N_19134,N_10790,N_10410);
or U19135 (N_19135,N_10508,N_13344);
or U19136 (N_19136,N_10241,N_11387);
and U19137 (N_19137,N_12060,N_11908);
or U19138 (N_19138,N_14292,N_13724);
or U19139 (N_19139,N_10278,N_10999);
or U19140 (N_19140,N_10339,N_14958);
xnor U19141 (N_19141,N_10322,N_14464);
nand U19142 (N_19142,N_10818,N_13096);
or U19143 (N_19143,N_11449,N_13437);
xnor U19144 (N_19144,N_11740,N_13623);
xnor U19145 (N_19145,N_12387,N_11851);
nor U19146 (N_19146,N_12283,N_12780);
nor U19147 (N_19147,N_11927,N_14038);
xor U19148 (N_19148,N_11118,N_10848);
xnor U19149 (N_19149,N_11233,N_10389);
xnor U19150 (N_19150,N_12311,N_13144);
or U19151 (N_19151,N_12090,N_13397);
and U19152 (N_19152,N_10753,N_12131);
and U19153 (N_19153,N_14153,N_13030);
xnor U19154 (N_19154,N_12156,N_14416);
xor U19155 (N_19155,N_13347,N_14943);
nor U19156 (N_19156,N_13962,N_13954);
or U19157 (N_19157,N_10336,N_14343);
or U19158 (N_19158,N_10025,N_12522);
xnor U19159 (N_19159,N_12718,N_14427);
xnor U19160 (N_19160,N_13864,N_12442);
or U19161 (N_19161,N_11911,N_13371);
and U19162 (N_19162,N_11414,N_10909);
xor U19163 (N_19163,N_14396,N_11086);
nand U19164 (N_19164,N_14307,N_13502);
nand U19165 (N_19165,N_10683,N_10754);
xor U19166 (N_19166,N_10987,N_12369);
and U19167 (N_19167,N_13121,N_12893);
nor U19168 (N_19168,N_11054,N_12083);
xnor U19169 (N_19169,N_12789,N_14207);
xor U19170 (N_19170,N_14488,N_14319);
nand U19171 (N_19171,N_10287,N_14024);
nor U19172 (N_19172,N_10683,N_10499);
xor U19173 (N_19173,N_12240,N_13449);
and U19174 (N_19174,N_10956,N_12914);
or U19175 (N_19175,N_13645,N_13720);
nor U19176 (N_19176,N_13036,N_13467);
xnor U19177 (N_19177,N_13869,N_12913);
nor U19178 (N_19178,N_14018,N_10947);
xnor U19179 (N_19179,N_11645,N_14344);
and U19180 (N_19180,N_14765,N_12627);
and U19181 (N_19181,N_12467,N_10511);
and U19182 (N_19182,N_10274,N_10086);
nor U19183 (N_19183,N_14347,N_12780);
or U19184 (N_19184,N_12816,N_12995);
nand U19185 (N_19185,N_10191,N_11130);
nand U19186 (N_19186,N_11852,N_13602);
nor U19187 (N_19187,N_12439,N_10470);
xnor U19188 (N_19188,N_12807,N_14821);
xnor U19189 (N_19189,N_10183,N_14387);
and U19190 (N_19190,N_10191,N_10432);
nor U19191 (N_19191,N_12605,N_12662);
or U19192 (N_19192,N_10593,N_10109);
and U19193 (N_19193,N_13853,N_14387);
or U19194 (N_19194,N_14602,N_10978);
nor U19195 (N_19195,N_11348,N_12218);
xnor U19196 (N_19196,N_10499,N_14630);
and U19197 (N_19197,N_12233,N_10470);
nor U19198 (N_19198,N_14843,N_12864);
xor U19199 (N_19199,N_13219,N_13000);
or U19200 (N_19200,N_10055,N_13226);
nor U19201 (N_19201,N_11903,N_12353);
or U19202 (N_19202,N_14518,N_14923);
or U19203 (N_19203,N_13408,N_14908);
xnor U19204 (N_19204,N_12564,N_14240);
xor U19205 (N_19205,N_14702,N_12560);
and U19206 (N_19206,N_10810,N_12837);
xor U19207 (N_19207,N_12652,N_12659);
xor U19208 (N_19208,N_14591,N_14636);
nand U19209 (N_19209,N_11568,N_12820);
and U19210 (N_19210,N_14853,N_13530);
or U19211 (N_19211,N_14258,N_10622);
or U19212 (N_19212,N_10687,N_13502);
and U19213 (N_19213,N_11344,N_13920);
nand U19214 (N_19214,N_11844,N_10662);
xnor U19215 (N_19215,N_14070,N_14916);
nand U19216 (N_19216,N_13043,N_11188);
xor U19217 (N_19217,N_14415,N_10854);
and U19218 (N_19218,N_11106,N_12374);
nand U19219 (N_19219,N_14015,N_10667);
or U19220 (N_19220,N_12824,N_13824);
nor U19221 (N_19221,N_12587,N_12483);
and U19222 (N_19222,N_13803,N_12812);
and U19223 (N_19223,N_11379,N_12155);
or U19224 (N_19224,N_13446,N_13088);
xor U19225 (N_19225,N_12803,N_14936);
and U19226 (N_19226,N_11901,N_14953);
or U19227 (N_19227,N_12548,N_11126);
nand U19228 (N_19228,N_14630,N_10032);
nand U19229 (N_19229,N_11543,N_14895);
nor U19230 (N_19230,N_12020,N_10191);
or U19231 (N_19231,N_13239,N_13582);
and U19232 (N_19232,N_13722,N_12086);
nand U19233 (N_19233,N_12023,N_14479);
xnor U19234 (N_19234,N_11932,N_14027);
and U19235 (N_19235,N_10035,N_11929);
xnor U19236 (N_19236,N_12079,N_10380);
xor U19237 (N_19237,N_11139,N_12085);
xor U19238 (N_19238,N_10325,N_14179);
xnor U19239 (N_19239,N_12030,N_13222);
or U19240 (N_19240,N_14649,N_12781);
nor U19241 (N_19241,N_11567,N_10600);
nand U19242 (N_19242,N_10229,N_11203);
xnor U19243 (N_19243,N_14015,N_12101);
nor U19244 (N_19244,N_12214,N_13052);
xor U19245 (N_19245,N_12028,N_10309);
nor U19246 (N_19246,N_12214,N_10678);
and U19247 (N_19247,N_12052,N_11191);
xor U19248 (N_19248,N_10969,N_11199);
nor U19249 (N_19249,N_10827,N_12135);
nand U19250 (N_19250,N_13631,N_10089);
nand U19251 (N_19251,N_13532,N_13097);
nor U19252 (N_19252,N_10272,N_10554);
nand U19253 (N_19253,N_10683,N_10424);
nor U19254 (N_19254,N_13766,N_11915);
nor U19255 (N_19255,N_14954,N_14437);
nand U19256 (N_19256,N_11596,N_12406);
and U19257 (N_19257,N_10775,N_11043);
and U19258 (N_19258,N_13118,N_10163);
xor U19259 (N_19259,N_10398,N_11536);
or U19260 (N_19260,N_14114,N_11738);
xor U19261 (N_19261,N_14522,N_10493);
xor U19262 (N_19262,N_10280,N_10334);
xnor U19263 (N_19263,N_10773,N_11826);
or U19264 (N_19264,N_13443,N_10919);
and U19265 (N_19265,N_14311,N_14820);
or U19266 (N_19266,N_14604,N_13653);
or U19267 (N_19267,N_14028,N_12463);
nor U19268 (N_19268,N_11151,N_10311);
and U19269 (N_19269,N_13837,N_10464);
and U19270 (N_19270,N_12447,N_14085);
xnor U19271 (N_19271,N_14920,N_11466);
nor U19272 (N_19272,N_14901,N_14973);
nand U19273 (N_19273,N_11501,N_12169);
nor U19274 (N_19274,N_12346,N_11348);
and U19275 (N_19275,N_12824,N_13058);
or U19276 (N_19276,N_10475,N_13239);
nand U19277 (N_19277,N_10900,N_13568);
xor U19278 (N_19278,N_13843,N_13695);
and U19279 (N_19279,N_10502,N_12022);
xnor U19280 (N_19280,N_12253,N_14050);
xnor U19281 (N_19281,N_12636,N_14182);
nand U19282 (N_19282,N_12030,N_14511);
and U19283 (N_19283,N_13583,N_13376);
nor U19284 (N_19284,N_12322,N_10415);
and U19285 (N_19285,N_13215,N_10147);
xor U19286 (N_19286,N_12619,N_13468);
nand U19287 (N_19287,N_11113,N_11654);
or U19288 (N_19288,N_10108,N_14561);
and U19289 (N_19289,N_13888,N_13752);
xor U19290 (N_19290,N_14616,N_11330);
nor U19291 (N_19291,N_10583,N_11639);
or U19292 (N_19292,N_11251,N_14147);
or U19293 (N_19293,N_13739,N_11381);
xor U19294 (N_19294,N_14025,N_13180);
nand U19295 (N_19295,N_11346,N_13128);
nor U19296 (N_19296,N_12311,N_11100);
or U19297 (N_19297,N_12684,N_10710);
nand U19298 (N_19298,N_12812,N_10101);
nand U19299 (N_19299,N_13118,N_11244);
nand U19300 (N_19300,N_13016,N_11890);
and U19301 (N_19301,N_12698,N_12956);
xor U19302 (N_19302,N_11588,N_10682);
and U19303 (N_19303,N_11984,N_12870);
nor U19304 (N_19304,N_12887,N_11992);
xnor U19305 (N_19305,N_14531,N_11253);
nor U19306 (N_19306,N_13568,N_11220);
nor U19307 (N_19307,N_10242,N_11353);
xnor U19308 (N_19308,N_12575,N_10069);
nand U19309 (N_19309,N_12001,N_12008);
xor U19310 (N_19310,N_14883,N_13076);
nand U19311 (N_19311,N_13331,N_12399);
or U19312 (N_19312,N_14590,N_11949);
or U19313 (N_19313,N_13091,N_12784);
or U19314 (N_19314,N_14902,N_14861);
xor U19315 (N_19315,N_12458,N_12420);
nand U19316 (N_19316,N_12329,N_14386);
nand U19317 (N_19317,N_11515,N_10990);
and U19318 (N_19318,N_10804,N_14012);
xnor U19319 (N_19319,N_10139,N_11314);
or U19320 (N_19320,N_14286,N_14666);
nand U19321 (N_19321,N_13535,N_14958);
and U19322 (N_19322,N_13414,N_14897);
and U19323 (N_19323,N_13275,N_10217);
nand U19324 (N_19324,N_12864,N_14014);
and U19325 (N_19325,N_11894,N_12837);
nor U19326 (N_19326,N_11016,N_13153);
nand U19327 (N_19327,N_14120,N_14122);
xor U19328 (N_19328,N_10260,N_10717);
nand U19329 (N_19329,N_11480,N_11294);
or U19330 (N_19330,N_10171,N_13027);
nor U19331 (N_19331,N_10116,N_12912);
xnor U19332 (N_19332,N_12782,N_14705);
nand U19333 (N_19333,N_14708,N_11185);
nand U19334 (N_19334,N_12738,N_11977);
xnor U19335 (N_19335,N_10662,N_14876);
nor U19336 (N_19336,N_10896,N_14707);
nor U19337 (N_19337,N_12605,N_12186);
or U19338 (N_19338,N_10211,N_13572);
xnor U19339 (N_19339,N_11031,N_11663);
nand U19340 (N_19340,N_10122,N_11580);
and U19341 (N_19341,N_12080,N_11803);
xnor U19342 (N_19342,N_14417,N_13865);
or U19343 (N_19343,N_10390,N_12553);
and U19344 (N_19344,N_11487,N_13361);
nor U19345 (N_19345,N_13089,N_12489);
and U19346 (N_19346,N_12034,N_14427);
xnor U19347 (N_19347,N_11052,N_11675);
or U19348 (N_19348,N_10929,N_12827);
or U19349 (N_19349,N_12726,N_14412);
nand U19350 (N_19350,N_12184,N_13345);
nor U19351 (N_19351,N_11464,N_10263);
nor U19352 (N_19352,N_12909,N_10414);
nor U19353 (N_19353,N_11747,N_10910);
nor U19354 (N_19354,N_14674,N_12151);
nor U19355 (N_19355,N_13288,N_12108);
xnor U19356 (N_19356,N_14644,N_10831);
and U19357 (N_19357,N_11233,N_11628);
or U19358 (N_19358,N_13503,N_14636);
and U19359 (N_19359,N_10284,N_11620);
nand U19360 (N_19360,N_13410,N_12484);
nand U19361 (N_19361,N_13478,N_14388);
and U19362 (N_19362,N_13093,N_13011);
xnor U19363 (N_19363,N_14111,N_13092);
xor U19364 (N_19364,N_14382,N_11730);
or U19365 (N_19365,N_12124,N_14911);
nor U19366 (N_19366,N_10092,N_12203);
nor U19367 (N_19367,N_10587,N_14397);
nand U19368 (N_19368,N_11122,N_11417);
nor U19369 (N_19369,N_12516,N_11062);
nor U19370 (N_19370,N_11464,N_11746);
xor U19371 (N_19371,N_13279,N_11999);
and U19372 (N_19372,N_14456,N_13915);
nor U19373 (N_19373,N_12166,N_14557);
nand U19374 (N_19374,N_11043,N_14577);
nand U19375 (N_19375,N_12485,N_13386);
nand U19376 (N_19376,N_11746,N_10266);
nor U19377 (N_19377,N_12971,N_13286);
nand U19378 (N_19378,N_14204,N_12152);
nor U19379 (N_19379,N_11774,N_11577);
nand U19380 (N_19380,N_11225,N_12635);
or U19381 (N_19381,N_14872,N_12521);
nor U19382 (N_19382,N_12379,N_12141);
nand U19383 (N_19383,N_13387,N_10951);
nor U19384 (N_19384,N_11384,N_13190);
nor U19385 (N_19385,N_14784,N_14612);
and U19386 (N_19386,N_11776,N_11512);
and U19387 (N_19387,N_13209,N_11489);
nand U19388 (N_19388,N_12758,N_14303);
or U19389 (N_19389,N_11761,N_13079);
and U19390 (N_19390,N_12942,N_10262);
nor U19391 (N_19391,N_12623,N_12271);
nor U19392 (N_19392,N_12115,N_11008);
and U19393 (N_19393,N_13252,N_13722);
and U19394 (N_19394,N_13696,N_10687);
and U19395 (N_19395,N_11597,N_14862);
nor U19396 (N_19396,N_12223,N_11845);
nand U19397 (N_19397,N_13825,N_13420);
or U19398 (N_19398,N_14136,N_12825);
xnor U19399 (N_19399,N_10153,N_13455);
nor U19400 (N_19400,N_11148,N_13241);
nand U19401 (N_19401,N_14923,N_12993);
nor U19402 (N_19402,N_13043,N_12220);
and U19403 (N_19403,N_11978,N_13353);
nor U19404 (N_19404,N_13807,N_14132);
xor U19405 (N_19405,N_10974,N_11720);
nand U19406 (N_19406,N_10258,N_12808);
nand U19407 (N_19407,N_14321,N_10076);
and U19408 (N_19408,N_12573,N_14030);
and U19409 (N_19409,N_14327,N_10292);
and U19410 (N_19410,N_14965,N_11526);
nand U19411 (N_19411,N_12779,N_10195);
and U19412 (N_19412,N_13549,N_13287);
nor U19413 (N_19413,N_11903,N_14690);
or U19414 (N_19414,N_11397,N_10564);
or U19415 (N_19415,N_14418,N_14579);
and U19416 (N_19416,N_11643,N_14077);
and U19417 (N_19417,N_10045,N_13597);
and U19418 (N_19418,N_12692,N_11836);
and U19419 (N_19419,N_10513,N_13725);
xnor U19420 (N_19420,N_11190,N_11782);
and U19421 (N_19421,N_14285,N_11252);
or U19422 (N_19422,N_12656,N_14548);
and U19423 (N_19423,N_11998,N_11293);
xor U19424 (N_19424,N_10324,N_12718);
nand U19425 (N_19425,N_14310,N_14749);
and U19426 (N_19426,N_11164,N_12798);
or U19427 (N_19427,N_11147,N_11781);
or U19428 (N_19428,N_10977,N_11397);
or U19429 (N_19429,N_14405,N_10240);
and U19430 (N_19430,N_10214,N_12014);
and U19431 (N_19431,N_14077,N_14940);
xor U19432 (N_19432,N_14400,N_12031);
nand U19433 (N_19433,N_14463,N_13694);
xnor U19434 (N_19434,N_11956,N_12388);
or U19435 (N_19435,N_10264,N_10880);
or U19436 (N_19436,N_12039,N_14436);
xnor U19437 (N_19437,N_14143,N_13811);
nor U19438 (N_19438,N_14199,N_10798);
xor U19439 (N_19439,N_14303,N_12378);
nand U19440 (N_19440,N_14360,N_10678);
xor U19441 (N_19441,N_13258,N_13718);
xnor U19442 (N_19442,N_13478,N_13698);
xnor U19443 (N_19443,N_10036,N_12619);
nor U19444 (N_19444,N_10228,N_13397);
xor U19445 (N_19445,N_14434,N_12963);
and U19446 (N_19446,N_12772,N_10670);
xnor U19447 (N_19447,N_13339,N_13930);
or U19448 (N_19448,N_13123,N_13824);
and U19449 (N_19449,N_13615,N_14625);
or U19450 (N_19450,N_10084,N_13679);
xor U19451 (N_19451,N_12207,N_10096);
nor U19452 (N_19452,N_11558,N_14769);
xor U19453 (N_19453,N_11727,N_14745);
nand U19454 (N_19454,N_14567,N_11526);
nand U19455 (N_19455,N_13300,N_12118);
nand U19456 (N_19456,N_12189,N_11471);
xor U19457 (N_19457,N_10632,N_11110);
xnor U19458 (N_19458,N_13636,N_11663);
or U19459 (N_19459,N_13554,N_13432);
or U19460 (N_19460,N_12927,N_10782);
or U19461 (N_19461,N_11882,N_12533);
nor U19462 (N_19462,N_10426,N_13088);
nand U19463 (N_19463,N_11211,N_11746);
and U19464 (N_19464,N_12113,N_13201);
and U19465 (N_19465,N_10657,N_11752);
and U19466 (N_19466,N_14766,N_11324);
nand U19467 (N_19467,N_12757,N_13727);
and U19468 (N_19468,N_14324,N_12287);
or U19469 (N_19469,N_14725,N_14748);
xnor U19470 (N_19470,N_10746,N_14607);
and U19471 (N_19471,N_13940,N_14174);
or U19472 (N_19472,N_10489,N_11711);
and U19473 (N_19473,N_11799,N_11563);
nor U19474 (N_19474,N_11359,N_12360);
nand U19475 (N_19475,N_12199,N_14528);
and U19476 (N_19476,N_11650,N_10931);
and U19477 (N_19477,N_14088,N_12936);
or U19478 (N_19478,N_13443,N_10889);
and U19479 (N_19479,N_14928,N_10123);
xor U19480 (N_19480,N_10499,N_12374);
or U19481 (N_19481,N_14731,N_14009);
xor U19482 (N_19482,N_14202,N_13192);
xnor U19483 (N_19483,N_11422,N_11344);
nand U19484 (N_19484,N_10009,N_12042);
nand U19485 (N_19485,N_12561,N_14134);
and U19486 (N_19486,N_12283,N_10678);
or U19487 (N_19487,N_13524,N_11985);
nor U19488 (N_19488,N_13871,N_10865);
nand U19489 (N_19489,N_11690,N_10510);
or U19490 (N_19490,N_12086,N_11111);
and U19491 (N_19491,N_13751,N_14148);
xnor U19492 (N_19492,N_14999,N_12538);
nand U19493 (N_19493,N_11614,N_13713);
and U19494 (N_19494,N_14195,N_13823);
xor U19495 (N_19495,N_11092,N_12972);
and U19496 (N_19496,N_12142,N_10567);
xor U19497 (N_19497,N_14330,N_11953);
xor U19498 (N_19498,N_14734,N_13438);
nor U19499 (N_19499,N_13399,N_12903);
and U19500 (N_19500,N_14974,N_11407);
nand U19501 (N_19501,N_14373,N_14155);
or U19502 (N_19502,N_11050,N_10112);
or U19503 (N_19503,N_13178,N_13703);
and U19504 (N_19504,N_11836,N_10085);
nand U19505 (N_19505,N_11545,N_13130);
nand U19506 (N_19506,N_11285,N_11648);
xor U19507 (N_19507,N_13122,N_10291);
or U19508 (N_19508,N_13206,N_14706);
and U19509 (N_19509,N_12855,N_13963);
nand U19510 (N_19510,N_10135,N_12704);
or U19511 (N_19511,N_14864,N_10020);
and U19512 (N_19512,N_14376,N_11747);
xnor U19513 (N_19513,N_13583,N_12894);
and U19514 (N_19514,N_14947,N_13939);
or U19515 (N_19515,N_12491,N_11151);
and U19516 (N_19516,N_11928,N_13799);
nand U19517 (N_19517,N_10182,N_14280);
and U19518 (N_19518,N_12589,N_12205);
xnor U19519 (N_19519,N_13053,N_12124);
nor U19520 (N_19520,N_14792,N_10957);
xor U19521 (N_19521,N_12044,N_13895);
or U19522 (N_19522,N_13552,N_11096);
nand U19523 (N_19523,N_11641,N_11995);
nand U19524 (N_19524,N_13954,N_11378);
or U19525 (N_19525,N_12406,N_11055);
xor U19526 (N_19526,N_14354,N_13961);
xnor U19527 (N_19527,N_12320,N_14442);
and U19528 (N_19528,N_14524,N_12214);
or U19529 (N_19529,N_11553,N_11977);
and U19530 (N_19530,N_10722,N_12253);
nor U19531 (N_19531,N_14228,N_10982);
or U19532 (N_19532,N_10451,N_10670);
nand U19533 (N_19533,N_14384,N_14885);
nor U19534 (N_19534,N_12413,N_14515);
or U19535 (N_19535,N_10858,N_13309);
nor U19536 (N_19536,N_11545,N_11801);
or U19537 (N_19537,N_13968,N_14660);
nand U19538 (N_19538,N_11795,N_10902);
xor U19539 (N_19539,N_10149,N_13294);
nand U19540 (N_19540,N_13784,N_12867);
xnor U19541 (N_19541,N_14368,N_14060);
or U19542 (N_19542,N_13075,N_14266);
and U19543 (N_19543,N_13162,N_14762);
xor U19544 (N_19544,N_12346,N_10444);
nand U19545 (N_19545,N_12749,N_13559);
nor U19546 (N_19546,N_14791,N_10887);
and U19547 (N_19547,N_10236,N_10048);
nand U19548 (N_19548,N_13275,N_11957);
nor U19549 (N_19549,N_10828,N_11349);
or U19550 (N_19550,N_14584,N_13042);
and U19551 (N_19551,N_12803,N_12337);
or U19552 (N_19552,N_12006,N_13488);
nand U19553 (N_19553,N_11300,N_11642);
nor U19554 (N_19554,N_14257,N_11295);
nor U19555 (N_19555,N_14774,N_10705);
nor U19556 (N_19556,N_10268,N_10281);
xor U19557 (N_19557,N_13748,N_10257);
nand U19558 (N_19558,N_13384,N_11578);
nor U19559 (N_19559,N_13651,N_11923);
and U19560 (N_19560,N_12615,N_10619);
nor U19561 (N_19561,N_11446,N_14550);
xnor U19562 (N_19562,N_12623,N_14112);
nand U19563 (N_19563,N_11448,N_13108);
nand U19564 (N_19564,N_10189,N_12343);
nand U19565 (N_19565,N_10536,N_10202);
and U19566 (N_19566,N_13003,N_12731);
nor U19567 (N_19567,N_13595,N_14235);
xor U19568 (N_19568,N_14572,N_14104);
or U19569 (N_19569,N_13898,N_10343);
and U19570 (N_19570,N_11687,N_13013);
nor U19571 (N_19571,N_13349,N_11796);
nand U19572 (N_19572,N_14679,N_11669);
or U19573 (N_19573,N_11987,N_11775);
and U19574 (N_19574,N_12439,N_12720);
nand U19575 (N_19575,N_11974,N_11318);
and U19576 (N_19576,N_11195,N_10181);
xor U19577 (N_19577,N_14133,N_14442);
xnor U19578 (N_19578,N_13478,N_12815);
nor U19579 (N_19579,N_12641,N_11440);
and U19580 (N_19580,N_12793,N_13043);
xnor U19581 (N_19581,N_12276,N_14881);
or U19582 (N_19582,N_13930,N_14573);
xor U19583 (N_19583,N_11959,N_13078);
and U19584 (N_19584,N_13041,N_12684);
xor U19585 (N_19585,N_11134,N_14701);
xnor U19586 (N_19586,N_13519,N_13019);
and U19587 (N_19587,N_10163,N_10784);
nand U19588 (N_19588,N_14821,N_13826);
xnor U19589 (N_19589,N_10338,N_14423);
nor U19590 (N_19590,N_10845,N_13781);
xnor U19591 (N_19591,N_10839,N_10057);
or U19592 (N_19592,N_13345,N_11046);
or U19593 (N_19593,N_12419,N_13133);
nand U19594 (N_19594,N_13158,N_11284);
or U19595 (N_19595,N_12937,N_13546);
xnor U19596 (N_19596,N_12887,N_11452);
xor U19597 (N_19597,N_11807,N_10479);
nor U19598 (N_19598,N_14318,N_11901);
nand U19599 (N_19599,N_14893,N_10422);
or U19600 (N_19600,N_14531,N_12281);
nor U19601 (N_19601,N_14165,N_13562);
or U19602 (N_19602,N_13788,N_10703);
nor U19603 (N_19603,N_11661,N_14623);
nor U19604 (N_19604,N_14486,N_13055);
nor U19605 (N_19605,N_11141,N_11542);
or U19606 (N_19606,N_12518,N_11275);
or U19607 (N_19607,N_14800,N_12908);
and U19608 (N_19608,N_14730,N_10557);
nand U19609 (N_19609,N_14722,N_11330);
xnor U19610 (N_19610,N_12848,N_12374);
nand U19611 (N_19611,N_10102,N_12219);
nor U19612 (N_19612,N_12921,N_10699);
and U19613 (N_19613,N_12305,N_10310);
nand U19614 (N_19614,N_10260,N_12739);
nand U19615 (N_19615,N_14217,N_14857);
nand U19616 (N_19616,N_11928,N_11589);
nand U19617 (N_19617,N_10664,N_10340);
or U19618 (N_19618,N_14223,N_11554);
or U19619 (N_19619,N_13653,N_12988);
nor U19620 (N_19620,N_10379,N_12885);
xor U19621 (N_19621,N_12153,N_14247);
nor U19622 (N_19622,N_13663,N_12461);
nor U19623 (N_19623,N_10358,N_14597);
or U19624 (N_19624,N_14401,N_12134);
nor U19625 (N_19625,N_12256,N_13132);
nor U19626 (N_19626,N_11390,N_12624);
and U19627 (N_19627,N_11068,N_12309);
and U19628 (N_19628,N_13526,N_12895);
and U19629 (N_19629,N_11703,N_10645);
nand U19630 (N_19630,N_13954,N_13777);
nor U19631 (N_19631,N_14823,N_14740);
and U19632 (N_19632,N_11303,N_13919);
xnor U19633 (N_19633,N_12448,N_10884);
nand U19634 (N_19634,N_14658,N_11359);
or U19635 (N_19635,N_11435,N_13196);
nand U19636 (N_19636,N_10690,N_11543);
nor U19637 (N_19637,N_13999,N_12696);
nand U19638 (N_19638,N_13548,N_10805);
nor U19639 (N_19639,N_10693,N_10465);
nor U19640 (N_19640,N_13933,N_11071);
and U19641 (N_19641,N_13493,N_10454);
xor U19642 (N_19642,N_11074,N_14486);
and U19643 (N_19643,N_12277,N_11891);
nor U19644 (N_19644,N_11910,N_14153);
or U19645 (N_19645,N_11751,N_14302);
nor U19646 (N_19646,N_14960,N_12824);
and U19647 (N_19647,N_11152,N_12330);
nand U19648 (N_19648,N_10759,N_12983);
or U19649 (N_19649,N_14686,N_13176);
or U19650 (N_19650,N_10472,N_11231);
or U19651 (N_19651,N_13550,N_10954);
nor U19652 (N_19652,N_12888,N_10048);
or U19653 (N_19653,N_12862,N_12726);
or U19654 (N_19654,N_10678,N_10683);
or U19655 (N_19655,N_14629,N_10701);
nand U19656 (N_19656,N_14682,N_11329);
xnor U19657 (N_19657,N_12315,N_11231);
nor U19658 (N_19658,N_14954,N_11520);
xor U19659 (N_19659,N_11774,N_12089);
nand U19660 (N_19660,N_14855,N_12115);
xor U19661 (N_19661,N_13139,N_12500);
xnor U19662 (N_19662,N_14649,N_14166);
nand U19663 (N_19663,N_12843,N_12480);
nand U19664 (N_19664,N_13665,N_11571);
xnor U19665 (N_19665,N_13025,N_13501);
xor U19666 (N_19666,N_14881,N_14030);
and U19667 (N_19667,N_14805,N_14561);
or U19668 (N_19668,N_13094,N_13514);
nor U19669 (N_19669,N_12113,N_13096);
and U19670 (N_19670,N_12069,N_10700);
nand U19671 (N_19671,N_10060,N_14126);
and U19672 (N_19672,N_10154,N_11553);
or U19673 (N_19673,N_10180,N_13274);
nor U19674 (N_19674,N_13838,N_14091);
nand U19675 (N_19675,N_11572,N_11779);
nand U19676 (N_19676,N_11470,N_14359);
or U19677 (N_19677,N_10269,N_10264);
and U19678 (N_19678,N_13279,N_11798);
xnor U19679 (N_19679,N_12630,N_14092);
and U19680 (N_19680,N_13376,N_14061);
nand U19681 (N_19681,N_14925,N_13753);
xnor U19682 (N_19682,N_10423,N_11420);
xor U19683 (N_19683,N_12514,N_11325);
nand U19684 (N_19684,N_11063,N_10200);
and U19685 (N_19685,N_12590,N_10407);
nand U19686 (N_19686,N_14625,N_12480);
xnor U19687 (N_19687,N_13210,N_11061);
nand U19688 (N_19688,N_14306,N_13866);
xnor U19689 (N_19689,N_14742,N_14751);
nand U19690 (N_19690,N_11212,N_11250);
xnor U19691 (N_19691,N_10773,N_14509);
or U19692 (N_19692,N_12464,N_10084);
xnor U19693 (N_19693,N_10951,N_10081);
nor U19694 (N_19694,N_13764,N_11021);
nor U19695 (N_19695,N_11136,N_12747);
or U19696 (N_19696,N_13762,N_12264);
nor U19697 (N_19697,N_12340,N_12210);
nor U19698 (N_19698,N_10178,N_12114);
nand U19699 (N_19699,N_13486,N_14413);
nand U19700 (N_19700,N_12517,N_14492);
and U19701 (N_19701,N_13962,N_10741);
nor U19702 (N_19702,N_10206,N_11626);
and U19703 (N_19703,N_14096,N_14674);
nor U19704 (N_19704,N_14052,N_12847);
or U19705 (N_19705,N_10257,N_14852);
nand U19706 (N_19706,N_13478,N_13919);
nand U19707 (N_19707,N_14732,N_13125);
or U19708 (N_19708,N_10886,N_12265);
or U19709 (N_19709,N_10127,N_11822);
and U19710 (N_19710,N_13631,N_11628);
and U19711 (N_19711,N_13525,N_14750);
and U19712 (N_19712,N_14044,N_12880);
xor U19713 (N_19713,N_11333,N_10603);
nand U19714 (N_19714,N_13264,N_12484);
nand U19715 (N_19715,N_11337,N_14471);
or U19716 (N_19716,N_14552,N_12105);
or U19717 (N_19717,N_12525,N_14503);
xnor U19718 (N_19718,N_14077,N_14788);
and U19719 (N_19719,N_10587,N_13631);
or U19720 (N_19720,N_10553,N_13399);
nand U19721 (N_19721,N_14070,N_10197);
or U19722 (N_19722,N_14575,N_12236);
nand U19723 (N_19723,N_12424,N_11557);
or U19724 (N_19724,N_10756,N_12520);
nand U19725 (N_19725,N_10525,N_13645);
nand U19726 (N_19726,N_13441,N_11518);
nor U19727 (N_19727,N_12842,N_14650);
xor U19728 (N_19728,N_12113,N_12530);
xnor U19729 (N_19729,N_13997,N_13996);
xnor U19730 (N_19730,N_13341,N_11247);
and U19731 (N_19731,N_13137,N_12172);
and U19732 (N_19732,N_10821,N_11370);
or U19733 (N_19733,N_13788,N_11583);
and U19734 (N_19734,N_10741,N_14617);
or U19735 (N_19735,N_14870,N_13941);
nor U19736 (N_19736,N_14801,N_10840);
and U19737 (N_19737,N_12517,N_13755);
xor U19738 (N_19738,N_11696,N_13921);
and U19739 (N_19739,N_11026,N_13637);
xnor U19740 (N_19740,N_12566,N_12742);
nor U19741 (N_19741,N_13798,N_10237);
nor U19742 (N_19742,N_14418,N_14090);
xor U19743 (N_19743,N_14491,N_11035);
xor U19744 (N_19744,N_12305,N_14410);
xnor U19745 (N_19745,N_10317,N_12402);
xor U19746 (N_19746,N_12790,N_13237);
nor U19747 (N_19747,N_14640,N_10475);
and U19748 (N_19748,N_12632,N_12058);
and U19749 (N_19749,N_13858,N_12316);
and U19750 (N_19750,N_11622,N_10328);
or U19751 (N_19751,N_14411,N_14833);
nand U19752 (N_19752,N_13473,N_13665);
nor U19753 (N_19753,N_12464,N_13235);
xor U19754 (N_19754,N_13852,N_13813);
and U19755 (N_19755,N_11909,N_12479);
xor U19756 (N_19756,N_11202,N_13087);
or U19757 (N_19757,N_11096,N_14230);
and U19758 (N_19758,N_11538,N_10587);
or U19759 (N_19759,N_11416,N_14834);
xnor U19760 (N_19760,N_11773,N_12205);
nor U19761 (N_19761,N_12313,N_14569);
nor U19762 (N_19762,N_12845,N_13644);
and U19763 (N_19763,N_14764,N_10966);
nor U19764 (N_19764,N_12752,N_14000);
xor U19765 (N_19765,N_10920,N_13221);
nand U19766 (N_19766,N_14691,N_13233);
nand U19767 (N_19767,N_10444,N_13612);
xor U19768 (N_19768,N_14599,N_13371);
xnor U19769 (N_19769,N_14179,N_13831);
xnor U19770 (N_19770,N_11449,N_10156);
xnor U19771 (N_19771,N_14339,N_13282);
and U19772 (N_19772,N_14670,N_12569);
and U19773 (N_19773,N_10396,N_14967);
or U19774 (N_19774,N_13603,N_12395);
nor U19775 (N_19775,N_14739,N_12018);
nor U19776 (N_19776,N_14097,N_12615);
nor U19777 (N_19777,N_12273,N_12600);
nand U19778 (N_19778,N_11713,N_10897);
nand U19779 (N_19779,N_14245,N_10139);
xnor U19780 (N_19780,N_13388,N_14161);
and U19781 (N_19781,N_11015,N_13270);
nand U19782 (N_19782,N_12425,N_11788);
nor U19783 (N_19783,N_14629,N_14225);
nand U19784 (N_19784,N_12097,N_13566);
nand U19785 (N_19785,N_10805,N_10640);
nand U19786 (N_19786,N_11404,N_11819);
or U19787 (N_19787,N_10786,N_12647);
or U19788 (N_19788,N_13533,N_11549);
nand U19789 (N_19789,N_12571,N_11574);
xnor U19790 (N_19790,N_12304,N_13265);
or U19791 (N_19791,N_13959,N_11641);
nand U19792 (N_19792,N_10329,N_14843);
nand U19793 (N_19793,N_12689,N_14268);
nor U19794 (N_19794,N_13220,N_13846);
xnor U19795 (N_19795,N_10534,N_11662);
or U19796 (N_19796,N_11046,N_11415);
and U19797 (N_19797,N_14718,N_14948);
xor U19798 (N_19798,N_11551,N_14404);
nor U19799 (N_19799,N_11341,N_14397);
xnor U19800 (N_19800,N_14540,N_10902);
nor U19801 (N_19801,N_14060,N_11751);
or U19802 (N_19802,N_11790,N_10148);
nand U19803 (N_19803,N_13939,N_12751);
xnor U19804 (N_19804,N_14237,N_12475);
and U19805 (N_19805,N_13263,N_10815);
and U19806 (N_19806,N_12012,N_13334);
or U19807 (N_19807,N_10553,N_14250);
and U19808 (N_19808,N_14120,N_14327);
nor U19809 (N_19809,N_14444,N_10596);
nor U19810 (N_19810,N_12414,N_10167);
and U19811 (N_19811,N_14251,N_13307);
xor U19812 (N_19812,N_14649,N_12498);
and U19813 (N_19813,N_10331,N_13089);
nand U19814 (N_19814,N_12645,N_12445);
xor U19815 (N_19815,N_14398,N_13717);
xnor U19816 (N_19816,N_12977,N_14783);
xor U19817 (N_19817,N_13267,N_11158);
or U19818 (N_19818,N_14590,N_12698);
nand U19819 (N_19819,N_10678,N_10578);
or U19820 (N_19820,N_10028,N_10455);
and U19821 (N_19821,N_12086,N_10029);
xor U19822 (N_19822,N_11705,N_14844);
nor U19823 (N_19823,N_13254,N_12164);
or U19824 (N_19824,N_10264,N_14133);
nor U19825 (N_19825,N_14396,N_12764);
and U19826 (N_19826,N_11137,N_13606);
nor U19827 (N_19827,N_14399,N_12846);
xor U19828 (N_19828,N_13386,N_13110);
and U19829 (N_19829,N_10864,N_11666);
nand U19830 (N_19830,N_11400,N_10804);
nand U19831 (N_19831,N_10279,N_10207);
xor U19832 (N_19832,N_13406,N_14315);
xor U19833 (N_19833,N_10551,N_11560);
nand U19834 (N_19834,N_14026,N_12048);
or U19835 (N_19835,N_12281,N_10028);
xor U19836 (N_19836,N_14446,N_10774);
and U19837 (N_19837,N_13726,N_13888);
nand U19838 (N_19838,N_10829,N_14138);
and U19839 (N_19839,N_13750,N_11351);
and U19840 (N_19840,N_14812,N_13875);
and U19841 (N_19841,N_10121,N_11782);
nor U19842 (N_19842,N_13698,N_11806);
nor U19843 (N_19843,N_14973,N_12404);
nand U19844 (N_19844,N_10003,N_14581);
and U19845 (N_19845,N_14295,N_14937);
and U19846 (N_19846,N_13652,N_13338);
nand U19847 (N_19847,N_10596,N_13829);
nor U19848 (N_19848,N_12715,N_14967);
nor U19849 (N_19849,N_12585,N_12231);
or U19850 (N_19850,N_11727,N_13668);
xnor U19851 (N_19851,N_14449,N_12889);
nand U19852 (N_19852,N_12914,N_11338);
nand U19853 (N_19853,N_10091,N_14717);
nor U19854 (N_19854,N_14550,N_13518);
nand U19855 (N_19855,N_14650,N_13789);
nand U19856 (N_19856,N_10748,N_13757);
or U19857 (N_19857,N_11077,N_12925);
nor U19858 (N_19858,N_13776,N_11680);
xor U19859 (N_19859,N_11645,N_13795);
nor U19860 (N_19860,N_11155,N_13184);
and U19861 (N_19861,N_10523,N_12471);
nor U19862 (N_19862,N_11059,N_13041);
and U19863 (N_19863,N_10573,N_13875);
and U19864 (N_19864,N_11687,N_12219);
nor U19865 (N_19865,N_13573,N_11741);
nor U19866 (N_19866,N_13167,N_12610);
nor U19867 (N_19867,N_12948,N_13773);
nand U19868 (N_19868,N_10161,N_10786);
nor U19869 (N_19869,N_13022,N_10982);
nand U19870 (N_19870,N_13882,N_11481);
nand U19871 (N_19871,N_11651,N_13888);
nand U19872 (N_19872,N_14906,N_13377);
nor U19873 (N_19873,N_11027,N_10116);
and U19874 (N_19874,N_14547,N_13156);
nand U19875 (N_19875,N_14475,N_12955);
and U19876 (N_19876,N_11276,N_10629);
xor U19877 (N_19877,N_14234,N_10553);
nor U19878 (N_19878,N_12844,N_12778);
nand U19879 (N_19879,N_13111,N_10175);
or U19880 (N_19880,N_13282,N_11235);
or U19881 (N_19881,N_10667,N_12049);
xnor U19882 (N_19882,N_13744,N_14562);
nor U19883 (N_19883,N_11796,N_10928);
and U19884 (N_19884,N_13236,N_11793);
nor U19885 (N_19885,N_12852,N_11171);
or U19886 (N_19886,N_13133,N_12303);
nand U19887 (N_19887,N_11682,N_14944);
nand U19888 (N_19888,N_13148,N_12724);
or U19889 (N_19889,N_14946,N_13209);
xnor U19890 (N_19890,N_12086,N_13545);
xnor U19891 (N_19891,N_14699,N_10675);
or U19892 (N_19892,N_11753,N_11446);
or U19893 (N_19893,N_10640,N_10511);
nor U19894 (N_19894,N_14293,N_11715);
nand U19895 (N_19895,N_11598,N_10960);
nor U19896 (N_19896,N_12241,N_10743);
or U19897 (N_19897,N_11960,N_12871);
xnor U19898 (N_19898,N_14299,N_13482);
nand U19899 (N_19899,N_12941,N_14595);
or U19900 (N_19900,N_14321,N_14130);
xnor U19901 (N_19901,N_13300,N_13916);
and U19902 (N_19902,N_14847,N_12083);
nor U19903 (N_19903,N_13361,N_10807);
xor U19904 (N_19904,N_14994,N_11756);
or U19905 (N_19905,N_11155,N_12050);
and U19906 (N_19906,N_10649,N_14540);
and U19907 (N_19907,N_14361,N_14455);
xor U19908 (N_19908,N_11378,N_13557);
xnor U19909 (N_19909,N_14555,N_13354);
or U19910 (N_19910,N_13222,N_12667);
and U19911 (N_19911,N_14121,N_13473);
and U19912 (N_19912,N_13478,N_12635);
nand U19913 (N_19913,N_14656,N_10167);
nand U19914 (N_19914,N_11053,N_10484);
or U19915 (N_19915,N_11445,N_11438);
or U19916 (N_19916,N_14506,N_11836);
nor U19917 (N_19917,N_13281,N_14092);
and U19918 (N_19918,N_10266,N_14362);
and U19919 (N_19919,N_10842,N_14012);
nand U19920 (N_19920,N_10514,N_12880);
nor U19921 (N_19921,N_12841,N_12800);
xnor U19922 (N_19922,N_13690,N_10213);
and U19923 (N_19923,N_12593,N_13462);
and U19924 (N_19924,N_13766,N_10404);
and U19925 (N_19925,N_13540,N_10854);
nor U19926 (N_19926,N_11029,N_13621);
xor U19927 (N_19927,N_14940,N_13733);
nor U19928 (N_19928,N_14841,N_11802);
or U19929 (N_19929,N_10425,N_13314);
xor U19930 (N_19930,N_10628,N_14601);
xnor U19931 (N_19931,N_12900,N_14523);
nor U19932 (N_19932,N_11148,N_12993);
and U19933 (N_19933,N_13712,N_10420);
and U19934 (N_19934,N_12746,N_14380);
nand U19935 (N_19935,N_14945,N_11396);
nor U19936 (N_19936,N_12216,N_11476);
xor U19937 (N_19937,N_14675,N_10527);
and U19938 (N_19938,N_14078,N_11250);
nand U19939 (N_19939,N_14653,N_14983);
nor U19940 (N_19940,N_12717,N_13976);
or U19941 (N_19941,N_10229,N_11463);
xnor U19942 (N_19942,N_12185,N_12312);
nand U19943 (N_19943,N_13847,N_13219);
or U19944 (N_19944,N_10285,N_12929);
xor U19945 (N_19945,N_13237,N_13896);
nor U19946 (N_19946,N_12801,N_12622);
and U19947 (N_19947,N_14404,N_14680);
xnor U19948 (N_19948,N_11244,N_14457);
xor U19949 (N_19949,N_10491,N_11928);
and U19950 (N_19950,N_10050,N_10652);
or U19951 (N_19951,N_11780,N_14223);
and U19952 (N_19952,N_12139,N_14863);
nor U19953 (N_19953,N_10160,N_14316);
xor U19954 (N_19954,N_13029,N_10494);
nor U19955 (N_19955,N_10097,N_12430);
nor U19956 (N_19956,N_10288,N_12437);
or U19957 (N_19957,N_11091,N_12096);
nand U19958 (N_19958,N_11144,N_12133);
and U19959 (N_19959,N_12472,N_14063);
and U19960 (N_19960,N_11696,N_12101);
nor U19961 (N_19961,N_13342,N_11752);
and U19962 (N_19962,N_11681,N_11409);
xor U19963 (N_19963,N_13144,N_12680);
nor U19964 (N_19964,N_13927,N_12506);
or U19965 (N_19965,N_10971,N_12783);
nand U19966 (N_19966,N_10923,N_14856);
and U19967 (N_19967,N_14103,N_10817);
and U19968 (N_19968,N_10320,N_12497);
nor U19969 (N_19969,N_14029,N_12182);
and U19970 (N_19970,N_13246,N_13388);
nand U19971 (N_19971,N_13016,N_11634);
xnor U19972 (N_19972,N_11528,N_11218);
and U19973 (N_19973,N_10411,N_11464);
nand U19974 (N_19974,N_13547,N_12096);
or U19975 (N_19975,N_12670,N_13564);
xnor U19976 (N_19976,N_10607,N_11818);
nand U19977 (N_19977,N_11499,N_13921);
and U19978 (N_19978,N_14455,N_13963);
xnor U19979 (N_19979,N_13683,N_14891);
nor U19980 (N_19980,N_13120,N_11722);
and U19981 (N_19981,N_11801,N_14787);
nor U19982 (N_19982,N_14151,N_11464);
or U19983 (N_19983,N_10198,N_10611);
and U19984 (N_19984,N_10504,N_12361);
nand U19985 (N_19985,N_10499,N_11164);
or U19986 (N_19986,N_12366,N_12771);
xor U19987 (N_19987,N_11502,N_12415);
and U19988 (N_19988,N_10631,N_10779);
or U19989 (N_19989,N_13437,N_12049);
or U19990 (N_19990,N_11566,N_14660);
nand U19991 (N_19991,N_13537,N_14605);
nand U19992 (N_19992,N_14283,N_13792);
nand U19993 (N_19993,N_11575,N_14123);
nand U19994 (N_19994,N_12861,N_14632);
xnor U19995 (N_19995,N_10916,N_10111);
or U19996 (N_19996,N_11168,N_11735);
xor U19997 (N_19997,N_11332,N_14587);
nand U19998 (N_19998,N_11533,N_14464);
and U19999 (N_19999,N_10328,N_12973);
and U20000 (N_20000,N_17527,N_19116);
nand U20001 (N_20001,N_17936,N_19058);
xnor U20002 (N_20002,N_19624,N_18898);
and U20003 (N_20003,N_16437,N_16869);
nor U20004 (N_20004,N_16423,N_18506);
or U20005 (N_20005,N_17723,N_19250);
nand U20006 (N_20006,N_15349,N_17658);
nand U20007 (N_20007,N_15407,N_15688);
or U20008 (N_20008,N_19488,N_15524);
xnor U20009 (N_20009,N_19996,N_19105);
or U20010 (N_20010,N_19211,N_16905);
and U20011 (N_20011,N_19885,N_16600);
and U20012 (N_20012,N_19103,N_19434);
nor U20013 (N_20013,N_19241,N_19337);
xnor U20014 (N_20014,N_16676,N_16695);
nor U20015 (N_20015,N_16808,N_19468);
or U20016 (N_20016,N_15387,N_15815);
nand U20017 (N_20017,N_18183,N_16907);
and U20018 (N_20018,N_16780,N_15911);
and U20019 (N_20019,N_16567,N_19338);
and U20020 (N_20020,N_17055,N_17119);
or U20021 (N_20021,N_19324,N_16860);
nor U20022 (N_20022,N_18235,N_18493);
and U20023 (N_20023,N_18788,N_17095);
or U20024 (N_20024,N_16652,N_17947);
or U20025 (N_20025,N_17970,N_19345);
or U20026 (N_20026,N_18239,N_18150);
xor U20027 (N_20027,N_17001,N_16852);
or U20028 (N_20028,N_18087,N_15164);
nor U20029 (N_20029,N_15880,N_16528);
xor U20030 (N_20030,N_17544,N_16443);
and U20031 (N_20031,N_15161,N_19965);
and U20032 (N_20032,N_16635,N_18306);
nor U20033 (N_20033,N_15490,N_18403);
or U20034 (N_20034,N_15998,N_18562);
nor U20035 (N_20035,N_15381,N_19010);
or U20036 (N_20036,N_18102,N_17386);
nor U20037 (N_20037,N_19493,N_16422);
nor U20038 (N_20038,N_19588,N_18495);
and U20039 (N_20039,N_17397,N_19879);
and U20040 (N_20040,N_19375,N_19939);
nor U20041 (N_20041,N_19296,N_16186);
and U20042 (N_20042,N_15293,N_19957);
nand U20043 (N_20043,N_17331,N_16468);
and U20044 (N_20044,N_17898,N_17135);
nand U20045 (N_20045,N_16448,N_16083);
or U20046 (N_20046,N_15104,N_15797);
or U20047 (N_20047,N_18074,N_16818);
and U20048 (N_20048,N_18244,N_16418);
xnor U20049 (N_20049,N_18508,N_16856);
and U20050 (N_20050,N_17372,N_18517);
and U20051 (N_20051,N_16775,N_15568);
or U20052 (N_20052,N_18600,N_18216);
nor U20053 (N_20053,N_17218,N_18546);
nor U20054 (N_20054,N_17539,N_19906);
xor U20055 (N_20055,N_18781,N_16883);
xor U20056 (N_20056,N_17863,N_17026);
or U20057 (N_20057,N_19796,N_17499);
nand U20058 (N_20058,N_19976,N_18370);
nand U20059 (N_20059,N_18939,N_18072);
or U20060 (N_20060,N_15320,N_15029);
nor U20061 (N_20061,N_16301,N_17392);
or U20062 (N_20062,N_18471,N_17146);
nand U20063 (N_20063,N_16628,N_19289);
and U20064 (N_20064,N_17513,N_19979);
and U20065 (N_20065,N_18443,N_19057);
nor U20066 (N_20066,N_18022,N_16704);
and U20067 (N_20067,N_18743,N_16784);
xnor U20068 (N_20068,N_15448,N_18585);
xor U20069 (N_20069,N_19706,N_15088);
nand U20070 (N_20070,N_19048,N_18573);
or U20071 (N_20071,N_19578,N_18490);
or U20072 (N_20072,N_16762,N_15890);
or U20073 (N_20073,N_16482,N_17102);
nor U20074 (N_20074,N_17620,N_16058);
nor U20075 (N_20075,N_16759,N_19328);
xnor U20076 (N_20076,N_18994,N_16892);
xor U20077 (N_20077,N_19964,N_18653);
nand U20078 (N_20078,N_16665,N_18956);
xnor U20079 (N_20079,N_17866,N_17576);
nor U20080 (N_20080,N_19688,N_15547);
nor U20081 (N_20081,N_15675,N_18934);
xor U20082 (N_20082,N_16006,N_16229);
xnor U20083 (N_20083,N_18854,N_17877);
xnor U20084 (N_20084,N_17188,N_17647);
and U20085 (N_20085,N_16539,N_19480);
nand U20086 (N_20086,N_18470,N_19650);
and U20087 (N_20087,N_16952,N_19862);
nor U20088 (N_20088,N_18207,N_16156);
nand U20089 (N_20089,N_18613,N_18619);
and U20090 (N_20090,N_17211,N_17213);
nor U20091 (N_20091,N_19034,N_18406);
or U20092 (N_20092,N_19625,N_15945);
nor U20093 (N_20093,N_17017,N_19658);
xor U20094 (N_20094,N_17548,N_18321);
nand U20095 (N_20095,N_17038,N_17064);
nor U20096 (N_20096,N_19270,N_17428);
nor U20097 (N_20097,N_15533,N_15232);
xor U20098 (N_20098,N_17651,N_16703);
or U20099 (N_20099,N_16134,N_17035);
nand U20100 (N_20100,N_19795,N_15722);
and U20101 (N_20101,N_16220,N_15868);
nor U20102 (N_20102,N_16497,N_16070);
xnor U20103 (N_20103,N_17821,N_15796);
and U20104 (N_20104,N_15076,N_16255);
nor U20105 (N_20105,N_15737,N_17785);
xor U20106 (N_20106,N_16767,N_16882);
and U20107 (N_20107,N_16458,N_17185);
or U20108 (N_20108,N_16021,N_17926);
or U20109 (N_20109,N_16467,N_16064);
nand U20110 (N_20110,N_18648,N_16178);
or U20111 (N_20111,N_18711,N_15431);
and U20112 (N_20112,N_18991,N_18430);
nand U20113 (N_20113,N_17087,N_19914);
or U20114 (N_20114,N_15379,N_15556);
nand U20115 (N_20115,N_15734,N_19497);
and U20116 (N_20116,N_18059,N_16701);
or U20117 (N_20117,N_17859,N_17644);
and U20118 (N_20118,N_18533,N_19644);
or U20119 (N_20119,N_17903,N_18132);
nor U20120 (N_20120,N_15565,N_19076);
xor U20121 (N_20121,N_15002,N_19776);
nor U20122 (N_20122,N_17393,N_17956);
or U20123 (N_20123,N_16316,N_18242);
and U20124 (N_20124,N_16823,N_19111);
nor U20125 (N_20125,N_17541,N_17429);
and U20126 (N_20126,N_17674,N_16077);
nand U20127 (N_20127,N_16126,N_15935);
or U20128 (N_20128,N_15714,N_16172);
nand U20129 (N_20129,N_16776,N_19504);
and U20130 (N_20130,N_15402,N_17816);
or U20131 (N_20131,N_15923,N_17965);
or U20132 (N_20132,N_15784,N_15738);
nand U20133 (N_20133,N_17130,N_18908);
nand U20134 (N_20134,N_19411,N_18067);
and U20135 (N_20135,N_18731,N_19100);
nor U20136 (N_20136,N_19155,N_17600);
nor U20137 (N_20137,N_19043,N_15500);
nand U20138 (N_20138,N_17118,N_15828);
or U20139 (N_20139,N_15649,N_18094);
nand U20140 (N_20140,N_16522,N_15783);
xor U20141 (N_20141,N_15212,N_17348);
xnor U20142 (N_20142,N_18276,N_16924);
and U20143 (N_20143,N_18825,N_16505);
xnor U20144 (N_20144,N_19843,N_19937);
and U20145 (N_20145,N_17356,N_16486);
nand U20146 (N_20146,N_17453,N_19192);
nor U20147 (N_20147,N_16867,N_17934);
nand U20148 (N_20148,N_15005,N_18549);
and U20149 (N_20149,N_18532,N_19593);
xor U20150 (N_20150,N_18817,N_18831);
and U20151 (N_20151,N_16460,N_18349);
xnor U20152 (N_20152,N_16000,N_18682);
nor U20153 (N_20153,N_19460,N_19581);
or U20154 (N_20154,N_18120,N_16597);
or U20155 (N_20155,N_17033,N_15944);
nor U20156 (N_20156,N_15888,N_19822);
nor U20157 (N_20157,N_17267,N_17341);
xor U20158 (N_20158,N_18886,N_19317);
or U20159 (N_20159,N_18620,N_16026);
or U20160 (N_20160,N_16292,N_18182);
nor U20161 (N_20161,N_15457,N_15021);
nor U20162 (N_20162,N_18123,N_19729);
nand U20163 (N_20163,N_15264,N_19037);
nor U20164 (N_20164,N_18221,N_17594);
xnor U20165 (N_20165,N_18547,N_16897);
nand U20166 (N_20166,N_16169,N_16039);
xor U20167 (N_20167,N_18425,N_18913);
or U20168 (N_20168,N_19871,N_15288);
nand U20169 (N_20169,N_16516,N_17925);
and U20170 (N_20170,N_16125,N_17769);
xnor U20171 (N_20171,N_17320,N_15598);
nand U20172 (N_20172,N_15985,N_15748);
or U20173 (N_20173,N_16215,N_19917);
or U20174 (N_20174,N_19304,N_18264);
nand U20175 (N_20175,N_19318,N_15501);
and U20176 (N_20176,N_19266,N_18372);
nor U20177 (N_20177,N_18286,N_15303);
and U20178 (N_20178,N_16661,N_16554);
or U20179 (N_20179,N_19558,N_17802);
nand U20180 (N_20180,N_19465,N_18259);
nand U20181 (N_20181,N_17333,N_17014);
nand U20182 (N_20182,N_17760,N_15643);
and U20183 (N_20183,N_18808,N_18971);
xnor U20184 (N_20184,N_15975,N_15658);
xor U20185 (N_20185,N_18899,N_17227);
xor U20186 (N_20186,N_15147,N_16806);
nand U20187 (N_20187,N_17291,N_19456);
or U20188 (N_20188,N_15419,N_15384);
nor U20189 (N_20189,N_18294,N_19055);
nand U20190 (N_20190,N_18659,N_16731);
xor U20191 (N_20191,N_15386,N_17044);
or U20192 (N_20192,N_17198,N_17707);
xnor U20193 (N_20193,N_15131,N_17791);
and U20194 (N_20194,N_18807,N_15909);
and U20195 (N_20195,N_16463,N_17959);
nand U20196 (N_20196,N_18924,N_18667);
and U20197 (N_20197,N_16471,N_16396);
or U20198 (N_20198,N_15703,N_18706);
xor U20199 (N_20199,N_17137,N_15258);
xor U20200 (N_20200,N_15889,N_15120);
or U20201 (N_20201,N_16283,N_16158);
xnor U20202 (N_20202,N_19606,N_15255);
and U20203 (N_20203,N_19394,N_16995);
or U20204 (N_20204,N_15862,N_19412);
and U20205 (N_20205,N_15018,N_15538);
and U20206 (N_20206,N_15509,N_19232);
xnor U20207 (N_20207,N_17706,N_19629);
or U20208 (N_20208,N_18401,N_16394);
or U20209 (N_20209,N_19319,N_16981);
nand U20210 (N_20210,N_18367,N_16304);
nand U20211 (N_20211,N_17603,N_19421);
xnor U20212 (N_20212,N_18487,N_15534);
and U20213 (N_20213,N_16576,N_15835);
xor U20214 (N_20214,N_19183,N_18023);
nor U20215 (N_20215,N_18029,N_16985);
and U20216 (N_20216,N_16097,N_16251);
xnor U20217 (N_20217,N_17986,N_16564);
or U20218 (N_20218,N_17729,N_18478);
and U20219 (N_20219,N_16433,N_19259);
nand U20220 (N_20220,N_15593,N_17011);
nor U20221 (N_20221,N_16876,N_16593);
xnor U20222 (N_20222,N_18290,N_19423);
xnor U20223 (N_20223,N_15199,N_15884);
and U20224 (N_20224,N_15251,N_15809);
and U20225 (N_20225,N_16138,N_16076);
and U20226 (N_20226,N_15248,N_19240);
xnor U20227 (N_20227,N_16520,N_15110);
nand U20228 (N_20228,N_17025,N_19522);
xnor U20229 (N_20229,N_17351,N_19785);
xnor U20230 (N_20230,N_16416,N_19739);
and U20231 (N_20231,N_19247,N_18890);
or U20232 (N_20232,N_15466,N_15771);
or U20233 (N_20233,N_19579,N_15388);
nand U20234 (N_20234,N_18694,N_19205);
and U20235 (N_20235,N_15152,N_18431);
nand U20236 (N_20236,N_16374,N_18677);
nand U20237 (N_20237,N_19027,N_18997);
nand U20238 (N_20238,N_16399,N_15261);
xor U20239 (N_20239,N_15220,N_15473);
and U20240 (N_20240,N_17426,N_15497);
nor U20241 (N_20241,N_17219,N_18379);
xor U20242 (N_20242,N_15892,N_19682);
nand U20243 (N_20243,N_17657,N_15361);
nor U20244 (N_20244,N_18993,N_15699);
xor U20245 (N_20245,N_15712,N_16562);
and U20246 (N_20246,N_17073,N_19128);
nand U20247 (N_20247,N_16609,N_15727);
xor U20248 (N_20248,N_19042,N_16559);
xnor U20249 (N_20249,N_15525,N_19640);
xnor U20250 (N_20250,N_17170,N_17566);
nand U20251 (N_20251,N_18842,N_18489);
nand U20252 (N_20252,N_18931,N_17085);
nor U20253 (N_20253,N_17324,N_15159);
and U20254 (N_20254,N_17759,N_19812);
nor U20255 (N_20255,N_15833,N_17493);
nor U20256 (N_20256,N_19334,N_16404);
and U20257 (N_20257,N_18553,N_16308);
nand U20258 (N_20258,N_16604,N_15958);
and U20259 (N_20259,N_19102,N_17475);
xor U20260 (N_20260,N_17988,N_15396);
nor U20261 (N_20261,N_19725,N_16713);
nor U20262 (N_20262,N_18103,N_15226);
and U20263 (N_20263,N_18577,N_15016);
nand U20264 (N_20264,N_15916,N_18423);
or U20265 (N_20265,N_17653,N_18346);
and U20266 (N_20266,N_16208,N_18737);
nand U20267 (N_20267,N_17983,N_17937);
or U20268 (N_20268,N_16734,N_18249);
nand U20269 (N_20269,N_18056,N_15539);
nor U20270 (N_20270,N_17103,N_16855);
and U20271 (N_20271,N_19370,N_18986);
or U20272 (N_20272,N_17784,N_19919);
and U20273 (N_20273,N_17672,N_15224);
nor U20274 (N_20274,N_19414,N_19182);
or U20275 (N_20275,N_15787,N_19613);
and U20276 (N_20276,N_19704,N_18334);
and U20277 (N_20277,N_19336,N_18247);
nor U20278 (N_20278,N_16903,N_18391);
nor U20279 (N_20279,N_15326,N_18757);
nor U20280 (N_20280,N_18829,N_16820);
xnor U20281 (N_20281,N_19889,N_19074);
or U20282 (N_20282,N_19791,N_19954);
xor U20283 (N_20283,N_16967,N_19782);
and U20284 (N_20284,N_17592,N_17003);
and U20285 (N_20285,N_16828,N_15461);
nand U20286 (N_20286,N_17865,N_15762);
xnor U20287 (N_20287,N_18734,N_16557);
xor U20288 (N_20288,N_15836,N_19217);
and U20289 (N_20289,N_18205,N_19741);
and U20290 (N_20290,N_15305,N_19462);
nand U20291 (N_20291,N_19966,N_18416);
nor U20292 (N_20292,N_15357,N_15124);
and U20293 (N_20293,N_15139,N_16387);
nand U20294 (N_20294,N_16645,N_17131);
xor U20295 (N_20295,N_17883,N_16618);
or U20296 (N_20296,N_17168,N_18881);
or U20297 (N_20297,N_17202,N_17890);
nand U20298 (N_20298,N_19632,N_18373);
nor U20299 (N_20299,N_16851,N_18267);
nand U20300 (N_20300,N_18970,N_19787);
xnor U20301 (N_20301,N_15700,N_18796);
nor U20302 (N_20302,N_19727,N_18536);
or U20303 (N_20303,N_18016,N_17590);
and U20304 (N_20304,N_15192,N_16027);
xnor U20305 (N_20305,N_18068,N_17161);
nand U20306 (N_20306,N_19672,N_15398);
and U20307 (N_20307,N_19904,N_16542);
nand U20308 (N_20308,N_15971,N_16878);
nand U20309 (N_20309,N_18771,N_19797);
nor U20310 (N_20310,N_16017,N_19285);
and U20311 (N_20311,N_16499,N_15749);
or U20312 (N_20312,N_17195,N_19988);
nand U20313 (N_20313,N_19784,N_18837);
or U20314 (N_20314,N_16356,N_15337);
and U20315 (N_20315,N_16581,N_19400);
nor U20316 (N_20316,N_18309,N_19515);
and U20317 (N_20317,N_18223,N_16674);
and U20318 (N_20318,N_18865,N_16222);
nand U20319 (N_20319,N_15195,N_19946);
nand U20320 (N_20320,N_18324,N_19348);
and U20321 (N_20321,N_16275,N_16466);
and U20322 (N_20322,N_18973,N_15200);
nand U20323 (N_20323,N_19267,N_15400);
xor U20324 (N_20324,N_17741,N_17379);
nand U20325 (N_20325,N_15670,N_18722);
nand U20326 (N_20326,N_18611,N_17854);
nor U20327 (N_20327,N_18998,N_16591);
xor U20328 (N_20328,N_19722,N_19150);
xor U20329 (N_20329,N_18154,N_19517);
and U20330 (N_20330,N_18541,N_17190);
nand U20331 (N_20331,N_15578,N_19449);
or U20332 (N_20332,N_18697,N_16577);
nand U20333 (N_20333,N_17323,N_19273);
and U20334 (N_20334,N_18586,N_17015);
nand U20335 (N_20335,N_18311,N_19086);
or U20336 (N_20336,N_15312,N_15070);
or U20337 (N_20337,N_18040,N_16190);
and U20338 (N_20338,N_18186,N_16580);
xnor U20339 (N_20339,N_18135,N_16485);
and U20340 (N_20340,N_17457,N_18287);
xor U20341 (N_20341,N_19179,N_16530);
and U20342 (N_20342,N_16699,N_18528);
and U20343 (N_20343,N_16085,N_19851);
or U20344 (N_20344,N_18462,N_15655);
or U20345 (N_20345,N_18785,N_19770);
nor U20346 (N_20346,N_17899,N_19368);
xor U20347 (N_20347,N_18894,N_18344);
nor U20348 (N_20348,N_18696,N_16957);
nor U20349 (N_20349,N_15352,N_16927);
or U20350 (N_20350,N_15959,N_19033);
or U20351 (N_20351,N_19853,N_15030);
or U20352 (N_20352,N_16153,N_19552);
nand U20353 (N_20353,N_16919,N_18962);
or U20354 (N_20354,N_19149,N_19135);
nand U20355 (N_20355,N_19516,N_17449);
or U20356 (N_20356,N_16365,N_17503);
and U20357 (N_20357,N_18901,N_17181);
nand U20358 (N_20358,N_16421,N_17133);
and U20359 (N_20359,N_16917,N_16062);
and U20360 (N_20360,N_18482,N_16265);
nand U20361 (N_20361,N_17160,N_15701);
nor U20362 (N_20362,N_15846,N_15845);
nor U20363 (N_20363,N_16477,N_16707);
nor U20364 (N_20364,N_18636,N_15507);
and U20365 (N_20365,N_15706,N_19991);
and U20366 (N_20366,N_19877,N_17418);
nand U20367 (N_20367,N_17906,N_17187);
xnor U20368 (N_20368,N_15709,N_18824);
and U20369 (N_20369,N_16096,N_17643);
nand U20370 (N_20370,N_16259,N_17610);
xor U20371 (N_20371,N_15066,N_17070);
nand U20372 (N_20372,N_17115,N_17282);
xor U20373 (N_20373,N_18735,N_15284);
nand U20374 (N_20374,N_15933,N_18310);
nor U20375 (N_20375,N_17650,N_18885);
xor U20376 (N_20376,N_17522,N_17430);
xor U20377 (N_20377,N_18503,N_15096);
nor U20378 (N_20378,N_16297,N_18250);
xnor U20379 (N_20379,N_16832,N_17432);
nand U20380 (N_20380,N_15742,N_16091);
nand U20381 (N_20381,N_15536,N_18599);
nand U20382 (N_20382,N_19555,N_18170);
xnor U20383 (N_20383,N_19185,N_19651);
or U20384 (N_20384,N_18882,N_19051);
nor U20385 (N_20385,N_16354,N_19845);
or U20386 (N_20386,N_17315,N_17414);
nor U20387 (N_20387,N_19333,N_15831);
or U20388 (N_20388,N_18245,N_15839);
nor U20389 (N_20389,N_15666,N_19035);
nand U20390 (N_20390,N_16045,N_16574);
or U20391 (N_20391,N_16073,N_17263);
nand U20392 (N_20392,N_19426,N_16601);
nand U20393 (N_20393,N_19294,N_18167);
and U20394 (N_20394,N_15947,N_16705);
nand U20395 (N_20395,N_19160,N_16960);
xor U20396 (N_20396,N_19882,N_15057);
nand U20397 (N_20397,N_17825,N_17357);
nand U20398 (N_20398,N_18277,N_16729);
xnor U20399 (N_20399,N_18494,N_15813);
nand U20400 (N_20400,N_15151,N_19909);
or U20401 (N_20401,N_15103,N_16269);
and U20402 (N_20402,N_17352,N_15427);
xnor U20403 (N_20403,N_19366,N_15963);
and U20404 (N_20404,N_18065,N_19117);
nand U20405 (N_20405,N_17270,N_17442);
nor U20406 (N_20406,N_17177,N_15537);
nand U20407 (N_20407,N_19013,N_19362);
or U20408 (N_20408,N_18328,N_15876);
nand U20409 (N_20409,N_15179,N_17604);
nor U20410 (N_20410,N_16901,N_17482);
or U20411 (N_20411,N_15572,N_19709);
or U20412 (N_20412,N_18836,N_17809);
or U20413 (N_20413,N_16053,N_18107);
nor U20414 (N_20414,N_15743,N_18369);
or U20415 (N_20415,N_19046,N_18670);
and U20416 (N_20416,N_18396,N_19393);
nor U20417 (N_20417,N_19507,N_18092);
nand U20418 (N_20418,N_15977,N_18165);
and U20419 (N_20419,N_16461,N_19742);
and U20420 (N_20420,N_17742,N_17728);
nor U20421 (N_20421,N_18121,N_16108);
nand U20422 (N_20422,N_17665,N_15456);
nand U20423 (N_20423,N_15084,N_17434);
nor U20424 (N_20424,N_15095,N_18362);
nor U20425 (N_20425,N_19595,N_19148);
xor U20426 (N_20426,N_15693,N_15882);
nor U20427 (N_20427,N_18448,N_18905);
xnor U20428 (N_20428,N_19886,N_16615);
xor U20429 (N_20429,N_19983,N_19575);
nor U20430 (N_20430,N_19808,N_16972);
or U20431 (N_20431,N_18858,N_15680);
nand U20432 (N_20432,N_19208,N_19069);
nor U20433 (N_20433,N_17750,N_19728);
nor U20434 (N_20434,N_19805,N_16513);
nor U20435 (N_20435,N_16464,N_17212);
nor U20436 (N_20436,N_16106,N_15136);
xor U20437 (N_20437,N_17952,N_18280);
or U20438 (N_20438,N_17498,N_18699);
or U20439 (N_20439,N_15127,N_18866);
or U20440 (N_20440,N_19082,N_15667);
xor U20441 (N_20441,N_17818,N_17030);
nor U20442 (N_20442,N_15955,N_17833);
xor U20443 (N_20443,N_18318,N_15395);
and U20444 (N_20444,N_16228,N_17364);
nor U20445 (N_20445,N_17958,N_16300);
or U20446 (N_20446,N_18215,N_17303);
or U20447 (N_20447,N_17327,N_16517);
and U20448 (N_20448,N_18412,N_17329);
nor U20449 (N_20449,N_16163,N_19170);
and U20450 (N_20450,N_17125,N_16555);
and U20451 (N_20451,N_17039,N_15843);
xnor U20452 (N_20452,N_17888,N_18459);
nand U20453 (N_20453,N_19880,N_19227);
and U20454 (N_20454,N_15778,N_17684);
nor U20455 (N_20455,N_16650,N_19373);
nor U20456 (N_20456,N_16997,N_18152);
or U20457 (N_20457,N_15596,N_15899);
nor U20458 (N_20458,N_17628,N_18199);
or U20459 (N_20459,N_18230,N_16336);
nor U20460 (N_20460,N_17796,N_17144);
nand U20461 (N_20461,N_18701,N_17147);
nand U20462 (N_20462,N_18384,N_17708);
xnor U20463 (N_20463,N_16446,N_18915);
xnor U20464 (N_20464,N_17365,N_16143);
nor U20465 (N_20465,N_18875,N_16671);
xor U20466 (N_20466,N_19761,N_15601);
nand U20467 (N_20467,N_18870,N_15587);
nor U20468 (N_20468,N_18397,N_17071);
xor U20469 (N_20469,N_17569,N_15271);
nor U20470 (N_20470,N_19162,N_18429);
nand U20471 (N_20471,N_17975,N_15552);
nor U20472 (N_20472,N_18254,N_15624);
xnor U20473 (N_20473,N_19015,N_19476);
xnor U20474 (N_20474,N_15588,N_17688);
nor U20475 (N_20475,N_19643,N_18990);
nor U20476 (N_20476,N_16059,N_19884);
and U20477 (N_20477,N_18233,N_19095);
and U20478 (N_20478,N_19809,N_16250);
nor U20479 (N_20479,N_17753,N_15409);
and U20480 (N_20480,N_17021,N_17246);
and U20481 (N_20481,N_19079,N_16738);
nor U20482 (N_20482,N_16947,N_17420);
nand U20483 (N_20483,N_19447,N_16225);
xor U20484 (N_20484,N_16926,N_16286);
nand U20485 (N_20485,N_15920,N_15335);
or U20486 (N_20486,N_18868,N_16605);
or U20487 (N_20487,N_19685,N_17695);
nor U20488 (N_20488,N_16692,N_17281);
and U20489 (N_20489,N_15717,N_18234);
or U20490 (N_20490,N_18030,N_17981);
xnor U20491 (N_20491,N_19733,N_19895);
nand U20492 (N_20492,N_18827,N_19836);
nand U20493 (N_20493,N_15766,N_16592);
nand U20494 (N_20494,N_16802,N_17174);
nor U20495 (N_20495,N_15049,N_16904);
xor U20496 (N_20496,N_19315,N_18687);
nor U20497 (N_20497,N_15840,N_16029);
and U20498 (N_20498,N_18929,N_17463);
and U20499 (N_20499,N_15472,N_17269);
or U20500 (N_20500,N_16685,N_17640);
nand U20501 (N_20501,N_17659,N_15330);
and U20502 (N_20502,N_16274,N_17156);
and U20503 (N_20503,N_18213,N_15993);
nor U20504 (N_20504,N_17157,N_15107);
nor U20505 (N_20505,N_18823,N_18758);
xor U20506 (N_20506,N_15652,N_16491);
xor U20507 (N_20507,N_18647,N_17940);
xnor U20508 (N_20508,N_19662,N_17391);
xor U20509 (N_20509,N_17524,N_15309);
nand U20510 (N_20510,N_18392,N_17835);
and U20511 (N_20511,N_17436,N_16318);
nor U20512 (N_20512,N_15505,N_17114);
nor U20513 (N_20513,N_17013,N_18927);
nand U20514 (N_20514,N_17469,N_18675);
nor U20515 (N_20515,N_17830,N_15039);
and U20516 (N_20516,N_15443,N_17902);
nand U20517 (N_20517,N_19008,N_17452);
xnor U20518 (N_20518,N_15557,N_15338);
nand U20519 (N_20519,N_18394,N_19671);
nand U20520 (N_20520,N_19313,N_18809);
or U20521 (N_20521,N_17954,N_19949);
xor U20522 (N_20522,N_15355,N_15117);
or U20523 (N_20523,N_16011,N_15341);
nand U20524 (N_20524,N_18279,N_18640);
xor U20525 (N_20525,N_18359,N_19798);
or U20526 (N_20526,N_15339,N_16603);
nor U20527 (N_20527,N_19299,N_18691);
nor U20528 (N_20528,N_16864,N_17961);
or U20529 (N_20529,N_17053,N_15079);
and U20530 (N_20530,N_19747,N_15054);
or U20531 (N_20531,N_18849,N_15968);
nand U20532 (N_20532,N_19527,N_17109);
or U20533 (N_20533,N_19283,N_19113);
nor U20534 (N_20534,N_16771,N_18864);
nand U20535 (N_20535,N_17691,N_18500);
nand U20536 (N_20536,N_15036,N_19311);
and U20537 (N_20537,N_19199,N_15878);
and U20538 (N_20538,N_18343,N_19252);
nor U20539 (N_20539,N_19018,N_18919);
or U20540 (N_20540,N_16563,N_19612);
nor U20541 (N_20541,N_15736,N_17294);
or U20542 (N_20542,N_17126,N_16649);
nor U20543 (N_20543,N_18399,N_19953);
or U20544 (N_20544,N_19970,N_19151);
nand U20545 (N_20545,N_19464,N_19374);
nand U20546 (N_20546,N_15938,N_19591);
nand U20547 (N_20547,N_17683,N_19410);
nor U20548 (N_20548,N_18521,N_15092);
or U20549 (N_20549,N_19532,N_17433);
nand U20550 (N_20550,N_15917,N_15754);
and U20551 (N_20551,N_17056,N_19164);
xor U20552 (N_20552,N_19006,N_15730);
nand U20553 (N_20553,N_19657,N_16347);
nand U20554 (N_20554,N_16929,N_18138);
and U20555 (N_20555,N_17558,N_16543);
xnor U20556 (N_20556,N_15223,N_15931);
or U20557 (N_20557,N_18830,N_19307);
nor U20558 (N_20558,N_16545,N_17250);
and U20559 (N_20559,N_17668,N_16980);
nand U20560 (N_20560,N_17220,N_17968);
or U20561 (N_20561,N_16352,N_19619);
nand U20562 (N_20562,N_19813,N_19523);
and U20563 (N_20563,N_17359,N_18921);
or U20564 (N_20564,N_18219,N_17296);
nor U20565 (N_20565,N_18810,N_16401);
nand U20566 (N_20566,N_17550,N_15751);
nand U20567 (N_20567,N_15932,N_17374);
xnor U20568 (N_20568,N_15984,N_15173);
nand U20569 (N_20569,N_19467,N_18840);
or U20570 (N_20570,N_16490,N_15969);
nor U20571 (N_20571,N_17384,N_17360);
and U20572 (N_20572,N_15351,N_19021);
xnor U20573 (N_20573,N_19901,N_17380);
nor U20574 (N_20574,N_19203,N_16141);
and U20575 (N_20575,N_17051,N_15163);
nor U20576 (N_20576,N_18910,N_19219);
xor U20577 (N_20577,N_18545,N_18017);
nor U20578 (N_20578,N_15385,N_18617);
or U20579 (N_20579,N_17142,N_15503);
nor U20580 (N_20580,N_15704,N_15896);
nand U20581 (N_20581,N_18237,N_18368);
nand U20582 (N_20582,N_18512,N_17705);
nor U20583 (N_20583,N_19881,N_18579);
nand U20584 (N_20584,N_15682,N_16339);
and U20585 (N_20585,N_19098,N_18683);
xnor U20586 (N_20586,N_18641,N_18556);
or U20587 (N_20587,N_19636,N_19019);
nand U20588 (N_20588,N_19865,N_19956);
nand U20589 (N_20589,N_19498,N_18447);
xor U20590 (N_20590,N_15553,N_15716);
and U20591 (N_20591,N_17630,N_18496);
xnor U20592 (N_20592,N_15803,N_19132);
and U20593 (N_20593,N_15435,N_17673);
xor U20594 (N_20594,N_19550,N_19239);
xor U20595 (N_20595,N_16012,N_18578);
or U20596 (N_20596,N_19123,N_16094);
nor U20597 (N_20597,N_19661,N_19978);
nand U20598 (N_20598,N_16964,N_15818);
or U20599 (N_20599,N_19676,N_19876);
and U20600 (N_20600,N_18896,N_19639);
and U20601 (N_20601,N_18454,N_15210);
nand U20602 (N_20602,N_16742,N_15207);
and U20603 (N_20603,N_15614,N_17476);
nor U20604 (N_20604,N_15964,N_15617);
nor U20605 (N_20605,N_16170,N_16410);
nand U20606 (N_20606,N_18895,N_18679);
xnor U20607 (N_20607,N_15992,N_19226);
nor U20608 (N_20608,N_19246,N_19277);
xnor U20609 (N_20609,N_18793,N_19980);
and U20610 (N_20610,N_19286,N_16983);
or U20611 (N_20611,N_18658,N_16546);
or U20612 (N_20612,N_19945,N_15496);
xnor U20613 (N_20613,N_15633,N_17893);
or U20614 (N_20614,N_16188,N_17892);
xor U20615 (N_20615,N_18071,N_18926);
xnor U20616 (N_20616,N_19260,N_16932);
nand U20617 (N_20617,N_17251,N_16859);
xor U20618 (N_20618,N_16669,N_17225);
nor U20619 (N_20619,N_19300,N_19450);
nor U20620 (N_20620,N_17853,N_17516);
and U20621 (N_20621,N_18531,N_15362);
nand U20622 (N_20622,N_16041,N_19794);
nand U20623 (N_20623,N_19134,N_18404);
nor U20624 (N_20624,N_19716,N_16719);
or U20625 (N_20625,N_15068,N_15297);
xnor U20626 (N_20626,N_19630,N_19793);
or U20627 (N_20627,N_19064,N_15157);
and U20628 (N_20628,N_19665,N_18060);
nor U20629 (N_20629,N_19180,N_19585);
and U20630 (N_20630,N_16614,N_16001);
and U20631 (N_20631,N_17172,N_16687);
or U20632 (N_20632,N_16092,N_16607);
or U20633 (N_20633,N_15042,N_15268);
and U20634 (N_20634,N_16970,N_19828);
nor U20635 (N_20635,N_17423,N_15040);
xor U20636 (N_20636,N_19934,N_18468);
and U20637 (N_20637,N_17306,N_17465);
or U20638 (N_20638,N_15249,N_16816);
and U20639 (N_20639,N_16821,N_19707);
nand U20640 (N_20640,N_16758,N_15015);
nor U20641 (N_20641,N_16831,N_16024);
nand U20642 (N_20642,N_17487,N_17454);
xor U20643 (N_20643,N_17072,N_17740);
nand U20644 (N_20644,N_17593,N_15528);
xor U20645 (N_20645,N_15188,N_15907);
xnor U20646 (N_20646,N_17941,N_16303);
xor U20647 (N_20647,N_18440,N_18904);
xnor U20648 (N_20648,N_17047,N_19620);
and U20649 (N_20649,N_16294,N_15559);
nor U20650 (N_20650,N_17209,N_19669);
and U20651 (N_20651,N_15834,N_17764);
nor U20652 (N_20652,N_16224,N_19188);
and U20653 (N_20653,N_15577,N_16140);
xnor U20654 (N_20654,N_16536,N_16965);
and U20655 (N_20655,N_18284,N_16406);
or U20656 (N_20656,N_18834,N_18777);
and U20657 (N_20657,N_16666,N_15368);
and U20658 (N_20658,N_17858,N_19960);
nor U20659 (N_20659,N_16060,N_17489);
nand U20660 (N_20660,N_18720,N_17811);
and U20661 (N_20661,N_19327,N_18288);
and U20662 (N_20662,N_16962,N_17381);
nand U20663 (N_20663,N_19864,N_19110);
nor U20664 (N_20664,N_19874,N_16372);
and U20665 (N_20665,N_18326,N_15295);
nor U20666 (N_20666,N_15181,N_16884);
and U20667 (N_20667,N_18769,N_16797);
and U20668 (N_20668,N_19985,N_17377);
or U20669 (N_20669,N_18316,N_18374);
or U20670 (N_20670,N_18211,N_15806);
or U20671 (N_20671,N_18090,N_15511);
nand U20672 (N_20672,N_16182,N_19850);
and U20673 (N_20673,N_18583,N_18356);
nor U20674 (N_20674,N_15741,N_15177);
nand U20675 (N_20675,N_19560,N_16009);
nand U20676 (N_20676,N_19952,N_19424);
nand U20677 (N_20677,N_18465,N_19003);
nand U20678 (N_20678,N_17197,N_17602);
nand U20679 (N_20679,N_16830,N_16500);
or U20680 (N_20680,N_16373,N_18897);
and U20681 (N_20681,N_17778,N_17416);
xor U20682 (N_20682,N_17611,N_17955);
or U20683 (N_20683,N_15894,N_18988);
or U20684 (N_20684,N_15174,N_17837);
nand U20685 (N_20685,N_17586,N_19868);
xnor U20686 (N_20686,N_17798,N_16768);
nor U20687 (N_20687,N_15424,N_17900);
or U20688 (N_20688,N_15924,N_18192);
or U20689 (N_20689,N_16602,N_15078);
or U20690 (N_20690,N_17664,N_15399);
xnor U20691 (N_20691,N_16754,N_17361);
nor U20692 (N_20692,N_17887,N_18143);
nand U20693 (N_20693,N_17661,N_18383);
nor U20694 (N_20694,N_16829,N_17207);
nand U20695 (N_20695,N_15850,N_17300);
nand U20696 (N_20696,N_16020,N_18805);
or U20697 (N_20697,N_19838,N_15026);
and U20698 (N_20698,N_17878,N_16777);
nand U20699 (N_20699,N_15007,N_19174);
or U20700 (N_20700,N_18618,N_15046);
and U20701 (N_20701,N_15990,N_15780);
or U20702 (N_20702,N_18021,N_19766);
nand U20703 (N_20703,N_19903,N_18477);
xor U20704 (N_20704,N_16202,N_17277);
or U20705 (N_20705,N_16589,N_18037);
nor U20706 (N_20706,N_16739,N_17155);
xor U20707 (N_20707,N_17621,N_15897);
nand U20708 (N_20708,N_18936,N_17553);
xor U20709 (N_20709,N_17545,N_19627);
nor U20710 (N_20710,N_16216,N_16690);
nor U20711 (N_20711,N_18937,N_15793);
xor U20712 (N_20712,N_17584,N_16146);
and U20713 (N_20713,N_17897,N_16238);
and U20714 (N_20714,N_18438,N_16572);
nand U20715 (N_20715,N_18698,N_17976);
xor U20716 (N_20716,N_17852,N_19660);
and U20717 (N_20717,N_15562,N_19175);
and U20718 (N_20718,N_15711,N_19503);
nor U20719 (N_20719,N_15657,N_16850);
xnor U20720 (N_20720,N_19989,N_19140);
and U20721 (N_20721,N_18801,N_19763);
and U20722 (N_20722,N_15239,N_15343);
nand U20723 (N_20723,N_15314,N_18702);
or U20724 (N_20724,N_17757,N_15989);
nor U20725 (N_20725,N_16746,N_17256);
xor U20726 (N_20726,N_16116,N_17529);
and U20727 (N_20727,N_15895,N_18592);
nand U20728 (N_20728,N_15486,N_17831);
nor U20729 (N_20729,N_18576,N_19648);
and U20730 (N_20730,N_17652,N_16912);
xnor U20731 (N_20731,N_16346,N_16987);
and U20732 (N_20732,N_17868,N_19428);
nor U20733 (N_20733,N_19559,N_15903);
or U20734 (N_20734,N_17235,N_17367);
nand U20735 (N_20735,N_17192,N_19890);
nor U20736 (N_20736,N_15439,N_18243);
and U20737 (N_20737,N_19119,N_16570);
and U20738 (N_20738,N_15886,N_17271);
xnor U20739 (N_20739,N_15654,N_15915);
and U20740 (N_20740,N_18332,N_15692);
xor U20741 (N_20741,N_16214,N_17577);
xor U20742 (N_20742,N_16348,N_18042);
or U20743 (N_20743,N_16281,N_19948);
nand U20744 (N_20744,N_19025,N_17689);
nand U20745 (N_20745,N_15438,N_15272);
and U20746 (N_20746,N_19769,N_19557);
xnor U20747 (N_20747,N_18228,N_16474);
and U20748 (N_20748,N_17971,N_19646);
nor U20749 (N_20749,N_17194,N_16008);
nor U20750 (N_20750,N_19212,N_18732);
or U20751 (N_20751,N_16873,N_17092);
or U20752 (N_20752,N_17501,N_17614);
nand U20753 (N_20753,N_19717,N_18061);
or U20754 (N_20754,N_16946,N_18417);
xnor U20755 (N_20755,N_19513,N_17995);
and U20756 (N_20756,N_15364,N_18948);
nor U20757 (N_20757,N_18450,N_16872);
or U20758 (N_20758,N_16005,N_15595);
nand U20759 (N_20759,N_19118,N_16249);
and U20760 (N_20760,N_18822,N_17677);
or U20761 (N_20761,N_15237,N_18315);
xor U20762 (N_20762,N_16328,N_16633);
or U20763 (N_20763,N_19652,N_18520);
or U20764 (N_20764,N_16928,N_15558);
or U20765 (N_20765,N_15939,N_19167);
nand U20766 (N_20766,N_15530,N_16313);
and U20767 (N_20767,N_17946,N_17169);
and U20768 (N_20768,N_17078,N_16069);
xnor U20769 (N_20769,N_17046,N_16428);
nor U20770 (N_20770,N_19255,N_19814);
xnor U20771 (N_20771,N_19365,N_19654);
nor U20772 (N_20772,N_18387,N_15111);
xor U20773 (N_20773,N_15346,N_15475);
nor U20774 (N_20774,N_17844,N_16748);
and U20775 (N_20775,N_16244,N_15085);
nand U20776 (N_20776,N_15452,N_18091);
xnor U20777 (N_20777,N_15687,N_15051);
xnor U20778 (N_20778,N_16891,N_15865);
xnor U20779 (N_20779,N_17507,N_19415);
or U20780 (N_20780,N_19533,N_15300);
nor U20781 (N_20781,N_15281,N_19887);
and U20782 (N_20782,N_15073,N_16353);
xnor U20783 (N_20783,N_19153,N_15921);
and U20784 (N_20784,N_15069,N_15866);
and U20785 (N_20785,N_19391,N_17456);
nand U20786 (N_20786,N_16192,N_19201);
nor U20787 (N_20787,N_18664,N_17531);
or U20788 (N_20788,N_19911,N_17536);
and U20789 (N_20789,N_18740,N_17285);
or U20790 (N_20790,N_18883,N_16658);
nor U20791 (N_20791,N_19981,N_19899);
and U20792 (N_20792,N_19099,N_16414);
nor U20793 (N_20793,N_15203,N_17979);
xor U20794 (N_20794,N_16121,N_15918);
and U20795 (N_20795,N_16393,N_15566);
nor U20796 (N_20796,N_16462,N_18437);
nor U20797 (N_20797,N_16098,N_15334);
xor U20798 (N_20798,N_15052,N_16044);
or U20799 (N_20799,N_17776,N_16956);
nor U20800 (N_20800,N_17974,N_19873);
nor U20801 (N_20801,N_16129,N_19198);
nand U20802 (N_20802,N_19641,N_16778);
nor U20803 (N_20803,N_16256,N_17260);
xor U20804 (N_20804,N_17288,N_18790);
or U20805 (N_20805,N_16114,N_16123);
or U20806 (N_20806,N_17690,N_16436);
or U20807 (N_20807,N_19121,N_15733);
xor U20808 (N_20808,N_19680,N_17121);
nand U20809 (N_20809,N_17894,N_17143);
nand U20810 (N_20810,N_16324,N_19216);
or U20811 (N_20811,N_19233,N_15492);
nand U20812 (N_20812,N_18289,N_18003);
xnor U20813 (N_20813,N_16755,N_16405);
xnor U20814 (N_20814,N_17856,N_15695);
xnor U20815 (N_20815,N_16717,N_18530);
nand U20816 (N_20816,N_16223,N_17514);
nand U20817 (N_20817,N_15176,N_17350);
or U20818 (N_20818,N_18933,N_16148);
xor U20819 (N_20819,N_15521,N_15582);
and U20820 (N_20820,N_16656,N_17108);
nor U20821 (N_20821,N_17960,N_19837);
or U20822 (N_20822,N_15285,N_19461);
nand U20823 (N_20823,N_18028,N_19379);
nor U20824 (N_20824,N_18148,N_19692);
or U20825 (N_20825,N_19249,N_15194);
and U20826 (N_20826,N_15128,N_17206);
nand U20827 (N_20827,N_18015,N_18749);
or U20828 (N_20828,N_18109,N_18625);
nand U20829 (N_20829,N_18922,N_18084);
nand U20830 (N_20830,N_19062,N_18045);
and U20831 (N_20831,N_15949,N_15631);
nor U20832 (N_20832,N_18772,N_17404);
xnor U20833 (N_20833,N_16978,N_18686);
or U20834 (N_20834,N_17580,N_16392);
xnor U20835 (N_20835,N_17074,N_15367);
nor U20836 (N_20836,N_17000,N_19854);
and U20837 (N_20837,N_16529,N_15615);
nand U20838 (N_20838,N_19404,N_15148);
nor U20839 (N_20839,N_18709,N_16803);
and U20840 (N_20840,N_19290,N_16310);
and U20841 (N_20841,N_17328,N_16684);
and U20842 (N_20842,N_17716,N_18716);
xor U20843 (N_20843,N_17088,N_16200);
or U20844 (N_20844,N_15792,N_19029);
xnor U20845 (N_20845,N_17623,N_16282);
nor U20846 (N_20846,N_15360,N_18158);
and U20847 (N_20847,N_17512,N_19012);
or U20848 (N_20848,N_18041,N_18166);
nor U20849 (N_20849,N_19332,N_17459);
nor U20850 (N_20850,N_18018,N_16145);
xor U20851 (N_20851,N_16086,N_16230);
xor U20852 (N_20852,N_17470,N_17783);
nand U20853 (N_20853,N_17918,N_17726);
or U20854 (N_20854,N_17004,N_18002);
and U20855 (N_20855,N_17441,N_19969);
and U20856 (N_20856,N_17189,N_19618);
or U20857 (N_20857,N_19542,N_15450);
or U20858 (N_20858,N_19920,N_19546);
or U20859 (N_20859,N_17967,N_17719);
nor U20860 (N_20860,N_16642,N_19556);
nand U20861 (N_20861,N_15238,N_17034);
and U20862 (N_20862,N_19196,N_19491);
or U20863 (N_20863,N_18043,N_15563);
xnor U20864 (N_20864,N_16682,N_15950);
and U20865 (N_20865,N_15340,N_19584);
and U20866 (N_20866,N_16955,N_15083);
and U20867 (N_20867,N_17625,N_19269);
nand U20868 (N_20868,N_17540,N_15777);
and U20869 (N_20869,N_18377,N_19284);
and U20870 (N_20870,N_17933,N_15729);
xnor U20871 (N_20871,N_18776,N_15669);
nor U20872 (N_20872,N_15391,N_17375);
or U20873 (N_20873,N_18903,N_18360);
and U20874 (N_20874,N_18202,N_15208);
nand U20875 (N_20875,N_18285,N_19416);
xor U20876 (N_20876,N_19126,N_18628);
xor U20877 (N_20877,N_15602,N_18323);
or U20878 (N_20878,N_17654,N_19628);
xor U20879 (N_20879,N_16049,N_19061);
nor U20880 (N_20880,N_16135,N_19633);
xor U20881 (N_20881,N_18767,N_19653);
nand U20882 (N_20882,N_19861,N_16470);
nand U20883 (N_20883,N_19496,N_19615);
nor U20884 (N_20884,N_17309,N_15211);
or U20885 (N_20885,N_15436,N_19041);
nor U20886 (N_20886,N_16866,N_15373);
and U20887 (N_20887,N_15725,N_18680);
and U20888 (N_20888,N_15019,N_18433);
nand U20889 (N_20889,N_19420,N_18820);
and U20890 (N_20890,N_18442,N_18811);
nand U20891 (N_20891,N_16568,N_17435);
xor U20892 (N_20892,N_15746,N_18597);
nand U20893 (N_20893,N_18632,N_17782);
xnor U20894 (N_20894,N_17100,N_18833);
and U20895 (N_20895,N_15997,N_18480);
and U20896 (N_20896,N_17388,N_19531);
or U20897 (N_20897,N_15826,N_16055);
xor U20898 (N_20898,N_19004,N_19663);
nand U20899 (N_20899,N_18928,N_15493);
xor U20900 (N_20900,N_18006,N_17424);
nand U20901 (N_20901,N_17660,N_18891);
nand U20902 (N_20902,N_19242,N_19724);
nand U20903 (N_20903,N_17747,N_15043);
nand U20904 (N_20904,N_15202,N_17244);
and U20905 (N_20905,N_19437,N_17042);
or U20906 (N_20906,N_15513,N_17624);
or U20907 (N_20907,N_15468,N_19353);
nand U20908 (N_20908,N_18765,N_16457);
nand U20909 (N_20909,N_18376,N_17509);
and U20910 (N_20910,N_17763,N_15319);
nand U20911 (N_20911,N_18571,N_17836);
and U20912 (N_20912,N_17107,N_16804);
xor U20913 (N_20913,N_17775,N_18491);
nand U20914 (N_20914,N_19258,N_18703);
xor U20915 (N_20915,N_18341,N_16206);
nor U20916 (N_20916,N_15807,N_15518);
nand U20917 (N_20917,N_15256,N_15752);
xor U20918 (N_20918,N_16694,N_18338);
and U20919 (N_20919,N_16367,N_19186);
or U20920 (N_20920,N_17334,N_16770);
nand U20921 (N_20921,N_19264,N_17287);
xor U20922 (N_20922,N_16982,N_19408);
or U20923 (N_20923,N_18569,N_19230);
or U20924 (N_20924,N_17237,N_16627);
nor U20925 (N_20925,N_17697,N_19576);
xnor U20926 (N_20926,N_15278,N_17082);
and U20927 (N_20927,N_19432,N_18780);
nand U20928 (N_20928,N_18196,N_19104);
and U20929 (N_20929,N_16056,N_18744);
xor U20930 (N_20930,N_15158,N_17325);
xor U20931 (N_20931,N_17720,N_17236);
nor U20932 (N_20932,N_18032,N_18710);
or U20933 (N_20933,N_19699,N_17977);
or U20934 (N_20934,N_19898,N_19536);
nor U20935 (N_20935,N_15668,N_18420);
nor U20936 (N_20936,N_15543,N_16359);
xor U20937 (N_20937,N_16906,N_16939);
nor U20938 (N_20938,N_17845,N_16254);
nor U20939 (N_20939,N_17140,N_18204);
xnor U20940 (N_20940,N_18455,N_18770);
nor U20941 (N_20941,N_18128,N_18814);
nand U20942 (N_20942,N_18181,N_17028);
xnor U20943 (N_20943,N_16887,N_15244);
xnor U20944 (N_20944,N_16807,N_17521);
nor U20945 (N_20945,N_16280,N_18161);
xor U20946 (N_20946,N_19698,N_16246);
xor U20947 (N_20947,N_19875,N_16842);
and U20948 (N_20948,N_19405,N_16524);
xnor U20949 (N_20949,N_18445,N_16325);
or U20950 (N_20950,N_19977,N_15485);
and U20951 (N_20951,N_18461,N_19161);
and U20952 (N_20952,N_15758,N_15166);
and U20953 (N_20953,N_18940,N_19352);
and U20954 (N_20954,N_19077,N_16078);
nand U20955 (N_20955,N_18449,N_17738);
nand U20956 (N_20956,N_19765,N_17787);
and U20957 (N_20957,N_16712,N_18631);
xor U20958 (N_20958,N_16333,N_18393);
xnor U20959 (N_20959,N_17166,N_17466);
nor U20960 (N_20960,N_16537,N_15800);
xnor U20961 (N_20961,N_16180,N_17780);
or U20962 (N_20962,N_18038,N_17376);
and U20963 (N_20963,N_15106,N_17838);
and U20964 (N_20964,N_15479,N_18020);
and U20965 (N_20965,N_18129,N_15647);
and U20966 (N_20966,N_15047,N_19923);
and U20967 (N_20967,N_17619,N_17910);
nand U20968 (N_20968,N_18876,N_16047);
nand U20969 (N_20969,N_17029,N_18612);
and U20970 (N_20970,N_18839,N_16877);
xor U20971 (N_20971,N_19635,N_16657);
and U20972 (N_20972,N_18402,N_17385);
nand U20973 (N_20973,N_19122,N_16341);
nor U20974 (N_20974,N_15515,N_18983);
nor U20975 (N_20975,N_19647,N_18502);
nand U20976 (N_20976,N_18013,N_19145);
nand U20977 (N_20977,N_16165,N_17552);
or U20978 (N_20978,N_15359,N_15411);
and U20979 (N_20979,N_15109,N_15764);
nand U20980 (N_20980,N_19528,N_18867);
and U20981 (N_20981,N_19136,N_18231);
xnor U20982 (N_20982,N_19959,N_16700);
nor U20983 (N_20983,N_16285,N_18902);
nor U20984 (N_20984,N_19036,N_18813);
nand U20985 (N_20985,N_18140,N_16370);
and U20986 (N_20986,N_17468,N_16198);
and U20987 (N_20987,N_17973,N_16827);
and U20988 (N_20988,N_16293,N_19081);
nor U20989 (N_20989,N_16305,N_16668);
nor U20990 (N_20990,N_15191,N_19438);
nand U20991 (N_20991,N_19089,N_16902);
nor U20992 (N_20992,N_19377,N_17467);
or U20993 (N_20993,N_19459,N_15451);
nand U20994 (N_20994,N_15254,N_16935);
and U20995 (N_20995,N_15458,N_18144);
xor U20996 (N_20996,N_19356,N_17183);
or U20997 (N_20997,N_17123,N_18914);
xnor U20998 (N_20998,N_19572,N_16507);
xor U20999 (N_20999,N_15906,N_16233);
xnor U21000 (N_21000,N_15410,N_18657);
nand U21001 (N_21001,N_17484,N_16824);
and U21002 (N_21002,N_18409,N_17713);
nor U21003 (N_21003,N_18481,N_17725);
and U21004 (N_21004,N_16397,N_18786);
nor U21005 (N_21005,N_18444,N_18093);
xor U21006 (N_21006,N_16409,N_18164);
or U21007 (N_21007,N_15215,N_15090);
or U21008 (N_21008,N_16331,N_16523);
xnor U21009 (N_21009,N_18863,N_16101);
or U21010 (N_21010,N_17638,N_19427);
nand U21011 (N_21011,N_15286,N_16834);
xnor U21012 (N_21012,N_16167,N_15618);
xor U21013 (N_21013,N_17876,N_16954);
nand U21014 (N_21014,N_16398,N_18117);
or U21015 (N_21015,N_19138,N_16667);
xnor U21016 (N_21016,N_15178,N_15801);
nand U21017 (N_21017,N_16102,N_17448);
xor U21018 (N_21018,N_17171,N_15429);
nand U21019 (N_21019,N_15823,N_17912);
nand U21020 (N_21020,N_16488,N_18000);
or U21021 (N_21021,N_19835,N_16276);
xnor U21022 (N_21022,N_15970,N_19448);
or U21023 (N_21023,N_18363,N_19291);
nand U21024 (N_21024,N_19346,N_16579);
xnor U21025 (N_21025,N_15745,N_15062);
or U21026 (N_21026,N_18352,N_15772);
and U21027 (N_21027,N_17895,N_15842);
and U21028 (N_21028,N_15252,N_15967);
and U21029 (N_21029,N_15469,N_18932);
and U21030 (N_21030,N_16252,N_15001);
nor U21031 (N_21031,N_18862,N_15162);
and U21032 (N_21032,N_17739,N_18802);
nand U21033 (N_21033,N_18422,N_18187);
nand U21034 (N_21034,N_15126,N_15265);
and U21035 (N_21035,N_15779,N_16582);
nand U21036 (N_21036,N_17820,N_19244);
nor U21037 (N_21037,N_18987,N_18008);
nor U21038 (N_21038,N_19254,N_19083);
and U21039 (N_21039,N_19381,N_19343);
xnor U21040 (N_21040,N_16766,N_15763);
nand U21041 (N_21041,N_15196,N_18039);
and U21042 (N_21042,N_18248,N_17336);
xor U21043 (N_21043,N_16168,N_15214);
nand U21044 (N_21044,N_18705,N_16362);
and U21045 (N_21045,N_15642,N_15476);
xnor U21046 (N_21046,N_19674,N_15634);
nand U21047 (N_21047,N_18077,N_17358);
xnor U21048 (N_21048,N_19440,N_18292);
nand U21049 (N_21049,N_17679,N_19279);
or U21050 (N_21050,N_15097,N_16723);
xor U21051 (N_21051,N_17186,N_18952);
and U21052 (N_21052,N_15756,N_18872);
and U21053 (N_21053,N_16454,N_18766);
nor U21054 (N_21054,N_19451,N_19802);
and U21055 (N_21055,N_16934,N_18819);
nand U21056 (N_21056,N_16361,N_18678);
nor U21057 (N_21057,N_19047,N_15227);
nand U21058 (N_21058,N_15371,N_19735);
xnor U21059 (N_21059,N_19715,N_18515);
nand U21060 (N_21060,N_16037,N_17167);
nand U21061 (N_21061,N_18498,N_15626);
nor U21062 (N_21062,N_19376,N_16968);
and U21063 (N_21063,N_16569,N_17901);
or U21064 (N_21064,N_17935,N_17962);
and U21065 (N_21065,N_19604,N_16844);
nand U21066 (N_21066,N_16641,N_19573);
or U21067 (N_21067,N_17427,N_16921);
or U21068 (N_21068,N_17129,N_16992);
or U21069 (N_21069,N_16584,N_15978);
nand U21070 (N_21070,N_15287,N_17258);
or U21071 (N_21071,N_19107,N_17065);
xor U21072 (N_21072,N_15713,N_15358);
nor U21073 (N_21073,N_19187,N_19070);
and U21074 (N_21074,N_17575,N_15625);
nor U21075 (N_21075,N_19968,N_19056);
nor U21076 (N_21076,N_17247,N_18714);
or U21077 (N_21077,N_16295,N_16363);
nor U21078 (N_21078,N_16632,N_18298);
or U21079 (N_21079,N_15639,N_17370);
or U21080 (N_21080,N_18262,N_16506);
and U21081 (N_21081,N_18974,N_16417);
or U21082 (N_21082,N_16971,N_16698);
and U21083 (N_21083,N_17389,N_19992);
xor U21084 (N_21084,N_17733,N_19384);
nor U21085 (N_21085,N_16082,N_16590);
nor U21086 (N_21086,N_15282,N_19441);
nor U21087 (N_21087,N_19038,N_18001);
or U21088 (N_21088,N_18598,N_15887);
nand U21089 (N_21089,N_16438,N_18194);
xor U21090 (N_21090,N_19551,N_17314);
and U21091 (N_21091,N_16587,N_18860);
nand U21092 (N_21092,N_18011,N_18949);
or U21093 (N_21093,N_19407,N_18708);
and U21094 (N_21094,N_18069,N_19078);
and U21095 (N_21095,N_18746,N_18335);
or U21096 (N_21096,N_17266,N_17310);
xor U21097 (N_21097,N_18081,N_15740);
nor U21098 (N_21098,N_16610,N_15653);
and U21099 (N_21099,N_16107,N_15408);
xor U21100 (N_21100,N_17399,N_15952);
or U21101 (N_21101,N_18570,N_18877);
nor U21102 (N_21102,N_18989,N_18818);
and U21103 (N_21103,N_19257,N_18019);
xnor U21104 (N_21104,N_16483,N_17297);
xnor U21105 (N_21105,N_15719,N_16411);
nand U21106 (N_21106,N_18388,N_17485);
nand U21107 (N_21107,N_17272,N_16052);
or U21108 (N_21108,N_16722,N_19413);
and U21109 (N_21109,N_19900,N_19736);
and U21110 (N_21110,N_16693,N_16721);
nand U21111 (N_21111,N_15313,N_16613);
nand U21112 (N_21112,N_19755,N_16986);
nor U21113 (N_21113,N_17402,N_19721);
nor U21114 (N_21114,N_16487,N_15517);
xnor U21115 (N_21115,N_19840,N_17128);
and U21116 (N_21116,N_17098,N_17528);
and U21117 (N_21117,N_17537,N_19608);
xnor U21118 (N_21118,N_17438,N_18787);
nand U21119 (N_21119,N_16643,N_19891);
nand U21120 (N_21120,N_17839,N_17779);
and U21121 (N_21121,N_19844,N_19753);
or U21122 (N_21122,N_16930,N_18101);
nand U21123 (N_21123,N_19470,N_18575);
nor U21124 (N_21124,N_18451,N_17069);
nand U21125 (N_21125,N_17525,N_19072);
and U21126 (N_21126,N_17867,N_17343);
nand U21127 (N_21127,N_17627,N_19779);
or U21128 (N_21128,N_19927,N_19616);
and U21129 (N_21129,N_17440,N_17765);
nand U21130 (N_21130,N_18474,N_18984);
xnor U21131 (N_21131,N_19463,N_19687);
nand U21132 (N_21132,N_17655,N_18779);
xnor U21133 (N_21133,N_17704,N_15470);
and U21134 (N_21134,N_17500,N_15962);
nand U21135 (N_21135,N_19189,N_15146);
nand U21136 (N_21136,N_16979,N_16531);
and U21137 (N_21137,N_15302,N_18347);
nor U21138 (N_21138,N_19936,N_15187);
or U21139 (N_21139,N_18587,N_16261);
nand U21140 (N_21140,N_15732,N_18650);
or U21141 (N_21141,N_18130,N_18080);
nor U21142 (N_21142,N_16697,N_17345);
or U21143 (N_21143,N_19210,N_19253);
and U21144 (N_21144,N_19908,N_17332);
and U21145 (N_21145,N_18965,N_17473);
or U21146 (N_21146,N_18669,N_17233);
nor U21147 (N_21147,N_17301,N_16284);
or U21148 (N_21148,N_17353,N_15347);
or U21149 (N_21149,N_18325,N_17164);
or U21150 (N_21150,N_17804,N_15245);
xnor U21151 (N_21151,N_16945,N_18961);
nor U21152 (N_21152,N_18841,N_16128);
or U21153 (N_21153,N_15506,N_18593);
nor U21154 (N_21154,N_18752,N_19237);
nor U21155 (N_21155,N_18171,N_16022);
nand U21156 (N_21156,N_17596,N_15805);
xnor U21157 (N_21157,N_18972,N_18713);
xnor U21158 (N_21158,N_15234,N_17259);
and U21159 (N_21159,N_16081,N_18329);
nor U21160 (N_21160,N_16072,N_17919);
or U21161 (N_21161,N_16439,N_15829);
nand U21162 (N_21162,N_16966,N_15567);
xor U21163 (N_21163,N_18313,N_16137);
xnor U21164 (N_21164,N_15860,N_18874);
nand U21165 (N_21165,N_19974,N_18715);
nand U21166 (N_21166,N_19780,N_19363);
and U21167 (N_21167,N_15554,N_17605);
and U21168 (N_21168,N_18884,N_19594);
xnor U21169 (N_21169,N_15394,N_16051);
nand U21170 (N_21170,N_15072,N_18004);
nor U21171 (N_21171,N_18226,N_15369);
xor U21172 (N_21172,N_15142,N_19144);
nor U21173 (N_21173,N_19092,N_15638);
and U21174 (N_21174,N_18981,N_19050);
xor U21175 (N_21175,N_15867,N_15628);
nand U21176 (N_21176,N_16175,N_16273);
nor U21177 (N_21177,N_18441,N_15487);
and U21178 (N_21178,N_18209,N_15266);
xor U21179 (N_21179,N_17698,N_19711);
or U21180 (N_21180,N_16958,N_17006);
xor U21181 (N_21181,N_19084,N_16616);
nand U21182 (N_21182,N_16088,N_15033);
or U21183 (N_21183,N_18775,N_18339);
nand U21184 (N_21184,N_17530,N_16115);
nor U21185 (N_21185,N_18156,N_15694);
nor U21186 (N_21186,N_15937,N_17945);
and U21187 (N_21187,N_17354,N_19141);
and U21188 (N_21188,N_19040,N_17581);
nand U21189 (N_21189,N_15873,N_15881);
or U21190 (N_21190,N_15661,N_16048);
xor U21191 (N_21191,N_16111,N_19063);
nand U21192 (N_21192,N_15233,N_16931);
or U21193 (N_21193,N_17232,N_16761);
nor U21194 (N_21194,N_18283,N_18024);
and U21195 (N_21195,N_18730,N_17730);
nand U21196 (N_21196,N_16670,N_16038);
nor U21197 (N_21197,N_17751,N_17368);
or U21198 (N_21198,N_18639,N_15900);
nand U21199 (N_21199,N_19941,N_15230);
or U21200 (N_21200,N_15213,N_15403);
nand U21201 (N_21201,N_19701,N_15747);
xnor U21202 (N_21202,N_18139,N_16740);
and U21203 (N_21203,N_19054,N_18812);
nor U21204 (N_21204,N_16130,N_15919);
or U21205 (N_21205,N_16042,N_16239);
nor U21206 (N_21206,N_19673,N_18389);
or U21207 (N_21207,N_17273,N_15031);
xor U21208 (N_21208,N_15038,N_15414);
nor U21209 (N_21209,N_19080,N_17505);
nor U21210 (N_21210,N_15760,N_17326);
or U21211 (N_21211,N_19888,N_17305);
and U21212 (N_21212,N_17656,N_18538);
xor U21213 (N_21213,N_16484,N_16327);
nor U21214 (N_21214,N_15491,N_15623);
nor U21215 (N_21215,N_18125,N_19726);
xnor U21216 (N_21216,N_15941,N_18308);
or U21217 (N_21217,N_15428,N_19599);
nor U21218 (N_21218,N_16763,N_19142);
and U21219 (N_21219,N_17928,N_15014);
xor U21220 (N_21220,N_18190,N_15065);
nand U21221 (N_21221,N_19248,N_15726);
nand U21222 (N_21222,N_18088,N_19349);
nor U21223 (N_21223,N_18610,N_16686);
and U21224 (N_21224,N_15922,N_16481);
and U21225 (N_21225,N_17792,N_19860);
or U21226 (N_21226,N_16154,N_19930);
xnor U21227 (N_21227,N_18614,N_19075);
or U21228 (N_21228,N_18850,N_18096);
xnor U21229 (N_21229,N_17703,N_19872);
and U21230 (N_21230,N_18415,N_17274);
or U21231 (N_21231,N_17241,N_19833);
nand U21232 (N_21232,N_19112,N_17491);
nor U21233 (N_21233,N_15761,N_19973);
xnor U21234 (N_21234,N_19372,N_18229);
xor U21235 (N_21235,N_16710,N_18134);
or U21236 (N_21236,N_15869,N_15678);
nor U21237 (N_21237,N_16752,N_15318);
xnor U21238 (N_21238,N_16953,N_19731);
nor U21239 (N_21239,N_18048,N_18293);
nor U21240 (N_21240,N_19371,N_19220);
nand U21241 (N_21241,N_19331,N_19571);
and U21242 (N_21242,N_18055,N_18063);
or U21243 (N_21243,N_19907,N_16054);
and U21244 (N_21244,N_15629,N_19443);
nand U21245 (N_21245,N_17162,N_18676);
xnor U21246 (N_21246,N_16660,N_18414);
xnor U21247 (N_21247,N_18296,N_19274);
or U21248 (N_21248,N_16258,N_18268);
nand U21249 (N_21249,N_15185,N_19690);
or U21250 (N_21250,N_15112,N_17810);
xor U21251 (N_21251,N_16164,N_15870);
xor U21252 (N_21252,N_16596,N_17024);
nor U21253 (N_21253,N_16152,N_17481);
and U21254 (N_21254,N_19222,N_19539);
or U21255 (N_21255,N_19268,N_17228);
xnor U21256 (N_21256,N_16810,N_15236);
nor U21257 (N_21257,N_18700,N_18095);
or U21258 (N_21258,N_17286,N_15635);
or U21259 (N_21259,N_17338,N_18336);
nor U21260 (N_21260,N_18434,N_18317);
xnor U21261 (N_21261,N_19849,N_19154);
nand U21262 (N_21262,N_18996,N_17371);
and U21263 (N_21263,N_19502,N_16790);
xnor U21264 (N_21264,N_18122,N_16857);
nor U21265 (N_21265,N_15488,N_15009);
xor U21266 (N_21266,N_15053,N_17722);
nor U21267 (N_21267,N_15061,N_18303);
nor U21268 (N_21268,N_19225,N_18567);
and U21269 (N_21269,N_17889,N_15946);
xnor U21270 (N_21270,N_19479,N_17567);
or U21271 (N_21271,N_18753,N_15697);
nand U21272 (N_21272,N_15665,N_15405);
nand U21273 (N_21273,N_18684,N_18642);
and U21274 (N_21274,N_18704,N_15926);
or U21275 (N_21275,N_16677,N_18179);
and U21276 (N_21276,N_18643,N_16769);
xor U21277 (N_21277,N_15184,N_15569);
and U21278 (N_21278,N_16063,N_19472);
nor U21279 (N_21279,N_18918,N_18564);
nor U21280 (N_21280,N_16232,N_17882);
or U21281 (N_21281,N_19921,N_17496);
nand U21282 (N_21282,N_15401,N_19403);
xor U21283 (N_21283,N_19955,N_16242);
and U21284 (N_21284,N_15190,N_17645);
xor U21285 (N_21285,N_18390,N_15306);
or U21286 (N_21286,N_18688,N_18064);
or U21287 (N_21287,N_17885,N_16751);
and U21288 (N_21288,N_18504,N_18419);
and U21289 (N_21289,N_18275,N_18655);
and U21290 (N_21290,N_16910,N_17649);
and U21291 (N_21291,N_18299,N_18195);
nand U21292 (N_21292,N_18366,N_19740);
or U21293 (N_21293,N_15948,N_16865);
or U21294 (N_21294,N_15006,N_18750);
nand U21295 (N_21295,N_17127,N_17734);
nor U21296 (N_21296,N_19666,N_19645);
and U21297 (N_21297,N_19065,N_17754);
nand U21298 (N_21298,N_18804,N_19799);
xnor U21299 (N_21299,N_19806,N_16306);
or U21300 (N_21300,N_16617,N_16773);
nor U21301 (N_21301,N_17676,N_18073);
xnor U21302 (N_21302,N_17579,N_16990);
nand U21303 (N_21303,N_17612,N_19541);
and U21304 (N_21304,N_17921,N_19803);
xnor U21305 (N_21305,N_17819,N_17964);
and U21306 (N_21306,N_19158,N_16991);
nor U21307 (N_21307,N_17089,N_16090);
xnor U21308 (N_21308,N_15273,N_17942);
xnor U21309 (N_21309,N_19783,N_19358);
and U21310 (N_21310,N_19124,N_19382);
xor U21311 (N_21311,N_19928,N_15644);
nand U21312 (N_21312,N_18909,N_15363);
nand U21313 (N_21313,N_16625,N_15325);
or U21314 (N_21314,N_19827,N_16492);
and U21315 (N_21315,N_19778,N_16993);
xor U21316 (N_21316,N_17862,N_17178);
nor U21317 (N_21317,N_18270,N_15728);
or U21318 (N_21318,N_18912,N_18563);
or U21319 (N_21319,N_17744,N_18622);
nand U21320 (N_21320,N_15217,N_17455);
nand U21321 (N_21321,N_18151,N_15242);
nand U21322 (N_21322,N_18364,N_19563);
nand U21323 (N_21323,N_17173,N_17999);
and U21324 (N_21324,N_15377,N_18543);
xor U21325 (N_21325,N_19314,N_18240);
and U21326 (N_21326,N_16840,N_16003);
xor U21327 (N_21327,N_19689,N_17773);
nor U21328 (N_21328,N_18175,N_18871);
nor U21329 (N_21329,N_18127,N_16782);
nor U21330 (N_21330,N_15674,N_15951);
nor U21331 (N_21331,N_16068,N_16112);
nand U21332 (N_21332,N_17460,N_18741);
xor U21333 (N_21333,N_17743,N_19610);
or U21334 (N_21334,N_16495,N_19929);
or U21335 (N_21335,N_18126,N_19505);
or U21336 (N_21336,N_19436,N_17248);
xnor U21337 (N_21337,N_17076,N_18305);
xnor U21338 (N_21338,N_15118,N_19341);
nand U21339 (N_21339,N_15115,N_17944);
nand U21340 (N_21340,N_15059,N_19697);
nor U21341 (N_21341,N_15616,N_17870);
or U21342 (N_21342,N_18066,N_17479);
and U21343 (N_21343,N_17701,N_16664);
xnor U21344 (N_21344,N_18499,N_18014);
or U21345 (N_21345,N_17699,N_16560);
nand U21346 (N_21346,N_18358,N_18149);
nand U21347 (N_21347,N_16243,N_16174);
nand U21348 (N_21348,N_16725,N_15134);
xor U21349 (N_21349,N_16634,N_16349);
or U21350 (N_21350,N_16672,N_15155);
nand U21351 (N_21351,N_19017,N_18220);
or U21352 (N_21352,N_18821,N_15739);
and U21353 (N_21353,N_17214,N_16036);
or U21354 (N_21354,N_19893,N_18816);
or U21355 (N_21355,N_16402,N_17304);
nand U21356 (N_21356,N_16159,N_15160);
nor U21357 (N_21357,N_19547,N_19918);
nor U21358 (N_21358,N_15606,N_16104);
xnor U21359 (N_21359,N_19361,N_15420);
or U21360 (N_21360,N_15331,N_19631);
and U21361 (N_21361,N_15942,N_19477);
nand U21362 (N_21362,N_19931,N_16588);
xnor U21363 (N_21363,N_17911,N_18079);
xnor U21364 (N_21364,N_17629,N_16424);
nor U21365 (N_21365,N_16307,N_19419);
xnor U21366 (N_21366,N_15630,N_15988);
nand U21367 (N_21367,N_15333,N_18012);
xor U21368 (N_21368,N_17335,N_19626);
xor U21369 (N_21369,N_17401,N_19425);
or U21370 (N_21370,N_18222,N_19133);
and U21371 (N_21371,N_19263,N_17062);
nand U21372 (N_21372,N_16659,N_15677);
or U21373 (N_21373,N_16496,N_16849);
xor U21374 (N_21374,N_16161,N_15956);
and U21375 (N_21375,N_15913,N_15791);
or U21376 (N_21376,N_19603,N_17050);
or U21377 (N_21377,N_19752,N_19695);
nor U21378 (N_21378,N_16407,N_17041);
xnor U21379 (N_21379,N_18112,N_18784);
nor U21380 (N_21380,N_17574,N_19184);
nand U21381 (N_21381,N_15660,N_19708);
nand U21382 (N_21382,N_19975,N_16788);
or U21383 (N_21383,N_16817,N_15545);
nand U21384 (N_21384,N_17875,N_19030);
nand U21385 (N_21385,N_18559,N_16419);
or U21386 (N_21386,N_15526,N_15412);
nor U21387 (N_21387,N_18046,N_16181);
and U21388 (N_21388,N_15980,N_15541);
nor U21389 (N_21389,N_19554,N_19693);
nand U21390 (N_21390,N_19430,N_19538);
nand U21391 (N_21391,N_18590,N_15332);
nand U21392 (N_21392,N_15627,N_15621);
or U21393 (N_21393,N_18717,N_17200);
nand U21394 (N_21394,N_15798,N_15564);
nor U21395 (N_21395,N_15849,N_17916);
xnor U21396 (N_21396,N_16575,N_16624);
or U21397 (N_21397,N_16779,N_15817);
or U21398 (N_21398,N_15489,N_18274);
nand U21399 (N_21399,N_19194,N_16533);
and U21400 (N_21400,N_18635,N_18851);
nor U21401 (N_21401,N_17678,N_19223);
and U21402 (N_21402,N_17848,N_18826);
or U21403 (N_21403,N_15465,N_18603);
xor U21404 (N_21404,N_19271,N_16279);
nand U21405 (N_21405,N_18663,N_18747);
nand U21406 (N_21406,N_18853,N_19213);
nor U21407 (N_21407,N_15397,N_19656);
or U21408 (N_21408,N_16248,N_19750);
nand U21409 (N_21409,N_17518,N_16794);
or U21410 (N_21410,N_15483,N_17148);
nor U21411 (N_21411,N_15231,N_16786);
or U21412 (N_21412,N_16726,N_15186);
xor U21413 (N_21413,N_17422,N_16247);
nor U21414 (N_21414,N_19272,N_18935);
xnor U21415 (N_21415,N_19444,N_17953);
xor U21416 (N_21416,N_19999,N_19534);
nor U21417 (N_21417,N_15153,N_18473);
and U21418 (N_21418,N_16961,N_17262);
nor U21419 (N_21419,N_17532,N_18320);
or U21420 (N_21420,N_19582,N_19094);
xor U21421 (N_21421,N_19602,N_16949);
and U21422 (N_21422,N_19580,N_17914);
xor U21423 (N_21423,N_17474,N_16278);
nor U21424 (N_21424,N_15020,N_18666);
xnor U21425 (N_21425,N_17096,N_16335);
nand U21426 (N_21426,N_17712,N_19197);
nand U21427 (N_21427,N_16765,N_17458);
nor U21428 (N_21428,N_18269,N_15877);
or U21429 (N_21429,N_15291,N_19320);
nor U21430 (N_21430,N_15824,N_19397);
nor U21431 (N_21431,N_16756,N_19870);
nor U21432 (N_21432,N_17662,N_18097);
xnor U21433 (N_21433,N_15004,N_16783);
nand U21434 (N_21434,N_17383,N_18197);
and U21435 (N_21435,N_17105,N_17904);
nand U21436 (N_21436,N_15028,N_18076);
and U21437 (N_21437,N_18673,N_17313);
xnor U21438 (N_21438,N_16087,N_17950);
nor U21439 (N_21439,N_15676,N_15940);
or U21440 (N_21440,N_18861,N_15861);
nand U21441 (N_21441,N_19367,N_16908);
or U21442 (N_21442,N_18189,N_17437);
nand U21443 (N_21443,N_19718,N_18848);
nor U21444 (N_21444,N_16959,N_15154);
and U21445 (N_21445,N_15247,N_17803);
nor U21446 (N_21446,N_18428,N_16449);
or U21447 (N_21447,N_17969,N_16109);
and U21448 (N_21448,N_18191,N_19494);
xor U21449 (N_21449,N_18900,N_18009);
xor U21450 (N_21450,N_18835,N_17943);
nor U21451 (N_21451,N_15441,N_17917);
nand U21452 (N_21452,N_19486,N_17344);
or U21453 (N_21453,N_19129,N_18561);
or U21454 (N_21454,N_17795,N_17471);
nand U21455 (N_21455,N_17824,N_15267);
xnor U21456 (N_21456,N_18751,N_19774);
nor U21457 (N_21457,N_17578,N_18337);
xor U21458 (N_21458,N_15432,N_17508);
nor U21459 (N_21459,N_19245,N_17534);
or U21460 (N_21460,N_17841,N_16342);
xnor U21461 (N_21461,N_15858,N_18892);
or U21462 (N_21462,N_17330,N_15453);
nor U21463 (N_21463,N_16241,N_19857);
nor U21464 (N_21464,N_15589,N_17972);
nand U21465 (N_21465,N_16400,N_15478);
and U21466 (N_21466,N_15197,N_17488);
xor U21467 (N_21467,N_15225,N_18070);
and U21468 (N_21468,N_19389,N_15168);
xor U21469 (N_21469,N_18345,N_15274);
or U21470 (N_21470,N_17275,N_15532);
nand U21471 (N_21471,N_16057,N_15135);
nor U21472 (N_21472,N_17020,N_19933);
nor U21473 (N_21473,N_15551,N_18557);
nor U21474 (N_21474,N_15442,N_19265);
or U21475 (N_21475,N_15169,N_19856);
xor U21476 (N_21476,N_17145,N_18660);
xnor U21477 (N_21477,N_17880,N_19564);
or U21478 (N_21478,N_19842,N_15705);
xnor U21479 (N_21479,N_15034,N_17951);
nor U21480 (N_21480,N_19466,N_18605);
and U21481 (N_21481,N_18424,N_16636);
nor U21482 (N_21482,N_18889,N_17322);
or U21483 (N_21483,N_15584,N_16015);
and U21484 (N_21484,N_18492,N_17768);
nor U21485 (N_21485,N_18278,N_15141);
nor U21486 (N_21486,N_16320,N_17588);
or U21487 (N_21487,N_16619,N_17622);
nor U21488 (N_21488,N_18695,N_16212);
and U21489 (N_21489,N_19492,N_15044);
nor U21490 (N_21490,N_15847,N_18911);
nor U21491 (N_21491,N_15099,N_15853);
or U21492 (N_21492,N_17066,N_19905);
or U21493 (N_21493,N_16950,N_16915);
or U21494 (N_21494,N_18251,N_15315);
or U21495 (N_21495,N_17349,N_15979);
nand U21496 (N_21496,N_15471,N_15219);
or U21497 (N_21497,N_16364,N_15875);
nor U21498 (N_21498,N_17318,N_15406);
nand U21499 (N_21499,N_17132,N_17431);
or U21500 (N_21500,N_16142,N_16996);
or U21501 (N_21501,N_15529,N_16315);
nor U21502 (N_21502,N_19298,N_17307);
or U21503 (N_21503,N_16071,N_16493);
and U21504 (N_21504,N_19786,N_16951);
or U21505 (N_21505,N_15269,N_17884);
and U21506 (N_21506,N_19984,N_18985);
or U21507 (N_21507,N_17208,N_18475);
nor U21508 (N_21508,N_16781,N_16525);
or U21509 (N_21509,N_15799,N_15445);
nand U21510 (N_21510,N_16540,N_19214);
nand U21511 (N_21511,N_19858,N_17681);
nand U21512 (N_21512,N_16689,N_16023);
xnor U21513 (N_21513,N_17797,N_16975);
and U21514 (N_21514,N_17283,N_18887);
xor U21515 (N_21515,N_15484,N_17215);
or U21516 (N_21516,N_15516,N_17408);
xnor U21517 (N_21517,N_17709,N_19406);
xor U21518 (N_21518,N_16586,N_17789);
nor U21519 (N_21519,N_18847,N_16654);
nor U21520 (N_21520,N_18733,N_17406);
and U21521 (N_21521,N_18544,N_16696);
or U21522 (N_21522,N_16384,N_17637);
nor U21523 (N_21523,N_15690,N_19166);
or U21524 (N_21524,N_19483,N_18353);
or U21525 (N_21525,N_19454,N_16940);
nand U21526 (N_21526,N_15936,N_16240);
nand U21527 (N_21527,N_18113,N_18034);
nor U21528 (N_21528,N_15354,N_15056);
nand U21529 (N_21529,N_17060,N_19378);
or U21530 (N_21530,N_19525,N_15576);
nand U21531 (N_21531,N_16494,N_18378);
or U21532 (N_21532,N_16105,N_16465);
or U21533 (N_21533,N_16825,N_19276);
nand U21534 (N_21534,N_19344,N_16538);
nand U21535 (N_21535,N_17419,N_15794);
nor U21536 (N_21536,N_17224,N_15205);
or U21537 (N_21537,N_15648,N_16653);
or U21538 (N_21538,N_15077,N_19067);
or U21539 (N_21539,N_17718,N_17755);
or U21540 (N_21540,N_16032,N_18594);
or U21541 (N_21541,N_17613,N_15037);
or U21542 (N_21542,N_16119,N_15976);
nand U21543 (N_21543,N_18410,N_15447);
xor U21544 (N_21544,N_18799,N_19330);
or U21545 (N_21545,N_18581,N_18616);
or U21546 (N_21546,N_19435,N_17339);
or U21547 (N_21547,N_16084,N_18027);
nand U21548 (N_21548,N_18111,N_19713);
or U21549 (N_21549,N_18674,N_15067);
and U21550 (N_21550,N_17443,N_16598);
or U21551 (N_21551,N_19130,N_17210);
nand U21552 (N_21552,N_19193,N_16290);
nor U21553 (N_21553,N_17685,N_16720);
nand U21554 (N_21554,N_18982,N_16435);
nor U21555 (N_21555,N_16709,N_17446);
nor U21556 (N_21556,N_16552,N_18049);
xnor U21557 (N_21557,N_18797,N_16899);
nand U21558 (N_21558,N_15064,N_17669);
xnor U21559 (N_21559,N_16452,N_16561);
nand U21560 (N_21560,N_19705,N_16343);
nand U21561 (N_21561,N_18906,N_15209);
nand U21562 (N_21562,N_18637,N_17199);
nand U21563 (N_21563,N_15294,N_18208);
or U21564 (N_21564,N_19422,N_15275);
or U21565 (N_21565,N_17568,N_15323);
or U21566 (N_21566,N_18479,N_15673);
nor U21567 (N_21567,N_16621,N_18566);
nor U21568 (N_21568,N_18609,N_18272);
xnor U21569 (N_21569,N_18232,N_16994);
xor U21570 (N_21570,N_18568,N_15240);
or U21571 (N_21571,N_18736,N_15710);
nand U21572 (N_21572,N_19146,N_18651);
or U21573 (N_21573,N_17403,N_16896);
and U21574 (N_21574,N_18188,N_19495);
and U21575 (N_21575,N_15811,N_15321);
nor U21576 (N_21576,N_16412,N_16431);
nor U21577 (N_21577,N_19177,N_19024);
and U21578 (N_21578,N_18261,N_17179);
xor U21579 (N_21579,N_19912,N_15656);
nand U21580 (N_21580,N_17872,N_15198);
or U21581 (N_21581,N_19417,N_17369);
nor U21582 (N_21582,N_19231,N_15350);
nor U21583 (N_21583,N_17686,N_17587);
nor U21584 (N_21584,N_15433,N_17032);
nor U21585 (N_21585,N_16612,N_19157);
and U21586 (N_21586,N_15425,N_18407);
nor U21587 (N_21587,N_18203,N_18395);
nor U21588 (N_21588,N_17646,N_16473);
or U21589 (N_21589,N_17851,N_18193);
or U21590 (N_21590,N_19044,N_17616);
nand U21591 (N_21591,N_15611,N_15961);
nor U21592 (N_21592,N_15508,N_16527);
nand U21593 (N_21593,N_18075,N_18880);
nand U21594 (N_21594,N_15781,N_16074);
xor U21595 (N_21595,N_15994,N_18958);
and U21596 (N_21596,N_19475,N_18795);
nor U21597 (N_21597,N_17957,N_18954);
nor U21598 (N_21598,N_17799,N_17815);
or U21599 (N_21599,N_18595,N_17526);
xnor U21600 (N_21600,N_16075,N_18815);
xnor U21601 (N_21601,N_16379,N_19859);
xor U21602 (N_21602,N_17770,N_19601);
nand U21603 (N_21603,N_16638,N_16237);
or U21604 (N_21604,N_17931,N_18435);
and U21605 (N_21605,N_16498,N_18010);
nor U21606 (N_21606,N_15613,N_17721);
and U21607 (N_21607,N_15851,N_18486);
nand U21608 (N_21608,N_15822,N_17648);
and U21609 (N_21609,N_16149,N_17996);
xor U21610 (N_21610,N_18995,N_18058);
xnor U21611 (N_21611,N_16162,N_17373);
xnor U21612 (N_21612,N_15329,N_16360);
nand U21613 (N_21613,N_15542,N_19847);
or U21614 (N_21614,N_16194,N_16553);
nand U21615 (N_21615,N_16226,N_19224);
and U21616 (N_21616,N_19310,N_15724);
or U21617 (N_21617,N_15222,N_18411);
nor U21618 (N_21618,N_18574,N_15814);
or U21619 (N_21619,N_15229,N_16518);
or U21620 (N_21620,N_16330,N_16984);
nor U21621 (N_21621,N_19256,N_17561);
xnor U21622 (N_21622,N_16189,N_15353);
or U21623 (N_21623,N_19634,N_15522);
xor U21624 (N_21624,N_18558,N_17480);
xor U21625 (N_21625,N_15000,N_18551);
xnor U21626 (N_21626,N_18408,N_18846);
and U21627 (N_21627,N_17805,N_19204);
nand U21628 (N_21628,N_15342,N_17022);
and U21629 (N_21629,N_18692,N_16558);
or U21630 (N_21630,N_15527,N_15810);
and U21631 (N_21631,N_17511,N_18106);
and U21632 (N_21632,N_19388,N_16826);
and U21633 (N_21633,N_16519,N_16888);
nor U21634 (N_21634,N_18252,N_16583);
and U21635 (N_21635,N_19234,N_15075);
nand U21636 (N_21636,N_19757,N_18331);
nor U21637 (N_21637,N_17930,N_18693);
nand U21638 (N_21638,N_17506,N_18307);
and U21639 (N_21639,N_19312,N_18053);
or U21640 (N_21640,N_19297,N_18690);
xor U21641 (N_21641,N_17873,N_18258);
and U21642 (N_21642,N_17342,N_15573);
xor U21643 (N_21643,N_17111,N_18712);
xnor U21644 (N_21644,N_18778,N_15943);
nor U21645 (N_21645,N_15819,N_19749);
or U21646 (N_21646,N_18146,N_19623);
and U21647 (N_21647,N_18601,N_15216);
nor U21648 (N_21648,N_15058,N_19810);
nor U21649 (N_21649,N_19961,N_19958);
nor U21650 (N_21650,N_17504,N_18845);
or U21651 (N_21651,N_17239,N_18089);
or U21652 (N_21652,N_16673,N_16724);
and U21653 (N_21653,N_19990,N_15789);
xor U21654 (N_21654,N_15149,N_19614);
xor U21655 (N_21655,N_15462,N_15327);
nor U21656 (N_21656,N_17502,N_16317);
nand U21657 (N_21657,N_19326,N_19710);
or U21658 (N_21658,N_18044,N_16549);
or U21659 (N_21659,N_18671,N_18469);
xor U21660 (N_21660,N_18381,N_15494);
nand U21661 (N_21661,N_16389,N_19200);
and U21662 (N_21662,N_15735,N_16430);
xnor U21663 (N_21663,N_18975,N_17366);
and U21664 (N_21664,N_18652,N_19932);
nand U21665 (N_21665,N_18124,N_17040);
nand U21666 (N_21666,N_16772,N_18281);
and U21667 (N_21667,N_15874,N_17355);
nand U21668 (N_21668,N_17929,N_17136);
nor U21669 (N_21669,N_16626,N_17255);
or U21670 (N_21670,N_17939,N_19764);
or U21671 (N_21671,N_17982,N_17842);
or U21672 (N_21672,N_17909,N_15560);
or U21673 (N_21673,N_19825,N_19383);
nor U21674 (N_21674,N_16534,N_16938);
nor U21675 (N_21675,N_17666,N_19788);
and U21676 (N_21676,N_17139,N_18100);
xnor U21677 (N_21677,N_19926,N_18460);
nor U21678 (N_21678,N_15954,N_19762);
xnor U21679 (N_21679,N_17409,N_17299);
xor U21680 (N_21680,N_18227,N_17762);
nor U21681 (N_21681,N_19567,N_18672);
xnor U21682 (N_21682,N_16326,N_16426);
or U21683 (N_21683,N_19066,N_17694);
and U21684 (N_21684,N_18723,N_16388);
xnor U21685 (N_21685,N_15960,N_16862);
or U21686 (N_21686,N_17966,N_15930);
or U21687 (N_21687,N_17149,N_15769);
nor U21688 (N_21688,N_18160,N_19308);
xor U21689 (N_21689,N_15023,N_17555);
and U21690 (N_21690,N_18198,N_17180);
xor U21691 (N_21691,N_15012,N_19176);
nand U21692 (N_21692,N_15891,N_15512);
nand U21693 (N_21693,N_17486,N_18057);
xnor U21694 (N_21694,N_18838,N_15599);
and U21695 (N_21695,N_19455,N_19487);
xor U21696 (N_21696,N_18789,N_16139);
nand U21697 (N_21697,N_19892,N_17292);
and U21698 (N_21698,N_15550,N_16728);
nand U21699 (N_21699,N_18330,N_16079);
and U21700 (N_21700,N_15856,N_15570);
nor U21701 (N_21701,N_17094,N_16067);
or U21702 (N_21702,N_18774,N_18725);
nor U21703 (N_21703,N_15137,N_16291);
nor U21704 (N_21704,N_17010,N_15421);
nand U21705 (N_21705,N_19638,N_18748);
and U21706 (N_21706,N_16745,N_15235);
or U21707 (N_21707,N_16089,N_15374);
or U21708 (N_21708,N_15650,N_19052);
or U21709 (N_21709,N_16371,N_17609);
and U21710 (N_21710,N_19402,N_18458);
and U21711 (N_21711,N_15767,N_15170);
or U21712 (N_21712,N_18260,N_15770);
nand U21713 (N_21713,N_17932,N_16093);
xnor U21714 (N_21714,N_19972,N_16332);
nand U21715 (N_21715,N_16314,N_15622);
and U21716 (N_21716,N_15017,N_19993);
or U21717 (N_21717,N_15546,N_15304);
nand U21718 (N_21718,N_17104,N_17849);
xor U21719 (N_21719,N_18646,N_16440);
or U21720 (N_21720,N_15982,N_18115);
and U21721 (N_21721,N_17254,N_19131);
xor U21722 (N_21722,N_18497,N_15679);
nand U21723 (N_21723,N_17346,N_16004);
and U21724 (N_21724,N_19357,N_15449);
or U21725 (N_21725,N_19060,N_15404);
and U21726 (N_21726,N_15348,N_18960);
nor U21727 (N_21727,N_17927,N_19947);
or U21728 (N_21728,N_18256,N_15263);
or U21729 (N_21729,N_18754,N_15708);
and U21730 (N_21730,N_19049,N_18964);
and U21731 (N_21731,N_19681,N_17860);
nor U21732 (N_21732,N_17714,N_18967);
nand U21733 (N_21733,N_17891,N_15604);
nand U21734 (N_21734,N_16296,N_17535);
and U21735 (N_21735,N_15707,N_16675);
nor U21736 (N_21736,N_17855,N_15953);
or U21737 (N_21737,N_16177,N_19347);
and U21738 (N_21738,N_19457,N_19867);
xor U21739 (N_21739,N_16236,N_15392);
or U21740 (N_21740,N_15510,N_18456);
nand U21741 (N_21741,N_18873,N_17390);
nand U21742 (N_21742,N_18980,N_15356);
or U21743 (N_21743,N_17618,N_18155);
and U21744 (N_21744,N_15974,N_17079);
nor U21745 (N_21745,N_16260,N_19683);
and U21746 (N_21746,N_16608,N_18745);
and U21747 (N_21747,N_19519,N_18920);
nand U21748 (N_21748,N_19442,N_15698);
and U21749 (N_21749,N_15132,N_17151);
nor U21750 (N_21750,N_16789,N_15790);
and U21751 (N_21751,N_16639,N_19014);
or U21752 (N_21752,N_19820,N_16622);
or U21753 (N_21753,N_16515,N_17204);
nor U21754 (N_21754,N_18054,N_19009);
xnor U21755 (N_21755,N_16573,N_17520);
or U21756 (N_21756,N_17152,N_16340);
nor U21757 (N_21757,N_15241,N_15102);
or U21758 (N_21758,N_15024,N_15983);
nand U21759 (N_21759,N_17249,N_16157);
xnor U21760 (N_21760,N_17746,N_17828);
and U21761 (N_21761,N_17120,N_18291);
nand U21762 (N_21762,N_19831,N_19537);
xnor U21763 (N_21763,N_17639,N_17052);
xnor U21764 (N_21764,N_16445,N_17191);
or U21765 (N_21765,N_19772,N_16861);
nand U21766 (N_21766,N_17886,N_17464);
nand U21767 (N_21767,N_16245,N_17563);
or U21768 (N_21768,N_15981,N_15607);
and U21769 (N_21769,N_17767,N_15175);
nand U21770 (N_21770,N_17572,N_17134);
nor U21771 (N_21771,N_19399,N_18755);
nand U21772 (N_21772,N_19026,N_17607);
and U21773 (N_21773,N_17570,N_18685);
or U21774 (N_21774,N_15972,N_16521);
or U21775 (N_21775,N_18026,N_15182);
and U21776 (N_21776,N_15123,N_18350);
xnor U21777 (N_21777,N_18116,N_17049);
xnor U21778 (N_21778,N_16871,N_17077);
nand U21779 (N_21779,N_19292,N_15910);
xor U21780 (N_21780,N_15259,N_19942);
and U21781 (N_21781,N_19481,N_17546);
nand U21782 (N_21782,N_15583,N_17632);
nand U21783 (N_21783,N_19091,N_19730);
or U21784 (N_21784,N_19570,N_18565);
nor U21785 (N_21785,N_16916,N_19207);
nor U21786 (N_21786,N_18518,N_17268);
nand U21787 (N_21787,N_18131,N_15848);
or U21788 (N_21788,N_19561,N_15035);
nand U21789 (N_21789,N_15296,N_17106);
and U21790 (N_21790,N_16489,N_18300);
xnor U21791 (N_21791,N_15498,N_18783);
and U21792 (N_21792,N_16511,N_18266);
nor U21793 (N_21793,N_17117,N_19940);
nor U21794 (N_21794,N_18185,N_18466);
or U21795 (N_21795,N_19173,N_18925);
nor U21796 (N_21796,N_19469,N_16478);
xnor U21797 (N_21797,N_15774,N_18238);
nor U21798 (N_21798,N_16822,N_18689);
and U21799 (N_21799,N_18843,N_17515);
nor U21800 (N_21800,N_19916,N_15098);
and U21801 (N_21801,N_16099,N_18938);
and U21802 (N_21802,N_17113,N_17585);
and U21803 (N_21803,N_17793,N_15365);
or U21804 (N_21804,N_19775,N_16150);
and U21805 (N_21805,N_17559,N_18483);
nor U21806 (N_21806,N_17412,N_18681);
nor U21807 (N_21807,N_15130,N_15795);
or U21808 (N_21808,N_18413,N_19732);
and U21809 (N_21809,N_15129,N_16272);
or U21810 (N_21810,N_18145,N_15504);
xor U21811 (N_21811,N_16151,N_19001);
or U21812 (N_21812,N_17949,N_15645);
or U21813 (N_21813,N_16378,N_16936);
or U21814 (N_21814,N_16880,N_19818);
or U21815 (N_21815,N_16812,N_17510);
and U21816 (N_21816,N_19863,N_18582);
nand U21817 (N_21817,N_18348,N_16514);
or U21818 (N_21818,N_18484,N_15600);
nor U21819 (N_21819,N_19303,N_16750);
or U21820 (N_21820,N_17226,N_16744);
and U21821 (N_21821,N_15825,N_15008);
xor U21822 (N_21822,N_16266,N_16383);
and U21823 (N_21823,N_18206,N_19396);
nand U21824 (N_21824,N_17444,N_18052);
nand U21825 (N_21825,N_16895,N_15773);
or U21826 (N_21826,N_17589,N_16620);
or U21827 (N_21827,N_19748,N_16205);
xnor U21828 (N_21828,N_19390,N_15344);
and U21829 (N_21829,N_17059,N_15086);
xnor U21830 (N_21830,N_19514,N_17099);
nand U21831 (N_21831,N_18943,N_19553);
xor U21832 (N_21832,N_17461,N_19172);
nor U21833 (N_21833,N_19022,N_17462);
xor U21834 (N_21834,N_17794,N_17122);
nor U21835 (N_21835,N_18201,N_19852);
xnor U21836 (N_21836,N_19607,N_15830);
or U21837 (N_21837,N_15415,N_17417);
xor U21838 (N_21838,N_18169,N_15292);
and U21839 (N_21839,N_19181,N_16853);
and U21840 (N_21840,N_17808,N_15289);
nand U21841 (N_21841,N_18476,N_17284);
or U21842 (N_21842,N_17826,N_19549);
or U21843 (N_21843,N_15893,N_16637);
nand U21844 (N_21844,N_19746,N_17671);
or U21845 (N_21845,N_18282,N_17257);
nor U21846 (N_21846,N_16648,N_19832);
or U21847 (N_21847,N_17710,N_19745);
nand U21848 (N_21848,N_19340,N_16503);
or U21849 (N_21849,N_15336,N_18400);
nor U21850 (N_21850,N_15966,N_15927);
or U21851 (N_21851,N_15283,N_15816);
and U21852 (N_21852,N_16881,N_18930);
xnor U21853 (N_21853,N_16544,N_19235);
nand U21854 (N_21854,N_19848,N_16683);
and U21855 (N_21855,N_16732,N_17597);
and U21856 (N_21856,N_18453,N_15119);
and U21857 (N_21857,N_18327,N_16217);
and U21858 (N_21858,N_19068,N_15370);
nand U21859 (N_21859,N_16270,N_16385);
nor U21860 (N_21860,N_18560,N_18627);
nor U21861 (N_21861,N_17874,N_17997);
nand U21862 (N_21862,N_15597,N_19586);
or U21863 (N_21863,N_16453,N_18542);
nand U21864 (N_21864,N_18398,N_19510);
nand U21865 (N_21865,N_19169,N_18630);
nor U21866 (N_21866,N_16479,N_16801);
xor U21867 (N_21867,N_17700,N_18516);
xor U21868 (N_21868,N_16197,N_15590);
and U21869 (N_21869,N_18806,N_16691);
and U21870 (N_21870,N_16846,N_19452);
xnor U21871 (N_21871,N_18791,N_17663);
or U21872 (N_21872,N_16480,N_16319);
xor U21873 (N_21873,N_16434,N_18969);
and U21874 (N_21874,N_17002,N_17861);
nand U21875 (N_21875,N_15925,N_19684);
xnor U21876 (N_21876,N_15571,N_16209);
xor U21877 (N_21877,N_18555,N_19897);
and U21878 (N_21878,N_19738,N_15905);
and U21879 (N_21879,N_17141,N_19101);
or U21880 (N_21880,N_16843,N_19392);
or U21881 (N_21881,N_19139,N_16191);
and U21882 (N_21882,N_17261,N_17362);
and U21883 (N_21883,N_15776,N_16210);
nor U21884 (N_21884,N_17984,N_16998);
and U21885 (N_21885,N_16345,N_15243);
xor U21886 (N_21886,N_16680,N_19935);
nor U21887 (N_21887,N_15480,N_16298);
xor U21888 (N_21888,N_16969,N_19734);
nand U21889 (N_21889,N_18047,N_18513);
and U21890 (N_21890,N_19243,N_16103);
xnor U21891 (N_21891,N_17711,N_15423);
or U21892 (N_21892,N_17554,N_19359);
nor U21893 (N_21893,N_17749,N_17633);
xor U21894 (N_21894,N_16442,N_17097);
xnor U21895 (N_21895,N_16447,N_17490);
nand U21896 (N_21896,N_18426,N_16623);
xnor U21897 (N_21897,N_18333,N_18852);
nor U21898 (N_21898,N_16879,N_19878);
nor U21899 (N_21899,N_19471,N_17340);
xnor U21900 (N_21900,N_18792,N_15183);
nand U21901 (N_21901,N_15328,N_19316);
and U21902 (N_21902,N_15681,N_18031);
xor U21903 (N_21903,N_16376,N_19409);
xor U21904 (N_21904,N_16173,N_16733);
or U21905 (N_21905,N_18721,N_19529);
and U21906 (N_21906,N_19696,N_18162);
xnor U21907 (N_21907,N_19773,N_19114);
and U21908 (N_21908,N_17067,N_16444);
and U21909 (N_21909,N_18141,N_17667);
nand U21910 (N_21910,N_16854,N_16973);
xor U21911 (N_21911,N_18976,N_15632);
nand U21912 (N_21912,N_19518,N_18539);
nor U21913 (N_21913,N_15145,N_18762);
and U21914 (N_21914,N_15854,N_19700);
or U21915 (N_21915,N_17278,N_15696);
or U21916 (N_21916,N_18828,N_18668);
nand U21917 (N_21917,N_16358,N_18271);
nor U21918 (N_21918,N_17772,N_18257);
nand U21919 (N_21919,N_15308,N_17116);
xor U21920 (N_21920,N_16629,N_15659);
or U21921 (N_21921,N_17163,N_16963);
or U21922 (N_21922,N_19351,N_16187);
xor U21923 (N_21923,N_15838,N_15114);
nor U21924 (N_21924,N_19592,N_16196);
or U21925 (N_21925,N_16727,N_16117);
xnor U21926 (N_21926,N_15535,N_19016);
nand U21927 (N_21927,N_18304,N_18963);
nor U21928 (N_21928,N_18255,N_15467);
and U21929 (N_21929,N_17400,N_16918);
nor U21930 (N_21930,N_16386,N_16708);
nand U21931 (N_21931,N_16455,N_19866);
and U21932 (N_21932,N_17682,N_17745);
nor U21933 (N_21933,N_18467,N_17533);
or U21934 (N_21934,N_17571,N_18535);
nand U21935 (N_21935,N_16800,N_15171);
xor U21936 (N_21936,N_18033,N_18947);
and U21937 (N_21937,N_18488,N_15827);
nor U21938 (N_21938,N_19228,N_19401);
nand U21939 (N_21939,N_19229,N_17347);
or U21940 (N_21940,N_19771,N_16203);
nand U21941 (N_21941,N_15027,N_16061);
nor U21942 (N_21942,N_15702,N_15555);
or U21943 (N_21943,N_17081,N_17316);
or U21944 (N_21944,N_17222,N_17080);
nor U21945 (N_21945,N_16179,N_19288);
nand U21946 (N_21946,N_17150,N_16183);
and U21947 (N_21947,N_19986,N_15437);
nand U21948 (N_21948,N_16551,N_15413);
nand U21949 (N_21949,N_19924,N_16469);
and U21950 (N_21950,N_15366,N_19938);
nor U21951 (N_21951,N_16976,N_16110);
or U21952 (N_21952,N_15011,N_17445);
or U21953 (N_21953,N_18957,N_19354);
nand U21954 (N_21954,N_17295,N_18979);
or U21955 (N_21955,N_17905,N_17415);
or U21956 (N_21956,N_17834,N_19031);
or U21957 (N_21957,N_19489,N_19520);
nand U21958 (N_21958,N_18302,N_18525);
or U21959 (N_21959,N_18800,N_19574);
and U21960 (N_21960,N_16889,N_18184);
or U21961 (N_21961,N_16837,N_16234);
nand U21962 (N_21962,N_18110,N_18719);
nor U21963 (N_21963,N_16155,N_19032);
nand U21964 (N_21964,N_16185,N_19568);
nand U21965 (N_21965,N_15898,N_15434);
or U21966 (N_21966,N_19841,N_15257);
or U21967 (N_21967,N_15715,N_19819);
nor U21968 (N_21968,N_18218,N_19398);
nor U21969 (N_21969,N_16556,N_16599);
nand U21970 (N_21970,N_15298,N_16606);
nand U21971 (N_21971,N_17308,N_18342);
and U21972 (N_21972,N_15755,N_17519);
or U21973 (N_21973,N_17290,N_15812);
or U21974 (N_21974,N_18726,N_19431);
xor U21975 (N_21975,N_16344,N_15883);
nor U21976 (N_21976,N_16002,N_16377);
and U21977 (N_21977,N_18645,N_19737);
and U21978 (N_21978,N_17781,N_19839);
nand U21979 (N_21979,N_16227,N_18661);
and U21980 (N_21980,N_16369,N_15372);
and U21981 (N_21981,N_18082,N_18742);
xor U21982 (N_21982,N_18236,N_18955);
and U21983 (N_21983,N_17766,N_15844);
or U21984 (N_21984,N_18724,N_18446);
or U21985 (N_21985,N_18118,N_18355);
and U21986 (N_21986,N_15093,N_19609);
or U21987 (N_21987,N_15080,N_19611);
and U21988 (N_21988,N_15150,N_18917);
and U21989 (N_21989,N_17543,N_15156);
and U21990 (N_21990,N_19679,N_15460);
nor U21991 (N_21991,N_16337,N_17396);
or U21992 (N_21992,N_19085,N_15663);
or U21993 (N_21993,N_17788,N_15686);
and U21994 (N_21994,N_18007,N_19987);
xor U21995 (N_21995,N_16819,N_18856);
or U21996 (N_21996,N_19127,N_18615);
nor U21997 (N_21997,N_18662,N_15605);
nand U21998 (N_21998,N_18522,N_16218);
and U21999 (N_21999,N_18136,N_15375);
and U22000 (N_22000,N_18153,N_18524);
or U22001 (N_22001,N_18421,N_15879);
xnor U22002 (N_22002,N_17823,N_16267);
nand U22003 (N_22003,N_18527,N_15087);
xnor U22004 (N_22004,N_18589,N_16799);
nor U22005 (N_22005,N_18794,N_17319);
nor U22006 (N_22006,N_19221,N_16287);
nor U22007 (N_22007,N_19152,N_17790);
or U22008 (N_22008,N_19589,N_16118);
xnor U22009 (N_22009,N_16885,N_16456);
xor U22010 (N_22010,N_15640,N_16814);
and U22011 (N_22011,N_16501,N_18978);
or U22012 (N_22012,N_16166,N_15105);
and U22013 (N_22013,N_16510,N_15672);
nor U22014 (N_22014,N_17091,N_19781);
xor U22015 (N_22015,N_17407,N_16989);
or U22016 (N_22016,N_17439,N_16100);
xnor U22017 (N_22017,N_18436,N_16944);
xor U22018 (N_22018,N_15636,N_19754);
or U22019 (N_22019,N_15440,N_15841);
nor U22020 (N_22020,N_15270,N_15262);
nor U22021 (N_22021,N_15928,N_16595);
and U22022 (N_22022,N_17317,N_16014);
and U22023 (N_22023,N_17045,N_17382);
xor U22024 (N_22024,N_15902,N_16870);
xor U22025 (N_22025,N_19490,N_18945);
nor U22026 (N_22026,N_18739,N_15094);
nor U22027 (N_22027,N_15165,N_17817);
nand U22028 (N_22028,N_18941,N_19600);
nand U22029 (N_22029,N_19039,N_17312);
or U22030 (N_22030,N_18968,N_18312);
nand U22031 (N_22031,N_15788,N_17138);
nor U22032 (N_22032,N_16839,N_15523);
nor U22033 (N_22033,N_18485,N_15246);
xnor U22034 (N_22034,N_19756,N_16350);
and U22035 (N_22035,N_18078,N_19678);
or U22036 (N_22036,N_16914,N_19165);
nor U22037 (N_22037,N_17907,N_19598);
nand U22038 (N_22038,N_16845,N_15619);
or U22039 (N_22039,N_17840,N_15228);
or U22040 (N_22040,N_15720,N_15561);
xnor U22041 (N_22041,N_17812,N_17252);
nor U22042 (N_22042,N_17411,N_19944);
and U22043 (N_22043,N_19191,N_15032);
and U22044 (N_22044,N_15041,N_15855);
and U22045 (N_22045,N_17998,N_15594);
or U22046 (N_22046,N_18035,N_19995);
or U22047 (N_22047,N_16526,N_18654);
or U22048 (N_22048,N_15280,N_16065);
xor U22049 (N_22049,N_15581,N_19445);
nor U22050 (N_22050,N_18157,N_18951);
nand U22051 (N_22051,N_16662,N_19792);
xor U22052 (N_22052,N_17675,N_16450);
nand U22053 (N_22053,N_19896,N_19760);
nand U22054 (N_22054,N_16863,N_18051);
or U22055 (N_22055,N_19106,N_18953);
nand U22056 (N_22056,N_17075,N_18523);
xor U22057 (N_22057,N_18621,N_18418);
or U22058 (N_22058,N_15378,N_16900);
nor U22059 (N_22059,N_17761,N_19501);
nor U22060 (N_22060,N_16289,N_19982);
xor U22061 (N_22061,N_19714,N_19387);
xor U22062 (N_22062,N_18439,N_17230);
or U22063 (N_22063,N_16716,N_17832);
or U22064 (N_22064,N_17786,N_19280);
nor U22065 (N_22065,N_19675,N_16311);
or U22066 (N_22066,N_18319,N_16028);
or U22067 (N_22067,N_15253,N_19521);
nand U22068 (N_22068,N_15685,N_17293);
nor U22069 (N_22069,N_17869,N_15417);
or U22070 (N_22070,N_17850,N_16922);
or U22071 (N_22071,N_16420,N_18427);
or U22072 (N_22072,N_19302,N_18534);
or U22073 (N_22073,N_15446,N_17680);
and U22074 (N_22074,N_15060,N_19751);
and U22075 (N_22075,N_15852,N_16886);
nand U22076 (N_22076,N_16911,N_17245);
nor U22077 (N_22077,N_18519,N_15520);
nor U22078 (N_22078,N_19824,N_17497);
nand U22079 (N_22079,N_16050,N_19702);
xor U22080 (N_22080,N_16875,N_15422);
or U22081 (N_22081,N_18098,N_18463);
and U22082 (N_22082,N_16207,N_16791);
or U22083 (N_22083,N_19005,N_16651);
nor U22084 (N_22084,N_19830,N_18803);
nand U22085 (N_22085,N_18946,N_18950);
xnor U22086 (N_22086,N_19380,N_15108);
and U22087 (N_22087,N_15481,N_18763);
and U22088 (N_22088,N_16268,N_16262);
nand U22089 (N_22089,N_15221,N_16193);
nand U22090 (N_22090,N_16611,N_16894);
nor U22091 (N_22091,N_18782,N_19913);
nand U22092 (N_22092,N_18728,N_16382);
xnor U22093 (N_22093,N_15464,N_19281);
nor U22094 (N_22094,N_16034,N_17693);
nor U22095 (N_22095,N_16113,N_17043);
nand U22096 (N_22096,N_19386,N_19500);
nor U22097 (N_22097,N_18888,N_16302);
xor U22098 (N_22098,N_17920,N_19309);
nand U22099 (N_22099,N_19902,N_17696);
nor U22100 (N_22100,N_16890,N_19000);
or U22101 (N_22101,N_16277,N_16509);
or U22102 (N_22102,N_16792,N_15996);
xor U22103 (N_22103,N_17636,N_16131);
nand U22104 (N_22104,N_16749,N_17687);
nand U22105 (N_22105,N_16679,N_17311);
and U22106 (N_22106,N_18764,N_19815);
xor U22107 (N_22107,N_16942,N_15531);
and U22108 (N_22108,N_15389,N_15912);
and U22109 (N_22109,N_19817,N_19007);
nor U22110 (N_22110,N_15864,N_19071);
and U22111 (N_22111,N_18142,N_19655);
and U22112 (N_22112,N_15122,N_18301);
nand U22113 (N_22113,N_15055,N_17027);
or U22114 (N_22114,N_15574,N_17276);
xnor U22115 (N_22115,N_16999,N_16640);
nor U22116 (N_22116,N_19096,N_18588);
xnor U22117 (N_22117,N_16231,N_17985);
or U22118 (N_22118,N_16753,N_18253);
or U22119 (N_22119,N_19125,N_19925);
nor U22120 (N_22120,N_19020,N_15821);
nor U22121 (N_22121,N_16221,N_19418);
and U22122 (N_22122,N_19801,N_19335);
or U22123 (N_22123,N_16974,N_17023);
nand U22124 (N_22124,N_18859,N_16309);
nor U22125 (N_22125,N_15592,N_18514);
xnor U22126 (N_22126,N_19011,N_19262);
or U22127 (N_22127,N_19950,N_15418);
and U22128 (N_22128,N_19621,N_19458);
nand U22129 (N_22129,N_19295,N_19478);
and U22130 (N_22130,N_19759,N_17595);
and U22131 (N_22131,N_17617,N_17242);
nor U22132 (N_22132,N_15454,N_16171);
nand U22133 (N_22133,N_18137,N_16741);
nand U22134 (N_22134,N_16432,N_17124);
nand U22135 (N_22135,N_16120,N_19482);
and U22136 (N_22136,N_19002,N_15125);
xnor U22137 (N_22137,N_18893,N_16288);
nand U22138 (N_22138,N_16571,N_15646);
xnor U22139 (N_22139,N_19540,N_17994);
xor U22140 (N_22140,N_17670,N_16380);
xor U22141 (N_22141,N_15585,N_16133);
nand U22142 (N_22142,N_19433,N_18224);
and U22143 (N_22143,N_17573,N_19321);
and U22144 (N_22144,N_17182,N_15802);
nand U22145 (N_22145,N_15723,N_18633);
xor U22146 (N_22146,N_15586,N_19637);
or U22147 (N_22147,N_19282,N_15999);
and U22148 (N_22148,N_17405,N_17908);
xor U22149 (N_22149,N_15063,N_18405);
nor U22150 (N_22150,N_15548,N_17016);
or U22151 (N_22151,N_18263,N_17692);
nor U22152 (N_22152,N_16796,N_19168);
xnor U22153 (N_22153,N_15808,N_19261);
nor U22154 (N_22154,N_19943,N_19834);
xor U22155 (N_22155,N_16030,N_17238);
or U22156 (N_22156,N_19159,N_16066);
and U22157 (N_22157,N_16688,N_15193);
nand U22158 (N_22158,N_19339,N_17615);
nand U22159 (N_22159,N_19963,N_16757);
nand U22160 (N_22160,N_15540,N_17264);
or U22161 (N_22161,N_15133,N_17175);
xor U22162 (N_22162,N_15138,N_19790);
or U22163 (N_22163,N_17829,N_18623);
nand U22164 (N_22164,N_15609,N_15544);
or U22165 (N_22165,N_18629,N_16550);
nor U22166 (N_22166,N_18025,N_17158);
or U22167 (N_22167,N_16663,N_19565);
nor U22168 (N_22168,N_16566,N_17752);
xnor U22169 (N_22169,N_19587,N_16033);
or U22170 (N_22170,N_15957,N_17395);
nand U22171 (N_22171,N_19816,N_19147);
or U22172 (N_22172,N_18108,N_16937);
or U22173 (N_22173,N_19720,N_17542);
and U22174 (N_22174,N_19218,N_16737);
or U22175 (N_22175,N_18550,N_16425);
and U22176 (N_22176,N_15775,N_17280);
and U22177 (N_22177,N_19087,N_19622);
nor U22178 (N_22178,N_16631,N_17176);
xnor U22179 (N_22179,N_15753,N_18178);
nand U22180 (N_22180,N_16747,N_16415);
and U22181 (N_22181,N_16147,N_16868);
nand U22182 (N_22182,N_19703,N_19971);
and U22183 (N_22183,N_15832,N_17387);
or U22184 (N_22184,N_19115,N_19789);
and U22185 (N_22185,N_19951,N_18604);
nand U22186 (N_22186,N_17447,N_17717);
xor U22187 (N_22187,N_17321,N_19997);
and U22188 (N_22188,N_16706,N_19156);
nand U22189 (N_22189,N_15495,N_18552);
nor U22190 (N_22190,N_16898,N_18212);
or U22191 (N_22191,N_19059,N_15718);
nor U22192 (N_22192,N_16211,N_19439);
nand U22193 (N_22193,N_19777,N_18086);
nand U22194 (N_22194,N_17813,N_16016);
xnor U22195 (N_22195,N_15620,N_17814);
xnor U22196 (N_22196,N_17547,N_19811);
nor U22197 (N_22197,N_15144,N_17774);
or U22198 (N_22198,N_15731,N_18241);
nand U22199 (N_22199,N_15277,N_16195);
and U22200 (N_22200,N_17279,N_16132);
xnor U22201 (N_22201,N_15857,N_15324);
xor U22202 (N_22202,N_19767,N_18992);
xnor U22203 (N_22203,N_19301,N_17093);
or U22204 (N_22204,N_17223,N_17084);
or U22205 (N_22205,N_19474,N_17410);
and U22206 (N_22206,N_17112,N_18626);
nand U22207 (N_22207,N_17879,N_17913);
and U22208 (N_22208,N_19719,N_16355);
xnor U22209 (N_22209,N_19922,N_16010);
nand U22210 (N_22210,N_18357,N_19473);
xnor U22211 (N_22211,N_16391,N_17302);
and U22212 (N_22212,N_15474,N_17591);
and U22213 (N_22213,N_18180,N_15575);
nor U22214 (N_22214,N_17398,N_16046);
nand U22215 (N_22215,N_19691,N_19967);
xor U22216 (N_22216,N_18050,N_18177);
nor U22217 (N_22217,N_18147,N_18738);
nor U22218 (N_22218,N_18432,N_15580);
nand U22219 (N_22219,N_15426,N_16787);
or U22220 (N_22220,N_17086,N_18602);
and U22221 (N_22221,N_18768,N_15204);
nand U22222 (N_22222,N_19962,N_19829);
nand U22223 (N_22223,N_16760,N_17154);
xnor U22224 (N_22224,N_15013,N_18062);
and U22225 (N_22225,N_17048,N_17483);
or U22226 (N_22226,N_16988,N_16735);
and U22227 (N_22227,N_16160,N_15416);
xnor U22228 (N_22228,N_17090,N_17801);
or U22229 (N_22229,N_17201,N_19238);
xnor U22230 (N_22230,N_16257,N_18511);
nand U22231 (N_22231,N_15768,N_16655);
xnor U22232 (N_22232,N_17771,N_15608);
and U22233 (N_22233,N_17538,N_16977);
xnor U22234 (N_22234,N_19883,N_17289);
or U22235 (N_22235,N_19998,N_17599);
nor U22236 (N_22236,N_18729,N_18529);
xnor U22237 (N_22237,N_18624,N_17737);
and U22238 (N_22238,N_19617,N_19535);
and U22239 (N_22239,N_15091,N_16043);
xor U22240 (N_22240,N_19306,N_16532);
and U22241 (N_22241,N_18322,N_15074);
nor U22242 (N_22242,N_18133,N_18727);
xor U22243 (N_22243,N_16813,N_17205);
or U22244 (N_22244,N_18507,N_19670);
or U22245 (N_22245,N_16798,N_17922);
nand U22246 (N_22246,N_19499,N_18760);
xor U22247 (N_22247,N_15121,N_18540);
and U22248 (N_22248,N_16913,N_17626);
xor U22249 (N_22249,N_18472,N_15872);
or U22250 (N_22250,N_17337,N_16711);
nor U22251 (N_22251,N_16271,N_17864);
xor U22252 (N_22252,N_16095,N_18665);
nand U22253 (N_22253,N_16321,N_15201);
xor U22254 (N_22254,N_18548,N_15885);
nand U22255 (N_22255,N_15750,N_16835);
xnor U22256 (N_22256,N_17598,N_17748);
xnor U22257 (N_22257,N_15499,N_17193);
xnor U22258 (N_22258,N_16127,N_18295);
and U22259 (N_22259,N_16815,N_17635);
nand U22260 (N_22260,N_18501,N_17556);
and U22261 (N_22261,N_18510,N_17221);
nand U22262 (N_22262,N_17063,N_17564);
nand U22263 (N_22263,N_15987,N_16833);
or U22264 (N_22264,N_19485,N_17777);
and U22265 (N_22265,N_15820,N_19744);
or U22266 (N_22266,N_19855,N_15691);
nand U22267 (N_22267,N_15113,N_15689);
xor U22268 (N_22268,N_17843,N_15430);
nor U22269 (N_22269,N_15757,N_19120);
nand U22270 (N_22270,N_17715,N_15514);
nor U22271 (N_22271,N_17978,N_18572);
nand U22272 (N_22272,N_15782,N_15871);
nor U22273 (N_22273,N_16459,N_16774);
and U22274 (N_22274,N_16508,N_16080);
xor U22275 (N_22275,N_15785,N_18375);
and U22276 (N_22276,N_18505,N_15786);
nand U22277 (N_22277,N_18537,N_17243);
and U22278 (N_22278,N_18591,N_16838);
or U22279 (N_22279,N_17009,N_15859);
nor U22280 (N_22280,N_17472,N_16322);
nor U22281 (N_22281,N_19453,N_16874);
and U22282 (N_22282,N_18857,N_15025);
nor U22283 (N_22283,N_16948,N_18464);
or U22284 (N_22284,N_18608,N_18217);
and U22285 (N_22285,N_16395,N_15290);
xor U22286 (N_22286,N_16136,N_17298);
xnor U22287 (N_22287,N_17727,N_17217);
xnor U22288 (N_22288,N_18959,N_16329);
and U22289 (N_22289,N_16204,N_17184);
or U22290 (N_22290,N_16678,N_19093);
nand U22291 (N_22291,N_16018,N_19667);
xor U22292 (N_22292,N_19073,N_16893);
nand U22293 (N_22293,N_19350,N_18855);
nand U22294 (N_22294,N_15637,N_19526);
nand U22295 (N_22295,N_19562,N_16502);
or U22296 (N_22296,N_17363,N_16351);
or U22297 (N_22297,N_19364,N_17378);
nand U22298 (N_22298,N_16736,N_15683);
and U22299 (N_22299,N_19915,N_18385);
xnor U22300 (N_22300,N_16630,N_17005);
xnor U22301 (N_22301,N_18869,N_16681);
xor U22302 (N_22302,N_15477,N_17583);
and U22303 (N_22303,N_16848,N_18761);
and U22304 (N_22304,N_17924,N_17758);
xor U22305 (N_22305,N_17007,N_19215);
nand U22306 (N_22306,N_19577,N_19143);
xor U22307 (N_22307,N_15101,N_16943);
or U22308 (N_22308,N_19023,N_15986);
xor U22309 (N_22309,N_16909,N_18365);
xor U22310 (N_22310,N_18105,N_16743);
nand U22311 (N_22311,N_15322,N_18707);
and U22312 (N_22312,N_17012,N_16702);
nor U22313 (N_22313,N_17800,N_16213);
or U22314 (N_22314,N_18297,N_16933);
xor U22315 (N_22315,N_18361,N_17110);
or U22316 (N_22316,N_16512,N_19659);
xnor U22317 (N_22317,N_15671,N_19804);
or U22318 (N_22318,N_18649,N_17265);
xor U22319 (N_22319,N_16124,N_15393);
xor U22320 (N_22320,N_17394,N_15804);
nand U22321 (N_22321,N_18172,N_17234);
nor U22322 (N_22322,N_15307,N_15482);
nor U22323 (N_22323,N_17923,N_19668);
or U22324 (N_22324,N_17450,N_19821);
or U22325 (N_22325,N_19512,N_15463);
nor U22326 (N_22326,N_18005,N_15081);
nor U22327 (N_22327,N_16809,N_17478);
or U22328 (N_22328,N_15863,N_18099);
and U22329 (N_22329,N_16122,N_17871);
nor U22330 (N_22330,N_15100,N_19548);
or U22331 (N_22331,N_18526,N_15022);
nor U22332 (N_22332,N_19088,N_15965);
and U22333 (N_22333,N_15603,N_17991);
xnor U22334 (N_22334,N_18879,N_17425);
and U22335 (N_22335,N_18832,N_18509);
or U22336 (N_22336,N_18314,N_17822);
and U22337 (N_22337,N_18878,N_19090);
xnor U22338 (N_22338,N_17915,N_17019);
nor U22339 (N_22339,N_15082,N_18457);
and U22340 (N_22340,N_18656,N_15299);
xor U22341 (N_22341,N_16472,N_19323);
nor U22342 (N_22342,N_19826,N_15455);
nor U22343 (N_22343,N_15765,N_16253);
nand U22344 (N_22344,N_16427,N_16144);
xnor U22345 (N_22345,N_15310,N_17203);
and U22346 (N_22346,N_15050,N_18798);
or U22347 (N_22347,N_15641,N_17551);
nor U22348 (N_22348,N_18083,N_16925);
or U22349 (N_22349,N_19596,N_18756);
nand U22350 (N_22350,N_17451,N_19686);
or U22351 (N_22351,N_19664,N_16368);
nor U22352 (N_22352,N_17847,N_15180);
xor U22353 (N_22353,N_16264,N_15934);
xnor U22354 (N_22354,N_19823,N_15914);
nand U22355 (N_22355,N_19807,N_18773);
nand U22356 (N_22356,N_17216,N_15502);
nor U22357 (N_22357,N_17702,N_18596);
xor U22358 (N_22358,N_17054,N_19524);
and U22359 (N_22359,N_19511,N_15549);
and U22360 (N_22360,N_16366,N_18085);
or U22361 (N_22361,N_15759,N_19846);
and U22362 (N_22362,N_19195,N_16923);
nor U22363 (N_22363,N_18176,N_19028);
nor U22364 (N_22364,N_17565,N_17240);
xnor U22365 (N_22365,N_19369,N_18718);
xnor U22366 (N_22366,N_17495,N_17990);
nand U22367 (N_22367,N_16035,N_17938);
or U22368 (N_22368,N_17732,N_15301);
or U22369 (N_22369,N_17736,N_15376);
nor U22370 (N_22370,N_16565,N_18354);
and U22371 (N_22371,N_16375,N_18225);
or U22372 (N_22372,N_18174,N_17477);
nor U22373 (N_22373,N_19723,N_19800);
nand U22374 (N_22374,N_19569,N_17229);
and U22375 (N_22375,N_17582,N_16031);
nand U22376 (N_22376,N_16714,N_18200);
and U22377 (N_22377,N_19163,N_15664);
or U22378 (N_22378,N_15837,N_16548);
and U22379 (N_22379,N_15189,N_15610);
and U22380 (N_22380,N_16403,N_19045);
or U22381 (N_22381,N_16413,N_15390);
nor U22382 (N_22382,N_17963,N_16920);
and U22383 (N_22383,N_18607,N_16019);
or U22384 (N_22384,N_16013,N_15380);
nand U22385 (N_22385,N_18644,N_16475);
and U22386 (N_22386,N_17068,N_19545);
or U22387 (N_22387,N_16841,N_15684);
nor U22388 (N_22388,N_16578,N_19894);
nand U22389 (N_22389,N_17517,N_19994);
nand U22390 (N_22390,N_16793,N_16941);
nand U22391 (N_22391,N_19322,N_17731);
or U22392 (N_22392,N_17061,N_19869);
nand U22393 (N_22393,N_16429,N_17608);
and U22394 (N_22394,N_17634,N_15744);
nor U22395 (N_22395,N_17724,N_19543);
and U22396 (N_22396,N_16201,N_18273);
or U22397 (N_22397,N_17031,N_17008);
and U22398 (N_22398,N_15218,N_16811);
nand U22399 (N_22399,N_17523,N_15383);
and U22400 (N_22400,N_15908,N_18606);
nand U22401 (N_22401,N_18214,N_15995);
nor U22402 (N_22402,N_17992,N_17987);
and U22403 (N_22403,N_16504,N_19209);
xor U22404 (N_22404,N_16795,N_17018);
xnor U22405 (N_22405,N_18999,N_15444);
xor U22406 (N_22406,N_17253,N_19597);
and U22407 (N_22407,N_17231,N_19694);
nand U22408 (N_22408,N_18386,N_16585);
and U22409 (N_22409,N_16184,N_16299);
and U22410 (N_22410,N_16646,N_18942);
xor U22411 (N_22411,N_16647,N_18104);
xor U22412 (N_22412,N_19544,N_15459);
nor U22413 (N_22413,N_17557,N_15143);
nand U22414 (N_22414,N_16730,N_17807);
or U22415 (N_22415,N_17562,N_15579);
nand U22416 (N_22416,N_18371,N_16007);
or U22417 (N_22417,N_16312,N_19171);
and U22418 (N_22418,N_19395,N_15382);
or U22419 (N_22419,N_19429,N_17948);
or U22420 (N_22420,N_18265,N_17101);
or U22421 (N_22421,N_17165,N_19484);
and U22422 (N_22422,N_17083,N_16847);
or U22423 (N_22423,N_17631,N_17827);
xnor U22424 (N_22424,N_18159,N_15279);
or U22425 (N_22425,N_19530,N_19360);
or U22426 (N_22426,N_17601,N_19097);
nand U22427 (N_22427,N_19590,N_16764);
nor U22428 (N_22428,N_17857,N_19325);
xnor U22429 (N_22429,N_15010,N_17560);
and U22430 (N_22430,N_17806,N_18584);
and U22431 (N_22431,N_19236,N_19677);
and U22432 (N_22432,N_18977,N_15519);
nand U22433 (N_22433,N_19137,N_18382);
nand U22434 (N_22434,N_16357,N_19605);
nor U22435 (N_22435,N_15003,N_15345);
or U22436 (N_22436,N_19305,N_16235);
or U22437 (N_22437,N_17641,N_17980);
and U22438 (N_22438,N_15140,N_19506);
or U22439 (N_22439,N_18452,N_16836);
nand U22440 (N_22440,N_15260,N_16715);
nand U22441 (N_22441,N_18173,N_16390);
nand U22442 (N_22442,N_18340,N_17756);
and U22443 (N_22443,N_19178,N_17549);
or U22444 (N_22444,N_15311,N_17735);
nor U22445 (N_22445,N_17413,N_16858);
xnor U22446 (N_22446,N_19566,N_16381);
nor U22447 (N_22447,N_15929,N_19355);
xor U22448 (N_22448,N_15904,N_19329);
and U22449 (N_22449,N_17642,N_16338);
or U22450 (N_22450,N_17846,N_19287);
and U22451 (N_22451,N_18966,N_15206);
xor U22452 (N_22452,N_18351,N_17881);
xnor U22453 (N_22453,N_19910,N_15651);
nor U22454 (N_22454,N_18580,N_17421);
xor U22455 (N_22455,N_16547,N_18554);
nand U22456 (N_22456,N_16323,N_19758);
xnor U22457 (N_22457,N_19446,N_15991);
nor U22458 (N_22458,N_16805,N_18944);
nor U22459 (N_22459,N_17993,N_19583);
xor U22460 (N_22460,N_17196,N_18923);
nor U22461 (N_22461,N_16334,N_15901);
nand U22462 (N_22462,N_16176,N_19202);
nor U22463 (N_22463,N_15045,N_17989);
and U22464 (N_22464,N_15316,N_18916);
nor U22465 (N_22465,N_18844,N_19649);
and U22466 (N_22466,N_17492,N_15317);
nor U22467 (N_22467,N_16718,N_16476);
and U22468 (N_22468,N_15071,N_18036);
nand U22469 (N_22469,N_16199,N_19642);
nand U22470 (N_22470,N_16535,N_15089);
xnor U22471 (N_22471,N_18246,N_16594);
xnor U22472 (N_22472,N_15591,N_19190);
nand U22473 (N_22473,N_17057,N_16263);
xor U22474 (N_22474,N_18210,N_19342);
and U22475 (N_22475,N_16441,N_18634);
and U22476 (N_22476,N_18638,N_18168);
xor U22477 (N_22477,N_17037,N_18163);
or U22478 (N_22478,N_19712,N_18119);
xor U22479 (N_22479,N_15612,N_19768);
nor U22480 (N_22480,N_17494,N_16785);
nand U22481 (N_22481,N_15973,N_19508);
xor U22482 (N_22482,N_19053,N_15721);
nand U22483 (N_22483,N_19293,N_19743);
nand U22484 (N_22484,N_17159,N_19108);
or U22485 (N_22485,N_16408,N_15250);
and U22486 (N_22486,N_19385,N_15048);
or U22487 (N_22487,N_17058,N_16219);
xnor U22488 (N_22488,N_19278,N_19275);
or U22489 (N_22489,N_15172,N_16644);
nor U22490 (N_22490,N_15662,N_16025);
and U22491 (N_22491,N_16040,N_18114);
xnor U22492 (N_22492,N_16541,N_18380);
or U22493 (N_22493,N_17153,N_15116);
and U22494 (N_22494,N_17036,N_18907);
xnor U22495 (N_22495,N_19251,N_16451);
xor U22496 (N_22496,N_17606,N_15167);
nor U22497 (N_22497,N_15276,N_19509);
nand U22498 (N_22498,N_18759,N_19109);
nand U22499 (N_22499,N_17896,N_19206);
xnor U22500 (N_22500,N_19555,N_15171);
nor U22501 (N_22501,N_18003,N_18347);
nor U22502 (N_22502,N_17538,N_19161);
nor U22503 (N_22503,N_18017,N_15972);
and U22504 (N_22504,N_16437,N_15849);
nor U22505 (N_22505,N_19796,N_19738);
nor U22506 (N_22506,N_19435,N_19312);
xor U22507 (N_22507,N_19148,N_16882);
and U22508 (N_22508,N_16156,N_15207);
xor U22509 (N_22509,N_16979,N_15596);
xor U22510 (N_22510,N_19985,N_17882);
nor U22511 (N_22511,N_18548,N_17645);
and U22512 (N_22512,N_19010,N_15886);
or U22513 (N_22513,N_15508,N_17365);
or U22514 (N_22514,N_16379,N_16904);
and U22515 (N_22515,N_18190,N_19317);
and U22516 (N_22516,N_19416,N_17211);
or U22517 (N_22517,N_16608,N_19789);
xnor U22518 (N_22518,N_18961,N_16097);
or U22519 (N_22519,N_19708,N_15547);
or U22520 (N_22520,N_16817,N_16068);
nor U22521 (N_22521,N_18821,N_16601);
nand U22522 (N_22522,N_16377,N_16481);
or U22523 (N_22523,N_16108,N_16613);
and U22524 (N_22524,N_19657,N_16004);
nor U22525 (N_22525,N_16516,N_19836);
nor U22526 (N_22526,N_15956,N_16875);
and U22527 (N_22527,N_16532,N_19571);
xor U22528 (N_22528,N_18389,N_19576);
or U22529 (N_22529,N_15694,N_19828);
nand U22530 (N_22530,N_15271,N_16703);
and U22531 (N_22531,N_16614,N_15659);
and U22532 (N_22532,N_17372,N_15240);
and U22533 (N_22533,N_18798,N_16186);
xnor U22534 (N_22534,N_19858,N_17500);
xor U22535 (N_22535,N_16913,N_19869);
xor U22536 (N_22536,N_18677,N_15075);
and U22537 (N_22537,N_18396,N_15385);
xnor U22538 (N_22538,N_17650,N_17107);
or U22539 (N_22539,N_18618,N_18248);
and U22540 (N_22540,N_15241,N_16626);
nor U22541 (N_22541,N_19127,N_15071);
or U22542 (N_22542,N_16325,N_19068);
and U22543 (N_22543,N_16182,N_15070);
nand U22544 (N_22544,N_17740,N_15040);
or U22545 (N_22545,N_17478,N_17217);
xor U22546 (N_22546,N_19173,N_15230);
and U22547 (N_22547,N_19640,N_19054);
nand U22548 (N_22548,N_18413,N_18132);
or U22549 (N_22549,N_17260,N_16227);
and U22550 (N_22550,N_19228,N_19571);
xnor U22551 (N_22551,N_19226,N_15577);
xor U22552 (N_22552,N_15191,N_18829);
and U22553 (N_22553,N_15179,N_16106);
and U22554 (N_22554,N_17462,N_17541);
nand U22555 (N_22555,N_18060,N_17503);
or U22556 (N_22556,N_15691,N_19306);
xnor U22557 (N_22557,N_15128,N_16128);
xnor U22558 (N_22558,N_19642,N_19728);
xor U22559 (N_22559,N_19681,N_19106);
nand U22560 (N_22560,N_15060,N_19314);
nand U22561 (N_22561,N_16537,N_16988);
or U22562 (N_22562,N_15721,N_17875);
and U22563 (N_22563,N_19241,N_19453);
nor U22564 (N_22564,N_18361,N_19552);
and U22565 (N_22565,N_19727,N_19734);
nor U22566 (N_22566,N_17322,N_15136);
and U22567 (N_22567,N_17007,N_18387);
or U22568 (N_22568,N_16238,N_19353);
nand U22569 (N_22569,N_18927,N_19244);
nand U22570 (N_22570,N_18335,N_16965);
nand U22571 (N_22571,N_16200,N_18787);
nor U22572 (N_22572,N_18796,N_17272);
xnor U22573 (N_22573,N_17449,N_16183);
and U22574 (N_22574,N_16736,N_18323);
xnor U22575 (N_22575,N_15012,N_18960);
or U22576 (N_22576,N_19422,N_19397);
or U22577 (N_22577,N_16360,N_18990);
nor U22578 (N_22578,N_16852,N_16466);
xor U22579 (N_22579,N_17446,N_17649);
and U22580 (N_22580,N_17231,N_16503);
xnor U22581 (N_22581,N_19818,N_19674);
and U22582 (N_22582,N_16975,N_15631);
nor U22583 (N_22583,N_15987,N_17858);
or U22584 (N_22584,N_19125,N_15447);
and U22585 (N_22585,N_18431,N_18550);
and U22586 (N_22586,N_19601,N_15271);
nand U22587 (N_22587,N_16701,N_18674);
nand U22588 (N_22588,N_15593,N_18790);
or U22589 (N_22589,N_17688,N_16077);
nand U22590 (N_22590,N_19893,N_16538);
and U22591 (N_22591,N_19991,N_17355);
or U22592 (N_22592,N_17845,N_16025);
or U22593 (N_22593,N_17913,N_16517);
nor U22594 (N_22594,N_18316,N_19351);
nand U22595 (N_22595,N_15663,N_17543);
nand U22596 (N_22596,N_17832,N_18129);
and U22597 (N_22597,N_16952,N_18218);
and U22598 (N_22598,N_15458,N_16531);
nor U22599 (N_22599,N_17637,N_18096);
nor U22600 (N_22600,N_18628,N_17759);
or U22601 (N_22601,N_16733,N_19361);
nor U22602 (N_22602,N_19620,N_19063);
nand U22603 (N_22603,N_15024,N_17760);
and U22604 (N_22604,N_17124,N_19695);
nand U22605 (N_22605,N_17883,N_18487);
nor U22606 (N_22606,N_17201,N_18930);
xor U22607 (N_22607,N_18802,N_17806);
xor U22608 (N_22608,N_17924,N_15627);
and U22609 (N_22609,N_18718,N_18368);
xor U22610 (N_22610,N_19387,N_18667);
or U22611 (N_22611,N_19770,N_16729);
and U22612 (N_22612,N_17517,N_15396);
xor U22613 (N_22613,N_18630,N_16671);
and U22614 (N_22614,N_18849,N_16231);
nand U22615 (N_22615,N_18415,N_15148);
nand U22616 (N_22616,N_15970,N_16138);
nand U22617 (N_22617,N_16873,N_15374);
nor U22618 (N_22618,N_16323,N_16793);
xor U22619 (N_22619,N_15616,N_17315);
or U22620 (N_22620,N_15796,N_17675);
nor U22621 (N_22621,N_18965,N_18624);
and U22622 (N_22622,N_16513,N_17107);
nor U22623 (N_22623,N_19758,N_15692);
or U22624 (N_22624,N_19773,N_16859);
nand U22625 (N_22625,N_19570,N_16416);
nor U22626 (N_22626,N_16466,N_16222);
or U22627 (N_22627,N_17736,N_18930);
and U22628 (N_22628,N_19176,N_18952);
nand U22629 (N_22629,N_19450,N_16366);
and U22630 (N_22630,N_17576,N_16310);
or U22631 (N_22631,N_18609,N_18036);
or U22632 (N_22632,N_18955,N_18361);
or U22633 (N_22633,N_18253,N_15407);
xor U22634 (N_22634,N_16691,N_18963);
nor U22635 (N_22635,N_18636,N_15776);
nand U22636 (N_22636,N_19576,N_17610);
nand U22637 (N_22637,N_16557,N_19067);
xor U22638 (N_22638,N_18592,N_17398);
nand U22639 (N_22639,N_17592,N_15124);
xnor U22640 (N_22640,N_16791,N_19958);
and U22641 (N_22641,N_19857,N_18514);
nor U22642 (N_22642,N_15074,N_18561);
or U22643 (N_22643,N_17376,N_15600);
nand U22644 (N_22644,N_15710,N_18902);
nand U22645 (N_22645,N_17419,N_15160);
xnor U22646 (N_22646,N_18260,N_17261);
nand U22647 (N_22647,N_16732,N_17099);
xnor U22648 (N_22648,N_16911,N_16525);
nand U22649 (N_22649,N_15099,N_19717);
nor U22650 (N_22650,N_16629,N_18204);
or U22651 (N_22651,N_15674,N_15940);
nor U22652 (N_22652,N_16162,N_16077);
nor U22653 (N_22653,N_16958,N_19152);
nand U22654 (N_22654,N_18217,N_15518);
and U22655 (N_22655,N_15397,N_18987);
nand U22656 (N_22656,N_17155,N_17686);
and U22657 (N_22657,N_16520,N_17410);
xor U22658 (N_22658,N_15890,N_16776);
nand U22659 (N_22659,N_19518,N_18242);
nand U22660 (N_22660,N_17087,N_16136);
xnor U22661 (N_22661,N_16471,N_16513);
nor U22662 (N_22662,N_17318,N_18938);
xor U22663 (N_22663,N_17649,N_19364);
and U22664 (N_22664,N_15128,N_19123);
and U22665 (N_22665,N_16738,N_17076);
or U22666 (N_22666,N_18591,N_18325);
or U22667 (N_22667,N_18026,N_16663);
nand U22668 (N_22668,N_18793,N_18750);
xnor U22669 (N_22669,N_18814,N_15899);
nand U22670 (N_22670,N_16245,N_15012);
or U22671 (N_22671,N_15821,N_19252);
or U22672 (N_22672,N_16573,N_15512);
nand U22673 (N_22673,N_18562,N_16534);
or U22674 (N_22674,N_17559,N_17461);
and U22675 (N_22675,N_19021,N_18426);
and U22676 (N_22676,N_18962,N_19618);
nand U22677 (N_22677,N_16997,N_18177);
xor U22678 (N_22678,N_15667,N_19626);
or U22679 (N_22679,N_16335,N_16871);
xor U22680 (N_22680,N_18449,N_17473);
or U22681 (N_22681,N_16082,N_17380);
or U22682 (N_22682,N_18679,N_15265);
nand U22683 (N_22683,N_19962,N_16863);
nand U22684 (N_22684,N_16627,N_19145);
nand U22685 (N_22685,N_19070,N_16809);
xnor U22686 (N_22686,N_16432,N_18997);
xnor U22687 (N_22687,N_19318,N_19705);
nand U22688 (N_22688,N_19735,N_18213);
or U22689 (N_22689,N_19111,N_18562);
xor U22690 (N_22690,N_16905,N_16264);
xnor U22691 (N_22691,N_15033,N_19416);
nor U22692 (N_22692,N_16515,N_18097);
nor U22693 (N_22693,N_19268,N_19382);
xor U22694 (N_22694,N_19012,N_15542);
xnor U22695 (N_22695,N_15364,N_17941);
nand U22696 (N_22696,N_19420,N_18876);
nand U22697 (N_22697,N_17902,N_16388);
nor U22698 (N_22698,N_18355,N_18124);
or U22699 (N_22699,N_18804,N_19497);
nor U22700 (N_22700,N_19705,N_16107);
and U22701 (N_22701,N_18060,N_16435);
and U22702 (N_22702,N_17133,N_15581);
and U22703 (N_22703,N_19675,N_17866);
xor U22704 (N_22704,N_17422,N_15985);
xor U22705 (N_22705,N_18426,N_18640);
nand U22706 (N_22706,N_17980,N_19529);
nor U22707 (N_22707,N_19540,N_17249);
and U22708 (N_22708,N_15739,N_17316);
nand U22709 (N_22709,N_18784,N_16374);
nand U22710 (N_22710,N_17938,N_16419);
or U22711 (N_22711,N_16159,N_17775);
nand U22712 (N_22712,N_19641,N_15961);
xor U22713 (N_22713,N_18864,N_19970);
xnor U22714 (N_22714,N_15477,N_16399);
xor U22715 (N_22715,N_15947,N_15116);
or U22716 (N_22716,N_15023,N_16610);
and U22717 (N_22717,N_15496,N_18481);
and U22718 (N_22718,N_18343,N_15702);
or U22719 (N_22719,N_15645,N_19532);
nand U22720 (N_22720,N_19581,N_17436);
or U22721 (N_22721,N_17402,N_16326);
or U22722 (N_22722,N_16052,N_15229);
nor U22723 (N_22723,N_15462,N_16565);
nor U22724 (N_22724,N_18567,N_16002);
or U22725 (N_22725,N_18948,N_16403);
nor U22726 (N_22726,N_17074,N_18164);
nand U22727 (N_22727,N_15569,N_16672);
xor U22728 (N_22728,N_18819,N_19669);
or U22729 (N_22729,N_18410,N_16047);
xnor U22730 (N_22730,N_17541,N_16423);
nor U22731 (N_22731,N_19665,N_15603);
nand U22732 (N_22732,N_19243,N_18147);
nor U22733 (N_22733,N_16971,N_17717);
nand U22734 (N_22734,N_19171,N_16649);
nor U22735 (N_22735,N_16404,N_16459);
nor U22736 (N_22736,N_15728,N_16441);
and U22737 (N_22737,N_18138,N_16603);
nand U22738 (N_22738,N_19445,N_16926);
nor U22739 (N_22739,N_19393,N_15145);
xor U22740 (N_22740,N_16211,N_19022);
xnor U22741 (N_22741,N_19581,N_16068);
xor U22742 (N_22742,N_15983,N_18278);
or U22743 (N_22743,N_18208,N_18879);
and U22744 (N_22744,N_16600,N_15444);
xor U22745 (N_22745,N_15914,N_18383);
or U22746 (N_22746,N_19722,N_15119);
or U22747 (N_22747,N_18555,N_15764);
xnor U22748 (N_22748,N_18459,N_19815);
nand U22749 (N_22749,N_15971,N_19338);
or U22750 (N_22750,N_15001,N_18168);
and U22751 (N_22751,N_18203,N_17420);
nor U22752 (N_22752,N_19577,N_19251);
or U22753 (N_22753,N_16645,N_19732);
and U22754 (N_22754,N_18422,N_15194);
nand U22755 (N_22755,N_17944,N_17177);
or U22756 (N_22756,N_18465,N_19372);
nand U22757 (N_22757,N_15595,N_18412);
or U22758 (N_22758,N_19136,N_17628);
nor U22759 (N_22759,N_15933,N_18665);
and U22760 (N_22760,N_18822,N_18541);
nand U22761 (N_22761,N_17147,N_16722);
xor U22762 (N_22762,N_15167,N_17599);
and U22763 (N_22763,N_18869,N_15093);
and U22764 (N_22764,N_17409,N_15944);
and U22765 (N_22765,N_17541,N_19442);
nor U22766 (N_22766,N_19041,N_18699);
nor U22767 (N_22767,N_15380,N_17109);
nor U22768 (N_22768,N_16636,N_18321);
or U22769 (N_22769,N_15867,N_19236);
or U22770 (N_22770,N_15741,N_18482);
nor U22771 (N_22771,N_16573,N_19687);
nand U22772 (N_22772,N_16920,N_15235);
or U22773 (N_22773,N_17348,N_17138);
and U22774 (N_22774,N_19468,N_16183);
or U22775 (N_22775,N_16075,N_17053);
xor U22776 (N_22776,N_18685,N_19779);
or U22777 (N_22777,N_15302,N_19776);
nand U22778 (N_22778,N_17727,N_15670);
nand U22779 (N_22779,N_19679,N_18228);
nand U22780 (N_22780,N_19149,N_18394);
and U22781 (N_22781,N_19471,N_18583);
xnor U22782 (N_22782,N_15277,N_16414);
or U22783 (N_22783,N_15951,N_17677);
and U22784 (N_22784,N_17314,N_17800);
and U22785 (N_22785,N_17163,N_16863);
or U22786 (N_22786,N_15032,N_17450);
nor U22787 (N_22787,N_18497,N_17639);
or U22788 (N_22788,N_17214,N_16535);
xnor U22789 (N_22789,N_18414,N_18245);
nand U22790 (N_22790,N_17869,N_16828);
nand U22791 (N_22791,N_15155,N_16453);
xor U22792 (N_22792,N_19673,N_15379);
xnor U22793 (N_22793,N_19657,N_17905);
and U22794 (N_22794,N_17396,N_17037);
and U22795 (N_22795,N_18113,N_15615);
and U22796 (N_22796,N_16222,N_16441);
or U22797 (N_22797,N_17360,N_17371);
xnor U22798 (N_22798,N_15122,N_17553);
xnor U22799 (N_22799,N_19332,N_17649);
nand U22800 (N_22800,N_17961,N_17592);
xnor U22801 (N_22801,N_17538,N_16249);
or U22802 (N_22802,N_17085,N_18686);
or U22803 (N_22803,N_18375,N_18362);
nand U22804 (N_22804,N_18236,N_17848);
xor U22805 (N_22805,N_18309,N_16485);
nor U22806 (N_22806,N_17683,N_19121);
or U22807 (N_22807,N_19362,N_16335);
or U22808 (N_22808,N_15132,N_18782);
or U22809 (N_22809,N_19747,N_19332);
nand U22810 (N_22810,N_19278,N_15842);
and U22811 (N_22811,N_16724,N_16046);
xor U22812 (N_22812,N_15133,N_15492);
nor U22813 (N_22813,N_15340,N_18760);
xor U22814 (N_22814,N_18585,N_18696);
and U22815 (N_22815,N_16353,N_17324);
and U22816 (N_22816,N_18125,N_16178);
and U22817 (N_22817,N_17495,N_17421);
nand U22818 (N_22818,N_19208,N_17731);
and U22819 (N_22819,N_17157,N_18541);
and U22820 (N_22820,N_19010,N_16071);
and U22821 (N_22821,N_17947,N_19640);
xnor U22822 (N_22822,N_17639,N_17622);
nand U22823 (N_22823,N_19290,N_16314);
nand U22824 (N_22824,N_15194,N_16343);
and U22825 (N_22825,N_19207,N_19777);
nor U22826 (N_22826,N_17569,N_16810);
and U22827 (N_22827,N_17342,N_19652);
or U22828 (N_22828,N_17590,N_15279);
or U22829 (N_22829,N_19189,N_15828);
and U22830 (N_22830,N_17979,N_15970);
and U22831 (N_22831,N_17532,N_15433);
nor U22832 (N_22832,N_16500,N_18186);
and U22833 (N_22833,N_19214,N_15244);
and U22834 (N_22834,N_15527,N_19907);
nor U22835 (N_22835,N_17511,N_18248);
nor U22836 (N_22836,N_18734,N_17288);
and U22837 (N_22837,N_19759,N_18834);
and U22838 (N_22838,N_15128,N_17454);
and U22839 (N_22839,N_15094,N_15229);
and U22840 (N_22840,N_17700,N_19916);
nand U22841 (N_22841,N_15906,N_19869);
xnor U22842 (N_22842,N_17176,N_19531);
xor U22843 (N_22843,N_19754,N_16474);
xor U22844 (N_22844,N_17876,N_17502);
and U22845 (N_22845,N_16008,N_19737);
xor U22846 (N_22846,N_19862,N_17142);
xnor U22847 (N_22847,N_19374,N_19325);
xnor U22848 (N_22848,N_19493,N_19910);
xor U22849 (N_22849,N_16740,N_18102);
nor U22850 (N_22850,N_17580,N_17918);
nor U22851 (N_22851,N_19470,N_19221);
and U22852 (N_22852,N_17134,N_16697);
and U22853 (N_22853,N_18866,N_17678);
and U22854 (N_22854,N_19723,N_16735);
and U22855 (N_22855,N_16081,N_16545);
nor U22856 (N_22856,N_15605,N_18357);
xor U22857 (N_22857,N_17383,N_15368);
nand U22858 (N_22858,N_19709,N_15942);
nor U22859 (N_22859,N_16650,N_19112);
nand U22860 (N_22860,N_16046,N_15217);
or U22861 (N_22861,N_18401,N_18653);
or U22862 (N_22862,N_17695,N_15448);
and U22863 (N_22863,N_19492,N_19917);
nor U22864 (N_22864,N_15875,N_19716);
nor U22865 (N_22865,N_16679,N_15726);
or U22866 (N_22866,N_18471,N_18224);
nor U22867 (N_22867,N_17888,N_16915);
and U22868 (N_22868,N_15560,N_17303);
xnor U22869 (N_22869,N_16664,N_17215);
and U22870 (N_22870,N_15951,N_16104);
or U22871 (N_22871,N_17641,N_16690);
nor U22872 (N_22872,N_18140,N_17526);
and U22873 (N_22873,N_19842,N_18908);
and U22874 (N_22874,N_17076,N_18050);
or U22875 (N_22875,N_15052,N_15911);
nand U22876 (N_22876,N_17242,N_18802);
xor U22877 (N_22877,N_19455,N_17884);
nor U22878 (N_22878,N_17568,N_18010);
nor U22879 (N_22879,N_16636,N_16719);
nand U22880 (N_22880,N_19478,N_18083);
nor U22881 (N_22881,N_19328,N_19324);
nand U22882 (N_22882,N_17092,N_17253);
nand U22883 (N_22883,N_17771,N_19137);
and U22884 (N_22884,N_18854,N_18291);
nor U22885 (N_22885,N_17965,N_17900);
or U22886 (N_22886,N_17811,N_16417);
xnor U22887 (N_22887,N_18100,N_16560);
and U22888 (N_22888,N_17756,N_18180);
nor U22889 (N_22889,N_19770,N_17996);
nand U22890 (N_22890,N_19253,N_18984);
xor U22891 (N_22891,N_19376,N_18546);
nand U22892 (N_22892,N_16903,N_18098);
nor U22893 (N_22893,N_16718,N_19652);
nand U22894 (N_22894,N_16102,N_17706);
and U22895 (N_22895,N_15847,N_15814);
and U22896 (N_22896,N_19208,N_17177);
or U22897 (N_22897,N_17013,N_16084);
xnor U22898 (N_22898,N_16126,N_15419);
nand U22899 (N_22899,N_17558,N_19981);
nand U22900 (N_22900,N_19960,N_17008);
nand U22901 (N_22901,N_19854,N_18992);
nor U22902 (N_22902,N_16150,N_15011);
nor U22903 (N_22903,N_18757,N_15666);
nand U22904 (N_22904,N_16990,N_16088);
xor U22905 (N_22905,N_19922,N_18755);
or U22906 (N_22906,N_16668,N_17228);
and U22907 (N_22907,N_19608,N_19853);
nand U22908 (N_22908,N_17841,N_16149);
nand U22909 (N_22909,N_16092,N_18824);
nor U22910 (N_22910,N_17337,N_15107);
or U22911 (N_22911,N_15970,N_18968);
nand U22912 (N_22912,N_19782,N_17189);
nor U22913 (N_22913,N_16975,N_18192);
or U22914 (N_22914,N_16802,N_19816);
xor U22915 (N_22915,N_18748,N_16752);
nand U22916 (N_22916,N_19204,N_18580);
nor U22917 (N_22917,N_15456,N_17290);
or U22918 (N_22918,N_15186,N_17560);
nand U22919 (N_22919,N_19735,N_16927);
nand U22920 (N_22920,N_18940,N_15724);
xnor U22921 (N_22921,N_18330,N_18561);
and U22922 (N_22922,N_16096,N_16905);
xnor U22923 (N_22923,N_17934,N_16789);
and U22924 (N_22924,N_15554,N_15124);
or U22925 (N_22925,N_16925,N_17438);
nand U22926 (N_22926,N_18404,N_18951);
or U22927 (N_22927,N_17375,N_15982);
nor U22928 (N_22928,N_15225,N_17975);
nand U22929 (N_22929,N_15441,N_15979);
or U22930 (N_22930,N_17526,N_16586);
nor U22931 (N_22931,N_17742,N_19500);
nor U22932 (N_22932,N_15063,N_19293);
xnor U22933 (N_22933,N_18807,N_19923);
or U22934 (N_22934,N_19284,N_17547);
or U22935 (N_22935,N_15197,N_16547);
and U22936 (N_22936,N_15973,N_16030);
or U22937 (N_22937,N_15249,N_16634);
xor U22938 (N_22938,N_17287,N_19309);
or U22939 (N_22939,N_18072,N_15118);
nor U22940 (N_22940,N_17213,N_19648);
xor U22941 (N_22941,N_17809,N_18881);
and U22942 (N_22942,N_16688,N_18692);
xnor U22943 (N_22943,N_16502,N_16525);
xnor U22944 (N_22944,N_15732,N_16426);
or U22945 (N_22945,N_15332,N_16491);
nor U22946 (N_22946,N_19230,N_16545);
nor U22947 (N_22947,N_19015,N_19143);
xor U22948 (N_22948,N_19432,N_16206);
nor U22949 (N_22949,N_15300,N_19233);
or U22950 (N_22950,N_18294,N_17529);
xnor U22951 (N_22951,N_15056,N_15623);
and U22952 (N_22952,N_19739,N_19594);
nand U22953 (N_22953,N_15391,N_18859);
or U22954 (N_22954,N_16090,N_19918);
nor U22955 (N_22955,N_19538,N_19180);
nand U22956 (N_22956,N_18100,N_15253);
nor U22957 (N_22957,N_16917,N_16590);
or U22958 (N_22958,N_19924,N_16185);
and U22959 (N_22959,N_15033,N_16548);
and U22960 (N_22960,N_15228,N_18661);
nor U22961 (N_22961,N_19563,N_15879);
nor U22962 (N_22962,N_17234,N_19668);
nand U22963 (N_22963,N_16861,N_18334);
xor U22964 (N_22964,N_17702,N_17536);
xnor U22965 (N_22965,N_19351,N_17212);
xor U22966 (N_22966,N_15483,N_16593);
nor U22967 (N_22967,N_17044,N_19145);
and U22968 (N_22968,N_18609,N_16155);
nor U22969 (N_22969,N_17370,N_17034);
or U22970 (N_22970,N_16673,N_16052);
or U22971 (N_22971,N_15272,N_18376);
nor U22972 (N_22972,N_15250,N_15728);
nor U22973 (N_22973,N_16487,N_19265);
nand U22974 (N_22974,N_18752,N_16713);
or U22975 (N_22975,N_19346,N_18989);
and U22976 (N_22976,N_18716,N_16698);
and U22977 (N_22977,N_15240,N_19342);
nor U22978 (N_22978,N_19193,N_18477);
or U22979 (N_22979,N_19779,N_17218);
and U22980 (N_22980,N_19811,N_19020);
xor U22981 (N_22981,N_15688,N_16390);
xor U22982 (N_22982,N_19117,N_16730);
and U22983 (N_22983,N_18863,N_16850);
or U22984 (N_22984,N_19072,N_19801);
nand U22985 (N_22985,N_18293,N_18615);
nand U22986 (N_22986,N_17619,N_19598);
and U22987 (N_22987,N_16989,N_16624);
xnor U22988 (N_22988,N_17754,N_19428);
nor U22989 (N_22989,N_17833,N_16103);
or U22990 (N_22990,N_18534,N_16989);
nand U22991 (N_22991,N_19889,N_16291);
nand U22992 (N_22992,N_16380,N_16315);
or U22993 (N_22993,N_16709,N_15378);
nand U22994 (N_22994,N_16628,N_19373);
nand U22995 (N_22995,N_19334,N_16775);
or U22996 (N_22996,N_15447,N_18332);
xor U22997 (N_22997,N_19521,N_18685);
nand U22998 (N_22998,N_17844,N_16366);
xor U22999 (N_22999,N_19278,N_18475);
or U23000 (N_23000,N_15052,N_16070);
and U23001 (N_23001,N_19554,N_19444);
nand U23002 (N_23002,N_19518,N_19048);
and U23003 (N_23003,N_17456,N_19324);
xor U23004 (N_23004,N_15901,N_17573);
and U23005 (N_23005,N_18813,N_16463);
nand U23006 (N_23006,N_17969,N_18714);
xnor U23007 (N_23007,N_18724,N_16071);
and U23008 (N_23008,N_17904,N_15601);
or U23009 (N_23009,N_18740,N_15941);
xor U23010 (N_23010,N_16275,N_16749);
xor U23011 (N_23011,N_17015,N_19714);
and U23012 (N_23012,N_18354,N_17396);
and U23013 (N_23013,N_17760,N_19228);
nor U23014 (N_23014,N_18687,N_17249);
nor U23015 (N_23015,N_15121,N_15766);
xnor U23016 (N_23016,N_15219,N_17966);
nor U23017 (N_23017,N_19760,N_16521);
nor U23018 (N_23018,N_16217,N_19586);
xnor U23019 (N_23019,N_17204,N_15006);
nand U23020 (N_23020,N_15307,N_17413);
xor U23021 (N_23021,N_19390,N_16748);
and U23022 (N_23022,N_15592,N_18012);
and U23023 (N_23023,N_17478,N_19194);
xnor U23024 (N_23024,N_16727,N_15648);
nor U23025 (N_23025,N_15745,N_19913);
nor U23026 (N_23026,N_18403,N_15303);
and U23027 (N_23027,N_18376,N_16546);
and U23028 (N_23028,N_19309,N_18760);
nand U23029 (N_23029,N_17203,N_16637);
and U23030 (N_23030,N_17227,N_15491);
xnor U23031 (N_23031,N_19962,N_19872);
and U23032 (N_23032,N_19106,N_17949);
nand U23033 (N_23033,N_17853,N_19574);
and U23034 (N_23034,N_16686,N_18524);
and U23035 (N_23035,N_17742,N_16302);
or U23036 (N_23036,N_16375,N_17847);
xor U23037 (N_23037,N_19180,N_15219);
nand U23038 (N_23038,N_18812,N_15911);
nor U23039 (N_23039,N_19667,N_19036);
or U23040 (N_23040,N_15403,N_19602);
or U23041 (N_23041,N_16460,N_15653);
nor U23042 (N_23042,N_16822,N_16920);
or U23043 (N_23043,N_18341,N_16877);
nand U23044 (N_23044,N_17713,N_17470);
and U23045 (N_23045,N_16972,N_17472);
or U23046 (N_23046,N_15893,N_15660);
xor U23047 (N_23047,N_18744,N_17134);
nor U23048 (N_23048,N_16669,N_17660);
and U23049 (N_23049,N_19227,N_19887);
or U23050 (N_23050,N_18261,N_16021);
nand U23051 (N_23051,N_16434,N_19749);
and U23052 (N_23052,N_18103,N_17878);
nand U23053 (N_23053,N_17839,N_16467);
or U23054 (N_23054,N_19160,N_19373);
or U23055 (N_23055,N_17718,N_15445);
nor U23056 (N_23056,N_18509,N_16990);
or U23057 (N_23057,N_16126,N_19280);
and U23058 (N_23058,N_16419,N_16846);
or U23059 (N_23059,N_16964,N_15751);
nor U23060 (N_23060,N_17436,N_15665);
or U23061 (N_23061,N_16808,N_18021);
nand U23062 (N_23062,N_17220,N_15444);
and U23063 (N_23063,N_19955,N_15800);
nand U23064 (N_23064,N_18086,N_16625);
and U23065 (N_23065,N_19538,N_19513);
nor U23066 (N_23066,N_16328,N_19512);
nor U23067 (N_23067,N_15848,N_19864);
nand U23068 (N_23068,N_19431,N_18202);
nor U23069 (N_23069,N_18485,N_15483);
xor U23070 (N_23070,N_18452,N_17810);
xnor U23071 (N_23071,N_17022,N_17619);
nor U23072 (N_23072,N_17545,N_18508);
or U23073 (N_23073,N_17727,N_18920);
nor U23074 (N_23074,N_17382,N_16843);
xor U23075 (N_23075,N_18591,N_15222);
and U23076 (N_23076,N_15189,N_16698);
xor U23077 (N_23077,N_17435,N_17862);
or U23078 (N_23078,N_16495,N_18137);
and U23079 (N_23079,N_16221,N_16689);
nor U23080 (N_23080,N_16269,N_19899);
nand U23081 (N_23081,N_19369,N_16202);
xor U23082 (N_23082,N_15979,N_18218);
xnor U23083 (N_23083,N_15444,N_16072);
nand U23084 (N_23084,N_19182,N_16649);
or U23085 (N_23085,N_19287,N_19147);
nand U23086 (N_23086,N_18580,N_18971);
xnor U23087 (N_23087,N_16134,N_18254);
nor U23088 (N_23088,N_16491,N_17814);
and U23089 (N_23089,N_19044,N_16829);
nand U23090 (N_23090,N_17184,N_18078);
xnor U23091 (N_23091,N_15983,N_15087);
xnor U23092 (N_23092,N_16569,N_19592);
xnor U23093 (N_23093,N_15046,N_16241);
xor U23094 (N_23094,N_19909,N_15370);
nor U23095 (N_23095,N_17258,N_18917);
xnor U23096 (N_23096,N_18255,N_16076);
nor U23097 (N_23097,N_19346,N_19010);
or U23098 (N_23098,N_16326,N_16688);
and U23099 (N_23099,N_16327,N_17290);
or U23100 (N_23100,N_16902,N_19657);
nand U23101 (N_23101,N_17911,N_19248);
and U23102 (N_23102,N_19290,N_16518);
nor U23103 (N_23103,N_17791,N_18434);
and U23104 (N_23104,N_17504,N_18859);
or U23105 (N_23105,N_18658,N_19686);
nor U23106 (N_23106,N_19955,N_17572);
nand U23107 (N_23107,N_16010,N_17996);
or U23108 (N_23108,N_19076,N_17734);
or U23109 (N_23109,N_18420,N_19471);
xor U23110 (N_23110,N_17717,N_17255);
or U23111 (N_23111,N_16763,N_15452);
xor U23112 (N_23112,N_15113,N_15493);
nor U23113 (N_23113,N_16520,N_16771);
or U23114 (N_23114,N_19529,N_16801);
and U23115 (N_23115,N_17027,N_18875);
nand U23116 (N_23116,N_17027,N_16850);
and U23117 (N_23117,N_19408,N_19289);
or U23118 (N_23118,N_19362,N_15516);
or U23119 (N_23119,N_19340,N_18003);
or U23120 (N_23120,N_17160,N_19122);
nor U23121 (N_23121,N_18931,N_15728);
nand U23122 (N_23122,N_15965,N_19483);
and U23123 (N_23123,N_19050,N_17718);
and U23124 (N_23124,N_16649,N_18604);
and U23125 (N_23125,N_19301,N_17005);
nand U23126 (N_23126,N_18202,N_18431);
xor U23127 (N_23127,N_17053,N_17811);
nand U23128 (N_23128,N_16496,N_15275);
and U23129 (N_23129,N_18359,N_17802);
and U23130 (N_23130,N_18075,N_17330);
or U23131 (N_23131,N_19768,N_15666);
and U23132 (N_23132,N_16426,N_15119);
nand U23133 (N_23133,N_15945,N_19643);
xnor U23134 (N_23134,N_15322,N_15635);
nand U23135 (N_23135,N_15710,N_17224);
nor U23136 (N_23136,N_19206,N_19407);
and U23137 (N_23137,N_17466,N_15053);
nor U23138 (N_23138,N_18294,N_16419);
xnor U23139 (N_23139,N_15946,N_16979);
or U23140 (N_23140,N_19947,N_17558);
nor U23141 (N_23141,N_16001,N_15237);
nand U23142 (N_23142,N_19590,N_19477);
xnor U23143 (N_23143,N_16123,N_15597);
and U23144 (N_23144,N_17044,N_18123);
nand U23145 (N_23145,N_18688,N_18383);
xor U23146 (N_23146,N_16233,N_15690);
and U23147 (N_23147,N_18477,N_17665);
or U23148 (N_23148,N_17561,N_17794);
nor U23149 (N_23149,N_17290,N_16588);
nor U23150 (N_23150,N_17958,N_17767);
and U23151 (N_23151,N_17537,N_16421);
xnor U23152 (N_23152,N_16214,N_18738);
xor U23153 (N_23153,N_17293,N_17558);
xnor U23154 (N_23154,N_18173,N_18417);
or U23155 (N_23155,N_19127,N_19812);
and U23156 (N_23156,N_15859,N_17795);
nor U23157 (N_23157,N_19682,N_16546);
xor U23158 (N_23158,N_15033,N_19072);
nand U23159 (N_23159,N_15553,N_18381);
xnor U23160 (N_23160,N_18305,N_19052);
and U23161 (N_23161,N_17826,N_17466);
or U23162 (N_23162,N_19516,N_19103);
xor U23163 (N_23163,N_15282,N_15057);
or U23164 (N_23164,N_15553,N_19760);
xnor U23165 (N_23165,N_17804,N_16367);
xor U23166 (N_23166,N_17055,N_18922);
xor U23167 (N_23167,N_15043,N_16722);
or U23168 (N_23168,N_16461,N_19994);
and U23169 (N_23169,N_19500,N_19010);
or U23170 (N_23170,N_18074,N_19381);
xnor U23171 (N_23171,N_19304,N_16934);
or U23172 (N_23172,N_16146,N_15093);
and U23173 (N_23173,N_15330,N_19251);
nand U23174 (N_23174,N_17407,N_17990);
xnor U23175 (N_23175,N_17647,N_16270);
xor U23176 (N_23176,N_18113,N_19940);
nand U23177 (N_23177,N_17037,N_19139);
or U23178 (N_23178,N_18686,N_16722);
nor U23179 (N_23179,N_15927,N_15253);
xnor U23180 (N_23180,N_18461,N_15345);
and U23181 (N_23181,N_18123,N_18485);
nand U23182 (N_23182,N_18698,N_18326);
nor U23183 (N_23183,N_16481,N_15748);
nand U23184 (N_23184,N_15712,N_16986);
or U23185 (N_23185,N_19757,N_19482);
xnor U23186 (N_23186,N_17443,N_18416);
xor U23187 (N_23187,N_16698,N_16071);
nand U23188 (N_23188,N_15711,N_19189);
and U23189 (N_23189,N_15980,N_15470);
or U23190 (N_23190,N_15232,N_18694);
or U23191 (N_23191,N_19112,N_18950);
xor U23192 (N_23192,N_18291,N_17100);
nand U23193 (N_23193,N_19175,N_17070);
and U23194 (N_23194,N_16000,N_19965);
and U23195 (N_23195,N_17464,N_16699);
nor U23196 (N_23196,N_15306,N_18912);
or U23197 (N_23197,N_15655,N_17540);
and U23198 (N_23198,N_17476,N_17296);
or U23199 (N_23199,N_19651,N_19188);
nor U23200 (N_23200,N_19073,N_15484);
and U23201 (N_23201,N_19976,N_15182);
and U23202 (N_23202,N_19772,N_17604);
and U23203 (N_23203,N_15355,N_17896);
nand U23204 (N_23204,N_19327,N_17354);
or U23205 (N_23205,N_18049,N_17481);
nand U23206 (N_23206,N_15384,N_19526);
and U23207 (N_23207,N_19816,N_18350);
and U23208 (N_23208,N_18007,N_19335);
nor U23209 (N_23209,N_15027,N_15746);
xor U23210 (N_23210,N_17764,N_16531);
nor U23211 (N_23211,N_15528,N_16066);
xnor U23212 (N_23212,N_18252,N_18937);
nand U23213 (N_23213,N_16215,N_17705);
or U23214 (N_23214,N_17704,N_15935);
nor U23215 (N_23215,N_16262,N_18005);
or U23216 (N_23216,N_19883,N_18295);
nor U23217 (N_23217,N_19421,N_17533);
and U23218 (N_23218,N_15811,N_17398);
xor U23219 (N_23219,N_18393,N_16464);
and U23220 (N_23220,N_17370,N_17420);
and U23221 (N_23221,N_18960,N_16656);
nand U23222 (N_23222,N_18804,N_18327);
xnor U23223 (N_23223,N_19858,N_15602);
nand U23224 (N_23224,N_19286,N_18351);
xor U23225 (N_23225,N_16524,N_15591);
nand U23226 (N_23226,N_17561,N_16130);
nor U23227 (N_23227,N_15251,N_17654);
nor U23228 (N_23228,N_16859,N_18704);
nor U23229 (N_23229,N_17803,N_15939);
nor U23230 (N_23230,N_16961,N_15844);
or U23231 (N_23231,N_15560,N_15624);
xnor U23232 (N_23232,N_16887,N_15664);
or U23233 (N_23233,N_16341,N_16707);
nand U23234 (N_23234,N_18140,N_18839);
and U23235 (N_23235,N_19713,N_16173);
xnor U23236 (N_23236,N_15287,N_15134);
or U23237 (N_23237,N_18740,N_19400);
xnor U23238 (N_23238,N_16111,N_18001);
and U23239 (N_23239,N_18956,N_16807);
nor U23240 (N_23240,N_16218,N_15764);
or U23241 (N_23241,N_15249,N_17850);
nand U23242 (N_23242,N_18440,N_18458);
nand U23243 (N_23243,N_15084,N_17070);
nor U23244 (N_23244,N_15359,N_18421);
xor U23245 (N_23245,N_18466,N_19527);
or U23246 (N_23246,N_16871,N_17147);
nor U23247 (N_23247,N_15386,N_19602);
nand U23248 (N_23248,N_18982,N_19776);
xor U23249 (N_23249,N_16123,N_19467);
nor U23250 (N_23250,N_16360,N_18991);
and U23251 (N_23251,N_18672,N_16359);
and U23252 (N_23252,N_19557,N_16128);
or U23253 (N_23253,N_16727,N_18246);
nand U23254 (N_23254,N_15258,N_17352);
xor U23255 (N_23255,N_16816,N_17849);
or U23256 (N_23256,N_19979,N_18246);
nor U23257 (N_23257,N_15401,N_16241);
or U23258 (N_23258,N_18660,N_16291);
nand U23259 (N_23259,N_15742,N_17664);
or U23260 (N_23260,N_18746,N_16407);
or U23261 (N_23261,N_17126,N_16627);
nand U23262 (N_23262,N_19199,N_16323);
and U23263 (N_23263,N_17377,N_18630);
xnor U23264 (N_23264,N_15111,N_18402);
or U23265 (N_23265,N_16591,N_16982);
nor U23266 (N_23266,N_17989,N_15643);
xor U23267 (N_23267,N_18825,N_19470);
and U23268 (N_23268,N_16650,N_17433);
and U23269 (N_23269,N_18807,N_17689);
or U23270 (N_23270,N_15812,N_17778);
xor U23271 (N_23271,N_16879,N_18721);
or U23272 (N_23272,N_15822,N_16450);
or U23273 (N_23273,N_18607,N_18066);
or U23274 (N_23274,N_15918,N_16566);
xor U23275 (N_23275,N_16606,N_16214);
and U23276 (N_23276,N_18150,N_17364);
or U23277 (N_23277,N_19069,N_17527);
or U23278 (N_23278,N_17108,N_19036);
nor U23279 (N_23279,N_19303,N_15176);
nand U23280 (N_23280,N_15235,N_17569);
nor U23281 (N_23281,N_18696,N_17389);
nor U23282 (N_23282,N_16839,N_16478);
nor U23283 (N_23283,N_19472,N_15495);
nor U23284 (N_23284,N_17396,N_19864);
nor U23285 (N_23285,N_16134,N_16408);
and U23286 (N_23286,N_17484,N_16191);
xor U23287 (N_23287,N_18422,N_16998);
or U23288 (N_23288,N_19496,N_16821);
xor U23289 (N_23289,N_15961,N_16761);
xnor U23290 (N_23290,N_16599,N_18666);
nor U23291 (N_23291,N_16991,N_17061);
or U23292 (N_23292,N_19826,N_18488);
and U23293 (N_23293,N_16779,N_15257);
nor U23294 (N_23294,N_17813,N_18603);
or U23295 (N_23295,N_17060,N_18980);
or U23296 (N_23296,N_15538,N_15831);
or U23297 (N_23297,N_16507,N_15136);
and U23298 (N_23298,N_16214,N_18571);
xnor U23299 (N_23299,N_16461,N_16115);
nor U23300 (N_23300,N_15172,N_19213);
or U23301 (N_23301,N_19056,N_17526);
nor U23302 (N_23302,N_19159,N_18908);
xnor U23303 (N_23303,N_17765,N_15321);
nor U23304 (N_23304,N_18696,N_18962);
nand U23305 (N_23305,N_18383,N_18580);
or U23306 (N_23306,N_15729,N_16018);
or U23307 (N_23307,N_18260,N_17434);
and U23308 (N_23308,N_18565,N_17114);
and U23309 (N_23309,N_17458,N_15488);
nand U23310 (N_23310,N_18021,N_17684);
nor U23311 (N_23311,N_15183,N_15293);
nand U23312 (N_23312,N_18774,N_18177);
or U23313 (N_23313,N_18879,N_15253);
nor U23314 (N_23314,N_17335,N_16959);
xnor U23315 (N_23315,N_19054,N_19100);
xor U23316 (N_23316,N_19095,N_15669);
nand U23317 (N_23317,N_15198,N_18627);
and U23318 (N_23318,N_15267,N_16877);
nand U23319 (N_23319,N_19356,N_16095);
or U23320 (N_23320,N_17156,N_18040);
nand U23321 (N_23321,N_18281,N_19540);
xnor U23322 (N_23322,N_19134,N_19871);
nand U23323 (N_23323,N_17219,N_17082);
and U23324 (N_23324,N_19382,N_16007);
xor U23325 (N_23325,N_18921,N_19125);
or U23326 (N_23326,N_19508,N_15671);
xor U23327 (N_23327,N_18981,N_16805);
or U23328 (N_23328,N_18401,N_15675);
and U23329 (N_23329,N_16745,N_16105);
and U23330 (N_23330,N_16428,N_17786);
or U23331 (N_23331,N_19098,N_19059);
nor U23332 (N_23332,N_18740,N_19694);
nor U23333 (N_23333,N_17375,N_18653);
nor U23334 (N_23334,N_17059,N_15937);
nor U23335 (N_23335,N_16766,N_17010);
xor U23336 (N_23336,N_18489,N_18165);
or U23337 (N_23337,N_19772,N_19723);
nor U23338 (N_23338,N_15897,N_15518);
and U23339 (N_23339,N_19823,N_18683);
and U23340 (N_23340,N_18175,N_16009);
nor U23341 (N_23341,N_15585,N_18421);
or U23342 (N_23342,N_19508,N_17654);
or U23343 (N_23343,N_18452,N_19891);
nand U23344 (N_23344,N_17448,N_15470);
and U23345 (N_23345,N_15707,N_16395);
or U23346 (N_23346,N_19026,N_15320);
and U23347 (N_23347,N_18826,N_16200);
nor U23348 (N_23348,N_16642,N_19295);
or U23349 (N_23349,N_15420,N_15124);
nor U23350 (N_23350,N_17064,N_19286);
nand U23351 (N_23351,N_15816,N_18275);
and U23352 (N_23352,N_17138,N_16999);
and U23353 (N_23353,N_15883,N_17653);
nand U23354 (N_23354,N_17274,N_18654);
nor U23355 (N_23355,N_15076,N_18421);
nor U23356 (N_23356,N_18036,N_15910);
and U23357 (N_23357,N_18349,N_19002);
and U23358 (N_23358,N_15794,N_17654);
nand U23359 (N_23359,N_16850,N_16647);
and U23360 (N_23360,N_17186,N_19092);
and U23361 (N_23361,N_19567,N_16803);
nor U23362 (N_23362,N_18836,N_17729);
or U23363 (N_23363,N_15634,N_17967);
and U23364 (N_23364,N_16334,N_18810);
xnor U23365 (N_23365,N_18502,N_19865);
xnor U23366 (N_23366,N_19560,N_15603);
and U23367 (N_23367,N_18721,N_19616);
or U23368 (N_23368,N_16601,N_18420);
and U23369 (N_23369,N_18485,N_18881);
or U23370 (N_23370,N_17956,N_17885);
nand U23371 (N_23371,N_15358,N_15422);
xnor U23372 (N_23372,N_19494,N_19780);
or U23373 (N_23373,N_17876,N_16076);
and U23374 (N_23374,N_16751,N_15096);
xor U23375 (N_23375,N_15007,N_17997);
nor U23376 (N_23376,N_15863,N_16913);
nor U23377 (N_23377,N_17990,N_17471);
and U23378 (N_23378,N_16064,N_17997);
nor U23379 (N_23379,N_19647,N_18620);
nor U23380 (N_23380,N_19527,N_18419);
or U23381 (N_23381,N_17293,N_19140);
and U23382 (N_23382,N_16176,N_18708);
xor U23383 (N_23383,N_19889,N_16510);
nor U23384 (N_23384,N_19736,N_19396);
or U23385 (N_23385,N_18363,N_15578);
nand U23386 (N_23386,N_17206,N_17260);
xnor U23387 (N_23387,N_19719,N_18298);
or U23388 (N_23388,N_19171,N_19513);
and U23389 (N_23389,N_19952,N_15361);
or U23390 (N_23390,N_17984,N_15748);
xor U23391 (N_23391,N_19790,N_18638);
nor U23392 (N_23392,N_16544,N_19608);
nor U23393 (N_23393,N_16404,N_15340);
nand U23394 (N_23394,N_15763,N_17063);
xnor U23395 (N_23395,N_16533,N_16823);
nor U23396 (N_23396,N_15427,N_18968);
and U23397 (N_23397,N_17759,N_18377);
nand U23398 (N_23398,N_15687,N_16167);
nand U23399 (N_23399,N_17365,N_18637);
nor U23400 (N_23400,N_16268,N_16188);
nor U23401 (N_23401,N_15127,N_17728);
xor U23402 (N_23402,N_15790,N_16410);
nand U23403 (N_23403,N_18786,N_15947);
or U23404 (N_23404,N_17102,N_19370);
xnor U23405 (N_23405,N_16518,N_17700);
nand U23406 (N_23406,N_15073,N_18895);
nand U23407 (N_23407,N_18988,N_18335);
and U23408 (N_23408,N_18774,N_18868);
and U23409 (N_23409,N_18032,N_19990);
or U23410 (N_23410,N_17568,N_15810);
nor U23411 (N_23411,N_16065,N_16074);
and U23412 (N_23412,N_18153,N_15296);
xnor U23413 (N_23413,N_17143,N_16556);
xnor U23414 (N_23414,N_19076,N_18262);
xnor U23415 (N_23415,N_15278,N_15609);
nor U23416 (N_23416,N_16826,N_19973);
nor U23417 (N_23417,N_19598,N_15292);
and U23418 (N_23418,N_19903,N_15450);
xor U23419 (N_23419,N_19366,N_15796);
xnor U23420 (N_23420,N_18562,N_18538);
nor U23421 (N_23421,N_16120,N_19267);
or U23422 (N_23422,N_16459,N_17572);
or U23423 (N_23423,N_16138,N_18305);
or U23424 (N_23424,N_19035,N_16029);
or U23425 (N_23425,N_17330,N_15256);
nor U23426 (N_23426,N_17303,N_15329);
nand U23427 (N_23427,N_15892,N_19569);
nand U23428 (N_23428,N_16411,N_16202);
or U23429 (N_23429,N_19424,N_15616);
or U23430 (N_23430,N_16031,N_19428);
nand U23431 (N_23431,N_17872,N_15731);
or U23432 (N_23432,N_17653,N_15368);
xnor U23433 (N_23433,N_18482,N_16179);
or U23434 (N_23434,N_19385,N_15207);
and U23435 (N_23435,N_18287,N_17672);
or U23436 (N_23436,N_17796,N_18403);
or U23437 (N_23437,N_16784,N_17892);
nand U23438 (N_23438,N_15742,N_15686);
xnor U23439 (N_23439,N_17976,N_15476);
xnor U23440 (N_23440,N_16462,N_17124);
nor U23441 (N_23441,N_17859,N_17514);
and U23442 (N_23442,N_18102,N_17998);
nor U23443 (N_23443,N_15343,N_15289);
nor U23444 (N_23444,N_18338,N_19672);
nor U23445 (N_23445,N_19260,N_17923);
nor U23446 (N_23446,N_19725,N_15675);
nor U23447 (N_23447,N_16834,N_16802);
or U23448 (N_23448,N_19874,N_18812);
xor U23449 (N_23449,N_15838,N_17488);
nand U23450 (N_23450,N_19886,N_19200);
nand U23451 (N_23451,N_16733,N_17461);
xor U23452 (N_23452,N_16743,N_15652);
and U23453 (N_23453,N_15945,N_19094);
or U23454 (N_23454,N_19022,N_17380);
or U23455 (N_23455,N_16174,N_15911);
and U23456 (N_23456,N_18397,N_16812);
xnor U23457 (N_23457,N_15517,N_16460);
nor U23458 (N_23458,N_15249,N_19848);
nand U23459 (N_23459,N_16035,N_17426);
nand U23460 (N_23460,N_19760,N_19267);
nor U23461 (N_23461,N_16264,N_18606);
xnor U23462 (N_23462,N_16191,N_18826);
nand U23463 (N_23463,N_16622,N_19260);
nor U23464 (N_23464,N_19726,N_19694);
or U23465 (N_23465,N_18265,N_16753);
and U23466 (N_23466,N_16766,N_15701);
or U23467 (N_23467,N_18861,N_15546);
nor U23468 (N_23468,N_16712,N_18340);
xor U23469 (N_23469,N_16744,N_16569);
and U23470 (N_23470,N_16549,N_19053);
nor U23471 (N_23471,N_16579,N_18032);
nand U23472 (N_23472,N_16675,N_17780);
and U23473 (N_23473,N_19000,N_19208);
xnor U23474 (N_23474,N_17628,N_16973);
nand U23475 (N_23475,N_15732,N_17815);
xnor U23476 (N_23476,N_18108,N_17129);
xor U23477 (N_23477,N_16176,N_17842);
nor U23478 (N_23478,N_18951,N_18369);
nand U23479 (N_23479,N_15085,N_16307);
nand U23480 (N_23480,N_18964,N_19289);
and U23481 (N_23481,N_15075,N_17550);
and U23482 (N_23482,N_15726,N_15354);
or U23483 (N_23483,N_15041,N_16910);
and U23484 (N_23484,N_17493,N_19348);
nand U23485 (N_23485,N_17396,N_19112);
xor U23486 (N_23486,N_18891,N_15573);
nand U23487 (N_23487,N_15382,N_17191);
nand U23488 (N_23488,N_16909,N_15254);
xnor U23489 (N_23489,N_18917,N_17567);
and U23490 (N_23490,N_15738,N_16097);
nor U23491 (N_23491,N_15601,N_15127);
or U23492 (N_23492,N_16461,N_16662);
or U23493 (N_23493,N_18361,N_16431);
nor U23494 (N_23494,N_17285,N_19601);
nor U23495 (N_23495,N_19913,N_15709);
nand U23496 (N_23496,N_18538,N_18805);
and U23497 (N_23497,N_15421,N_16661);
nand U23498 (N_23498,N_19859,N_18202);
and U23499 (N_23499,N_17388,N_15568);
xnor U23500 (N_23500,N_15576,N_18733);
and U23501 (N_23501,N_18411,N_17604);
xor U23502 (N_23502,N_19756,N_19148);
or U23503 (N_23503,N_19086,N_17172);
or U23504 (N_23504,N_17981,N_17903);
or U23505 (N_23505,N_17276,N_17802);
and U23506 (N_23506,N_16601,N_18427);
nand U23507 (N_23507,N_19200,N_17504);
and U23508 (N_23508,N_15874,N_18457);
xnor U23509 (N_23509,N_17038,N_18284);
xnor U23510 (N_23510,N_19965,N_18240);
nand U23511 (N_23511,N_18778,N_17028);
nand U23512 (N_23512,N_15905,N_17151);
xor U23513 (N_23513,N_18339,N_16652);
nand U23514 (N_23514,N_19421,N_19868);
or U23515 (N_23515,N_17437,N_16791);
and U23516 (N_23516,N_19306,N_15637);
xor U23517 (N_23517,N_17957,N_15151);
nor U23518 (N_23518,N_18398,N_19563);
nand U23519 (N_23519,N_15701,N_17473);
and U23520 (N_23520,N_16300,N_15065);
and U23521 (N_23521,N_15947,N_18090);
nor U23522 (N_23522,N_17631,N_18693);
nor U23523 (N_23523,N_15827,N_16787);
and U23524 (N_23524,N_18237,N_15505);
and U23525 (N_23525,N_19246,N_17574);
nor U23526 (N_23526,N_17560,N_17382);
xor U23527 (N_23527,N_18027,N_17329);
and U23528 (N_23528,N_16888,N_16971);
or U23529 (N_23529,N_15350,N_15973);
nor U23530 (N_23530,N_19068,N_16765);
xor U23531 (N_23531,N_16502,N_15103);
nand U23532 (N_23532,N_19262,N_15055);
xnor U23533 (N_23533,N_19336,N_19511);
nor U23534 (N_23534,N_18902,N_19101);
or U23535 (N_23535,N_17771,N_19729);
or U23536 (N_23536,N_15548,N_16620);
and U23537 (N_23537,N_17667,N_19653);
nand U23538 (N_23538,N_15580,N_18129);
xnor U23539 (N_23539,N_17290,N_19010);
xnor U23540 (N_23540,N_17105,N_16941);
nand U23541 (N_23541,N_17528,N_17847);
or U23542 (N_23542,N_19300,N_18206);
xor U23543 (N_23543,N_15582,N_15424);
nor U23544 (N_23544,N_15130,N_17769);
or U23545 (N_23545,N_19437,N_19974);
nand U23546 (N_23546,N_17931,N_18331);
and U23547 (N_23547,N_15809,N_15792);
or U23548 (N_23548,N_17863,N_18441);
or U23549 (N_23549,N_18866,N_17353);
and U23550 (N_23550,N_16624,N_18047);
or U23551 (N_23551,N_17349,N_15617);
or U23552 (N_23552,N_17226,N_18185);
xor U23553 (N_23553,N_16608,N_19671);
or U23554 (N_23554,N_18600,N_15856);
nor U23555 (N_23555,N_16955,N_15947);
and U23556 (N_23556,N_15671,N_16965);
nand U23557 (N_23557,N_17625,N_16928);
and U23558 (N_23558,N_16398,N_18601);
nor U23559 (N_23559,N_18502,N_18004);
xor U23560 (N_23560,N_18708,N_18579);
xnor U23561 (N_23561,N_16897,N_19727);
xnor U23562 (N_23562,N_16443,N_15384);
or U23563 (N_23563,N_16756,N_18477);
nor U23564 (N_23564,N_16642,N_18794);
or U23565 (N_23565,N_19187,N_15634);
nand U23566 (N_23566,N_17779,N_19488);
xor U23567 (N_23567,N_17492,N_16066);
nor U23568 (N_23568,N_15598,N_19363);
nor U23569 (N_23569,N_15982,N_16571);
nand U23570 (N_23570,N_16712,N_17148);
and U23571 (N_23571,N_17596,N_15934);
and U23572 (N_23572,N_18040,N_18942);
nand U23573 (N_23573,N_18047,N_17687);
nor U23574 (N_23574,N_18537,N_18226);
nand U23575 (N_23575,N_16711,N_17630);
xor U23576 (N_23576,N_18935,N_17850);
nand U23577 (N_23577,N_18034,N_15331);
and U23578 (N_23578,N_15725,N_15421);
nand U23579 (N_23579,N_16650,N_19757);
xor U23580 (N_23580,N_19675,N_16048);
nand U23581 (N_23581,N_18584,N_15369);
and U23582 (N_23582,N_18716,N_15636);
xor U23583 (N_23583,N_16651,N_16831);
nor U23584 (N_23584,N_19351,N_19215);
and U23585 (N_23585,N_16262,N_18158);
nor U23586 (N_23586,N_19831,N_18753);
nand U23587 (N_23587,N_16397,N_16056);
nand U23588 (N_23588,N_17136,N_19257);
and U23589 (N_23589,N_15001,N_18523);
nand U23590 (N_23590,N_19689,N_16565);
nor U23591 (N_23591,N_16767,N_15416);
xor U23592 (N_23592,N_18581,N_15507);
or U23593 (N_23593,N_18445,N_19139);
or U23594 (N_23594,N_15218,N_15262);
xnor U23595 (N_23595,N_15815,N_19315);
and U23596 (N_23596,N_16351,N_17487);
and U23597 (N_23597,N_16769,N_16286);
nand U23598 (N_23598,N_19045,N_17835);
or U23599 (N_23599,N_18786,N_15763);
and U23600 (N_23600,N_16709,N_18482);
or U23601 (N_23601,N_18050,N_16103);
xor U23602 (N_23602,N_18361,N_15837);
xor U23603 (N_23603,N_18289,N_19387);
or U23604 (N_23604,N_19294,N_15155);
nor U23605 (N_23605,N_17187,N_19140);
nor U23606 (N_23606,N_18593,N_15944);
nand U23607 (N_23607,N_15303,N_16986);
and U23608 (N_23608,N_18650,N_19746);
xor U23609 (N_23609,N_18355,N_18566);
and U23610 (N_23610,N_15408,N_17693);
or U23611 (N_23611,N_17355,N_18565);
xnor U23612 (N_23612,N_19752,N_17333);
and U23613 (N_23613,N_15571,N_17681);
or U23614 (N_23614,N_17817,N_16846);
or U23615 (N_23615,N_15498,N_16262);
or U23616 (N_23616,N_17716,N_18221);
and U23617 (N_23617,N_19299,N_17050);
and U23618 (N_23618,N_18834,N_16885);
or U23619 (N_23619,N_15042,N_17224);
or U23620 (N_23620,N_16289,N_16150);
nor U23621 (N_23621,N_15458,N_15776);
and U23622 (N_23622,N_15514,N_18483);
nand U23623 (N_23623,N_17171,N_19799);
nor U23624 (N_23624,N_19368,N_17850);
or U23625 (N_23625,N_19150,N_16629);
and U23626 (N_23626,N_17832,N_17487);
xnor U23627 (N_23627,N_18396,N_19500);
xor U23628 (N_23628,N_16915,N_19649);
nand U23629 (N_23629,N_18692,N_16911);
and U23630 (N_23630,N_15049,N_19393);
nand U23631 (N_23631,N_18848,N_16499);
or U23632 (N_23632,N_16285,N_19747);
or U23633 (N_23633,N_19845,N_17542);
or U23634 (N_23634,N_17498,N_15298);
nand U23635 (N_23635,N_15365,N_19249);
nor U23636 (N_23636,N_16044,N_16636);
nand U23637 (N_23637,N_16005,N_19771);
and U23638 (N_23638,N_19580,N_16797);
and U23639 (N_23639,N_18575,N_17393);
nor U23640 (N_23640,N_17746,N_18009);
and U23641 (N_23641,N_16799,N_17456);
or U23642 (N_23642,N_16662,N_19730);
and U23643 (N_23643,N_16942,N_15836);
nor U23644 (N_23644,N_15000,N_17860);
xnor U23645 (N_23645,N_19864,N_15902);
xnor U23646 (N_23646,N_18912,N_18111);
xor U23647 (N_23647,N_17393,N_15844);
nand U23648 (N_23648,N_17190,N_17894);
and U23649 (N_23649,N_17122,N_16346);
or U23650 (N_23650,N_15566,N_17255);
nand U23651 (N_23651,N_16533,N_18485);
nor U23652 (N_23652,N_16348,N_17257);
nand U23653 (N_23653,N_19803,N_17857);
xor U23654 (N_23654,N_15499,N_17837);
nor U23655 (N_23655,N_16993,N_19885);
and U23656 (N_23656,N_17662,N_18705);
or U23657 (N_23657,N_15343,N_18591);
or U23658 (N_23658,N_19939,N_18738);
or U23659 (N_23659,N_15417,N_15288);
or U23660 (N_23660,N_17646,N_17521);
and U23661 (N_23661,N_16813,N_18438);
xor U23662 (N_23662,N_17633,N_17716);
or U23663 (N_23663,N_19858,N_15161);
xnor U23664 (N_23664,N_16550,N_15924);
nand U23665 (N_23665,N_18994,N_16159);
or U23666 (N_23666,N_15361,N_16893);
nand U23667 (N_23667,N_19526,N_19116);
nand U23668 (N_23668,N_19526,N_16748);
nand U23669 (N_23669,N_15955,N_16598);
nor U23670 (N_23670,N_16985,N_18338);
nand U23671 (N_23671,N_17203,N_16281);
nand U23672 (N_23672,N_19532,N_19180);
or U23673 (N_23673,N_16682,N_15367);
nand U23674 (N_23674,N_15973,N_16610);
nand U23675 (N_23675,N_17555,N_17447);
or U23676 (N_23676,N_15501,N_18749);
nand U23677 (N_23677,N_16860,N_16978);
or U23678 (N_23678,N_15597,N_19243);
nor U23679 (N_23679,N_15800,N_18258);
nor U23680 (N_23680,N_17442,N_18192);
or U23681 (N_23681,N_18788,N_15169);
nor U23682 (N_23682,N_16414,N_18635);
nand U23683 (N_23683,N_15506,N_18964);
xnor U23684 (N_23684,N_19110,N_17291);
nand U23685 (N_23685,N_15303,N_19896);
xor U23686 (N_23686,N_17615,N_15583);
nand U23687 (N_23687,N_17753,N_17379);
nand U23688 (N_23688,N_17227,N_16391);
or U23689 (N_23689,N_17362,N_15214);
nand U23690 (N_23690,N_16613,N_17630);
xnor U23691 (N_23691,N_18440,N_17041);
xnor U23692 (N_23692,N_16402,N_15705);
nor U23693 (N_23693,N_18902,N_16441);
and U23694 (N_23694,N_17445,N_17850);
nor U23695 (N_23695,N_17039,N_19165);
and U23696 (N_23696,N_18336,N_15964);
nor U23697 (N_23697,N_15321,N_16033);
xor U23698 (N_23698,N_15715,N_18931);
and U23699 (N_23699,N_16265,N_19441);
or U23700 (N_23700,N_16753,N_15490);
nand U23701 (N_23701,N_15903,N_18192);
nor U23702 (N_23702,N_17125,N_18195);
nand U23703 (N_23703,N_17669,N_15379);
and U23704 (N_23704,N_15510,N_15315);
nor U23705 (N_23705,N_18217,N_16803);
or U23706 (N_23706,N_17966,N_18479);
nor U23707 (N_23707,N_15955,N_17750);
nor U23708 (N_23708,N_16941,N_17988);
and U23709 (N_23709,N_19183,N_19950);
nand U23710 (N_23710,N_18855,N_16622);
and U23711 (N_23711,N_18738,N_19349);
and U23712 (N_23712,N_17320,N_15939);
or U23713 (N_23713,N_17870,N_17279);
xor U23714 (N_23714,N_18436,N_16406);
xnor U23715 (N_23715,N_16871,N_15726);
or U23716 (N_23716,N_19866,N_15371);
xnor U23717 (N_23717,N_16554,N_19039);
nand U23718 (N_23718,N_17724,N_16203);
or U23719 (N_23719,N_19838,N_16778);
xnor U23720 (N_23720,N_15091,N_15867);
or U23721 (N_23721,N_19715,N_16688);
nor U23722 (N_23722,N_17533,N_18394);
and U23723 (N_23723,N_17980,N_19869);
and U23724 (N_23724,N_18699,N_18108);
nor U23725 (N_23725,N_15273,N_18923);
or U23726 (N_23726,N_17428,N_18894);
nor U23727 (N_23727,N_16994,N_17950);
nor U23728 (N_23728,N_17727,N_15803);
xor U23729 (N_23729,N_19889,N_19098);
and U23730 (N_23730,N_16059,N_19022);
or U23731 (N_23731,N_15537,N_15695);
nor U23732 (N_23732,N_18665,N_17583);
nor U23733 (N_23733,N_16952,N_16365);
and U23734 (N_23734,N_18719,N_16369);
nand U23735 (N_23735,N_18646,N_15833);
or U23736 (N_23736,N_15407,N_17132);
nand U23737 (N_23737,N_19811,N_15815);
nor U23738 (N_23738,N_15264,N_16257);
nand U23739 (N_23739,N_17070,N_16417);
and U23740 (N_23740,N_15035,N_18727);
and U23741 (N_23741,N_17781,N_18994);
or U23742 (N_23742,N_18952,N_15846);
or U23743 (N_23743,N_17131,N_19188);
xnor U23744 (N_23744,N_16585,N_15507);
and U23745 (N_23745,N_18426,N_15450);
nor U23746 (N_23746,N_15271,N_15831);
xnor U23747 (N_23747,N_15180,N_17307);
nand U23748 (N_23748,N_16961,N_18932);
and U23749 (N_23749,N_18970,N_15488);
and U23750 (N_23750,N_17080,N_18077);
xor U23751 (N_23751,N_18162,N_18066);
nand U23752 (N_23752,N_18007,N_18917);
xnor U23753 (N_23753,N_16297,N_15463);
nand U23754 (N_23754,N_19193,N_19682);
or U23755 (N_23755,N_16072,N_18328);
nor U23756 (N_23756,N_16966,N_16414);
and U23757 (N_23757,N_15580,N_19963);
nand U23758 (N_23758,N_19075,N_16012);
nand U23759 (N_23759,N_18461,N_16412);
and U23760 (N_23760,N_17761,N_17337);
xnor U23761 (N_23761,N_17406,N_18667);
xnor U23762 (N_23762,N_17792,N_19267);
xor U23763 (N_23763,N_18814,N_17484);
and U23764 (N_23764,N_17520,N_19006);
xor U23765 (N_23765,N_18567,N_17862);
and U23766 (N_23766,N_15616,N_15733);
and U23767 (N_23767,N_18745,N_18934);
nand U23768 (N_23768,N_15588,N_16811);
and U23769 (N_23769,N_16031,N_16724);
or U23770 (N_23770,N_16954,N_17320);
nand U23771 (N_23771,N_17861,N_19155);
or U23772 (N_23772,N_19596,N_19629);
or U23773 (N_23773,N_19947,N_17145);
nor U23774 (N_23774,N_15013,N_16798);
nor U23775 (N_23775,N_18268,N_18311);
or U23776 (N_23776,N_17724,N_19148);
or U23777 (N_23777,N_17519,N_19100);
and U23778 (N_23778,N_16618,N_16413);
nor U23779 (N_23779,N_19141,N_19553);
and U23780 (N_23780,N_15585,N_17595);
or U23781 (N_23781,N_15157,N_19853);
and U23782 (N_23782,N_18890,N_19173);
and U23783 (N_23783,N_17711,N_15935);
nor U23784 (N_23784,N_15541,N_19189);
and U23785 (N_23785,N_16266,N_15099);
nor U23786 (N_23786,N_19261,N_15694);
nand U23787 (N_23787,N_15379,N_15199);
nor U23788 (N_23788,N_17619,N_19023);
or U23789 (N_23789,N_18461,N_18609);
nor U23790 (N_23790,N_18339,N_15967);
nand U23791 (N_23791,N_16341,N_16062);
nor U23792 (N_23792,N_16347,N_18880);
nor U23793 (N_23793,N_16846,N_17447);
nand U23794 (N_23794,N_18776,N_18307);
nor U23795 (N_23795,N_19953,N_19281);
xor U23796 (N_23796,N_19136,N_19338);
nor U23797 (N_23797,N_19627,N_17255);
nor U23798 (N_23798,N_18113,N_17254);
or U23799 (N_23799,N_19147,N_19987);
nand U23800 (N_23800,N_15256,N_17466);
or U23801 (N_23801,N_18072,N_15929);
and U23802 (N_23802,N_18787,N_17406);
nor U23803 (N_23803,N_17507,N_16071);
and U23804 (N_23804,N_17408,N_15153);
nor U23805 (N_23805,N_15080,N_19780);
xor U23806 (N_23806,N_16719,N_15082);
or U23807 (N_23807,N_17900,N_19585);
nor U23808 (N_23808,N_16178,N_15766);
xor U23809 (N_23809,N_18396,N_17920);
nor U23810 (N_23810,N_19898,N_19032);
nor U23811 (N_23811,N_16586,N_15759);
nand U23812 (N_23812,N_18450,N_18193);
nor U23813 (N_23813,N_17077,N_15148);
nor U23814 (N_23814,N_18194,N_17841);
xnor U23815 (N_23815,N_16133,N_15177);
or U23816 (N_23816,N_16925,N_17589);
nand U23817 (N_23817,N_16741,N_18790);
or U23818 (N_23818,N_16497,N_17018);
nor U23819 (N_23819,N_16994,N_15450);
nand U23820 (N_23820,N_17773,N_16617);
nand U23821 (N_23821,N_17696,N_19442);
nand U23822 (N_23822,N_15212,N_19144);
xnor U23823 (N_23823,N_16975,N_15071);
or U23824 (N_23824,N_16517,N_18883);
nor U23825 (N_23825,N_18148,N_15922);
nor U23826 (N_23826,N_18711,N_16117);
or U23827 (N_23827,N_19800,N_17958);
nor U23828 (N_23828,N_19259,N_18952);
xnor U23829 (N_23829,N_18660,N_19084);
or U23830 (N_23830,N_17236,N_19733);
nor U23831 (N_23831,N_17414,N_15106);
nand U23832 (N_23832,N_15488,N_15840);
nand U23833 (N_23833,N_16321,N_17996);
nand U23834 (N_23834,N_15348,N_16450);
and U23835 (N_23835,N_15425,N_18114);
and U23836 (N_23836,N_19541,N_18963);
nand U23837 (N_23837,N_17462,N_19560);
or U23838 (N_23838,N_17079,N_18604);
xnor U23839 (N_23839,N_17874,N_19900);
nor U23840 (N_23840,N_17271,N_15633);
and U23841 (N_23841,N_19232,N_15467);
or U23842 (N_23842,N_19651,N_16638);
nor U23843 (N_23843,N_16070,N_17326);
xnor U23844 (N_23844,N_15592,N_16401);
nand U23845 (N_23845,N_16395,N_17191);
nor U23846 (N_23846,N_18277,N_15636);
nand U23847 (N_23847,N_18477,N_17401);
nor U23848 (N_23848,N_16223,N_17702);
and U23849 (N_23849,N_15419,N_15496);
and U23850 (N_23850,N_17665,N_18479);
or U23851 (N_23851,N_17134,N_15864);
nand U23852 (N_23852,N_18447,N_18621);
and U23853 (N_23853,N_18905,N_19919);
and U23854 (N_23854,N_15282,N_16740);
and U23855 (N_23855,N_16416,N_15564);
or U23856 (N_23856,N_19828,N_18009);
nand U23857 (N_23857,N_16982,N_19701);
xor U23858 (N_23858,N_18106,N_16933);
or U23859 (N_23859,N_18327,N_19636);
and U23860 (N_23860,N_16038,N_15074);
xnor U23861 (N_23861,N_18859,N_17836);
nand U23862 (N_23862,N_15262,N_16793);
xor U23863 (N_23863,N_18137,N_15848);
and U23864 (N_23864,N_17926,N_15383);
and U23865 (N_23865,N_19068,N_19698);
xnor U23866 (N_23866,N_15684,N_17624);
xnor U23867 (N_23867,N_18557,N_16209);
nand U23868 (N_23868,N_17658,N_19662);
nor U23869 (N_23869,N_18676,N_15605);
or U23870 (N_23870,N_19331,N_18704);
nor U23871 (N_23871,N_19319,N_15930);
nand U23872 (N_23872,N_17387,N_19009);
or U23873 (N_23873,N_17852,N_16119);
or U23874 (N_23874,N_18889,N_18649);
and U23875 (N_23875,N_17446,N_16326);
or U23876 (N_23876,N_19758,N_19707);
or U23877 (N_23877,N_15749,N_19897);
or U23878 (N_23878,N_17437,N_19746);
nand U23879 (N_23879,N_15767,N_15280);
nor U23880 (N_23880,N_19415,N_19204);
or U23881 (N_23881,N_19150,N_16293);
or U23882 (N_23882,N_17540,N_18258);
and U23883 (N_23883,N_19975,N_18011);
nor U23884 (N_23884,N_18440,N_18170);
xor U23885 (N_23885,N_18954,N_18673);
xnor U23886 (N_23886,N_18748,N_18621);
or U23887 (N_23887,N_15031,N_19197);
or U23888 (N_23888,N_15132,N_19237);
nor U23889 (N_23889,N_16544,N_18360);
or U23890 (N_23890,N_19361,N_15571);
nand U23891 (N_23891,N_15241,N_18975);
or U23892 (N_23892,N_15085,N_18113);
nand U23893 (N_23893,N_17109,N_16982);
nand U23894 (N_23894,N_18361,N_17917);
xor U23895 (N_23895,N_19542,N_17840);
xor U23896 (N_23896,N_19685,N_17114);
nand U23897 (N_23897,N_18970,N_18615);
xnor U23898 (N_23898,N_16144,N_16486);
xor U23899 (N_23899,N_15734,N_15243);
or U23900 (N_23900,N_17753,N_18384);
xor U23901 (N_23901,N_19987,N_16503);
or U23902 (N_23902,N_18798,N_18510);
or U23903 (N_23903,N_15138,N_16136);
nor U23904 (N_23904,N_16621,N_17582);
and U23905 (N_23905,N_17578,N_18700);
nor U23906 (N_23906,N_18607,N_16567);
or U23907 (N_23907,N_15723,N_19098);
and U23908 (N_23908,N_19012,N_16305);
nand U23909 (N_23909,N_18964,N_19106);
and U23910 (N_23910,N_15829,N_18566);
xnor U23911 (N_23911,N_18971,N_19403);
xor U23912 (N_23912,N_18911,N_19242);
nand U23913 (N_23913,N_18458,N_15736);
or U23914 (N_23914,N_15512,N_19863);
xor U23915 (N_23915,N_17399,N_15468);
or U23916 (N_23916,N_16452,N_17491);
or U23917 (N_23917,N_16037,N_15200);
or U23918 (N_23918,N_17777,N_19505);
xor U23919 (N_23919,N_16603,N_19825);
or U23920 (N_23920,N_17723,N_18115);
nor U23921 (N_23921,N_16507,N_18150);
xnor U23922 (N_23922,N_15263,N_17683);
nor U23923 (N_23923,N_17437,N_17236);
or U23924 (N_23924,N_15113,N_18264);
nor U23925 (N_23925,N_15714,N_15373);
nand U23926 (N_23926,N_16100,N_19564);
xnor U23927 (N_23927,N_18946,N_16540);
xor U23928 (N_23928,N_19901,N_15496);
or U23929 (N_23929,N_17412,N_17175);
xnor U23930 (N_23930,N_15563,N_15884);
nand U23931 (N_23931,N_16071,N_18400);
xor U23932 (N_23932,N_15848,N_18791);
and U23933 (N_23933,N_18937,N_18591);
nor U23934 (N_23934,N_17840,N_16244);
nor U23935 (N_23935,N_16624,N_19747);
xor U23936 (N_23936,N_18187,N_16772);
xnor U23937 (N_23937,N_15872,N_17504);
or U23938 (N_23938,N_17711,N_16113);
or U23939 (N_23939,N_18568,N_19977);
nor U23940 (N_23940,N_17081,N_18294);
and U23941 (N_23941,N_16690,N_15296);
or U23942 (N_23942,N_18618,N_17841);
nor U23943 (N_23943,N_15088,N_18517);
and U23944 (N_23944,N_18108,N_19580);
nor U23945 (N_23945,N_16791,N_16048);
nor U23946 (N_23946,N_15717,N_18066);
xnor U23947 (N_23947,N_18541,N_17525);
nand U23948 (N_23948,N_16211,N_17151);
or U23949 (N_23949,N_15551,N_19126);
nor U23950 (N_23950,N_15873,N_19953);
or U23951 (N_23951,N_15883,N_19519);
and U23952 (N_23952,N_16159,N_19941);
xnor U23953 (N_23953,N_16811,N_19898);
nor U23954 (N_23954,N_15978,N_17970);
and U23955 (N_23955,N_16473,N_16795);
and U23956 (N_23956,N_19404,N_19088);
xor U23957 (N_23957,N_16276,N_16645);
xor U23958 (N_23958,N_15540,N_18675);
or U23959 (N_23959,N_19700,N_19019);
xor U23960 (N_23960,N_19769,N_17767);
or U23961 (N_23961,N_15646,N_19338);
nand U23962 (N_23962,N_16904,N_18613);
nand U23963 (N_23963,N_15924,N_16251);
nand U23964 (N_23964,N_16041,N_15569);
nor U23965 (N_23965,N_17351,N_18866);
nand U23966 (N_23966,N_17942,N_19009);
and U23967 (N_23967,N_18126,N_16769);
or U23968 (N_23968,N_15710,N_15265);
or U23969 (N_23969,N_16468,N_18487);
nor U23970 (N_23970,N_17844,N_19919);
nand U23971 (N_23971,N_17801,N_17833);
xor U23972 (N_23972,N_18143,N_16348);
xor U23973 (N_23973,N_17518,N_18450);
or U23974 (N_23974,N_18479,N_15220);
xnor U23975 (N_23975,N_18021,N_18380);
nor U23976 (N_23976,N_18913,N_15464);
xor U23977 (N_23977,N_15561,N_18265);
or U23978 (N_23978,N_18110,N_18132);
and U23979 (N_23979,N_15433,N_18960);
nor U23980 (N_23980,N_18195,N_15670);
or U23981 (N_23981,N_17690,N_18430);
nand U23982 (N_23982,N_16606,N_19772);
and U23983 (N_23983,N_18794,N_17705);
or U23984 (N_23984,N_18428,N_15852);
xnor U23985 (N_23985,N_15052,N_15828);
nor U23986 (N_23986,N_16897,N_18807);
or U23987 (N_23987,N_18024,N_18530);
nor U23988 (N_23988,N_15702,N_18430);
nand U23989 (N_23989,N_16983,N_15498);
xnor U23990 (N_23990,N_16749,N_17549);
nand U23991 (N_23991,N_16893,N_19912);
nand U23992 (N_23992,N_18525,N_15407);
nand U23993 (N_23993,N_15075,N_19720);
nand U23994 (N_23994,N_16852,N_15865);
nand U23995 (N_23995,N_17329,N_17075);
xnor U23996 (N_23996,N_17888,N_18741);
nor U23997 (N_23997,N_17872,N_18338);
nand U23998 (N_23998,N_16558,N_15594);
xnor U23999 (N_23999,N_15510,N_15514);
nand U24000 (N_24000,N_17581,N_19138);
xor U24001 (N_24001,N_18346,N_17095);
xor U24002 (N_24002,N_19910,N_16957);
nor U24003 (N_24003,N_17701,N_15847);
nor U24004 (N_24004,N_19359,N_17673);
or U24005 (N_24005,N_17611,N_18149);
or U24006 (N_24006,N_16029,N_17802);
nand U24007 (N_24007,N_19919,N_19149);
nand U24008 (N_24008,N_15701,N_19900);
and U24009 (N_24009,N_18549,N_18851);
or U24010 (N_24010,N_16321,N_15832);
nand U24011 (N_24011,N_15093,N_15726);
nor U24012 (N_24012,N_19014,N_15560);
nand U24013 (N_24013,N_19973,N_16377);
or U24014 (N_24014,N_16000,N_19649);
nor U24015 (N_24015,N_19338,N_18515);
nor U24016 (N_24016,N_19392,N_19246);
or U24017 (N_24017,N_16830,N_19469);
nor U24018 (N_24018,N_18332,N_18718);
nor U24019 (N_24019,N_16306,N_19027);
nor U24020 (N_24020,N_19707,N_17719);
nand U24021 (N_24021,N_15789,N_18064);
and U24022 (N_24022,N_19287,N_17611);
and U24023 (N_24023,N_19976,N_16181);
nor U24024 (N_24024,N_16552,N_18263);
nor U24025 (N_24025,N_18202,N_18782);
nand U24026 (N_24026,N_16119,N_15720);
nand U24027 (N_24027,N_16528,N_19017);
nand U24028 (N_24028,N_18878,N_15585);
or U24029 (N_24029,N_18450,N_19024);
nand U24030 (N_24030,N_19314,N_16633);
and U24031 (N_24031,N_19594,N_17761);
xor U24032 (N_24032,N_15704,N_19351);
xnor U24033 (N_24033,N_16153,N_16998);
nor U24034 (N_24034,N_17590,N_16262);
nand U24035 (N_24035,N_16733,N_19974);
or U24036 (N_24036,N_16646,N_15467);
and U24037 (N_24037,N_15199,N_16979);
nand U24038 (N_24038,N_19909,N_17532);
xnor U24039 (N_24039,N_15789,N_18218);
or U24040 (N_24040,N_19468,N_15072);
and U24041 (N_24041,N_18012,N_19691);
or U24042 (N_24042,N_17305,N_15701);
nor U24043 (N_24043,N_19150,N_18672);
nand U24044 (N_24044,N_17907,N_18614);
and U24045 (N_24045,N_19507,N_19595);
nand U24046 (N_24046,N_16252,N_19420);
nor U24047 (N_24047,N_17926,N_17665);
and U24048 (N_24048,N_15116,N_15893);
xor U24049 (N_24049,N_15344,N_18332);
nor U24050 (N_24050,N_18056,N_17852);
nand U24051 (N_24051,N_17385,N_18267);
nor U24052 (N_24052,N_18719,N_17386);
and U24053 (N_24053,N_16796,N_17594);
and U24054 (N_24054,N_15826,N_17953);
xor U24055 (N_24055,N_18752,N_18787);
or U24056 (N_24056,N_16879,N_18306);
and U24057 (N_24057,N_17126,N_17238);
nand U24058 (N_24058,N_18939,N_18354);
nor U24059 (N_24059,N_19212,N_16977);
or U24060 (N_24060,N_17552,N_15818);
xor U24061 (N_24061,N_19190,N_15864);
nor U24062 (N_24062,N_17957,N_17643);
nand U24063 (N_24063,N_15824,N_19633);
nor U24064 (N_24064,N_16333,N_15185);
nor U24065 (N_24065,N_16490,N_16501);
xnor U24066 (N_24066,N_16745,N_16989);
or U24067 (N_24067,N_18826,N_17691);
and U24068 (N_24068,N_15340,N_19891);
and U24069 (N_24069,N_19491,N_18367);
xnor U24070 (N_24070,N_17258,N_15291);
nand U24071 (N_24071,N_19681,N_16235);
and U24072 (N_24072,N_18335,N_15811);
nand U24073 (N_24073,N_18609,N_15121);
nor U24074 (N_24074,N_18714,N_15212);
xor U24075 (N_24075,N_16614,N_15765);
xnor U24076 (N_24076,N_17166,N_15771);
xor U24077 (N_24077,N_19883,N_17579);
and U24078 (N_24078,N_18513,N_19151);
nor U24079 (N_24079,N_17810,N_17401);
and U24080 (N_24080,N_15026,N_17869);
nand U24081 (N_24081,N_19562,N_18788);
nand U24082 (N_24082,N_15352,N_19259);
xor U24083 (N_24083,N_15613,N_18696);
or U24084 (N_24084,N_19824,N_18196);
and U24085 (N_24085,N_19385,N_17209);
xor U24086 (N_24086,N_15149,N_15733);
nor U24087 (N_24087,N_17149,N_17130);
nor U24088 (N_24088,N_16521,N_15519);
and U24089 (N_24089,N_16427,N_18854);
and U24090 (N_24090,N_17029,N_16798);
xor U24091 (N_24091,N_16984,N_15928);
xnor U24092 (N_24092,N_19762,N_16518);
nand U24093 (N_24093,N_17888,N_17835);
and U24094 (N_24094,N_17974,N_15415);
xnor U24095 (N_24095,N_18021,N_17215);
xor U24096 (N_24096,N_18335,N_17332);
nor U24097 (N_24097,N_15162,N_17314);
nand U24098 (N_24098,N_15572,N_18117);
nor U24099 (N_24099,N_18405,N_16781);
nor U24100 (N_24100,N_15174,N_17933);
and U24101 (N_24101,N_19665,N_17718);
or U24102 (N_24102,N_18582,N_17177);
nor U24103 (N_24103,N_15147,N_16000);
xor U24104 (N_24104,N_15475,N_15113);
xnor U24105 (N_24105,N_19107,N_18317);
nand U24106 (N_24106,N_15222,N_18766);
nand U24107 (N_24107,N_17286,N_15423);
or U24108 (N_24108,N_17407,N_19534);
nor U24109 (N_24109,N_17184,N_16212);
or U24110 (N_24110,N_18148,N_15742);
and U24111 (N_24111,N_19462,N_15832);
nor U24112 (N_24112,N_18407,N_17324);
nor U24113 (N_24113,N_16832,N_19973);
nand U24114 (N_24114,N_16492,N_18358);
or U24115 (N_24115,N_18304,N_17997);
and U24116 (N_24116,N_16012,N_17627);
and U24117 (N_24117,N_19993,N_19992);
nand U24118 (N_24118,N_15086,N_18906);
or U24119 (N_24119,N_16542,N_16835);
nand U24120 (N_24120,N_16278,N_16575);
nand U24121 (N_24121,N_15350,N_19760);
nand U24122 (N_24122,N_19526,N_16070);
nor U24123 (N_24123,N_16265,N_16211);
nor U24124 (N_24124,N_15705,N_15399);
and U24125 (N_24125,N_18369,N_18099);
and U24126 (N_24126,N_15799,N_17983);
nand U24127 (N_24127,N_18252,N_19492);
nor U24128 (N_24128,N_19884,N_16192);
nor U24129 (N_24129,N_16296,N_17123);
nor U24130 (N_24130,N_16612,N_19143);
xor U24131 (N_24131,N_18055,N_18387);
or U24132 (N_24132,N_19057,N_19719);
nor U24133 (N_24133,N_18936,N_17386);
nor U24134 (N_24134,N_15811,N_19608);
xor U24135 (N_24135,N_15592,N_16475);
nand U24136 (N_24136,N_15737,N_15012);
and U24137 (N_24137,N_19140,N_17419);
xnor U24138 (N_24138,N_18683,N_16960);
or U24139 (N_24139,N_18819,N_17526);
or U24140 (N_24140,N_17142,N_17447);
nand U24141 (N_24141,N_17391,N_17893);
nand U24142 (N_24142,N_17621,N_19704);
nand U24143 (N_24143,N_15636,N_15295);
and U24144 (N_24144,N_16477,N_16301);
nand U24145 (N_24145,N_15407,N_19686);
xnor U24146 (N_24146,N_18984,N_18726);
nand U24147 (N_24147,N_16094,N_18655);
and U24148 (N_24148,N_17057,N_18368);
nor U24149 (N_24149,N_17044,N_16436);
xnor U24150 (N_24150,N_17659,N_16104);
and U24151 (N_24151,N_18828,N_15981);
xnor U24152 (N_24152,N_17044,N_17805);
xor U24153 (N_24153,N_17254,N_18740);
xnor U24154 (N_24154,N_18834,N_19086);
nor U24155 (N_24155,N_18314,N_15815);
xnor U24156 (N_24156,N_17958,N_18547);
and U24157 (N_24157,N_18106,N_17035);
nor U24158 (N_24158,N_16902,N_15856);
nand U24159 (N_24159,N_17910,N_17008);
or U24160 (N_24160,N_19634,N_19420);
or U24161 (N_24161,N_19657,N_17846);
and U24162 (N_24162,N_15186,N_18592);
and U24163 (N_24163,N_19748,N_19391);
nor U24164 (N_24164,N_17014,N_18699);
and U24165 (N_24165,N_15222,N_19025);
and U24166 (N_24166,N_19417,N_15313);
or U24167 (N_24167,N_18350,N_18058);
nand U24168 (N_24168,N_15072,N_19682);
xor U24169 (N_24169,N_19157,N_17788);
nand U24170 (N_24170,N_15064,N_15703);
xor U24171 (N_24171,N_17874,N_19624);
xnor U24172 (N_24172,N_17293,N_17374);
nand U24173 (N_24173,N_17880,N_15595);
or U24174 (N_24174,N_16012,N_19947);
and U24175 (N_24175,N_19973,N_15634);
and U24176 (N_24176,N_16198,N_18743);
or U24177 (N_24177,N_16007,N_18677);
xnor U24178 (N_24178,N_19741,N_17882);
or U24179 (N_24179,N_16517,N_16250);
xnor U24180 (N_24180,N_16468,N_16756);
or U24181 (N_24181,N_16335,N_16079);
nor U24182 (N_24182,N_15727,N_18113);
and U24183 (N_24183,N_17760,N_18541);
and U24184 (N_24184,N_19056,N_17019);
nor U24185 (N_24185,N_15111,N_18129);
or U24186 (N_24186,N_15238,N_18491);
xnor U24187 (N_24187,N_17873,N_18016);
nor U24188 (N_24188,N_18988,N_17400);
and U24189 (N_24189,N_15454,N_15644);
or U24190 (N_24190,N_18828,N_16629);
and U24191 (N_24191,N_17305,N_19794);
nor U24192 (N_24192,N_19266,N_19611);
xnor U24193 (N_24193,N_16838,N_19011);
xor U24194 (N_24194,N_19986,N_19966);
or U24195 (N_24195,N_17784,N_16657);
nor U24196 (N_24196,N_16785,N_16921);
xnor U24197 (N_24197,N_18979,N_19948);
or U24198 (N_24198,N_18963,N_19702);
or U24199 (N_24199,N_15550,N_16132);
and U24200 (N_24200,N_19075,N_17204);
xnor U24201 (N_24201,N_17727,N_18997);
xor U24202 (N_24202,N_18544,N_16146);
nor U24203 (N_24203,N_18849,N_19785);
xor U24204 (N_24204,N_17972,N_18480);
xor U24205 (N_24205,N_16004,N_15748);
and U24206 (N_24206,N_19841,N_19491);
and U24207 (N_24207,N_16938,N_16764);
nand U24208 (N_24208,N_18116,N_19660);
or U24209 (N_24209,N_19014,N_18607);
or U24210 (N_24210,N_18154,N_18279);
and U24211 (N_24211,N_18255,N_15773);
nand U24212 (N_24212,N_18863,N_17280);
or U24213 (N_24213,N_18595,N_18431);
xnor U24214 (N_24214,N_17970,N_15198);
and U24215 (N_24215,N_17548,N_18838);
nand U24216 (N_24216,N_15372,N_18604);
nor U24217 (N_24217,N_17261,N_16566);
or U24218 (N_24218,N_16865,N_16211);
or U24219 (N_24219,N_15924,N_19377);
xnor U24220 (N_24220,N_16256,N_17335);
or U24221 (N_24221,N_15218,N_19450);
nor U24222 (N_24222,N_19291,N_15492);
nor U24223 (N_24223,N_15138,N_19420);
or U24224 (N_24224,N_19277,N_17275);
xnor U24225 (N_24225,N_19466,N_18687);
nand U24226 (N_24226,N_16646,N_19904);
nor U24227 (N_24227,N_16233,N_16711);
xor U24228 (N_24228,N_16507,N_16672);
xnor U24229 (N_24229,N_15563,N_15786);
nand U24230 (N_24230,N_18972,N_18683);
nor U24231 (N_24231,N_15688,N_19905);
nand U24232 (N_24232,N_18871,N_15066);
nand U24233 (N_24233,N_17645,N_17894);
xor U24234 (N_24234,N_18405,N_15604);
or U24235 (N_24235,N_17499,N_16155);
and U24236 (N_24236,N_15076,N_15186);
or U24237 (N_24237,N_16903,N_18903);
nor U24238 (N_24238,N_17042,N_19988);
nand U24239 (N_24239,N_15849,N_16511);
or U24240 (N_24240,N_15926,N_17359);
and U24241 (N_24241,N_16891,N_18881);
or U24242 (N_24242,N_16082,N_16567);
or U24243 (N_24243,N_15311,N_19332);
and U24244 (N_24244,N_16043,N_15663);
and U24245 (N_24245,N_16255,N_18027);
and U24246 (N_24246,N_19231,N_15925);
xnor U24247 (N_24247,N_17360,N_19634);
nand U24248 (N_24248,N_17770,N_19653);
nor U24249 (N_24249,N_19937,N_18205);
xnor U24250 (N_24250,N_15174,N_15282);
nand U24251 (N_24251,N_16403,N_18601);
xnor U24252 (N_24252,N_18664,N_15632);
nand U24253 (N_24253,N_18136,N_16270);
nor U24254 (N_24254,N_15710,N_18821);
nor U24255 (N_24255,N_16809,N_18476);
or U24256 (N_24256,N_15022,N_15918);
xor U24257 (N_24257,N_16651,N_17928);
nand U24258 (N_24258,N_19366,N_18457);
nor U24259 (N_24259,N_19843,N_16175);
nor U24260 (N_24260,N_18913,N_17172);
and U24261 (N_24261,N_17188,N_15571);
or U24262 (N_24262,N_17415,N_16087);
or U24263 (N_24263,N_18031,N_15367);
xnor U24264 (N_24264,N_19677,N_17908);
nor U24265 (N_24265,N_16963,N_15605);
nand U24266 (N_24266,N_19248,N_16646);
xor U24267 (N_24267,N_18379,N_18554);
nand U24268 (N_24268,N_15405,N_18440);
nor U24269 (N_24269,N_15062,N_19133);
nor U24270 (N_24270,N_16652,N_16184);
nand U24271 (N_24271,N_19375,N_15520);
and U24272 (N_24272,N_19961,N_18854);
nand U24273 (N_24273,N_17654,N_19739);
or U24274 (N_24274,N_17699,N_18968);
and U24275 (N_24275,N_17853,N_18220);
nand U24276 (N_24276,N_16947,N_17008);
xor U24277 (N_24277,N_17026,N_16451);
and U24278 (N_24278,N_15953,N_17246);
xor U24279 (N_24279,N_17253,N_15007);
nand U24280 (N_24280,N_19439,N_18187);
and U24281 (N_24281,N_16251,N_17865);
nor U24282 (N_24282,N_17466,N_15833);
nand U24283 (N_24283,N_18079,N_16908);
nand U24284 (N_24284,N_19013,N_18414);
or U24285 (N_24285,N_16156,N_17629);
or U24286 (N_24286,N_17391,N_18355);
nor U24287 (N_24287,N_17615,N_19123);
nor U24288 (N_24288,N_18559,N_15503);
nand U24289 (N_24289,N_18085,N_16472);
xor U24290 (N_24290,N_17277,N_16179);
nor U24291 (N_24291,N_17618,N_17083);
nor U24292 (N_24292,N_18695,N_18796);
and U24293 (N_24293,N_16235,N_18208);
or U24294 (N_24294,N_19810,N_17079);
xor U24295 (N_24295,N_16436,N_19449);
or U24296 (N_24296,N_16303,N_15001);
nand U24297 (N_24297,N_16987,N_17058);
nand U24298 (N_24298,N_19979,N_18724);
nand U24299 (N_24299,N_15726,N_17444);
or U24300 (N_24300,N_17542,N_17380);
and U24301 (N_24301,N_16037,N_15483);
or U24302 (N_24302,N_19637,N_15045);
and U24303 (N_24303,N_16811,N_16027);
xnor U24304 (N_24304,N_16270,N_18155);
nand U24305 (N_24305,N_16592,N_16572);
or U24306 (N_24306,N_18034,N_19481);
xor U24307 (N_24307,N_17374,N_15067);
and U24308 (N_24308,N_17714,N_19275);
or U24309 (N_24309,N_17535,N_17921);
or U24310 (N_24310,N_15763,N_17408);
nor U24311 (N_24311,N_19564,N_16669);
nor U24312 (N_24312,N_19707,N_19339);
nand U24313 (N_24313,N_19437,N_16233);
nand U24314 (N_24314,N_15986,N_16792);
and U24315 (N_24315,N_19229,N_18996);
nor U24316 (N_24316,N_15555,N_16002);
or U24317 (N_24317,N_15240,N_17656);
or U24318 (N_24318,N_18753,N_16766);
or U24319 (N_24319,N_15515,N_15907);
nand U24320 (N_24320,N_17152,N_15086);
and U24321 (N_24321,N_15433,N_16218);
or U24322 (N_24322,N_15121,N_19442);
nand U24323 (N_24323,N_16684,N_17389);
or U24324 (N_24324,N_18649,N_15224);
xor U24325 (N_24325,N_17284,N_17456);
or U24326 (N_24326,N_19820,N_19879);
and U24327 (N_24327,N_16860,N_17117);
or U24328 (N_24328,N_18903,N_18575);
and U24329 (N_24329,N_16470,N_16094);
xor U24330 (N_24330,N_19181,N_18857);
nor U24331 (N_24331,N_17694,N_18145);
xor U24332 (N_24332,N_18616,N_16494);
xnor U24333 (N_24333,N_19021,N_15682);
and U24334 (N_24334,N_15146,N_15471);
nand U24335 (N_24335,N_19062,N_16055);
and U24336 (N_24336,N_18736,N_19106);
or U24337 (N_24337,N_16081,N_17244);
nand U24338 (N_24338,N_19088,N_17187);
or U24339 (N_24339,N_16387,N_17868);
xor U24340 (N_24340,N_17355,N_18685);
nor U24341 (N_24341,N_19149,N_19895);
or U24342 (N_24342,N_19995,N_15547);
or U24343 (N_24343,N_16802,N_19095);
nor U24344 (N_24344,N_16866,N_16331);
xnor U24345 (N_24345,N_17160,N_16157);
nand U24346 (N_24346,N_16478,N_19910);
xnor U24347 (N_24347,N_15197,N_16333);
xnor U24348 (N_24348,N_18066,N_19783);
and U24349 (N_24349,N_19980,N_18573);
xor U24350 (N_24350,N_15430,N_17496);
or U24351 (N_24351,N_18053,N_16446);
xnor U24352 (N_24352,N_16945,N_19957);
nand U24353 (N_24353,N_19362,N_19118);
xnor U24354 (N_24354,N_16001,N_15990);
xnor U24355 (N_24355,N_16691,N_19502);
nor U24356 (N_24356,N_19721,N_15509);
xnor U24357 (N_24357,N_17652,N_15339);
or U24358 (N_24358,N_18829,N_15454);
nand U24359 (N_24359,N_18594,N_16002);
and U24360 (N_24360,N_19281,N_18126);
nor U24361 (N_24361,N_16552,N_18792);
nor U24362 (N_24362,N_18474,N_17327);
nand U24363 (N_24363,N_17830,N_16772);
or U24364 (N_24364,N_19918,N_19916);
xor U24365 (N_24365,N_18825,N_19145);
xor U24366 (N_24366,N_15659,N_16920);
nor U24367 (N_24367,N_17031,N_17003);
or U24368 (N_24368,N_15179,N_18673);
nor U24369 (N_24369,N_18476,N_18400);
xor U24370 (N_24370,N_19545,N_17111);
nand U24371 (N_24371,N_15980,N_17820);
nor U24372 (N_24372,N_15365,N_19280);
nor U24373 (N_24373,N_19472,N_16727);
and U24374 (N_24374,N_16507,N_15523);
nand U24375 (N_24375,N_16308,N_18240);
or U24376 (N_24376,N_19644,N_15329);
and U24377 (N_24377,N_16529,N_19571);
xnor U24378 (N_24378,N_16138,N_15413);
and U24379 (N_24379,N_17081,N_15198);
or U24380 (N_24380,N_16935,N_15444);
nor U24381 (N_24381,N_17926,N_18397);
nor U24382 (N_24382,N_18789,N_16260);
nor U24383 (N_24383,N_18769,N_17811);
or U24384 (N_24384,N_19810,N_16034);
nand U24385 (N_24385,N_17442,N_19666);
xnor U24386 (N_24386,N_18341,N_17195);
nand U24387 (N_24387,N_15923,N_16429);
nand U24388 (N_24388,N_18932,N_15030);
nand U24389 (N_24389,N_19582,N_15799);
and U24390 (N_24390,N_19319,N_15019);
or U24391 (N_24391,N_19808,N_15195);
nor U24392 (N_24392,N_17689,N_15057);
and U24393 (N_24393,N_15743,N_15256);
xnor U24394 (N_24394,N_19341,N_15126);
or U24395 (N_24395,N_15972,N_19780);
or U24396 (N_24396,N_18452,N_16835);
nor U24397 (N_24397,N_16752,N_17263);
or U24398 (N_24398,N_18048,N_18138);
xnor U24399 (N_24399,N_17696,N_15487);
and U24400 (N_24400,N_19529,N_19705);
nand U24401 (N_24401,N_19125,N_18395);
or U24402 (N_24402,N_15147,N_17943);
nor U24403 (N_24403,N_16210,N_18770);
nor U24404 (N_24404,N_18027,N_18803);
nand U24405 (N_24405,N_17793,N_19436);
nor U24406 (N_24406,N_17535,N_16831);
or U24407 (N_24407,N_17889,N_17003);
and U24408 (N_24408,N_17129,N_15522);
nand U24409 (N_24409,N_19650,N_19351);
xnor U24410 (N_24410,N_17358,N_16495);
or U24411 (N_24411,N_16082,N_15507);
nor U24412 (N_24412,N_16716,N_18633);
xnor U24413 (N_24413,N_16731,N_16752);
and U24414 (N_24414,N_17163,N_15859);
or U24415 (N_24415,N_19509,N_15375);
nor U24416 (N_24416,N_18485,N_18920);
or U24417 (N_24417,N_18285,N_18111);
nor U24418 (N_24418,N_15617,N_19988);
and U24419 (N_24419,N_19564,N_16957);
xor U24420 (N_24420,N_19827,N_18315);
nor U24421 (N_24421,N_16415,N_17192);
and U24422 (N_24422,N_15546,N_19367);
or U24423 (N_24423,N_18622,N_16931);
or U24424 (N_24424,N_19067,N_15158);
xnor U24425 (N_24425,N_18584,N_17016);
and U24426 (N_24426,N_15297,N_17288);
and U24427 (N_24427,N_18165,N_19826);
or U24428 (N_24428,N_17683,N_17424);
xnor U24429 (N_24429,N_16916,N_18552);
nor U24430 (N_24430,N_16952,N_19762);
or U24431 (N_24431,N_17492,N_18216);
and U24432 (N_24432,N_16894,N_17071);
xnor U24433 (N_24433,N_17843,N_16158);
and U24434 (N_24434,N_19144,N_15046);
xor U24435 (N_24435,N_19923,N_17805);
and U24436 (N_24436,N_18713,N_17628);
nand U24437 (N_24437,N_19880,N_16256);
xnor U24438 (N_24438,N_19173,N_19594);
nand U24439 (N_24439,N_16260,N_19406);
nor U24440 (N_24440,N_18985,N_16261);
or U24441 (N_24441,N_16609,N_18492);
xor U24442 (N_24442,N_15121,N_15978);
or U24443 (N_24443,N_19916,N_19355);
or U24444 (N_24444,N_19356,N_19120);
nand U24445 (N_24445,N_15163,N_16037);
nor U24446 (N_24446,N_17024,N_15481);
and U24447 (N_24447,N_19954,N_18966);
nor U24448 (N_24448,N_17737,N_17367);
and U24449 (N_24449,N_17936,N_17642);
nor U24450 (N_24450,N_16999,N_18680);
or U24451 (N_24451,N_18205,N_15450);
nor U24452 (N_24452,N_17331,N_19068);
or U24453 (N_24453,N_15108,N_18913);
nand U24454 (N_24454,N_15539,N_19923);
nor U24455 (N_24455,N_16361,N_19476);
xor U24456 (N_24456,N_16385,N_19828);
or U24457 (N_24457,N_16630,N_19725);
nor U24458 (N_24458,N_19672,N_15910);
or U24459 (N_24459,N_17136,N_17095);
xor U24460 (N_24460,N_18264,N_18607);
nor U24461 (N_24461,N_16218,N_17314);
and U24462 (N_24462,N_15478,N_19896);
nor U24463 (N_24463,N_19709,N_18427);
and U24464 (N_24464,N_15459,N_18281);
nand U24465 (N_24465,N_16134,N_17378);
nor U24466 (N_24466,N_15265,N_17065);
nor U24467 (N_24467,N_16013,N_19850);
or U24468 (N_24468,N_16330,N_18332);
nor U24469 (N_24469,N_18370,N_18381);
xor U24470 (N_24470,N_17752,N_18525);
or U24471 (N_24471,N_15488,N_16564);
nand U24472 (N_24472,N_18338,N_16055);
and U24473 (N_24473,N_19086,N_19839);
nand U24474 (N_24474,N_17987,N_16775);
and U24475 (N_24475,N_19433,N_15581);
or U24476 (N_24476,N_18960,N_17702);
xor U24477 (N_24477,N_19014,N_16392);
xor U24478 (N_24478,N_15154,N_15457);
or U24479 (N_24479,N_16249,N_16272);
xor U24480 (N_24480,N_19507,N_19061);
xnor U24481 (N_24481,N_15148,N_15909);
or U24482 (N_24482,N_17783,N_16883);
nor U24483 (N_24483,N_18131,N_19207);
xor U24484 (N_24484,N_19076,N_15079);
or U24485 (N_24485,N_15191,N_16735);
and U24486 (N_24486,N_15398,N_19945);
and U24487 (N_24487,N_15746,N_19216);
nand U24488 (N_24488,N_16923,N_16473);
nand U24489 (N_24489,N_19736,N_16632);
nor U24490 (N_24490,N_19829,N_19434);
nor U24491 (N_24491,N_16206,N_18168);
and U24492 (N_24492,N_17093,N_17329);
xnor U24493 (N_24493,N_18480,N_18629);
and U24494 (N_24494,N_19841,N_18604);
and U24495 (N_24495,N_18581,N_16683);
or U24496 (N_24496,N_16494,N_19352);
and U24497 (N_24497,N_19181,N_17861);
and U24498 (N_24498,N_15516,N_16157);
and U24499 (N_24499,N_17507,N_17657);
or U24500 (N_24500,N_16738,N_17722);
and U24501 (N_24501,N_15562,N_18763);
nor U24502 (N_24502,N_18044,N_15842);
or U24503 (N_24503,N_19522,N_19646);
xor U24504 (N_24504,N_15563,N_19059);
nor U24505 (N_24505,N_15474,N_17778);
xor U24506 (N_24506,N_18031,N_19229);
xnor U24507 (N_24507,N_16725,N_15729);
or U24508 (N_24508,N_17416,N_17930);
xnor U24509 (N_24509,N_17020,N_19527);
nor U24510 (N_24510,N_16111,N_19834);
or U24511 (N_24511,N_18104,N_15218);
and U24512 (N_24512,N_17222,N_17404);
or U24513 (N_24513,N_18794,N_17431);
or U24514 (N_24514,N_16789,N_19326);
and U24515 (N_24515,N_17018,N_17887);
xor U24516 (N_24516,N_15974,N_15126);
xor U24517 (N_24517,N_15956,N_15952);
nor U24518 (N_24518,N_19237,N_18407);
nand U24519 (N_24519,N_15100,N_17049);
xnor U24520 (N_24520,N_17662,N_15853);
nand U24521 (N_24521,N_17438,N_16457);
or U24522 (N_24522,N_18631,N_16538);
and U24523 (N_24523,N_16280,N_16347);
or U24524 (N_24524,N_15257,N_17477);
xor U24525 (N_24525,N_16624,N_19589);
or U24526 (N_24526,N_15395,N_19467);
nand U24527 (N_24527,N_18462,N_19258);
xor U24528 (N_24528,N_19111,N_18179);
xor U24529 (N_24529,N_17730,N_16596);
or U24530 (N_24530,N_18179,N_18783);
or U24531 (N_24531,N_16981,N_19313);
or U24532 (N_24532,N_18304,N_16547);
or U24533 (N_24533,N_19478,N_15489);
or U24534 (N_24534,N_18215,N_16161);
or U24535 (N_24535,N_19415,N_15790);
nor U24536 (N_24536,N_16932,N_15201);
or U24537 (N_24537,N_18982,N_16220);
nand U24538 (N_24538,N_15562,N_18224);
nor U24539 (N_24539,N_19979,N_17256);
or U24540 (N_24540,N_17657,N_19231);
or U24541 (N_24541,N_17546,N_19723);
nand U24542 (N_24542,N_17012,N_17286);
nand U24543 (N_24543,N_17887,N_19171);
and U24544 (N_24544,N_17039,N_15062);
and U24545 (N_24545,N_17815,N_19001);
xnor U24546 (N_24546,N_15284,N_18438);
nor U24547 (N_24547,N_16009,N_16204);
xor U24548 (N_24548,N_18937,N_18525);
and U24549 (N_24549,N_18654,N_18414);
xnor U24550 (N_24550,N_17521,N_16434);
nor U24551 (N_24551,N_15939,N_18514);
nor U24552 (N_24552,N_15682,N_15103);
nor U24553 (N_24553,N_17371,N_19606);
and U24554 (N_24554,N_15421,N_15320);
and U24555 (N_24555,N_15316,N_15320);
and U24556 (N_24556,N_17489,N_15958);
nand U24557 (N_24557,N_15723,N_18587);
and U24558 (N_24558,N_18973,N_16953);
xor U24559 (N_24559,N_18413,N_16333);
and U24560 (N_24560,N_17610,N_18250);
nor U24561 (N_24561,N_18165,N_15585);
and U24562 (N_24562,N_17517,N_16540);
nor U24563 (N_24563,N_17905,N_16515);
nor U24564 (N_24564,N_17067,N_15350);
and U24565 (N_24565,N_18513,N_17867);
or U24566 (N_24566,N_16225,N_19824);
and U24567 (N_24567,N_17875,N_15535);
nor U24568 (N_24568,N_19597,N_16349);
or U24569 (N_24569,N_19748,N_17917);
or U24570 (N_24570,N_16069,N_19671);
or U24571 (N_24571,N_18423,N_19395);
nor U24572 (N_24572,N_17815,N_19833);
xnor U24573 (N_24573,N_15820,N_16920);
or U24574 (N_24574,N_15827,N_18068);
nor U24575 (N_24575,N_18620,N_18034);
xnor U24576 (N_24576,N_19628,N_18215);
and U24577 (N_24577,N_18887,N_18405);
or U24578 (N_24578,N_18246,N_17456);
and U24579 (N_24579,N_16311,N_15934);
nor U24580 (N_24580,N_16258,N_19407);
nor U24581 (N_24581,N_16064,N_15177);
nor U24582 (N_24582,N_19289,N_18476);
nand U24583 (N_24583,N_15107,N_18395);
or U24584 (N_24584,N_15529,N_15614);
nand U24585 (N_24585,N_16561,N_16896);
xnor U24586 (N_24586,N_17885,N_17407);
nand U24587 (N_24587,N_19944,N_19556);
nor U24588 (N_24588,N_18232,N_16394);
nor U24589 (N_24589,N_18067,N_17096);
and U24590 (N_24590,N_16019,N_17926);
xnor U24591 (N_24591,N_17260,N_18210);
or U24592 (N_24592,N_18522,N_18046);
nor U24593 (N_24593,N_17585,N_18402);
nand U24594 (N_24594,N_15876,N_17559);
xnor U24595 (N_24595,N_18170,N_15782);
xnor U24596 (N_24596,N_19927,N_18409);
nand U24597 (N_24597,N_18052,N_18494);
and U24598 (N_24598,N_15108,N_15701);
xor U24599 (N_24599,N_15337,N_15656);
or U24600 (N_24600,N_17416,N_18953);
nand U24601 (N_24601,N_16588,N_19664);
or U24602 (N_24602,N_18824,N_18750);
xnor U24603 (N_24603,N_16176,N_15508);
or U24604 (N_24604,N_19672,N_16825);
xor U24605 (N_24605,N_15154,N_15906);
or U24606 (N_24606,N_16824,N_19763);
and U24607 (N_24607,N_16773,N_17874);
nand U24608 (N_24608,N_19670,N_19704);
xnor U24609 (N_24609,N_18847,N_17881);
xnor U24610 (N_24610,N_15300,N_15880);
or U24611 (N_24611,N_18842,N_16456);
nor U24612 (N_24612,N_18772,N_15623);
xor U24613 (N_24613,N_15944,N_15812);
and U24614 (N_24614,N_19573,N_18407);
and U24615 (N_24615,N_17575,N_17694);
xor U24616 (N_24616,N_17413,N_16406);
or U24617 (N_24617,N_18261,N_15853);
or U24618 (N_24618,N_16162,N_15625);
or U24619 (N_24619,N_19305,N_18882);
nor U24620 (N_24620,N_18004,N_15366);
xnor U24621 (N_24621,N_15835,N_17962);
nor U24622 (N_24622,N_17388,N_18993);
and U24623 (N_24623,N_17967,N_16171);
nor U24624 (N_24624,N_15265,N_19868);
xnor U24625 (N_24625,N_19472,N_19843);
nand U24626 (N_24626,N_15635,N_18875);
nor U24627 (N_24627,N_17565,N_16484);
nor U24628 (N_24628,N_17512,N_18204);
or U24629 (N_24629,N_16303,N_15075);
xnor U24630 (N_24630,N_17922,N_18207);
and U24631 (N_24631,N_17001,N_16421);
nand U24632 (N_24632,N_19938,N_18557);
or U24633 (N_24633,N_17534,N_17551);
nand U24634 (N_24634,N_15699,N_19802);
and U24635 (N_24635,N_19943,N_19254);
nor U24636 (N_24636,N_17793,N_16948);
nand U24637 (N_24637,N_18418,N_19831);
or U24638 (N_24638,N_18261,N_18689);
or U24639 (N_24639,N_18513,N_18139);
nor U24640 (N_24640,N_18574,N_18358);
nor U24641 (N_24641,N_17545,N_18434);
or U24642 (N_24642,N_18137,N_17122);
nand U24643 (N_24643,N_19080,N_18539);
nand U24644 (N_24644,N_16908,N_17981);
xnor U24645 (N_24645,N_17366,N_19377);
xnor U24646 (N_24646,N_19620,N_15477);
and U24647 (N_24647,N_15688,N_19276);
nor U24648 (N_24648,N_16882,N_17594);
xor U24649 (N_24649,N_19376,N_19144);
or U24650 (N_24650,N_19638,N_19851);
or U24651 (N_24651,N_18948,N_19072);
and U24652 (N_24652,N_16747,N_18555);
and U24653 (N_24653,N_19981,N_19961);
nor U24654 (N_24654,N_18318,N_17846);
nor U24655 (N_24655,N_15038,N_16324);
nor U24656 (N_24656,N_16537,N_18658);
nand U24657 (N_24657,N_18450,N_15173);
nor U24658 (N_24658,N_17214,N_16965);
and U24659 (N_24659,N_16048,N_18904);
nand U24660 (N_24660,N_17718,N_15438);
and U24661 (N_24661,N_18666,N_17222);
or U24662 (N_24662,N_18346,N_17795);
xor U24663 (N_24663,N_17961,N_16258);
and U24664 (N_24664,N_18369,N_19963);
xor U24665 (N_24665,N_17548,N_18900);
nand U24666 (N_24666,N_17794,N_17119);
nand U24667 (N_24667,N_17698,N_16852);
xor U24668 (N_24668,N_15517,N_19826);
or U24669 (N_24669,N_15287,N_18617);
and U24670 (N_24670,N_15790,N_17649);
and U24671 (N_24671,N_19815,N_15779);
and U24672 (N_24672,N_19181,N_17032);
or U24673 (N_24673,N_19119,N_19656);
nand U24674 (N_24674,N_19438,N_17843);
nor U24675 (N_24675,N_19415,N_19297);
and U24676 (N_24676,N_15442,N_16194);
xnor U24677 (N_24677,N_15475,N_17564);
xor U24678 (N_24678,N_19543,N_16020);
xor U24679 (N_24679,N_17031,N_17818);
nand U24680 (N_24680,N_18438,N_17106);
and U24681 (N_24681,N_16764,N_15711);
xnor U24682 (N_24682,N_17654,N_19894);
nor U24683 (N_24683,N_18946,N_15536);
xor U24684 (N_24684,N_16008,N_18814);
nor U24685 (N_24685,N_17594,N_16498);
and U24686 (N_24686,N_16131,N_17095);
nand U24687 (N_24687,N_17087,N_17293);
xnor U24688 (N_24688,N_15410,N_19278);
xor U24689 (N_24689,N_15658,N_16194);
xnor U24690 (N_24690,N_17232,N_17148);
nand U24691 (N_24691,N_19443,N_19195);
or U24692 (N_24692,N_18165,N_18804);
and U24693 (N_24693,N_17447,N_19716);
nand U24694 (N_24694,N_15185,N_19271);
or U24695 (N_24695,N_16250,N_19418);
or U24696 (N_24696,N_16179,N_19957);
nor U24697 (N_24697,N_16615,N_18638);
xor U24698 (N_24698,N_18728,N_16589);
or U24699 (N_24699,N_16691,N_18242);
nor U24700 (N_24700,N_16533,N_19584);
or U24701 (N_24701,N_19582,N_19357);
xnor U24702 (N_24702,N_18742,N_18496);
xnor U24703 (N_24703,N_16818,N_17055);
and U24704 (N_24704,N_17267,N_16034);
or U24705 (N_24705,N_17473,N_15256);
nand U24706 (N_24706,N_18576,N_17822);
nand U24707 (N_24707,N_18385,N_19956);
nor U24708 (N_24708,N_15217,N_17873);
and U24709 (N_24709,N_19262,N_18674);
xor U24710 (N_24710,N_16431,N_19344);
nor U24711 (N_24711,N_15093,N_15510);
nand U24712 (N_24712,N_15128,N_17010);
or U24713 (N_24713,N_16095,N_19473);
xor U24714 (N_24714,N_17810,N_15487);
nand U24715 (N_24715,N_15922,N_17474);
xor U24716 (N_24716,N_17564,N_19154);
or U24717 (N_24717,N_16016,N_18264);
or U24718 (N_24718,N_16107,N_16285);
nor U24719 (N_24719,N_18440,N_16936);
or U24720 (N_24720,N_17637,N_15885);
or U24721 (N_24721,N_16507,N_19242);
nor U24722 (N_24722,N_18644,N_16946);
xnor U24723 (N_24723,N_19704,N_17277);
xnor U24724 (N_24724,N_17245,N_17209);
or U24725 (N_24725,N_15560,N_19561);
nor U24726 (N_24726,N_18915,N_15287);
or U24727 (N_24727,N_18530,N_18227);
xnor U24728 (N_24728,N_19446,N_17556);
nand U24729 (N_24729,N_15924,N_15302);
xor U24730 (N_24730,N_19423,N_19712);
nor U24731 (N_24731,N_18544,N_15698);
nor U24732 (N_24732,N_19076,N_19393);
nor U24733 (N_24733,N_16811,N_19753);
nor U24734 (N_24734,N_17888,N_17379);
xnor U24735 (N_24735,N_18050,N_18423);
nand U24736 (N_24736,N_15327,N_15488);
xor U24737 (N_24737,N_15463,N_15228);
and U24738 (N_24738,N_18268,N_16708);
and U24739 (N_24739,N_15877,N_19475);
or U24740 (N_24740,N_15343,N_19111);
nand U24741 (N_24741,N_18140,N_18842);
xor U24742 (N_24742,N_15400,N_18253);
and U24743 (N_24743,N_15118,N_16152);
nand U24744 (N_24744,N_18984,N_19222);
nand U24745 (N_24745,N_18097,N_19802);
nor U24746 (N_24746,N_19077,N_17577);
or U24747 (N_24747,N_17580,N_19482);
or U24748 (N_24748,N_15488,N_19099);
nor U24749 (N_24749,N_18027,N_16703);
nand U24750 (N_24750,N_18902,N_16651);
nor U24751 (N_24751,N_16382,N_15018);
or U24752 (N_24752,N_17655,N_16808);
and U24753 (N_24753,N_16643,N_19802);
nor U24754 (N_24754,N_15070,N_18120);
and U24755 (N_24755,N_19622,N_17687);
or U24756 (N_24756,N_18423,N_15158);
and U24757 (N_24757,N_17246,N_16278);
and U24758 (N_24758,N_19568,N_16786);
or U24759 (N_24759,N_16257,N_18472);
xnor U24760 (N_24760,N_19833,N_19401);
or U24761 (N_24761,N_18833,N_17397);
or U24762 (N_24762,N_18699,N_18479);
and U24763 (N_24763,N_19450,N_19382);
or U24764 (N_24764,N_16359,N_15722);
xor U24765 (N_24765,N_19633,N_18859);
xor U24766 (N_24766,N_16064,N_17811);
nor U24767 (N_24767,N_18252,N_15688);
xor U24768 (N_24768,N_16421,N_19135);
nor U24769 (N_24769,N_18357,N_16780);
nand U24770 (N_24770,N_18335,N_19354);
nor U24771 (N_24771,N_16706,N_18580);
xnor U24772 (N_24772,N_19360,N_15207);
nor U24773 (N_24773,N_15205,N_16133);
xnor U24774 (N_24774,N_15851,N_15193);
xor U24775 (N_24775,N_18645,N_18174);
or U24776 (N_24776,N_18931,N_16601);
nor U24777 (N_24777,N_15291,N_18720);
and U24778 (N_24778,N_19606,N_17789);
xor U24779 (N_24779,N_19951,N_19836);
nor U24780 (N_24780,N_17108,N_15204);
nor U24781 (N_24781,N_17385,N_18309);
xnor U24782 (N_24782,N_16837,N_17000);
xor U24783 (N_24783,N_18092,N_18569);
nor U24784 (N_24784,N_19430,N_16862);
xor U24785 (N_24785,N_19626,N_15882);
or U24786 (N_24786,N_17674,N_16209);
xnor U24787 (N_24787,N_15767,N_18423);
nor U24788 (N_24788,N_19496,N_17618);
nand U24789 (N_24789,N_17247,N_18686);
xnor U24790 (N_24790,N_16341,N_19881);
and U24791 (N_24791,N_18699,N_15360);
nand U24792 (N_24792,N_17461,N_19486);
and U24793 (N_24793,N_19476,N_17005);
nor U24794 (N_24794,N_16681,N_18044);
nor U24795 (N_24795,N_17809,N_19855);
nor U24796 (N_24796,N_17304,N_15960);
nor U24797 (N_24797,N_15977,N_18964);
or U24798 (N_24798,N_16325,N_16045);
and U24799 (N_24799,N_17019,N_18962);
or U24800 (N_24800,N_18793,N_18492);
xnor U24801 (N_24801,N_16196,N_18738);
and U24802 (N_24802,N_16120,N_15849);
or U24803 (N_24803,N_15312,N_19025);
or U24804 (N_24804,N_18429,N_16673);
nor U24805 (N_24805,N_18871,N_16279);
nor U24806 (N_24806,N_15395,N_19847);
nand U24807 (N_24807,N_15878,N_18096);
xnor U24808 (N_24808,N_16849,N_19264);
or U24809 (N_24809,N_18726,N_16376);
xor U24810 (N_24810,N_16411,N_19694);
nand U24811 (N_24811,N_18136,N_16704);
or U24812 (N_24812,N_19939,N_18071);
or U24813 (N_24813,N_16655,N_15538);
nor U24814 (N_24814,N_18866,N_17269);
and U24815 (N_24815,N_15859,N_16995);
nand U24816 (N_24816,N_19613,N_17074);
nand U24817 (N_24817,N_15523,N_16443);
and U24818 (N_24818,N_17735,N_16269);
nand U24819 (N_24819,N_15824,N_15987);
and U24820 (N_24820,N_16890,N_17041);
xor U24821 (N_24821,N_17825,N_17475);
and U24822 (N_24822,N_16448,N_19431);
or U24823 (N_24823,N_17831,N_17099);
and U24824 (N_24824,N_17078,N_18897);
or U24825 (N_24825,N_15814,N_17558);
xor U24826 (N_24826,N_16761,N_17708);
or U24827 (N_24827,N_16978,N_19500);
nor U24828 (N_24828,N_18206,N_15494);
and U24829 (N_24829,N_18893,N_19065);
or U24830 (N_24830,N_15393,N_16105);
and U24831 (N_24831,N_18638,N_17610);
nand U24832 (N_24832,N_15599,N_18854);
or U24833 (N_24833,N_18780,N_18217);
xnor U24834 (N_24834,N_15597,N_19623);
nor U24835 (N_24835,N_18386,N_17247);
and U24836 (N_24836,N_16768,N_19320);
nor U24837 (N_24837,N_15972,N_15156);
nor U24838 (N_24838,N_16171,N_19272);
xnor U24839 (N_24839,N_16206,N_17185);
nand U24840 (N_24840,N_16560,N_16188);
or U24841 (N_24841,N_18610,N_15520);
or U24842 (N_24842,N_17945,N_16068);
xor U24843 (N_24843,N_15563,N_16773);
nor U24844 (N_24844,N_15216,N_15418);
xnor U24845 (N_24845,N_17042,N_18600);
nor U24846 (N_24846,N_18174,N_19382);
xnor U24847 (N_24847,N_15250,N_19776);
and U24848 (N_24848,N_16265,N_16650);
or U24849 (N_24849,N_17047,N_19736);
or U24850 (N_24850,N_15029,N_17315);
xnor U24851 (N_24851,N_15143,N_18701);
or U24852 (N_24852,N_16918,N_18201);
nand U24853 (N_24853,N_19930,N_15306);
nor U24854 (N_24854,N_17144,N_17690);
nor U24855 (N_24855,N_18989,N_16290);
xnor U24856 (N_24856,N_17876,N_17587);
nor U24857 (N_24857,N_15815,N_17345);
nand U24858 (N_24858,N_16175,N_18211);
nand U24859 (N_24859,N_18131,N_15263);
nand U24860 (N_24860,N_17591,N_18827);
nand U24861 (N_24861,N_15730,N_17396);
nand U24862 (N_24862,N_19682,N_19142);
and U24863 (N_24863,N_15147,N_16183);
and U24864 (N_24864,N_18175,N_17102);
or U24865 (N_24865,N_16309,N_18355);
and U24866 (N_24866,N_18673,N_15776);
or U24867 (N_24867,N_17544,N_19869);
or U24868 (N_24868,N_19256,N_16550);
nor U24869 (N_24869,N_18338,N_16140);
nand U24870 (N_24870,N_16620,N_19961);
or U24871 (N_24871,N_18712,N_18681);
xnor U24872 (N_24872,N_17821,N_17614);
nor U24873 (N_24873,N_17140,N_15992);
and U24874 (N_24874,N_16938,N_19372);
and U24875 (N_24875,N_18170,N_15185);
or U24876 (N_24876,N_19024,N_19574);
nand U24877 (N_24877,N_18146,N_19095);
or U24878 (N_24878,N_15597,N_19982);
nor U24879 (N_24879,N_18984,N_18314);
nand U24880 (N_24880,N_16391,N_17872);
and U24881 (N_24881,N_15672,N_19980);
or U24882 (N_24882,N_19515,N_15075);
xnor U24883 (N_24883,N_17790,N_17272);
xnor U24884 (N_24884,N_16269,N_15293);
xor U24885 (N_24885,N_17891,N_15212);
nand U24886 (N_24886,N_15013,N_16425);
nand U24887 (N_24887,N_19152,N_18708);
xor U24888 (N_24888,N_16420,N_19155);
or U24889 (N_24889,N_19733,N_18693);
or U24890 (N_24890,N_15429,N_18950);
nand U24891 (N_24891,N_19048,N_16229);
nor U24892 (N_24892,N_18729,N_16377);
nor U24893 (N_24893,N_17627,N_15914);
nor U24894 (N_24894,N_16937,N_19076);
nand U24895 (N_24895,N_17547,N_18851);
xnor U24896 (N_24896,N_19640,N_16481);
xnor U24897 (N_24897,N_16956,N_19289);
or U24898 (N_24898,N_19620,N_17932);
xnor U24899 (N_24899,N_17377,N_19926);
and U24900 (N_24900,N_19450,N_16558);
nor U24901 (N_24901,N_15180,N_16554);
and U24902 (N_24902,N_15608,N_19225);
and U24903 (N_24903,N_16082,N_15981);
xor U24904 (N_24904,N_15963,N_19518);
xnor U24905 (N_24905,N_16943,N_19119);
nand U24906 (N_24906,N_19801,N_15435);
nor U24907 (N_24907,N_17511,N_17149);
and U24908 (N_24908,N_19139,N_18290);
xor U24909 (N_24909,N_15023,N_17738);
or U24910 (N_24910,N_19523,N_15302);
nor U24911 (N_24911,N_16652,N_16277);
nand U24912 (N_24912,N_16483,N_18206);
xor U24913 (N_24913,N_15286,N_15471);
nand U24914 (N_24914,N_19708,N_19178);
nor U24915 (N_24915,N_17132,N_19839);
xnor U24916 (N_24916,N_15051,N_15594);
xnor U24917 (N_24917,N_18392,N_19301);
and U24918 (N_24918,N_15875,N_15129);
and U24919 (N_24919,N_18935,N_18770);
nor U24920 (N_24920,N_17971,N_19464);
xor U24921 (N_24921,N_15524,N_17438);
nand U24922 (N_24922,N_16271,N_17757);
or U24923 (N_24923,N_18790,N_18299);
or U24924 (N_24924,N_17498,N_18422);
and U24925 (N_24925,N_16604,N_17583);
xor U24926 (N_24926,N_19770,N_15700);
xor U24927 (N_24927,N_15581,N_16247);
nor U24928 (N_24928,N_18832,N_19422);
nand U24929 (N_24929,N_17568,N_17986);
and U24930 (N_24930,N_16805,N_16862);
nand U24931 (N_24931,N_15550,N_19585);
and U24932 (N_24932,N_18261,N_16381);
nor U24933 (N_24933,N_17541,N_17074);
xor U24934 (N_24934,N_16745,N_15010);
xnor U24935 (N_24935,N_15143,N_15390);
nand U24936 (N_24936,N_16719,N_18135);
nor U24937 (N_24937,N_18127,N_18941);
or U24938 (N_24938,N_18614,N_15396);
nand U24939 (N_24939,N_18945,N_19904);
and U24940 (N_24940,N_15313,N_15739);
or U24941 (N_24941,N_17910,N_18508);
or U24942 (N_24942,N_16149,N_16464);
xnor U24943 (N_24943,N_18385,N_19340);
nand U24944 (N_24944,N_15156,N_16785);
or U24945 (N_24945,N_18651,N_18787);
or U24946 (N_24946,N_19097,N_19161);
nand U24947 (N_24947,N_15476,N_16580);
and U24948 (N_24948,N_16390,N_15387);
nand U24949 (N_24949,N_16280,N_15991);
and U24950 (N_24950,N_15382,N_17990);
xor U24951 (N_24951,N_17517,N_19491);
or U24952 (N_24952,N_19495,N_19587);
xnor U24953 (N_24953,N_19496,N_19581);
and U24954 (N_24954,N_16254,N_17261);
nand U24955 (N_24955,N_18179,N_15710);
and U24956 (N_24956,N_16937,N_17262);
xnor U24957 (N_24957,N_17136,N_19830);
or U24958 (N_24958,N_18152,N_17965);
and U24959 (N_24959,N_15262,N_16179);
xnor U24960 (N_24960,N_17224,N_18828);
nor U24961 (N_24961,N_16701,N_16477);
or U24962 (N_24962,N_16736,N_18119);
or U24963 (N_24963,N_18899,N_15984);
nand U24964 (N_24964,N_15963,N_19962);
and U24965 (N_24965,N_19522,N_16624);
nor U24966 (N_24966,N_15300,N_15913);
or U24967 (N_24967,N_17482,N_15436);
nand U24968 (N_24968,N_16214,N_17625);
nor U24969 (N_24969,N_19503,N_19053);
or U24970 (N_24970,N_18037,N_17732);
and U24971 (N_24971,N_16720,N_15659);
or U24972 (N_24972,N_15653,N_15797);
nand U24973 (N_24973,N_16120,N_15983);
and U24974 (N_24974,N_16371,N_17708);
or U24975 (N_24975,N_15575,N_18273);
nor U24976 (N_24976,N_17446,N_19306);
xor U24977 (N_24977,N_15413,N_15469);
xnor U24978 (N_24978,N_18784,N_18196);
or U24979 (N_24979,N_19093,N_17199);
xnor U24980 (N_24980,N_16826,N_16434);
nor U24981 (N_24981,N_18747,N_19328);
nand U24982 (N_24982,N_16898,N_15189);
nor U24983 (N_24983,N_17675,N_17070);
xor U24984 (N_24984,N_15904,N_17409);
nand U24985 (N_24985,N_18230,N_19836);
xnor U24986 (N_24986,N_17524,N_17208);
and U24987 (N_24987,N_15430,N_16863);
nor U24988 (N_24988,N_17902,N_19363);
or U24989 (N_24989,N_15530,N_19033);
and U24990 (N_24990,N_16577,N_19714);
xnor U24991 (N_24991,N_19273,N_18844);
or U24992 (N_24992,N_18131,N_19197);
xnor U24993 (N_24993,N_19483,N_15230);
or U24994 (N_24994,N_15095,N_19627);
nand U24995 (N_24995,N_17564,N_19160);
nor U24996 (N_24996,N_16554,N_19599);
and U24997 (N_24997,N_15409,N_15411);
xor U24998 (N_24998,N_17709,N_18497);
nand U24999 (N_24999,N_16482,N_19546);
xor U25000 (N_25000,N_21977,N_21800);
nand U25001 (N_25001,N_22086,N_20551);
and U25002 (N_25002,N_21118,N_21584);
and U25003 (N_25003,N_22590,N_21703);
xnor U25004 (N_25004,N_21120,N_23997);
xor U25005 (N_25005,N_22288,N_22687);
nor U25006 (N_25006,N_21032,N_22025);
or U25007 (N_25007,N_22990,N_24838);
and U25008 (N_25008,N_21166,N_21681);
or U25009 (N_25009,N_23360,N_20645);
xnor U25010 (N_25010,N_20557,N_23575);
and U25011 (N_25011,N_24138,N_23647);
xnor U25012 (N_25012,N_20313,N_20742);
or U25013 (N_25013,N_23762,N_23929);
nor U25014 (N_25014,N_21980,N_22319);
nand U25015 (N_25015,N_23534,N_22854);
and U25016 (N_25016,N_22313,N_22029);
or U25017 (N_25017,N_20496,N_21250);
nand U25018 (N_25018,N_21184,N_24526);
nand U25019 (N_25019,N_24034,N_21914);
nand U25020 (N_25020,N_21633,N_21056);
or U25021 (N_25021,N_23112,N_22382);
nor U25022 (N_25022,N_20994,N_24864);
nand U25023 (N_25023,N_21626,N_24994);
and U25024 (N_25024,N_21135,N_23644);
nor U25025 (N_25025,N_20656,N_23837);
and U25026 (N_25026,N_22176,N_22519);
nor U25027 (N_25027,N_20217,N_20368);
or U25028 (N_25028,N_21875,N_23808);
and U25029 (N_25029,N_22484,N_20930);
xnor U25030 (N_25030,N_20278,N_21234);
or U25031 (N_25031,N_21946,N_21768);
xor U25032 (N_25032,N_24287,N_24230);
and U25033 (N_25033,N_22035,N_21030);
nor U25034 (N_25034,N_22435,N_23803);
nor U25035 (N_25035,N_23556,N_21782);
nor U25036 (N_25036,N_22521,N_21867);
or U25037 (N_25037,N_24750,N_21085);
nand U25038 (N_25038,N_20296,N_22381);
and U25039 (N_25039,N_24854,N_20195);
and U25040 (N_25040,N_20956,N_24359);
nand U25041 (N_25041,N_21669,N_24078);
xor U25042 (N_25042,N_21422,N_24350);
xnor U25043 (N_25043,N_22424,N_24384);
and U25044 (N_25044,N_22306,N_21581);
nand U25045 (N_25045,N_22820,N_23405);
and U25046 (N_25046,N_21114,N_20820);
nand U25047 (N_25047,N_20934,N_20796);
or U25048 (N_25048,N_21452,N_21022);
or U25049 (N_25049,N_21677,N_20522);
xnor U25050 (N_25050,N_20276,N_20580);
nand U25051 (N_25051,N_23468,N_23527);
nand U25052 (N_25052,N_22165,N_22123);
xnor U25053 (N_25053,N_20570,N_20733);
and U25054 (N_25054,N_20248,N_22146);
nand U25055 (N_25055,N_23311,N_20401);
and U25056 (N_25056,N_20176,N_24159);
and U25057 (N_25057,N_22623,N_22103);
or U25058 (N_25058,N_21215,N_20170);
or U25059 (N_25059,N_23028,N_24153);
or U25060 (N_25060,N_23267,N_24024);
nand U25061 (N_25061,N_24545,N_22612);
xor U25062 (N_25062,N_22981,N_20443);
nand U25063 (N_25063,N_20495,N_24115);
nor U25064 (N_25064,N_21941,N_23503);
nand U25065 (N_25065,N_22971,N_23895);
and U25066 (N_25066,N_21722,N_21792);
nor U25067 (N_25067,N_20397,N_22143);
or U25068 (N_25068,N_24829,N_20130);
nor U25069 (N_25069,N_21299,N_23716);
nor U25070 (N_25070,N_21212,N_22752);
xor U25071 (N_25071,N_23023,N_24665);
nor U25072 (N_25072,N_20494,N_23707);
and U25073 (N_25073,N_22802,N_21053);
nand U25074 (N_25074,N_22145,N_23865);
xor U25075 (N_25075,N_22371,N_22336);
nor U25076 (N_25076,N_23990,N_23072);
xnor U25077 (N_25077,N_21610,N_23806);
xnor U25078 (N_25078,N_20970,N_20197);
and U25079 (N_25079,N_21658,N_22104);
xnor U25080 (N_25080,N_21324,N_22586);
nor U25081 (N_25081,N_20751,N_24587);
and U25082 (N_25082,N_21006,N_22005);
or U25083 (N_25083,N_22046,N_23443);
and U25084 (N_25084,N_22679,N_21932);
or U25085 (N_25085,N_22642,N_20345);
or U25086 (N_25086,N_24174,N_20892);
nand U25087 (N_25087,N_24134,N_23768);
xnor U25088 (N_25088,N_24708,N_21544);
xnor U25089 (N_25089,N_20663,N_21576);
or U25090 (N_25090,N_20490,N_21958);
and U25091 (N_25091,N_24530,N_21121);
xnor U25092 (N_25092,N_21442,N_22106);
or U25093 (N_25093,N_24289,N_23886);
nor U25094 (N_25094,N_20251,N_24692);
xnor U25095 (N_25095,N_24327,N_24308);
nand U25096 (N_25096,N_22727,N_23129);
nand U25097 (N_25097,N_24978,N_24171);
nor U25098 (N_25098,N_21163,N_21758);
or U25099 (N_25099,N_21638,N_21865);
nand U25100 (N_25100,N_21690,N_23827);
xnor U25101 (N_25101,N_20372,N_24787);
or U25102 (N_25102,N_20953,N_24229);
xnor U25103 (N_25103,N_22048,N_21027);
xor U25104 (N_25104,N_21819,N_23348);
xor U25105 (N_25105,N_21482,N_20469);
nor U25106 (N_25106,N_24993,N_24248);
xnor U25107 (N_25107,N_23027,N_23275);
nand U25108 (N_25108,N_24463,N_23152);
nand U25109 (N_25109,N_24756,N_21298);
or U25110 (N_25110,N_20291,N_24728);
nand U25111 (N_25111,N_20936,N_22002);
nor U25112 (N_25112,N_24443,N_22461);
nand U25113 (N_25113,N_23935,N_24607);
xor U25114 (N_25114,N_24555,N_22695);
nor U25115 (N_25115,N_20132,N_21582);
nand U25116 (N_25116,N_21892,N_22865);
and U25117 (N_25117,N_23001,N_20019);
nand U25118 (N_25118,N_21940,N_20428);
or U25119 (N_25119,N_23227,N_21833);
or U25120 (N_25120,N_21342,N_21099);
and U25121 (N_25121,N_21090,N_23045);
xor U25122 (N_25122,N_24210,N_22677);
and U25123 (N_25123,N_23614,N_20235);
nor U25124 (N_25124,N_22648,N_22730);
and U25125 (N_25125,N_24638,N_22515);
nand U25126 (N_25126,N_22600,N_20288);
and U25127 (N_25127,N_22208,N_23479);
and U25128 (N_25128,N_24066,N_20491);
nand U25129 (N_25129,N_24346,N_21534);
nand U25130 (N_25130,N_24061,N_23943);
nor U25131 (N_25131,N_21232,N_20593);
nand U25132 (N_25132,N_22894,N_20875);
and U25133 (N_25133,N_22417,N_23453);
nand U25134 (N_25134,N_20781,N_21469);
nor U25135 (N_25135,N_21919,N_20531);
xor U25136 (N_25136,N_24619,N_20754);
nand U25137 (N_25137,N_24431,N_20699);
nand U25138 (N_25138,N_22090,N_20894);
nor U25139 (N_25139,N_24893,N_21315);
nor U25140 (N_25140,N_23113,N_23344);
or U25141 (N_25141,N_20436,N_23017);
nor U25142 (N_25142,N_20358,N_24533);
xor U25143 (N_25143,N_20474,N_24483);
nor U25144 (N_25144,N_23870,N_24591);
and U25145 (N_25145,N_22310,N_21850);
nand U25146 (N_25146,N_20701,N_23298);
xor U25147 (N_25147,N_24840,N_22431);
xor U25148 (N_25148,N_23730,N_20745);
xor U25149 (N_25149,N_21297,N_23821);
xor U25150 (N_25150,N_22693,N_23628);
or U25151 (N_25151,N_22668,N_21441);
xor U25152 (N_25152,N_20838,N_21578);
or U25153 (N_25153,N_22523,N_21730);
nor U25154 (N_25154,N_23334,N_20339);
and U25155 (N_25155,N_23277,N_24490);
nor U25156 (N_25156,N_22560,N_20383);
nand U25157 (N_25157,N_20918,N_23752);
nor U25158 (N_25158,N_24070,N_23799);
xnor U25159 (N_25159,N_22286,N_24405);
and U25160 (N_25160,N_20660,N_21087);
xnor U25161 (N_25161,N_23502,N_20691);
nand U25162 (N_25162,N_20343,N_24075);
xor U25163 (N_25163,N_24570,N_20211);
and U25164 (N_25164,N_24636,N_20074);
or U25165 (N_25165,N_23914,N_23404);
and U25166 (N_25166,N_20560,N_23018);
nand U25167 (N_25167,N_20878,N_20695);
and U25168 (N_25168,N_22979,N_23492);
xor U25169 (N_25169,N_24107,N_21863);
nand U25170 (N_25170,N_20434,N_22657);
nand U25171 (N_25171,N_24009,N_22229);
nor U25172 (N_25172,N_20135,N_22446);
or U25173 (N_25173,N_20033,N_20402);
xor U25174 (N_25174,N_23535,N_24317);
nor U25175 (N_25175,N_24047,N_22798);
xor U25176 (N_25176,N_23209,N_23498);
nor U25177 (N_25177,N_24554,N_23412);
nand U25178 (N_25178,N_23450,N_20737);
xnor U25179 (N_25179,N_20566,N_24195);
nand U25180 (N_25180,N_22686,N_22060);
xor U25181 (N_25181,N_24960,N_20206);
or U25182 (N_25182,N_20225,N_20629);
xor U25183 (N_25183,N_22643,N_24778);
or U25184 (N_25184,N_23048,N_22154);
or U25185 (N_25185,N_20022,N_20117);
and U25186 (N_25186,N_21507,N_22673);
nand U25187 (N_25187,N_23156,N_23099);
xnor U25188 (N_25188,N_21778,N_23121);
or U25189 (N_25189,N_23012,N_23847);
nor U25190 (N_25190,N_23949,N_20308);
xor U25191 (N_25191,N_23733,N_24017);
nand U25192 (N_25192,N_20384,N_24509);
nor U25193 (N_25193,N_24858,N_21779);
nand U25194 (N_25194,N_24576,N_23473);
or U25195 (N_25195,N_24358,N_24502);
nor U25196 (N_25196,N_21585,N_24725);
nand U25197 (N_25197,N_23105,N_21304);
nor U25198 (N_25198,N_22869,N_22985);
nand U25199 (N_25199,N_23223,N_20046);
and U25200 (N_25200,N_23153,N_22471);
or U25201 (N_25201,N_20957,N_22770);
or U25202 (N_25202,N_22287,N_22557);
nor U25203 (N_25203,N_22055,N_23608);
and U25204 (N_25204,N_20357,N_23258);
nand U25205 (N_25205,N_22181,N_24727);
nor U25206 (N_25206,N_22159,N_24142);
xnor U25207 (N_25207,N_22924,N_22934);
xor U25208 (N_25208,N_20649,N_24455);
xnor U25209 (N_25209,N_22082,N_22066);
xor U25210 (N_25210,N_21489,N_22353);
nand U25211 (N_25211,N_21479,N_20342);
and U25212 (N_25212,N_22380,N_20855);
nand U25213 (N_25213,N_22716,N_24713);
nand U25214 (N_25214,N_24139,N_20785);
or U25215 (N_25215,N_24785,N_24808);
nand U25216 (N_25216,N_23236,N_24557);
and U25217 (N_25217,N_23703,N_23470);
nand U25218 (N_25218,N_22737,N_21186);
or U25219 (N_25219,N_20452,N_20584);
nand U25220 (N_25220,N_21628,N_22290);
nor U25221 (N_25221,N_21216,N_22470);
or U25222 (N_25222,N_22553,N_23335);
xor U25223 (N_25223,N_21895,N_24300);
or U25224 (N_25224,N_22121,N_21123);
and U25225 (N_25225,N_21765,N_21648);
nand U25226 (N_25226,N_23967,N_21495);
xor U25227 (N_25227,N_23930,N_24241);
xnor U25228 (N_25228,N_20836,N_21143);
xor U25229 (N_25229,N_21321,N_21876);
or U25230 (N_25230,N_21359,N_21011);
nor U25231 (N_25231,N_23230,N_22655);
or U25232 (N_25232,N_24933,N_20616);
nand U25233 (N_25233,N_20827,N_21275);
xor U25234 (N_25234,N_22087,N_21897);
and U25235 (N_25235,N_23651,N_23588);
xnor U25236 (N_25236,N_23096,N_24745);
or U25237 (N_25237,N_23330,N_22621);
nand U25238 (N_25238,N_21427,N_23970);
nand U25239 (N_25239,N_23228,N_23579);
xor U25240 (N_25240,N_22913,N_22428);
nor U25241 (N_25241,N_22000,N_23071);
or U25242 (N_25242,N_22163,N_22853);
xnor U25243 (N_25243,N_21246,N_23869);
or U25244 (N_25244,N_23325,N_22749);
or U25245 (N_25245,N_23781,N_22567);
or U25246 (N_25246,N_20377,N_22721);
xnor U25247 (N_25247,N_23260,N_21725);
and U25248 (N_25248,N_22626,N_20112);
and U25249 (N_25249,N_23370,N_22469);
nand U25250 (N_25250,N_24562,N_24328);
nand U25251 (N_25251,N_23904,N_22710);
and U25252 (N_25252,N_22440,N_23116);
nand U25253 (N_25253,N_21686,N_20548);
nand U25254 (N_25254,N_21645,N_22303);
nor U25255 (N_25255,N_24222,N_20529);
xnor U25256 (N_25256,N_20344,N_22045);
nor U25257 (N_25257,N_24190,N_24668);
nand U25258 (N_25258,N_24313,N_22624);
xor U25259 (N_25259,N_22312,N_21075);
and U25260 (N_25260,N_24495,N_23905);
nor U25261 (N_25261,N_20488,N_23994);
or U25262 (N_25262,N_20067,N_20035);
xnor U25263 (N_25263,N_20111,N_22806);
nor U25264 (N_25264,N_22453,N_23823);
nor U25265 (N_25265,N_21004,N_20741);
nand U25266 (N_25266,N_24296,N_23771);
nor U25267 (N_25267,N_21860,N_23235);
nor U25268 (N_25268,N_22191,N_20779);
xor U25269 (N_25269,N_22351,N_20614);
nor U25270 (N_25270,N_23415,N_24506);
or U25271 (N_25271,N_24039,N_22972);
xor U25272 (N_25272,N_21367,N_22615);
nand U25273 (N_25273,N_20724,N_24802);
nor U25274 (N_25274,N_23124,N_22199);
or U25275 (N_25275,N_20759,N_24236);
or U25276 (N_25276,N_23397,N_24322);
or U25277 (N_25277,N_23119,N_22348);
xnor U25278 (N_25278,N_20350,N_23182);
or U25279 (N_25279,N_21404,N_22040);
nand U25280 (N_25280,N_20194,N_24771);
nor U25281 (N_25281,N_24501,N_23368);
or U25282 (N_25282,N_23142,N_20030);
xnor U25283 (N_25283,N_22999,N_21437);
xor U25284 (N_25284,N_21736,N_20743);
nand U25285 (N_25285,N_21459,N_20347);
and U25286 (N_25286,N_20872,N_24967);
and U25287 (N_25287,N_21943,N_24408);
or U25288 (N_25288,N_23437,N_24003);
and U25289 (N_25289,N_23778,N_24605);
and U25290 (N_25290,N_21222,N_21912);
or U25291 (N_25291,N_20250,N_20861);
xor U25292 (N_25292,N_22747,N_23463);
xnor U25293 (N_25293,N_21844,N_23438);
or U25294 (N_25294,N_23361,N_22337);
or U25295 (N_25295,N_20240,N_24564);
nand U25296 (N_25296,N_20230,N_24887);
or U25297 (N_25297,N_20232,N_24321);
nor U25298 (N_25298,N_21365,N_21134);
and U25299 (N_25299,N_22361,N_24970);
and U25300 (N_25300,N_22980,N_23871);
and U25301 (N_25301,N_24316,N_20795);
or U25302 (N_25302,N_20717,N_24228);
or U25303 (N_25303,N_22259,N_23441);
or U25304 (N_25304,N_24611,N_22463);
nand U25305 (N_25305,N_24029,N_22734);
nand U25306 (N_25306,N_20025,N_20858);
nand U25307 (N_25307,N_24733,N_20059);
xor U25308 (N_25308,N_20245,N_21543);
nor U25309 (N_25309,N_21629,N_21732);
and U25310 (N_25310,N_20830,N_23559);
xor U25311 (N_25311,N_23585,N_20804);
or U25312 (N_25312,N_20416,N_20806);
nor U25313 (N_25313,N_22292,N_22606);
or U25314 (N_25314,N_24467,N_24176);
or U25315 (N_25315,N_22868,N_24238);
or U25316 (N_25316,N_24233,N_23478);
xnor U25317 (N_25317,N_22419,N_24937);
nor U25318 (N_25318,N_22033,N_20601);
and U25319 (N_25319,N_21081,N_22161);
nand U25320 (N_25320,N_22534,N_21557);
nor U25321 (N_25321,N_21862,N_21453);
or U25322 (N_25322,N_20281,N_21682);
nor U25323 (N_25323,N_23369,N_20845);
or U25324 (N_25324,N_21711,N_22038);
nand U25325 (N_25325,N_22438,N_21999);
nor U25326 (N_25326,N_21942,N_20465);
xor U25327 (N_25327,N_20047,N_23154);
or U25328 (N_25328,N_22363,N_22877);
or U25329 (N_25329,N_24684,N_20193);
xor U25330 (N_25330,N_22723,N_20640);
nand U25331 (N_25331,N_22340,N_23067);
nand U25332 (N_25332,N_23328,N_21073);
nand U25333 (N_25333,N_21068,N_22284);
nand U25334 (N_25334,N_23723,N_21513);
nand U25335 (N_25335,N_22997,N_23576);
nand U25336 (N_25336,N_20951,N_20773);
nor U25337 (N_25337,N_21806,N_23798);
or U25338 (N_25338,N_23489,N_20846);
and U25339 (N_25339,N_22758,N_22549);
xnor U25340 (N_25340,N_24199,N_20776);
nor U25341 (N_25341,N_24675,N_20188);
or U25342 (N_25342,N_24215,N_20774);
or U25343 (N_25343,N_21036,N_24439);
nor U25344 (N_25344,N_23593,N_21530);
nor U25345 (N_25345,N_21088,N_23831);
nand U25346 (N_25346,N_24757,N_22575);
nand U25347 (N_25347,N_21928,N_22358);
nor U25348 (N_25348,N_24342,N_23046);
xnor U25349 (N_25349,N_22269,N_22239);
and U25350 (N_25350,N_21592,N_24433);
and U25351 (N_25351,N_20935,N_22119);
nand U25352 (N_25352,N_24486,N_23237);
and U25353 (N_25353,N_20317,N_20987);
nor U25354 (N_25354,N_20627,N_22539);
nand U25355 (N_25355,N_22374,N_22212);
xnor U25356 (N_25356,N_22091,N_20760);
nor U25357 (N_25357,N_22230,N_20700);
or U25358 (N_25358,N_20068,N_23530);
or U25359 (N_25359,N_20532,N_24069);
nand U25360 (N_25360,N_22840,N_24453);
or U25361 (N_25361,N_22681,N_24044);
nor U25362 (N_25362,N_20525,N_22728);
nor U25363 (N_25363,N_20139,N_24451);
nand U25364 (N_25364,N_24318,N_20438);
xnor U25365 (N_25365,N_21559,N_23175);
nor U25366 (N_25366,N_22244,N_20221);
or U25367 (N_25367,N_24381,N_20018);
xnor U25368 (N_25368,N_21655,N_24830);
xnor U25369 (N_25369,N_24147,N_22225);
xnor U25370 (N_25370,N_21458,N_21745);
nor U25371 (N_25371,N_21107,N_22291);
xnor U25372 (N_25372,N_24773,N_21522);
nor U25373 (N_25373,N_20198,N_23688);
nand U25374 (N_25374,N_21301,N_20307);
nor U25375 (N_25375,N_22079,N_22878);
xor U25376 (N_25376,N_20683,N_20455);
nor U25377 (N_25377,N_20052,N_23190);
nor U25378 (N_25378,N_23711,N_20320);
nand U25379 (N_25379,N_21751,N_21370);
and U25380 (N_25380,N_24989,N_23747);
xor U25381 (N_25381,N_24052,N_20723);
nor U25382 (N_25382,N_23891,N_21277);
nor U25383 (N_25383,N_22334,N_24437);
and U25384 (N_25384,N_22335,N_22430);
nand U25385 (N_25385,N_22107,N_21937);
nor U25386 (N_25386,N_22565,N_23481);
or U25387 (N_25387,N_23801,N_22186);
nand U25388 (N_25388,N_23381,N_21217);
and U25389 (N_25389,N_20355,N_24632);
nand U25390 (N_25390,N_23898,N_24064);
and U25391 (N_25391,N_23972,N_23064);
or U25392 (N_25392,N_20429,N_23138);
xnor U25393 (N_25393,N_24946,N_22318);
and U25394 (N_25394,N_23954,N_22187);
nor U25395 (N_25395,N_22860,N_24374);
or U25396 (N_25396,N_20937,N_23329);
nor U25397 (N_25397,N_20422,N_24444);
xnor U25398 (N_25398,N_21790,N_21274);
xor U25399 (N_25399,N_23186,N_22366);
nor U25400 (N_25400,N_23336,N_22058);
nand U25401 (N_25401,N_22157,N_24097);
and U25402 (N_25402,N_23996,N_20991);
nor U25403 (N_25403,N_23777,N_23735);
nand U25404 (N_25404,N_22164,N_20579);
or U25405 (N_25405,N_23928,N_22569);
or U25406 (N_25406,N_23517,N_20254);
and U25407 (N_25407,N_22817,N_24341);
nand U25408 (N_25408,N_21033,N_20406);
nor U25409 (N_25409,N_20088,N_22684);
or U25410 (N_25410,N_23849,N_24677);
or U25411 (N_25411,N_21480,N_21352);
and U25412 (N_25412,N_22257,N_21858);
nor U25413 (N_25413,N_24376,N_21188);
or U25414 (N_25414,N_22432,N_23496);
nand U25415 (N_25415,N_24456,N_24368);
nor U25416 (N_25416,N_23571,N_24247);
xor U25417 (N_25417,N_22509,N_21528);
xor U25418 (N_25418,N_22698,N_23308);
nand U25419 (N_25419,N_24340,N_20376);
nand U25420 (N_25420,N_23592,N_20228);
and U25421 (N_25421,N_21938,N_24105);
nor U25422 (N_25422,N_24286,N_24538);
nor U25423 (N_25423,N_22405,N_24415);
and U25424 (N_25424,N_20405,N_24759);
or U25425 (N_25425,N_22881,N_23856);
xnor U25426 (N_25426,N_23456,N_24901);
xor U25427 (N_25427,N_21093,N_22604);
or U25428 (N_25428,N_22576,N_21335);
or U25429 (N_25429,N_24655,N_20910);
or U25430 (N_25430,N_23565,N_21735);
and U25431 (N_25431,N_23003,N_22670);
nor U25432 (N_25432,N_21089,N_20960);
xnor U25433 (N_25433,N_21696,N_22571);
nor U25434 (N_25434,N_20972,N_23459);
or U25435 (N_25435,N_20899,N_23538);
xor U25436 (N_25436,N_24478,N_22421);
and U25437 (N_25437,N_20905,N_24053);
and U25438 (N_25438,N_24001,N_23818);
xnor U25439 (N_25439,N_21096,N_23695);
nand U25440 (N_25440,N_21925,N_20694);
xor U25441 (N_25441,N_23514,N_24984);
nand U25442 (N_25442,N_23687,N_20702);
or U25443 (N_25443,N_20369,N_24481);
xnor U25444 (N_25444,N_20886,N_22426);
and U25445 (N_25445,N_21969,N_20044);
or U25446 (N_25446,N_23766,N_20908);
nand U25447 (N_25447,N_21287,N_21380);
and U25448 (N_25448,N_23761,N_24109);
nand U25449 (N_25449,N_21260,N_24323);
nor U25450 (N_25450,N_23050,N_21181);
nand U25451 (N_25451,N_23399,N_23937);
xnor U25452 (N_25452,N_22732,N_23518);
xor U25453 (N_25453,N_23155,N_24649);
nor U25454 (N_25454,N_21041,N_20985);
xnor U25455 (N_25455,N_21891,N_24315);
and U25456 (N_25456,N_22513,N_24312);
nand U25457 (N_25457,N_24098,N_22117);
and U25458 (N_25458,N_23342,N_24263);
nor U25459 (N_25459,N_24461,N_20750);
and U25460 (N_25460,N_21464,N_24599);
nand U25461 (N_25461,N_22053,N_23097);
xnor U25462 (N_25462,N_23109,N_21944);
nand U25463 (N_25463,N_20940,N_23650);
and U25464 (N_25464,N_24423,N_22849);
xor U25465 (N_25465,N_21278,N_24297);
nand U25466 (N_25466,N_21237,N_24640);
nand U25467 (N_25467,N_22198,N_23805);
and U25468 (N_25468,N_20187,N_21547);
and U25469 (N_25469,N_21069,N_24542);
or U25470 (N_25470,N_22021,N_23157);
xor U25471 (N_25471,N_23875,N_24399);
or U25472 (N_25472,N_21151,N_23120);
or U25473 (N_25473,N_21265,N_22299);
nor U25474 (N_25474,N_21071,N_22378);
or U25475 (N_25475,N_24087,N_20208);
or U25476 (N_25476,N_21018,N_22223);
nand U25477 (N_25477,N_20562,N_23883);
or U25478 (N_25478,N_23881,N_23901);
nor U25479 (N_25479,N_22388,N_20105);
or U25480 (N_25480,N_20965,N_21887);
and U25481 (N_25481,N_24927,N_24332);
and U25482 (N_25482,N_22221,N_23697);
and U25483 (N_25483,N_24696,N_23991);
nand U25484 (N_25484,N_21492,N_24791);
or U25485 (N_25485,N_22905,N_24569);
nand U25486 (N_25486,N_23522,N_23266);
or U25487 (N_25487,N_23379,N_20658);
and U25488 (N_25488,N_21175,N_23654);
nand U25489 (N_25489,N_21567,N_20073);
and U25490 (N_25490,N_21490,N_23164);
or U25491 (N_25491,N_23084,N_23341);
nand U25492 (N_25492,N_23739,N_20564);
nand U25493 (N_25493,N_23378,N_22540);
nand U25494 (N_25494,N_20484,N_22759);
nand U25495 (N_25495,N_21001,N_24352);
nand U25496 (N_25496,N_21227,N_21811);
or U25497 (N_25497,N_23621,N_21383);
or U25498 (N_25498,N_23957,N_20120);
and U25499 (N_25499,N_21025,N_23410);
nor U25500 (N_25500,N_24432,N_22715);
and U25501 (N_25501,N_20466,N_20698);
nand U25502 (N_25502,N_23835,N_21047);
nor U25503 (N_25503,N_20541,N_20444);
xnor U25504 (N_25504,N_23758,N_24906);
xor U25505 (N_25505,N_20950,N_21804);
xnor U25506 (N_25506,N_24843,N_22731);
or U25507 (N_25507,N_24251,N_24084);
nor U25508 (N_25508,N_21094,N_23216);
or U25509 (N_25509,N_20995,N_24211);
and U25510 (N_25510,N_24491,N_21727);
xnor U25511 (N_25511,N_23065,N_21408);
nand U25512 (N_25512,N_24577,N_22462);
nand U25513 (N_25513,N_23965,N_20516);
nor U25514 (N_25514,N_23310,N_24111);
xnor U25515 (N_25515,N_23826,N_21385);
and U25516 (N_25516,N_23429,N_20255);
nor U25517 (N_25517,N_23900,N_22138);
and U25518 (N_25518,N_24380,N_23272);
nor U25519 (N_25519,N_23276,N_22653);
xor U25520 (N_25520,N_23389,N_21063);
xor U25521 (N_25521,N_21760,N_20267);
and U25522 (N_25522,N_22692,N_23477);
xor U25523 (N_25523,N_21009,N_23192);
nor U25524 (N_25524,N_22773,N_23917);
or U25525 (N_25525,N_24119,N_22132);
nor U25526 (N_25526,N_20744,N_21542);
and U25527 (N_25527,N_24307,N_20302);
nand U25528 (N_25528,N_22506,N_20093);
and U25529 (N_25529,N_21201,N_20076);
or U25530 (N_25530,N_20437,N_21809);
and U25531 (N_25531,N_23961,N_24285);
nand U25532 (N_25532,N_22874,N_24742);
and U25533 (N_25533,N_20642,N_21660);
nor U25534 (N_25534,N_21323,N_23167);
or U25535 (N_25535,N_20622,N_23103);
or U25536 (N_25536,N_21900,N_20041);
nand U25537 (N_25537,N_23743,N_21712);
nor U25538 (N_25538,N_24716,N_21243);
nand U25539 (N_25539,N_23583,N_20080);
and U25540 (N_25540,N_23832,N_23791);
or U25541 (N_25541,N_20400,N_24637);
and U25542 (N_25542,N_22986,N_24353);
or U25543 (N_25543,N_21653,N_22264);
and U25544 (N_25544,N_23061,N_21264);
and U25545 (N_25545,N_20843,N_22184);
nor U25546 (N_25546,N_20293,N_22476);
and U25547 (N_25547,N_23364,N_20274);
xnor U25548 (N_25548,N_23128,N_20097);
and U25549 (N_25549,N_20721,N_20923);
xor U25550 (N_25550,N_21931,N_24827);
nand U25551 (N_25551,N_22599,N_23487);
xnor U25552 (N_25552,N_21616,N_23613);
nor U25553 (N_25553,N_21601,N_20761);
xor U25554 (N_25554,N_21837,N_20822);
and U25555 (N_25555,N_24008,N_24013);
xor U25556 (N_25556,N_21622,N_20175);
and U25557 (N_25557,N_20440,N_21689);
or U25558 (N_25558,N_23147,N_22270);
or U25559 (N_25559,N_20471,N_22963);
nand U25560 (N_25560,N_23127,N_24831);
nor U25561 (N_25561,N_21256,N_22783);
nand U25562 (N_25562,N_23446,N_21621);
nand U25563 (N_25563,N_20056,N_22527);
or U25564 (N_25564,N_22831,N_23981);
or U25565 (N_25565,N_21406,N_20381);
nand U25566 (N_25566,N_22751,N_23353);
and U25567 (N_25567,N_24760,N_20420);
or U25568 (N_25568,N_21326,N_23963);
nor U25569 (N_25569,N_20454,N_20749);
nand U25570 (N_25570,N_23885,N_23908);
nor U25571 (N_25571,N_21410,N_24744);
or U25572 (N_25572,N_20083,N_23811);
and U25573 (N_25573,N_21074,N_24406);
xor U25574 (N_25574,N_24398,N_22397);
and U25575 (N_25575,N_24413,N_20898);
and U25576 (N_25576,N_20199,N_21329);
nor U25577 (N_25577,N_21477,N_20902);
or U25578 (N_25578,N_21921,N_21426);
nand U25579 (N_25579,N_20478,N_23394);
or U25580 (N_25580,N_23385,N_24594);
or U25581 (N_25581,N_23757,N_24110);
nor U25582 (N_25582,N_24096,N_20222);
xnor U25583 (N_25583,N_20708,N_21906);
or U25584 (N_25584,N_24268,N_23528);
nor U25585 (N_25585,N_21774,N_23737);
nand U25586 (N_25586,N_23682,N_20353);
or U25587 (N_25587,N_20263,N_21614);
xor U25588 (N_25588,N_20962,N_22795);
xor U25589 (N_25589,N_23889,N_22762);
or U25590 (N_25590,N_22810,N_23025);
nand U25591 (N_25591,N_21634,N_20998);
nand U25592 (N_25592,N_20714,N_20613);
and U25593 (N_25593,N_20361,N_20718);
nor U25594 (N_25594,N_24687,N_23131);
and U25595 (N_25595,N_24707,N_22850);
or U25596 (N_25596,N_23658,N_20356);
nand U25597 (N_25597,N_24644,N_24730);
or U25598 (N_25598,N_21369,N_24180);
nor U25599 (N_25599,N_21572,N_23140);
or U25600 (N_25600,N_22131,N_23497);
xor U25601 (N_25601,N_21664,N_21117);
and U25602 (N_25602,N_23547,N_21608);
nor U25603 (N_25603,N_24197,N_23767);
nand U25604 (N_25604,N_24265,N_21684);
or U25605 (N_25605,N_20223,N_23178);
xor U25606 (N_25606,N_20048,N_21780);
nand U25607 (N_25607,N_20655,N_21148);
nand U25608 (N_25608,N_20857,N_24661);
xnor U25609 (N_25609,N_24216,N_20511);
and U25610 (N_25610,N_21202,N_21555);
nor U25611 (N_25611,N_22992,N_22280);
and U25612 (N_25612,N_23525,N_23657);
nor U25613 (N_25613,N_20860,N_21874);
xor U25614 (N_25614,N_20021,N_21501);
and U25615 (N_25615,N_22733,N_20262);
or U25616 (N_25616,N_23104,N_22638);
xnor U25617 (N_25617,N_24348,N_23738);
or U25618 (N_25618,N_21854,N_22617);
and U25619 (N_25619,N_21158,N_20968);
and U25620 (N_25620,N_23617,N_20338);
xor U25621 (N_25621,N_24749,N_21827);
xnor U25622 (N_25622,N_24705,N_22220);
nand U25623 (N_25623,N_22251,N_20647);
nand U25624 (N_25624,N_20520,N_21954);
or U25625 (N_25625,N_21662,N_22375);
nor U25626 (N_25626,N_24974,N_22819);
xnor U25627 (N_25627,N_22898,N_23595);
nand U25628 (N_25628,N_24896,N_24043);
nor U25629 (N_25629,N_24442,N_24130);
or U25630 (N_25630,N_23727,N_23822);
nand U25631 (N_25631,N_20094,N_20949);
nand U25632 (N_25632,N_22625,N_20877);
nor U25633 (N_25633,N_20837,N_23203);
nand U25634 (N_25634,N_23148,N_22634);
or U25635 (N_25635,N_23347,N_22811);
nand U25636 (N_25636,N_20807,N_20644);
or U25637 (N_25637,N_24604,N_20391);
xnor U25638 (N_25638,N_23372,N_22784);
and U25639 (N_25639,N_23349,N_24969);
and U25640 (N_25640,N_23176,N_23696);
and U25641 (N_25641,N_24860,N_23611);
nor U25642 (N_25642,N_20004,N_22794);
and U25643 (N_25643,N_21144,N_21208);
or U25644 (N_25644,N_20713,N_23944);
and U25645 (N_25645,N_20127,N_23618);
nand U25646 (N_25646,N_21035,N_23989);
nor U25647 (N_25647,N_20390,N_22799);
nor U25648 (N_25648,N_23988,N_21325);
or U25649 (N_25649,N_23548,N_20706);
nand U25650 (N_25650,N_21893,N_24962);
nand U25651 (N_25651,N_21007,N_20553);
nor U25652 (N_25652,N_23597,N_20417);
or U25653 (N_25653,N_23243,N_24489);
xnor U25654 (N_25654,N_21153,N_20147);
xnor U25655 (N_25655,N_22152,N_21788);
or U25656 (N_25656,N_24979,N_23683);
xor U25657 (N_25657,N_24574,N_20890);
and U25658 (N_25658,N_20947,N_22276);
and U25659 (N_25659,N_21444,N_20166);
nor U25660 (N_25660,N_24218,N_20136);
or U25661 (N_25661,N_21600,N_20791);
xnor U25662 (N_25662,N_22051,N_21095);
nor U25663 (N_25663,N_21218,N_24279);
and U25664 (N_25664,N_21607,N_20696);
or U25665 (N_25665,N_22763,N_23572);
nor U25666 (N_25666,N_23137,N_22873);
nor U25667 (N_25667,N_22110,N_21116);
xor U25668 (N_25668,N_20289,N_23923);
xor U25669 (N_25669,N_21643,N_24578);
xnor U25670 (N_25670,N_21783,N_22073);
nor U25671 (N_25671,N_24683,N_20850);
nor U25672 (N_25672,N_22650,N_23263);
and U25673 (N_25673,N_22036,N_21034);
and U25674 (N_25674,N_23386,N_21569);
and U25675 (N_25675,N_24522,N_24242);
or U25676 (N_25676,N_23852,N_24226);
xor U25677 (N_25677,N_22888,N_20816);
or U25678 (N_25678,N_23476,N_20243);
xnor U25679 (N_25679,N_21726,N_22968);
nor U25680 (N_25680,N_22742,N_20792);
and U25681 (N_25681,N_20458,N_20456);
and U25682 (N_25682,N_23884,N_24532);
nor U25683 (N_25683,N_22858,N_23985);
nor U25684 (N_25684,N_22823,N_20264);
or U25685 (N_25685,N_22365,N_23173);
and U25686 (N_25686,N_24612,N_24435);
nor U25687 (N_25687,N_20330,N_21042);
or U25688 (N_25688,N_21587,N_23913);
nor U25689 (N_25689,N_21756,N_21397);
xor U25690 (N_25690,N_22807,N_21594);
nor U25691 (N_25691,N_21272,N_24427);
nand U25692 (N_25692,N_23195,N_23206);
nand U25693 (N_25693,N_24309,N_20722);
nand U25694 (N_25694,N_24904,N_22266);
and U25695 (N_25695,N_21432,N_20337);
or U25696 (N_25696,N_23144,N_22088);
nor U25697 (N_25697,N_20503,N_21671);
xor U25698 (N_25698,N_22169,N_21976);
nor U25699 (N_25699,N_20070,N_22489);
nand U25700 (N_25700,N_21674,N_21657);
xor U25701 (N_25701,N_24375,N_24942);
nor U25702 (N_25702,N_22701,N_20573);
nand U25703 (N_25703,N_24973,N_24775);
xnor U25704 (N_25704,N_24634,N_21909);
and U25705 (N_25705,N_24162,N_21322);
nor U25706 (N_25706,N_24571,N_23281);
and U25707 (N_25707,N_21564,N_21092);
or U25708 (N_25708,N_23993,N_20399);
nor U25709 (N_25709,N_24523,N_20729);
nand U25710 (N_25710,N_22141,N_20277);
and U25711 (N_25711,N_22326,N_21142);
xor U25712 (N_25712,N_22134,N_24543);
and U25713 (N_25713,N_21249,N_24189);
and U25714 (N_25714,N_21884,N_24653);
and U25715 (N_25715,N_21762,N_22568);
xor U25716 (N_25716,N_20316,N_22645);
nand U25717 (N_25717,N_22834,N_22907);
xor U25718 (N_25718,N_20589,N_22596);
xor U25719 (N_25719,N_24524,N_20191);
nand U25720 (N_25720,N_24959,N_20988);
nand U25721 (N_25721,N_24351,N_22736);
and U25722 (N_25722,N_24438,N_20233);
and U25723 (N_25723,N_24807,N_21057);
nor U25724 (N_25724,N_24339,N_23909);
or U25725 (N_25725,N_23638,N_22379);
nor U25726 (N_25726,N_23541,N_24471);
xnor U25727 (N_25727,N_24895,N_24363);
nor U25728 (N_25728,N_20385,N_22441);
and U25729 (N_25729,N_22308,N_22510);
nor U25730 (N_25730,N_20505,N_23262);
and U25731 (N_25731,N_23800,N_21353);
and U25732 (N_25732,N_20266,N_23318);
or U25733 (N_25733,N_24020,N_24809);
or U25734 (N_25734,N_21591,N_24792);
nand U25735 (N_25735,N_24584,N_20912);
nor U25736 (N_25736,N_22884,N_23987);
or U25737 (N_25737,N_23393,N_23734);
or U25738 (N_25738,N_22433,N_21992);
or U25739 (N_25739,N_22183,N_23448);
nand U25740 (N_25740,N_21831,N_21598);
nor U25741 (N_25741,N_24608,N_21915);
and U25742 (N_25742,N_23845,N_21786);
or U25743 (N_25743,N_23666,N_24202);
nor U25744 (N_25744,N_23751,N_24871);
nand U25745 (N_25745,N_20530,N_24622);
or U25746 (N_25746,N_22578,N_22329);
nor U25747 (N_25747,N_20259,N_20349);
nand U25748 (N_25748,N_21562,N_21508);
and U25749 (N_25749,N_21663,N_21282);
xor U25750 (N_25750,N_20341,N_22028);
nand U25751 (N_25751,N_23020,N_22636);
and U25752 (N_25752,N_20600,N_21529);
nand U25753 (N_25753,N_22411,N_23846);
nor U25754 (N_25754,N_22864,N_23691);
xor U25755 (N_25755,N_20367,N_24821);
or U25756 (N_25756,N_21411,N_24445);
or U25757 (N_25757,N_23934,N_22178);
and U25758 (N_25758,N_20057,N_21247);
xor U25759 (N_25759,N_23274,N_22829);
nand U25760 (N_25760,N_24269,N_20574);
nor U25761 (N_25761,N_21003,N_24715);
xnor U25762 (N_25762,N_21966,N_24695);
and U25763 (N_25763,N_23079,N_24186);
nand U25764 (N_25764,N_24485,N_20835);
xnor U25765 (N_25765,N_22320,N_24278);
nand U25766 (N_25766,N_22393,N_22554);
xnor U25767 (N_25767,N_22133,N_22137);
nor U25768 (N_25768,N_23653,N_22516);
nor U25769 (N_25769,N_24091,N_21602);
or U25770 (N_25770,N_22587,N_23877);
xor U25771 (N_25771,N_23772,N_22719);
xnor U25772 (N_25772,N_22003,N_24618);
nor U25773 (N_25773,N_23375,N_22482);
xnor U25774 (N_25774,N_23893,N_23663);
and U25775 (N_25775,N_20648,N_24992);
and U25776 (N_25776,N_23674,N_20597);
or U25777 (N_25777,N_22300,N_21455);
nor U25778 (N_25778,N_20295,N_22305);
nand U25779 (N_25779,N_23232,N_22442);
or U25780 (N_25780,N_24299,N_21289);
nor U25781 (N_25781,N_23491,N_20621);
or U25782 (N_25782,N_21721,N_23011);
nor U25783 (N_25783,N_24922,N_23060);
nand U25784 (N_25784,N_21418,N_20866);
nor U25785 (N_25785,N_20231,N_21266);
nand U25786 (N_25786,N_24627,N_20922);
nand U25787 (N_25787,N_21901,N_22434);
nand U25788 (N_25788,N_23295,N_22215);
xor U25789 (N_25789,N_21924,N_24295);
nor U25790 (N_25790,N_23075,N_24867);
nor U25791 (N_25791,N_21590,N_24964);
nand U25792 (N_25792,N_22013,N_21168);
xor U25793 (N_25793,N_22918,N_24184);
nor U25794 (N_25794,N_22098,N_24231);
or U25795 (N_25795,N_24869,N_24585);
and U25796 (N_25796,N_23755,N_21113);
nor U25797 (N_25797,N_24390,N_20829);
nand U25798 (N_25798,N_23495,N_24862);
nor U25799 (N_25799,N_22911,N_22032);
xnor U25800 (N_25800,N_21494,N_24006);
or U25801 (N_25801,N_21577,N_22049);
nor U25802 (N_25802,N_21694,N_20138);
nand U25803 (N_25803,N_24528,N_20029);
xor U25804 (N_25804,N_23829,N_21750);
xnor U25805 (N_25805,N_20054,N_23264);
nand U25806 (N_25806,N_23207,N_23507);
xnor U25807 (N_25807,N_24049,N_21384);
and U25808 (N_25808,N_22260,N_23091);
or U25809 (N_25809,N_20679,N_23855);
or U25810 (N_25810,N_23357,N_20084);
nor U25811 (N_25811,N_20183,N_20874);
xnor U25812 (N_25812,N_21106,N_23672);
or U25813 (N_25813,N_20888,N_24763);
nor U25814 (N_25814,N_24420,N_20913);
or U25815 (N_25815,N_23704,N_24473);
xor U25816 (N_25816,N_23685,N_22943);
or U25817 (N_25817,N_23490,N_23117);
xnor U25818 (N_25818,N_21652,N_24911);
nor U25819 (N_25819,N_21899,N_21379);
xnor U25820 (N_25820,N_23786,N_20637);
or U25821 (N_25821,N_21767,N_24616);
nor U25822 (N_25822,N_22099,N_24476);
nor U25823 (N_25823,N_24735,N_21139);
nor U25824 (N_25824,N_20290,N_21228);
or U25825 (N_25825,N_24479,N_24765);
xnor U25826 (N_25826,N_20955,N_23726);
or U25827 (N_25827,N_22207,N_23317);
nor U25828 (N_25828,N_23729,N_22202);
nand U25829 (N_25829,N_24112,N_21259);
or U25830 (N_25830,N_20632,N_20518);
and U25831 (N_25831,N_22857,N_24600);
nand U25832 (N_25832,N_24366,N_23784);
nand U25833 (N_25833,N_21425,N_24302);
nand U25834 (N_25834,N_23110,N_23159);
and U25835 (N_25835,N_24129,N_23742);
xnor U25836 (N_25836,N_20028,N_20182);
nand U25837 (N_25837,N_24168,N_21207);
nand U25838 (N_25838,N_23745,N_21889);
and U25839 (N_25839,N_24157,N_22192);
xnor U25840 (N_25840,N_20389,N_23290);
nand U25841 (N_25841,N_23366,N_23975);
nor U25842 (N_25842,N_24038,N_23472);
nand U25843 (N_25843,N_21235,N_20595);
nor U25844 (N_25844,N_24054,N_21520);
and U25845 (N_25845,N_22680,N_22451);
and U25846 (N_25846,N_20148,N_24460);
xor U25847 (N_25847,N_23062,N_21440);
or U25848 (N_25848,N_21841,N_22917);
and U25849 (N_25849,N_22808,N_22603);
xnor U25850 (N_25850,N_22503,N_22652);
nor U25851 (N_25851,N_22785,N_23442);
nor U25852 (N_25852,N_23291,N_24648);
nor U25853 (N_25853,N_23035,N_23196);
nand U25854 (N_25854,N_21350,N_23022);
nor U25855 (N_25855,N_23873,N_20684);
nand U25856 (N_25856,N_23567,N_20104);
xnor U25857 (N_25857,N_24356,N_22828);
xor U25858 (N_25858,N_21998,N_22331);
xor U25859 (N_25859,N_21761,N_24934);
xnor U25860 (N_25860,N_23897,N_24581);
nand U25861 (N_25861,N_23024,N_24899);
nand U25862 (N_25862,N_23607,N_22893);
xor U25863 (N_25863,N_20467,N_20306);
nor U25864 (N_25864,N_23251,N_23645);
nand U25865 (N_25865,N_24551,N_21104);
nor U25866 (N_25866,N_23108,N_21454);
nand U25867 (N_25867,N_23278,N_21647);
nand U25868 (N_25868,N_24198,N_22975);
and U25869 (N_25869,N_24975,N_22237);
nor U25870 (N_25870,N_20547,N_24588);
nand U25871 (N_25871,N_22350,N_21885);
or U25872 (N_25872,N_22042,N_21796);
xor U25873 (N_25873,N_24201,N_20944);
xor U25874 (N_25874,N_22203,N_22283);
nand U25875 (N_25875,N_22781,N_22194);
xnor U25876 (N_25876,N_21620,N_21503);
nor U25877 (N_25877,N_23982,N_20212);
xnor U25878 (N_25878,N_20973,N_21403);
and U25879 (N_25879,N_24515,N_20146);
nor U25880 (N_25880,N_20847,N_21401);
nor U25881 (N_25881,N_21642,N_21066);
nor U25882 (N_25882,N_22882,N_23590);
nand U25883 (N_25883,N_22899,N_24395);
nand U25884 (N_25884,N_21752,N_22595);
nor U25885 (N_25885,N_20100,N_24335);
and U25886 (N_25886,N_21609,N_23649);
and U25887 (N_25887,N_24736,N_21704);
nor U25888 (N_25888,N_23959,N_24499);
and U25889 (N_25889,N_24235,N_20764);
xnor U25890 (N_25890,N_20360,N_22948);
nand U25891 (N_25891,N_23601,N_21196);
xnor U25892 (N_25892,N_21498,N_20287);
xor U25893 (N_25893,N_24718,N_24536);
or U25894 (N_25894,N_21292,N_22780);
or U25895 (N_25895,N_21824,N_23633);
nand U25896 (N_25896,N_20062,N_22120);
xnor U25897 (N_25897,N_20650,N_20374);
or U25898 (N_25898,N_21446,N_20122);
xnor U25899 (N_25899,N_24257,N_22741);
and U25900 (N_25900,N_22792,N_23785);
and U25901 (N_25901,N_23358,N_23499);
xor U25902 (N_25902,N_23537,N_20325);
xnor U25903 (N_25903,N_20045,N_22030);
nand U25904 (N_25904,N_21245,N_21574);
xnor U25905 (N_25905,N_24912,N_23201);
nor U25906 (N_25906,N_21450,N_22916);
nor U25907 (N_25907,N_21670,N_22518);
nand U25908 (N_25908,N_24089,N_20919);
nand U25909 (N_25909,N_20378,N_21072);
nand U25910 (N_25910,N_23668,N_22635);
and U25911 (N_25911,N_21523,N_22666);
or U25912 (N_25912,N_22352,N_24062);
nand U25913 (N_25913,N_22436,N_21061);
nor U25914 (N_25914,N_24178,N_22156);
xnor U25915 (N_25915,N_22410,N_20340);
nand U25916 (N_25916,N_23213,N_20790);
xor U25917 (N_25917,N_23631,N_21169);
nand U25918 (N_25918,N_24583,N_22841);
and U25919 (N_25919,N_23639,N_22987);
nand U25920 (N_25920,N_20975,N_24468);
nor U25921 (N_25921,N_20149,N_23189);
and U25922 (N_25922,N_24511,N_24848);
nor U25923 (N_25923,N_23656,N_20418);
nor U25924 (N_25924,N_20020,N_22481);
xor U25925 (N_25925,N_21777,N_22148);
or U25926 (N_25926,N_21052,N_23319);
nor U25927 (N_25927,N_20286,N_21157);
and U25928 (N_25928,N_24449,N_21665);
xor U25929 (N_25929,N_24949,N_20483);
nand U25930 (N_25930,N_20669,N_21185);
and U25931 (N_25931,N_24940,N_20802);
or U25932 (N_25932,N_22369,N_24626);
and U25933 (N_25933,N_20241,N_21923);
or U25934 (N_25934,N_21927,N_23722);
and U25935 (N_25935,N_23323,N_21994);
xnor U25936 (N_25936,N_22903,N_24320);
nand U25937 (N_25937,N_22095,N_24945);
nand U25938 (N_25938,N_24337,N_23625);
or U25939 (N_25939,N_22304,N_24947);
xnor U25940 (N_25940,N_23007,N_21154);
or U25941 (N_25941,N_21880,N_21412);
nand U25942 (N_25942,N_21271,N_20319);
xnor U25943 (N_25943,N_21308,N_22342);
xor U25944 (N_25944,N_23840,N_21251);
and U25945 (N_25945,N_21130,N_20275);
nand U25946 (N_25946,N_21825,N_24290);
nor U25947 (N_25947,N_24741,N_20924);
or U25948 (N_25948,N_24148,N_24200);
and U25949 (N_25949,N_24334,N_24518);
and U25950 (N_25950,N_20907,N_23280);
and U25951 (N_25951,N_21152,N_20003);
or U25952 (N_25952,N_23940,N_22052);
and U25953 (N_25953,N_20772,N_22629);
nor U25954 (N_25954,N_20552,N_23681);
nor U25955 (N_25955,N_22897,N_20398);
nor U25956 (N_25956,N_24081,N_21341);
nor U25957 (N_25957,N_22158,N_22445);
and U25958 (N_25958,N_21496,N_23552);
nor U25959 (N_25959,N_22279,N_24493);
or U25960 (N_25960,N_21828,N_23008);
xnor U25961 (N_25961,N_22993,N_24656);
xnor U25962 (N_25962,N_23916,N_21688);
and U25963 (N_25963,N_22439,N_22037);
xnor U25964 (N_25964,N_20116,N_22589);
or U25965 (N_25965,N_21623,N_20034);
nand U25966 (N_25966,N_24534,N_22958);
nand U25967 (N_25967,N_23692,N_24997);
and U25968 (N_25968,N_22092,N_21067);
or U25969 (N_25969,N_20414,N_23146);
xor U25970 (N_25970,N_21024,N_23878);
or U25971 (N_25971,N_22344,N_21434);
nand U25972 (N_25972,N_22647,N_24693);
or U25973 (N_25973,N_23351,N_24022);
and U25974 (N_25974,N_23098,N_23760);
nor U25975 (N_25975,N_21333,N_21160);
xnor U25976 (N_25976,N_24680,N_21054);
or U25977 (N_25977,N_24093,N_23557);
xnor U25978 (N_25978,N_24076,N_21473);
xor U25979 (N_25979,N_24204,N_24392);
or U25980 (N_25980,N_22717,N_21907);
nor U25981 (N_25981,N_20881,N_20559);
xnor U25982 (N_25982,N_22498,N_23861);
nand U25983 (N_25983,N_24919,N_20304);
xor U25984 (N_25984,N_24373,N_21970);
or U25985 (N_25985,N_22620,N_24652);
xnor U25986 (N_25986,N_22338,N_21646);
or U25987 (N_25987,N_20784,N_24488);
and U25988 (N_25988,N_23053,N_20005);
nor U25989 (N_25989,N_24681,N_22776);
nand U25990 (N_25990,N_24173,N_20775);
xnor U25991 (N_25991,N_23717,N_22522);
xnor U25992 (N_25992,N_20408,N_24593);
or U25993 (N_25993,N_20659,N_22706);
or U25994 (N_25994,N_22977,N_20184);
nor U25995 (N_25995,N_24738,N_24751);
or U25996 (N_25996,N_21540,N_22271);
or U25997 (N_25997,N_24219,N_24249);
nand U25998 (N_25998,N_21233,N_23859);
nor U25999 (N_25999,N_23002,N_21424);
or U26000 (N_26000,N_22413,N_21702);
nand U26001 (N_26001,N_20180,N_24282);
and U26002 (N_26002,N_24203,N_20862);
xor U26003 (N_26003,N_22061,N_21295);
nor U26004 (N_26004,N_21102,N_24428);
or U26005 (N_26005,N_23581,N_21749);
nor U26006 (N_26006,N_20114,N_24610);
nor U26007 (N_26007,N_21525,N_21855);
nor U26008 (N_26008,N_21604,N_24469);
xor U26009 (N_26009,N_22185,N_21759);
and U26010 (N_26010,N_23150,N_21378);
and U26011 (N_26011,N_20351,N_21351);
nand U26012 (N_26012,N_20863,N_24726);
or U26013 (N_26013,N_22170,N_24898);
xor U26014 (N_26014,N_24246,N_23779);
and U26015 (N_26015,N_20575,N_22454);
xor U26016 (N_26016,N_22724,N_20782);
or U26017 (N_26017,N_24790,N_22961);
nor U26018 (N_26018,N_21883,N_24050);
or U26019 (N_26019,N_23769,N_22418);
nor U26020 (N_26020,N_24950,N_20410);
nand U26021 (N_26021,N_21904,N_21757);
and U26022 (N_26022,N_24961,N_21729);
or U26023 (N_26023,N_22856,N_21870);
and U26024 (N_26024,N_20766,N_24719);
or U26025 (N_26025,N_23995,N_23143);
xnor U26026 (N_26026,N_22538,N_20900);
and U26027 (N_26027,N_21226,N_20162);
or U26028 (N_26028,N_21580,N_21465);
nand U26029 (N_26029,N_21268,N_22976);
xor U26030 (N_26030,N_21257,N_21083);
or U26031 (N_26031,N_20158,N_23106);
xor U26032 (N_26032,N_23083,N_22105);
nand U26033 (N_26033,N_20732,N_22839);
and U26034 (N_26034,N_21176,N_24410);
or U26035 (N_26035,N_24319,N_21818);
nor U26036 (N_26036,N_24643,N_23764);
nor U26037 (N_26037,N_24876,N_20624);
nor U26038 (N_26038,N_24065,N_22531);
and U26039 (N_26039,N_24819,N_24691);
nor U26040 (N_26040,N_22517,N_22801);
nand U26041 (N_26041,N_24430,N_24999);
xnor U26042 (N_26042,N_21049,N_22536);
nor U26043 (N_26043,N_23371,N_24568);
nand U26044 (N_26044,N_21019,N_23427);
and U26045 (N_26045,N_22745,N_20439);
nand U26046 (N_26046,N_22735,N_22277);
nor U26047 (N_26047,N_22129,N_22236);
and U26048 (N_26048,N_24253,N_23531);
and U26049 (N_26049,N_21164,N_20292);
and U26050 (N_26050,N_24464,N_23842);
or U26051 (N_26051,N_24586,N_20799);
nor U26052 (N_26052,N_23305,N_23430);
xor U26053 (N_26053,N_20329,N_21640);
xor U26054 (N_26054,N_23713,N_22268);
nor U26055 (N_26055,N_20154,N_24721);
nor U26056 (N_26056,N_20619,N_24085);
and U26057 (N_26057,N_20603,N_21606);
and U26058 (N_26058,N_22285,N_24344);
and U26059 (N_26059,N_22872,N_22307);
nor U26060 (N_26060,N_22391,N_20755);
xnor U26061 (N_26061,N_22707,N_20459);
and U26062 (N_26062,N_20424,N_24676);
or U26063 (N_26063,N_20103,N_24458);
xnor U26064 (N_26064,N_22139,N_21695);
and U26065 (N_26065,N_20279,N_24514);
xnor U26066 (N_26066,N_22396,N_23465);
or U26067 (N_26067,N_21214,N_20324);
nor U26068 (N_26068,N_21541,N_21155);
xnor U26069 (N_26069,N_24378,N_23486);
and U26070 (N_26070,N_22109,N_23461);
or U26071 (N_26071,N_20387,N_24777);
or U26072 (N_26072,N_23684,N_24505);
or U26073 (N_26073,N_21084,N_21334);
or U26074 (N_26074,N_22662,N_23233);
and U26075 (N_26075,N_22422,N_22880);
xor U26076 (N_26076,N_23417,N_24549);
nand U26077 (N_26077,N_24734,N_24849);
and U26078 (N_26078,N_21672,N_24155);
or U26079 (N_26079,N_22669,N_22922);
xnor U26080 (N_26080,N_24620,N_20539);
nand U26081 (N_26081,N_21717,N_21979);
or U26082 (N_26082,N_23445,N_22218);
nand U26083 (N_26083,N_24852,N_20586);
nand U26084 (N_26084,N_20945,N_21849);
or U26085 (N_26085,N_23218,N_24349);
and U26086 (N_26086,N_21829,N_24877);
and U26087 (N_26087,N_22316,N_22297);
nor U26088 (N_26088,N_22437,N_21476);
and U26089 (N_26089,N_24646,N_22962);
nand U26090 (N_26090,N_23562,N_24851);
nand U26091 (N_26091,N_22659,N_22298);
nor U26092 (N_26092,N_22765,N_23352);
nand U26093 (N_26093,N_21922,N_20065);
or U26094 (N_26094,N_22594,N_21023);
nor U26095 (N_26095,N_20294,N_22384);
and U26096 (N_26096,N_22957,N_23033);
nor U26097 (N_26097,N_22346,N_23551);
and U26098 (N_26098,N_23401,N_22790);
xnor U26099 (N_26099,N_23516,N_20786);
nand U26100 (N_26100,N_22952,N_23980);
nand U26101 (N_26101,N_24916,N_21028);
nand U26102 (N_26102,N_20085,N_22149);
xnor U26103 (N_26103,N_21474,N_22699);
or U26104 (N_26104,N_24404,N_21358);
and U26105 (N_26105,N_24647,N_20746);
xnor U26106 (N_26106,N_24149,N_20921);
or U26107 (N_26107,N_24855,N_20419);
nand U26108 (N_26108,N_21685,N_21894);
nand U26109 (N_26109,N_22151,N_23133);
and U26110 (N_26110,N_22627,N_20013);
xnor U26111 (N_26111,N_23467,N_20150);
and U26112 (N_26112,N_21965,N_24372);
nand U26113 (N_26113,N_24572,N_22022);
xnor U26114 (N_26114,N_23013,N_21755);
nor U26115 (N_26115,N_22588,N_20633);
nor U26116 (N_26116,N_22425,N_21112);
xor U26117 (N_26117,N_24280,N_24407);
and U26118 (N_26118,N_24382,N_23824);
nand U26119 (N_26119,N_21902,N_23782);
nor U26120 (N_26120,N_24628,N_24672);
nor U26121 (N_26121,N_20594,N_23759);
and U26122 (N_26122,N_23809,N_24552);
and U26123 (N_26123,N_24609,N_21167);
and U26124 (N_26124,N_20710,N_24952);
nor U26125 (N_26125,N_21388,N_24995);
nor U26126 (N_26126,N_24164,N_22775);
and U26127 (N_26127,N_24484,N_20446);
nand U26128 (N_26128,N_21617,N_24664);
nor U26129 (N_26129,N_20335,N_22478);
nor U26130 (N_26130,N_21532,N_21842);
and U26131 (N_26131,N_22994,N_21535);
xnor U26132 (N_26132,N_22423,N_24362);
and U26133 (N_26133,N_21518,N_20963);
nand U26134 (N_26134,N_24915,N_23655);
nor U26135 (N_26135,N_21813,N_23539);
xor U26136 (N_26136,N_24206,N_23257);
and U26137 (N_26137,N_23089,N_23555);
nand U26138 (N_26138,N_20092,N_21423);
or U26139 (N_26139,N_20082,N_22989);
xnor U26140 (N_26140,N_24063,N_22200);
nand U26141 (N_26141,N_22116,N_22906);
and U26142 (N_26142,N_24364,N_22912);
nor U26143 (N_26143,N_22124,N_23844);
or U26144 (N_26144,N_20055,N_21491);
xor U26145 (N_26145,N_23217,N_20583);
nand U26146 (N_26146,N_20787,N_24846);
nand U26147 (N_26147,N_23183,N_24579);
xor U26148 (N_26148,N_24417,N_23049);
nand U26149 (N_26149,N_23390,N_21549);
xor U26150 (N_26150,N_23765,N_22102);
and U26151 (N_26151,N_21431,N_21046);
nor U26152 (N_26152,N_21627,N_21252);
xor U26153 (N_26153,N_21784,N_21656);
nand U26154 (N_26154,N_22700,N_20931);
nand U26155 (N_26155,N_24099,N_23088);
nor U26156 (N_26156,N_24058,N_20246);
nand U26157 (N_26157,N_20190,N_24774);
nor U26158 (N_26158,N_23609,N_22373);
nand U26159 (N_26159,N_20853,N_24674);
xnor U26160 (N_26160,N_21199,N_21463);
and U26161 (N_26161,N_24747,N_22939);
xnor U26162 (N_26162,N_22664,N_20157);
xnor U26163 (N_26163,N_24274,N_23208);
xor U26164 (N_26164,N_24923,N_24779);
nand U26165 (N_26165,N_23947,N_21683);
or U26166 (N_26166,N_20997,N_20219);
and U26167 (N_26167,N_23172,N_23193);
or U26168 (N_26168,N_21556,N_20599);
nand U26169 (N_26169,N_20268,N_23238);
nor U26170 (N_26170,N_21738,N_23673);
xor U26171 (N_26171,N_21270,N_22674);
xor U26172 (N_26172,N_20303,N_20126);
or U26173 (N_26173,N_24220,N_22940);
or U26174 (N_26174,N_20704,N_24958);
or U26175 (N_26175,N_22330,N_23199);
nor U26176 (N_26176,N_21550,N_24475);
and U26177 (N_26177,N_20952,N_20171);
or U26178 (N_26178,N_21838,N_23068);
and U26179 (N_26179,N_22996,N_24908);
nor U26180 (N_26180,N_20379,N_23174);
xor U26181 (N_26181,N_22017,N_20312);
or U26182 (N_26182,N_20585,N_20252);
nor U26183 (N_26183,N_21680,N_24601);
nor U26184 (N_26184,N_20554,N_22879);
and U26185 (N_26185,N_20703,N_22201);
or U26186 (N_26186,N_24623,N_23180);
or U26187 (N_26187,N_22738,N_21209);
or U26188 (N_26188,N_23485,N_20605);
or U26189 (N_26189,N_20667,N_24294);
xor U26190 (N_26190,N_23014,N_23998);
nand U26191 (N_26191,N_21595,N_24245);
xnor U26192 (N_26192,N_24010,N_21336);
or U26193 (N_26193,N_24527,N_21472);
and U26194 (N_26194,N_23973,N_21128);
nor U26195 (N_26195,N_20946,N_23333);
nor U26196 (N_26196,N_23460,N_24370);
and U26197 (N_26197,N_24067,N_23259);
nand U26198 (N_26198,N_20298,N_23076);
xnor U26199 (N_26199,N_23903,N_24980);
nand U26200 (N_26200,N_22547,N_20961);
or U26201 (N_26201,N_20662,N_22757);
xnor U26202 (N_26202,N_24820,N_22671);
nand U26203 (N_26203,N_22555,N_24845);
or U26204 (N_26204,N_24434,N_22217);
nor U26205 (N_26205,N_23205,N_23968);
and U26206 (N_26206,N_21775,N_23471);
or U26207 (N_26207,N_20322,N_20145);
nor U26208 (N_26208,N_21859,N_22548);
nor U26209 (N_26209,N_22960,N_21420);
and U26210 (N_26210,N_24252,N_20533);
or U26211 (N_26211,N_23032,N_24941);
xor U26212 (N_26212,N_22125,N_20770);
nand U26213 (N_26213,N_21963,N_24311);
nand U26214 (N_26214,N_23561,N_20752);
or U26215 (N_26215,N_20938,N_20404);
and U26216 (N_26216,N_21314,N_22895);
nor U26217 (N_26217,N_23612,N_20412);
xnor U26218 (N_26218,N_21720,N_23421);
and U26219 (N_26219,N_24223,N_21055);
nor U26220 (N_26220,N_23574,N_23090);
xnor U26221 (N_26221,N_20727,N_20728);
and U26222 (N_26222,N_20224,N_20842);
and U26223 (N_26223,N_24573,N_20581);
nand U26224 (N_26224,N_20037,N_24880);
or U26225 (N_26225,N_24221,N_24121);
xnor U26226 (N_26226,N_24596,N_22832);
and U26227 (N_26227,N_22607,N_21253);
nand U26228 (N_26228,N_24550,N_20272);
or U26229 (N_26229,N_22153,N_24698);
xor U26230 (N_26230,N_21797,N_23134);
nand U26231 (N_26231,N_22800,N_22323);
xor U26232 (N_26232,N_23282,N_24764);
and U26233 (N_26233,N_23509,N_21744);
or U26234 (N_26234,N_22392,N_20954);
nor U26235 (N_26235,N_24183,N_20101);
or U26236 (N_26236,N_22034,N_22821);
nor U26237 (N_26237,N_24127,N_20480);
nand U26238 (N_26238,N_23396,N_21395);
and U26239 (N_26239,N_23513,N_23549);
and U26240 (N_26240,N_20920,N_20630);
nand U26241 (N_26241,N_20797,N_23783);
nand U26242 (N_26242,N_22753,N_24714);
and U26243 (N_26243,N_22796,N_24803);
xnor U26244 (N_26244,N_21781,N_21346);
and U26245 (N_26245,N_22408,N_22168);
and U26246 (N_26246,N_24441,N_20333);
or U26247 (N_26247,N_24789,N_20485);
and U26248 (N_26248,N_24095,N_23095);
and U26249 (N_26249,N_23241,N_21147);
and U26250 (N_26250,N_20978,N_21240);
or U26251 (N_26251,N_24291,N_20365);
nor U26252 (N_26252,N_22718,N_22836);
xnor U26253 (N_26253,N_20392,N_24347);
nand U26254 (N_26254,N_23197,N_21545);
and U26255 (N_26255,N_21429,N_23279);
and U26256 (N_26256,N_21957,N_21619);
nor U26257 (N_26257,N_23253,N_21511);
xor U26258 (N_26258,N_24272,N_24926);
and U26259 (N_26259,N_24517,N_23292);
nand U26260 (N_26260,N_21981,N_23866);
or U26261 (N_26261,N_24697,N_22846);
and U26262 (N_26262,N_22177,N_24472);
xnor U26263 (N_26263,N_20882,N_23724);
or U26264 (N_26264,N_21527,N_24181);
and U26265 (N_26265,N_22507,N_23667);
nand U26266 (N_26266,N_21060,N_22459);
xor U26267 (N_26267,N_23066,N_21839);
or U26268 (N_26268,N_20540,N_21413);
or U26269 (N_26269,N_23636,N_22552);
nand U26270 (N_26270,N_23640,N_21935);
nand U26271 (N_26271,N_22998,N_20051);
or U26272 (N_26272,N_23398,N_21363);
xnor U26273 (N_26273,N_20588,N_20543);
or U26274 (N_26274,N_23679,N_21364);
xnor U26275 (N_26275,N_20309,N_20981);
xnor U26276 (N_26276,N_23834,N_24224);
and U26277 (N_26277,N_24128,N_21905);
nor U26278 (N_26278,N_24270,N_21330);
nor U26279 (N_26279,N_23339,N_23420);
or U26280 (N_26280,N_20270,N_23426);
or U26281 (N_26281,N_20623,N_20508);
nand U26282 (N_26282,N_23676,N_22598);
nor U26283 (N_26283,N_21438,N_21661);
and U26284 (N_26284,N_24872,N_21399);
nand U26285 (N_26285,N_20328,N_21563);
and U26286 (N_26286,N_23204,N_22245);
xor U26287 (N_26287,N_20990,N_22809);
nand U26288 (N_26288,N_20558,N_21133);
xnor U26289 (N_26289,N_21170,N_20332);
nand U26290 (N_26290,N_23964,N_24028);
nand U26291 (N_26291,N_24766,N_21558);
nor U26292 (N_26292,N_20726,N_23604);
nor U26293 (N_26293,N_21593,N_21366);
or U26294 (N_26294,N_21165,N_20072);
and U26295 (N_26295,N_23670,N_21810);
nor U26296 (N_26296,N_20036,N_23960);
nand U26297 (N_26297,N_22341,N_22479);
nand U26298 (N_26298,N_20536,N_21394);
or U26299 (N_26299,N_23454,N_22631);
xnor U26300 (N_26300,N_24931,N_24448);
nor U26301 (N_26301,N_22472,N_23170);
and U26302 (N_26302,N_23919,N_24179);
and U26303 (N_26303,N_24217,N_22720);
and U26304 (N_26304,N_24663,N_21499);
nor U26305 (N_26305,N_22233,N_20993);
nand U26306 (N_26306,N_21173,N_24752);
nor U26307 (N_26307,N_23480,N_21161);
nor U26308 (N_26308,N_22761,N_21573);
or U26309 (N_26309,N_23587,N_22078);
or U26310 (N_26310,N_24797,N_20499);
xnor U26311 (N_26311,N_22359,N_24383);
nand U26312 (N_26312,N_21517,N_23736);
and U26313 (N_26313,N_24436,N_24972);
and U26314 (N_26314,N_23787,N_20682);
and U26315 (N_26315,N_24597,N_22866);
or U26316 (N_26316,N_23069,N_24385);
nor U26317 (N_26317,N_23122,N_22691);
nand U26318 (N_26318,N_24072,N_20382);
xor U26319 (N_26319,N_21773,N_22532);
nand U26320 (N_26320,N_24810,N_22675);
nand U26321 (N_26321,N_22685,N_21903);
and U26322 (N_26322,N_24642,N_22537);
and U26323 (N_26323,N_22278,N_23792);
or U26324 (N_26324,N_21949,N_22708);
or U26325 (N_26325,N_21229,N_22409);
nand U26326 (N_26326,N_20423,N_20976);
or U26327 (N_26327,N_24669,N_22891);
and U26328 (N_26328,N_24746,N_24844);
and U26329 (N_26329,N_23544,N_24654);
xnor U26330 (N_26330,N_21486,N_20606);
nor U26331 (N_26331,N_24881,N_23748);
xnor U26332 (N_26332,N_23151,N_22188);
and U26333 (N_26333,N_20571,N_21140);
xor U26334 (N_26334,N_23892,N_22561);
or U26335 (N_26335,N_23484,N_23698);
nand U26336 (N_26336,N_24833,N_20652);
nand U26337 (N_26337,N_22004,N_21197);
xor U26338 (N_26338,N_22926,N_24987);
nand U26339 (N_26339,N_21392,N_20769);
and U26340 (N_26340,N_20069,N_20192);
or U26341 (N_26341,N_21821,N_23455);
xor U26342 (N_26342,N_24447,N_23926);
nor U26343 (N_26343,N_20284,N_22591);
and U26344 (N_26344,N_22654,N_24679);
and U26345 (N_26345,N_22354,N_23042);
nor U26346 (N_26346,N_24925,N_22835);
and U26347 (N_26347,N_21300,N_24260);
nand U26348 (N_26348,N_22232,N_21795);
or U26349 (N_26349,N_23858,N_21076);
nor U26350 (N_26350,N_24857,N_22562);
xor U26351 (N_26351,N_21972,N_24910);
and U26352 (N_26352,N_21754,N_21787);
nand U26353 (N_26353,N_20833,N_20798);
nor U26354 (N_26354,N_21851,N_21651);
nand U26355 (N_26355,N_24800,N_22317);
and U26356 (N_26356,N_23226,N_20549);
or U26357 (N_26357,N_22545,N_23773);
xor U26358 (N_26358,N_23402,N_22429);
nand U26359 (N_26359,N_23864,N_21122);
and U26360 (N_26360,N_20854,N_24921);
xnor U26361 (N_26361,N_21127,N_21051);
xor U26362 (N_26362,N_24811,N_22113);
and U26363 (N_26363,N_24131,N_21823);
and U26364 (N_26364,N_22771,N_24355);
xnor U26365 (N_26365,N_21415,N_23373);
nand U26366 (N_26366,N_21017,N_23966);
nor U26367 (N_26367,N_20098,N_23540);
nand U26368 (N_26368,N_22908,N_21571);
or U26369 (N_26369,N_21890,N_21872);
nor U26370 (N_26370,N_20486,N_21254);
or U26371 (N_26371,N_24412,N_21659);
or U26372 (N_26372,N_24060,N_24498);
nand U26373 (N_26373,N_24426,N_23030);
xnor U26374 (N_26374,N_20665,N_21039);
or U26375 (N_26375,N_24048,N_22467);
xnor U26376 (N_26376,N_21255,N_24582);
nor U26377 (N_26377,N_23074,N_22597);
or U26378 (N_26378,N_22486,N_20808);
or U26379 (N_26379,N_23111,N_22900);
or U26380 (N_26380,N_21219,N_22564);
and U26381 (N_26381,N_21583,N_20282);
xor U26382 (N_26382,N_24000,N_23756);
nand U26383 (N_26383,N_20388,N_22949);
xnor U26384 (N_26384,N_21059,N_23408);
nand U26385 (N_26385,N_24136,N_23435);
and U26386 (N_26386,N_20959,N_23139);
or U26387 (N_26387,N_23021,N_21331);
and U26388 (N_26388,N_20596,N_23177);
nand U26389 (N_26389,N_23234,N_20634);
xor U26390 (N_26390,N_23246,N_20081);
nor U26391 (N_26391,N_21189,N_21993);
nand U26392 (N_26392,N_22068,N_24930);
xor U26393 (N_26393,N_23932,N_23078);
xnor U26394 (N_26394,N_21740,N_22085);
xnor U26395 (N_26395,N_22162,N_21381);
or U26396 (N_26396,N_22851,N_24023);
nor U26397 (N_26397,N_24558,N_20375);
and U26398 (N_26398,N_22797,N_20253);
nor U26399 (N_26399,N_21320,N_21045);
or U26400 (N_26400,N_22764,N_21280);
nor U26401 (N_26401,N_24768,N_22492);
nor U26402 (N_26402,N_23862,N_21193);
and U26403 (N_26403,N_22814,N_24419);
xnor U26404 (N_26404,N_23946,N_23324);
or U26405 (N_26405,N_21978,N_23268);
nand U26406 (N_26406,N_22644,N_22493);
and U26407 (N_26407,N_24165,N_22859);
xor U26408 (N_26408,N_24755,N_22228);
or U26409 (N_26409,N_22754,N_20757);
nand U26410 (N_26410,N_21706,N_23788);
nor U26411 (N_26411,N_20828,N_22130);
and U26412 (N_26412,N_21387,N_22197);
nor U26413 (N_26413,N_20725,N_20887);
xor U26414 (N_26414,N_22128,N_21983);
or U26415 (N_26415,N_22936,N_23220);
nand U26416 (N_26416,N_20124,N_23031);
or U26417 (N_26417,N_24657,N_20334);
and U26418 (N_26418,N_24396,N_20783);
and U26419 (N_26419,N_20812,N_22027);
nand U26420 (N_26420,N_21183,N_21419);
nor U26421 (N_26421,N_20514,N_21710);
nor U26422 (N_26422,N_23297,N_21632);
xnor U26423 (N_26423,N_21635,N_24055);
and U26424 (N_26424,N_23255,N_20731);
and U26425 (N_26425,N_21012,N_24225);
xor U26426 (N_26426,N_22311,N_24977);
nor U26427 (N_26427,N_24903,N_24955);
or U26428 (N_26428,N_20762,N_22750);
and U26429 (N_26429,N_21785,N_21589);
and U26430 (N_26430,N_24160,N_20768);
nand U26431 (N_26431,N_24379,N_20815);
nor U26432 (N_26432,N_22546,N_22487);
nand U26433 (N_26433,N_24386,N_24793);
xor U26434 (N_26434,N_20283,N_21206);
nand U26435 (N_26435,N_20203,N_23040);
nor U26436 (N_26436,N_21666,N_23794);
xnor U26437 (N_26437,N_22573,N_21764);
xor U26438 (N_26438,N_20817,N_21930);
and U26439 (N_26439,N_23876,N_20314);
nor U26440 (N_26440,N_23605,N_24377);
nor U26441 (N_26441,N_22450,N_24324);
nand U26442 (N_26442,N_24592,N_22016);
and U26443 (N_26443,N_20011,N_20865);
xor U26444 (N_26444,N_20996,N_23413);
nand U26445 (N_26445,N_20576,N_21008);
xor U26446 (N_26446,N_24815,N_21510);
xnor U26447 (N_26447,N_23483,N_24835);
xnor U26448 (N_26448,N_21951,N_21808);
and U26449 (N_26449,N_22530,N_20506);
nor U26450 (N_26450,N_24630,N_24965);
xor U26451 (N_26451,N_23853,N_20811);
xor U26452 (N_26452,N_23242,N_23830);
xor U26453 (N_26453,N_23977,N_22633);
nor U26454 (N_26454,N_24575,N_20492);
or U26455 (N_26455,N_23294,N_21613);
nor U26456 (N_26456,N_24737,N_21313);
xnor U26457 (N_26457,N_24712,N_20448);
and U26458 (N_26458,N_23087,N_21293);
xnor U26459 (N_26459,N_24645,N_21290);
and U26460 (N_26460,N_22195,N_24670);
xor U26461 (N_26461,N_23009,N_20280);
or U26462 (N_26462,N_24753,N_23029);
nand U26463 (N_26463,N_24907,N_22744);
xnor U26464 (N_26464,N_21405,N_23314);
nand U26465 (N_26465,N_22155,N_22063);
nor U26466 (N_26466,N_23436,N_24650);
or U26467 (N_26467,N_20914,N_20740);
or U26468 (N_26468,N_22006,N_20026);
nor U26469 (N_26469,N_21136,N_24357);
nor U26470 (N_26470,N_20415,N_20053);
nand U26471 (N_26471,N_24816,N_22452);
and U26472 (N_26472,N_20736,N_22394);
nor U26473 (N_26473,N_22500,N_20134);
nand U26474 (N_26474,N_21934,N_23316);
or U26475 (N_26475,N_20777,N_23126);
xor U26476 (N_26476,N_23660,N_23047);
nand U26477 (N_26477,N_22386,N_23493);
or U26478 (N_26478,N_22777,N_20569);
nand U26479 (N_26479,N_20256,N_23553);
and U26480 (N_26480,N_23416,N_23776);
nand U26481 (N_26481,N_21037,N_23839);
nor U26482 (N_26482,N_24520,N_21044);
or U26483 (N_26483,N_22301,N_22097);
and U26484 (N_26484,N_22070,N_21714);
nand U26485 (N_26485,N_22937,N_20693);
nor U26486 (N_26486,N_22769,N_21987);
xor U26487 (N_26487,N_22966,N_20654);
or U26488 (N_26488,N_22416,N_23918);
and U26489 (N_26489,N_21497,N_23313);
and U26490 (N_26490,N_24710,N_21328);
nor U26491 (N_26491,N_22883,N_22242);
nor U26492 (N_26492,N_20173,N_22542);
nor U26493 (N_26493,N_23346,N_20323);
nand U26494 (N_26494,N_23214,N_24529);
and U26495 (N_26495,N_20479,N_24207);
and U26496 (N_26496,N_20421,N_24166);
or U26497 (N_26497,N_20926,N_24277);
nand U26498 (N_26498,N_23578,N_24939);
and U26499 (N_26499,N_23836,N_24393);
and U26500 (N_26500,N_22923,N_21748);
nand U26501 (N_26501,N_22901,N_22550);
nand U26502 (N_26502,N_20810,N_23245);
or U26503 (N_26503,N_23418,N_22174);
xor U26504 (N_26504,N_22135,N_23797);
nor U26505 (N_26505,N_24275,N_24090);
nor U26506 (N_26506,N_20163,N_23086);
xnor U26507 (N_26507,N_22321,N_22015);
nand U26508 (N_26508,N_21848,N_23584);
nor U26509 (N_26509,N_23141,N_21551);
nand U26510 (N_26510,N_21376,N_22204);
and U26511 (N_26511,N_20393,N_20868);
and U26512 (N_26512,N_22009,N_20977);
and U26513 (N_26513,N_20869,N_21162);
and U26514 (N_26514,N_20238,N_22240);
or U26515 (N_26515,N_24411,N_23718);
nor U26516 (N_26516,N_22661,N_24935);
xnor U26517 (N_26517,N_23181,N_22855);
and U26518 (N_26518,N_24983,N_23942);
nand U26519 (N_26519,N_20331,N_20310);
nor U26520 (N_26520,N_23403,N_24678);
and U26521 (N_26521,N_24624,N_21439);
and U26522 (N_26522,N_23712,N_21579);
or U26523 (N_26523,N_24421,N_24243);
and U26524 (N_26524,N_23976,N_24553);
or U26525 (N_26525,N_20685,N_23063);
and U26526 (N_26526,N_23984,N_23586);
or U26527 (N_26527,N_24883,N_22100);
and U26528 (N_26528,N_23950,N_24859);
and U26529 (N_26529,N_24124,N_23322);
and U26530 (N_26530,N_24617,N_24512);
and U26531 (N_26531,N_22333,N_20651);
xnor U26532 (N_26532,N_23992,N_23520);
xor U26533 (N_26533,N_21421,N_23922);
or U26534 (N_26534,N_21349,N_24539);
nor U26535 (N_26535,N_22585,N_20470);
and U26536 (N_26536,N_23546,N_21815);
and U26537 (N_26537,N_22065,N_22984);
and U26538 (N_26538,N_22826,N_23915);
nand U26539 (N_26539,N_22672,N_23327);
or U26540 (N_26540,N_22845,N_21537);
nand U26541 (N_26541,N_24104,N_24261);
nor U26542 (N_26542,N_24556,N_21955);
or U26543 (N_26543,N_23457,N_24783);
nor U26544 (N_26544,N_21230,N_21345);
xor U26545 (N_26545,N_21262,N_24776);
xor U26546 (N_26546,N_21236,N_22688);
and U26547 (N_26547,N_21475,N_24535);
xor U26548 (N_26548,N_24847,N_23414);
nand U26549 (N_26549,N_24450,N_24122);
and U26550 (N_26550,N_23603,N_20567);
or U26551 (N_26551,N_24689,N_21086);
nand U26552 (N_26552,N_20687,N_20517);
nor U26553 (N_26553,N_23345,N_21560);
and U26554 (N_26554,N_21505,N_23300);
xnor U26555 (N_26555,N_21362,N_22020);
nor U26556 (N_26556,N_24429,N_21225);
and U26557 (N_26557,N_23034,N_20664);
nor U26558 (N_26558,N_20141,N_20507);
and U26559 (N_26559,N_24563,N_20542);
nand U26560 (N_26560,N_21043,N_21911);
nor U26561 (N_26561,N_24150,N_22057);
or U26562 (N_26562,N_21371,N_20123);
nand U26563 (N_26563,N_21488,N_22101);
and U26564 (N_26564,N_22827,N_23907);
xor U26565 (N_26565,N_21402,N_24824);
and U26566 (N_26566,N_22093,N_22368);
nand U26567 (N_26567,N_22614,N_24740);
or U26568 (N_26568,N_24516,N_20039);
or U26569 (N_26569,N_23591,N_20705);
nand U26570 (N_26570,N_23795,N_20582);
nand U26571 (N_26571,N_23971,N_22480);
nand U26572 (N_26572,N_21565,N_21267);
xor U26573 (N_26573,N_24135,N_20537);
and U26574 (N_26574,N_21521,N_23221);
or U26575 (N_26575,N_20578,N_22729);
or U26576 (N_26576,N_21747,N_23802);
or U26577 (N_26577,N_21493,N_20897);
or U26578 (N_26578,N_22502,N_20061);
nand U26579 (N_26579,N_22892,N_23702);
or U26580 (N_26580,N_21568,N_21305);
and U26581 (N_26581,N_23451,N_21132);
nor U26582 (N_26582,N_21223,N_22182);
nand U26583 (N_26583,N_21137,N_23145);
and U26584 (N_26584,N_22226,N_21597);
nand U26585 (N_26585,N_23077,N_22755);
or U26586 (N_26586,N_24271,N_22023);
or U26587 (N_26587,N_21471,N_20929);
xnor U26588 (N_26588,N_20618,N_20611);
xor U26589 (N_26589,N_21065,N_20636);
nand U26590 (N_26590,N_23200,N_20697);
or U26591 (N_26591,N_21131,N_24477);
nor U26592 (N_26592,N_24863,N_22144);
and U26593 (N_26593,N_22056,N_20189);
and U26594 (N_26594,N_21174,N_21753);
nor U26595 (N_26595,N_20880,N_21141);
nand U26596 (N_26596,N_23043,N_20364);
nand U26597 (N_26597,N_21374,N_22115);
xor U26598 (N_26598,N_23194,N_22743);
nand U26599 (N_26599,N_22231,N_22281);
and U26600 (N_26600,N_23825,N_21952);
and U26601 (N_26601,N_23419,N_20545);
and U26602 (N_26602,N_23187,N_23168);
nor U26603 (N_26603,N_24537,N_22325);
or U26604 (N_26604,N_24123,N_21588);
xnor U26605 (N_26605,N_23026,N_22059);
and U26606 (N_26606,N_21596,N_23629);
and U26607 (N_26607,N_22108,N_21273);
nor U26608 (N_26608,N_24011,N_22529);
nor U26609 (N_26609,N_24365,N_24281);
xnor U26610 (N_26610,N_23952,N_21108);
nor U26611 (N_26611,N_23162,N_21644);
and U26612 (N_26612,N_24748,N_20178);
nor U26613 (N_26613,N_20602,N_23431);
or U26614 (N_26614,N_22067,N_21816);
nor U26615 (N_26615,N_21276,N_24036);
nor U26616 (N_26616,N_23677,N_21390);
xnor U26617 (N_26617,N_20407,N_20871);
and U26618 (N_26618,N_23974,N_22415);
xnor U26619 (N_26619,N_24953,N_22272);
xnor U26620 (N_26620,N_24018,N_24425);
or U26621 (N_26621,N_20177,N_23659);
xnor U26622 (N_26622,N_23706,N_22889);
and U26623 (N_26623,N_24154,N_20064);
nand U26624 (N_26624,N_23569,N_20590);
xnor U26625 (N_26625,N_22610,N_23464);
or U26626 (N_26626,N_24208,N_22345);
xnor U26627 (N_26627,N_20164,N_20980);
nand U26628 (N_26628,N_24892,N_20673);
nor U26629 (N_26629,N_24106,N_20504);
nor U26630 (N_26630,N_22676,N_24040);
and U26631 (N_26631,N_22525,N_23566);
nor U26632 (N_26632,N_23054,N_21279);
or U26633 (N_26633,N_22611,N_24662);
xor U26634 (N_26634,N_23160,N_22909);
nor U26635 (N_26635,N_23678,N_22167);
and U26636 (N_26636,N_20519,N_20425);
xnor U26637 (N_26637,N_23006,N_23123);
nor U26638 (N_26638,N_21678,N_21435);
and U26639 (N_26639,N_20102,N_20523);
or U26640 (N_26640,N_22041,N_23365);
nand U26641 (N_26641,N_21281,N_20346);
nand U26642 (N_26642,N_23343,N_22211);
xor U26643 (N_26643,N_20824,N_23293);
or U26644 (N_26644,N_23887,N_24273);
or U26645 (N_26645,N_23851,N_22072);
nor U26646 (N_26646,N_20911,N_24254);
nor U26647 (N_26647,N_24446,N_24704);
nand U26648 (N_26648,N_22274,N_24033);
and U26649 (N_26649,N_21805,N_23945);
xnor U26650 (N_26650,N_20509,N_22558);
nand U26651 (N_26651,N_21675,N_23367);
or U26652 (N_26652,N_24388,N_22136);
and U26653 (N_26653,N_22581,N_20301);
xor U26654 (N_26654,N_22190,N_21178);
nand U26655 (N_26655,N_20909,N_21500);
xor U26656 (N_26656,N_21461,N_20071);
and U26657 (N_26657,N_21649,N_24012);
nor U26658 (N_26658,N_23406,N_23377);
xnor U26659 (N_26659,N_21220,N_23500);
and U26660 (N_26660,N_21016,N_20515);
nor U26661 (N_26661,N_23073,N_20000);
xnor U26662 (N_26662,N_20521,N_24140);
nand U26663 (N_26663,N_23671,N_24232);
or U26664 (N_26664,N_21667,N_23244);
or U26665 (N_26665,N_23620,N_24343);
or U26666 (N_26666,N_24007,N_24101);
or U26667 (N_26667,N_24114,N_20715);
xnor U26668 (N_26668,N_22511,N_24724);
xor U26669 (N_26669,N_20273,N_23166);
and U26670 (N_26670,N_24146,N_20964);
nand U26671 (N_26671,N_24416,N_23662);
xor U26672 (N_26672,N_22842,N_24795);
or U26673 (N_26673,N_24531,N_21975);
nor U26674 (N_26674,N_22663,N_22490);
or U26675 (N_26675,N_22609,N_24014);
nand U26676 (N_26676,N_21327,N_22616);
nand U26677 (N_26677,N_23523,N_21728);
xnor U26678 (N_26678,N_24507,N_24913);
nor U26679 (N_26679,N_23019,N_22639);
nor U26680 (N_26680,N_24966,N_21462);
nor U26681 (N_26681,N_22928,N_24205);
or U26682 (N_26682,N_23978,N_21715);
or U26683 (N_26683,N_22327,N_20631);
nor U26684 (N_26684,N_21343,N_21146);
nand U26685 (N_26685,N_21487,N_21650);
nand U26686 (N_26686,N_24402,N_20017);
nor U26687 (N_26687,N_22867,N_23725);
and U26688 (N_26688,N_23596,N_24839);
xor U26689 (N_26689,N_23093,N_23296);
xnor U26690 (N_26690,N_21673,N_24264);
and U26691 (N_26691,N_20617,N_20242);
nor U26692 (N_26692,N_21150,N_24957);
or U26693 (N_26693,N_23719,N_20591);
xor U26694 (N_26694,N_23354,N_23564);
or U26695 (N_26695,N_24565,N_20125);
xnor U26696 (N_26696,N_22112,N_24865);
xnor U26697 (N_26697,N_22458,N_21386);
xnor U26698 (N_26698,N_21393,N_24823);
nor U26699 (N_26699,N_22324,N_20906);
xor U26700 (N_26700,N_21840,N_21724);
xnor U26701 (N_26701,N_24262,N_21910);
nor U26702 (N_26702,N_21794,N_23956);
nor U26703 (N_26703,N_24152,N_23326);
or U26704 (N_26704,N_22064,N_21917);
xor U26705 (N_26705,N_22224,N_20638);
or U26706 (N_26706,N_22173,N_23812);
nand U26707 (N_26707,N_22347,N_22683);
and U26708 (N_26708,N_24418,N_21516);
xor U26709 (N_26709,N_24703,N_24500);
nor U26710 (N_26710,N_21679,N_22205);
xor U26711 (N_26711,N_20885,N_23508);
xor U26712 (N_26712,N_23447,N_22955);
or U26713 (N_26713,N_24496,N_21959);
or U26714 (N_26714,N_21618,N_24874);
and U26715 (N_26715,N_24814,N_22582);
xnor U26716 (N_26716,N_20690,N_23770);
xnor U26717 (N_26717,N_23249,N_22399);
or U26718 (N_26718,N_20561,N_23927);
and U26719 (N_26719,N_21624,N_23912);
and U26720 (N_26720,N_21933,N_22475);
xor U26721 (N_26721,N_24345,N_24948);
or U26722 (N_26722,N_23215,N_21407);
nor U26723 (N_26723,N_22402,N_22514);
xor U26724 (N_26724,N_20615,N_20984);
or U26725 (N_26725,N_20087,N_20674);
nor U26726 (N_26726,N_23359,N_20608);
or U26727 (N_26727,N_20535,N_24685);
and U26728 (N_26728,N_22953,N_21539);
and U26729 (N_26729,N_22267,N_22407);
nor U26730 (N_26730,N_22579,N_20550);
nand U26731 (N_26731,N_24991,N_21967);
or U26732 (N_26732,N_20160,N_22118);
nand U26733 (N_26733,N_21561,N_20205);
nor U26734 (N_26734,N_20524,N_24310);
and U26735 (N_26735,N_24754,N_21830);
xor U26736 (N_26736,N_23754,N_22786);
nor U26737 (N_26737,N_21791,N_24918);
and U26738 (N_26738,N_24891,N_24602);
nor U26739 (N_26739,N_24641,N_24041);
and U26740 (N_26740,N_23920,N_23624);
and U26741 (N_26741,N_20078,N_24361);
and U26742 (N_26742,N_21125,N_20967);
or U26743 (N_26743,N_23568,N_21309);
nand U26744 (N_26744,N_21603,N_22535);
nand U26745 (N_26745,N_21939,N_23482);
or U26746 (N_26746,N_22166,N_21040);
nor U26747 (N_26747,N_24143,N_23198);
nand U26748 (N_26748,N_24784,N_20411);
nor U26749 (N_26749,N_22920,N_24329);
nor U26750 (N_26750,N_22443,N_20641);
xnor U26751 (N_26751,N_22448,N_24606);
nand U26752 (N_26752,N_24772,N_24659);
xnor U26753 (N_26753,N_21263,N_22008);
xnor U26754 (N_26754,N_24508,N_21852);
and U26755 (N_26755,N_23114,N_23184);
and U26756 (N_26756,N_24561,N_21416);
nor U26757 (N_26757,N_20352,N_21460);
and U26758 (N_26758,N_21436,N_24990);
and U26759 (N_26759,N_24788,N_21945);
nand U26760 (N_26760,N_23686,N_21820);
nor U26761 (N_26761,N_23573,N_20903);
nor U26762 (N_26762,N_22941,N_21101);
and U26763 (N_26763,N_21080,N_22651);
and U26764 (N_26764,N_22896,N_23309);
xnor U26765 (N_26765,N_20265,N_20681);
and U26766 (N_26766,N_24213,N_24403);
or U26767 (N_26767,N_20373,N_23015);
or U26768 (N_26768,N_21737,N_22533);
nand U26769 (N_26769,N_20089,N_23107);
nand U26770 (N_26770,N_23506,N_24882);
and U26771 (N_26771,N_21731,N_22871);
xor U26772 (N_26772,N_22618,N_22241);
nand U26773 (N_26773,N_24885,N_21984);
xnor U26774 (N_26774,N_22696,N_21000);
xor U26775 (N_26775,N_20763,N_24276);
xnor U26776 (N_26776,N_24566,N_21524);
and U26777 (N_26777,N_21718,N_23637);
xnor U26778 (N_26778,N_24487,N_20038);
nand U26779 (N_26779,N_20214,N_20107);
xnor U26780 (N_26780,N_24951,N_21389);
xor U26781 (N_26781,N_23252,N_23577);
nor U26782 (N_26782,N_20639,N_22071);
xor U26783 (N_26783,N_20476,N_20027);
and U26784 (N_26784,N_22768,N_20635);
xnor U26785 (N_26785,N_23699,N_22504);
nand U26786 (N_26786,N_21746,N_21177);
xor U26787 (N_26787,N_20427,N_21078);
nor U26788 (N_26788,N_24711,N_23924);
and U26789 (N_26789,N_20023,N_22690);
nand U26790 (N_26790,N_22890,N_20489);
nand U26791 (N_26791,N_20119,N_21417);
and U26792 (N_26792,N_23841,N_24660);
nor U26793 (N_26793,N_20735,N_22818);
xnor U26794 (N_26794,N_21509,N_22447);
or U26795 (N_26795,N_24694,N_23910);
xnor U26796 (N_26796,N_21317,N_21430);
or U26797 (N_26797,N_23136,N_21126);
or U26798 (N_26798,N_22460,N_22689);
or U26799 (N_26799,N_23356,N_21504);
xor U26800 (N_26800,N_20966,N_21956);
nand U26801 (N_26801,N_22196,N_22302);
nor U26802 (N_26802,N_20889,N_21002);
nand U26803 (N_26803,N_22362,N_21611);
or U26804 (N_26804,N_20016,N_24255);
or U26805 (N_26805,N_23130,N_24873);
and U26806 (N_26806,N_23102,N_21771);
and U26807 (N_26807,N_21194,N_23598);
xor U26808 (N_26808,N_22189,N_22512);
nor U26809 (N_26809,N_20359,N_24151);
nand U26810 (N_26810,N_23240,N_20457);
xnor U26811 (N_26811,N_20321,N_23474);
nor U26812 (N_26812,N_23092,N_21936);
nor U26813 (N_26813,N_24633,N_20814);
xnor U26814 (N_26814,N_22929,N_22075);
nor U26815 (N_26815,N_24894,N_23936);
xnor U26816 (N_26816,N_22656,N_20747);
nor U26817 (N_26817,N_24452,N_24177);
or U26818 (N_26818,N_21693,N_22577);
xnor U26819 (N_26819,N_21318,N_21294);
xnor U26820 (N_26820,N_20271,N_22593);
and U26821 (N_26821,N_20620,N_20992);
or U26822 (N_26822,N_21048,N_23701);
nor U26823 (N_26823,N_21554,N_20915);
xnor U26824 (N_26824,N_23057,N_24758);
and U26825 (N_26825,N_20153,N_24796);
nor U26826 (N_26826,N_24059,N_20152);
nand U26827 (N_26827,N_20501,N_24590);
or U26828 (N_26828,N_23744,N_24828);
or U26829 (N_26829,N_20050,N_22328);
or U26830 (N_26830,N_20748,N_23505);
nand U26831 (N_26831,N_21447,N_22915);
nand U26832 (N_26832,N_21109,N_22011);
nor U26833 (N_26833,N_22838,N_24544);
nor U26834 (N_26834,N_21637,N_20688);
nand U26835 (N_26835,N_24306,N_21224);
and U26836 (N_26836,N_23331,N_20826);
and U26837 (N_26837,N_23270,N_23082);
nand U26838 (N_26838,N_21570,N_23070);
nand U26839 (N_26839,N_20730,N_23449);
and U26840 (N_26840,N_21182,N_23433);
and U26841 (N_26841,N_22332,N_20653);
xor U26842 (N_26842,N_20592,N_21091);
nand U26843 (N_26843,N_20463,N_24331);
and U26844 (N_26844,N_21519,N_21156);
xor U26845 (N_26845,N_21700,N_20143);
or U26846 (N_26846,N_24806,N_22254);
xnor U26847 (N_26847,N_23016,N_22414);
and U26848 (N_26848,N_24519,N_24397);
or U26849 (N_26849,N_20989,N_21575);
xnor U26850 (N_26850,N_21817,N_24706);
or U26851 (N_26851,N_22262,N_22885);
xor U26852 (N_26852,N_21302,N_20969);
nor U26853 (N_26853,N_22263,N_23705);
nor U26854 (N_26854,N_23780,N_22714);
and U26855 (N_26855,N_22944,N_20468);
xnor U26856 (N_26856,N_24298,N_23921);
or U26857 (N_26857,N_22466,N_22726);
nand U26858 (N_26858,N_21210,N_21845);
and U26859 (N_26859,N_23321,N_24303);
and U26860 (N_26860,N_20363,N_22127);
nor U26861 (N_26861,N_23059,N_22711);
or U26862 (N_26862,N_23817,N_23931);
nor U26863 (N_26863,N_23790,N_21997);
nor U26864 (N_26864,N_24175,N_23690);
nor U26865 (N_26865,N_22010,N_22420);
nand U26866 (N_26866,N_24799,N_24325);
or U26867 (N_26867,N_24682,N_22524);
nor U26868 (N_26868,N_23642,N_21789);
or U26869 (N_26869,N_23850,N_20442);
nor U26870 (N_26870,N_21733,N_21414);
or U26871 (N_26871,N_22160,N_23055);
or U26872 (N_26872,N_23432,N_20789);
nor U26873 (N_26873,N_22914,N_22951);
and U26874 (N_26874,N_21886,N_23953);
or U26875 (N_26875,N_22074,N_22150);
and U26876 (N_26876,N_21021,N_23789);
or U26877 (N_26877,N_22180,N_21835);
and U26878 (N_26878,N_21159,N_22982);
nand U26879 (N_26879,N_23287,N_22465);
nor U26880 (N_26880,N_22640,N_23814);
xnor U26881 (N_26881,N_21514,N_24686);
or U26882 (N_26882,N_21312,N_22356);
xnor U26883 (N_26883,N_24234,N_20901);
and U26884 (N_26884,N_23542,N_23165);
nor U26885 (N_26885,N_20348,N_23044);
xor U26886 (N_26886,N_24897,N_24192);
or U26887 (N_26887,N_24256,N_21871);
and U26888 (N_26888,N_23212,N_20151);
or U26889 (N_26889,N_24971,N_20527);
xnor U26890 (N_26890,N_24956,N_23269);
nor U26891 (N_26891,N_23440,N_23188);
or U26892 (N_26892,N_21020,N_20121);
nand U26893 (N_26893,N_24030,N_20831);
nor U26894 (N_26894,N_21869,N_22965);
nand U26895 (N_26895,N_23052,N_21668);
xor U26896 (N_26896,N_20435,N_24879);
xnor U26897 (N_26897,N_20711,N_24214);
xnor U26898 (N_26898,N_22294,N_21481);
or U26899 (N_26899,N_20413,N_24156);
nor U26900 (N_26900,N_20823,N_22398);
or U26901 (N_26901,N_24905,N_23301);
and U26902 (N_26902,N_21244,N_22694);
and U26903 (N_26903,N_24301,N_22026);
xor U26904 (N_26904,N_22499,N_22837);
xnor U26905 (N_26905,N_23504,N_22494);
xor U26906 (N_26906,N_23606,N_24482);
or U26907 (N_26907,N_23594,N_22613);
or U26908 (N_26908,N_20497,N_23288);
and U26909 (N_26909,N_20236,N_21630);
and U26910 (N_26910,N_22355,N_24194);
or U26911 (N_26911,N_24172,N_24853);
and U26912 (N_26912,N_23622,N_20803);
or U26913 (N_26913,N_22501,N_20140);
nand U26914 (N_26914,N_20299,N_21286);
xor U26915 (N_26915,N_24920,N_20675);
and U26916 (N_26916,N_20778,N_21705);
nand U26917 (N_26917,N_20318,N_24133);
and U26918 (N_26918,N_23363,N_23894);
xnor U26919 (N_26919,N_21485,N_24890);
or U26920 (N_26920,N_24389,N_22400);
and U26921 (N_26921,N_20610,N_20161);
or U26922 (N_26922,N_21348,N_23925);
or U26923 (N_26923,N_20771,N_22050);
and U26924 (N_26924,N_23289,N_20200);
nor U26925 (N_26925,N_20108,N_20904);
xnor U26926 (N_26926,N_22945,N_20670);
or U26927 (N_26927,N_22570,N_24615);
xnor U26928 (N_26928,N_22403,N_24804);
nand U26929 (N_26929,N_20009,N_21211);
xnor U26930 (N_26930,N_24936,N_21213);
nand U26931 (N_26931,N_21929,N_21950);
and U26932 (N_26932,N_23383,N_24709);
and U26933 (N_26933,N_22243,N_23041);
or U26934 (N_26934,N_23710,N_22508);
nand U26935 (N_26935,N_22697,N_23036);
nand U26936 (N_26936,N_22069,N_23694);
and U26937 (N_26937,N_21763,N_22919);
and U26938 (N_26938,N_24560,N_22252);
nand U26939 (N_26939,N_21832,N_24850);
nand U26940 (N_26940,N_21238,N_20060);
nand U26941 (N_26941,N_22019,N_20572);
and U26942 (N_26942,N_20449,N_21015);
nor U26943 (N_26943,N_22140,N_24120);
nand U26944 (N_26944,N_20891,N_23005);
and U26945 (N_26945,N_20237,N_20079);
and U26946 (N_26946,N_20692,N_22370);
or U26947 (N_26947,N_22457,N_20788);
or U26948 (N_26948,N_24548,N_24884);
xnor U26949 (N_26949,N_22014,N_24651);
and U26950 (N_26950,N_23600,N_21261);
nand U26951 (N_26951,N_22248,N_24761);
xnor U26952 (N_26952,N_20249,N_24360);
xnor U26953 (N_26953,N_23337,N_20686);
xnor U26954 (N_26954,N_24631,N_20884);
nand U26955 (N_26955,N_20933,N_24842);
nand U26956 (N_26956,N_24266,N_21187);
nand U26957 (N_26957,N_20825,N_21868);
and U26958 (N_26958,N_22740,N_20472);
xnor U26959 (N_26959,N_21347,N_22039);
nand U26960 (N_26960,N_21467,N_23038);
and U26961 (N_26961,N_22622,N_24996);
or U26962 (N_26962,N_24141,N_22497);
nor U26963 (N_26963,N_20239,N_22289);
xnor U26964 (N_26964,N_22682,N_21822);
or U26965 (N_26965,N_24132,N_21005);
and U26966 (N_26966,N_24188,N_23211);
nand U26967 (N_26967,N_21947,N_22206);
and U26968 (N_26968,N_24480,N_24454);
xor U26969 (N_26969,N_22360,N_20229);
xnor U26970 (N_26970,N_23338,N_24666);
or U26971 (N_26971,N_23010,N_21908);
nand U26972 (N_26972,N_21882,N_24510);
nor U26973 (N_26973,N_22314,N_20451);
and U26974 (N_26974,N_24079,N_23100);
and U26975 (N_26975,N_21636,N_23810);
or U26976 (N_26976,N_22526,N_22089);
and U26977 (N_26977,N_23510,N_24103);
nand U26978 (N_26978,N_20668,N_20794);
and U26979 (N_26979,N_21776,N_22574);
and U26980 (N_26980,N_24100,N_20109);
nand U26981 (N_26981,N_21231,N_22983);
xnor U26982 (N_26982,N_24621,N_22978);
or U26983 (N_26983,N_22702,N_22608);
xor U26984 (N_26984,N_21248,N_22315);
or U26985 (N_26985,N_23306,N_20513);
or U26986 (N_26986,N_23428,N_23132);
xor U26987 (N_26987,N_24917,N_22722);
nor U26988 (N_26988,N_24503,N_22081);
and U26989 (N_26989,N_22322,N_24459);
or U26990 (N_26990,N_23979,N_23731);
xnor U26991 (N_26991,N_23661,N_24051);
and U26992 (N_26992,N_21698,N_23619);
or U26993 (N_26993,N_22935,N_24837);
or U26994 (N_26994,N_20207,N_22772);
and U26995 (N_26995,N_20849,N_21742);
xnor U26996 (N_26996,N_22875,N_23890);
nor U26997 (N_26997,N_21029,N_22791);
or U26998 (N_26998,N_20986,N_20168);
nand U26999 (N_26999,N_23868,N_20852);
nand U27000 (N_27000,N_20305,N_20226);
nand U27001 (N_27001,N_22852,N_23163);
nor U27002 (N_27002,N_22833,N_21974);
nor U27003 (N_27003,N_24117,N_23708);
or U27004 (N_27004,N_24077,N_20851);
and U27005 (N_27005,N_20144,N_23149);
nand U27006 (N_27006,N_20260,N_24613);
or U27007 (N_27007,N_23320,N_23158);
nand U27008 (N_27008,N_23424,N_22925);
and U27009 (N_27009,N_22844,N_23185);
nor U27010 (N_27010,N_21013,N_24731);
nor U27011 (N_27011,N_20300,N_22389);
and U27012 (N_27012,N_24440,N_24658);
or U27013 (N_27013,N_23828,N_22760);
xnor U27014 (N_27014,N_23171,N_24391);
nor U27015 (N_27015,N_23202,N_21241);
nor U27016 (N_27016,N_21149,N_24163);
xor U27017 (N_27017,N_20958,N_20473);
nor U27018 (N_27018,N_20879,N_21807);
and U27019 (N_27019,N_22031,N_20137);
or U27020 (N_27020,N_24603,N_20801);
nor U27021 (N_27021,N_21913,N_20870);
xor U27022 (N_27022,N_21953,N_24976);
nand U27023 (N_27023,N_24193,N_22477);
nor U27024 (N_27024,N_20462,N_24982);
or U27025 (N_27025,N_24998,N_20844);
and U27026 (N_27026,N_21064,N_24635);
or U27027 (N_27027,N_22464,N_22214);
or U27028 (N_27028,N_20202,N_21538);
nor U27029 (N_27029,N_24688,N_21916);
or U27030 (N_27030,N_22805,N_21713);
nand U27031 (N_27031,N_22756,N_23466);
and U27032 (N_27032,N_21466,N_22967);
nand U27033 (N_27033,N_21739,N_24094);
nand U27034 (N_27034,N_20244,N_23225);
xnor U27035 (N_27035,N_20565,N_22235);
nor U27036 (N_27036,N_24743,N_20209);
xnor U27037 (N_27037,N_23796,N_21716);
nand U27038 (N_27038,N_22847,N_21586);
xor U27039 (N_27039,N_23051,N_20939);
xor U27040 (N_27040,N_24671,N_22142);
or U27041 (N_27041,N_21802,N_20819);
xnor U27042 (N_27042,N_23746,N_22083);
nor U27043 (N_27043,N_21356,N_23224);
xor U27044 (N_27044,N_22843,N_24813);
and U27045 (N_27045,N_20999,N_22739);
nor U27046 (N_27046,N_20464,N_23229);
and U27047 (N_27047,N_24832,N_24781);
or U27048 (N_27048,N_21203,N_23037);
and U27049 (N_27049,N_20063,N_20738);
nor U27050 (N_27050,N_20433,N_22255);
nor U27051 (N_27051,N_24717,N_20370);
and U27052 (N_27052,N_24466,N_21303);
and U27053 (N_27053,N_22822,N_21515);
or U27054 (N_27054,N_22930,N_23532);
nand U27055 (N_27055,N_24227,N_23860);
xnor U27056 (N_27056,N_22630,N_22767);
and U27057 (N_27057,N_20475,N_21391);
and U27058 (N_27058,N_21355,N_20213);
nor U27059 (N_27059,N_20609,N_21625);
nand U27060 (N_27060,N_21864,N_24504);
nand U27061 (N_27061,N_21138,N_24902);
xor U27062 (N_27062,N_22973,N_20461);
xnor U27063 (N_27063,N_22619,N_24161);
or U27064 (N_27064,N_22947,N_22725);
nor U27065 (N_27065,N_21451,N_22946);
or U27066 (N_27066,N_24032,N_20106);
and U27067 (N_27067,N_24723,N_22942);
and U27068 (N_27068,N_21283,N_20131);
and U27069 (N_27069,N_24387,N_23627);
xnor U27070 (N_27070,N_21205,N_20556);
nor U27071 (N_27071,N_23986,N_20896);
nor U27072 (N_27072,N_21926,N_21843);
nand U27073 (N_27073,N_21982,N_23582);
nor U27074 (N_27074,N_24288,N_22779);
nor U27075 (N_27075,N_21502,N_21098);
or U27076 (N_27076,N_22543,N_23958);
nor U27077 (N_27077,N_22076,N_21701);
nor U27078 (N_27078,N_20925,N_23857);
and U27079 (N_27079,N_20864,N_21985);
or U27080 (N_27080,N_20734,N_23911);
xor U27081 (N_27081,N_20075,N_24954);
xnor U27082 (N_27082,N_24782,N_23843);
nor U27083 (N_27083,N_24547,N_22357);
nor U27084 (N_27084,N_21398,N_21368);
or U27085 (N_27085,N_21548,N_23750);
nand U27086 (N_27086,N_23896,N_21709);
or U27087 (N_27087,N_22921,N_21881);
xor U27088 (N_27088,N_23815,N_23728);
nor U27089 (N_27089,N_21382,N_21918);
nand U27090 (N_27090,N_24474,N_23804);
and U27091 (N_27091,N_20185,N_24354);
nor U27092 (N_27092,N_20409,N_23879);
nor U27093 (N_27093,N_24886,N_20805);
xnor U27094 (N_27094,N_24580,N_21988);
or U27095 (N_27095,N_23271,N_21793);
and U27096 (N_27096,N_24988,N_22250);
xor U27097 (N_27097,N_21986,N_20598);
xnor U27098 (N_27098,N_24673,N_24125);
xnor U27099 (N_27099,N_24700,N_24690);
nand U27100 (N_27100,N_22473,N_23863);
and U27101 (N_27101,N_24944,N_20441);
nor U27102 (N_27102,N_21339,N_24924);
and U27103 (N_27103,N_22122,N_21734);
xor U27104 (N_27104,N_21692,N_23962);
nand U27105 (N_27105,N_20712,N_20196);
nor U27106 (N_27106,N_22096,N_23395);
nor U27107 (N_27107,N_22520,N_22551);
nor U27108 (N_27108,N_23721,N_24258);
and U27109 (N_27109,N_22667,N_22904);
nor U27110 (N_27110,N_21861,N_23340);
and U27111 (N_27111,N_24336,N_24929);
or U27112 (N_27112,N_23819,N_22234);
and U27113 (N_27113,N_23115,N_24401);
nor U27114 (N_27114,N_24082,N_22803);
xor U27115 (N_27115,N_22969,N_20676);
xor U27116 (N_27116,N_21361,N_23469);
or U27117 (N_27117,N_23955,N_23740);
nand U27118 (N_27118,N_22605,N_24589);
or U27119 (N_27119,N_24769,N_23648);
xor U27120 (N_27120,N_21526,N_22488);
xor U27121 (N_27121,N_23626,N_23610);
or U27122 (N_27122,N_21812,N_24465);
nor U27123 (N_27123,N_22249,N_24212);
nand U27124 (N_27124,N_22592,N_23838);
xnor U27125 (N_27125,N_24470,N_24244);
or U27126 (N_27126,N_20544,N_23570);
nor U27127 (N_27127,N_23874,N_22080);
xnor U27128 (N_27128,N_22601,N_23273);
and U27129 (N_27129,N_23362,N_24086);
nand U27130 (N_27130,N_23774,N_24701);
nor U27131 (N_27131,N_23254,N_23283);
nor U27132 (N_27132,N_23948,N_21242);
and U27133 (N_27133,N_20767,N_22444);
or U27134 (N_27134,N_20204,N_22219);
or U27135 (N_27135,N_23423,N_24729);
or U27136 (N_27136,N_21449,N_20941);
nand U27137 (N_27137,N_22932,N_22959);
or U27138 (N_27138,N_20096,N_23641);
nand U27139 (N_27139,N_23680,N_20186);
nand U27140 (N_27140,N_21478,N_24293);
or U27141 (N_27141,N_21357,N_21506);
and U27142 (N_27142,N_21847,N_21553);
nand U27143 (N_27143,N_22824,N_23169);
and U27144 (N_27144,N_24333,N_24818);
nand U27145 (N_27145,N_20118,N_21445);
nor U27146 (N_27146,N_24861,N_23813);
or U27147 (N_27147,N_20386,N_23161);
or U27148 (N_27148,N_22709,N_24817);
nand U27149 (N_27149,N_22505,N_20834);
and U27150 (N_27150,N_20661,N_22210);
nand U27151 (N_27151,N_21344,N_21340);
and U27152 (N_27152,N_23599,N_22830);
or U27153 (N_27153,N_23284,N_22660);
and U27154 (N_27154,N_23135,N_24986);
or U27155 (N_27155,N_20066,N_24240);
xnor U27156 (N_27156,N_23543,N_24250);
nand U27157 (N_27157,N_20058,N_24367);
nor U27158 (N_27158,N_22704,N_22848);
nor U27159 (N_27159,N_23652,N_20577);
nor U27160 (N_27160,N_21079,N_22628);
and U27161 (N_27161,N_20091,N_20227);
and U27162 (N_27162,N_22541,N_23391);
nand U27163 (N_27163,N_21100,N_20948);
xor U27164 (N_27164,N_23634,N_23616);
and U27165 (N_27165,N_21707,N_22273);
nor U27166 (N_27166,N_20002,N_20974);
xor U27167 (N_27167,N_21070,N_20155);
or U27168 (N_27168,N_23558,N_24330);
nand U27169 (N_27169,N_23388,N_20719);
xor U27170 (N_27170,N_24170,N_22412);
nand U27171 (N_27171,N_21612,N_20528);
xor U27172 (N_27172,N_20677,N_24525);
nand U27173 (N_27173,N_20671,N_21172);
nand U27174 (N_27174,N_23646,N_22406);
nand U27175 (N_27175,N_22956,N_24812);
nand U27176 (N_27176,N_24909,N_23999);
and U27177 (N_27177,N_24780,N_21360);
nand U27178 (N_27178,N_23434,N_24080);
xor U27179 (N_27179,N_23444,N_23902);
nor U27180 (N_27180,N_22862,N_23374);
and U27181 (N_27181,N_20840,N_20942);
nor U27182 (N_27182,N_20657,N_24019);
nand U27183 (N_27183,N_21103,N_20689);
xor U27184 (N_27184,N_23589,N_22970);
nor U27185 (N_27185,N_20015,N_23521);
xnor U27186 (N_27186,N_22782,N_21082);
xor U27187 (N_27187,N_22495,N_20447);
or U27188 (N_27188,N_23425,N_21124);
or U27189 (N_27189,N_23511,N_23261);
xnor U27190 (N_27190,N_24092,N_20110);
nor U27191 (N_27191,N_24767,N_22746);
nand U27192 (N_27192,N_24798,N_22641);
and U27193 (N_27193,N_23219,N_23125);
or U27194 (N_27194,N_24073,N_23256);
xnor U27195 (N_27195,N_22077,N_20167);
nand U27196 (N_27196,N_23906,N_21332);
and U27197 (N_27197,N_23179,N_22383);
and U27198 (N_27198,N_20500,N_22902);
xor U27199 (N_27199,N_20032,N_23462);
nor U27200 (N_27200,N_24786,N_20859);
nand U27201 (N_27201,N_21615,N_20460);
xor U27202 (N_27202,N_21605,N_22813);
nor U27203 (N_27203,N_23524,N_23545);
nor U27204 (N_27204,N_20403,N_22427);
and U27205 (N_27205,N_24521,N_21433);
nor U27206 (N_27206,N_20979,N_20916);
nand U27207 (N_27207,N_23000,N_22566);
or U27208 (N_27208,N_22649,N_22385);
or U27209 (N_27209,N_23376,N_24045);
and U27210 (N_27210,N_21654,N_23560);
or U27211 (N_27211,N_22387,N_20873);
or U27212 (N_27212,N_23458,N_20534);
nor U27213 (N_27213,N_22580,N_20090);
or U27214 (N_27214,N_23720,N_21483);
nor U27215 (N_27215,N_24414,N_23632);
and U27216 (N_27216,N_21038,N_20362);
nand U27217 (N_27217,N_22339,N_20563);
xnor U27218 (N_27218,N_23452,N_22559);
or U27219 (N_27219,N_24875,N_22007);
or U27220 (N_27220,N_20201,N_20883);
nor U27221 (N_27221,N_24027,N_20396);
or U27222 (N_27222,N_22094,N_22703);
and U27223 (N_27223,N_24239,N_22265);
and U27224 (N_27224,N_20487,N_20169);
or U27225 (N_27225,N_21866,N_20643);
and U27226 (N_27226,N_24042,N_24409);
nor U27227 (N_27227,N_21964,N_21306);
or U27228 (N_27228,N_24900,N_21878);
xnor U27229 (N_27229,N_21533,N_24259);
and U27230 (N_27230,N_22766,N_22863);
xor U27231 (N_27231,N_23554,N_21316);
nand U27232 (N_27232,N_21639,N_24068);
nand U27233 (N_27233,N_22774,N_24722);
or U27234 (N_27234,N_20159,N_23623);
xnor U27235 (N_27235,N_21198,N_24494);
xnor U27236 (N_27236,N_21310,N_20445);
or U27237 (N_27237,N_24914,N_24167);
nor U27238 (N_27238,N_22988,N_21258);
xnor U27239 (N_27239,N_20395,N_23302);
nand U27240 (N_27240,N_23848,N_22974);
or U27241 (N_27241,N_20800,N_23529);
and U27242 (N_27242,N_23411,N_20832);
and U27243 (N_27243,N_24035,N_24292);
nor U27244 (N_27244,N_21990,N_20014);
xor U27245 (N_27245,N_21311,N_21470);
and U27246 (N_27246,N_23191,N_24629);
and U27247 (N_27247,N_23867,N_22927);
xor U27248 (N_27248,N_22376,N_21443);
and U27249 (N_27249,N_23700,N_22712);
and U27250 (N_27250,N_24889,N_22705);
nor U27251 (N_27251,N_23933,N_22491);
or U27252 (N_27252,N_22789,N_21354);
nor U27253 (N_27253,N_23299,N_24943);
nand U27254 (N_27254,N_24371,N_22275);
nor U27255 (N_27255,N_22193,N_20371);
nor U27256 (N_27256,N_24422,N_21097);
nand U27257 (N_27257,N_20928,N_22886);
or U27258 (N_27258,N_21180,N_21723);
and U27259 (N_27259,N_22485,N_24185);
nor U27260 (N_27260,N_23286,N_23494);
xor U27261 (N_27261,N_22910,N_20716);
nand U27262 (N_27262,N_23899,N_24424);
nand U27263 (N_27263,N_21836,N_24002);
nor U27264 (N_27264,N_24182,N_20568);
nor U27265 (N_27265,N_22216,N_21239);
and U27266 (N_27266,N_20086,N_20040);
and U27267 (N_27267,N_23439,N_24267);
nor U27268 (N_27268,N_20477,N_21766);
nand U27269 (N_27269,N_20012,N_23512);
xor U27270 (N_27270,N_23094,N_20327);
or U27271 (N_27271,N_21221,N_20917);
nand U27272 (N_27272,N_20354,N_24856);
and U27273 (N_27273,N_20893,N_23882);
xnor U27274 (N_27274,N_20453,N_22456);
xnor U27275 (N_27275,N_24108,N_22001);
and U27276 (N_27276,N_22175,N_23715);
and U27277 (N_27277,N_24305,N_23239);
xnor U27278 (N_27278,N_24968,N_22147);
or U27279 (N_27279,N_20380,N_21960);
and U27280 (N_27280,N_24513,N_24801);
or U27281 (N_27281,N_20430,N_21769);
and U27282 (N_27282,N_24016,N_22111);
or U27283 (N_27283,N_21962,N_24932);
nor U27284 (N_27284,N_24794,N_21708);
nor U27285 (N_27285,N_23951,N_20502);
and U27286 (N_27286,N_23519,N_22778);
or U27287 (N_27287,N_24540,N_20315);
and U27288 (N_27288,N_23669,N_22665);
and U27289 (N_27289,N_20142,N_21119);
nor U27290 (N_27290,N_20678,N_24326);
or U27291 (N_27291,N_23422,N_22367);
and U27292 (N_27292,N_22222,N_23635);
xnor U27293 (N_27293,N_24209,N_21879);
and U27294 (N_27294,N_21050,N_21269);
xor U27295 (N_27295,N_22253,N_21898);
nor U27296 (N_27296,N_22247,N_22295);
nand U27297 (N_27297,N_20756,N_21995);
and U27298 (N_27298,N_21772,N_20666);
and U27299 (N_27299,N_21971,N_24057);
and U27300 (N_27300,N_20181,N_22364);
nor U27301 (N_27301,N_24187,N_23355);
nand U27302 (N_27302,N_20215,N_24981);
or U27303 (N_27303,N_23816,N_22812);
nand U27304 (N_27304,N_21014,N_20510);
xor U27305 (N_27305,N_21856,N_24394);
or U27306 (N_27306,N_20210,N_22991);
nand U27307 (N_27307,N_20257,N_23265);
nor U27308 (N_27308,N_24126,N_20129);
nor U27309 (N_27309,N_21991,N_24037);
xor U27310 (N_27310,N_24074,N_24567);
xnor U27311 (N_27311,N_20482,N_24888);
nand U27312 (N_27312,N_23058,N_22054);
xnor U27313 (N_27313,N_21296,N_22870);
and U27314 (N_27314,N_24739,N_21195);
or U27315 (N_27315,N_21968,N_24598);
or U27316 (N_27316,N_21484,N_20031);
or U27317 (N_27317,N_23580,N_20876);
nor U27318 (N_27318,N_23384,N_20006);
xnor U27319 (N_27319,N_20758,N_21989);
and U27320 (N_27320,N_23248,N_21741);
nand U27321 (N_27321,N_24559,N_24878);
and U27322 (N_27322,N_24237,N_20932);
and U27323 (N_27323,N_21031,N_23807);
and U27324 (N_27324,N_22658,N_22238);
and U27325 (N_27325,N_23250,N_21200);
and U27326 (N_27326,N_21456,N_23793);
xor U27327 (N_27327,N_23039,N_21631);
and U27328 (N_27328,N_21372,N_22213);
or U27329 (N_27329,N_22748,N_24191);
xor U27330 (N_27330,N_24836,N_24462);
or U27331 (N_27331,N_21375,N_22474);
xor U27332 (N_27332,N_21192,N_23409);
nand U27333 (N_27333,N_21288,N_21973);
and U27334 (N_27334,N_22637,N_23536);
xnor U27335 (N_27335,N_23941,N_24457);
nand U27336 (N_27336,N_21512,N_24639);
nand U27337 (N_27337,N_21743,N_24868);
xor U27338 (N_27338,N_21920,N_24732);
xor U27339 (N_27339,N_21770,N_21338);
xor U27340 (N_27340,N_22995,N_21204);
and U27341 (N_27341,N_22468,N_22372);
xor U27342 (N_27342,N_21687,N_20366);
nor U27343 (N_27343,N_20971,N_21896);
and U27344 (N_27344,N_23820,N_20431);
xor U27345 (N_27345,N_20261,N_23387);
nand U27346 (N_27346,N_23983,N_20646);
or U27347 (N_27347,N_22172,N_20793);
or U27348 (N_27348,N_22062,N_24400);
xor U27349 (N_27349,N_21111,N_21468);
and U27350 (N_27350,N_20983,N_24026);
nand U27351 (N_27351,N_23210,N_22246);
nor U27352 (N_27352,N_23304,N_22583);
xnor U27353 (N_27353,N_20269,N_22258);
or U27354 (N_27354,N_20809,N_21077);
nand U27355 (N_27355,N_20247,N_21337);
nor U27356 (N_27356,N_24284,N_21961);
xnor U27357 (N_27357,N_20077,N_24834);
or U27358 (N_27358,N_20432,N_21145);
and U27359 (N_27359,N_23888,N_20927);
nor U27360 (N_27360,N_23004,N_20672);
nor U27361 (N_27361,N_20720,N_24667);
or U27362 (N_27362,N_21996,N_20394);
or U27363 (N_27363,N_20839,N_21058);
and U27364 (N_27364,N_21877,N_23303);
xor U27365 (N_27365,N_20042,N_22256);
xnor U27366 (N_27366,N_21010,N_22528);
xor U27367 (N_27367,N_21676,N_20426);
nand U27368 (N_27368,N_23693,N_24546);
nor U27369 (N_27369,N_20680,N_20707);
or U27370 (N_27370,N_20008,N_24492);
nor U27371 (N_27371,N_22931,N_23085);
xnor U27372 (N_27372,N_23689,N_21105);
or U27373 (N_27373,N_20753,N_21826);
nand U27374 (N_27374,N_20113,N_22343);
nand U27375 (N_27375,N_22455,N_22390);
nor U27376 (N_27376,N_23714,N_22815);
xnor U27377 (N_27377,N_22449,N_23475);
or U27378 (N_27378,N_24625,N_23749);
and U27379 (N_27379,N_22395,N_24497);
xor U27380 (N_27380,N_20818,N_21457);
xnor U27381 (N_27381,N_22556,N_20133);
or U27382 (N_27382,N_23332,N_20867);
nor U27383 (N_27383,N_21536,N_23675);
and U27384 (N_27384,N_22954,N_24720);
or U27385 (N_27385,N_23222,N_22563);
and U27386 (N_27386,N_20010,N_20049);
xnor U27387 (N_27387,N_20115,N_20285);
nor U27388 (N_27388,N_22293,N_22964);
nor U27389 (N_27389,N_20628,N_20043);
or U27390 (N_27390,N_21409,N_24021);
nand U27391 (N_27391,N_21179,N_20095);
and U27392 (N_27392,N_23350,N_24314);
or U27393 (N_27393,N_23382,N_24283);
nor U27394 (N_27394,N_24870,N_21566);
and U27395 (N_27395,N_22861,N_22713);
nand U27396 (N_27396,N_22012,N_20821);
and U27397 (N_27397,N_22572,N_22282);
xnor U27398 (N_27398,N_20258,N_20311);
nor U27399 (N_27399,N_22887,N_20813);
nand U27400 (N_27400,N_23247,N_21291);
and U27401 (N_27401,N_22816,N_20174);
and U27402 (N_27402,N_22114,N_21191);
nor U27403 (N_27403,N_22404,N_20165);
and U27404 (N_27404,N_20538,N_24938);
nor U27405 (N_27405,N_22024,N_20128);
nor U27406 (N_27406,N_20625,N_20218);
nand U27407 (N_27407,N_20297,N_24338);
nor U27408 (N_27408,N_21641,N_20007);
xor U27409 (N_27409,N_24822,N_22084);
xor U27410 (N_27410,N_24866,N_24137);
xnor U27411 (N_27411,N_24046,N_24595);
nand U27412 (N_27412,N_23515,N_22126);
nand U27413 (N_27413,N_23285,N_21396);
or U27414 (N_27414,N_20001,N_20765);
nand U27415 (N_27415,N_23307,N_24083);
and U27416 (N_27416,N_21699,N_22825);
nand U27417 (N_27417,N_21319,N_21400);
and U27418 (N_27418,N_20841,N_20156);
nand U27419 (N_27419,N_20024,N_24118);
and U27420 (N_27420,N_23833,N_21171);
nand U27421 (N_27421,N_20607,N_21888);
and U27422 (N_27422,N_24005,N_24841);
or U27423 (N_27423,N_20555,N_21373);
nand U27424 (N_27424,N_23709,N_21284);
or U27425 (N_27425,N_24088,N_22938);
xor U27426 (N_27426,N_22227,N_23872);
or U27427 (N_27427,N_21948,N_22950);
nor U27428 (N_27428,N_21377,N_24928);
or U27429 (N_27429,N_23081,N_20526);
nand U27430 (N_27430,N_23400,N_23312);
nand U27431 (N_27431,N_23501,N_20179);
or U27432 (N_27432,N_21803,N_20498);
nand U27433 (N_27433,N_23763,N_24004);
and U27434 (N_27434,N_24145,N_23741);
and U27435 (N_27435,N_23407,N_20856);
xnor U27436 (N_27436,N_22584,N_22261);
nand U27437 (N_27437,N_23118,N_24805);
and U27438 (N_27438,N_24770,N_24169);
nand U27439 (N_27439,N_20982,N_23665);
nand U27440 (N_27440,N_21285,N_24985);
nand U27441 (N_27441,N_23854,N_24056);
or U27442 (N_27442,N_24541,N_23488);
nor U27443 (N_27443,N_23938,N_24826);
nor U27444 (N_27444,N_21814,N_24031);
nor U27445 (N_27445,N_22602,N_22793);
nand U27446 (N_27446,N_20943,N_23101);
or U27447 (N_27447,N_21448,N_21697);
or U27448 (N_27448,N_22632,N_20326);
or U27449 (N_27449,N_22678,N_24071);
nor U27450 (N_27450,N_23533,N_23526);
or U27451 (N_27451,N_23969,N_23775);
or U27452 (N_27452,N_22496,N_20848);
or U27453 (N_27453,N_20587,N_24699);
or U27454 (N_27454,N_22544,N_24113);
or U27455 (N_27455,N_21552,N_20234);
nor U27456 (N_27456,N_24614,N_23392);
or U27457 (N_27457,N_20626,N_20216);
and U27458 (N_27458,N_21834,N_22483);
and U27459 (N_27459,N_20604,N_24102);
nand U27460 (N_27460,N_23643,N_20481);
and U27461 (N_27461,N_21853,N_23550);
and U27462 (N_27462,N_23753,N_23630);
nand U27463 (N_27463,N_23664,N_24025);
or U27464 (N_27464,N_22349,N_22309);
nor U27465 (N_27465,N_21857,N_21428);
and U27466 (N_27466,N_23231,N_22401);
nor U27467 (N_27467,N_23080,N_21190);
and U27468 (N_27468,N_22047,N_21873);
or U27469 (N_27469,N_22804,N_24304);
nand U27470 (N_27470,N_24963,N_21531);
nor U27471 (N_27471,N_23380,N_21546);
and U27472 (N_27472,N_21691,N_23315);
and U27473 (N_27473,N_21799,N_20099);
nand U27474 (N_27474,N_20336,N_23056);
nor U27475 (N_27475,N_22788,N_24762);
or U27476 (N_27476,N_24158,N_20546);
nor U27477 (N_27477,N_20709,N_23602);
xnor U27478 (N_27478,N_21062,N_21846);
or U27479 (N_27479,N_21307,N_22933);
nor U27480 (N_27480,N_23615,N_22171);
or U27481 (N_27481,N_22018,N_22787);
nor U27482 (N_27482,N_21115,N_20493);
nor U27483 (N_27483,N_23732,N_21719);
or U27484 (N_27484,N_20220,N_21110);
and U27485 (N_27485,N_22043,N_22876);
and U27486 (N_27486,N_21026,N_24015);
or U27487 (N_27487,N_22646,N_24144);
and U27488 (N_27488,N_22044,N_20612);
xnor U27489 (N_27489,N_22296,N_24196);
xor U27490 (N_27490,N_21599,N_20512);
nand U27491 (N_27491,N_24369,N_21801);
and U27492 (N_27492,N_21798,N_20895);
nor U27493 (N_27493,N_20780,N_21129);
or U27494 (N_27494,N_23939,N_24116);
nand U27495 (N_27495,N_22209,N_23880);
and U27496 (N_27496,N_24702,N_22179);
nand U27497 (N_27497,N_23563,N_22377);
xor U27498 (N_27498,N_20450,N_20172);
nor U27499 (N_27499,N_20739,N_24825);
or U27500 (N_27500,N_20150,N_20504);
nor U27501 (N_27501,N_23429,N_21475);
and U27502 (N_27502,N_22279,N_23281);
nor U27503 (N_27503,N_24912,N_21949);
or U27504 (N_27504,N_24484,N_22296);
nor U27505 (N_27505,N_20949,N_22953);
or U27506 (N_27506,N_21950,N_20955);
xor U27507 (N_27507,N_22539,N_24585);
xor U27508 (N_27508,N_23051,N_23021);
and U27509 (N_27509,N_20718,N_21503);
nand U27510 (N_27510,N_23251,N_22879);
nand U27511 (N_27511,N_22831,N_20458);
nor U27512 (N_27512,N_24566,N_24014);
xor U27513 (N_27513,N_20870,N_23377);
nor U27514 (N_27514,N_23097,N_20539);
or U27515 (N_27515,N_23478,N_21256);
xnor U27516 (N_27516,N_24006,N_21388);
nand U27517 (N_27517,N_21666,N_22325);
nor U27518 (N_27518,N_22757,N_20097);
or U27519 (N_27519,N_23435,N_21671);
nor U27520 (N_27520,N_20807,N_21821);
xor U27521 (N_27521,N_23221,N_23546);
and U27522 (N_27522,N_21674,N_24938);
nor U27523 (N_27523,N_24723,N_20507);
and U27524 (N_27524,N_22499,N_20754);
xnor U27525 (N_27525,N_24280,N_20471);
nor U27526 (N_27526,N_20505,N_20837);
xnor U27527 (N_27527,N_20438,N_23655);
xor U27528 (N_27528,N_24305,N_24444);
or U27529 (N_27529,N_24887,N_22424);
and U27530 (N_27530,N_20960,N_20969);
or U27531 (N_27531,N_23960,N_24025);
nand U27532 (N_27532,N_22052,N_21398);
or U27533 (N_27533,N_23553,N_24959);
and U27534 (N_27534,N_21402,N_23732);
nor U27535 (N_27535,N_21770,N_22621);
nand U27536 (N_27536,N_21585,N_22892);
nor U27537 (N_27537,N_22380,N_21289);
or U27538 (N_27538,N_24217,N_22768);
or U27539 (N_27539,N_22372,N_24025);
and U27540 (N_27540,N_22669,N_21873);
or U27541 (N_27541,N_24912,N_20668);
nor U27542 (N_27542,N_21258,N_22809);
and U27543 (N_27543,N_23607,N_24099);
nand U27544 (N_27544,N_23013,N_23521);
or U27545 (N_27545,N_23722,N_20659);
and U27546 (N_27546,N_22403,N_22814);
nand U27547 (N_27547,N_20356,N_20927);
xor U27548 (N_27548,N_20366,N_21674);
nor U27549 (N_27549,N_24948,N_23184);
xor U27550 (N_27550,N_24215,N_21092);
xor U27551 (N_27551,N_22601,N_20398);
nand U27552 (N_27552,N_20609,N_24738);
or U27553 (N_27553,N_20257,N_23536);
nor U27554 (N_27554,N_22458,N_21189);
or U27555 (N_27555,N_23574,N_20552);
or U27556 (N_27556,N_24502,N_24616);
or U27557 (N_27557,N_24483,N_21033);
xnor U27558 (N_27558,N_20280,N_21769);
nor U27559 (N_27559,N_20871,N_24954);
and U27560 (N_27560,N_23688,N_22457);
nand U27561 (N_27561,N_21207,N_21896);
xor U27562 (N_27562,N_22623,N_20398);
xnor U27563 (N_27563,N_23771,N_20767);
nor U27564 (N_27564,N_23600,N_20546);
xor U27565 (N_27565,N_24128,N_22476);
nor U27566 (N_27566,N_21529,N_24115);
and U27567 (N_27567,N_24513,N_21231);
xnor U27568 (N_27568,N_21940,N_22255);
and U27569 (N_27569,N_21540,N_23203);
nor U27570 (N_27570,N_20843,N_22253);
or U27571 (N_27571,N_21795,N_23856);
nand U27572 (N_27572,N_20031,N_22432);
nand U27573 (N_27573,N_21303,N_23220);
nand U27574 (N_27574,N_24949,N_23741);
or U27575 (N_27575,N_21500,N_23573);
nand U27576 (N_27576,N_21660,N_23074);
or U27577 (N_27577,N_24774,N_20294);
xor U27578 (N_27578,N_23148,N_23153);
and U27579 (N_27579,N_23129,N_22295);
or U27580 (N_27580,N_21744,N_22222);
or U27581 (N_27581,N_22497,N_21077);
nand U27582 (N_27582,N_20285,N_20942);
or U27583 (N_27583,N_23070,N_22397);
and U27584 (N_27584,N_20796,N_23309);
nand U27585 (N_27585,N_21858,N_23808);
or U27586 (N_27586,N_23969,N_23313);
nand U27587 (N_27587,N_23062,N_22454);
nor U27588 (N_27588,N_21960,N_24557);
or U27589 (N_27589,N_20829,N_24673);
nand U27590 (N_27590,N_22204,N_22599);
or U27591 (N_27591,N_22540,N_21843);
xor U27592 (N_27592,N_24914,N_21132);
nor U27593 (N_27593,N_23239,N_20531);
nand U27594 (N_27594,N_24800,N_24942);
nor U27595 (N_27595,N_20533,N_22977);
nor U27596 (N_27596,N_24111,N_23752);
xnor U27597 (N_27597,N_23141,N_24984);
and U27598 (N_27598,N_22723,N_22984);
xor U27599 (N_27599,N_20791,N_20907);
and U27600 (N_27600,N_20042,N_22014);
or U27601 (N_27601,N_24268,N_23820);
nand U27602 (N_27602,N_22353,N_22306);
or U27603 (N_27603,N_23720,N_20931);
and U27604 (N_27604,N_24952,N_24566);
or U27605 (N_27605,N_21377,N_24360);
xnor U27606 (N_27606,N_24201,N_21011);
or U27607 (N_27607,N_20484,N_24910);
xnor U27608 (N_27608,N_21171,N_22589);
nor U27609 (N_27609,N_21016,N_23165);
or U27610 (N_27610,N_22953,N_24455);
and U27611 (N_27611,N_20606,N_23914);
nor U27612 (N_27612,N_20867,N_22618);
and U27613 (N_27613,N_23655,N_22272);
xnor U27614 (N_27614,N_20777,N_21709);
xor U27615 (N_27615,N_22745,N_23271);
nand U27616 (N_27616,N_24862,N_24481);
and U27617 (N_27617,N_24022,N_20643);
and U27618 (N_27618,N_20397,N_20829);
xor U27619 (N_27619,N_21993,N_21856);
xor U27620 (N_27620,N_20260,N_24640);
xor U27621 (N_27621,N_20729,N_21211);
or U27622 (N_27622,N_24796,N_24846);
nand U27623 (N_27623,N_21808,N_24594);
nand U27624 (N_27624,N_20262,N_24053);
nand U27625 (N_27625,N_24623,N_23873);
or U27626 (N_27626,N_22192,N_24960);
xor U27627 (N_27627,N_22336,N_23693);
nand U27628 (N_27628,N_21151,N_20994);
and U27629 (N_27629,N_22917,N_22595);
nor U27630 (N_27630,N_20807,N_24942);
or U27631 (N_27631,N_22328,N_20536);
or U27632 (N_27632,N_20558,N_21249);
or U27633 (N_27633,N_24039,N_20223);
xor U27634 (N_27634,N_21192,N_24624);
or U27635 (N_27635,N_24341,N_22462);
xor U27636 (N_27636,N_20992,N_24057);
or U27637 (N_27637,N_21738,N_22211);
nor U27638 (N_27638,N_20927,N_21235);
nand U27639 (N_27639,N_23515,N_20416);
nand U27640 (N_27640,N_20041,N_24333);
xnor U27641 (N_27641,N_21144,N_21345);
and U27642 (N_27642,N_22450,N_23153);
nor U27643 (N_27643,N_21706,N_21807);
and U27644 (N_27644,N_22548,N_23095);
xor U27645 (N_27645,N_23502,N_23107);
and U27646 (N_27646,N_20101,N_23177);
xor U27647 (N_27647,N_24461,N_24742);
xor U27648 (N_27648,N_23756,N_22272);
or U27649 (N_27649,N_21329,N_21231);
and U27650 (N_27650,N_21835,N_22379);
nor U27651 (N_27651,N_20072,N_21226);
or U27652 (N_27652,N_24343,N_21355);
nor U27653 (N_27653,N_21095,N_24213);
xnor U27654 (N_27654,N_23164,N_22471);
nand U27655 (N_27655,N_22024,N_20812);
nand U27656 (N_27656,N_22607,N_23560);
nand U27657 (N_27657,N_20743,N_23862);
or U27658 (N_27658,N_20000,N_20357);
xnor U27659 (N_27659,N_24165,N_20946);
or U27660 (N_27660,N_20963,N_21946);
or U27661 (N_27661,N_20849,N_21058);
nor U27662 (N_27662,N_22880,N_24360);
xor U27663 (N_27663,N_22786,N_20878);
nor U27664 (N_27664,N_23935,N_21414);
and U27665 (N_27665,N_24929,N_22595);
or U27666 (N_27666,N_24795,N_20830);
and U27667 (N_27667,N_24450,N_20129);
and U27668 (N_27668,N_20076,N_24443);
or U27669 (N_27669,N_24051,N_22337);
nor U27670 (N_27670,N_20387,N_20386);
or U27671 (N_27671,N_20565,N_23404);
nand U27672 (N_27672,N_23982,N_24319);
xnor U27673 (N_27673,N_24286,N_24378);
and U27674 (N_27674,N_21902,N_21403);
and U27675 (N_27675,N_24118,N_22751);
nor U27676 (N_27676,N_22993,N_22213);
nor U27677 (N_27677,N_21179,N_22757);
and U27678 (N_27678,N_22343,N_24595);
xnor U27679 (N_27679,N_21426,N_23395);
nor U27680 (N_27680,N_23113,N_22108);
nand U27681 (N_27681,N_21738,N_20105);
nor U27682 (N_27682,N_20427,N_23715);
nand U27683 (N_27683,N_20603,N_20611);
nand U27684 (N_27684,N_22967,N_20642);
nand U27685 (N_27685,N_20945,N_20251);
and U27686 (N_27686,N_24591,N_23826);
nand U27687 (N_27687,N_23043,N_21315);
nor U27688 (N_27688,N_23506,N_24053);
nand U27689 (N_27689,N_20772,N_20672);
nor U27690 (N_27690,N_22293,N_23266);
nor U27691 (N_27691,N_24675,N_22741);
xor U27692 (N_27692,N_21745,N_22861);
nor U27693 (N_27693,N_23765,N_24433);
and U27694 (N_27694,N_23825,N_21498);
nor U27695 (N_27695,N_20407,N_20605);
nand U27696 (N_27696,N_22266,N_21065);
or U27697 (N_27697,N_21789,N_20146);
nand U27698 (N_27698,N_20697,N_23827);
xnor U27699 (N_27699,N_20621,N_20021);
nor U27700 (N_27700,N_23473,N_21320);
xnor U27701 (N_27701,N_21993,N_20881);
or U27702 (N_27702,N_24806,N_22709);
or U27703 (N_27703,N_24821,N_20163);
and U27704 (N_27704,N_22411,N_21308);
nand U27705 (N_27705,N_22469,N_22145);
and U27706 (N_27706,N_23471,N_24817);
and U27707 (N_27707,N_22540,N_20487);
or U27708 (N_27708,N_21592,N_23334);
and U27709 (N_27709,N_21047,N_21689);
xnor U27710 (N_27710,N_20859,N_21285);
nor U27711 (N_27711,N_24146,N_24055);
xnor U27712 (N_27712,N_21387,N_24567);
or U27713 (N_27713,N_21117,N_23770);
nor U27714 (N_27714,N_20915,N_21389);
nor U27715 (N_27715,N_20115,N_23573);
or U27716 (N_27716,N_23523,N_22924);
and U27717 (N_27717,N_21080,N_24313);
xor U27718 (N_27718,N_21611,N_21906);
nand U27719 (N_27719,N_20840,N_24063);
and U27720 (N_27720,N_24777,N_24486);
nand U27721 (N_27721,N_24916,N_24694);
or U27722 (N_27722,N_24434,N_22302);
or U27723 (N_27723,N_24600,N_23775);
xor U27724 (N_27724,N_20322,N_24961);
and U27725 (N_27725,N_23343,N_23278);
xor U27726 (N_27726,N_21429,N_22456);
and U27727 (N_27727,N_22068,N_21570);
xor U27728 (N_27728,N_23831,N_22911);
nand U27729 (N_27729,N_21146,N_21323);
xor U27730 (N_27730,N_21230,N_23001);
nand U27731 (N_27731,N_22957,N_21365);
or U27732 (N_27732,N_24455,N_23443);
or U27733 (N_27733,N_21194,N_20997);
and U27734 (N_27734,N_20175,N_23498);
or U27735 (N_27735,N_22374,N_23828);
and U27736 (N_27736,N_20322,N_24763);
nor U27737 (N_27737,N_22648,N_24810);
and U27738 (N_27738,N_20927,N_24165);
nand U27739 (N_27739,N_20773,N_23272);
or U27740 (N_27740,N_23196,N_24724);
and U27741 (N_27741,N_20386,N_20924);
xor U27742 (N_27742,N_22437,N_22403);
nor U27743 (N_27743,N_21640,N_22077);
nand U27744 (N_27744,N_24254,N_21223);
xnor U27745 (N_27745,N_20662,N_24897);
or U27746 (N_27746,N_24943,N_23297);
nand U27747 (N_27747,N_23417,N_20217);
nand U27748 (N_27748,N_24774,N_22854);
xor U27749 (N_27749,N_22734,N_23696);
or U27750 (N_27750,N_22121,N_21845);
or U27751 (N_27751,N_21199,N_24228);
nand U27752 (N_27752,N_22163,N_23278);
xnor U27753 (N_27753,N_20173,N_24903);
xnor U27754 (N_27754,N_21281,N_22277);
xor U27755 (N_27755,N_21377,N_24197);
nor U27756 (N_27756,N_24645,N_21163);
nand U27757 (N_27757,N_20865,N_24522);
nand U27758 (N_27758,N_20523,N_20446);
and U27759 (N_27759,N_21192,N_20880);
or U27760 (N_27760,N_21701,N_24080);
xor U27761 (N_27761,N_21148,N_24707);
or U27762 (N_27762,N_20138,N_22762);
xnor U27763 (N_27763,N_24850,N_20865);
and U27764 (N_27764,N_22411,N_20645);
nand U27765 (N_27765,N_21776,N_20846);
and U27766 (N_27766,N_20552,N_20917);
xnor U27767 (N_27767,N_24649,N_23216);
or U27768 (N_27768,N_22361,N_24563);
nor U27769 (N_27769,N_21297,N_23525);
nand U27770 (N_27770,N_21912,N_20634);
xor U27771 (N_27771,N_22807,N_24763);
xnor U27772 (N_27772,N_23664,N_23298);
nand U27773 (N_27773,N_21348,N_21080);
and U27774 (N_27774,N_23022,N_23406);
nor U27775 (N_27775,N_21230,N_24801);
and U27776 (N_27776,N_23348,N_22692);
and U27777 (N_27777,N_22367,N_22279);
or U27778 (N_27778,N_23604,N_21841);
nand U27779 (N_27779,N_22454,N_23442);
nand U27780 (N_27780,N_24751,N_21828);
or U27781 (N_27781,N_24366,N_23093);
and U27782 (N_27782,N_22344,N_20211);
nor U27783 (N_27783,N_22781,N_21851);
and U27784 (N_27784,N_23382,N_22102);
and U27785 (N_27785,N_20102,N_24209);
nand U27786 (N_27786,N_20178,N_23088);
xnor U27787 (N_27787,N_22082,N_23947);
nor U27788 (N_27788,N_24402,N_21052);
nand U27789 (N_27789,N_21977,N_20879);
nand U27790 (N_27790,N_20751,N_24977);
nor U27791 (N_27791,N_23673,N_21262);
xnor U27792 (N_27792,N_22201,N_23549);
xor U27793 (N_27793,N_23686,N_22171);
nand U27794 (N_27794,N_20004,N_22613);
nor U27795 (N_27795,N_24244,N_24895);
and U27796 (N_27796,N_21027,N_24614);
nand U27797 (N_27797,N_23176,N_23914);
nand U27798 (N_27798,N_21719,N_24988);
nand U27799 (N_27799,N_20707,N_24486);
and U27800 (N_27800,N_22539,N_20458);
nand U27801 (N_27801,N_21307,N_23681);
or U27802 (N_27802,N_20870,N_23075);
nand U27803 (N_27803,N_21106,N_24880);
or U27804 (N_27804,N_21589,N_22640);
nand U27805 (N_27805,N_21178,N_22762);
and U27806 (N_27806,N_22539,N_22214);
nor U27807 (N_27807,N_23824,N_21039);
nand U27808 (N_27808,N_23623,N_23401);
nor U27809 (N_27809,N_24122,N_22471);
nor U27810 (N_27810,N_24851,N_22278);
and U27811 (N_27811,N_24454,N_23835);
nand U27812 (N_27812,N_20926,N_24748);
or U27813 (N_27813,N_20183,N_21562);
and U27814 (N_27814,N_24906,N_22586);
nor U27815 (N_27815,N_23211,N_23457);
or U27816 (N_27816,N_20075,N_20907);
xnor U27817 (N_27817,N_21886,N_23560);
nor U27818 (N_27818,N_23972,N_24401);
xnor U27819 (N_27819,N_20719,N_24880);
xor U27820 (N_27820,N_23251,N_23939);
nand U27821 (N_27821,N_23369,N_24859);
or U27822 (N_27822,N_23484,N_23478);
nor U27823 (N_27823,N_21493,N_20275);
or U27824 (N_27824,N_24340,N_24233);
nor U27825 (N_27825,N_20093,N_23477);
xnor U27826 (N_27826,N_20845,N_22715);
nor U27827 (N_27827,N_21995,N_20854);
nand U27828 (N_27828,N_24274,N_20323);
and U27829 (N_27829,N_23660,N_21206);
xnor U27830 (N_27830,N_24106,N_22953);
xnor U27831 (N_27831,N_23811,N_22477);
xor U27832 (N_27832,N_22820,N_23790);
nand U27833 (N_27833,N_21106,N_23126);
nor U27834 (N_27834,N_23710,N_22371);
nor U27835 (N_27835,N_23759,N_20175);
nand U27836 (N_27836,N_21277,N_22000);
and U27837 (N_27837,N_21613,N_23669);
and U27838 (N_27838,N_20054,N_22009);
xor U27839 (N_27839,N_24036,N_20979);
nor U27840 (N_27840,N_20332,N_20243);
and U27841 (N_27841,N_23574,N_23541);
nor U27842 (N_27842,N_24405,N_23322);
and U27843 (N_27843,N_24273,N_23211);
nand U27844 (N_27844,N_23766,N_24787);
nor U27845 (N_27845,N_23795,N_22572);
and U27846 (N_27846,N_22838,N_21986);
nor U27847 (N_27847,N_21366,N_22875);
or U27848 (N_27848,N_24451,N_21680);
or U27849 (N_27849,N_24047,N_22142);
xnor U27850 (N_27850,N_20998,N_20970);
nand U27851 (N_27851,N_24395,N_23423);
nor U27852 (N_27852,N_22660,N_20275);
nor U27853 (N_27853,N_23425,N_23656);
nand U27854 (N_27854,N_23179,N_20686);
xnor U27855 (N_27855,N_22852,N_21282);
nand U27856 (N_27856,N_20247,N_23755);
and U27857 (N_27857,N_21475,N_20224);
xnor U27858 (N_27858,N_23808,N_21486);
nor U27859 (N_27859,N_23561,N_22922);
or U27860 (N_27860,N_23019,N_22879);
nand U27861 (N_27861,N_22757,N_22095);
or U27862 (N_27862,N_23348,N_20836);
nor U27863 (N_27863,N_24815,N_22109);
or U27864 (N_27864,N_24985,N_22306);
xnor U27865 (N_27865,N_20262,N_22529);
and U27866 (N_27866,N_24073,N_23862);
nand U27867 (N_27867,N_24456,N_21229);
and U27868 (N_27868,N_24002,N_22230);
xor U27869 (N_27869,N_20692,N_23240);
or U27870 (N_27870,N_20911,N_21998);
and U27871 (N_27871,N_22439,N_24160);
nor U27872 (N_27872,N_20411,N_23058);
nand U27873 (N_27873,N_22469,N_23382);
nor U27874 (N_27874,N_21438,N_22502);
and U27875 (N_27875,N_22429,N_21953);
and U27876 (N_27876,N_23983,N_20389);
nand U27877 (N_27877,N_21630,N_20309);
nor U27878 (N_27878,N_23402,N_21898);
nor U27879 (N_27879,N_24186,N_21404);
and U27880 (N_27880,N_23984,N_21318);
or U27881 (N_27881,N_21321,N_24243);
nand U27882 (N_27882,N_21203,N_23016);
xor U27883 (N_27883,N_22487,N_20003);
xor U27884 (N_27884,N_24313,N_23693);
nand U27885 (N_27885,N_24381,N_21120);
nor U27886 (N_27886,N_21961,N_20214);
xor U27887 (N_27887,N_21695,N_20726);
and U27888 (N_27888,N_20968,N_24015);
nor U27889 (N_27889,N_20801,N_20469);
xnor U27890 (N_27890,N_20791,N_22008);
xnor U27891 (N_27891,N_20919,N_23173);
nand U27892 (N_27892,N_22630,N_22325);
or U27893 (N_27893,N_24909,N_23589);
or U27894 (N_27894,N_21545,N_21506);
nor U27895 (N_27895,N_24844,N_20541);
nor U27896 (N_27896,N_20711,N_22444);
and U27897 (N_27897,N_21298,N_23593);
xor U27898 (N_27898,N_20515,N_24708);
nor U27899 (N_27899,N_22599,N_20122);
or U27900 (N_27900,N_23284,N_22579);
nand U27901 (N_27901,N_23491,N_21860);
xor U27902 (N_27902,N_21042,N_21152);
nand U27903 (N_27903,N_23408,N_24999);
xor U27904 (N_27904,N_22267,N_20192);
nand U27905 (N_27905,N_21173,N_20214);
or U27906 (N_27906,N_21267,N_23387);
nor U27907 (N_27907,N_20681,N_24016);
and U27908 (N_27908,N_20956,N_22254);
and U27909 (N_27909,N_22692,N_23521);
or U27910 (N_27910,N_20849,N_21298);
nand U27911 (N_27911,N_22518,N_24129);
nor U27912 (N_27912,N_23533,N_24646);
or U27913 (N_27913,N_20387,N_23093);
and U27914 (N_27914,N_21563,N_21840);
nor U27915 (N_27915,N_21366,N_20641);
xnor U27916 (N_27916,N_24405,N_23979);
xor U27917 (N_27917,N_24582,N_20914);
nor U27918 (N_27918,N_20943,N_20076);
and U27919 (N_27919,N_23430,N_22071);
xnor U27920 (N_27920,N_21550,N_24505);
and U27921 (N_27921,N_21643,N_23560);
or U27922 (N_27922,N_23491,N_22247);
nand U27923 (N_27923,N_24138,N_20107);
xor U27924 (N_27924,N_21989,N_24611);
nor U27925 (N_27925,N_20715,N_22687);
nor U27926 (N_27926,N_22252,N_23347);
and U27927 (N_27927,N_23347,N_20973);
or U27928 (N_27928,N_22931,N_21431);
nor U27929 (N_27929,N_22108,N_23590);
nand U27930 (N_27930,N_20023,N_24827);
or U27931 (N_27931,N_24796,N_21591);
xor U27932 (N_27932,N_24872,N_24054);
and U27933 (N_27933,N_24839,N_24381);
and U27934 (N_27934,N_21479,N_21918);
and U27935 (N_27935,N_22438,N_22204);
nand U27936 (N_27936,N_20021,N_20278);
and U27937 (N_27937,N_22506,N_24516);
and U27938 (N_27938,N_20898,N_20534);
or U27939 (N_27939,N_20072,N_22330);
xor U27940 (N_27940,N_20880,N_21712);
nor U27941 (N_27941,N_20440,N_24328);
or U27942 (N_27942,N_20479,N_20465);
xnor U27943 (N_27943,N_24853,N_24753);
or U27944 (N_27944,N_23326,N_22448);
or U27945 (N_27945,N_24982,N_23888);
or U27946 (N_27946,N_20486,N_23347);
nand U27947 (N_27947,N_23613,N_21475);
and U27948 (N_27948,N_20072,N_23669);
and U27949 (N_27949,N_21071,N_23374);
nor U27950 (N_27950,N_21012,N_23843);
nand U27951 (N_27951,N_22305,N_22066);
nand U27952 (N_27952,N_24502,N_22098);
xnor U27953 (N_27953,N_21269,N_24064);
nor U27954 (N_27954,N_21518,N_22068);
xor U27955 (N_27955,N_23088,N_22069);
nand U27956 (N_27956,N_24264,N_20819);
xor U27957 (N_27957,N_24347,N_21352);
nor U27958 (N_27958,N_24712,N_21220);
and U27959 (N_27959,N_23462,N_20077);
xor U27960 (N_27960,N_23614,N_20011);
nand U27961 (N_27961,N_24654,N_20275);
xor U27962 (N_27962,N_22400,N_21717);
nor U27963 (N_27963,N_23279,N_24825);
nand U27964 (N_27964,N_20630,N_20537);
xor U27965 (N_27965,N_23386,N_21162);
nand U27966 (N_27966,N_24782,N_20002);
xnor U27967 (N_27967,N_20446,N_21107);
or U27968 (N_27968,N_22269,N_23127);
xnor U27969 (N_27969,N_23562,N_23619);
or U27970 (N_27970,N_23056,N_24225);
or U27971 (N_27971,N_24897,N_24330);
xor U27972 (N_27972,N_23945,N_23957);
and U27973 (N_27973,N_23957,N_20572);
nor U27974 (N_27974,N_22028,N_20037);
and U27975 (N_27975,N_22497,N_22136);
nor U27976 (N_27976,N_24170,N_22254);
nor U27977 (N_27977,N_21925,N_21924);
or U27978 (N_27978,N_24237,N_23626);
and U27979 (N_27979,N_21921,N_24862);
nand U27980 (N_27980,N_22870,N_23701);
nand U27981 (N_27981,N_21622,N_20485);
and U27982 (N_27982,N_22466,N_20363);
nor U27983 (N_27983,N_21905,N_20205);
and U27984 (N_27984,N_24770,N_24323);
nor U27985 (N_27985,N_21736,N_20038);
or U27986 (N_27986,N_24087,N_20493);
and U27987 (N_27987,N_22683,N_24123);
nand U27988 (N_27988,N_20988,N_24404);
xor U27989 (N_27989,N_20490,N_22392);
nand U27990 (N_27990,N_21685,N_24900);
and U27991 (N_27991,N_22255,N_21600);
or U27992 (N_27992,N_22201,N_23888);
xnor U27993 (N_27993,N_23567,N_24069);
and U27994 (N_27994,N_24569,N_20378);
xor U27995 (N_27995,N_22982,N_21379);
and U27996 (N_27996,N_22603,N_20702);
or U27997 (N_27997,N_21561,N_24288);
or U27998 (N_27998,N_23855,N_21506);
nor U27999 (N_27999,N_22100,N_20046);
nor U28000 (N_28000,N_23232,N_23352);
xor U28001 (N_28001,N_21406,N_20549);
and U28002 (N_28002,N_23451,N_22359);
or U28003 (N_28003,N_22176,N_24973);
and U28004 (N_28004,N_23694,N_22315);
nand U28005 (N_28005,N_23661,N_22499);
nand U28006 (N_28006,N_24903,N_22001);
xnor U28007 (N_28007,N_20451,N_20536);
and U28008 (N_28008,N_23251,N_23738);
or U28009 (N_28009,N_21638,N_22288);
or U28010 (N_28010,N_24273,N_23965);
or U28011 (N_28011,N_21829,N_22049);
and U28012 (N_28012,N_23049,N_21818);
or U28013 (N_28013,N_24809,N_22813);
xor U28014 (N_28014,N_20492,N_20584);
and U28015 (N_28015,N_22031,N_22330);
xnor U28016 (N_28016,N_21923,N_22629);
nor U28017 (N_28017,N_23748,N_20708);
or U28018 (N_28018,N_22822,N_21813);
xor U28019 (N_28019,N_23814,N_23893);
nand U28020 (N_28020,N_24879,N_23292);
and U28021 (N_28021,N_22912,N_23050);
and U28022 (N_28022,N_21848,N_23487);
nand U28023 (N_28023,N_23339,N_24568);
or U28024 (N_28024,N_24035,N_22388);
nor U28025 (N_28025,N_24873,N_23606);
nor U28026 (N_28026,N_20760,N_24568);
or U28027 (N_28027,N_21217,N_21708);
xnor U28028 (N_28028,N_23633,N_21023);
and U28029 (N_28029,N_20363,N_20340);
xnor U28030 (N_28030,N_24572,N_20366);
xnor U28031 (N_28031,N_20163,N_24375);
and U28032 (N_28032,N_24287,N_24002);
xor U28033 (N_28033,N_22515,N_24662);
nand U28034 (N_28034,N_24909,N_22257);
xnor U28035 (N_28035,N_20707,N_22050);
or U28036 (N_28036,N_21451,N_21650);
nand U28037 (N_28037,N_21962,N_24667);
xnor U28038 (N_28038,N_21388,N_24036);
nor U28039 (N_28039,N_21075,N_22758);
xnor U28040 (N_28040,N_20280,N_20521);
xnor U28041 (N_28041,N_24121,N_24350);
nand U28042 (N_28042,N_21472,N_22442);
nor U28043 (N_28043,N_21214,N_21959);
or U28044 (N_28044,N_24076,N_22701);
nor U28045 (N_28045,N_24631,N_23484);
and U28046 (N_28046,N_20271,N_23483);
and U28047 (N_28047,N_23059,N_21305);
nor U28048 (N_28048,N_21728,N_24202);
and U28049 (N_28049,N_23515,N_22249);
or U28050 (N_28050,N_23564,N_21924);
xnor U28051 (N_28051,N_24390,N_24233);
and U28052 (N_28052,N_23851,N_24043);
xnor U28053 (N_28053,N_23801,N_24487);
or U28054 (N_28054,N_23625,N_22805);
nor U28055 (N_28055,N_21178,N_21106);
nand U28056 (N_28056,N_21118,N_23651);
nor U28057 (N_28057,N_22923,N_23906);
xnor U28058 (N_28058,N_21598,N_20899);
or U28059 (N_28059,N_22277,N_24144);
or U28060 (N_28060,N_20038,N_21183);
and U28061 (N_28061,N_22578,N_21527);
nand U28062 (N_28062,N_23544,N_22067);
and U28063 (N_28063,N_22633,N_20955);
or U28064 (N_28064,N_20605,N_20299);
and U28065 (N_28065,N_20237,N_20019);
nand U28066 (N_28066,N_21278,N_23093);
nand U28067 (N_28067,N_20755,N_22219);
and U28068 (N_28068,N_20651,N_20091);
and U28069 (N_28069,N_21081,N_20721);
and U28070 (N_28070,N_21563,N_21172);
or U28071 (N_28071,N_24271,N_20745);
nor U28072 (N_28072,N_21013,N_23261);
xnor U28073 (N_28073,N_23722,N_24133);
nand U28074 (N_28074,N_22875,N_24040);
and U28075 (N_28075,N_21080,N_21304);
xnor U28076 (N_28076,N_20460,N_22992);
nand U28077 (N_28077,N_22875,N_23058);
xnor U28078 (N_28078,N_20931,N_23951);
nand U28079 (N_28079,N_20196,N_23048);
nand U28080 (N_28080,N_21290,N_24206);
or U28081 (N_28081,N_23603,N_24197);
xnor U28082 (N_28082,N_24249,N_20393);
xnor U28083 (N_28083,N_22394,N_24462);
nor U28084 (N_28084,N_22524,N_24773);
and U28085 (N_28085,N_24200,N_22542);
nand U28086 (N_28086,N_23241,N_21985);
nor U28087 (N_28087,N_24056,N_23681);
nand U28088 (N_28088,N_22327,N_21140);
or U28089 (N_28089,N_24148,N_22206);
and U28090 (N_28090,N_23557,N_20816);
xor U28091 (N_28091,N_22592,N_20126);
and U28092 (N_28092,N_22855,N_20462);
nand U28093 (N_28093,N_24334,N_20147);
nand U28094 (N_28094,N_20219,N_23812);
nand U28095 (N_28095,N_21413,N_21936);
or U28096 (N_28096,N_23756,N_23490);
nand U28097 (N_28097,N_23876,N_23101);
and U28098 (N_28098,N_20091,N_20010);
nor U28099 (N_28099,N_24508,N_22523);
xor U28100 (N_28100,N_20635,N_24652);
xnor U28101 (N_28101,N_22605,N_23257);
nand U28102 (N_28102,N_20875,N_24571);
or U28103 (N_28103,N_24250,N_22410);
and U28104 (N_28104,N_21321,N_22591);
and U28105 (N_28105,N_24806,N_21539);
and U28106 (N_28106,N_20758,N_24524);
nand U28107 (N_28107,N_23582,N_23651);
and U28108 (N_28108,N_20409,N_21676);
or U28109 (N_28109,N_22212,N_21803);
xor U28110 (N_28110,N_20162,N_20472);
nand U28111 (N_28111,N_22811,N_22847);
xor U28112 (N_28112,N_21207,N_21969);
nor U28113 (N_28113,N_22409,N_20670);
and U28114 (N_28114,N_20288,N_23445);
nand U28115 (N_28115,N_23018,N_23769);
or U28116 (N_28116,N_22519,N_23100);
nor U28117 (N_28117,N_23473,N_20646);
nand U28118 (N_28118,N_23173,N_20934);
and U28119 (N_28119,N_20126,N_20963);
nor U28120 (N_28120,N_20328,N_20457);
xnor U28121 (N_28121,N_20026,N_24286);
or U28122 (N_28122,N_23591,N_21125);
and U28123 (N_28123,N_20292,N_20676);
nand U28124 (N_28124,N_22469,N_21743);
xnor U28125 (N_28125,N_23667,N_24323);
nand U28126 (N_28126,N_20730,N_22336);
and U28127 (N_28127,N_20133,N_22491);
nand U28128 (N_28128,N_22173,N_24547);
or U28129 (N_28129,N_22165,N_21152);
and U28130 (N_28130,N_23444,N_24633);
xnor U28131 (N_28131,N_23189,N_23464);
and U28132 (N_28132,N_23097,N_24198);
nand U28133 (N_28133,N_22045,N_21073);
nor U28134 (N_28134,N_20337,N_21419);
xnor U28135 (N_28135,N_22893,N_22544);
xor U28136 (N_28136,N_21389,N_23424);
nand U28137 (N_28137,N_23735,N_20828);
nor U28138 (N_28138,N_24008,N_20287);
and U28139 (N_28139,N_22787,N_20518);
and U28140 (N_28140,N_20308,N_22061);
or U28141 (N_28141,N_21355,N_20174);
and U28142 (N_28142,N_22190,N_21622);
or U28143 (N_28143,N_22602,N_22162);
nor U28144 (N_28144,N_21144,N_20079);
or U28145 (N_28145,N_23280,N_21125);
nand U28146 (N_28146,N_20150,N_20556);
nand U28147 (N_28147,N_24094,N_20700);
nand U28148 (N_28148,N_24847,N_22330);
and U28149 (N_28149,N_21799,N_21125);
nor U28150 (N_28150,N_24807,N_24851);
or U28151 (N_28151,N_23296,N_22803);
nor U28152 (N_28152,N_24389,N_24925);
nor U28153 (N_28153,N_23210,N_24847);
or U28154 (N_28154,N_24604,N_22230);
nand U28155 (N_28155,N_20183,N_20941);
or U28156 (N_28156,N_21761,N_23401);
and U28157 (N_28157,N_23896,N_20547);
nand U28158 (N_28158,N_20611,N_20490);
nor U28159 (N_28159,N_20378,N_23984);
or U28160 (N_28160,N_21160,N_24284);
and U28161 (N_28161,N_21734,N_22194);
and U28162 (N_28162,N_24110,N_20723);
and U28163 (N_28163,N_20533,N_24592);
and U28164 (N_28164,N_21175,N_20690);
nor U28165 (N_28165,N_20588,N_20966);
or U28166 (N_28166,N_22559,N_21774);
or U28167 (N_28167,N_22458,N_24808);
xor U28168 (N_28168,N_22930,N_23595);
or U28169 (N_28169,N_22449,N_22259);
and U28170 (N_28170,N_20468,N_20592);
or U28171 (N_28171,N_22043,N_24731);
and U28172 (N_28172,N_21421,N_20813);
nor U28173 (N_28173,N_21046,N_24569);
nor U28174 (N_28174,N_22143,N_23800);
nand U28175 (N_28175,N_22891,N_20352);
xnor U28176 (N_28176,N_21691,N_24466);
xor U28177 (N_28177,N_22433,N_24930);
or U28178 (N_28178,N_20885,N_22384);
nor U28179 (N_28179,N_22741,N_22387);
nor U28180 (N_28180,N_21994,N_20957);
or U28181 (N_28181,N_20441,N_23540);
and U28182 (N_28182,N_24532,N_24124);
nor U28183 (N_28183,N_22913,N_22591);
and U28184 (N_28184,N_24760,N_22351);
and U28185 (N_28185,N_22518,N_21026);
nor U28186 (N_28186,N_21327,N_20823);
nor U28187 (N_28187,N_20729,N_22870);
or U28188 (N_28188,N_21610,N_24801);
nor U28189 (N_28189,N_20162,N_24209);
and U28190 (N_28190,N_24227,N_21583);
nor U28191 (N_28191,N_21573,N_24655);
xor U28192 (N_28192,N_22377,N_23678);
and U28193 (N_28193,N_24831,N_22474);
nor U28194 (N_28194,N_23313,N_22935);
or U28195 (N_28195,N_21468,N_24428);
or U28196 (N_28196,N_20200,N_21849);
nor U28197 (N_28197,N_24736,N_23493);
or U28198 (N_28198,N_21124,N_22391);
or U28199 (N_28199,N_24793,N_20863);
nand U28200 (N_28200,N_21343,N_22104);
nand U28201 (N_28201,N_20506,N_23914);
or U28202 (N_28202,N_23375,N_20887);
nand U28203 (N_28203,N_24180,N_22905);
and U28204 (N_28204,N_21586,N_21562);
nand U28205 (N_28205,N_23390,N_20220);
xnor U28206 (N_28206,N_22416,N_23549);
nor U28207 (N_28207,N_21276,N_20833);
nor U28208 (N_28208,N_21609,N_20312);
nand U28209 (N_28209,N_20052,N_22389);
nor U28210 (N_28210,N_24688,N_21211);
xnor U28211 (N_28211,N_20876,N_23818);
or U28212 (N_28212,N_22888,N_21023);
xor U28213 (N_28213,N_24202,N_22483);
and U28214 (N_28214,N_22538,N_23263);
nor U28215 (N_28215,N_23173,N_21634);
nor U28216 (N_28216,N_24381,N_24241);
and U28217 (N_28217,N_22292,N_23581);
nand U28218 (N_28218,N_23849,N_21459);
or U28219 (N_28219,N_23153,N_20898);
and U28220 (N_28220,N_20114,N_24739);
nand U28221 (N_28221,N_20970,N_24400);
or U28222 (N_28222,N_20584,N_20170);
xnor U28223 (N_28223,N_24077,N_20935);
and U28224 (N_28224,N_23948,N_24144);
and U28225 (N_28225,N_23671,N_20919);
nand U28226 (N_28226,N_21872,N_23656);
nor U28227 (N_28227,N_22551,N_21827);
or U28228 (N_28228,N_21018,N_23627);
xnor U28229 (N_28229,N_22089,N_20193);
and U28230 (N_28230,N_20945,N_20289);
or U28231 (N_28231,N_22618,N_23112);
nand U28232 (N_28232,N_21211,N_23089);
nor U28233 (N_28233,N_20875,N_20964);
xor U28234 (N_28234,N_23246,N_22282);
or U28235 (N_28235,N_23023,N_21203);
or U28236 (N_28236,N_24477,N_23485);
xnor U28237 (N_28237,N_24015,N_24271);
or U28238 (N_28238,N_22325,N_24042);
nor U28239 (N_28239,N_21785,N_20677);
and U28240 (N_28240,N_21162,N_22027);
nor U28241 (N_28241,N_20370,N_20021);
nor U28242 (N_28242,N_20672,N_23907);
and U28243 (N_28243,N_20490,N_23097);
xor U28244 (N_28244,N_20500,N_23959);
and U28245 (N_28245,N_22425,N_21916);
xnor U28246 (N_28246,N_21844,N_22262);
nand U28247 (N_28247,N_23696,N_20299);
nor U28248 (N_28248,N_22511,N_20864);
nand U28249 (N_28249,N_20092,N_22535);
nand U28250 (N_28250,N_22103,N_23218);
or U28251 (N_28251,N_20560,N_24650);
or U28252 (N_28252,N_23727,N_22283);
nor U28253 (N_28253,N_20786,N_21719);
xor U28254 (N_28254,N_21974,N_23083);
or U28255 (N_28255,N_21508,N_23325);
nor U28256 (N_28256,N_20762,N_21521);
nand U28257 (N_28257,N_20747,N_21633);
nor U28258 (N_28258,N_22265,N_22288);
nor U28259 (N_28259,N_23877,N_23283);
xor U28260 (N_28260,N_23618,N_23423);
xor U28261 (N_28261,N_23730,N_22655);
xor U28262 (N_28262,N_24659,N_21577);
nand U28263 (N_28263,N_21666,N_20468);
xnor U28264 (N_28264,N_20590,N_22814);
nor U28265 (N_28265,N_20283,N_24683);
or U28266 (N_28266,N_22591,N_23656);
xnor U28267 (N_28267,N_22397,N_23071);
xor U28268 (N_28268,N_21415,N_20610);
and U28269 (N_28269,N_23282,N_23813);
nand U28270 (N_28270,N_22212,N_23645);
nor U28271 (N_28271,N_21440,N_20341);
nand U28272 (N_28272,N_22077,N_22931);
or U28273 (N_28273,N_20192,N_21074);
and U28274 (N_28274,N_21715,N_23478);
or U28275 (N_28275,N_21110,N_21915);
and U28276 (N_28276,N_24889,N_21328);
or U28277 (N_28277,N_20318,N_24878);
nand U28278 (N_28278,N_21541,N_24693);
nor U28279 (N_28279,N_22947,N_20569);
xor U28280 (N_28280,N_23318,N_23794);
xnor U28281 (N_28281,N_24139,N_20146);
and U28282 (N_28282,N_22162,N_23727);
or U28283 (N_28283,N_21749,N_20407);
xnor U28284 (N_28284,N_21749,N_24755);
and U28285 (N_28285,N_22136,N_23617);
or U28286 (N_28286,N_20153,N_24635);
xnor U28287 (N_28287,N_23403,N_23810);
nand U28288 (N_28288,N_21053,N_23959);
and U28289 (N_28289,N_21369,N_23989);
nor U28290 (N_28290,N_23944,N_20385);
or U28291 (N_28291,N_20197,N_23466);
xnor U28292 (N_28292,N_23054,N_20775);
xor U28293 (N_28293,N_20883,N_23786);
xor U28294 (N_28294,N_20160,N_23063);
or U28295 (N_28295,N_24910,N_22910);
xor U28296 (N_28296,N_20696,N_23693);
nand U28297 (N_28297,N_22226,N_23785);
or U28298 (N_28298,N_20880,N_22826);
nor U28299 (N_28299,N_22932,N_20427);
and U28300 (N_28300,N_22927,N_23394);
nor U28301 (N_28301,N_20816,N_24434);
or U28302 (N_28302,N_22605,N_20387);
xor U28303 (N_28303,N_22864,N_22479);
xor U28304 (N_28304,N_23471,N_22415);
and U28305 (N_28305,N_24529,N_21605);
nand U28306 (N_28306,N_20693,N_22406);
or U28307 (N_28307,N_22153,N_24191);
nand U28308 (N_28308,N_22607,N_23395);
nand U28309 (N_28309,N_23356,N_23134);
xnor U28310 (N_28310,N_21088,N_21477);
or U28311 (N_28311,N_24051,N_20254);
nand U28312 (N_28312,N_22593,N_23150);
or U28313 (N_28313,N_22116,N_21837);
xor U28314 (N_28314,N_23449,N_21010);
or U28315 (N_28315,N_22812,N_22297);
nand U28316 (N_28316,N_24369,N_21470);
nor U28317 (N_28317,N_20661,N_20071);
and U28318 (N_28318,N_20727,N_24764);
xor U28319 (N_28319,N_24698,N_23342);
or U28320 (N_28320,N_23159,N_23664);
nor U28321 (N_28321,N_20295,N_24179);
or U28322 (N_28322,N_20696,N_23389);
xor U28323 (N_28323,N_21964,N_20442);
and U28324 (N_28324,N_20016,N_20865);
nor U28325 (N_28325,N_23443,N_20349);
xor U28326 (N_28326,N_22457,N_21377);
nand U28327 (N_28327,N_23717,N_20495);
xor U28328 (N_28328,N_22931,N_22367);
nor U28329 (N_28329,N_20399,N_23384);
xor U28330 (N_28330,N_24938,N_22414);
xnor U28331 (N_28331,N_24000,N_21439);
nor U28332 (N_28332,N_22329,N_21664);
or U28333 (N_28333,N_22098,N_22333);
and U28334 (N_28334,N_22911,N_22125);
xor U28335 (N_28335,N_20476,N_23505);
and U28336 (N_28336,N_21630,N_20857);
and U28337 (N_28337,N_24080,N_23782);
xor U28338 (N_28338,N_22724,N_20443);
and U28339 (N_28339,N_24755,N_22837);
and U28340 (N_28340,N_23062,N_20137);
or U28341 (N_28341,N_21377,N_24253);
nor U28342 (N_28342,N_23440,N_21193);
xor U28343 (N_28343,N_20602,N_21808);
or U28344 (N_28344,N_24572,N_21210);
nand U28345 (N_28345,N_20572,N_22615);
nand U28346 (N_28346,N_21849,N_24482);
nor U28347 (N_28347,N_21779,N_20965);
nor U28348 (N_28348,N_20375,N_21376);
xor U28349 (N_28349,N_21690,N_21067);
or U28350 (N_28350,N_23263,N_22634);
and U28351 (N_28351,N_20015,N_23161);
nor U28352 (N_28352,N_24529,N_21201);
xnor U28353 (N_28353,N_21197,N_21409);
and U28354 (N_28354,N_24399,N_24230);
nand U28355 (N_28355,N_20465,N_24406);
nand U28356 (N_28356,N_20234,N_24791);
xnor U28357 (N_28357,N_21339,N_24569);
nor U28358 (N_28358,N_23687,N_24979);
and U28359 (N_28359,N_20139,N_24380);
nor U28360 (N_28360,N_20133,N_20515);
nand U28361 (N_28361,N_23916,N_21119);
nor U28362 (N_28362,N_22272,N_23452);
xnor U28363 (N_28363,N_22511,N_23675);
xnor U28364 (N_28364,N_23903,N_20447);
nor U28365 (N_28365,N_20099,N_24762);
or U28366 (N_28366,N_21946,N_23917);
or U28367 (N_28367,N_24409,N_22822);
nor U28368 (N_28368,N_22557,N_21014);
nand U28369 (N_28369,N_21414,N_24291);
or U28370 (N_28370,N_21584,N_21724);
nand U28371 (N_28371,N_24180,N_22455);
or U28372 (N_28372,N_20168,N_21143);
and U28373 (N_28373,N_22451,N_22345);
nand U28374 (N_28374,N_23602,N_21177);
nand U28375 (N_28375,N_22079,N_20491);
nor U28376 (N_28376,N_24107,N_23468);
or U28377 (N_28377,N_22969,N_21415);
or U28378 (N_28378,N_23015,N_20096);
or U28379 (N_28379,N_24117,N_23952);
and U28380 (N_28380,N_20482,N_22394);
xnor U28381 (N_28381,N_22689,N_24584);
nand U28382 (N_28382,N_24482,N_22343);
or U28383 (N_28383,N_24006,N_20174);
and U28384 (N_28384,N_23065,N_20848);
nor U28385 (N_28385,N_20981,N_20528);
and U28386 (N_28386,N_24656,N_21143);
nor U28387 (N_28387,N_21442,N_21579);
nand U28388 (N_28388,N_22919,N_23688);
nor U28389 (N_28389,N_23665,N_23943);
xor U28390 (N_28390,N_24807,N_21651);
or U28391 (N_28391,N_24577,N_23261);
xor U28392 (N_28392,N_24719,N_24387);
nand U28393 (N_28393,N_23792,N_21736);
xnor U28394 (N_28394,N_21404,N_24323);
or U28395 (N_28395,N_21860,N_23319);
xor U28396 (N_28396,N_23876,N_23643);
nor U28397 (N_28397,N_24193,N_20082);
xor U28398 (N_28398,N_24588,N_24334);
nor U28399 (N_28399,N_21010,N_24887);
xor U28400 (N_28400,N_21221,N_24464);
or U28401 (N_28401,N_24342,N_21647);
or U28402 (N_28402,N_24673,N_23682);
and U28403 (N_28403,N_24794,N_24962);
and U28404 (N_28404,N_24058,N_23194);
or U28405 (N_28405,N_24598,N_21757);
and U28406 (N_28406,N_24314,N_20195);
and U28407 (N_28407,N_20702,N_21006);
nand U28408 (N_28408,N_22127,N_24115);
and U28409 (N_28409,N_21197,N_24698);
or U28410 (N_28410,N_21680,N_22546);
nor U28411 (N_28411,N_21128,N_23137);
nor U28412 (N_28412,N_22484,N_21766);
nor U28413 (N_28413,N_24691,N_20678);
nor U28414 (N_28414,N_20147,N_24145);
nand U28415 (N_28415,N_21025,N_22098);
nor U28416 (N_28416,N_22646,N_23050);
xor U28417 (N_28417,N_21754,N_22345);
nand U28418 (N_28418,N_22019,N_20147);
nand U28419 (N_28419,N_22726,N_24313);
or U28420 (N_28420,N_20201,N_24799);
or U28421 (N_28421,N_22262,N_21767);
or U28422 (N_28422,N_20005,N_24242);
or U28423 (N_28423,N_21216,N_21311);
nand U28424 (N_28424,N_23920,N_20234);
nor U28425 (N_28425,N_22305,N_21610);
and U28426 (N_28426,N_20065,N_20752);
xnor U28427 (N_28427,N_21344,N_22299);
or U28428 (N_28428,N_20592,N_23878);
or U28429 (N_28429,N_21895,N_21276);
xor U28430 (N_28430,N_20408,N_20365);
nand U28431 (N_28431,N_24844,N_23214);
xnor U28432 (N_28432,N_23215,N_20668);
or U28433 (N_28433,N_24304,N_24307);
nand U28434 (N_28434,N_24346,N_20108);
or U28435 (N_28435,N_23594,N_22577);
nand U28436 (N_28436,N_21861,N_24190);
or U28437 (N_28437,N_23474,N_21086);
and U28438 (N_28438,N_22575,N_22861);
or U28439 (N_28439,N_24333,N_23770);
xor U28440 (N_28440,N_20148,N_22090);
nand U28441 (N_28441,N_24721,N_24143);
xor U28442 (N_28442,N_20363,N_24068);
or U28443 (N_28443,N_20804,N_24200);
nor U28444 (N_28444,N_21397,N_23655);
nand U28445 (N_28445,N_20971,N_20244);
and U28446 (N_28446,N_20798,N_23432);
nor U28447 (N_28447,N_20360,N_21119);
and U28448 (N_28448,N_22702,N_22559);
xor U28449 (N_28449,N_21021,N_24132);
nor U28450 (N_28450,N_23054,N_21001);
nor U28451 (N_28451,N_22933,N_21037);
nand U28452 (N_28452,N_22672,N_21075);
and U28453 (N_28453,N_23617,N_21871);
xor U28454 (N_28454,N_20466,N_20589);
xor U28455 (N_28455,N_21164,N_20479);
or U28456 (N_28456,N_24545,N_22051);
nor U28457 (N_28457,N_24788,N_21471);
nor U28458 (N_28458,N_22414,N_24049);
xnor U28459 (N_28459,N_20240,N_24144);
nor U28460 (N_28460,N_22714,N_20699);
nand U28461 (N_28461,N_23184,N_21260);
or U28462 (N_28462,N_22293,N_20609);
xnor U28463 (N_28463,N_24923,N_24817);
nor U28464 (N_28464,N_20466,N_24141);
nor U28465 (N_28465,N_21957,N_20997);
nand U28466 (N_28466,N_21328,N_22137);
and U28467 (N_28467,N_22779,N_20258);
or U28468 (N_28468,N_24878,N_21835);
nor U28469 (N_28469,N_23403,N_20345);
nand U28470 (N_28470,N_21587,N_22996);
or U28471 (N_28471,N_24139,N_21887);
xor U28472 (N_28472,N_22573,N_20047);
xnor U28473 (N_28473,N_20183,N_22430);
xnor U28474 (N_28474,N_20123,N_24078);
or U28475 (N_28475,N_20185,N_22852);
nor U28476 (N_28476,N_23630,N_21821);
or U28477 (N_28477,N_23706,N_24395);
or U28478 (N_28478,N_23526,N_24377);
nand U28479 (N_28479,N_21585,N_22169);
nor U28480 (N_28480,N_23131,N_20801);
nand U28481 (N_28481,N_21085,N_24234);
and U28482 (N_28482,N_21425,N_21334);
or U28483 (N_28483,N_22811,N_20350);
and U28484 (N_28484,N_20917,N_21603);
and U28485 (N_28485,N_22589,N_23002);
or U28486 (N_28486,N_20536,N_23815);
and U28487 (N_28487,N_24601,N_22401);
nand U28488 (N_28488,N_20233,N_21153);
xnor U28489 (N_28489,N_23004,N_21679);
and U28490 (N_28490,N_23070,N_23824);
nor U28491 (N_28491,N_24760,N_20241);
nor U28492 (N_28492,N_20595,N_22911);
xnor U28493 (N_28493,N_22881,N_22282);
or U28494 (N_28494,N_22357,N_22959);
nor U28495 (N_28495,N_21164,N_24530);
and U28496 (N_28496,N_22175,N_23646);
xnor U28497 (N_28497,N_22730,N_21001);
and U28498 (N_28498,N_22366,N_23612);
and U28499 (N_28499,N_21173,N_23222);
nand U28500 (N_28500,N_23058,N_24841);
nand U28501 (N_28501,N_20453,N_24367);
nor U28502 (N_28502,N_24640,N_23836);
nand U28503 (N_28503,N_21694,N_24338);
nor U28504 (N_28504,N_23352,N_22382);
nor U28505 (N_28505,N_22007,N_23536);
xnor U28506 (N_28506,N_20040,N_23758);
and U28507 (N_28507,N_22286,N_21749);
and U28508 (N_28508,N_22718,N_20439);
or U28509 (N_28509,N_21032,N_20900);
and U28510 (N_28510,N_24609,N_23302);
xnor U28511 (N_28511,N_24037,N_24465);
nand U28512 (N_28512,N_22654,N_23320);
xnor U28513 (N_28513,N_24271,N_20615);
or U28514 (N_28514,N_23127,N_24509);
and U28515 (N_28515,N_22821,N_21831);
nor U28516 (N_28516,N_23891,N_21491);
nor U28517 (N_28517,N_22534,N_20991);
and U28518 (N_28518,N_20826,N_21220);
xor U28519 (N_28519,N_21348,N_23754);
xnor U28520 (N_28520,N_24682,N_24105);
and U28521 (N_28521,N_24241,N_22564);
or U28522 (N_28522,N_20351,N_21049);
nand U28523 (N_28523,N_22246,N_20216);
nor U28524 (N_28524,N_23392,N_23709);
xnor U28525 (N_28525,N_23773,N_20991);
and U28526 (N_28526,N_21189,N_22017);
or U28527 (N_28527,N_23583,N_21351);
nor U28528 (N_28528,N_21926,N_20810);
or U28529 (N_28529,N_22379,N_22862);
and U28530 (N_28530,N_22203,N_21573);
nand U28531 (N_28531,N_20680,N_24468);
and U28532 (N_28532,N_23137,N_23463);
and U28533 (N_28533,N_23504,N_23784);
and U28534 (N_28534,N_20205,N_24943);
nor U28535 (N_28535,N_24697,N_20053);
nor U28536 (N_28536,N_24609,N_20322);
nor U28537 (N_28537,N_24757,N_21095);
and U28538 (N_28538,N_21899,N_23026);
and U28539 (N_28539,N_23809,N_22113);
nor U28540 (N_28540,N_20865,N_22345);
nor U28541 (N_28541,N_24726,N_22950);
nor U28542 (N_28542,N_21157,N_24107);
xnor U28543 (N_28543,N_23453,N_22679);
and U28544 (N_28544,N_20746,N_22288);
xnor U28545 (N_28545,N_24072,N_24908);
xor U28546 (N_28546,N_23581,N_20476);
nand U28547 (N_28547,N_24679,N_20185);
and U28548 (N_28548,N_24177,N_20675);
xor U28549 (N_28549,N_24287,N_23436);
nor U28550 (N_28550,N_22834,N_21341);
nor U28551 (N_28551,N_24415,N_23932);
nand U28552 (N_28552,N_20796,N_22734);
and U28553 (N_28553,N_20111,N_23894);
and U28554 (N_28554,N_24457,N_24215);
xnor U28555 (N_28555,N_20721,N_24944);
or U28556 (N_28556,N_23735,N_24297);
nor U28557 (N_28557,N_24193,N_23780);
and U28558 (N_28558,N_24616,N_24642);
nand U28559 (N_28559,N_24796,N_23566);
or U28560 (N_28560,N_24833,N_24750);
nand U28561 (N_28561,N_22511,N_24040);
xor U28562 (N_28562,N_23751,N_23105);
and U28563 (N_28563,N_21914,N_23387);
and U28564 (N_28564,N_24551,N_24671);
or U28565 (N_28565,N_24664,N_22191);
nor U28566 (N_28566,N_22168,N_22205);
xnor U28567 (N_28567,N_24193,N_23546);
nand U28568 (N_28568,N_21200,N_21445);
nand U28569 (N_28569,N_22170,N_21797);
and U28570 (N_28570,N_23033,N_21061);
nand U28571 (N_28571,N_20266,N_23023);
nand U28572 (N_28572,N_24095,N_24512);
and U28573 (N_28573,N_23999,N_23394);
and U28574 (N_28574,N_24654,N_20804);
or U28575 (N_28575,N_23754,N_23790);
xnor U28576 (N_28576,N_21659,N_23625);
nand U28577 (N_28577,N_23025,N_24571);
nor U28578 (N_28578,N_22072,N_21653);
nand U28579 (N_28579,N_20731,N_21074);
xor U28580 (N_28580,N_24800,N_20547);
and U28581 (N_28581,N_21252,N_24427);
and U28582 (N_28582,N_24442,N_23895);
nor U28583 (N_28583,N_20474,N_23815);
nor U28584 (N_28584,N_24853,N_22832);
xnor U28585 (N_28585,N_22311,N_21629);
nand U28586 (N_28586,N_20954,N_23087);
or U28587 (N_28587,N_24306,N_23581);
and U28588 (N_28588,N_20874,N_22769);
nor U28589 (N_28589,N_23773,N_22016);
nand U28590 (N_28590,N_21690,N_24639);
or U28591 (N_28591,N_24763,N_24219);
nor U28592 (N_28592,N_22482,N_24129);
nor U28593 (N_28593,N_23616,N_24581);
and U28594 (N_28594,N_22076,N_21832);
xor U28595 (N_28595,N_20881,N_21107);
nor U28596 (N_28596,N_23052,N_24063);
nor U28597 (N_28597,N_22444,N_22326);
nand U28598 (N_28598,N_21670,N_23671);
or U28599 (N_28599,N_24628,N_23890);
or U28600 (N_28600,N_22785,N_21336);
or U28601 (N_28601,N_22329,N_21892);
or U28602 (N_28602,N_22939,N_20025);
nor U28603 (N_28603,N_24536,N_20621);
nand U28604 (N_28604,N_24692,N_22392);
or U28605 (N_28605,N_24490,N_24624);
or U28606 (N_28606,N_21827,N_22197);
and U28607 (N_28607,N_22961,N_23064);
or U28608 (N_28608,N_23568,N_21906);
xor U28609 (N_28609,N_23458,N_23425);
and U28610 (N_28610,N_21060,N_20445);
xor U28611 (N_28611,N_22918,N_23907);
and U28612 (N_28612,N_22155,N_20357);
and U28613 (N_28613,N_23692,N_23629);
or U28614 (N_28614,N_24667,N_23013);
xor U28615 (N_28615,N_21757,N_20935);
or U28616 (N_28616,N_21319,N_21688);
or U28617 (N_28617,N_21293,N_21498);
nor U28618 (N_28618,N_23541,N_24748);
or U28619 (N_28619,N_20631,N_23160);
xnor U28620 (N_28620,N_22197,N_23008);
nand U28621 (N_28621,N_24917,N_23457);
and U28622 (N_28622,N_23247,N_23693);
nor U28623 (N_28623,N_21702,N_24063);
and U28624 (N_28624,N_24101,N_24748);
or U28625 (N_28625,N_20090,N_22591);
and U28626 (N_28626,N_22642,N_20233);
nor U28627 (N_28627,N_24038,N_20396);
nand U28628 (N_28628,N_20727,N_23371);
xor U28629 (N_28629,N_20576,N_22665);
nand U28630 (N_28630,N_23424,N_23146);
or U28631 (N_28631,N_22359,N_24075);
nor U28632 (N_28632,N_23291,N_20805);
nor U28633 (N_28633,N_21761,N_23450);
xnor U28634 (N_28634,N_21379,N_23774);
nor U28635 (N_28635,N_21246,N_23666);
or U28636 (N_28636,N_23621,N_20040);
nand U28637 (N_28637,N_24616,N_21807);
nand U28638 (N_28638,N_23306,N_21430);
nand U28639 (N_28639,N_23759,N_20419);
or U28640 (N_28640,N_23430,N_20114);
and U28641 (N_28641,N_20475,N_21581);
or U28642 (N_28642,N_20742,N_21831);
nand U28643 (N_28643,N_22107,N_20095);
nand U28644 (N_28644,N_22607,N_24783);
nand U28645 (N_28645,N_21443,N_21257);
nand U28646 (N_28646,N_23186,N_21026);
xor U28647 (N_28647,N_20281,N_24777);
and U28648 (N_28648,N_24303,N_22484);
and U28649 (N_28649,N_20635,N_20676);
and U28650 (N_28650,N_24354,N_23518);
and U28651 (N_28651,N_21737,N_23019);
nor U28652 (N_28652,N_20088,N_23349);
and U28653 (N_28653,N_24894,N_23715);
xor U28654 (N_28654,N_24782,N_20261);
nand U28655 (N_28655,N_20595,N_20200);
nand U28656 (N_28656,N_24936,N_23839);
and U28657 (N_28657,N_20283,N_23389);
nor U28658 (N_28658,N_22267,N_21623);
xnor U28659 (N_28659,N_22200,N_22203);
xnor U28660 (N_28660,N_23029,N_21089);
xor U28661 (N_28661,N_21519,N_22042);
or U28662 (N_28662,N_21367,N_23219);
nand U28663 (N_28663,N_22439,N_24848);
xor U28664 (N_28664,N_22746,N_24037);
or U28665 (N_28665,N_22215,N_22494);
nor U28666 (N_28666,N_21180,N_21545);
or U28667 (N_28667,N_24537,N_24435);
xnor U28668 (N_28668,N_23282,N_23080);
or U28669 (N_28669,N_21219,N_23618);
nand U28670 (N_28670,N_24514,N_22807);
nor U28671 (N_28671,N_22270,N_20904);
or U28672 (N_28672,N_21246,N_23980);
or U28673 (N_28673,N_24969,N_24454);
or U28674 (N_28674,N_23143,N_20481);
nor U28675 (N_28675,N_22594,N_20589);
nor U28676 (N_28676,N_24139,N_20644);
xor U28677 (N_28677,N_20203,N_21522);
nand U28678 (N_28678,N_21383,N_22514);
and U28679 (N_28679,N_23061,N_21608);
nand U28680 (N_28680,N_20048,N_23337);
nor U28681 (N_28681,N_22882,N_24814);
nor U28682 (N_28682,N_23033,N_24888);
or U28683 (N_28683,N_22489,N_24687);
or U28684 (N_28684,N_23448,N_20384);
and U28685 (N_28685,N_21666,N_21534);
and U28686 (N_28686,N_20904,N_24760);
nand U28687 (N_28687,N_24100,N_21252);
nor U28688 (N_28688,N_23609,N_21425);
xor U28689 (N_28689,N_20456,N_23895);
and U28690 (N_28690,N_22775,N_22199);
or U28691 (N_28691,N_21207,N_20564);
nor U28692 (N_28692,N_23496,N_21898);
nor U28693 (N_28693,N_23853,N_20412);
nand U28694 (N_28694,N_23513,N_22972);
and U28695 (N_28695,N_20551,N_24154);
nor U28696 (N_28696,N_22835,N_23164);
xnor U28697 (N_28697,N_24856,N_24005);
and U28698 (N_28698,N_20306,N_24766);
nand U28699 (N_28699,N_23602,N_24915);
or U28700 (N_28700,N_20201,N_24772);
and U28701 (N_28701,N_24866,N_24655);
xnor U28702 (N_28702,N_22308,N_21542);
nand U28703 (N_28703,N_23848,N_23466);
nand U28704 (N_28704,N_22859,N_21675);
xor U28705 (N_28705,N_24929,N_24310);
nor U28706 (N_28706,N_21539,N_21404);
xnor U28707 (N_28707,N_21539,N_20452);
and U28708 (N_28708,N_22002,N_22029);
or U28709 (N_28709,N_20912,N_24705);
xnor U28710 (N_28710,N_21722,N_24295);
and U28711 (N_28711,N_21098,N_21435);
xor U28712 (N_28712,N_21308,N_22273);
nand U28713 (N_28713,N_24838,N_20047);
and U28714 (N_28714,N_24317,N_24459);
and U28715 (N_28715,N_21797,N_24514);
or U28716 (N_28716,N_20688,N_23796);
nor U28717 (N_28717,N_24374,N_23001);
or U28718 (N_28718,N_23097,N_24004);
and U28719 (N_28719,N_24945,N_23485);
nand U28720 (N_28720,N_22737,N_21417);
nor U28721 (N_28721,N_24340,N_21895);
or U28722 (N_28722,N_24830,N_21289);
nand U28723 (N_28723,N_21622,N_21199);
or U28724 (N_28724,N_24702,N_22921);
nor U28725 (N_28725,N_22801,N_20500);
and U28726 (N_28726,N_24103,N_24251);
and U28727 (N_28727,N_20702,N_23314);
and U28728 (N_28728,N_22779,N_20169);
nor U28729 (N_28729,N_23869,N_22780);
nand U28730 (N_28730,N_23263,N_24813);
nor U28731 (N_28731,N_22954,N_21834);
nand U28732 (N_28732,N_23276,N_21842);
xnor U28733 (N_28733,N_22189,N_20152);
and U28734 (N_28734,N_20230,N_21420);
or U28735 (N_28735,N_24338,N_23863);
nand U28736 (N_28736,N_20493,N_24813);
xnor U28737 (N_28737,N_23999,N_24949);
nor U28738 (N_28738,N_24279,N_20117);
xor U28739 (N_28739,N_22230,N_22896);
or U28740 (N_28740,N_20010,N_22393);
or U28741 (N_28741,N_24543,N_22312);
nor U28742 (N_28742,N_23492,N_22954);
or U28743 (N_28743,N_24683,N_21079);
nor U28744 (N_28744,N_24516,N_20146);
nand U28745 (N_28745,N_21968,N_21540);
nand U28746 (N_28746,N_20452,N_24722);
xnor U28747 (N_28747,N_22242,N_22396);
and U28748 (N_28748,N_20479,N_21879);
or U28749 (N_28749,N_22340,N_24938);
nand U28750 (N_28750,N_20983,N_22389);
nand U28751 (N_28751,N_20161,N_23792);
or U28752 (N_28752,N_20998,N_21330);
and U28753 (N_28753,N_22688,N_21182);
nor U28754 (N_28754,N_20168,N_22543);
nand U28755 (N_28755,N_23347,N_21902);
or U28756 (N_28756,N_23312,N_24492);
and U28757 (N_28757,N_20056,N_22935);
or U28758 (N_28758,N_20175,N_20229);
nand U28759 (N_28759,N_23454,N_20182);
and U28760 (N_28760,N_21928,N_20502);
and U28761 (N_28761,N_21605,N_21673);
nor U28762 (N_28762,N_23163,N_20645);
xnor U28763 (N_28763,N_24895,N_20602);
xnor U28764 (N_28764,N_23433,N_23668);
nor U28765 (N_28765,N_23848,N_22271);
xnor U28766 (N_28766,N_24278,N_22274);
xnor U28767 (N_28767,N_20936,N_22302);
xnor U28768 (N_28768,N_23099,N_23839);
and U28769 (N_28769,N_24209,N_23201);
nor U28770 (N_28770,N_20090,N_22034);
nand U28771 (N_28771,N_23587,N_21414);
nand U28772 (N_28772,N_22151,N_23694);
nand U28773 (N_28773,N_24914,N_23157);
nor U28774 (N_28774,N_20340,N_21813);
xnor U28775 (N_28775,N_22067,N_21986);
xor U28776 (N_28776,N_22636,N_22775);
or U28777 (N_28777,N_23140,N_21123);
xor U28778 (N_28778,N_20201,N_21985);
nand U28779 (N_28779,N_20199,N_20374);
and U28780 (N_28780,N_20756,N_20667);
xnor U28781 (N_28781,N_24706,N_21387);
or U28782 (N_28782,N_20957,N_23700);
nor U28783 (N_28783,N_23974,N_20504);
or U28784 (N_28784,N_24988,N_23268);
and U28785 (N_28785,N_20968,N_24220);
nor U28786 (N_28786,N_21186,N_20238);
or U28787 (N_28787,N_24662,N_24474);
xor U28788 (N_28788,N_22342,N_21008);
nand U28789 (N_28789,N_22287,N_20174);
xnor U28790 (N_28790,N_21949,N_24516);
and U28791 (N_28791,N_21087,N_23572);
or U28792 (N_28792,N_22695,N_23059);
and U28793 (N_28793,N_24597,N_20765);
xnor U28794 (N_28794,N_24823,N_23234);
and U28795 (N_28795,N_20499,N_21456);
and U28796 (N_28796,N_24685,N_20952);
xnor U28797 (N_28797,N_20647,N_24744);
or U28798 (N_28798,N_23186,N_20168);
nand U28799 (N_28799,N_24408,N_24411);
nand U28800 (N_28800,N_24318,N_21203);
and U28801 (N_28801,N_24924,N_22013);
or U28802 (N_28802,N_20626,N_23696);
or U28803 (N_28803,N_24036,N_23528);
and U28804 (N_28804,N_22757,N_23714);
and U28805 (N_28805,N_20516,N_22663);
nor U28806 (N_28806,N_24469,N_20807);
nand U28807 (N_28807,N_20826,N_23074);
nand U28808 (N_28808,N_24529,N_24082);
nor U28809 (N_28809,N_24099,N_22944);
nand U28810 (N_28810,N_22836,N_21134);
and U28811 (N_28811,N_23524,N_22988);
xor U28812 (N_28812,N_23387,N_20052);
nor U28813 (N_28813,N_22013,N_22878);
and U28814 (N_28814,N_21943,N_21647);
nand U28815 (N_28815,N_22458,N_24397);
and U28816 (N_28816,N_21374,N_20935);
xnor U28817 (N_28817,N_23031,N_22256);
or U28818 (N_28818,N_23944,N_23840);
xor U28819 (N_28819,N_24589,N_24946);
xnor U28820 (N_28820,N_21003,N_23437);
and U28821 (N_28821,N_24376,N_22221);
nand U28822 (N_28822,N_24854,N_20562);
nand U28823 (N_28823,N_22904,N_20283);
nor U28824 (N_28824,N_21800,N_22022);
nand U28825 (N_28825,N_21373,N_24132);
nand U28826 (N_28826,N_21756,N_24368);
nor U28827 (N_28827,N_20228,N_24682);
and U28828 (N_28828,N_24683,N_24604);
nand U28829 (N_28829,N_23102,N_22452);
nand U28830 (N_28830,N_23775,N_21035);
and U28831 (N_28831,N_20071,N_22409);
xnor U28832 (N_28832,N_21779,N_21933);
nand U28833 (N_28833,N_23464,N_21731);
or U28834 (N_28834,N_21169,N_23817);
or U28835 (N_28835,N_23352,N_24225);
or U28836 (N_28836,N_24098,N_21324);
nand U28837 (N_28837,N_20674,N_23859);
nor U28838 (N_28838,N_20030,N_22218);
xnor U28839 (N_28839,N_23996,N_22658);
nand U28840 (N_28840,N_23160,N_24409);
nand U28841 (N_28841,N_21934,N_23912);
nor U28842 (N_28842,N_23363,N_22906);
nor U28843 (N_28843,N_23391,N_23031);
nor U28844 (N_28844,N_24315,N_24626);
nand U28845 (N_28845,N_22116,N_20561);
or U28846 (N_28846,N_23707,N_20349);
xnor U28847 (N_28847,N_23939,N_24986);
or U28848 (N_28848,N_22683,N_24420);
or U28849 (N_28849,N_22791,N_22256);
xor U28850 (N_28850,N_21318,N_24895);
nand U28851 (N_28851,N_20475,N_21187);
nor U28852 (N_28852,N_22090,N_20881);
or U28853 (N_28853,N_22921,N_22046);
nor U28854 (N_28854,N_20430,N_23509);
nand U28855 (N_28855,N_20272,N_20128);
nor U28856 (N_28856,N_20013,N_20646);
and U28857 (N_28857,N_20498,N_24442);
and U28858 (N_28858,N_24272,N_23940);
nor U28859 (N_28859,N_22575,N_20612);
or U28860 (N_28860,N_20702,N_22940);
nand U28861 (N_28861,N_22398,N_22302);
nor U28862 (N_28862,N_20675,N_23540);
or U28863 (N_28863,N_23269,N_22840);
nand U28864 (N_28864,N_20647,N_23926);
xor U28865 (N_28865,N_20881,N_24977);
and U28866 (N_28866,N_20444,N_22011);
nor U28867 (N_28867,N_23218,N_23088);
xor U28868 (N_28868,N_20966,N_22039);
and U28869 (N_28869,N_23089,N_23929);
nand U28870 (N_28870,N_23933,N_21846);
nand U28871 (N_28871,N_22386,N_21827);
and U28872 (N_28872,N_23560,N_22422);
or U28873 (N_28873,N_21447,N_21514);
nor U28874 (N_28874,N_21842,N_23899);
xnor U28875 (N_28875,N_23919,N_24827);
nand U28876 (N_28876,N_20919,N_21769);
nand U28877 (N_28877,N_20503,N_21532);
xnor U28878 (N_28878,N_20778,N_20051);
nor U28879 (N_28879,N_22231,N_20123);
nor U28880 (N_28880,N_22567,N_23623);
nand U28881 (N_28881,N_21570,N_22059);
or U28882 (N_28882,N_21508,N_22174);
or U28883 (N_28883,N_23875,N_24509);
and U28884 (N_28884,N_23506,N_24253);
xor U28885 (N_28885,N_20442,N_23673);
and U28886 (N_28886,N_20054,N_22615);
or U28887 (N_28887,N_24751,N_24157);
or U28888 (N_28888,N_23947,N_24585);
nor U28889 (N_28889,N_23189,N_24286);
nand U28890 (N_28890,N_21936,N_24924);
and U28891 (N_28891,N_23343,N_23026);
nor U28892 (N_28892,N_20386,N_21502);
and U28893 (N_28893,N_20811,N_22915);
and U28894 (N_28894,N_24410,N_23873);
or U28895 (N_28895,N_20856,N_21863);
nor U28896 (N_28896,N_24538,N_21986);
or U28897 (N_28897,N_20839,N_23607);
and U28898 (N_28898,N_23389,N_21519);
nor U28899 (N_28899,N_24450,N_21217);
and U28900 (N_28900,N_20565,N_22939);
nand U28901 (N_28901,N_24079,N_24028);
nor U28902 (N_28902,N_22676,N_23420);
nand U28903 (N_28903,N_22403,N_20984);
or U28904 (N_28904,N_20113,N_21070);
xnor U28905 (N_28905,N_20778,N_20867);
nor U28906 (N_28906,N_24001,N_24756);
nor U28907 (N_28907,N_22403,N_21819);
or U28908 (N_28908,N_21690,N_24689);
nor U28909 (N_28909,N_20164,N_24496);
nand U28910 (N_28910,N_24125,N_23180);
xnor U28911 (N_28911,N_20991,N_22157);
or U28912 (N_28912,N_24019,N_24487);
xor U28913 (N_28913,N_20125,N_23205);
nand U28914 (N_28914,N_24069,N_23355);
xnor U28915 (N_28915,N_21162,N_24974);
or U28916 (N_28916,N_24552,N_23068);
and U28917 (N_28917,N_21439,N_22938);
xor U28918 (N_28918,N_21930,N_20289);
xnor U28919 (N_28919,N_20824,N_22694);
nand U28920 (N_28920,N_22850,N_23947);
nand U28921 (N_28921,N_21866,N_23494);
nor U28922 (N_28922,N_23482,N_23622);
or U28923 (N_28923,N_20574,N_23264);
and U28924 (N_28924,N_22352,N_20826);
and U28925 (N_28925,N_23927,N_22732);
nand U28926 (N_28926,N_24080,N_22380);
nand U28927 (N_28927,N_22173,N_21950);
or U28928 (N_28928,N_23372,N_23552);
or U28929 (N_28929,N_20088,N_24869);
nor U28930 (N_28930,N_21590,N_20700);
nor U28931 (N_28931,N_20490,N_24151);
nor U28932 (N_28932,N_22653,N_23783);
xor U28933 (N_28933,N_23105,N_20905);
nand U28934 (N_28934,N_23735,N_20387);
nand U28935 (N_28935,N_20318,N_20753);
nand U28936 (N_28936,N_21450,N_24523);
xnor U28937 (N_28937,N_21129,N_20660);
xnor U28938 (N_28938,N_20644,N_24990);
nand U28939 (N_28939,N_20359,N_20667);
and U28940 (N_28940,N_23333,N_21427);
xor U28941 (N_28941,N_20345,N_23852);
nor U28942 (N_28942,N_23994,N_24737);
nand U28943 (N_28943,N_22494,N_21873);
nand U28944 (N_28944,N_22822,N_22812);
nand U28945 (N_28945,N_22940,N_22810);
nor U28946 (N_28946,N_23913,N_20012);
and U28947 (N_28947,N_24227,N_24519);
xor U28948 (N_28948,N_23650,N_20110);
nor U28949 (N_28949,N_22925,N_24603);
nor U28950 (N_28950,N_24571,N_22019);
and U28951 (N_28951,N_20753,N_20596);
nor U28952 (N_28952,N_24425,N_21926);
or U28953 (N_28953,N_21333,N_23379);
nor U28954 (N_28954,N_22401,N_20976);
and U28955 (N_28955,N_22674,N_21335);
and U28956 (N_28956,N_22637,N_20753);
nor U28957 (N_28957,N_23368,N_22493);
xor U28958 (N_28958,N_23070,N_24418);
or U28959 (N_28959,N_24954,N_23840);
xor U28960 (N_28960,N_21950,N_20933);
nand U28961 (N_28961,N_23711,N_23402);
nor U28962 (N_28962,N_22777,N_20729);
xor U28963 (N_28963,N_21546,N_22599);
or U28964 (N_28964,N_21296,N_22509);
or U28965 (N_28965,N_22536,N_23332);
or U28966 (N_28966,N_22795,N_20769);
nand U28967 (N_28967,N_23677,N_23771);
and U28968 (N_28968,N_22756,N_22071);
or U28969 (N_28969,N_23454,N_21033);
and U28970 (N_28970,N_24329,N_20394);
xnor U28971 (N_28971,N_24471,N_21216);
xor U28972 (N_28972,N_24538,N_24384);
nand U28973 (N_28973,N_22213,N_20716);
or U28974 (N_28974,N_23689,N_21522);
nand U28975 (N_28975,N_23043,N_21526);
nor U28976 (N_28976,N_20109,N_23101);
xnor U28977 (N_28977,N_21981,N_22323);
and U28978 (N_28978,N_23187,N_20899);
and U28979 (N_28979,N_24317,N_23560);
nand U28980 (N_28980,N_23954,N_23207);
xnor U28981 (N_28981,N_20453,N_21242);
and U28982 (N_28982,N_24865,N_20631);
nand U28983 (N_28983,N_20810,N_21795);
xor U28984 (N_28984,N_21676,N_22644);
xor U28985 (N_28985,N_23315,N_20702);
xor U28986 (N_28986,N_22514,N_24943);
nor U28987 (N_28987,N_23965,N_23747);
and U28988 (N_28988,N_23648,N_24437);
nor U28989 (N_28989,N_24686,N_20404);
nand U28990 (N_28990,N_22265,N_22999);
xor U28991 (N_28991,N_21478,N_22348);
or U28992 (N_28992,N_23786,N_23886);
and U28993 (N_28993,N_20825,N_22641);
nand U28994 (N_28994,N_23348,N_23912);
or U28995 (N_28995,N_22153,N_20181);
xor U28996 (N_28996,N_22012,N_21643);
xnor U28997 (N_28997,N_23006,N_20019);
nand U28998 (N_28998,N_24434,N_22326);
nor U28999 (N_28999,N_24022,N_21419);
xnor U29000 (N_29000,N_24432,N_23496);
and U29001 (N_29001,N_21343,N_23059);
nand U29002 (N_29002,N_20812,N_20663);
nor U29003 (N_29003,N_22617,N_21988);
and U29004 (N_29004,N_23400,N_22445);
nand U29005 (N_29005,N_24816,N_24041);
and U29006 (N_29006,N_22844,N_23590);
nand U29007 (N_29007,N_22227,N_21045);
nor U29008 (N_29008,N_22116,N_20495);
nand U29009 (N_29009,N_23578,N_23782);
xor U29010 (N_29010,N_20573,N_20184);
xnor U29011 (N_29011,N_22669,N_23786);
and U29012 (N_29012,N_20688,N_20617);
nand U29013 (N_29013,N_23532,N_21027);
nand U29014 (N_29014,N_21333,N_21971);
xor U29015 (N_29015,N_24839,N_20427);
and U29016 (N_29016,N_22335,N_20706);
nor U29017 (N_29017,N_22123,N_20215);
and U29018 (N_29018,N_24596,N_21270);
nand U29019 (N_29019,N_24512,N_23598);
nand U29020 (N_29020,N_20133,N_21531);
nand U29021 (N_29021,N_24171,N_20079);
xnor U29022 (N_29022,N_22633,N_24872);
xor U29023 (N_29023,N_21845,N_21686);
nand U29024 (N_29024,N_23058,N_23003);
and U29025 (N_29025,N_24118,N_24149);
or U29026 (N_29026,N_20225,N_22610);
xor U29027 (N_29027,N_20032,N_24195);
nand U29028 (N_29028,N_21990,N_22245);
or U29029 (N_29029,N_22182,N_20151);
xnor U29030 (N_29030,N_20346,N_23894);
xor U29031 (N_29031,N_24815,N_24647);
or U29032 (N_29032,N_23497,N_22561);
nor U29033 (N_29033,N_20064,N_21011);
or U29034 (N_29034,N_23185,N_21255);
nor U29035 (N_29035,N_23350,N_20566);
nor U29036 (N_29036,N_24173,N_20111);
xor U29037 (N_29037,N_22329,N_21582);
xor U29038 (N_29038,N_21513,N_20951);
and U29039 (N_29039,N_20604,N_24813);
xor U29040 (N_29040,N_24947,N_24689);
and U29041 (N_29041,N_21666,N_22413);
and U29042 (N_29042,N_23729,N_21921);
xor U29043 (N_29043,N_21119,N_20835);
nand U29044 (N_29044,N_22286,N_23149);
xnor U29045 (N_29045,N_21743,N_22217);
or U29046 (N_29046,N_20633,N_24816);
nor U29047 (N_29047,N_20933,N_24149);
or U29048 (N_29048,N_22212,N_22233);
nor U29049 (N_29049,N_24987,N_20011);
nand U29050 (N_29050,N_21487,N_23893);
nand U29051 (N_29051,N_20223,N_21630);
and U29052 (N_29052,N_22280,N_20387);
xor U29053 (N_29053,N_20113,N_21108);
nand U29054 (N_29054,N_21112,N_22673);
nor U29055 (N_29055,N_22596,N_23655);
and U29056 (N_29056,N_21041,N_21600);
xnor U29057 (N_29057,N_23827,N_21777);
nor U29058 (N_29058,N_22528,N_22053);
or U29059 (N_29059,N_21822,N_23715);
xor U29060 (N_29060,N_23633,N_24339);
nor U29061 (N_29061,N_22766,N_20356);
and U29062 (N_29062,N_22476,N_24535);
and U29063 (N_29063,N_24017,N_20584);
or U29064 (N_29064,N_22674,N_21066);
or U29065 (N_29065,N_20540,N_24723);
nand U29066 (N_29066,N_23290,N_23337);
xnor U29067 (N_29067,N_24788,N_24309);
nor U29068 (N_29068,N_23572,N_24349);
and U29069 (N_29069,N_24724,N_22052);
nand U29070 (N_29070,N_21303,N_23448);
nor U29071 (N_29071,N_24772,N_22745);
or U29072 (N_29072,N_21893,N_22496);
or U29073 (N_29073,N_23074,N_21457);
nor U29074 (N_29074,N_21663,N_20947);
nand U29075 (N_29075,N_22765,N_21042);
and U29076 (N_29076,N_24293,N_20536);
and U29077 (N_29077,N_20386,N_22372);
xor U29078 (N_29078,N_24411,N_24386);
and U29079 (N_29079,N_22749,N_24806);
and U29080 (N_29080,N_22548,N_20653);
and U29081 (N_29081,N_23216,N_24185);
and U29082 (N_29082,N_23849,N_23561);
and U29083 (N_29083,N_20174,N_24778);
xnor U29084 (N_29084,N_24069,N_22565);
or U29085 (N_29085,N_24225,N_23969);
nand U29086 (N_29086,N_20473,N_21591);
or U29087 (N_29087,N_22530,N_20372);
nand U29088 (N_29088,N_22399,N_20962);
nor U29089 (N_29089,N_20161,N_22398);
or U29090 (N_29090,N_22205,N_20188);
or U29091 (N_29091,N_20901,N_21491);
nand U29092 (N_29092,N_24093,N_21156);
nor U29093 (N_29093,N_23536,N_20298);
and U29094 (N_29094,N_23276,N_20657);
or U29095 (N_29095,N_23017,N_24077);
nand U29096 (N_29096,N_24564,N_24632);
nor U29097 (N_29097,N_24941,N_21950);
xor U29098 (N_29098,N_22997,N_21001);
nand U29099 (N_29099,N_22900,N_23082);
nor U29100 (N_29100,N_24747,N_24288);
or U29101 (N_29101,N_23897,N_22684);
or U29102 (N_29102,N_22886,N_21749);
xor U29103 (N_29103,N_21402,N_23232);
nand U29104 (N_29104,N_22320,N_21649);
xor U29105 (N_29105,N_21623,N_23577);
nor U29106 (N_29106,N_21929,N_24986);
xnor U29107 (N_29107,N_24118,N_21475);
nor U29108 (N_29108,N_22825,N_24468);
and U29109 (N_29109,N_21532,N_20400);
nand U29110 (N_29110,N_22632,N_21415);
xor U29111 (N_29111,N_20785,N_22910);
nand U29112 (N_29112,N_20709,N_24125);
or U29113 (N_29113,N_24654,N_21268);
or U29114 (N_29114,N_22274,N_20206);
nor U29115 (N_29115,N_24252,N_22537);
xnor U29116 (N_29116,N_24579,N_24382);
xor U29117 (N_29117,N_20498,N_23517);
xnor U29118 (N_29118,N_24219,N_23071);
nor U29119 (N_29119,N_21132,N_24980);
nand U29120 (N_29120,N_23272,N_21062);
nand U29121 (N_29121,N_21857,N_20270);
nand U29122 (N_29122,N_23239,N_21154);
nand U29123 (N_29123,N_23294,N_21686);
xor U29124 (N_29124,N_21674,N_23796);
nor U29125 (N_29125,N_21101,N_21022);
and U29126 (N_29126,N_22169,N_21394);
nor U29127 (N_29127,N_21193,N_24958);
nand U29128 (N_29128,N_20119,N_20502);
nor U29129 (N_29129,N_21699,N_20946);
nand U29130 (N_29130,N_22348,N_24174);
or U29131 (N_29131,N_22029,N_23424);
xor U29132 (N_29132,N_20170,N_23987);
and U29133 (N_29133,N_21733,N_22376);
and U29134 (N_29134,N_24430,N_20235);
or U29135 (N_29135,N_24936,N_20596);
nor U29136 (N_29136,N_24897,N_21920);
and U29137 (N_29137,N_22671,N_21508);
xnor U29138 (N_29138,N_20392,N_23474);
xnor U29139 (N_29139,N_24712,N_21938);
or U29140 (N_29140,N_24401,N_24760);
nand U29141 (N_29141,N_24292,N_20571);
nand U29142 (N_29142,N_24276,N_21401);
and U29143 (N_29143,N_22596,N_21170);
nor U29144 (N_29144,N_22437,N_22778);
xnor U29145 (N_29145,N_21320,N_21557);
nor U29146 (N_29146,N_22890,N_22687);
nor U29147 (N_29147,N_21716,N_21305);
nand U29148 (N_29148,N_22789,N_20791);
and U29149 (N_29149,N_23488,N_23201);
nor U29150 (N_29150,N_21912,N_20854);
nor U29151 (N_29151,N_22756,N_20185);
nand U29152 (N_29152,N_20383,N_23638);
nor U29153 (N_29153,N_21112,N_21798);
and U29154 (N_29154,N_21681,N_24402);
xnor U29155 (N_29155,N_20035,N_24696);
xor U29156 (N_29156,N_21966,N_20855);
and U29157 (N_29157,N_22558,N_23612);
and U29158 (N_29158,N_21535,N_23880);
nor U29159 (N_29159,N_23195,N_22715);
and U29160 (N_29160,N_24726,N_23763);
xor U29161 (N_29161,N_21873,N_23681);
or U29162 (N_29162,N_23002,N_21154);
or U29163 (N_29163,N_21306,N_22765);
xnor U29164 (N_29164,N_24763,N_23062);
nor U29165 (N_29165,N_23695,N_22499);
or U29166 (N_29166,N_23312,N_24107);
xor U29167 (N_29167,N_22727,N_24294);
or U29168 (N_29168,N_21140,N_24439);
nor U29169 (N_29169,N_20287,N_22030);
nor U29170 (N_29170,N_22746,N_21356);
or U29171 (N_29171,N_24639,N_20882);
nor U29172 (N_29172,N_20417,N_21071);
nor U29173 (N_29173,N_23626,N_20614);
xor U29174 (N_29174,N_23993,N_23602);
nor U29175 (N_29175,N_22630,N_21120);
nand U29176 (N_29176,N_22138,N_21489);
nand U29177 (N_29177,N_21235,N_23383);
xor U29178 (N_29178,N_21425,N_20959);
nor U29179 (N_29179,N_21083,N_24772);
xor U29180 (N_29180,N_24345,N_22038);
nor U29181 (N_29181,N_22136,N_24323);
or U29182 (N_29182,N_24102,N_22331);
nor U29183 (N_29183,N_21938,N_24272);
xnor U29184 (N_29184,N_22935,N_20365);
and U29185 (N_29185,N_21295,N_24455);
xnor U29186 (N_29186,N_23570,N_21502);
or U29187 (N_29187,N_22749,N_24873);
xnor U29188 (N_29188,N_22179,N_22901);
or U29189 (N_29189,N_22243,N_24522);
nor U29190 (N_29190,N_20127,N_24283);
or U29191 (N_29191,N_21316,N_20262);
nand U29192 (N_29192,N_21772,N_24957);
xnor U29193 (N_29193,N_24896,N_21622);
or U29194 (N_29194,N_24729,N_21120);
xnor U29195 (N_29195,N_23257,N_20423);
and U29196 (N_29196,N_21413,N_22155);
nor U29197 (N_29197,N_23057,N_21566);
nor U29198 (N_29198,N_22845,N_23994);
nor U29199 (N_29199,N_23525,N_23871);
nor U29200 (N_29200,N_21060,N_24115);
nor U29201 (N_29201,N_22456,N_24452);
or U29202 (N_29202,N_22868,N_22016);
and U29203 (N_29203,N_21985,N_21203);
nor U29204 (N_29204,N_20641,N_22281);
and U29205 (N_29205,N_20015,N_20345);
and U29206 (N_29206,N_20878,N_23544);
xor U29207 (N_29207,N_21525,N_20348);
xnor U29208 (N_29208,N_20160,N_21495);
nand U29209 (N_29209,N_24875,N_23770);
xnor U29210 (N_29210,N_24873,N_22252);
or U29211 (N_29211,N_21888,N_23472);
xor U29212 (N_29212,N_24814,N_22079);
or U29213 (N_29213,N_23574,N_22432);
xor U29214 (N_29214,N_22826,N_21003);
or U29215 (N_29215,N_20680,N_21112);
and U29216 (N_29216,N_23925,N_22597);
xnor U29217 (N_29217,N_23383,N_22194);
nand U29218 (N_29218,N_20563,N_22399);
xnor U29219 (N_29219,N_24051,N_21878);
nor U29220 (N_29220,N_22366,N_23800);
or U29221 (N_29221,N_23809,N_20008);
nor U29222 (N_29222,N_22872,N_21164);
or U29223 (N_29223,N_22307,N_23892);
nor U29224 (N_29224,N_21903,N_24821);
and U29225 (N_29225,N_21364,N_22971);
or U29226 (N_29226,N_22143,N_22429);
nor U29227 (N_29227,N_21599,N_21449);
or U29228 (N_29228,N_20372,N_20627);
and U29229 (N_29229,N_24217,N_23626);
xor U29230 (N_29230,N_20713,N_24220);
or U29231 (N_29231,N_23837,N_23854);
or U29232 (N_29232,N_24876,N_24725);
and U29233 (N_29233,N_23067,N_21887);
nand U29234 (N_29234,N_21637,N_24611);
and U29235 (N_29235,N_24779,N_22567);
nor U29236 (N_29236,N_20073,N_21176);
and U29237 (N_29237,N_24058,N_21004);
nor U29238 (N_29238,N_21923,N_24635);
and U29239 (N_29239,N_23029,N_21226);
or U29240 (N_29240,N_22791,N_20619);
nor U29241 (N_29241,N_20481,N_22946);
and U29242 (N_29242,N_21758,N_24948);
xnor U29243 (N_29243,N_22868,N_23361);
nor U29244 (N_29244,N_21093,N_22277);
xor U29245 (N_29245,N_23816,N_21251);
or U29246 (N_29246,N_21524,N_23230);
nor U29247 (N_29247,N_22357,N_21414);
or U29248 (N_29248,N_23524,N_23656);
nand U29249 (N_29249,N_22760,N_22237);
nor U29250 (N_29250,N_24552,N_20916);
nor U29251 (N_29251,N_23542,N_22179);
nand U29252 (N_29252,N_23308,N_20959);
nand U29253 (N_29253,N_23002,N_23396);
or U29254 (N_29254,N_24297,N_20044);
or U29255 (N_29255,N_23086,N_22679);
nor U29256 (N_29256,N_24125,N_21339);
nand U29257 (N_29257,N_20231,N_22692);
nor U29258 (N_29258,N_23575,N_24053);
nor U29259 (N_29259,N_21741,N_23854);
nor U29260 (N_29260,N_20339,N_23654);
or U29261 (N_29261,N_24047,N_20145);
or U29262 (N_29262,N_24847,N_22024);
xor U29263 (N_29263,N_24040,N_24174);
nor U29264 (N_29264,N_23547,N_23894);
or U29265 (N_29265,N_21752,N_24112);
nor U29266 (N_29266,N_20600,N_21265);
and U29267 (N_29267,N_23973,N_20067);
nor U29268 (N_29268,N_21731,N_23069);
or U29269 (N_29269,N_24003,N_21636);
or U29270 (N_29270,N_22664,N_24881);
or U29271 (N_29271,N_22389,N_21358);
nand U29272 (N_29272,N_24688,N_20344);
nand U29273 (N_29273,N_22355,N_20122);
nand U29274 (N_29274,N_24801,N_23460);
and U29275 (N_29275,N_20042,N_21060);
or U29276 (N_29276,N_22499,N_22374);
xor U29277 (N_29277,N_24195,N_24110);
nor U29278 (N_29278,N_21365,N_22900);
and U29279 (N_29279,N_24631,N_24279);
nor U29280 (N_29280,N_22258,N_20511);
xor U29281 (N_29281,N_24820,N_21158);
nand U29282 (N_29282,N_20877,N_23377);
and U29283 (N_29283,N_22504,N_22677);
or U29284 (N_29284,N_20573,N_22345);
or U29285 (N_29285,N_23609,N_22535);
xnor U29286 (N_29286,N_23791,N_22006);
nand U29287 (N_29287,N_20876,N_24405);
and U29288 (N_29288,N_22132,N_23905);
nor U29289 (N_29289,N_24586,N_21109);
xor U29290 (N_29290,N_24033,N_21358);
and U29291 (N_29291,N_20569,N_23358);
or U29292 (N_29292,N_24894,N_21207);
or U29293 (N_29293,N_20566,N_21629);
and U29294 (N_29294,N_20903,N_22995);
or U29295 (N_29295,N_20165,N_21759);
xor U29296 (N_29296,N_21827,N_23171);
or U29297 (N_29297,N_24883,N_23112);
nor U29298 (N_29298,N_22997,N_21254);
and U29299 (N_29299,N_22319,N_24705);
and U29300 (N_29300,N_20919,N_23969);
and U29301 (N_29301,N_24300,N_22891);
nor U29302 (N_29302,N_21668,N_21339);
xor U29303 (N_29303,N_21026,N_23597);
xnor U29304 (N_29304,N_20244,N_22889);
nand U29305 (N_29305,N_22649,N_23858);
nor U29306 (N_29306,N_22823,N_21516);
nand U29307 (N_29307,N_20885,N_21257);
nand U29308 (N_29308,N_21783,N_20191);
nor U29309 (N_29309,N_21425,N_21149);
xnor U29310 (N_29310,N_23239,N_23123);
xnor U29311 (N_29311,N_21925,N_23894);
xor U29312 (N_29312,N_22179,N_21265);
and U29313 (N_29313,N_24384,N_23809);
or U29314 (N_29314,N_20890,N_24388);
and U29315 (N_29315,N_20960,N_20459);
xnor U29316 (N_29316,N_20418,N_20481);
nand U29317 (N_29317,N_21323,N_20707);
nand U29318 (N_29318,N_23928,N_24169);
nor U29319 (N_29319,N_24314,N_22030);
or U29320 (N_29320,N_23105,N_20514);
and U29321 (N_29321,N_23044,N_23288);
xor U29322 (N_29322,N_22904,N_21081);
xor U29323 (N_29323,N_22368,N_24045);
and U29324 (N_29324,N_22425,N_22731);
and U29325 (N_29325,N_21293,N_20640);
and U29326 (N_29326,N_24824,N_21318);
and U29327 (N_29327,N_24981,N_21850);
nor U29328 (N_29328,N_22208,N_24672);
nor U29329 (N_29329,N_21532,N_23895);
nand U29330 (N_29330,N_23997,N_23708);
or U29331 (N_29331,N_22797,N_23605);
or U29332 (N_29332,N_24157,N_22270);
or U29333 (N_29333,N_23762,N_21186);
or U29334 (N_29334,N_20684,N_22697);
nand U29335 (N_29335,N_23002,N_24556);
nor U29336 (N_29336,N_21866,N_23648);
xnor U29337 (N_29337,N_22935,N_23725);
nor U29338 (N_29338,N_21592,N_22342);
xnor U29339 (N_29339,N_20603,N_24520);
or U29340 (N_29340,N_20737,N_23566);
xnor U29341 (N_29341,N_23976,N_23816);
and U29342 (N_29342,N_24924,N_22851);
and U29343 (N_29343,N_23454,N_24095);
or U29344 (N_29344,N_20221,N_23835);
xor U29345 (N_29345,N_20592,N_22775);
xnor U29346 (N_29346,N_22607,N_23318);
nand U29347 (N_29347,N_24829,N_20035);
xor U29348 (N_29348,N_24975,N_23257);
and U29349 (N_29349,N_24440,N_21167);
or U29350 (N_29350,N_24482,N_23756);
xor U29351 (N_29351,N_20875,N_23159);
nand U29352 (N_29352,N_22431,N_20625);
xnor U29353 (N_29353,N_21611,N_20938);
nand U29354 (N_29354,N_20791,N_22382);
xnor U29355 (N_29355,N_24293,N_20053);
nand U29356 (N_29356,N_20070,N_21273);
xor U29357 (N_29357,N_22953,N_21646);
nand U29358 (N_29358,N_21388,N_23509);
nor U29359 (N_29359,N_24816,N_24667);
and U29360 (N_29360,N_24818,N_24062);
nand U29361 (N_29361,N_21581,N_21034);
and U29362 (N_29362,N_23448,N_24133);
xnor U29363 (N_29363,N_23835,N_20627);
nor U29364 (N_29364,N_20412,N_24479);
and U29365 (N_29365,N_23219,N_20911);
nor U29366 (N_29366,N_24151,N_20955);
nand U29367 (N_29367,N_21915,N_22348);
nand U29368 (N_29368,N_24191,N_24149);
or U29369 (N_29369,N_24984,N_24929);
nor U29370 (N_29370,N_24378,N_22342);
or U29371 (N_29371,N_22593,N_20965);
and U29372 (N_29372,N_21497,N_23501);
and U29373 (N_29373,N_24086,N_21489);
xor U29374 (N_29374,N_23571,N_22637);
and U29375 (N_29375,N_21414,N_23648);
nand U29376 (N_29376,N_21809,N_22556);
and U29377 (N_29377,N_23426,N_21215);
nor U29378 (N_29378,N_21623,N_21700);
nand U29379 (N_29379,N_24381,N_24376);
and U29380 (N_29380,N_22952,N_23585);
or U29381 (N_29381,N_23785,N_22221);
xnor U29382 (N_29382,N_21387,N_21451);
or U29383 (N_29383,N_21352,N_20388);
nor U29384 (N_29384,N_22107,N_21565);
xnor U29385 (N_29385,N_23889,N_23777);
xnor U29386 (N_29386,N_21662,N_22651);
and U29387 (N_29387,N_24855,N_21277);
or U29388 (N_29388,N_22881,N_23017);
nand U29389 (N_29389,N_22524,N_20976);
nand U29390 (N_29390,N_22742,N_23612);
and U29391 (N_29391,N_23360,N_23259);
nand U29392 (N_29392,N_23400,N_22365);
nand U29393 (N_29393,N_22874,N_23390);
or U29394 (N_29394,N_23166,N_22294);
nand U29395 (N_29395,N_23094,N_24496);
and U29396 (N_29396,N_23275,N_22571);
or U29397 (N_29397,N_22634,N_23319);
nand U29398 (N_29398,N_24376,N_20860);
nor U29399 (N_29399,N_23378,N_23792);
or U29400 (N_29400,N_22950,N_21608);
nor U29401 (N_29401,N_23926,N_22100);
or U29402 (N_29402,N_21890,N_22177);
xor U29403 (N_29403,N_22376,N_22799);
xor U29404 (N_29404,N_22119,N_24409);
nand U29405 (N_29405,N_24087,N_20094);
nand U29406 (N_29406,N_24519,N_23560);
and U29407 (N_29407,N_21366,N_24257);
nand U29408 (N_29408,N_23328,N_23662);
and U29409 (N_29409,N_21809,N_22203);
and U29410 (N_29410,N_20920,N_24383);
xnor U29411 (N_29411,N_23213,N_22400);
nor U29412 (N_29412,N_24323,N_24235);
nand U29413 (N_29413,N_20836,N_21587);
nand U29414 (N_29414,N_23518,N_24890);
nand U29415 (N_29415,N_20319,N_20266);
or U29416 (N_29416,N_20808,N_21224);
and U29417 (N_29417,N_22036,N_24672);
or U29418 (N_29418,N_24122,N_24200);
and U29419 (N_29419,N_24430,N_24103);
nand U29420 (N_29420,N_20191,N_22720);
nand U29421 (N_29421,N_23071,N_22782);
nand U29422 (N_29422,N_21914,N_24418);
nand U29423 (N_29423,N_23070,N_24616);
xnor U29424 (N_29424,N_24743,N_21353);
xor U29425 (N_29425,N_24329,N_21433);
xor U29426 (N_29426,N_23572,N_20946);
and U29427 (N_29427,N_24380,N_24696);
and U29428 (N_29428,N_21911,N_24036);
or U29429 (N_29429,N_21069,N_20100);
nand U29430 (N_29430,N_23539,N_23352);
nand U29431 (N_29431,N_20308,N_23520);
nor U29432 (N_29432,N_20518,N_21661);
xnor U29433 (N_29433,N_23197,N_22148);
nor U29434 (N_29434,N_24434,N_20139);
nand U29435 (N_29435,N_22901,N_22371);
or U29436 (N_29436,N_23699,N_20256);
nand U29437 (N_29437,N_20290,N_22350);
or U29438 (N_29438,N_23727,N_20681);
xnor U29439 (N_29439,N_21135,N_22516);
nand U29440 (N_29440,N_22691,N_24559);
nor U29441 (N_29441,N_20840,N_24218);
and U29442 (N_29442,N_24144,N_21905);
nand U29443 (N_29443,N_22983,N_22156);
or U29444 (N_29444,N_22159,N_23271);
nor U29445 (N_29445,N_24420,N_20884);
or U29446 (N_29446,N_24089,N_20184);
nor U29447 (N_29447,N_20075,N_20594);
and U29448 (N_29448,N_22060,N_21689);
nand U29449 (N_29449,N_24941,N_22279);
nor U29450 (N_29450,N_23258,N_22203);
and U29451 (N_29451,N_23907,N_24316);
xnor U29452 (N_29452,N_21072,N_21521);
and U29453 (N_29453,N_20811,N_23019);
nand U29454 (N_29454,N_20421,N_21631);
or U29455 (N_29455,N_20926,N_24668);
and U29456 (N_29456,N_22707,N_24815);
or U29457 (N_29457,N_20805,N_21491);
and U29458 (N_29458,N_22650,N_22862);
xnor U29459 (N_29459,N_20615,N_22271);
and U29460 (N_29460,N_21563,N_22051);
xnor U29461 (N_29461,N_21183,N_24370);
and U29462 (N_29462,N_21703,N_23384);
and U29463 (N_29463,N_23069,N_22966);
and U29464 (N_29464,N_20480,N_23502);
nor U29465 (N_29465,N_23946,N_20716);
nand U29466 (N_29466,N_23251,N_24741);
or U29467 (N_29467,N_23003,N_24755);
nor U29468 (N_29468,N_24498,N_22086);
nor U29469 (N_29469,N_20848,N_21693);
and U29470 (N_29470,N_24678,N_22234);
or U29471 (N_29471,N_20048,N_24635);
nor U29472 (N_29472,N_23336,N_21009);
xor U29473 (N_29473,N_21371,N_23967);
and U29474 (N_29474,N_22774,N_20392);
or U29475 (N_29475,N_20190,N_21259);
and U29476 (N_29476,N_22243,N_20515);
and U29477 (N_29477,N_22467,N_21985);
and U29478 (N_29478,N_22870,N_22514);
or U29479 (N_29479,N_21458,N_23903);
or U29480 (N_29480,N_22092,N_22641);
or U29481 (N_29481,N_21901,N_21496);
nor U29482 (N_29482,N_21977,N_23721);
xnor U29483 (N_29483,N_21156,N_21016);
nor U29484 (N_29484,N_24207,N_21664);
xnor U29485 (N_29485,N_22236,N_24868);
or U29486 (N_29486,N_24653,N_20397);
xor U29487 (N_29487,N_22947,N_24102);
nand U29488 (N_29488,N_22802,N_24057);
nor U29489 (N_29489,N_20247,N_21148);
or U29490 (N_29490,N_21811,N_22899);
and U29491 (N_29491,N_24356,N_20884);
nor U29492 (N_29492,N_24820,N_23741);
and U29493 (N_29493,N_20685,N_20207);
or U29494 (N_29494,N_21917,N_22072);
xnor U29495 (N_29495,N_23530,N_22639);
nand U29496 (N_29496,N_23432,N_20573);
xor U29497 (N_29497,N_20340,N_20123);
and U29498 (N_29498,N_23545,N_21066);
and U29499 (N_29499,N_22044,N_20912);
or U29500 (N_29500,N_22269,N_22330);
xnor U29501 (N_29501,N_22473,N_23570);
nor U29502 (N_29502,N_23292,N_21076);
and U29503 (N_29503,N_23926,N_22478);
or U29504 (N_29504,N_22689,N_24237);
nor U29505 (N_29505,N_20754,N_20164);
nor U29506 (N_29506,N_23368,N_24309);
or U29507 (N_29507,N_20740,N_24668);
or U29508 (N_29508,N_24527,N_24228);
and U29509 (N_29509,N_24083,N_21379);
nand U29510 (N_29510,N_24717,N_20191);
nor U29511 (N_29511,N_22116,N_24376);
nor U29512 (N_29512,N_22338,N_20844);
xor U29513 (N_29513,N_20867,N_20682);
nor U29514 (N_29514,N_20930,N_23332);
and U29515 (N_29515,N_21451,N_20562);
nand U29516 (N_29516,N_24582,N_21235);
xnor U29517 (N_29517,N_21229,N_23759);
and U29518 (N_29518,N_21179,N_23635);
nand U29519 (N_29519,N_24503,N_22224);
or U29520 (N_29520,N_20810,N_22566);
nor U29521 (N_29521,N_24436,N_22229);
xnor U29522 (N_29522,N_23127,N_24421);
nand U29523 (N_29523,N_23967,N_22003);
or U29524 (N_29524,N_24650,N_23587);
xor U29525 (N_29525,N_22367,N_23888);
and U29526 (N_29526,N_21700,N_23810);
or U29527 (N_29527,N_22323,N_23683);
or U29528 (N_29528,N_21588,N_22907);
xnor U29529 (N_29529,N_22064,N_20715);
nor U29530 (N_29530,N_23165,N_21525);
and U29531 (N_29531,N_22946,N_20288);
xnor U29532 (N_29532,N_24362,N_20064);
and U29533 (N_29533,N_21531,N_24695);
xor U29534 (N_29534,N_21731,N_23978);
or U29535 (N_29535,N_23817,N_24271);
nand U29536 (N_29536,N_20030,N_21542);
nor U29537 (N_29537,N_22273,N_22062);
xnor U29538 (N_29538,N_20763,N_21198);
or U29539 (N_29539,N_24580,N_23409);
and U29540 (N_29540,N_23201,N_20423);
or U29541 (N_29541,N_22486,N_21809);
or U29542 (N_29542,N_22062,N_20518);
or U29543 (N_29543,N_23395,N_22375);
and U29544 (N_29544,N_24084,N_22668);
nand U29545 (N_29545,N_22845,N_20666);
or U29546 (N_29546,N_24475,N_20412);
and U29547 (N_29547,N_23039,N_22621);
and U29548 (N_29548,N_24142,N_24805);
and U29549 (N_29549,N_20420,N_22743);
and U29550 (N_29550,N_23849,N_24917);
and U29551 (N_29551,N_24479,N_23727);
nor U29552 (N_29552,N_22615,N_23620);
xor U29553 (N_29553,N_23960,N_21373);
nand U29554 (N_29554,N_23481,N_23148);
nand U29555 (N_29555,N_20383,N_20615);
nand U29556 (N_29556,N_23658,N_22498);
nand U29557 (N_29557,N_21644,N_24679);
xor U29558 (N_29558,N_22966,N_22288);
nand U29559 (N_29559,N_22161,N_20823);
or U29560 (N_29560,N_24010,N_21120);
nor U29561 (N_29561,N_23327,N_21577);
nor U29562 (N_29562,N_22651,N_22905);
nand U29563 (N_29563,N_21394,N_23787);
and U29564 (N_29564,N_22709,N_23373);
nand U29565 (N_29565,N_23234,N_21050);
and U29566 (N_29566,N_20036,N_23774);
and U29567 (N_29567,N_23712,N_23318);
xnor U29568 (N_29568,N_23862,N_24045);
and U29569 (N_29569,N_20663,N_23910);
xnor U29570 (N_29570,N_22547,N_20520);
xnor U29571 (N_29571,N_22871,N_22331);
or U29572 (N_29572,N_23146,N_22632);
nand U29573 (N_29573,N_22918,N_24120);
nand U29574 (N_29574,N_22546,N_23078);
nand U29575 (N_29575,N_20542,N_24533);
nand U29576 (N_29576,N_20562,N_21920);
and U29577 (N_29577,N_24883,N_20819);
or U29578 (N_29578,N_21566,N_23292);
or U29579 (N_29579,N_23449,N_20510);
xor U29580 (N_29580,N_22283,N_20845);
nand U29581 (N_29581,N_24456,N_20288);
or U29582 (N_29582,N_20387,N_23254);
nand U29583 (N_29583,N_20028,N_22514);
nand U29584 (N_29584,N_23671,N_20239);
xor U29585 (N_29585,N_22367,N_23026);
and U29586 (N_29586,N_24475,N_21354);
xor U29587 (N_29587,N_23178,N_21375);
and U29588 (N_29588,N_20691,N_21111);
and U29589 (N_29589,N_21029,N_20239);
or U29590 (N_29590,N_21836,N_21177);
xor U29591 (N_29591,N_21584,N_22308);
nand U29592 (N_29592,N_21288,N_21779);
nand U29593 (N_29593,N_21506,N_21277);
xnor U29594 (N_29594,N_21473,N_22393);
or U29595 (N_29595,N_21036,N_24566);
or U29596 (N_29596,N_23702,N_23231);
nor U29597 (N_29597,N_24638,N_20244);
or U29598 (N_29598,N_22612,N_23721);
nor U29599 (N_29599,N_24385,N_23796);
nor U29600 (N_29600,N_21474,N_24450);
nand U29601 (N_29601,N_20524,N_20022);
nor U29602 (N_29602,N_23990,N_23604);
or U29603 (N_29603,N_24377,N_22618);
nand U29604 (N_29604,N_24367,N_20004);
and U29605 (N_29605,N_24241,N_21118);
nand U29606 (N_29606,N_20553,N_20203);
xor U29607 (N_29607,N_24562,N_24262);
or U29608 (N_29608,N_21938,N_23964);
nand U29609 (N_29609,N_20243,N_23985);
nor U29610 (N_29610,N_20646,N_21989);
and U29611 (N_29611,N_21448,N_21567);
nor U29612 (N_29612,N_24090,N_21109);
and U29613 (N_29613,N_24502,N_21857);
or U29614 (N_29614,N_24143,N_20671);
nor U29615 (N_29615,N_21032,N_20898);
nand U29616 (N_29616,N_24285,N_24703);
or U29617 (N_29617,N_23386,N_23324);
or U29618 (N_29618,N_23419,N_21543);
and U29619 (N_29619,N_23585,N_21517);
and U29620 (N_29620,N_20355,N_22615);
or U29621 (N_29621,N_21989,N_20023);
or U29622 (N_29622,N_24073,N_24220);
nand U29623 (N_29623,N_23229,N_21331);
nor U29624 (N_29624,N_20001,N_23480);
and U29625 (N_29625,N_20075,N_23710);
nand U29626 (N_29626,N_23436,N_21208);
and U29627 (N_29627,N_24635,N_24753);
xor U29628 (N_29628,N_22290,N_22324);
and U29629 (N_29629,N_24726,N_23077);
xnor U29630 (N_29630,N_24802,N_22571);
nand U29631 (N_29631,N_23516,N_24820);
or U29632 (N_29632,N_24645,N_20180);
nor U29633 (N_29633,N_24181,N_21983);
xor U29634 (N_29634,N_21086,N_21858);
or U29635 (N_29635,N_22620,N_24033);
nor U29636 (N_29636,N_20654,N_24323);
or U29637 (N_29637,N_23562,N_23416);
or U29638 (N_29638,N_23161,N_21059);
and U29639 (N_29639,N_22289,N_24493);
xor U29640 (N_29640,N_22445,N_20941);
and U29641 (N_29641,N_20507,N_20136);
xor U29642 (N_29642,N_23964,N_22829);
nor U29643 (N_29643,N_23880,N_22225);
xor U29644 (N_29644,N_24443,N_21845);
or U29645 (N_29645,N_24522,N_23372);
nand U29646 (N_29646,N_21672,N_22793);
xor U29647 (N_29647,N_21482,N_23539);
and U29648 (N_29648,N_22774,N_21185);
or U29649 (N_29649,N_22950,N_20354);
nor U29650 (N_29650,N_20283,N_23105);
xnor U29651 (N_29651,N_20951,N_24266);
or U29652 (N_29652,N_24952,N_23611);
and U29653 (N_29653,N_20007,N_23580);
or U29654 (N_29654,N_24535,N_23783);
xnor U29655 (N_29655,N_23349,N_20624);
and U29656 (N_29656,N_23738,N_23934);
and U29657 (N_29657,N_24892,N_22443);
nor U29658 (N_29658,N_20506,N_22980);
nand U29659 (N_29659,N_24301,N_23110);
nor U29660 (N_29660,N_21274,N_23943);
or U29661 (N_29661,N_22463,N_21904);
or U29662 (N_29662,N_21396,N_23497);
and U29663 (N_29663,N_23265,N_22756);
and U29664 (N_29664,N_20528,N_21473);
xor U29665 (N_29665,N_20431,N_21055);
and U29666 (N_29666,N_21900,N_20971);
or U29667 (N_29667,N_22109,N_24921);
or U29668 (N_29668,N_20052,N_22499);
nand U29669 (N_29669,N_20483,N_24906);
and U29670 (N_29670,N_23291,N_24289);
and U29671 (N_29671,N_24629,N_22854);
nor U29672 (N_29672,N_22698,N_23675);
or U29673 (N_29673,N_23949,N_23735);
nor U29674 (N_29674,N_23113,N_23358);
or U29675 (N_29675,N_24794,N_22694);
or U29676 (N_29676,N_21196,N_23488);
nor U29677 (N_29677,N_22124,N_23259);
and U29678 (N_29678,N_23793,N_24108);
xor U29679 (N_29679,N_23913,N_22439);
nor U29680 (N_29680,N_24796,N_20756);
nor U29681 (N_29681,N_24948,N_20583);
and U29682 (N_29682,N_22735,N_21443);
or U29683 (N_29683,N_23861,N_23242);
and U29684 (N_29684,N_24782,N_23543);
xnor U29685 (N_29685,N_20564,N_20235);
or U29686 (N_29686,N_23344,N_24322);
xnor U29687 (N_29687,N_22557,N_24687);
xor U29688 (N_29688,N_20230,N_21235);
xor U29689 (N_29689,N_24212,N_24108);
nor U29690 (N_29690,N_21022,N_21353);
nor U29691 (N_29691,N_20402,N_22321);
nand U29692 (N_29692,N_24646,N_20156);
xnor U29693 (N_29693,N_21648,N_22632);
and U29694 (N_29694,N_23652,N_22768);
and U29695 (N_29695,N_22963,N_23159);
nand U29696 (N_29696,N_24376,N_21731);
or U29697 (N_29697,N_23530,N_22857);
nand U29698 (N_29698,N_23212,N_24055);
nand U29699 (N_29699,N_21107,N_21995);
nand U29700 (N_29700,N_24910,N_23182);
xnor U29701 (N_29701,N_24139,N_24190);
xnor U29702 (N_29702,N_23360,N_23254);
nor U29703 (N_29703,N_21780,N_24877);
or U29704 (N_29704,N_20071,N_20473);
and U29705 (N_29705,N_22473,N_23530);
nand U29706 (N_29706,N_21950,N_23227);
nor U29707 (N_29707,N_24703,N_24751);
or U29708 (N_29708,N_23716,N_24337);
or U29709 (N_29709,N_22977,N_24733);
xor U29710 (N_29710,N_24046,N_24733);
and U29711 (N_29711,N_24021,N_22713);
and U29712 (N_29712,N_22528,N_24574);
nor U29713 (N_29713,N_22989,N_22239);
nor U29714 (N_29714,N_24247,N_23520);
xnor U29715 (N_29715,N_21186,N_20368);
or U29716 (N_29716,N_21311,N_22118);
or U29717 (N_29717,N_21294,N_22953);
nor U29718 (N_29718,N_24543,N_24721);
xnor U29719 (N_29719,N_21676,N_23876);
and U29720 (N_29720,N_22281,N_24702);
nor U29721 (N_29721,N_20174,N_23331);
nor U29722 (N_29722,N_24791,N_24066);
nor U29723 (N_29723,N_23831,N_23546);
xnor U29724 (N_29724,N_20894,N_22229);
nand U29725 (N_29725,N_21954,N_22530);
xor U29726 (N_29726,N_24947,N_24807);
nand U29727 (N_29727,N_22482,N_24952);
and U29728 (N_29728,N_21506,N_20265);
xor U29729 (N_29729,N_24705,N_22965);
and U29730 (N_29730,N_23593,N_23412);
nand U29731 (N_29731,N_24468,N_20311);
nor U29732 (N_29732,N_21273,N_22831);
nand U29733 (N_29733,N_24816,N_22253);
or U29734 (N_29734,N_22814,N_24732);
nand U29735 (N_29735,N_20738,N_21356);
xnor U29736 (N_29736,N_23951,N_20840);
nand U29737 (N_29737,N_22492,N_23757);
nor U29738 (N_29738,N_24948,N_23203);
and U29739 (N_29739,N_22769,N_21371);
nor U29740 (N_29740,N_23494,N_24823);
xor U29741 (N_29741,N_21063,N_23856);
and U29742 (N_29742,N_20953,N_23611);
xor U29743 (N_29743,N_24582,N_23243);
nand U29744 (N_29744,N_21774,N_24687);
nor U29745 (N_29745,N_20020,N_23444);
nand U29746 (N_29746,N_24464,N_22945);
and U29747 (N_29747,N_22269,N_22035);
and U29748 (N_29748,N_23606,N_23029);
and U29749 (N_29749,N_21198,N_23207);
nor U29750 (N_29750,N_22082,N_21352);
nand U29751 (N_29751,N_21318,N_23529);
nor U29752 (N_29752,N_20442,N_20206);
nor U29753 (N_29753,N_21583,N_24928);
nand U29754 (N_29754,N_23336,N_23100);
nand U29755 (N_29755,N_20359,N_23532);
nor U29756 (N_29756,N_20114,N_24465);
nand U29757 (N_29757,N_20107,N_24019);
and U29758 (N_29758,N_21135,N_24347);
nor U29759 (N_29759,N_20697,N_24325);
and U29760 (N_29760,N_20874,N_22702);
nand U29761 (N_29761,N_23993,N_22712);
nor U29762 (N_29762,N_24379,N_20459);
and U29763 (N_29763,N_20568,N_21888);
xnor U29764 (N_29764,N_21055,N_21370);
or U29765 (N_29765,N_20081,N_24203);
and U29766 (N_29766,N_24341,N_20648);
nand U29767 (N_29767,N_21440,N_23181);
and U29768 (N_29768,N_20052,N_20760);
and U29769 (N_29769,N_21028,N_22078);
and U29770 (N_29770,N_24220,N_23307);
xnor U29771 (N_29771,N_22676,N_23504);
xnor U29772 (N_29772,N_24142,N_22572);
xnor U29773 (N_29773,N_22592,N_22966);
nor U29774 (N_29774,N_21232,N_24894);
nand U29775 (N_29775,N_24529,N_21589);
or U29776 (N_29776,N_23002,N_20458);
nor U29777 (N_29777,N_20663,N_24292);
nor U29778 (N_29778,N_20189,N_20850);
nor U29779 (N_29779,N_22457,N_22742);
and U29780 (N_29780,N_23479,N_21595);
nand U29781 (N_29781,N_21832,N_23811);
or U29782 (N_29782,N_22986,N_23556);
or U29783 (N_29783,N_23962,N_22894);
and U29784 (N_29784,N_20104,N_20307);
and U29785 (N_29785,N_21348,N_24901);
xor U29786 (N_29786,N_21625,N_23338);
nand U29787 (N_29787,N_22771,N_24401);
nor U29788 (N_29788,N_24049,N_24812);
xor U29789 (N_29789,N_21213,N_24634);
xnor U29790 (N_29790,N_21320,N_22552);
nor U29791 (N_29791,N_21975,N_20809);
nor U29792 (N_29792,N_20985,N_22990);
or U29793 (N_29793,N_24798,N_21370);
and U29794 (N_29794,N_21277,N_24932);
or U29795 (N_29795,N_23793,N_20720);
nand U29796 (N_29796,N_24483,N_20032);
nor U29797 (N_29797,N_23984,N_20906);
nand U29798 (N_29798,N_20944,N_21889);
or U29799 (N_29799,N_22663,N_21018);
xor U29800 (N_29800,N_21753,N_22186);
and U29801 (N_29801,N_23271,N_23454);
and U29802 (N_29802,N_22450,N_23637);
xnor U29803 (N_29803,N_23811,N_22487);
nor U29804 (N_29804,N_24365,N_20662);
nor U29805 (N_29805,N_23890,N_22768);
and U29806 (N_29806,N_24000,N_21150);
xor U29807 (N_29807,N_20015,N_24242);
or U29808 (N_29808,N_22181,N_20931);
or U29809 (N_29809,N_20267,N_22395);
or U29810 (N_29810,N_21183,N_20741);
nand U29811 (N_29811,N_20707,N_21948);
and U29812 (N_29812,N_23526,N_24361);
or U29813 (N_29813,N_23818,N_20824);
nor U29814 (N_29814,N_24558,N_23588);
xor U29815 (N_29815,N_21219,N_20743);
xor U29816 (N_29816,N_22300,N_20280);
nand U29817 (N_29817,N_23656,N_24676);
nor U29818 (N_29818,N_21946,N_20870);
nor U29819 (N_29819,N_23773,N_23272);
xnor U29820 (N_29820,N_23164,N_20458);
and U29821 (N_29821,N_24177,N_24062);
nor U29822 (N_29822,N_20914,N_20169);
xor U29823 (N_29823,N_24462,N_20237);
and U29824 (N_29824,N_21270,N_21747);
and U29825 (N_29825,N_23475,N_20273);
xnor U29826 (N_29826,N_22829,N_20852);
nor U29827 (N_29827,N_24385,N_22909);
and U29828 (N_29828,N_21976,N_23025);
or U29829 (N_29829,N_22491,N_22577);
nor U29830 (N_29830,N_21903,N_23943);
xnor U29831 (N_29831,N_20346,N_21109);
nand U29832 (N_29832,N_20758,N_20068);
nor U29833 (N_29833,N_20829,N_21396);
nor U29834 (N_29834,N_20242,N_23718);
and U29835 (N_29835,N_23450,N_20035);
and U29836 (N_29836,N_23702,N_20394);
and U29837 (N_29837,N_24302,N_24558);
or U29838 (N_29838,N_21885,N_21936);
and U29839 (N_29839,N_20768,N_21234);
nand U29840 (N_29840,N_21711,N_23126);
and U29841 (N_29841,N_21670,N_23477);
xnor U29842 (N_29842,N_20172,N_23696);
or U29843 (N_29843,N_21063,N_21400);
xor U29844 (N_29844,N_20577,N_21215);
nand U29845 (N_29845,N_24809,N_24093);
nand U29846 (N_29846,N_24164,N_24647);
xnor U29847 (N_29847,N_24269,N_23369);
nand U29848 (N_29848,N_21948,N_23763);
and U29849 (N_29849,N_22411,N_22178);
and U29850 (N_29850,N_21441,N_20056);
and U29851 (N_29851,N_20106,N_20055);
or U29852 (N_29852,N_24237,N_20167);
or U29853 (N_29853,N_22729,N_20591);
or U29854 (N_29854,N_22633,N_20037);
and U29855 (N_29855,N_20597,N_20715);
nor U29856 (N_29856,N_20522,N_24063);
nand U29857 (N_29857,N_24204,N_22082);
or U29858 (N_29858,N_22370,N_22561);
nor U29859 (N_29859,N_21649,N_21574);
or U29860 (N_29860,N_24533,N_22935);
or U29861 (N_29861,N_23695,N_21497);
xnor U29862 (N_29862,N_22796,N_21555);
and U29863 (N_29863,N_23887,N_21181);
nor U29864 (N_29864,N_21023,N_24047);
or U29865 (N_29865,N_22766,N_23051);
or U29866 (N_29866,N_20094,N_24301);
xor U29867 (N_29867,N_24904,N_22727);
nand U29868 (N_29868,N_23096,N_23758);
or U29869 (N_29869,N_20354,N_20976);
nand U29870 (N_29870,N_22673,N_24762);
nor U29871 (N_29871,N_23064,N_20133);
xnor U29872 (N_29872,N_23306,N_22639);
or U29873 (N_29873,N_24813,N_23652);
nand U29874 (N_29874,N_23870,N_21877);
or U29875 (N_29875,N_23985,N_21995);
nor U29876 (N_29876,N_24886,N_22122);
and U29877 (N_29877,N_20820,N_21675);
nand U29878 (N_29878,N_20110,N_20476);
nand U29879 (N_29879,N_20996,N_23593);
and U29880 (N_29880,N_20646,N_21664);
and U29881 (N_29881,N_24109,N_21871);
nor U29882 (N_29882,N_20030,N_23862);
nand U29883 (N_29883,N_24056,N_24521);
nand U29884 (N_29884,N_20999,N_21608);
and U29885 (N_29885,N_24781,N_20566);
xor U29886 (N_29886,N_20675,N_23212);
xnor U29887 (N_29887,N_22629,N_23722);
and U29888 (N_29888,N_20314,N_20688);
nand U29889 (N_29889,N_21884,N_23850);
nand U29890 (N_29890,N_22067,N_21767);
nor U29891 (N_29891,N_23847,N_22587);
nor U29892 (N_29892,N_23026,N_21099);
xnor U29893 (N_29893,N_22545,N_24916);
nand U29894 (N_29894,N_24013,N_20971);
nand U29895 (N_29895,N_23061,N_23038);
nor U29896 (N_29896,N_20321,N_24837);
nor U29897 (N_29897,N_22436,N_24247);
nor U29898 (N_29898,N_22547,N_24427);
nor U29899 (N_29899,N_21646,N_22460);
or U29900 (N_29900,N_23030,N_22177);
nand U29901 (N_29901,N_21810,N_20022);
nand U29902 (N_29902,N_21406,N_22244);
nand U29903 (N_29903,N_20019,N_24425);
nor U29904 (N_29904,N_23548,N_22874);
xnor U29905 (N_29905,N_21115,N_21436);
or U29906 (N_29906,N_20145,N_21990);
nand U29907 (N_29907,N_21703,N_21378);
and U29908 (N_29908,N_24827,N_22117);
xnor U29909 (N_29909,N_23501,N_21646);
or U29910 (N_29910,N_22929,N_21495);
xor U29911 (N_29911,N_22414,N_20548);
nor U29912 (N_29912,N_24042,N_24936);
and U29913 (N_29913,N_21626,N_24539);
nor U29914 (N_29914,N_23301,N_22352);
nor U29915 (N_29915,N_23287,N_23464);
nand U29916 (N_29916,N_24848,N_23319);
xor U29917 (N_29917,N_21240,N_20758);
nor U29918 (N_29918,N_20986,N_22174);
or U29919 (N_29919,N_20093,N_21445);
and U29920 (N_29920,N_21481,N_21922);
or U29921 (N_29921,N_21132,N_20222);
or U29922 (N_29922,N_22307,N_23341);
or U29923 (N_29923,N_20476,N_23602);
xnor U29924 (N_29924,N_23831,N_22770);
and U29925 (N_29925,N_24524,N_23959);
and U29926 (N_29926,N_20473,N_20686);
and U29927 (N_29927,N_21858,N_21111);
xnor U29928 (N_29928,N_23600,N_20040);
and U29929 (N_29929,N_21775,N_22979);
xor U29930 (N_29930,N_22496,N_20215);
nor U29931 (N_29931,N_21203,N_24485);
and U29932 (N_29932,N_23845,N_24310);
and U29933 (N_29933,N_23692,N_21958);
and U29934 (N_29934,N_23647,N_21511);
nand U29935 (N_29935,N_21404,N_22243);
or U29936 (N_29936,N_21400,N_24138);
nor U29937 (N_29937,N_24908,N_20290);
and U29938 (N_29938,N_24045,N_21134);
and U29939 (N_29939,N_22390,N_21387);
or U29940 (N_29940,N_24286,N_24341);
or U29941 (N_29941,N_23798,N_21282);
nand U29942 (N_29942,N_22594,N_23499);
nor U29943 (N_29943,N_20049,N_23727);
xor U29944 (N_29944,N_21797,N_20261);
and U29945 (N_29945,N_23826,N_24984);
nor U29946 (N_29946,N_21010,N_24008);
nand U29947 (N_29947,N_22948,N_22539);
and U29948 (N_29948,N_21123,N_23849);
or U29949 (N_29949,N_22422,N_23701);
nand U29950 (N_29950,N_22133,N_21987);
and U29951 (N_29951,N_22809,N_22781);
nand U29952 (N_29952,N_24457,N_22609);
or U29953 (N_29953,N_24397,N_20986);
and U29954 (N_29954,N_20871,N_22282);
xor U29955 (N_29955,N_24621,N_22073);
nor U29956 (N_29956,N_23938,N_21604);
and U29957 (N_29957,N_20883,N_24197);
nor U29958 (N_29958,N_20627,N_22710);
nand U29959 (N_29959,N_21067,N_21861);
xor U29960 (N_29960,N_23800,N_20103);
nor U29961 (N_29961,N_23637,N_24884);
and U29962 (N_29962,N_21940,N_22463);
nor U29963 (N_29963,N_20471,N_23940);
nand U29964 (N_29964,N_23635,N_20726);
nor U29965 (N_29965,N_22690,N_23214);
nor U29966 (N_29966,N_24959,N_20556);
xor U29967 (N_29967,N_24878,N_22310);
or U29968 (N_29968,N_23287,N_22340);
xnor U29969 (N_29969,N_24729,N_24794);
or U29970 (N_29970,N_22940,N_21214);
and U29971 (N_29971,N_24668,N_24352);
nand U29972 (N_29972,N_23247,N_24104);
nor U29973 (N_29973,N_21370,N_24550);
or U29974 (N_29974,N_21933,N_21445);
and U29975 (N_29975,N_23655,N_20615);
xor U29976 (N_29976,N_24523,N_23737);
nand U29977 (N_29977,N_21877,N_21745);
nand U29978 (N_29978,N_24247,N_21742);
and U29979 (N_29979,N_24620,N_20253);
and U29980 (N_29980,N_21025,N_24160);
xor U29981 (N_29981,N_20464,N_22913);
or U29982 (N_29982,N_20671,N_21310);
xnor U29983 (N_29983,N_22485,N_22642);
and U29984 (N_29984,N_21609,N_20845);
nor U29985 (N_29985,N_22979,N_24964);
xnor U29986 (N_29986,N_23211,N_24280);
xor U29987 (N_29987,N_24218,N_23702);
nor U29988 (N_29988,N_22233,N_23796);
and U29989 (N_29989,N_20231,N_22323);
and U29990 (N_29990,N_22798,N_22060);
nand U29991 (N_29991,N_24708,N_22245);
and U29992 (N_29992,N_23983,N_22148);
nor U29993 (N_29993,N_20518,N_21406);
or U29994 (N_29994,N_23876,N_21040);
nor U29995 (N_29995,N_21625,N_22215);
xnor U29996 (N_29996,N_24248,N_23043);
nor U29997 (N_29997,N_20729,N_21841);
nor U29998 (N_29998,N_20655,N_20520);
or U29999 (N_29999,N_23198,N_24794);
nand U30000 (N_30000,N_27187,N_26776);
nor U30001 (N_30001,N_27182,N_28714);
or U30002 (N_30002,N_26634,N_29714);
and U30003 (N_30003,N_28951,N_28547);
nor U30004 (N_30004,N_25616,N_29237);
or U30005 (N_30005,N_29069,N_25848);
xnor U30006 (N_30006,N_27419,N_25420);
or U30007 (N_30007,N_25439,N_25106);
nand U30008 (N_30008,N_25510,N_27003);
or U30009 (N_30009,N_28398,N_27408);
or U30010 (N_30010,N_27903,N_26720);
and U30011 (N_30011,N_29864,N_25746);
or U30012 (N_30012,N_26402,N_27467);
xor U30013 (N_30013,N_28595,N_29632);
or U30014 (N_30014,N_25727,N_27781);
nand U30015 (N_30015,N_29268,N_26509);
nor U30016 (N_30016,N_28655,N_29269);
nor U30017 (N_30017,N_25118,N_26407);
xnor U30018 (N_30018,N_27483,N_29961);
xnor U30019 (N_30019,N_28414,N_29896);
nor U30020 (N_30020,N_29034,N_26123);
or U30021 (N_30021,N_25661,N_27193);
or U30022 (N_30022,N_28337,N_29169);
or U30023 (N_30023,N_27041,N_26583);
nand U30024 (N_30024,N_26263,N_27212);
nand U30025 (N_30025,N_28639,N_26164);
nor U30026 (N_30026,N_26086,N_25315);
nand U30027 (N_30027,N_27090,N_29182);
and U30028 (N_30028,N_27963,N_29854);
xnor U30029 (N_30029,N_29634,N_27162);
and U30030 (N_30030,N_26243,N_29425);
xnor U30031 (N_30031,N_29151,N_25790);
nor U30032 (N_30032,N_27753,N_27073);
xnor U30033 (N_30033,N_25016,N_28095);
nor U30034 (N_30034,N_25429,N_28966);
nor U30035 (N_30035,N_28082,N_28188);
xnor U30036 (N_30036,N_29116,N_28368);
or U30037 (N_30037,N_26866,N_25302);
nor U30038 (N_30038,N_29023,N_28142);
or U30039 (N_30039,N_26721,N_28262);
and U30040 (N_30040,N_29444,N_29316);
xnor U30041 (N_30041,N_29000,N_25215);
nor U30042 (N_30042,N_25276,N_28111);
nor U30043 (N_30043,N_27884,N_29903);
and U30044 (N_30044,N_26248,N_26745);
xor U30045 (N_30045,N_29476,N_26504);
or U30046 (N_30046,N_25541,N_28464);
nand U30047 (N_30047,N_29304,N_26681);
xnor U30048 (N_30048,N_28386,N_26194);
and U30049 (N_30049,N_25651,N_29134);
xor U30050 (N_30050,N_27678,N_28164);
nand U30051 (N_30051,N_27831,N_26047);
nor U30052 (N_30052,N_25702,N_29335);
nor U30053 (N_30053,N_27733,N_28751);
xnor U30054 (N_30054,N_28820,N_27420);
nand U30055 (N_30055,N_25239,N_29489);
xor U30056 (N_30056,N_27741,N_28850);
xor U30057 (N_30057,N_28048,N_27142);
or U30058 (N_30058,N_25491,N_29306);
nor U30059 (N_30059,N_29996,N_29827);
xor U30060 (N_30060,N_28287,N_25299);
nand U30061 (N_30061,N_26452,N_29581);
nand U30062 (N_30062,N_25354,N_27308);
nand U30063 (N_30063,N_26110,N_25117);
and U30064 (N_30064,N_28317,N_26840);
nor U30065 (N_30065,N_26401,N_29358);
nand U30066 (N_30066,N_25130,N_26844);
nor U30067 (N_30067,N_29437,N_28955);
nor U30068 (N_30068,N_25447,N_26804);
and U30069 (N_30069,N_26961,N_25151);
or U30070 (N_30070,N_28072,N_28681);
nor U30071 (N_30071,N_27621,N_29064);
and U30072 (N_30072,N_25278,N_26555);
nor U30073 (N_30073,N_28268,N_29748);
nand U30074 (N_30074,N_28073,N_26307);
or U30075 (N_30075,N_27188,N_26706);
xor U30076 (N_30076,N_27439,N_28663);
nor U30077 (N_30077,N_27024,N_27786);
xor U30078 (N_30078,N_26601,N_26169);
or U30079 (N_30079,N_28996,N_25891);
nand U30080 (N_30080,N_25163,N_29041);
nor U30081 (N_30081,N_27295,N_28774);
nor U30082 (N_30082,N_28668,N_27471);
xnor U30083 (N_30083,N_25542,N_27201);
or U30084 (N_30084,N_29014,N_29773);
and U30085 (N_30085,N_29716,N_28030);
xnor U30086 (N_30086,N_25546,N_26682);
and U30087 (N_30087,N_25578,N_26995);
xnor U30088 (N_30088,N_27738,N_28447);
nand U30089 (N_30089,N_27102,N_28840);
nand U30090 (N_30090,N_27320,N_26278);
and U30091 (N_30091,N_27055,N_25935);
nor U30092 (N_30092,N_26136,N_26620);
or U30093 (N_30093,N_26596,N_29969);
xor U30094 (N_30094,N_25605,N_25360);
nand U30095 (N_30095,N_26696,N_27424);
nand U30096 (N_30096,N_28504,N_28146);
nor U30097 (N_30097,N_28734,N_27523);
nand U30098 (N_30098,N_28785,N_27402);
xnor U30099 (N_30099,N_26349,N_27821);
and U30100 (N_30100,N_28068,N_27005);
or U30101 (N_30101,N_26111,N_26815);
or U30102 (N_30102,N_26109,N_27986);
nor U30103 (N_30103,N_25824,N_26965);
and U30104 (N_30104,N_26883,N_27018);
nor U30105 (N_30105,N_25960,N_26606);
nand U30106 (N_30106,N_27338,N_27504);
nor U30107 (N_30107,N_27575,N_29627);
xor U30108 (N_30108,N_28715,N_25703);
xor U30109 (N_30109,N_27530,N_28586);
and U30110 (N_30110,N_29541,N_25245);
and U30111 (N_30111,N_26004,N_26302);
nor U30112 (N_30112,N_28013,N_28281);
or U30113 (N_30113,N_27353,N_27837);
nand U30114 (N_30114,N_27877,N_26030);
nand U30115 (N_30115,N_26912,N_29689);
or U30116 (N_30116,N_28390,N_29284);
xor U30117 (N_30117,N_26587,N_26808);
or U30118 (N_30118,N_28041,N_27694);
or U30119 (N_30119,N_28837,N_29641);
or U30120 (N_30120,N_27956,N_26408);
or U30121 (N_30121,N_29285,N_29510);
xnor U30122 (N_30122,N_28454,N_26143);
nand U30123 (N_30123,N_29668,N_26257);
or U30124 (N_30124,N_26638,N_25431);
xor U30125 (N_30125,N_26385,N_29958);
or U30126 (N_30126,N_27568,N_27824);
nor U30127 (N_30127,N_27836,N_25224);
and U30128 (N_30128,N_29338,N_28886);
nand U30129 (N_30129,N_29520,N_26274);
and U30130 (N_30130,N_29110,N_26919);
xnor U30131 (N_30131,N_29068,N_26898);
or U30132 (N_30132,N_29459,N_26035);
xnor U30133 (N_30133,N_29382,N_29059);
nand U30134 (N_30134,N_26139,N_25309);
nand U30135 (N_30135,N_25059,N_29652);
or U30136 (N_30136,N_26201,N_27995);
nor U30137 (N_30137,N_29712,N_29238);
nor U30138 (N_30138,N_26911,N_29600);
and U30139 (N_30139,N_27199,N_27728);
and U30140 (N_30140,N_25248,N_28669);
or U30141 (N_30141,N_27748,N_26447);
nor U30142 (N_30142,N_28144,N_28795);
nor U30143 (N_30143,N_25110,N_28508);
nor U30144 (N_30144,N_25346,N_25290);
xnor U30145 (N_30145,N_28762,N_28677);
xor U30146 (N_30146,N_29767,N_28309);
nor U30147 (N_30147,N_28129,N_27131);
or U30148 (N_30148,N_28989,N_27804);
or U30149 (N_30149,N_25197,N_25619);
xnor U30150 (N_30150,N_27885,N_28195);
nand U30151 (N_30151,N_29163,N_27444);
and U30152 (N_30152,N_29149,N_27448);
or U30153 (N_30153,N_28744,N_26099);
or U30154 (N_30154,N_25580,N_28573);
and U30155 (N_30155,N_26070,N_26975);
or U30156 (N_30156,N_25018,N_27239);
nand U30157 (N_30157,N_27278,N_26531);
xnor U30158 (N_30158,N_27640,N_27426);
and U30159 (N_30159,N_29988,N_27503);
or U30160 (N_30160,N_25423,N_28786);
or U30161 (N_30161,N_26432,N_26842);
nor U30162 (N_30162,N_28849,N_27272);
nand U30163 (N_30163,N_28599,N_29575);
xor U30164 (N_30164,N_28866,N_29866);
nand U30165 (N_30165,N_26137,N_28884);
nor U30166 (N_30166,N_29620,N_27019);
nand U30167 (N_30167,N_29883,N_25774);
or U30168 (N_30168,N_26865,N_26737);
nand U30169 (N_30169,N_26436,N_29914);
or U30170 (N_30170,N_26183,N_29047);
or U30171 (N_30171,N_25020,N_25052);
nor U30172 (N_30172,N_29667,N_26062);
and U30173 (N_30173,N_26803,N_28332);
and U30174 (N_30174,N_27729,N_25840);
or U30175 (N_30175,N_26065,N_28151);
or U30176 (N_30176,N_27871,N_26314);
nor U30177 (N_30177,N_28721,N_25187);
nand U30178 (N_30178,N_27985,N_25630);
xor U30179 (N_30179,N_26820,N_29891);
or U30180 (N_30180,N_27259,N_27511);
and U30181 (N_30181,N_29131,N_29192);
nor U30182 (N_30182,N_29436,N_27614);
nor U30183 (N_30183,N_27765,N_27153);
xnor U30184 (N_30184,N_29043,N_27326);
xor U30185 (N_30185,N_26202,N_25701);
xor U30186 (N_30186,N_29421,N_25126);
and U30187 (N_30187,N_25634,N_25484);
and U30188 (N_30188,N_25000,N_28790);
nand U30189 (N_30189,N_28781,N_28004);
xnor U30190 (N_30190,N_29823,N_29953);
nor U30191 (N_30191,N_29533,N_29884);
xor U30192 (N_30192,N_26569,N_27542);
or U30193 (N_30193,N_29147,N_27442);
xor U30194 (N_30194,N_28661,N_25244);
xnor U30195 (N_30195,N_29579,N_25709);
xor U30196 (N_30196,N_25614,N_27251);
or U30197 (N_30197,N_25322,N_26417);
or U30198 (N_30198,N_28415,N_29647);
or U30199 (N_30199,N_29311,N_28127);
nand U30200 (N_30200,N_27797,N_25228);
or U30201 (N_30201,N_25767,N_25449);
nand U30202 (N_30202,N_26433,N_29949);
nor U30203 (N_30203,N_29056,N_27715);
xnor U30204 (N_30204,N_28488,N_27709);
xor U30205 (N_30205,N_25919,N_29152);
xnor U30206 (N_30206,N_26541,N_27888);
or U30207 (N_30207,N_26480,N_28024);
xnor U30208 (N_30208,N_27927,N_26394);
nor U30209 (N_30209,N_25738,N_28394);
nor U30210 (N_30210,N_26625,N_27116);
or U30211 (N_30211,N_25850,N_25008);
xor U30212 (N_30212,N_25168,N_28061);
nand U30213 (N_30213,N_25830,N_27100);
or U30214 (N_30214,N_25178,N_28437);
nand U30215 (N_30215,N_26933,N_25185);
nand U30216 (N_30216,N_28301,N_27834);
nor U30217 (N_30217,N_28474,N_28374);
xnor U30218 (N_30218,N_26475,N_27565);
or U30219 (N_30219,N_25035,N_26585);
xor U30220 (N_30220,N_27793,N_28456);
nor U30221 (N_30221,N_26337,N_29099);
nand U30222 (N_30222,N_25789,N_25582);
nand U30223 (N_30223,N_27016,N_25623);
nor U30224 (N_30224,N_27304,N_29591);
and U30225 (N_30225,N_25895,N_28703);
or U30226 (N_30226,N_27132,N_25884);
nor U30227 (N_30227,N_29720,N_27384);
nand U30228 (N_30228,N_28887,N_25921);
nor U30229 (N_30229,N_28376,N_26484);
and U30230 (N_30230,N_25109,N_28308);
nand U30231 (N_30231,N_27790,N_29211);
and U30232 (N_30232,N_29951,N_28888);
xor U30233 (N_30233,N_29062,N_29010);
and U30234 (N_30234,N_28355,N_25162);
and U30235 (N_30235,N_25900,N_25535);
or U30236 (N_30236,N_26542,N_28701);
nor U30237 (N_30237,N_27962,N_28782);
nand U30238 (N_30238,N_29474,N_29717);
xor U30239 (N_30239,N_26594,N_27763);
xor U30240 (N_30240,N_25877,N_29218);
nand U30241 (N_30241,N_29628,N_28286);
nor U30242 (N_30242,N_29126,N_25441);
nand U30243 (N_30243,N_29747,N_27250);
nor U30244 (N_30244,N_27128,N_28976);
or U30245 (N_30245,N_25514,N_25913);
or U30246 (N_30246,N_27161,N_27376);
nand U30247 (N_30247,N_27436,N_25385);
and U30248 (N_30248,N_25205,N_26930);
nor U30249 (N_30249,N_27261,N_26879);
nand U30250 (N_30250,N_26245,N_26695);
nand U30251 (N_30251,N_25656,N_29550);
or U30252 (N_30252,N_28426,N_26175);
nor U30253 (N_30253,N_28618,N_27996);
xor U30254 (N_30254,N_25925,N_28865);
or U30255 (N_30255,N_27392,N_26896);
and U30256 (N_30256,N_25140,N_25355);
nand U30257 (N_30257,N_26924,N_28333);
xor U30258 (N_30258,N_27566,N_28638);
nor U30259 (N_30259,N_27064,N_29181);
nor U30260 (N_30260,N_29097,N_27777);
xnor U30261 (N_30261,N_27737,N_26294);
nor U30262 (N_30262,N_27076,N_27668);
or U30263 (N_30263,N_25881,N_25133);
nand U30264 (N_30264,N_27011,N_29426);
or U30265 (N_30265,N_29763,N_25032);
nand U30266 (N_30266,N_29721,N_27157);
or U30267 (N_30267,N_28771,N_25089);
and U30268 (N_30268,N_28830,N_26464);
xor U30269 (N_30269,N_27158,N_26161);
xnor U30270 (N_30270,N_29992,N_25287);
xor U30271 (N_30271,N_27519,N_25395);
and U30272 (N_30272,N_27110,N_25515);
xnor U30273 (N_30273,N_27688,N_27817);
xnor U30274 (N_30274,N_26619,N_28657);
or U30275 (N_30275,N_26665,N_28484);
and U30276 (N_30276,N_28174,N_28620);
nor U30277 (N_30277,N_29815,N_27262);
nand U30278 (N_30278,N_29402,N_25161);
nor U30279 (N_30279,N_28876,N_28846);
and U30280 (N_30280,N_29658,N_28838);
nand U30281 (N_30281,N_29089,N_29878);
nand U30282 (N_30282,N_28975,N_25506);
nor U30283 (N_30283,N_26182,N_27275);
and U30284 (N_30284,N_28383,N_28208);
and U30285 (N_30285,N_25643,N_27172);
and U30286 (N_30286,N_27659,N_29715);
xor U30287 (N_30287,N_29963,N_26783);
nor U30288 (N_30288,N_27724,N_28043);
and U30289 (N_30289,N_25403,N_28014);
or U30290 (N_30290,N_27121,N_27905);
and U30291 (N_30291,N_28184,N_27412);
or U30292 (N_30292,N_26254,N_27257);
xor U30293 (N_30293,N_27510,N_25771);
xor U30294 (N_30294,N_25152,N_25872);
and U30295 (N_30295,N_29995,N_27354);
nor U30296 (N_30296,N_27313,N_26670);
or U30297 (N_30297,N_26105,N_28788);
nor U30298 (N_30298,N_25351,N_26604);
xnor U30299 (N_30299,N_29655,N_25617);
and U30300 (N_30300,N_29244,N_27292);
or U30301 (N_30301,N_29983,N_28803);
and U30302 (N_30302,N_29880,N_27204);
nand U30303 (N_30303,N_27274,N_25138);
or U30304 (N_30304,N_27109,N_27665);
nor U30305 (N_30305,N_27581,N_26557);
nor U30306 (N_30306,N_25524,N_28823);
or U30307 (N_30307,N_25470,N_25268);
nor U30308 (N_30308,N_27855,N_26704);
xnor U30309 (N_30309,N_28834,N_29725);
xnor U30310 (N_30310,N_29569,N_29494);
nor U30311 (N_30311,N_27206,N_28557);
nor U30312 (N_30312,N_29220,N_25868);
xor U30313 (N_30313,N_25815,N_27909);
nand U30314 (N_30314,N_29463,N_26240);
and U30315 (N_30315,N_29556,N_26693);
nor U30316 (N_30316,N_28101,N_28676);
xnor U30317 (N_30317,N_29378,N_26171);
nand U30318 (N_30318,N_26528,N_27049);
or U30319 (N_30319,N_29932,N_26468);
nand U30320 (N_30320,N_28360,N_29075);
nor U30321 (N_30321,N_26869,N_25832);
nor U30322 (N_30322,N_29329,N_27938);
nand U30323 (N_30323,N_26396,N_26688);
or U30324 (N_30324,N_26074,N_29241);
or U30325 (N_30325,N_28583,N_26441);
or U30326 (N_30326,N_26451,N_25838);
and U30327 (N_30327,N_25038,N_29330);
nor U30328 (N_30328,N_28239,N_29873);
nand U30329 (N_30329,N_27755,N_26567);
xor U30330 (N_30330,N_28224,N_27437);
xnor U30331 (N_30331,N_29230,N_29362);
nand U30332 (N_30332,N_26185,N_27900);
or U30333 (N_30333,N_26729,N_29613);
xor U30334 (N_30334,N_27258,N_29607);
and U30335 (N_30335,N_29177,N_26717);
xor U30336 (N_30336,N_29824,N_29841);
and U30337 (N_30337,N_29319,N_25834);
xor U30338 (N_30338,N_25749,N_28336);
nand U30339 (N_30339,N_25673,N_25496);
and U30340 (N_30340,N_25487,N_27331);
nand U30341 (N_30341,N_27291,N_25766);
nor U30342 (N_30342,N_28025,N_28568);
nand U30343 (N_30343,N_28939,N_27409);
nor U30344 (N_30344,N_28040,N_25912);
nor U30345 (N_30345,N_25862,N_25034);
and U30346 (N_30346,N_25548,N_29595);
and U30347 (N_30347,N_29538,N_26205);
or U30348 (N_30348,N_28187,N_26999);
nor U30349 (N_30349,N_26649,N_28369);
xor U30350 (N_30350,N_27949,N_27929);
nand U30351 (N_30351,N_27997,N_28956);
or U30352 (N_30352,N_27864,N_27191);
and U30353 (N_30353,N_27764,N_29803);
and U30354 (N_30354,N_29555,N_28152);
nor U30355 (N_30355,N_27410,N_28382);
nor U30356 (N_30356,N_25885,N_26053);
or U30357 (N_30357,N_27217,N_28633);
and U30358 (N_30358,N_27653,N_26444);
and U30359 (N_30359,N_27805,N_28660);
and U30360 (N_30360,N_26725,N_26224);
xor U30361 (N_30361,N_27641,N_26559);
xor U30362 (N_30362,N_28864,N_29624);
nand U30363 (N_30363,N_28986,N_25029);
or U30364 (N_30364,N_27070,N_26425);
nor U30365 (N_30365,N_28123,N_25902);
and U30366 (N_30366,N_29571,N_29930);
xnor U30367 (N_30367,N_25589,N_27335);
and U30368 (N_30368,N_26945,N_29165);
nor U30369 (N_30369,N_27247,N_26229);
nand U30370 (N_30370,N_25947,N_29265);
nand U30371 (N_30371,N_27446,N_26295);
nor U30372 (N_30372,N_25365,N_29452);
and U30373 (N_30373,N_28154,N_25467);
or U30374 (N_30374,N_26976,N_28284);
nand U30375 (N_30375,N_25367,N_26671);
or U30376 (N_30376,N_28628,N_27447);
xor U30377 (N_30377,N_25579,N_25056);
nand U30378 (N_30378,N_26722,N_28299);
nand U30379 (N_30379,N_25626,N_29923);
nand U30380 (N_30380,N_29419,N_26899);
nor U30381 (N_30381,N_25425,N_25143);
and U30382 (N_30382,N_28760,N_29172);
and U30383 (N_30383,N_26216,N_28310);
or U30384 (N_30384,N_26217,N_25375);
nor U30385 (N_30385,N_26701,N_25896);
nor U30386 (N_30386,N_29907,N_28571);
nor U30387 (N_30387,N_29310,N_26923);
nand U30388 (N_30388,N_27012,N_25972);
and U30389 (N_30389,N_29999,N_29281);
or U30390 (N_30390,N_26546,N_25583);
nor U30391 (N_30391,N_29527,N_29947);
nor U30392 (N_30392,N_25171,N_25334);
and U30393 (N_30393,N_27245,N_29375);
xnor U30394 (N_30394,N_27774,N_28926);
nor U30395 (N_30395,N_26104,N_25691);
nand U30396 (N_30396,N_29057,N_26520);
xnor U30397 (N_30397,N_28562,N_25773);
nand U30398 (N_30398,N_25587,N_26233);
nor U30399 (N_30399,N_27642,N_29698);
and U30400 (N_30400,N_26756,N_26437);
and U30401 (N_30401,N_25723,N_27279);
nand U30402 (N_30402,N_26998,N_27861);
and U30403 (N_30403,N_27571,N_29360);
nand U30404 (N_30404,N_27925,N_27567);
xnor U30405 (N_30405,N_28552,N_28155);
nor U30406 (N_30406,N_25554,N_29117);
and U30407 (N_30407,N_28326,N_27117);
nor U30408 (N_30408,N_28249,N_27229);
nand U30409 (N_30409,N_25221,N_25033);
nor U30410 (N_30410,N_25124,N_27707);
nor U30411 (N_30411,N_28783,N_27492);
xnor U30412 (N_30412,N_27159,N_26303);
xor U30413 (N_30413,N_25389,N_25167);
nor U30414 (N_30414,N_29998,N_25995);
xnor U30415 (N_30415,N_27355,N_26458);
and U30416 (N_30416,N_27429,N_29127);
or U30417 (N_30417,N_26948,N_25776);
and U30418 (N_30418,N_29570,N_26636);
nand U30419 (N_30419,N_25464,N_26347);
xor U30420 (N_30420,N_29386,N_28363);
xor U30421 (N_30421,N_28377,N_25319);
and U30422 (N_30422,N_29167,N_26789);
or U30423 (N_30423,N_25588,N_28083);
or U30424 (N_30424,N_29389,N_28543);
and U30425 (N_30425,N_29288,N_27319);
xnor U30426 (N_30426,N_25843,N_29380);
or U30427 (N_30427,N_28269,N_26718);
and U30428 (N_30428,N_26777,N_29313);
and U30429 (N_30429,N_28798,N_29816);
nand U30430 (N_30430,N_29994,N_26614);
and U30431 (N_30431,N_28828,N_29597);
and U30432 (N_30432,N_27990,N_27549);
xnor U30433 (N_30433,N_29029,N_27405);
or U30434 (N_30434,N_25608,N_28847);
nand U30435 (N_30435,N_25424,N_29843);
nor U30436 (N_30436,N_28226,N_28036);
xor U30437 (N_30437,N_29657,N_25141);
nand U30438 (N_30438,N_25883,N_25865);
or U30439 (N_30439,N_28613,N_29321);
and U30440 (N_30440,N_25945,N_29576);
xnor U30441 (N_30441,N_25223,N_25666);
xor U30442 (N_30442,N_27303,N_27538);
xnor U30443 (N_30443,N_28577,N_27886);
and U30444 (N_30444,N_26949,N_25706);
xor U30445 (N_30445,N_27666,N_25069);
or U30446 (N_30446,N_27311,N_27720);
nand U30447 (N_30447,N_29013,N_28278);
nor U30448 (N_30448,N_29905,N_26550);
nor U30449 (N_30449,N_25561,N_26969);
nand U30450 (N_30450,N_26648,N_28460);
xor U30451 (N_30451,N_29525,N_27866);
nand U30452 (N_30452,N_27403,N_28728);
xor U30453 (N_30453,N_27381,N_26656);
and U30454 (N_30454,N_25407,N_28058);
or U30455 (N_30455,N_27052,N_26518);
or U30456 (N_30456,N_27149,N_29587);
nor U30457 (N_30457,N_26511,N_28679);
nor U30458 (N_30458,N_29333,N_28959);
xnor U30459 (N_30459,N_29610,N_26120);
xor U30460 (N_30460,N_29544,N_26960);
xor U30461 (N_30461,N_26145,N_26612);
nand U30462 (N_30462,N_27890,N_28104);
xor U30463 (N_30463,N_26106,N_26101);
nor U30464 (N_30464,N_27035,N_29677);
nand U30465 (N_30465,N_26011,N_28439);
or U30466 (N_30466,N_26381,N_25120);
or U30467 (N_30467,N_27754,N_29801);
or U30468 (N_30468,N_28396,N_25363);
or U30469 (N_30469,N_29140,N_27238);
xnor U30470 (N_30470,N_26525,N_29183);
xnor U30471 (N_30471,N_26764,N_29559);
and U30472 (N_30472,N_26913,N_27225);
or U30473 (N_30473,N_29482,N_28037);
nand U30474 (N_30474,N_26069,N_26855);
or U30475 (N_30475,N_27306,N_28766);
and U30476 (N_30476,N_28235,N_26689);
nor U30477 (N_30477,N_25641,N_25473);
nor U30478 (N_30478,N_25298,N_29124);
and U30479 (N_30479,N_29888,N_25466);
nand U30480 (N_30480,N_29155,N_26873);
nand U30481 (N_30481,N_25505,N_26060);
or U30482 (N_30482,N_26784,N_29552);
xor U30483 (N_30483,N_26079,N_27414);
and U30484 (N_30484,N_27456,N_26005);
nor U30485 (N_30485,N_25784,N_26027);
nand U30486 (N_30486,N_28913,N_28066);
or U30487 (N_30487,N_29173,N_26699);
nand U30488 (N_30488,N_29295,N_27502);
and U30489 (N_30489,N_25647,N_29564);
or U30490 (N_30490,N_29722,N_25938);
nand U30491 (N_30491,N_26147,N_28687);
xnor U30492 (N_30492,N_27819,N_25211);
and U30493 (N_30493,N_27550,N_25176);
nand U30494 (N_30494,N_25886,N_27803);
nand U30495 (N_30495,N_29400,N_27431);
xnor U30496 (N_30496,N_28988,N_26677);
nor U30497 (N_30497,N_29616,N_26685);
nand U30498 (N_30498,N_27256,N_27108);
nand U30499 (N_30499,N_27349,N_28328);
or U30500 (N_30500,N_26055,N_26795);
nor U30501 (N_30501,N_29954,N_27499);
nand U30502 (N_30502,N_26523,N_29536);
and U30503 (N_30503,N_28219,N_28202);
nor U30504 (N_30504,N_29245,N_26212);
xor U30505 (N_30505,N_29032,N_26893);
xnor U30506 (N_30506,N_28453,N_25183);
or U30507 (N_30507,N_28455,N_28160);
and U30508 (N_30508,N_28228,N_25882);
and U30509 (N_30509,N_26095,N_28475);
nand U30510 (N_30510,N_25530,N_26702);
or U30511 (N_30511,N_25154,N_25009);
and U30512 (N_30512,N_26344,N_27254);
and U30513 (N_30513,N_27673,N_25053);
xor U30514 (N_30514,N_26463,N_25970);
nand U30515 (N_30515,N_29524,N_28692);
and U30516 (N_30516,N_29781,N_25193);
and U30517 (N_30517,N_26087,N_28797);
nand U30518 (N_30518,N_28522,N_28248);
nor U30519 (N_30519,N_25679,N_25708);
or U30520 (N_30520,N_28331,N_28404);
nand U30521 (N_30521,N_27421,N_26987);
and U30522 (N_30522,N_28023,N_27366);
or U30523 (N_30523,N_27369,N_25480);
and U30524 (N_30524,N_27263,N_29535);
or U30525 (N_30525,N_28600,N_27318);
nand U30526 (N_30526,N_26419,N_27271);
and U30527 (N_30527,N_26521,N_27170);
and U30528 (N_30528,N_25603,N_27185);
nand U30529 (N_30529,N_27242,N_26056);
nor U30530 (N_30530,N_27716,N_29844);
nand U30531 (N_30531,N_25169,N_29911);
nor U30532 (N_30532,N_29738,N_26438);
nand U30533 (N_30533,N_28912,N_28558);
nor U30534 (N_30534,N_27651,N_29809);
or U30535 (N_30535,N_26421,N_25220);
and U30536 (N_30536,N_29833,N_28880);
and U30537 (N_30537,N_27594,N_26131);
nor U30538 (N_30538,N_26172,N_29692);
nor U30539 (N_30539,N_25194,N_28486);
nor U30540 (N_30540,N_28005,N_27481);
xor U30541 (N_30541,N_27545,N_26631);
or U30542 (N_30542,N_26686,N_27357);
xor U30543 (N_30543,N_28792,N_26916);
nor U30544 (N_30544,N_25050,N_25135);
and U30545 (N_30545,N_26340,N_27609);
or U30546 (N_30546,N_29012,N_26622);
or U30547 (N_30547,N_26621,N_27582);
nand U30548 (N_30548,N_28063,N_28277);
or U30549 (N_30549,N_29184,N_26496);
or U30550 (N_30550,N_25669,N_29484);
xor U30551 (N_30551,N_28452,N_26097);
nand U30552 (N_30552,N_29122,N_26028);
nand U30553 (N_30553,N_28497,N_25260);
nand U30554 (N_30554,N_26498,N_26561);
xor U30555 (N_30555,N_27034,N_28379);
or U30556 (N_30556,N_27887,N_27865);
or U30557 (N_30557,N_29625,N_26012);
and U30558 (N_30558,N_25750,N_26386);
nand U30559 (N_30559,N_27039,N_26020);
xor U30560 (N_30560,N_27989,N_25160);
and U30561 (N_30561,N_28627,N_27486);
nor U30562 (N_30562,N_28015,N_25863);
nor U30563 (N_30563,N_29125,N_26607);
nand U30564 (N_30564,N_25768,N_28361);
or U30565 (N_30565,N_27682,N_25404);
xnor U30566 (N_30566,N_25087,N_29631);
or U30567 (N_30567,N_25036,N_27506);
nor U30568 (N_30568,N_27517,N_26098);
xor U30569 (N_30569,N_28727,N_28231);
or U30570 (N_30570,N_29035,N_29204);
xor U30571 (N_30571,N_25237,N_26816);
and U30572 (N_30572,N_28672,N_25388);
xnor U30573 (N_30573,N_28033,N_28917);
and U30574 (N_30574,N_29233,N_27243);
xor U30575 (N_30575,N_29810,N_28819);
xnor U30576 (N_30576,N_29812,N_27061);
or U30577 (N_30577,N_25752,N_25637);
or U30578 (N_30578,N_28984,N_28499);
nand U30579 (N_30579,N_29424,N_28156);
xor U30580 (N_30580,N_26346,N_25571);
nand U30581 (N_30581,N_27736,N_29428);
nor U30582 (N_30582,N_28252,N_25905);
or U30583 (N_30583,N_26361,N_28724);
nand U30584 (N_30584,N_29495,N_28943);
and U30585 (N_30585,N_25381,N_27345);
xor U30586 (N_30586,N_29696,N_27543);
and U30587 (N_30587,N_29795,N_28292);
nor U30588 (N_30588,N_25967,N_27082);
nand U30589 (N_30589,N_29519,N_29621);
and U30590 (N_30590,N_25783,N_27163);
xnor U30591 (N_30591,N_28517,N_26424);
or U30592 (N_30592,N_25332,N_29411);
nor U30593 (N_30593,N_26928,N_26483);
nor U30594 (N_30594,N_26910,N_29753);
or U30595 (N_30595,N_25421,N_26318);
or U30596 (N_30596,N_29584,N_25485);
xor U30597 (N_30597,N_27558,N_26968);
nand U30598 (N_30598,N_29429,N_29394);
nor U30599 (N_30599,N_29308,N_29351);
nor U30600 (N_30600,N_26179,N_28468);
and U30601 (N_30601,N_29193,N_25188);
xor U30602 (N_30602,N_27951,N_27112);
nand U30603 (N_30603,N_27536,N_25063);
xnor U30604 (N_30604,N_28438,N_27181);
and U30605 (N_30605,N_26711,N_26057);
xor U30606 (N_30606,N_26651,N_29077);
nand U30607 (N_30607,N_29877,N_27378);
nand U30608 (N_30608,N_26574,N_26174);
and U30609 (N_30609,N_29079,N_29931);
and U30610 (N_30610,N_29132,N_26533);
or U30611 (N_30611,N_29414,N_27868);
and U30612 (N_30612,N_28738,N_28902);
nand U30613 (N_30613,N_27521,N_26929);
or U30614 (N_30614,N_26932,N_28067);
or U30615 (N_30615,N_29979,N_29415);
nand U30616 (N_30616,N_27348,N_28177);
and U30617 (N_30617,N_26431,N_26871);
or U30618 (N_30618,N_25932,N_25787);
xnor U30619 (N_30619,N_26971,N_26637);
xor U30620 (N_30620,N_28954,N_29670);
xnor U30621 (N_30621,N_29853,N_28294);
nand U30622 (N_30622,N_26306,N_29212);
nor U30623 (N_30623,N_29920,N_25944);
or U30624 (N_30624,N_29160,N_28450);
or U30625 (N_30625,N_29705,N_26673);
xor U30626 (N_30626,N_26411,N_29693);
nor U30627 (N_30627,N_29290,N_29372);
nand U30628 (N_30628,N_25820,N_26796);
and U30629 (N_30629,N_28012,N_25410);
xnor U30630 (N_30630,N_25181,N_29434);
nand U30631 (N_30631,N_29418,N_27051);
or U30632 (N_30632,N_29750,N_28075);
xnor U30633 (N_30633,N_28780,N_28594);
nor U30634 (N_30634,N_28860,N_28826);
xor U30635 (N_30635,N_25270,N_25642);
nor U30636 (N_30636,N_29326,N_27177);
or U30637 (N_30637,N_27676,N_28705);
or U30638 (N_30638,N_28443,N_28282);
xor U30639 (N_30639,N_29959,N_26917);
xnor U30640 (N_30640,N_27654,N_26886);
nor U30641 (N_30641,N_29094,N_26178);
nand U30642 (N_30642,N_25468,N_28746);
nand U30643 (N_30643,N_25074,N_29819);
or U30644 (N_30644,N_26825,N_25428);
xnor U30645 (N_30645,N_29095,N_27950);
nor U30646 (N_30646,N_25699,N_28132);
nand U30647 (N_30647,N_27782,N_27600);
or U30648 (N_30648,N_28211,N_25736);
or U30649 (N_30649,N_25527,N_27717);
or U30650 (N_30650,N_28733,N_25928);
xnor U30651 (N_30651,N_28907,N_25338);
or U30652 (N_30652,N_28634,N_29573);
nor U30653 (N_30653,N_25083,N_29608);
and U30654 (N_30654,N_27607,N_26149);
or U30655 (N_30655,N_25172,N_26125);
nor U30656 (N_30656,N_26885,N_28233);
nor U30657 (N_30657,N_28042,N_29708);
nor U30658 (N_30658,N_25442,N_28283);
or U30659 (N_30659,N_29471,N_26470);
or U30660 (N_30660,N_26678,N_27228);
and U30661 (N_30661,N_26204,N_28490);
nor U30662 (N_30662,N_26489,N_25672);
xnor U30663 (N_30663,N_27891,N_29135);
and U30664 (N_30664,N_28942,N_25180);
and U30665 (N_30665,N_25025,N_27548);
xnor U30666 (N_30666,N_29465,N_29522);
xnor U30667 (N_30667,N_25317,N_25292);
or U30668 (N_30668,N_26526,N_29618);
xnor U30669 (N_30669,N_27411,N_29078);
xor U30670 (N_30670,N_27552,N_29865);
xnor U30671 (N_30671,N_28393,N_28532);
and U30672 (N_30672,N_26151,N_26395);
or U30673 (N_30673,N_27327,N_28719);
xor U30674 (N_30674,N_29820,N_25566);
or U30675 (N_30675,N_28559,N_27352);
or U30676 (N_30676,N_29283,N_27882);
or U30677 (N_30677,N_26359,N_28997);
and U30678 (N_30678,N_28428,N_29449);
and U30679 (N_30679,N_27179,N_29455);
nor U30680 (N_30680,N_26369,N_29240);
nor U30681 (N_30681,N_25937,N_27050);
xnor U30682 (N_30682,N_29746,N_28615);
and U30683 (N_30683,N_29917,N_25609);
xnor U30684 (N_30684,N_26049,N_29206);
nand U30685 (N_30685,N_25357,N_29325);
nor U30686 (N_30686,N_27508,N_26168);
and U30687 (N_30687,N_27813,N_28590);
and U30688 (N_30688,N_25528,N_26491);
and U30689 (N_30689,N_29390,N_26117);
and U30690 (N_30690,N_25127,N_27712);
nand U30691 (N_30691,N_28047,N_28261);
nand U30692 (N_30692,N_25611,N_27309);
nand U30693 (N_30693,N_26530,N_29687);
xnor U30694 (N_30694,N_25722,N_26635);
or U30695 (N_30695,N_28905,N_25624);
and U30696 (N_30696,N_28347,N_29847);
and U30697 (N_30697,N_26310,N_26457);
nor U30698 (N_30698,N_29989,N_28653);
nor U30699 (N_30699,N_27343,N_27912);
and U30700 (N_30700,N_27487,N_29236);
nand U30701 (N_30701,N_28300,N_29457);
nand U30702 (N_30702,N_26460,N_26114);
xnor U30703 (N_30703,N_26195,N_25818);
nand U30704 (N_30704,N_27462,N_27340);
nor U30705 (N_30705,N_28915,N_26223);
nor U30706 (N_30706,N_25567,N_27359);
nor U30707 (N_30707,N_25380,N_26287);
xor U30708 (N_30708,N_27841,N_29063);
nor U30709 (N_30709,N_27015,N_27124);
nor U30710 (N_30710,N_25599,N_28567);
xor U30711 (N_30711,N_29370,N_27649);
and U30712 (N_30712,N_25422,N_28632);
or U30713 (N_30713,N_28784,N_25014);
nand U30714 (N_30714,N_26754,N_29256);
and U30715 (N_30715,N_26128,N_27305);
nor U30716 (N_30716,N_28135,N_26751);
or U30717 (N_30717,N_25654,N_28879);
and U30718 (N_30718,N_29580,N_29838);
xnor U30719 (N_30719,N_26354,N_29557);
nor U30720 (N_30720,N_28643,N_29825);
nor U30721 (N_30721,N_28109,N_29439);
xor U30722 (N_30722,N_29623,N_28011);
xnor U30723 (N_30723,N_26547,N_25569);
xnor U30724 (N_30724,N_25356,N_28340);
or U30725 (N_30725,N_28533,N_29501);
nor U30726 (N_30726,N_25978,N_25811);
and U30727 (N_30727,N_25894,N_26277);
nand U30728 (N_30728,N_26293,N_25289);
nor U30729 (N_30729,N_25376,N_27048);
or U30730 (N_30730,N_29651,N_27060);
nor U30731 (N_30731,N_25760,N_25954);
nand U30732 (N_30732,N_27086,N_26782);
or U30733 (N_30733,N_28895,N_27939);
and U30734 (N_30734,N_25688,N_26093);
nor U30735 (N_30735,N_25775,N_26582);
nand U30736 (N_30736,N_26786,N_27572);
nor U30737 (N_30737,N_28362,N_25806);
or U30738 (N_30738,N_27874,N_25294);
xnor U30739 (N_30739,N_26332,N_25210);
and U30740 (N_30740,N_29409,N_26867);
and U30741 (N_30741,N_28425,N_29451);
xnor U30742 (N_30742,N_27959,N_28608);
nand U30743 (N_30743,N_29076,N_27913);
xnor U30744 (N_30744,N_27760,N_27252);
and U30745 (N_30745,N_28832,N_26112);
nand U30746 (N_30746,N_29935,N_29247);
xor U30747 (N_30747,N_29589,N_25131);
and U30748 (N_30748,N_28121,N_27092);
or U30749 (N_30749,N_28491,N_29656);
and U30750 (N_30750,N_27827,N_28021);
nor U30751 (N_30751,N_28133,N_26586);
xnor U30752 (N_30752,N_26445,N_25108);
nor U30753 (N_30753,N_26645,N_29171);
and U30754 (N_30754,N_27236,N_28502);
nor U30755 (N_30755,N_29141,N_26363);
or U30756 (N_30756,N_29363,N_27324);
nor U30757 (N_30757,N_26023,N_29084);
nor U30758 (N_30758,N_27965,N_29470);
nand U30759 (N_30759,N_28685,N_29365);
nand U30760 (N_30760,N_29786,N_26962);
and U30761 (N_30761,N_25648,N_25700);
and U30762 (N_30762,N_26297,N_25917);
or U30763 (N_30763,N_29837,N_29275);
or U30764 (N_30764,N_29440,N_25799);
xnor U30765 (N_30765,N_29203,N_26281);
xor U30766 (N_30766,N_29546,N_27580);
and U30767 (N_30767,N_25324,N_27526);
nand U30768 (N_30768,N_28175,N_28868);
or U30769 (N_30769,N_26734,N_26345);
xnor U30770 (N_30770,N_25073,N_27430);
nand U30771 (N_30771,N_26156,N_27629);
nor U30772 (N_30772,N_26905,N_26562);
nor U30773 (N_30773,N_29373,N_25352);
nor U30774 (N_30774,N_26502,N_25372);
nor U30775 (N_30775,N_29282,N_28076);
and U30776 (N_30776,N_28896,N_28086);
or U30777 (N_30777,N_25204,N_27146);
xnor U30778 (N_30778,N_26512,N_29793);
and U30779 (N_30779,N_29249,N_28016);
or U30780 (N_30780,N_25714,N_28316);
xnor U30781 (N_30781,N_29427,N_25904);
xnor U30782 (N_30782,N_27053,N_25387);
nor U30783 (N_30783,N_26990,N_25413);
or U30784 (N_30784,N_25481,N_26835);
or U30785 (N_30785,N_26357,N_28843);
xnor U30786 (N_30786,N_28658,N_29016);
xor U30787 (N_30787,N_28815,N_26193);
and U30788 (N_30788,N_25693,N_25364);
nand U30789 (N_30789,N_26875,N_28273);
and U30790 (N_30790,N_25213,N_27105);
and U30791 (N_30791,N_25989,N_26746);
xor U30792 (N_30792,N_29606,N_27516);
nand U30793 (N_30793,N_29120,N_29446);
xnor U30794 (N_30794,N_28467,N_25158);
xnor U30795 (N_30795,N_27209,N_25844);
xor U30796 (N_30796,N_26166,N_25725);
and U30797 (N_30797,N_28965,N_25501);
or U30798 (N_30798,N_26793,N_29396);
nor U30799 (N_30799,N_26261,N_25956);
xnor U30800 (N_30800,N_28243,N_28752);
or U30801 (N_30801,N_29111,N_28509);
nand U30802 (N_30802,N_28540,N_27505);
xnor U30803 (N_30803,N_27541,N_25246);
or U30804 (N_30804,N_25851,N_28624);
nor U30805 (N_30805,N_25719,N_25225);
nor U30806 (N_30806,N_28334,N_29950);
and U30807 (N_30807,N_29893,N_27603);
xor U30808 (N_30808,N_27626,N_25288);
nand U30809 (N_30809,N_27356,N_25539);
nand U30810 (N_30810,N_28971,N_29898);
or U30811 (N_30811,N_28168,N_26107);
xnor U30812 (N_30812,N_28527,N_25071);
nor U30813 (N_30813,N_27083,N_27285);
xnor U30814 (N_30814,N_28789,N_27166);
or U30815 (N_30815,N_26897,N_29770);
xor U30816 (N_30816,N_29272,N_27843);
xor U30817 (N_30817,N_28863,N_29867);
nor U30818 (N_30818,N_26507,N_25010);
nor U30819 (N_30819,N_29291,N_26597);
xnor U30820 (N_30820,N_25846,N_29500);
xnor U30821 (N_30821,N_25829,N_29188);
and U30822 (N_30822,N_29784,N_28617);
xnor U30823 (N_30823,N_28476,N_28857);
nor U30824 (N_30824,N_25476,N_29279);
or U30825 (N_30825,N_27759,N_27878);
and U30826 (N_30826,N_27731,N_29904);
nand U30827 (N_30827,N_26045,N_29253);
and U30828 (N_30828,N_27844,N_29936);
nand U30829 (N_30829,N_26861,N_29179);
and U30830 (N_30830,N_25711,N_26943);
and U30831 (N_30831,N_26694,N_28867);
nor U30832 (N_30832,N_27907,N_29694);
and U30833 (N_30833,N_25157,N_25507);
or U30834 (N_30834,N_25296,N_25490);
nand U30835 (N_30835,N_26080,N_27856);
nor U30836 (N_30836,N_26247,N_27454);
nand U30837 (N_30837,N_29910,N_25003);
xnor U30838 (N_30838,N_28950,N_29105);
nor U30839 (N_30839,N_25875,N_27286);
nand U30840 (N_30840,N_29025,N_26488);
xor U30841 (N_30841,N_26977,N_25119);
xor U30842 (N_30842,N_28466,N_27165);
nor U30843 (N_30843,N_27260,N_29860);
nand U30844 (N_30844,N_25030,N_25282);
xor U30845 (N_30845,N_25874,N_29971);
and U30846 (N_30846,N_25860,N_28113);
nor U30847 (N_30847,N_26829,N_28159);
nor U30848 (N_30848,N_27638,N_27758);
nor U30849 (N_30849,N_27144,N_29195);
nor U30850 (N_30850,N_25839,N_25024);
nor U30851 (N_30851,N_29399,N_29159);
xor U30852 (N_30852,N_27169,N_29811);
and U30853 (N_30853,N_27030,N_25990);
and U30854 (N_30854,N_25048,N_26406);
xnor U30855 (N_30855,N_27393,N_25392);
or U30856 (N_30856,N_27879,N_28463);
xor U30857 (N_30857,N_27529,N_28805);
nor U30858 (N_30858,N_29565,N_29190);
or U30859 (N_30859,N_28892,N_26416);
nor U30860 (N_30860,N_29176,N_25051);
or U30861 (N_30861,N_26581,N_26926);
and U30862 (N_30862,N_28859,N_26330);
xor U30863 (N_30863,N_27219,N_26429);
or U30864 (N_30864,N_28835,N_27244);
nor U30865 (N_30865,N_27636,N_27130);
and U30866 (N_30866,N_26220,N_27198);
nor U30867 (N_30867,N_26311,N_28973);
and U30868 (N_30868,N_26534,N_28542);
nand U30869 (N_30869,N_26992,N_29643);
nand U30870 (N_30870,N_26994,N_26129);
or U30871 (N_30871,N_28970,N_29970);
nand U30872 (N_30872,N_28329,N_26935);
nand U30873 (N_30873,N_29785,N_28038);
nand U30874 (N_30874,N_28656,N_25068);
or U30875 (N_30875,N_28720,N_28032);
or U30876 (N_30876,N_25663,N_25819);
nor U30877 (N_30877,N_28220,N_27952);
and U30878 (N_30878,N_27391,N_28344);
xnor U30879 (N_30879,N_26788,N_27889);
and U30880 (N_30880,N_25628,N_27148);
nand U30881 (N_30881,N_29129,N_25920);
xor U30882 (N_30882,N_26333,N_25992);
nor U30883 (N_30883,N_28726,N_25757);
nand U30884 (N_30884,N_25216,N_29136);
nor U30885 (N_30885,N_25632,N_29848);
nand U30886 (N_30886,N_26162,N_25888);
nor U30887 (N_30887,N_26780,N_27401);
xnor U30888 (N_30888,N_28578,N_28141);
and U30889 (N_30889,N_25961,N_29509);
nand U30890 (N_30890,N_26382,N_29648);
nor U30891 (N_30891,N_26133,N_28003);
xor U30892 (N_30892,N_25958,N_29780);
and U30893 (N_30893,N_25867,N_26951);
xnor U30894 (N_30894,N_25993,N_27389);
nand U30895 (N_30895,N_27438,N_27687);
or U30896 (N_30896,N_25615,N_25411);
and U30897 (N_30897,N_28730,N_25659);
xnor U30898 (N_30898,N_27358,N_28045);
xor U30899 (N_30899,N_28759,N_29130);
or U30900 (N_30900,N_29940,N_26032);
xor U30901 (N_30901,N_28576,N_27809);
or U30902 (N_30902,N_29515,N_26736);
and U30903 (N_30903,N_25415,N_28647);
and U30904 (N_30904,N_26652,N_26213);
nand U30905 (N_30905,N_27847,N_27273);
nor U30906 (N_30906,N_27880,N_25765);
xor U30907 (N_30907,N_29644,N_26040);
or U30908 (N_30908,N_25730,N_26379);
nand U30909 (N_30909,N_28709,N_27232);
nand U30910 (N_30910,N_28749,N_28775);
and U30911 (N_30911,N_28079,N_26246);
xor U30912 (N_30912,N_27362,N_25924);
or U30913 (N_30913,N_27968,N_25235);
xnor U30914 (N_30914,N_27337,N_25075);
xor U30915 (N_30915,N_29251,N_27867);
and U30916 (N_30916,N_26997,N_27851);
or U30917 (N_30917,N_25705,N_25361);
xnor U30918 (N_30918,N_25293,N_29517);
or U30919 (N_30919,N_28419,N_29196);
and U30920 (N_30920,N_28919,N_29661);
xnor U30921 (N_30921,N_28873,N_28189);
nor U30922 (N_30922,N_26984,N_26707);
nand U30923 (N_30923,N_29614,N_27531);
or U30924 (N_30924,N_27014,N_28920);
nand U30925 (N_30925,N_28345,N_25233);
nand U30926 (N_30926,N_25513,N_28645);
nand U30927 (N_30927,N_29232,N_25694);
or U30928 (N_30928,N_27178,N_25596);
nand U30929 (N_30929,N_29919,N_25553);
nor U30930 (N_30930,N_27767,N_26096);
and U30931 (N_30931,N_26907,N_29270);
and U30932 (N_30932,N_25146,N_29435);
nor U30933 (N_30933,N_27497,N_25308);
or U30934 (N_30934,N_28126,N_28210);
nor U30935 (N_30935,N_29857,N_29083);
or U30936 (N_30936,N_27186,N_26221);
nand U30937 (N_30937,N_29590,N_25103);
and U30938 (N_30938,N_27849,N_28769);
or U30939 (N_30939,N_29227,N_28397);
and U30940 (N_30940,N_28199,N_26716);
or U30941 (N_30941,N_29082,N_26135);
nor U30942 (N_30942,N_27601,N_28114);
nor U30943 (N_30943,N_29085,N_28511);
or U30944 (N_30944,N_28507,N_28569);
xnor U30945 (N_30945,N_25923,N_26891);
xor U30946 (N_30946,N_26071,N_26724);
or U30947 (N_30947,N_27160,N_27029);
xnor U30948 (N_30948,N_26571,N_25504);
nor U30949 (N_30949,N_27476,N_27814);
nand U30950 (N_30950,N_26791,N_27415);
xnor U30951 (N_30951,N_26772,N_27727);
or U30952 (N_30952,N_25745,N_27046);
nand U30953 (N_30953,N_25646,N_26856);
nand U30954 (N_30954,N_25942,N_28346);
nand U30955 (N_30955,N_29531,N_25519);
xor U30956 (N_30956,N_25453,N_29391);
nor U30957 (N_30957,N_28978,N_26335);
xor U30958 (N_30958,N_26770,N_28185);
nor U30959 (N_30959,N_28448,N_29480);
or U30960 (N_30960,N_27719,N_26593);
nor U30961 (N_30961,N_29487,N_28105);
and U30962 (N_30962,N_26538,N_25452);
or U30963 (N_30963,N_27557,N_28858);
nand U30964 (N_30964,N_28667,N_28215);
nor U30965 (N_30965,N_25408,N_28304);
nand U30966 (N_30966,N_26181,N_27205);
nor U30967 (N_30967,N_29379,N_26148);
nor U30968 (N_30968,N_29635,N_25077);
nor U30969 (N_30969,N_28465,N_28564);
xnor U30970 (N_30970,N_28579,N_27570);
nor U30971 (N_30971,N_29802,N_26048);
nand U30972 (N_30972,N_25948,N_26903);
xor U30973 (N_30973,N_25159,N_25795);
or U30974 (N_30974,N_29913,N_29831);
nor U30975 (N_30975,N_25436,N_25281);
and U30976 (N_30976,N_26609,N_25348);
and U30977 (N_30977,N_25716,N_28247);
xnor U30978 (N_30978,N_29060,N_27416);
and U30979 (N_30979,N_26446,N_25532);
or U30980 (N_30980,N_25737,N_27711);
and U30981 (N_30981,N_29977,N_28861);
xnor U30982 (N_30982,N_26368,N_25122);
or U30983 (N_30983,N_28883,N_25987);
nand U30984 (N_30984,N_28444,N_29065);
nand U30985 (N_30985,N_28173,N_26238);
or U30986 (N_30986,N_29080,N_27002);
xor U30987 (N_30987,N_28410,N_27078);
and U30988 (N_30988,N_27518,N_29566);
nand U30989 (N_30989,N_26465,N_25521);
xnor U30990 (N_30990,N_28513,N_29855);
nor U30991 (N_30991,N_27677,N_29318);
xnor U30992 (N_30992,N_27940,N_25707);
xor U30993 (N_30993,N_25342,N_28898);
or U30994 (N_30994,N_25081,N_27089);
nor U30995 (N_30995,N_27972,N_27267);
nor U30996 (N_30996,N_29346,N_26301);
and U30997 (N_30997,N_28431,N_27351);
xor U30998 (N_30998,N_26315,N_25207);
xor U30999 (N_30999,N_25409,N_26611);
or U31000 (N_31000,N_27120,N_26050);
or U31001 (N_31001,N_27452,N_25011);
and U31002 (N_31002,N_25994,N_27474);
nand U31003 (N_31003,N_25262,N_26397);
nand U31004 (N_31004,N_26766,N_28069);
nand U31005 (N_31005,N_25639,N_29133);
xnor U31006 (N_31006,N_28699,N_29962);
xnor U31007 (N_31007,N_27739,N_28207);
or U31008 (N_31008,N_27098,N_29344);
xnor U31009 (N_31009,N_27284,N_25635);
nor U31010 (N_31010,N_28603,N_25586);
nand U31011 (N_31011,N_25988,N_28652);
xor U31012 (N_31012,N_29783,N_26863);
xnor U31013 (N_31013,N_29201,N_25498);
and U31014 (N_31014,N_28518,N_25739);
nand U31015 (N_31015,N_28354,N_26226);
nand U31016 (N_31016,N_27922,N_26009);
or U31017 (N_31017,N_27000,N_26747);
or U31018 (N_31018,N_26450,N_29483);
xor U31019 (N_31019,N_26755,N_29438);
or U31020 (N_31020,N_27791,N_25337);
xor U31021 (N_31021,N_28494,N_25941);
nand U31022 (N_31022,N_26206,N_27801);
and U31023 (N_31023,N_29561,N_26895);
nor U31024 (N_31024,N_28234,N_27898);
and U31025 (N_31025,N_28162,N_28909);
or U31026 (N_31026,N_28225,N_29928);
and U31027 (N_31027,N_29973,N_29118);
nand U31028 (N_31028,N_26768,N_25533);
and U31029 (N_31029,N_27979,N_27031);
or U31030 (N_31030,N_28848,N_29453);
and U31031 (N_31031,N_29381,N_28696);
xnor U31032 (N_31032,N_27776,N_26426);
nand U31033 (N_31033,N_29475,N_25879);
and U31034 (N_31034,N_27745,N_28312);
and U31035 (N_31035,N_26362,N_25004);
and U31036 (N_31036,N_28977,N_28493);
and U31037 (N_31037,N_26100,N_29353);
nand U31038 (N_31038,N_28581,N_25558);
and U31039 (N_31039,N_28240,N_25540);
and U31040 (N_31040,N_27382,N_28257);
nand U31041 (N_31041,N_28521,N_27514);
nand U31042 (N_31042,N_27115,N_28218);
or U31043 (N_31043,N_26922,N_28244);
nor U31044 (N_31044,N_25946,N_26598);
or U31045 (N_31045,N_29139,N_25852);
nor U31046 (N_31046,N_29724,N_27634);
nand U31047 (N_31047,N_25326,N_27080);
xor U31048 (N_31048,N_25478,N_27383);
and U31049 (N_31049,N_27314,N_25713);
and U31050 (N_31050,N_26225,N_26207);
or U31051 (N_31051,N_28548,N_27368);
xnor U31052 (N_31052,N_27290,N_25559);
xor U31053 (N_31053,N_25683,N_25132);
nand U31054 (N_31054,N_27069,N_25283);
xnor U31055 (N_31055,N_25926,N_27652);
nor U31056 (N_31056,N_26235,N_26486);
and U31057 (N_31057,N_27625,N_29432);
xnor U31058 (N_31058,N_29529,N_28831);
xnor U31059 (N_31059,N_27613,N_27265);
or U31060 (N_31060,N_29410,N_26953);
and U31061 (N_31061,N_26579,N_28107);
or U31062 (N_31062,N_28665,N_27099);
or U31063 (N_31063,N_28712,N_26304);
nor U31064 (N_31064,N_27934,N_29757);
or U31065 (N_31065,N_26200,N_27595);
xnor U31066 (N_31066,N_26163,N_27701);
and U31067 (N_31067,N_25525,N_28584);
xnor U31068 (N_31068,N_26506,N_28206);
or U31069 (N_31069,N_26578,N_28001);
xnor U31070 (N_31070,N_26471,N_25975);
or U31071 (N_31071,N_28143,N_27210);
and U31072 (N_31072,N_29485,N_25998);
xnor U31073 (N_31073,N_26309,N_28356);
and U31074 (N_31074,N_29166,N_28471);
xnor U31075 (N_31075,N_28302,N_28417);
xnor U31076 (N_31076,N_29547,N_26710);
xnor U31077 (N_31077,N_27293,N_25692);
xnor U31078 (N_31078,N_28387,N_28203);
nor U31079 (N_31079,N_26284,N_28602);
or U31080 (N_31080,N_27576,N_25512);
and U31081 (N_31081,N_27928,N_29869);
and U31082 (N_31082,N_27010,N_28948);
nand U31083 (N_31083,N_25377,N_27943);
or U31084 (N_31084,N_29539,N_27367);
nor U31085 (N_31085,N_25362,N_25823);
nor U31086 (N_31086,N_28524,N_26908);
or U31087 (N_31087,N_25208,N_25316);
and U31088 (N_31088,N_26537,N_27118);
or U31089 (N_31089,N_29974,N_29051);
and U31090 (N_31090,N_26700,N_26549);
or U31091 (N_31091,N_27224,N_25323);
nor U31092 (N_31092,N_27655,N_27141);
xnor U31093 (N_31093,N_27407,N_28851);
nor U31094 (N_31094,N_29123,N_28555);
xor U31095 (N_31095,N_26192,N_26167);
nand U31096 (N_31096,N_28307,N_29302);
nor U31097 (N_31097,N_28716,N_25371);
and U31098 (N_31098,N_26152,N_26774);
nand U31099 (N_31099,N_26626,N_25231);
nor U31100 (N_31100,N_29665,N_28130);
and U31101 (N_31101,N_29498,N_25037);
nor U31102 (N_31102,N_25781,N_28585);
nand U31103 (N_31103,N_29186,N_29908);
nand U31104 (N_31104,N_26592,N_26481);
xnor U31105 (N_31105,N_28349,N_25070);
nand U31106 (N_31106,N_26811,N_29986);
nand U31107 (N_31107,N_28666,N_29324);
nor U31108 (N_31108,N_27901,N_25275);
and U31109 (N_31109,N_26409,N_29981);
nand U31110 (N_31110,N_29813,N_29387);
or U31111 (N_31111,N_27897,N_29170);
and U31112 (N_31112,N_29301,N_25222);
and U31113 (N_31113,N_29504,N_25417);
nor U31114 (N_31114,N_28263,N_26092);
xnor U31115 (N_31115,N_29807,N_29567);
or U31116 (N_31116,N_28842,N_25128);
xnor U31117 (N_31117,N_27551,N_29946);
or U31118 (N_31118,N_27982,N_28800);
nor U31119 (N_31119,N_28812,N_29108);
xnor U31120 (N_31120,N_25250,N_25254);
and U31121 (N_31121,N_25563,N_27858);
nor U31122 (N_31122,N_26267,N_29235);
and U31123 (N_31123,N_27341,N_27135);
and U31124 (N_31124,N_25729,N_27569);
or U31125 (N_31125,N_25712,N_28351);
nand U31126 (N_31126,N_25328,N_26839);
xnor U31127 (N_31127,N_26830,N_26708);
nor U31128 (N_31128,N_29683,N_28186);
xor U31129 (N_31129,N_27679,N_25985);
or U31130 (N_31130,N_25095,N_29663);
or U31131 (N_31131,N_26552,N_28291);
and U31132 (N_31132,N_29028,N_28960);
nand U31133 (N_31133,N_26002,N_29822);
xor U31134 (N_31134,N_29407,N_25461);
xor U31135 (N_31135,N_26418,N_27006);
nor U31136 (N_31136,N_25704,N_29736);
xnor U31137 (N_31137,N_29828,N_28039);
nor U31138 (N_31138,N_27406,N_29530);
nor U31139 (N_31139,N_29761,N_26319);
nor U31140 (N_31140,N_29337,N_28122);
and U31141 (N_31141,N_26448,N_28808);
nand U31142 (N_31142,N_29458,N_27455);
nor U31143 (N_31143,N_27747,N_25531);
nand U31144 (N_31144,N_26750,N_25847);
nor U31145 (N_31145,N_27380,N_25497);
nand U31146 (N_31146,N_26985,N_28968);
or U31147 (N_31147,N_25191,N_28944);
nand U31148 (N_31148,N_27441,N_25345);
nand U31149 (N_31149,N_28539,N_28995);
xnor U31150 (N_31150,N_25536,N_26950);
and U31151 (N_31151,N_27893,N_27590);
xnor U31152 (N_31152,N_25099,N_27269);
and U31153 (N_31153,N_25241,N_28641);
and U31154 (N_31154,N_29357,N_29528);
nor U31155 (N_31155,N_29492,N_29145);
and U31156 (N_31156,N_25543,N_26244);
xnor U31157 (N_31157,N_29090,N_28607);
xnor U31158 (N_31158,N_28298,N_27683);
xor U31159 (N_31159,N_26952,N_27333);
xnor U31160 (N_31160,N_25922,N_27749);
nor U31161 (N_31161,N_26430,N_28022);
xnor U31162 (N_31162,N_25149,N_27321);
or U31163 (N_31163,N_26996,N_27264);
nand U31164 (N_31164,N_28182,N_26374);
or U31165 (N_31165,N_26749,N_27592);
or U31166 (N_31166,N_28545,N_29537);
nor U31167 (N_31167,N_26270,N_28449);
or U31168 (N_31168,N_28606,N_25043);
nand U31169 (N_31169,N_26841,N_26119);
xnor U31170 (N_31170,N_25841,N_28406);
nor U31171 (N_31171,N_28689,N_29619);
nor U31172 (N_31172,N_29072,N_26022);
or U31173 (N_31173,N_29776,N_28432);
nand U31174 (N_31174,N_25472,N_26155);
or U31175 (N_31175,N_26388,N_25264);
nand U31176 (N_31176,N_29260,N_25618);
or U31177 (N_31177,N_28274,N_28034);
and U31178 (N_31178,N_29242,N_25255);
or U31179 (N_31179,N_27766,N_28181);
or U31180 (N_31180,N_26723,N_27168);
or U31181 (N_31181,N_29158,N_28191);
or U31182 (N_31182,N_27838,N_26599);
nand U31183 (N_31183,N_25955,N_29209);
xor U31184 (N_31184,N_29700,N_26008);
and U31185 (N_31185,N_28238,N_26499);
or U31186 (N_31186,N_29713,N_27919);
nand U31187 (N_31187,N_26365,N_27910);
xnor U31188 (N_31188,N_25203,N_26376);
nor U31189 (N_31189,N_27137,N_25983);
or U31190 (N_31190,N_27632,N_26742);
or U31191 (N_31191,N_28852,N_29185);
or U31192 (N_31192,N_25715,N_26031);
nor U31193 (N_31193,N_25526,N_29296);
or U31194 (N_31194,N_26957,N_29486);
nor U31195 (N_31195,N_29011,N_29734);
and U31196 (N_31196,N_25927,N_29568);
nand U31197 (N_31197,N_29604,N_29703);
nand U31198 (N_31198,N_26643,N_29194);
nor U31199 (N_31199,N_26186,N_29968);
xnor U31200 (N_31200,N_27202,N_27547);
xor U31201 (N_31201,N_27184,N_28729);
or U31202 (N_31202,N_27075,N_26524);
xor U31203 (N_31203,N_27088,N_27875);
nand U31204 (N_31204,N_27975,N_29267);
xor U31205 (N_31205,N_28259,N_26837);
nand U31206 (N_31206,N_26094,N_27266);
nor U31207 (N_31207,N_28204,N_25306);
xor U31208 (N_31208,N_29516,N_26864);
nand U31209 (N_31209,N_28171,N_26591);
nand U31210 (N_31210,N_25940,N_26655);
and U31211 (N_31211,N_28596,N_25256);
nor U31212 (N_31212,N_25080,N_29274);
and U31213 (N_31213,N_25549,N_25640);
or U31214 (N_31214,N_25434,N_28741);
or U31215 (N_31215,N_27140,N_28935);
nor U31216 (N_31216,N_29653,N_27775);
nand U31217 (N_31217,N_25502,N_25797);
nor U31218 (N_31218,N_28297,N_28899);
and U31219 (N_31219,N_27960,N_27983);
nor U31220 (N_31220,N_26355,N_28266);
nor U31221 (N_31221,N_26797,N_28489);
or U31222 (N_31222,N_27937,N_26209);
nor U31223 (N_31223,N_29870,N_25831);
nor U31224 (N_31224,N_25682,N_28869);
nor U31225 (N_31225,N_25584,N_25463);
xnor U31226 (N_31226,N_28288,N_29814);
nand U31227 (N_31227,N_27620,N_25325);
or U31228 (N_31228,N_25139,N_29915);
or U31229 (N_31229,N_29100,N_25778);
and U31230 (N_31230,N_28501,N_26420);
or U31231 (N_31231,N_26343,N_28373);
xor U31232 (N_31232,N_28985,N_29377);
nand U31233 (N_31233,N_29768,N_28357);
or U31234 (N_31234,N_27540,N_27633);
xor U31235 (N_31235,N_27004,N_29022);
nand U31236 (N_31236,N_27059,N_26285);
nor U31237 (N_31237,N_26691,N_29723);
nand U31238 (N_31238,N_28137,N_29067);
and U31239 (N_31239,N_29926,N_25028);
nand U31240 (N_31240,N_28609,N_28761);
nand U31241 (N_31241,N_27126,N_26947);
nand U31242 (N_31242,N_27280,N_29991);
nor U31243 (N_31243,N_25111,N_27203);
nor U31244 (N_31244,N_28822,N_25475);
nor U31245 (N_31245,N_25590,N_29901);
and U31246 (N_31246,N_26568,N_29420);
xor U31247 (N_31247,N_27299,N_26904);
xor U31248 (N_31248,N_27435,N_28200);
xnor U31249 (N_31249,N_28350,N_25664);
nor U31250 (N_31250,N_25930,N_27779);
and U31251 (N_31251,N_28227,N_29818);
xnor U31252 (N_31252,N_28172,N_25115);
xor U31253 (N_31253,N_28904,N_25769);
or U31254 (N_31254,N_25058,N_29790);
and U31255 (N_31255,N_26787,N_27255);
nand U31256 (N_31256,N_28813,N_28526);
and U31257 (N_31257,N_27794,N_27883);
or U31258 (N_31258,N_29900,N_29637);
or U31259 (N_31259,N_27174,N_27087);
and U31260 (N_31260,N_26459,N_28591);
or U31261 (N_31261,N_28725,N_28659);
and U31262 (N_31262,N_26954,N_26176);
and U31263 (N_31263,N_25174,N_26659);
nor U31264 (N_31264,N_29096,N_25591);
and U31265 (N_31265,N_25398,N_26632);
or U31266 (N_31266,N_29849,N_28516);
nor U31267 (N_31267,N_27525,N_27585);
nor U31268 (N_31268,N_27056,N_28906);
xnor U31269 (N_31269,N_26000,N_28764);
xnor U31270 (N_31270,N_25914,N_25150);
or U31271 (N_31271,N_28794,N_26752);
or U31272 (N_31272,N_27579,N_25560);
nor U31273 (N_31273,N_27036,N_25426);
and U31274 (N_31274,N_27725,N_26536);
nor U31275 (N_31275,N_25976,N_25427);
nand U31276 (N_31276,N_26478,N_28874);
nor U31277 (N_31277,N_25503,N_26398);
xor U31278 (N_31278,N_25871,N_25717);
or U31279 (N_31279,N_26821,N_25114);
nor U31280 (N_31280,N_26329,N_25489);
or U31281 (N_31281,N_29615,N_27145);
or U31282 (N_31282,N_29582,N_27127);
or U31283 (N_31283,N_26564,N_28093);
nand U31284 (N_31284,N_28469,N_27648);
or U31285 (N_31285,N_29805,N_26153);
xor U31286 (N_31286,N_28824,N_26610);
nor U31287 (N_31287,N_28872,N_29348);
or U31288 (N_31288,N_29638,N_26794);
and U31289 (N_31289,N_28167,N_28392);
xnor U31290 (N_31290,N_27850,N_29002);
xnor U31291 (N_31291,N_28056,N_29406);
nor U31292 (N_31292,N_27852,N_25086);
or U31293 (N_31293,N_26108,N_28050);
and U31294 (N_31294,N_26801,N_27892);
nand U31295 (N_31295,N_26068,N_26616);
or U31296 (N_31296,N_26203,N_29404);
and U31297 (N_31297,N_27911,N_25557);
or U31298 (N_31298,N_28440,N_25331);
or U31299 (N_31299,N_29364,N_25303);
and U31300 (N_31300,N_28695,N_27622);
and U31301 (N_31301,N_26320,N_26391);
nor U31302 (N_31302,N_27881,N_26366);
or U31303 (N_31303,N_26377,N_28409);
nor U31304 (N_31304,N_25817,N_25555);
nor U31305 (N_31305,N_27328,N_28402);
nand U31306 (N_31306,N_26972,N_25906);
nand U31307 (N_31307,N_27013,N_27740);
nand U31308 (N_31308,N_27294,N_29423);
xnor U31309 (N_31309,N_25382,N_25057);
nor U31310 (N_31310,N_27953,N_27539);
or U31311 (N_31311,N_25631,N_28934);
xnor U31312 (N_31312,N_29518,N_25094);
and U31313 (N_31313,N_28092,N_28949);
nor U31314 (N_31314,N_29154,N_28707);
nand U31315 (N_31315,N_26771,N_28358);
or U31316 (N_31316,N_27297,N_26219);
and U31317 (N_31317,N_25931,N_27107);
xnor U31318 (N_31318,N_26570,N_28967);
xor U31319 (N_31319,N_29688,N_27695);
nor U31320 (N_31320,N_25212,N_28544);
or U31321 (N_31321,N_28957,N_29473);
and U31322 (N_31322,N_27270,N_29340);
nand U31323 (N_31323,N_29664,N_29960);
nand U31324 (N_31324,N_25022,N_27555);
nand U31325 (N_31325,N_26566,N_29943);
and U31326 (N_31326,N_27465,N_28178);
nand U31327 (N_31327,N_29369,N_26497);
xor U31328 (N_31328,N_25853,N_25822);
xnor U31329 (N_31329,N_26190,N_25042);
nor U31330 (N_31330,N_27125,N_25192);
or U31331 (N_31331,N_25104,N_29277);
nor U31332 (N_31332,N_27032,N_29754);
nor U31333 (N_31333,N_27619,N_29297);
nor U31334 (N_31334,N_28049,N_29037);
xor U31335 (N_31335,N_28691,N_25650);
xor U31336 (N_31336,N_27802,N_26580);
or U31337 (N_31337,N_25764,N_26979);
xnor U31338 (N_31338,N_26414,N_25907);
or U31339 (N_31339,N_27346,N_26927);
nand U31340 (N_31340,N_27045,N_28179);
xnor U31341 (N_31341,N_26894,N_28802);
or U31342 (N_31342,N_26802,N_27991);
and U31343 (N_31343,N_26556,N_25678);
nor U31344 (N_31344,N_29017,N_26231);
and U31345 (N_31345,N_28087,N_26831);
or U31346 (N_31346,N_28758,N_29681);
nand U31347 (N_31347,N_27287,N_29678);
nand U31348 (N_31348,N_26472,N_26058);
or U31349 (N_31349,N_27826,N_28893);
nand U31350 (N_31350,N_25091,N_25695);
nor U31351 (N_31351,N_26662,N_26252);
xor U31352 (N_31352,N_26959,N_25189);
or U31353 (N_31353,N_27945,N_26615);
xnor U31354 (N_31354,N_28342,N_26938);
and U31355 (N_31355,N_26282,N_28320);
or U31356 (N_31356,N_28580,N_29554);
nor U31357 (N_31357,N_26760,N_25258);
and U31358 (N_31358,N_27240,N_28736);
or U31359 (N_31359,N_25199,N_28407);
xor U31360 (N_31360,N_26513,N_29450);
and U31361 (N_31361,N_27752,N_25950);
or U31362 (N_31362,N_28442,N_29388);
nand U31363 (N_31363,N_26041,N_28436);
xnor U31364 (N_31364,N_25593,N_27104);
nor U31365 (N_31365,N_29682,N_25155);
nor U31366 (N_31366,N_26753,N_29137);
xnor U31367 (N_31367,N_28991,N_27932);
or U31368 (N_31368,N_29273,N_28303);
xnor U31369 (N_31369,N_25045,N_29336);
and U31370 (N_31370,N_27091,N_27987);
xnor U31371 (N_31371,N_29430,N_28280);
nor U31372 (N_31372,N_29331,N_26956);
xor U31373 (N_31373,N_29322,N_28221);
or U31374 (N_31374,N_29756,N_26140);
nand U31375 (N_31375,N_26348,N_27726);
and U31376 (N_31376,N_26576,N_27223);
and U31377 (N_31377,N_26016,N_27370);
xor U31378 (N_31378,N_29990,N_26184);
nand U31379 (N_31379,N_28100,N_26222);
or U31380 (N_31380,N_29985,N_27513);
nand U31381 (N_31381,N_27509,N_28931);
xnor U31382 (N_31382,N_26832,N_28938);
and U31383 (N_31383,N_26853,N_27961);
nand U31384 (N_31384,N_27044,N_26544);
or U31385 (N_31385,N_25153,N_25963);
xnor U31386 (N_31386,N_29840,N_25092);
nand U31387 (N_31387,N_29808,N_28818);
xnor U31388 (N_31388,N_26380,N_26423);
nand U31389 (N_31389,N_27822,N_28770);
or U31390 (N_31390,N_25598,N_26142);
nand U31391 (N_31391,N_28364,N_26495);
nand U31392 (N_31392,N_27788,N_29104);
xnor U31393 (N_31393,N_29772,N_29342);
nor U31394 (N_31394,N_29030,N_25898);
and U31395 (N_31395,N_27872,N_28829);
and U31396 (N_31396,N_27915,N_25876);
nor U31397 (N_31397,N_28078,N_26051);
nand U31398 (N_31398,N_26600,N_25314);
xnor U31399 (N_31399,N_26215,N_29464);
or U31400 (N_31400,N_25803,N_25219);
nand U31401 (N_31401,N_27746,N_27347);
nor U31402 (N_31402,N_29719,N_26088);
nand U31403 (N_31403,N_28825,N_26590);
nor U31404 (N_31404,N_26138,N_29850);
xor U31405 (N_31405,N_27114,N_25190);
nand U31406 (N_31406,N_27721,N_27008);
nor U31407 (N_31407,N_25455,N_26037);
nor U31408 (N_31408,N_28914,N_27627);
and U31409 (N_31409,N_25202,N_29040);
and U31410 (N_31410,N_28901,N_29294);
and U31411 (N_31411,N_26469,N_28503);
xnor U31412 (N_31412,N_27964,N_26177);
nand U31413 (N_31413,N_28682,N_29821);
or U31414 (N_31414,N_27667,N_25430);
or U31415 (N_31415,N_27344,N_28756);
or U31416 (N_31416,N_28929,N_25366);
nor U31417 (N_31417,N_26288,N_26259);
and U31418 (N_31418,N_28983,N_27398);
nor U31419 (N_31419,N_29092,N_28592);
nand U31420 (N_31420,N_29669,N_28145);
nor U31421 (N_31421,N_28470,N_27671);
nor U31422 (N_31422,N_28339,N_25845);
nor U31423 (N_31423,N_29695,N_28754);
or U31424 (N_31424,N_25728,N_28124);
nor U31425 (N_31425,N_25570,N_27189);
nor U31426 (N_31426,N_27139,N_25658);
nand U31427 (N_31427,N_25046,N_26854);
xor U31428 (N_31428,N_27469,N_25477);
and U31429 (N_31429,N_26249,N_26519);
nand U31430 (N_31430,N_27608,N_28538);
xor U31431 (N_31431,N_28052,N_27498);
or U31432 (N_31432,N_29526,N_28314);
or U31433 (N_31433,N_28371,N_29469);
or U31434 (N_31434,N_29180,N_29412);
or U31435 (N_31435,N_26081,N_25794);
and U31436 (N_31436,N_29592,N_26763);
nor U31437 (N_31437,N_27007,N_26850);
xor U31438 (N_31438,N_29315,N_25492);
xnor U31439 (N_31439,N_29393,N_28217);
or U31440 (N_31440,N_28690,N_27692);
or U31441 (N_31441,N_27697,N_26822);
and U31442 (N_31442,N_29699,N_26980);
nand U31443 (N_31443,N_25670,N_25604);
and U31444 (N_31444,N_28000,N_27023);
nand U31445 (N_31445,N_26824,N_27310);
nand U31446 (N_31446,N_28616,N_28814);
or U31447 (N_31447,N_28952,N_27496);
nand U31448 (N_31448,N_28999,N_25085);
nor U31449 (N_31449,N_25636,N_26964);
or U31450 (N_31450,N_27283,N_25689);
xor U31451 (N_31451,N_25733,N_27097);
and U31452 (N_31452,N_26628,N_29806);
or U31453 (N_31453,N_26868,N_26697);
xnor U31454 (N_31454,N_29797,N_28811);
or U31455 (N_31455,N_25084,N_25516);
or U31456 (N_31456,N_26692,N_25318);
and U31457 (N_31457,N_27787,N_29707);
xor U31458 (N_31458,N_26738,N_25866);
nor U31459 (N_31459,N_27361,N_26373);
or U31460 (N_31460,N_29543,N_25966);
xor U31461 (N_31461,N_26308,N_27643);
or U31462 (N_31462,N_26410,N_28046);
nor U31463 (N_31463,N_29217,N_27869);
xnor U31464 (N_31464,N_27537,N_29876);
nand U31465 (N_31465,N_28593,N_29742);
xnor U31466 (N_31466,N_28446,N_29685);
nor U31467 (N_31467,N_25339,N_28947);
xor U31468 (N_31468,N_25201,N_27732);
or U31469 (N_31469,N_27605,N_26228);
or U31470 (N_31470,N_28008,N_27635);
nand U31471 (N_31471,N_25980,N_25585);
or U31472 (N_31472,N_28881,N_25105);
xor U31473 (N_31473,N_25952,N_28554);
and U31474 (N_31474,N_27675,N_27065);
nor U31475 (N_31475,N_29264,N_28496);
or U31476 (N_31476,N_27433,N_27554);
and U31477 (N_31477,N_29341,N_28193);
and U31478 (N_31478,N_27372,N_25474);
nor U31479 (N_31479,N_25538,N_27268);
and U31480 (N_31480,N_25756,N_28359);
xor U31481 (N_31481,N_25660,N_27084);
nand U31482 (N_31482,N_28412,N_28923);
nor U31483 (N_31483,N_25013,N_25788);
and U31484 (N_31484,N_27577,N_26790);
and U31485 (N_31485,N_26300,N_28258);
nand U31486 (N_31486,N_28753,N_26553);
nor U31487 (N_31487,N_25238,N_29066);
nor U31488 (N_31488,N_26838,N_27472);
or U31489 (N_31489,N_27524,N_28408);
or U31490 (N_31490,N_29320,N_29359);
or U31491 (N_31491,N_29804,N_25911);
nand U31492 (N_31492,N_26902,N_26514);
or U31493 (N_31493,N_25471,N_28882);
xnor U31494 (N_31494,N_28711,N_26920);
nand U31495 (N_31495,N_26942,N_25798);
or U31496 (N_31496,N_27133,N_28862);
nor U31497 (N_31497,N_28961,N_28529);
or U31498 (N_31498,N_28318,N_27670);
and U31499 (N_31499,N_28473,N_29447);
or U31500 (N_31500,N_27757,N_29662);
and U31501 (N_31501,N_26714,N_28370);
xnor U31502 (N_31502,N_27681,N_29466);
or U31503 (N_31503,N_29292,N_28807);
nand U31504 (N_31504,N_28212,N_27068);
or U31505 (N_31505,N_26474,N_29611);
xnor U31506 (N_31506,N_27095,N_26251);
and U31507 (N_31507,N_26769,N_29093);
or U31508 (N_31508,N_28877,N_29675);
nor U31509 (N_31509,N_27839,N_25957);
and U31510 (N_31510,N_27129,N_27386);
xnor U31511 (N_31511,N_28149,N_25368);
nand U31512 (N_31512,N_28702,N_25939);
xnor U31513 (N_31513,N_26013,N_27610);
and U31514 (N_31514,N_28793,N_28480);
or U31515 (N_31515,N_25148,N_26558);
and U31516 (N_31516,N_26807,N_26851);
xnor U31517 (N_31517,N_28427,N_29846);
or U31518 (N_31518,N_29461,N_25718);
nor U31519 (N_31519,N_28323,N_28306);
nor U31520 (N_31520,N_26779,N_28250);
nor U31521 (N_31521,N_25286,N_28779);
nor U31522 (N_31522,N_27432,N_26018);
xnor U31523 (N_31523,N_28839,N_29491);
nand U31524 (N_31524,N_29762,N_26387);
xor U31525 (N_31525,N_25751,N_25755);
xor U31526 (N_31526,N_25758,N_26360);
or U31527 (N_31527,N_29503,N_25601);
nand U31528 (N_31528,N_27458,N_26317);
nand U31529 (N_31529,N_26180,N_27918);
xor U31530 (N_31530,N_29735,N_27628);
nand U31531 (N_31531,N_26227,N_26761);
nor U31532 (N_31532,N_28128,N_25116);
or U31533 (N_31533,N_29562,N_27546);
or U31534 (N_31534,N_25564,N_29909);
xor U31535 (N_31535,N_27325,N_28587);
nor U31536 (N_31536,N_27810,N_26963);
nand U31537 (N_31537,N_25826,N_28563);
or U31538 (N_31538,N_29899,N_27233);
or U31539 (N_31539,N_25458,N_29852);
or U31540 (N_31540,N_29027,N_29042);
or U31541 (N_31541,N_25804,N_28684);
nor U31542 (N_31542,N_25681,N_27001);
or U31543 (N_31543,N_28158,N_29416);
nor U31544 (N_31544,N_28604,N_27624);
and U31545 (N_31545,N_25620,N_27136);
and U31546 (N_31546,N_28422,N_25265);
or U31547 (N_31547,N_26236,N_28099);
and U31548 (N_31548,N_27698,N_25653);
and U31549 (N_31549,N_28057,N_25964);
and U31550 (N_31550,N_25645,N_26130);
and U31551 (N_31551,N_29472,N_29202);
nand U31552 (N_31552,N_29280,N_29508);
nand U31553 (N_31553,N_28481,N_27742);
and U31554 (N_31554,N_28311,N_28071);
xor U31555 (N_31555,N_28116,N_28621);
and U31556 (N_31556,N_28505,N_25440);
or U31557 (N_31557,N_27222,N_26860);
and U31558 (N_31558,N_29751,N_26503);
nand U31559 (N_31559,N_29199,N_27339);
nand U31560 (N_31560,N_27379,N_25785);
nand U31561 (N_31561,N_26255,N_29287);
and U31562 (N_31562,N_28120,N_29558);
nand U31563 (N_31563,N_29058,N_29895);
nor U31564 (N_31564,N_27113,N_26232);
and U31565 (N_31565,N_27615,N_25147);
nand U31566 (N_31566,N_27123,N_26482);
xnor U31567 (N_31567,N_28232,N_27981);
nand U31568 (N_31568,N_27761,N_27493);
and U31569 (N_31569,N_26392,N_25625);
xnor U31570 (N_31570,N_27818,N_29727);
nor U31571 (N_31571,N_28060,N_29454);
or U31572 (N_31572,N_27966,N_27876);
or U31573 (N_31573,N_26276,N_27920);
or U31574 (N_31574,N_28214,N_25401);
or U31575 (N_31575,N_28401,N_25962);
nand U31576 (N_31576,N_26715,N_25655);
nand U31577 (N_31577,N_26955,N_27690);
nor U31578 (N_31578,N_29506,N_29221);
nor U31579 (N_31579,N_26668,N_28353);
and U31580 (N_31580,N_27459,N_26602);
xor U31581 (N_31581,N_26757,N_27147);
or U31582 (N_31582,N_28640,N_26024);
and U31583 (N_31583,N_28327,N_25280);
nand U31584 (N_31584,N_26477,N_29488);
nand U31585 (N_31585,N_25508,N_25017);
nor U31586 (N_31586,N_26991,N_26299);
or U31587 (N_31587,N_28190,N_29376);
xnor U31588 (N_31588,N_29307,N_25997);
nand U31589 (N_31589,N_28400,N_25234);
or U31590 (N_31590,N_25060,N_27770);
xor U31591 (N_31591,N_29119,N_29368);
and U31592 (N_31592,N_26672,N_29231);
and U31593 (N_31593,N_27533,N_28183);
nor U31594 (N_31594,N_25878,N_26762);
and U31595 (N_31595,N_25353,N_25097);
and U31596 (N_31596,N_29897,N_25227);
or U31597 (N_31597,N_29826,N_28525);
and U31598 (N_31598,N_29371,N_27374);
nor U31599 (N_31599,N_29686,N_28605);
nand U31600 (N_31600,N_27829,N_25170);
and U31601 (N_31601,N_25499,N_26393);
xor U31602 (N_31602,N_28102,N_26044);
nor U31603 (N_31603,N_29572,N_28267);
or U31604 (N_31604,N_25667,N_29460);
nor U31605 (N_31605,N_29691,N_28550);
nand U31606 (N_31606,N_29398,N_29261);
nand U31607 (N_31607,N_27489,N_25810);
or U31608 (N_31608,N_29630,N_25973);
xnor U31609 (N_31609,N_25545,N_26731);
nand U31610 (N_31610,N_26848,N_25435);
nor U31611 (N_31611,N_28411,N_29829);
xor U31612 (N_31612,N_29697,N_28953);
and U31613 (N_31613,N_29189,N_26375);
or U31614 (N_31614,N_27443,N_29015);
or U31615 (N_31615,N_27828,N_27063);
xnor U31616 (N_31616,N_29254,N_25574);
or U31617 (N_31617,N_27230,N_26033);
xor U31618 (N_31618,N_26350,N_26253);
or U31619 (N_31619,N_26015,N_25638);
nor U31620 (N_31620,N_26258,N_29788);
nor U31621 (N_31621,N_29941,N_26256);
nand U31622 (N_31622,N_28272,N_27096);
nand U31623 (N_31623,N_29585,N_26073);
nor U31624 (N_31624,N_26748,N_27553);
or U31625 (N_31625,N_28115,N_26170);
nand U31626 (N_31626,N_26732,N_25573);
xnor U31627 (N_31627,N_27862,N_26501);
nand U31628 (N_31628,N_28246,N_28936);
nor U31629 (N_31629,N_28108,N_28932);
nand U31630 (N_31630,N_25373,N_26325);
nor U31631 (N_31631,N_29706,N_25271);
and U31632 (N_31632,N_29403,N_27573);
xnor U31633 (N_31633,N_28870,N_28885);
nand U31634 (N_31634,N_25552,N_27453);
nor U31635 (N_31635,N_25550,N_28103);
nand U31636 (N_31636,N_27930,N_29945);
and U31637 (N_31637,N_25686,N_26007);
xor U31638 (N_31638,N_27823,N_27047);
xnor U31639 (N_31639,N_26077,N_26189);
nand U31640 (N_31640,N_26966,N_26627);
nor U31641 (N_31641,N_29045,N_28010);
and U31642 (N_31642,N_28928,N_29026);
nand U31643 (N_31643,N_29874,N_26817);
nand U31644 (N_31644,N_25735,N_28732);
or U31645 (N_31645,N_27475,N_26812);
nor U31646 (N_31646,N_25465,N_26719);
nand U31647 (N_31647,N_28903,N_25854);
xnor U31648 (N_31648,N_26453,N_26115);
and U31649 (N_31649,N_26740,N_28223);
and U31650 (N_31650,N_29601,N_25801);
and U31651 (N_31651,N_26563,N_25627);
xor U31652 (N_31652,N_25918,N_28140);
nand U31653 (N_31653,N_27025,N_25816);
nor U31654 (N_31654,N_28878,N_28768);
nor U31655 (N_31655,N_25748,N_28062);
nor U31656 (N_31656,N_29892,N_25836);
nand U31657 (N_31657,N_28698,N_28980);
xor U31658 (N_31658,N_26462,N_25261);
or U31659 (N_31659,N_27564,N_28642);
or U31660 (N_31660,N_26588,N_29512);
and U31661 (N_31661,N_27706,N_27315);
or U31662 (N_31662,N_28325,N_27249);
and U31663 (N_31663,N_25007,N_28649);
xor U31664 (N_31664,N_28925,N_27896);
nand U31665 (N_31665,N_27152,N_28927);
nand U31666 (N_31666,N_25229,N_28429);
nor U31667 (N_31667,N_29197,N_26765);
nand U31668 (N_31668,N_26654,N_25386);
and U31669 (N_31669,N_28635,N_25379);
xnor U31670 (N_31670,N_27460,N_28575);
or U31671 (N_31671,N_28582,N_29073);
nor U31672 (N_31672,N_28031,N_28708);
or U31673 (N_31673,N_26575,N_25671);
nor U31674 (N_31674,N_29271,N_29599);
or U31675 (N_31675,N_25873,N_27713);
nor U31676 (N_31676,N_28515,N_27532);
and U31677 (N_31677,N_29007,N_27859);
nand U31678 (N_31678,N_29205,N_25971);
and U31679 (N_31679,N_25674,N_25761);
nand U31680 (N_31680,N_26709,N_29832);
or U31681 (N_31681,N_27214,N_29799);
xnor U31682 (N_31682,N_27833,N_27167);
nor U31683 (N_31683,N_27853,N_26160);
nor U31684 (N_31684,N_27647,N_27180);
nand U31685 (N_31685,N_28855,N_26283);
or U31686 (N_31686,N_25300,N_28836);
and U31687 (N_31687,N_25101,N_29774);
or U31688 (N_31688,N_29886,N_26467);
and U31689 (N_31689,N_27150,N_25054);
and U31690 (N_31690,N_28993,N_29005);
nor U31691 (N_31691,N_27656,N_26843);
or U31692 (N_31692,N_26370,N_28338);
nand U31693 (N_31693,N_28536,N_25974);
nor U31694 (N_31694,N_25049,N_27528);
nand U31695 (N_31695,N_29493,N_28875);
or U31696 (N_31696,N_28026,N_26529);
nor U31697 (N_31697,N_27194,N_27451);
and U31698 (N_31698,N_28423,N_25493);
nor U31699 (N_31699,N_25915,N_26014);
nor U31700 (N_31700,N_26946,N_26454);
nor U31701 (N_31701,N_27494,N_28574);
nor U31702 (N_31702,N_29872,N_29048);
xnor U31703 (N_31703,N_25607,N_25454);
nor U31704 (N_31704,N_27835,N_25629);
nor U31705 (N_31705,N_25835,N_27423);
or U31706 (N_31706,N_27134,N_29361);
or U31707 (N_31707,N_27969,N_28065);
and U31708 (N_31708,N_26810,N_28570);
nand U31709 (N_31709,N_28520,N_25562);
xnor U31710 (N_31710,N_28148,N_29481);
or U31711 (N_31711,N_25509,N_26399);
and U31712 (N_31712,N_28510,N_28117);
or U31713 (N_31713,N_28343,N_25893);
nand U31714 (N_31714,N_27428,N_25652);
nor U31715 (N_31715,N_27195,N_29798);
nor U31716 (N_31716,N_28176,N_27512);
nor U31717 (N_31717,N_29933,N_25772);
nand U31718 (N_31718,N_27021,N_27307);
xor U31719 (N_31719,N_28891,N_25680);
and U31720 (N_31720,N_29542,N_26262);
or U31721 (N_31721,N_29024,N_28933);
nand U31722 (N_31722,N_26767,N_28776);
xnor U31723 (N_31723,N_29626,N_26508);
nand U31724 (N_31724,N_27296,N_28157);
nor U31725 (N_31725,N_29787,N_28614);
and U31726 (N_31726,N_28530,N_29532);
xor U31727 (N_31727,N_26906,N_27598);
nor U31728 (N_31728,N_26001,N_25418);
nand U31729 (N_31729,N_28150,N_29603);
and U31730 (N_31730,N_26630,N_28094);
nor U31731 (N_31731,N_29228,N_29743);
and U31732 (N_31732,N_26650,N_29039);
nand U31733 (N_31733,N_26847,N_25511);
nand U31734 (N_31734,N_29778,N_25397);
and U31735 (N_31735,N_25343,N_27923);
xnor U31736 (N_31736,N_29332,N_26061);
or U31737 (N_31737,N_28009,N_29858);
nand U31738 (N_31738,N_25400,N_25518);
xor U31739 (N_31739,N_25005,N_25633);
xor U31740 (N_31740,N_26939,N_29349);
xor U31741 (N_31741,N_27466,N_28637);
and U31742 (N_31742,N_25145,N_29442);
and U31743 (N_31743,N_26608,N_28209);
or U31744 (N_31744,N_29513,N_26584);
nor U31745 (N_31745,N_26828,N_29219);
nor U31746 (N_31746,N_25253,N_26449);
nand U31747 (N_31747,N_29588,N_29710);
or U31748 (N_31748,N_25792,N_26124);
and U31749 (N_31749,N_29305,N_26605);
nor U31750 (N_31750,N_29740,N_28324);
and U31751 (N_31751,N_28315,N_26312);
and U31752 (N_31752,N_27800,N_27302);
and U31753 (N_31753,N_28821,N_28610);
or U31754 (N_31754,N_25406,N_26039);
or U31755 (N_31755,N_25732,N_29263);
and U31756 (N_31756,N_25901,N_27215);
nand U31757 (N_31757,N_26687,N_29769);
and U31758 (N_31758,N_26342,N_25805);
or U31759 (N_31759,N_27593,N_25273);
nor U31760 (N_31760,N_28755,N_28541);
and U31761 (N_31761,N_25259,N_27895);
xor U31762 (N_31762,N_29213,N_29327);
nand U31763 (N_31763,N_29210,N_25240);
xnor U31764 (N_31764,N_28686,N_28251);
nor U31765 (N_31765,N_28718,N_25335);
nor U31766 (N_31766,N_27994,N_28945);
or U31767 (N_31767,N_25055,N_28245);
and U31768 (N_31768,N_26268,N_26532);
xnor U31769 (N_31769,N_27735,N_29286);
nand U31770 (N_31770,N_26884,N_26400);
xnor U31771 (N_31771,N_28131,N_27815);
nor U31772 (N_31772,N_29150,N_27914);
and U31773 (N_31773,N_25984,N_29702);
and U31774 (N_31774,N_28170,N_29215);
nand U31775 (N_31775,N_28027,N_28742);
xor U31776 (N_31776,N_25864,N_28972);
nand U31777 (N_31777,N_28458,N_27704);
nor U31778 (N_31778,N_28165,N_29262);
nand U31779 (N_31779,N_28433,N_29009);
or U31780 (N_31780,N_28229,N_25581);
nand U31781 (N_31781,N_27515,N_27926);
or U31782 (N_31782,N_25500,N_26826);
and U31783 (N_31783,N_25359,N_25301);
nand U31784 (N_31784,N_28236,N_29984);
nor U31785 (N_31785,N_29660,N_27464);
xor U31786 (N_31786,N_25341,N_27534);
nand U31787 (N_31787,N_28743,N_25534);
nand U31788 (N_31788,N_27388,N_29672);
and U31789 (N_31789,N_25443,N_27705);
xor U31790 (N_31790,N_28077,N_25347);
xor U31791 (N_31791,N_28697,N_26683);
and U31792 (N_31792,N_28395,N_25892);
and U31793 (N_31793,N_28565,N_25861);
and U31794 (N_31794,N_26116,N_26540);
nor U31795 (N_31795,N_27980,N_27350);
or U31796 (N_31796,N_25134,N_26684);
xor U31797 (N_31797,N_28110,N_27611);
xor U31798 (N_31798,N_25166,N_29366);
nand U31799 (N_31799,N_29642,N_28675);
and U31800 (N_31800,N_25445,N_29718);
xor U31801 (N_31801,N_29916,N_27281);
and U31802 (N_31802,N_27612,N_28611);
and U31803 (N_31803,N_26617,N_28255);
or U31804 (N_31804,N_27902,N_28276);
xor U31805 (N_31805,N_26336,N_26646);
and U31806 (N_31806,N_26623,N_27043);
nand U31807 (N_31807,N_28662,N_25802);
or U31808 (N_31808,N_27999,N_29617);
nor U31809 (N_31809,N_25517,N_27520);
xnor U31810 (N_31810,N_26743,N_29098);
nor U31811 (N_31811,N_25782,N_25495);
nand U31812 (N_31812,N_26741,N_27967);
nand U31813 (N_31813,N_25675,N_28097);
and U31814 (N_31814,N_27500,N_25164);
or U31815 (N_31815,N_25469,N_25857);
nor U31816 (N_31816,N_26146,N_27846);
nand U31817 (N_31817,N_27562,N_27156);
and U31818 (N_31818,N_29605,N_26973);
nor U31819 (N_31819,N_26674,N_28237);
nor U31820 (N_31820,N_26882,N_27674);
and U31821 (N_31821,N_27213,N_29019);
xnor U31822 (N_31822,N_28205,N_28589);
xor U31823 (N_31823,N_28791,N_27026);
nand U31824 (N_31824,N_27033,N_28531);
nor U31825 (N_31825,N_26102,N_27599);
nand U31826 (N_31826,N_28461,N_28194);
and U31827 (N_31827,N_25814,N_26739);
and U31828 (N_31828,N_26914,N_28674);
xor U31829 (N_31829,N_29654,N_28688);
and U31830 (N_31830,N_26390,N_26324);
nand U31831 (N_31831,N_26250,N_26517);
nand U31832 (N_31832,N_27899,N_26679);
xnor U31833 (N_31833,N_26026,N_25044);
xor U31834 (N_31834,N_29882,N_29115);
nand U31835 (N_31835,N_27413,N_29156);
nand U31836 (N_31836,N_28147,N_25457);
nor U31837 (N_31837,N_29577,N_29383);
or U31838 (N_31838,N_27364,N_25800);
nand U31839 (N_31839,N_29684,N_26010);
nor U31840 (N_31840,N_29405,N_28341);
and U31841 (N_31841,N_25644,N_29842);
nor U31842 (N_31842,N_27750,N_26813);
and U31843 (N_31843,N_28537,N_28381);
nor U31844 (N_31844,N_28706,N_26836);
xnor U31845 (N_31845,N_26230,N_29835);
and U31846 (N_31846,N_28962,N_27461);
or U31847 (N_31847,N_29478,N_29252);
xor U31848 (N_31848,N_27197,N_27691);
or U31849 (N_31849,N_28138,N_25419);
nand U31850 (N_31850,N_25486,N_28070);
and U31851 (N_31851,N_25724,N_28081);
nand U31852 (N_31852,N_27978,N_27730);
nand U31853 (N_31853,N_25226,N_29792);
and U31854 (N_31854,N_27301,N_27623);
and U31855 (N_31855,N_29417,N_25002);
nor U31856 (N_31856,N_26859,N_27661);
xnor U31857 (N_31857,N_28911,N_29018);
and U31858 (N_31858,N_25066,N_28654);
nor U31859 (N_31859,N_27445,N_25252);
nand U31860 (N_31860,N_29987,N_29980);
nand U31861 (N_31861,N_28335,N_29345);
or U31862 (N_31862,N_26618,N_26038);
nor U31863 (N_31863,N_28748,N_29759);
and U31864 (N_31864,N_28871,N_27561);
or U31865 (N_31865,N_28275,N_29239);
nor U31866 (N_31866,N_26892,N_27085);
nor U31867 (N_31867,N_28051,N_29650);
and U31868 (N_31868,N_26199,N_29730);
and U31869 (N_31869,N_27955,N_26113);
xor U31870 (N_31870,N_28801,N_29207);
nor U31871 (N_31871,N_29922,N_29395);
nor U31872 (N_31872,N_26075,N_29918);
or U31873 (N_31873,N_25291,N_27330);
nand U31874 (N_31874,N_27371,N_26239);
and U31875 (N_31875,N_27072,N_26434);
and U31876 (N_31876,N_28810,N_25100);
and U31877 (N_31877,N_27282,N_26264);
nand U31878 (N_31878,N_28671,N_26657);
or U31879 (N_31879,N_26127,N_26466);
and U31880 (N_31880,N_27916,N_26122);
and U31881 (N_31881,N_26021,N_26134);
nor U31882 (N_31882,N_29354,N_27820);
xor U31883 (N_31883,N_29462,N_27840);
or U31884 (N_31884,N_25793,N_29198);
xnor U31885 (N_31885,N_27778,N_27825);
xnor U31886 (N_31886,N_26527,N_28462);
nand U31887 (N_31887,N_29545,N_27192);
nand U31888 (N_31888,N_25909,N_26076);
nor U31889 (N_31889,N_27101,N_29794);
nand U31890 (N_31890,N_26653,N_27373);
nor U31891 (N_31891,N_26159,N_27020);
nand U31892 (N_31892,N_29674,N_25887);
or U31893 (N_31893,N_25102,N_26154);
nor U31894 (N_31894,N_28806,N_27332);
or U31895 (N_31895,N_28723,N_29894);
and U31896 (N_31896,N_27863,N_26705);
and U31897 (N_31897,N_28330,N_28006);
and U31898 (N_31898,N_29830,N_27422);
nor U31899 (N_31899,N_29938,N_26565);
or U31900 (N_31900,N_29112,N_26384);
nand U31901 (N_31901,N_27578,N_26208);
nor U31902 (N_31902,N_28492,N_28413);
nor U31903 (N_31903,N_26661,N_27288);
xnor U31904 (N_31904,N_25710,N_26845);
nor U31905 (N_31905,N_27970,N_26378);
nand U31906 (N_31906,N_26487,N_28139);
xor U31907 (N_31907,N_27176,N_26833);
or U31908 (N_31908,N_25575,N_27479);
xnor U31909 (N_31909,N_25236,N_26988);
nand U31910 (N_31910,N_25078,N_27587);
nand U31911 (N_31911,N_29293,N_25572);
xor U31912 (N_31912,N_29101,N_27449);
xnor U31913 (N_31913,N_25446,N_25200);
xnor U31914 (N_31914,N_25827,N_26937);
and U31915 (N_31915,N_28485,N_28631);
or U31916 (N_31916,N_27792,N_28528);
nor U31917 (N_31917,N_27196,N_27317);
nor U31918 (N_31918,N_28385,N_29350);
or U31919 (N_31919,N_27799,N_25206);
xnor U31920 (N_31920,N_27672,N_26298);
nor U31921 (N_31921,N_28384,N_29551);
nand U31922 (N_31922,N_29701,N_28998);
or U31923 (N_31923,N_25112,N_27480);
xnor U31924 (N_31924,N_25196,N_27400);
xnor U31925 (N_31925,N_26958,N_28704);
and U31926 (N_31926,N_25544,N_26870);
nor U31927 (N_31927,N_27657,N_29006);
nand U31928 (N_31928,N_28731,N_26046);
nor U31929 (N_31929,N_27935,N_26218);
xor U31930 (N_31930,N_29549,N_27710);
or U31931 (N_31931,N_25855,N_27848);
nand U31932 (N_31932,N_27604,N_28816);
and U31933 (N_31933,N_28678,N_28700);
xor U31934 (N_31934,N_29765,N_29234);
and U31935 (N_31935,N_26577,N_29020);
or U31936 (N_31936,N_26921,N_25929);
or U31937 (N_31937,N_27501,N_29074);
and U31938 (N_31938,N_29259,N_27207);
or U31939 (N_31939,N_26639,N_26647);
nand U31940 (N_31940,N_25041,N_26890);
or U31941 (N_31941,N_28560,N_27208);
nand U31942 (N_31942,N_25330,N_27857);
or U31943 (N_31943,N_25165,N_26548);
nand U31944 (N_31944,N_26405,N_25384);
or U31945 (N_31945,N_27785,N_27703);
nor U31946 (N_31946,N_26196,N_25742);
nor U31947 (N_31947,N_29187,N_27028);
or U31948 (N_31948,N_27094,N_25416);
nand U31949 (N_31949,N_27660,N_27081);
or U31950 (N_31950,N_27684,N_26305);
or U31951 (N_31951,N_26271,N_25979);
nand U31952 (N_31952,N_29966,N_29598);
nand U31953 (N_31953,N_27957,N_28969);
or U31954 (N_31954,N_28626,N_27942);
or U31955 (N_31955,N_25015,N_29081);
or U31956 (N_31956,N_28403,N_25412);
or U31957 (N_31957,N_25568,N_26727);
nand U31958 (N_31958,N_29680,N_27544);
xnor U31959 (N_31959,N_28421,N_28673);
nor U31960 (N_31960,N_26479,N_26874);
xor U31961 (N_31961,N_28090,N_27235);
or U31962 (N_31962,N_26712,N_29676);
nor U31963 (N_31963,N_28958,N_25459);
nor U31964 (N_31964,N_28535,N_25251);
nand U31965 (N_31965,N_28856,N_26880);
nand U31966 (N_31966,N_25676,N_28028);
or U31967 (N_31967,N_25565,N_29208);
and U31968 (N_31968,N_29912,N_28241);
and U31969 (N_31969,N_27143,N_27071);
or U31970 (N_31970,N_26862,N_29071);
and U31971 (N_31971,N_26422,N_28125);
or U31972 (N_31972,N_25313,N_25121);
nor U31973 (N_31973,N_27054,N_29146);
nand U31974 (N_31974,N_29760,N_25383);
xor U31975 (N_31975,N_25186,N_26364);
nand U31976 (N_31976,N_25432,N_26878);
and U31977 (N_31977,N_29008,N_25777);
nor U31978 (N_31978,N_25981,N_28018);
xor U31979 (N_31979,N_26573,N_25982);
xnor U31980 (N_31980,N_29050,N_25488);
and U31981 (N_31981,N_25369,N_25333);
nand U31982 (N_31982,N_27936,N_27744);
nand U31983 (N_31983,N_29934,N_29875);
and U31984 (N_31984,N_28169,N_29003);
and U31985 (N_31985,N_28519,N_26280);
or U31986 (N_31986,N_25968,N_27022);
or U31987 (N_31987,N_27645,N_27241);
or U31988 (N_31988,N_27175,N_26572);
and U31989 (N_31989,N_28561,N_29729);
nor U31990 (N_31990,N_29222,N_27322);
xor U31991 (N_31991,N_26827,N_26187);
xnor U31992 (N_31992,N_26234,N_25047);
or U31993 (N_31993,N_27482,N_25144);
nand U31994 (N_31994,N_25062,N_25592);
xor U31995 (N_31995,N_25537,N_26603);
nor U31996 (N_31996,N_29243,N_29574);
nor U31997 (N_31997,N_26667,N_29602);
and U31998 (N_31998,N_28435,N_25064);
nor U31999 (N_31999,N_28088,N_26881);
nand U32000 (N_32000,N_29629,N_28196);
xor U32001 (N_32001,N_28420,N_25378);
nor U32002 (N_32002,N_29834,N_28921);
and U32003 (N_32003,N_25594,N_25350);
xor U32004 (N_32004,N_27906,N_28740);
nand U32005 (N_32005,N_26296,N_29964);
nor U32006 (N_32006,N_27490,N_25460);
nor U32007 (N_32007,N_26967,N_29496);
or U32008 (N_32008,N_25916,N_26059);
xnor U32009 (N_32009,N_26624,N_27066);
or U32010 (N_32010,N_28180,N_25808);
and U32011 (N_32011,N_29298,N_26091);
nor U32012 (N_32012,N_26273,N_26003);
nand U32013 (N_32013,N_29223,N_29737);
xor U32014 (N_32014,N_29594,N_29952);
or U32015 (N_32015,N_29741,N_29103);
or U32016 (N_32016,N_28293,N_27973);
nand U32017 (N_32017,N_25031,N_29070);
nor U32018 (N_32018,N_29128,N_28556);
nor U32019 (N_32019,N_27637,N_26799);
xor U32020 (N_32020,N_25285,N_28625);
or U32021 (N_32021,N_25479,N_26535);
or U32022 (N_32022,N_29278,N_25320);
or U32023 (N_32023,N_29088,N_27463);
nor U32024 (N_32024,N_25494,N_25890);
nand U32025 (N_32025,N_25903,N_29303);
nand U32026 (N_32026,N_28321,N_26289);
and U32027 (N_32027,N_28553,N_26901);
nor U32028 (N_32028,N_25433,N_26758);
and U32029 (N_32029,N_26141,N_29339);
or U32030 (N_32030,N_29771,N_26266);
xor U32031 (N_32031,N_29317,N_27151);
nor U32032 (N_32032,N_29258,N_28546);
and U32033 (N_32033,N_26690,N_29690);
or U32034 (N_32034,N_27984,N_27457);
or U32035 (N_32035,N_26456,N_29612);
xor U32036 (N_32036,N_29031,N_27216);
nand U32037 (N_32037,N_27806,N_25006);
xor U32038 (N_32038,N_27574,N_29091);
nor U32039 (N_32039,N_27556,N_26641);
or U32040 (N_32040,N_29521,N_25269);
or U32041 (N_32041,N_26485,N_27484);
nand U32042 (N_32042,N_25825,N_25936);
nand U32043 (N_32043,N_28763,N_25610);
nor U32044 (N_32044,N_28198,N_25665);
nor U32045 (N_32045,N_28551,N_28670);
nand U32046 (N_32046,N_26660,N_25807);
xnor U32047 (N_32047,N_29563,N_26173);
xnor U32048 (N_32048,N_26188,N_29250);
xnor U32049 (N_32049,N_28900,N_25668);
or U32050 (N_32050,N_26083,N_25870);
and U32051 (N_32051,N_29153,N_25266);
and U32052 (N_32052,N_28457,N_29666);
xnor U32053 (N_32053,N_28845,N_28372);
or U32054 (N_32054,N_27693,N_28279);
xor U32055 (N_32055,N_25267,N_28619);
xor U32056 (N_32056,N_28472,N_25450);
and U32057 (N_32057,N_25606,N_26339);
or U32058 (N_32058,N_26925,N_25175);
nand U32059 (N_32059,N_29749,N_29955);
xnor U32060 (N_32060,N_28717,N_28296);
or U32061 (N_32061,N_27630,N_26211);
or U32062 (N_32062,N_28964,N_28495);
nor U32063 (N_32063,N_29468,N_28378);
xor U32064 (N_32064,N_26823,N_27017);
xor U32065 (N_32065,N_25026,N_29967);
nand U32066 (N_32066,N_28055,N_26121);
nand U32067 (N_32067,N_29299,N_26290);
or U32068 (N_32068,N_25740,N_27696);
nand U32069 (N_32069,N_29889,N_25842);
nand U32070 (N_32070,N_25349,N_29413);
nor U32071 (N_32071,N_28091,N_28007);
xnor U32072 (N_32072,N_25065,N_29036);
xnor U32073 (N_32073,N_27762,N_25129);
and U32074 (N_32074,N_27946,N_28254);
and U32075 (N_32075,N_26327,N_29106);
xor U32076 (N_32076,N_26595,N_25444);
and U32077 (N_32077,N_28044,N_26265);
xor U32078 (N_32078,N_27237,N_26090);
or U32079 (N_32079,N_28430,N_26210);
or U32080 (N_32080,N_29752,N_25123);
or U32081 (N_32081,N_28264,N_28963);
and U32082 (N_32082,N_25482,N_25889);
nor U32083 (N_32083,N_25405,N_26982);
or U32084 (N_32084,N_29583,N_27589);
nor U32085 (N_32085,N_25040,N_28841);
xnor U32086 (N_32086,N_27842,N_25880);
nand U32087 (N_32087,N_26165,N_25399);
or U32088 (N_32088,N_26291,N_26351);
and U32089 (N_32089,N_25304,N_25027);
or U32090 (N_32090,N_28777,N_26237);
nand U32091 (N_32091,N_29497,N_25284);
or U32092 (N_32092,N_26341,N_29467);
or U32093 (N_32093,N_26440,N_29352);
xnor U32094 (N_32094,N_29433,N_25934);
nand U32095 (N_32095,N_25721,N_28650);
or U32096 (N_32096,N_25965,N_29972);
xor U32097 (N_32097,N_27227,N_28612);
nand U32098 (N_32098,N_25684,N_25393);
and U32099 (N_32099,N_29514,N_27417);
or U32100 (N_32100,N_28974,N_27226);
xnor U32101 (N_32101,N_26872,N_25079);
nand U32102 (N_32102,N_25943,N_29499);
or U32103 (N_32103,N_25209,N_28434);
xnor U32104 (N_32104,N_25394,N_28319);
and U32105 (N_32105,N_27921,N_28601);
and U32106 (N_32106,N_25173,N_26191);
nand U32107 (N_32107,N_28271,N_29004);
nand U32108 (N_32108,N_28946,N_29191);
nor U32109 (N_32109,N_27375,N_27663);
xor U32110 (N_32110,N_29046,N_27917);
nand U32111 (N_32111,N_29997,N_25021);
or U32112 (N_32112,N_25813,N_26089);
or U32113 (N_32113,N_28844,N_29671);
xnor U32114 (N_32114,N_29144,N_25217);
xor U32115 (N_32115,N_26389,N_28512);
nand U32116 (N_32116,N_26877,N_27122);
xnor U32117 (N_32117,N_27173,N_25899);
or U32118 (N_32118,N_26067,N_27807);
nand U32119 (N_32119,N_29956,N_29976);
xnor U32120 (N_32120,N_27992,N_25529);
nor U32121 (N_32121,N_27507,N_26427);
nor U32122 (N_32122,N_25602,N_28918);
nor U32123 (N_32123,N_29385,N_27342);
and U32124 (N_32124,N_27588,N_28778);
and U32125 (N_32125,N_29456,N_28163);
nor U32126 (N_32126,N_25837,N_29924);
nor U32127 (N_32127,N_25833,N_28987);
nor U32128 (N_32128,N_28588,N_29782);
and U32129 (N_32129,N_29356,N_27037);
and U32130 (N_32130,N_26792,N_29033);
and U32131 (N_32131,N_26857,N_28737);
nor U32132 (N_32132,N_29879,N_29479);
nor U32133 (N_32133,N_29726,N_27669);
nor U32134 (N_32134,N_25039,N_26064);
xnor U32135 (N_32135,N_27067,N_26834);
xor U32136 (N_32136,N_27190,N_27365);
nor U32137 (N_32137,N_27218,N_28804);
nand U32138 (N_32138,N_26286,N_26241);
or U32139 (N_32139,N_26989,N_25012);
xor U32140 (N_32140,N_26461,N_27103);
xor U32141 (N_32141,N_27584,N_28136);
and U32142 (N_32142,N_29636,N_27246);
nand U32143 (N_32143,N_26889,N_26818);
nor U32144 (N_32144,N_25996,N_27478);
or U32145 (N_32145,N_26805,N_28418);
or U32146 (N_32146,N_27586,N_29965);
nor U32147 (N_32147,N_28630,N_27248);
nor U32148 (N_32148,N_29902,N_29868);
or U32149 (N_32149,N_27631,N_27527);
xor U32150 (N_32150,N_29086,N_28498);
nor U32151 (N_32151,N_29764,N_28941);
xor U32152 (N_32152,N_28366,N_25249);
nand U32153 (N_32153,N_27931,N_27394);
xor U32154 (N_32154,N_29309,N_29622);
nand U32155 (N_32155,N_28017,N_28134);
nand U32156 (N_32156,N_28622,N_26042);
nor U32157 (N_32157,N_27200,N_25437);
nor U32158 (N_32158,N_25754,N_28305);
and U32159 (N_32159,N_29560,N_25770);
and U32160 (N_32160,N_29733,N_29948);
or U32161 (N_32161,N_29392,N_29871);
and U32162 (N_32162,N_25991,N_26778);
xnor U32163 (N_32163,N_28981,N_27042);
or U32164 (N_32164,N_28096,N_27789);
and U32165 (N_32165,N_29408,N_27363);
nand U32166 (N_32166,N_25230,N_26888);
nor U32167 (N_32167,N_26915,N_25743);
nand U32168 (N_32168,N_26713,N_29138);
nand U32169 (N_32169,N_28924,N_29021);
xor U32170 (N_32170,N_28119,N_29443);
xor U32171 (N_32171,N_26944,N_25696);
or U32172 (N_32172,N_25329,N_25520);
or U32173 (N_32173,N_27395,N_27768);
and U32174 (N_32174,N_25821,N_26560);
or U32175 (N_32175,N_29502,N_26150);
nand U32176 (N_32176,N_29845,N_26680);
xnor U32177 (N_32177,N_26157,N_28365);
nand U32178 (N_32178,N_25999,N_27714);
nand U32179 (N_32179,N_28161,N_26383);
or U32180 (N_32180,N_25612,N_26666);
nand U32181 (N_32181,N_29548,N_26132);
nor U32182 (N_32182,N_25762,N_27334);
nand U32183 (N_32183,N_27769,N_28572);
or U32184 (N_32184,N_25600,N_27231);
nand U32185 (N_32185,N_26698,N_25076);
xor U32186 (N_32186,N_27664,N_26025);
nand U32187 (N_32187,N_27111,N_28853);
nand U32188 (N_32188,N_27954,N_29200);
or U32189 (N_32189,N_27289,N_28680);
or U32190 (N_32190,N_27618,N_28644);
and U32191 (N_32191,N_26494,N_29957);
or U32192 (N_32192,N_28459,N_27662);
or U32193 (N_32193,N_25214,N_29343);
and U32194 (N_32194,N_26036,N_26703);
nor U32195 (N_32195,N_28322,N_28930);
nor U32196 (N_32196,N_28020,N_29593);
nand U32197 (N_32197,N_27784,N_25522);
xor U32198 (N_32198,N_25067,N_26806);
nand U32199 (N_32199,N_26372,N_26404);
and U32200 (N_32200,N_28817,N_29578);
nand U32201 (N_32201,N_29640,N_27164);
or U32202 (N_32202,N_28441,N_28029);
nand U32203 (N_32203,N_27093,N_28230);
xnor U32204 (N_32204,N_25023,N_25812);
xor U32205 (N_32205,N_28827,N_27385);
nor U32206 (N_32206,N_26941,N_26353);
nand U32207 (N_32207,N_29679,N_26640);
or U32208 (N_32208,N_27933,N_28285);
xor U32209 (N_32209,N_26118,N_26676);
or U32210 (N_32210,N_26158,N_28922);
or U32211 (N_32211,N_25933,N_27947);
xnor U32212 (N_32212,N_25098,N_26852);
or U32213 (N_32213,N_29114,N_29975);
nand U32214 (N_32214,N_27908,N_29162);
or U32215 (N_32215,N_28477,N_29224);
nor U32216 (N_32216,N_28694,N_29906);
and U32217 (N_32217,N_27058,N_29553);
nor U32218 (N_32218,N_25577,N_26198);
or U32219 (N_32219,N_27894,N_29490);
or U32220 (N_32220,N_25959,N_27606);
nand U32221 (N_32221,N_29744,N_25088);
xor U32222 (N_32222,N_26900,N_27559);
xor U32223 (N_32223,N_25177,N_28482);
nand U32224 (N_32224,N_26443,N_29745);
nand U32225 (N_32225,N_29817,N_25414);
and U32226 (N_32226,N_27873,N_28483);
xnor U32227 (N_32227,N_29257,N_29312);
and U32228 (N_32228,N_29861,N_25744);
and U32229 (N_32229,N_27434,N_25391);
and U32230 (N_32230,N_27924,N_26043);
nor U32231 (N_32231,N_29246,N_26978);
xnor U32232 (N_32232,N_25908,N_28739);
xor U32233 (N_32233,N_25677,N_26006);
nand U32234 (N_32234,N_25082,N_28683);
or U32235 (N_32235,N_26326,N_26589);
or U32236 (N_32236,N_28416,N_27440);
nand U32237 (N_32237,N_27644,N_27425);
and U32238 (N_32238,N_25791,N_25113);
and U32239 (N_32239,N_29178,N_25763);
nor U32240 (N_32240,N_29038,N_27597);
nand U32241 (N_32241,N_27686,N_25136);
and U32242 (N_32242,N_25279,N_28270);
nand U32243 (N_32243,N_28064,N_28598);
nor U32244 (N_32244,N_29161,N_27602);
nand U32245 (N_32245,N_29174,N_28910);
and U32246 (N_32246,N_29355,N_29226);
or U32247 (N_32247,N_28451,N_27473);
xor U32248 (N_32248,N_29728,N_29731);
xor U32249 (N_32249,N_28745,N_25779);
xor U32250 (N_32250,N_25307,N_25897);
or U32251 (N_32251,N_26476,N_27027);
and U32252 (N_32252,N_27220,N_27470);
or U32253 (N_32253,N_25613,N_27702);
or U32254 (N_32254,N_26728,N_26403);
xor U32255 (N_32255,N_25859,N_26554);
nand U32256 (N_32256,N_25698,N_27450);
nor U32257 (N_32257,N_25321,N_25295);
nand U32258 (N_32258,N_25858,N_25310);
xor U32259 (N_32259,N_26819,N_29523);
and U32260 (N_32260,N_27336,N_26981);
nand U32261 (N_32261,N_28089,N_27396);
and U32262 (N_32262,N_26773,N_29659);
or U32263 (N_32263,N_27808,N_28854);
nand U32264 (N_32264,N_29384,N_29300);
or U32265 (N_32265,N_29143,N_25731);
and U32266 (N_32266,N_26063,N_25019);
and U32267 (N_32267,N_27390,N_25856);
nand U32268 (N_32268,N_28990,N_25786);
nor U32269 (N_32269,N_25305,N_29397);
xnor U32270 (N_32270,N_29863,N_28636);
nand U32271 (N_32271,N_26733,N_28002);
or U32272 (N_32272,N_25649,N_26876);
nand U32273 (N_32273,N_27870,N_26986);
or U32274 (N_32274,N_25462,N_26214);
nor U32275 (N_32275,N_26909,N_28222);
or U32276 (N_32276,N_25759,N_26439);
xor U32277 (N_32277,N_27399,N_25336);
nor U32278 (N_32278,N_28080,N_29401);
xnor U32279 (N_32279,N_29431,N_29755);
or U32280 (N_32280,N_25272,N_28597);
xor U32281 (N_32281,N_29890,N_29157);
or U32282 (N_32282,N_29053,N_28265);
xnor U32283 (N_32283,N_27074,N_28787);
nand U32284 (N_32284,N_29314,N_27253);
xor U32285 (N_32285,N_25483,N_29266);
and U32286 (N_32286,N_27617,N_27860);
and U32287 (N_32287,N_25597,N_25093);
nor U32288 (N_32288,N_28216,N_25370);
or U32289 (N_32289,N_28106,N_25448);
nand U32290 (N_32290,N_28085,N_27488);
and U32291 (N_32291,N_26675,N_29885);
nand U32292 (N_32292,N_26034,N_29214);
and U32293 (N_32293,N_26936,N_28735);
and U32294 (N_32294,N_29942,N_26316);
or U32295 (N_32295,N_25986,N_28809);
nor U32296 (N_32296,N_25061,N_28757);
nor U32297 (N_32297,N_27751,N_27944);
or U32298 (N_32298,N_29921,N_29939);
and U32299 (N_32299,N_29633,N_28773);
or U32300 (N_32300,N_25969,N_29639);
and U32301 (N_32301,N_26500,N_26428);
nand U32302 (N_32302,N_27904,N_27300);
xor U32303 (N_32303,N_27708,N_25595);
nor U32304 (N_32304,N_29649,N_27387);
and U32305 (N_32305,N_29791,N_26515);
nor U32306 (N_32306,N_28623,N_29087);
or U32307 (N_32307,N_28391,N_25257);
xor U32308 (N_32308,N_29505,N_27418);
or U32309 (N_32309,N_29374,N_26629);
nor U32310 (N_32310,N_29148,N_28084);
xnor U32311 (N_32311,N_29862,N_25869);
or U32312 (N_32312,N_25622,N_27993);
nor U32313 (N_32313,N_28389,N_26292);
nand U32314 (N_32314,N_28765,N_25780);
nor U32315 (N_32315,N_29507,N_28313);
or U32316 (N_32316,N_26442,N_27404);
xor U32317 (N_32317,N_27832,N_29276);
or U32318 (N_32318,N_26455,N_26775);
xor U32319 (N_32319,N_27796,N_28201);
or U32320 (N_32320,N_29982,N_25657);
xnor U32321 (N_32321,N_25277,N_28112);
or U32322 (N_32322,N_26322,N_25247);
or U32323 (N_32323,N_26510,N_28940);
nor U32324 (N_32324,N_27397,N_26356);
nand U32325 (N_32325,N_26260,N_27183);
xnor U32326 (N_32326,N_29225,N_28424);
nand U32327 (N_32327,N_26078,N_27948);
nand U32328 (N_32328,N_28253,N_26918);
xnor U32329 (N_32329,N_27689,N_27977);
nand U32330 (N_32330,N_27811,N_25828);
nor U32331 (N_32331,N_28074,N_27773);
and U32332 (N_32332,N_28059,N_26323);
and U32333 (N_32333,N_25390,N_28166);
nand U32334 (N_32334,N_27057,N_27771);
or U32335 (N_32335,N_27316,N_28648);
nor U32336 (N_32336,N_26144,N_28890);
xor U32337 (N_32337,N_29477,N_27062);
xnor U32338 (N_32338,N_26269,N_27040);
or U32339 (N_32339,N_29534,N_25720);
xor U32340 (N_32340,N_28833,N_26275);
nand U32341 (N_32341,N_29255,N_29367);
nand U32342 (N_32342,N_25340,N_25687);
nor U32343 (N_32343,N_26082,N_28054);
nor U32344 (N_32344,N_27211,N_26522);
or U32345 (N_32345,N_25451,N_27468);
nand U32346 (N_32346,N_29422,N_27650);
xor U32347 (N_32347,N_26072,N_26313);
nor U32348 (N_32348,N_29054,N_26052);
nand U32349 (N_32349,N_26934,N_27780);
nor U32350 (N_32350,N_28405,N_26516);
nor U32351 (N_32351,N_26084,N_27485);
and U32352 (N_32352,N_29800,N_28019);
or U32353 (N_32353,N_27377,N_27535);
xor U32354 (N_32354,N_28295,N_26279);
nor U32355 (N_32355,N_25753,N_28549);
xor U32356 (N_32356,N_29102,N_27998);
and U32357 (N_32357,N_29001,N_27323);
or U32358 (N_32358,N_28664,N_25456);
or U32359 (N_32359,N_27756,N_29248);
nor U32360 (N_32360,N_29175,N_27685);
nor U32361 (N_32361,N_28478,N_25438);
nor U32362 (N_32362,N_25137,N_27958);
nor U32363 (N_32363,N_25697,N_25396);
nor U32364 (N_32364,N_26658,N_28445);
xor U32365 (N_32365,N_27743,N_27658);
and U32366 (N_32366,N_26663,N_27522);
nor U32367 (N_32367,N_28772,N_27596);
nor U32368 (N_32368,N_25232,N_29993);
xor U32369 (N_32369,N_27477,N_29049);
xor U32370 (N_32370,N_29859,N_28487);
nor U32371 (N_32371,N_26029,N_26633);
xor U32372 (N_32372,N_25734,N_26367);
xnor U32373 (N_32373,N_27699,N_29775);
nand U32374 (N_32374,N_27312,N_26730);
nand U32375 (N_32375,N_26435,N_27138);
nand U32376 (N_32376,N_27560,N_25142);
and U32377 (N_32377,N_25327,N_27646);
and U32378 (N_32378,N_27830,N_26334);
or U32379 (N_32379,N_27155,N_29839);
and U32380 (N_32380,N_26545,N_28693);
nand U32381 (N_32381,N_25551,N_27680);
xnor U32382 (N_32382,N_27718,N_28367);
xnor U32383 (N_32383,N_29323,N_25910);
nand U32384 (N_32384,N_29777,N_26473);
and U32385 (N_32385,N_29836,N_28750);
or U32386 (N_32386,N_27734,N_25179);
nor U32387 (N_32387,N_28722,N_26800);
xnor U32388 (N_32388,N_28894,N_25001);
or U32389 (N_32389,N_29168,N_26085);
nor U32390 (N_32390,N_26785,N_27772);
and U32391 (N_32391,N_28646,N_28937);
and U32392 (N_32392,N_28651,N_26328);
xor U32393 (N_32393,N_28629,N_28375);
nand U32394 (N_32394,N_29229,N_25242);
xnor U32395 (N_32395,N_28197,N_29758);
or U32396 (N_32396,N_26338,N_28118);
nand U32397 (N_32397,N_28290,N_29766);
or U32398 (N_32398,N_28916,N_26551);
and U32399 (N_32399,N_26490,N_25523);
or U32400 (N_32400,N_25096,N_26543);
xnor U32401 (N_32401,N_29347,N_29289);
xnor U32402 (N_32402,N_27009,N_27491);
or U32403 (N_32403,N_29704,N_29925);
and U32404 (N_32404,N_27079,N_26983);
or U32405 (N_32405,N_27495,N_28523);
or U32406 (N_32406,N_26358,N_29789);
nand U32407 (N_32407,N_29445,N_26993);
nand U32408 (N_32408,N_29732,N_25195);
nor U32409 (N_32409,N_27298,N_29328);
xor U32410 (N_32410,N_26735,N_28213);
nand U32411 (N_32411,N_28767,N_25312);
and U32412 (N_32412,N_25547,N_26371);
xor U32413 (N_32413,N_27591,N_28799);
nor U32414 (N_32414,N_25274,N_26644);
and U32415 (N_32415,N_27563,N_29586);
or U32416 (N_32416,N_26846,N_29887);
nor U32417 (N_32417,N_25726,N_28710);
nor U32418 (N_32418,N_29142,N_28897);
xor U32419 (N_32419,N_26019,N_28035);
nand U32420 (N_32420,N_28982,N_25198);
nand U32421 (N_32421,N_29448,N_26412);
nor U32422 (N_32422,N_26744,N_27941);
nor U32423 (N_32423,N_26726,N_28260);
nand U32424 (N_32424,N_27221,N_29927);
nand U32425 (N_32425,N_25344,N_28192);
nor U32426 (N_32426,N_27845,N_25263);
xnor U32427 (N_32427,N_27988,N_26814);
nor U32428 (N_32428,N_27276,N_27077);
and U32429 (N_32429,N_26798,N_28153);
nand U32430 (N_32430,N_27816,N_26781);
and U32431 (N_32431,N_29645,N_29044);
nor U32432 (N_32432,N_25556,N_25358);
or U32433 (N_32433,N_29109,N_28352);
xnor U32434 (N_32434,N_27723,N_27171);
or U32435 (N_32435,N_25977,N_29609);
nand U32436 (N_32436,N_27329,N_25243);
nand U32437 (N_32437,N_28994,N_27234);
nand U32438 (N_32438,N_27974,N_25156);
xnor U32439 (N_32439,N_26887,N_28713);
xnor U32440 (N_32440,N_29055,N_27360);
xnor U32441 (N_32441,N_26126,N_27616);
nor U32442 (N_32442,N_29121,N_27038);
and U32443 (N_32443,N_28506,N_26054);
nand U32444 (N_32444,N_28242,N_25072);
nand U32445 (N_32445,N_28992,N_25685);
nand U32446 (N_32446,N_25402,N_26103);
or U32447 (N_32447,N_25747,N_25090);
nor U32448 (N_32448,N_27639,N_28566);
and U32449 (N_32449,N_26669,N_29107);
nor U32450 (N_32450,N_29937,N_25953);
or U32451 (N_32451,N_26759,N_25311);
or U32452 (N_32452,N_27795,N_27106);
and U32453 (N_32453,N_28348,N_26974);
or U32454 (N_32454,N_26321,N_28500);
nor U32455 (N_32455,N_26272,N_29511);
xnor U32456 (N_32456,N_28388,N_28053);
or U32457 (N_32457,N_25374,N_25107);
or U32458 (N_32458,N_28889,N_27583);
nor U32459 (N_32459,N_29113,N_29164);
nand U32460 (N_32460,N_28399,N_29441);
xnor U32461 (N_32461,N_26066,N_25184);
and U32462 (N_32462,N_26931,N_25796);
nor U32463 (N_32463,N_29709,N_26352);
or U32464 (N_32464,N_26642,N_28908);
xnor U32465 (N_32465,N_26505,N_26858);
or U32466 (N_32466,N_29673,N_28514);
and U32467 (N_32467,N_25125,N_25951);
and U32468 (N_32468,N_26970,N_29334);
or U32469 (N_32469,N_25949,N_29052);
nor U32470 (N_32470,N_29856,N_26197);
nand U32471 (N_32471,N_25662,N_25576);
nand U32472 (N_32472,N_29851,N_27154);
nor U32473 (N_32473,N_26242,N_28256);
nand U32474 (N_32474,N_27783,N_29739);
or U32475 (N_32475,N_25218,N_27971);
xor U32476 (N_32476,N_29540,N_26809);
and U32477 (N_32477,N_26017,N_26613);
nand U32478 (N_32478,N_28479,N_27854);
nand U32479 (N_32479,N_26413,N_26940);
nor U32480 (N_32480,N_25849,N_28289);
nor U32481 (N_32481,N_27976,N_26539);
or U32482 (N_32482,N_29779,N_25741);
nand U32483 (N_32483,N_28534,N_28747);
and U32484 (N_32484,N_25297,N_27119);
or U32485 (N_32485,N_29978,N_26664);
and U32486 (N_32486,N_25621,N_25809);
or U32487 (N_32487,N_29711,N_27722);
and U32488 (N_32488,N_27700,N_28098);
or U32489 (N_32489,N_29929,N_27277);
or U32490 (N_32490,N_29061,N_28796);
nor U32491 (N_32491,N_26331,N_27812);
nor U32492 (N_32492,N_29796,N_28979);
xnor U32493 (N_32493,N_25690,N_26849);
nor U32494 (N_32494,N_27798,N_29646);
or U32495 (N_32495,N_28380,N_27427);
and U32496 (N_32496,N_29216,N_26415);
nor U32497 (N_32497,N_26492,N_25182);
nand U32498 (N_32498,N_26493,N_29944);
and U32499 (N_32499,N_29596,N_29881);
nor U32500 (N_32500,N_29866,N_27630);
or U32501 (N_32501,N_25261,N_25458);
and U32502 (N_32502,N_28590,N_27894);
nand U32503 (N_32503,N_29067,N_26593);
nor U32504 (N_32504,N_26921,N_25933);
nand U32505 (N_32505,N_25829,N_27663);
xor U32506 (N_32506,N_26481,N_29647);
nand U32507 (N_32507,N_28791,N_25562);
or U32508 (N_32508,N_25609,N_29984);
or U32509 (N_32509,N_29202,N_27086);
and U32510 (N_32510,N_27650,N_26642);
or U32511 (N_32511,N_28471,N_27352);
xnor U32512 (N_32512,N_26137,N_25192);
nand U32513 (N_32513,N_25901,N_28866);
nand U32514 (N_32514,N_25442,N_28045);
or U32515 (N_32515,N_29442,N_25568);
and U32516 (N_32516,N_26071,N_28299);
nand U32517 (N_32517,N_29473,N_26284);
nand U32518 (N_32518,N_29223,N_29662);
nor U32519 (N_32519,N_28274,N_26308);
nand U32520 (N_32520,N_29049,N_29176);
or U32521 (N_32521,N_29966,N_26236);
and U32522 (N_32522,N_26775,N_28503);
xor U32523 (N_32523,N_25490,N_29161);
or U32524 (N_32524,N_28625,N_26604);
nor U32525 (N_32525,N_27789,N_27947);
and U32526 (N_32526,N_27663,N_26424);
nor U32527 (N_32527,N_28151,N_26351);
nand U32528 (N_32528,N_26000,N_26134);
or U32529 (N_32529,N_28024,N_26808);
and U32530 (N_32530,N_28390,N_26374);
nor U32531 (N_32531,N_28318,N_29782);
and U32532 (N_32532,N_27050,N_27102);
xor U32533 (N_32533,N_26112,N_28122);
or U32534 (N_32534,N_25611,N_26276);
nand U32535 (N_32535,N_27305,N_25729);
xor U32536 (N_32536,N_28230,N_28256);
and U32537 (N_32537,N_27908,N_28440);
xnor U32538 (N_32538,N_26634,N_25438);
nor U32539 (N_32539,N_27502,N_27044);
nand U32540 (N_32540,N_26641,N_28645);
or U32541 (N_32541,N_25922,N_28326);
nor U32542 (N_32542,N_25522,N_27653);
and U32543 (N_32543,N_26823,N_27884);
xnor U32544 (N_32544,N_28074,N_29285);
and U32545 (N_32545,N_28366,N_28575);
and U32546 (N_32546,N_26183,N_26510);
or U32547 (N_32547,N_27276,N_29662);
or U32548 (N_32548,N_25179,N_27264);
and U32549 (N_32549,N_27679,N_26040);
xor U32550 (N_32550,N_25595,N_27618);
nand U32551 (N_32551,N_29619,N_27886);
xor U32552 (N_32552,N_27208,N_27717);
nand U32553 (N_32553,N_27205,N_29633);
and U32554 (N_32554,N_29511,N_28014);
or U32555 (N_32555,N_28963,N_25820);
or U32556 (N_32556,N_25090,N_27534);
nand U32557 (N_32557,N_26899,N_28469);
and U32558 (N_32558,N_28318,N_28473);
nand U32559 (N_32559,N_26059,N_26904);
nor U32560 (N_32560,N_26544,N_28307);
or U32561 (N_32561,N_26755,N_26671);
nor U32562 (N_32562,N_28459,N_26630);
xnor U32563 (N_32563,N_27776,N_25583);
or U32564 (N_32564,N_27491,N_26341);
xnor U32565 (N_32565,N_26417,N_26620);
or U32566 (N_32566,N_28689,N_29216);
nor U32567 (N_32567,N_28034,N_27940);
and U32568 (N_32568,N_29695,N_29256);
xor U32569 (N_32569,N_26957,N_28785);
nand U32570 (N_32570,N_25917,N_27635);
xnor U32571 (N_32571,N_25793,N_29342);
nor U32572 (N_32572,N_28422,N_29559);
xor U32573 (N_32573,N_28981,N_25390);
or U32574 (N_32574,N_27838,N_26880);
or U32575 (N_32575,N_28065,N_26630);
and U32576 (N_32576,N_25467,N_25797);
and U32577 (N_32577,N_25929,N_28263);
nand U32578 (N_32578,N_26581,N_26148);
and U32579 (N_32579,N_29679,N_27675);
nor U32580 (N_32580,N_26525,N_25412);
xnor U32581 (N_32581,N_26787,N_26410);
or U32582 (N_32582,N_29917,N_27998);
nand U32583 (N_32583,N_29433,N_25417);
or U32584 (N_32584,N_29676,N_28827);
nand U32585 (N_32585,N_27775,N_25608);
nand U32586 (N_32586,N_28300,N_25050);
nand U32587 (N_32587,N_27036,N_27498);
nor U32588 (N_32588,N_28166,N_29574);
and U32589 (N_32589,N_28222,N_27061);
nand U32590 (N_32590,N_26534,N_27942);
and U32591 (N_32591,N_25165,N_28514);
and U32592 (N_32592,N_26150,N_28751);
or U32593 (N_32593,N_25496,N_27413);
xnor U32594 (N_32594,N_25634,N_26889);
or U32595 (N_32595,N_26989,N_29555);
and U32596 (N_32596,N_27235,N_25526);
or U32597 (N_32597,N_29495,N_26599);
xor U32598 (N_32598,N_29993,N_25177);
and U32599 (N_32599,N_29156,N_27596);
or U32600 (N_32600,N_26694,N_28592);
or U32601 (N_32601,N_27730,N_25555);
nand U32602 (N_32602,N_26508,N_27271);
nor U32603 (N_32603,N_29655,N_25086);
nor U32604 (N_32604,N_27138,N_26571);
and U32605 (N_32605,N_29183,N_28696);
xor U32606 (N_32606,N_26644,N_29641);
nor U32607 (N_32607,N_26475,N_26178);
xor U32608 (N_32608,N_28109,N_29120);
and U32609 (N_32609,N_27328,N_28630);
and U32610 (N_32610,N_26942,N_28270);
xnor U32611 (N_32611,N_28127,N_28835);
and U32612 (N_32612,N_25455,N_26462);
nor U32613 (N_32613,N_28800,N_26542);
nand U32614 (N_32614,N_26358,N_29182);
or U32615 (N_32615,N_29397,N_29983);
and U32616 (N_32616,N_26987,N_27939);
xnor U32617 (N_32617,N_25377,N_26256);
nand U32618 (N_32618,N_25452,N_28792);
xor U32619 (N_32619,N_27316,N_28072);
xnor U32620 (N_32620,N_26619,N_25814);
nand U32621 (N_32621,N_26470,N_25872);
xnor U32622 (N_32622,N_28763,N_27649);
or U32623 (N_32623,N_28091,N_28474);
or U32624 (N_32624,N_27725,N_26496);
and U32625 (N_32625,N_26063,N_25751);
nand U32626 (N_32626,N_28182,N_25823);
xnor U32627 (N_32627,N_27213,N_26384);
or U32628 (N_32628,N_25907,N_26826);
xor U32629 (N_32629,N_28095,N_26122);
xnor U32630 (N_32630,N_27984,N_28267);
nor U32631 (N_32631,N_29633,N_27882);
and U32632 (N_32632,N_28681,N_29019);
and U32633 (N_32633,N_26190,N_28293);
and U32634 (N_32634,N_28132,N_28794);
xnor U32635 (N_32635,N_29541,N_25906);
nor U32636 (N_32636,N_26138,N_26453);
nand U32637 (N_32637,N_26321,N_26156);
and U32638 (N_32638,N_26336,N_25803);
or U32639 (N_32639,N_27820,N_29514);
or U32640 (N_32640,N_28602,N_26002);
nor U32641 (N_32641,N_29964,N_28203);
xnor U32642 (N_32642,N_26095,N_25120);
or U32643 (N_32643,N_28335,N_27672);
and U32644 (N_32644,N_25703,N_27097);
xnor U32645 (N_32645,N_27398,N_28257);
xor U32646 (N_32646,N_26850,N_25233);
and U32647 (N_32647,N_28225,N_27518);
or U32648 (N_32648,N_28031,N_25307);
or U32649 (N_32649,N_27383,N_27534);
xor U32650 (N_32650,N_25205,N_25826);
xnor U32651 (N_32651,N_25885,N_29736);
or U32652 (N_32652,N_29005,N_25599);
nand U32653 (N_32653,N_28540,N_25029);
and U32654 (N_32654,N_29973,N_29671);
nand U32655 (N_32655,N_27869,N_29177);
and U32656 (N_32656,N_28732,N_29207);
xor U32657 (N_32657,N_29911,N_25149);
and U32658 (N_32658,N_29004,N_25454);
nand U32659 (N_32659,N_26313,N_27822);
and U32660 (N_32660,N_28472,N_28931);
xor U32661 (N_32661,N_27139,N_27331);
and U32662 (N_32662,N_29485,N_26342);
nand U32663 (N_32663,N_29160,N_27614);
nand U32664 (N_32664,N_29640,N_29603);
nor U32665 (N_32665,N_29498,N_26813);
xnor U32666 (N_32666,N_25651,N_28519);
or U32667 (N_32667,N_25889,N_27166);
and U32668 (N_32668,N_28264,N_28020);
or U32669 (N_32669,N_28671,N_27365);
nand U32670 (N_32670,N_29137,N_29498);
nand U32671 (N_32671,N_26155,N_28944);
nand U32672 (N_32672,N_28926,N_26264);
xor U32673 (N_32673,N_28454,N_27282);
or U32674 (N_32674,N_27296,N_26354);
xor U32675 (N_32675,N_28169,N_26048);
nand U32676 (N_32676,N_26046,N_26708);
nand U32677 (N_32677,N_29438,N_28957);
nand U32678 (N_32678,N_29346,N_27940);
nor U32679 (N_32679,N_28448,N_25676);
xor U32680 (N_32680,N_27959,N_29096);
and U32681 (N_32681,N_26270,N_27154);
nand U32682 (N_32682,N_27365,N_25897);
or U32683 (N_32683,N_27276,N_28159);
and U32684 (N_32684,N_25517,N_29158);
nor U32685 (N_32685,N_25155,N_29531);
and U32686 (N_32686,N_25483,N_29714);
and U32687 (N_32687,N_28898,N_26259);
nand U32688 (N_32688,N_28738,N_28866);
xnor U32689 (N_32689,N_27669,N_26337);
and U32690 (N_32690,N_28386,N_29039);
nor U32691 (N_32691,N_28860,N_26338);
nand U32692 (N_32692,N_25851,N_26234);
nor U32693 (N_32693,N_25977,N_25749);
nor U32694 (N_32694,N_28616,N_25433);
or U32695 (N_32695,N_29570,N_29964);
nand U32696 (N_32696,N_25738,N_25806);
nor U32697 (N_32697,N_29741,N_26494);
xnor U32698 (N_32698,N_26919,N_28235);
or U32699 (N_32699,N_27862,N_25940);
nand U32700 (N_32700,N_28792,N_26959);
nor U32701 (N_32701,N_28124,N_25505);
xnor U32702 (N_32702,N_29282,N_28894);
and U32703 (N_32703,N_25161,N_25243);
or U32704 (N_32704,N_26985,N_29307);
xor U32705 (N_32705,N_27195,N_26208);
and U32706 (N_32706,N_29265,N_25294);
and U32707 (N_32707,N_28141,N_25270);
nor U32708 (N_32708,N_29260,N_25525);
or U32709 (N_32709,N_27016,N_29705);
or U32710 (N_32710,N_25598,N_28755);
or U32711 (N_32711,N_28001,N_27787);
xnor U32712 (N_32712,N_28629,N_25885);
or U32713 (N_32713,N_26551,N_25697);
and U32714 (N_32714,N_27536,N_27406);
or U32715 (N_32715,N_25983,N_25383);
nor U32716 (N_32716,N_29892,N_28262);
nand U32717 (N_32717,N_26783,N_25065);
and U32718 (N_32718,N_29257,N_27371);
or U32719 (N_32719,N_25941,N_26534);
and U32720 (N_32720,N_25678,N_27597);
and U32721 (N_32721,N_26331,N_27581);
xor U32722 (N_32722,N_26444,N_29530);
nor U32723 (N_32723,N_27040,N_26402);
and U32724 (N_32724,N_28505,N_26276);
or U32725 (N_32725,N_29456,N_27137);
and U32726 (N_32726,N_26880,N_29352);
nor U32727 (N_32727,N_25092,N_26308);
and U32728 (N_32728,N_26034,N_27068);
nand U32729 (N_32729,N_28556,N_29795);
xnor U32730 (N_32730,N_25059,N_26639);
or U32731 (N_32731,N_26870,N_28792);
nor U32732 (N_32732,N_27495,N_29077);
or U32733 (N_32733,N_28562,N_29750);
nand U32734 (N_32734,N_28290,N_26903);
and U32735 (N_32735,N_25317,N_27986);
or U32736 (N_32736,N_29705,N_28867);
xnor U32737 (N_32737,N_28166,N_29916);
nand U32738 (N_32738,N_27875,N_25674);
xnor U32739 (N_32739,N_25136,N_27389);
and U32740 (N_32740,N_26983,N_27734);
nor U32741 (N_32741,N_25713,N_28190);
xor U32742 (N_32742,N_28454,N_27934);
nand U32743 (N_32743,N_26013,N_29964);
xor U32744 (N_32744,N_27193,N_26683);
or U32745 (N_32745,N_26465,N_29048);
or U32746 (N_32746,N_27813,N_28141);
nand U32747 (N_32747,N_26333,N_26884);
or U32748 (N_32748,N_27819,N_27707);
xnor U32749 (N_32749,N_25450,N_29211);
nor U32750 (N_32750,N_29558,N_29081);
nand U32751 (N_32751,N_26581,N_26284);
nor U32752 (N_32752,N_27289,N_26684);
or U32753 (N_32753,N_28551,N_29614);
xor U32754 (N_32754,N_28634,N_28438);
and U32755 (N_32755,N_28085,N_28332);
nor U32756 (N_32756,N_26148,N_26098);
nand U32757 (N_32757,N_25271,N_29348);
xor U32758 (N_32758,N_29105,N_28820);
nand U32759 (N_32759,N_26671,N_29792);
nand U32760 (N_32760,N_25439,N_27613);
xnor U32761 (N_32761,N_27147,N_29449);
or U32762 (N_32762,N_25168,N_28478);
and U32763 (N_32763,N_29956,N_25393);
nor U32764 (N_32764,N_28007,N_25407);
and U32765 (N_32765,N_25254,N_25115);
nand U32766 (N_32766,N_29236,N_26293);
xnor U32767 (N_32767,N_27394,N_25277);
xnor U32768 (N_32768,N_27846,N_25310);
nand U32769 (N_32769,N_28913,N_26395);
xor U32770 (N_32770,N_29129,N_25832);
nor U32771 (N_32771,N_28572,N_25952);
nand U32772 (N_32772,N_25897,N_25900);
and U32773 (N_32773,N_29960,N_27129);
or U32774 (N_32774,N_28747,N_29044);
and U32775 (N_32775,N_28531,N_26163);
nor U32776 (N_32776,N_26745,N_25523);
nand U32777 (N_32777,N_28816,N_27146);
nor U32778 (N_32778,N_27480,N_28458);
and U32779 (N_32779,N_29058,N_25255);
nand U32780 (N_32780,N_28845,N_25321);
nor U32781 (N_32781,N_25320,N_26588);
or U32782 (N_32782,N_28803,N_27242);
and U32783 (N_32783,N_28145,N_27801);
or U32784 (N_32784,N_29675,N_29159);
and U32785 (N_32785,N_29924,N_25698);
and U32786 (N_32786,N_26971,N_27183);
xor U32787 (N_32787,N_25886,N_25505);
or U32788 (N_32788,N_29948,N_28706);
xor U32789 (N_32789,N_25443,N_25546);
or U32790 (N_32790,N_26472,N_26614);
and U32791 (N_32791,N_28506,N_26439);
and U32792 (N_32792,N_25324,N_25824);
or U32793 (N_32793,N_27137,N_25885);
and U32794 (N_32794,N_29792,N_26843);
or U32795 (N_32795,N_25678,N_25832);
nand U32796 (N_32796,N_26336,N_28460);
nor U32797 (N_32797,N_25016,N_29801);
xor U32798 (N_32798,N_26303,N_25758);
and U32799 (N_32799,N_25696,N_25636);
xor U32800 (N_32800,N_27778,N_26165);
and U32801 (N_32801,N_29449,N_27843);
nand U32802 (N_32802,N_27512,N_26677);
nor U32803 (N_32803,N_26587,N_26602);
nor U32804 (N_32804,N_26293,N_25192);
and U32805 (N_32805,N_26436,N_27201);
nand U32806 (N_32806,N_26169,N_26850);
or U32807 (N_32807,N_28877,N_27129);
xor U32808 (N_32808,N_26159,N_28961);
nor U32809 (N_32809,N_27419,N_27739);
or U32810 (N_32810,N_28348,N_25945);
or U32811 (N_32811,N_27544,N_27740);
and U32812 (N_32812,N_28196,N_29355);
and U32813 (N_32813,N_28932,N_29334);
and U32814 (N_32814,N_26743,N_29006);
or U32815 (N_32815,N_25209,N_25189);
xor U32816 (N_32816,N_27073,N_27757);
nor U32817 (N_32817,N_26117,N_28562);
nor U32818 (N_32818,N_28762,N_28298);
nor U32819 (N_32819,N_26435,N_26184);
and U32820 (N_32820,N_25303,N_25254);
and U32821 (N_32821,N_26174,N_27928);
nand U32822 (N_32822,N_27897,N_29251);
or U32823 (N_32823,N_25108,N_27824);
nor U32824 (N_32824,N_29502,N_26650);
or U32825 (N_32825,N_28533,N_27721);
and U32826 (N_32826,N_27532,N_29915);
nand U32827 (N_32827,N_26300,N_28230);
nor U32828 (N_32828,N_26564,N_29815);
nand U32829 (N_32829,N_29388,N_29350);
or U32830 (N_32830,N_26772,N_28487);
nor U32831 (N_32831,N_25156,N_26825);
nor U32832 (N_32832,N_29543,N_28161);
nor U32833 (N_32833,N_26946,N_27466);
nor U32834 (N_32834,N_28475,N_25624);
xnor U32835 (N_32835,N_25829,N_29098);
or U32836 (N_32836,N_28435,N_25716);
nor U32837 (N_32837,N_28643,N_27259);
nor U32838 (N_32838,N_26855,N_25092);
and U32839 (N_32839,N_25429,N_26214);
nand U32840 (N_32840,N_26700,N_27975);
and U32841 (N_32841,N_27461,N_25068);
xnor U32842 (N_32842,N_25493,N_25204);
xnor U32843 (N_32843,N_27727,N_27676);
nor U32844 (N_32844,N_29032,N_25522);
and U32845 (N_32845,N_27922,N_29791);
or U32846 (N_32846,N_26820,N_29927);
xnor U32847 (N_32847,N_29635,N_25976);
or U32848 (N_32848,N_28244,N_29867);
or U32849 (N_32849,N_29296,N_26684);
nand U32850 (N_32850,N_25519,N_25815);
and U32851 (N_32851,N_29870,N_25712);
xnor U32852 (N_32852,N_26362,N_29763);
xor U32853 (N_32853,N_29066,N_25411);
or U32854 (N_32854,N_27149,N_27881);
nor U32855 (N_32855,N_27068,N_26922);
nand U32856 (N_32856,N_26728,N_28425);
and U32857 (N_32857,N_27152,N_29435);
xor U32858 (N_32858,N_25197,N_28373);
nor U32859 (N_32859,N_25246,N_27400);
nand U32860 (N_32860,N_27320,N_28477);
and U32861 (N_32861,N_26552,N_28340);
nand U32862 (N_32862,N_28062,N_25414);
nand U32863 (N_32863,N_27971,N_29851);
and U32864 (N_32864,N_28862,N_27566);
nor U32865 (N_32865,N_26132,N_26302);
and U32866 (N_32866,N_28928,N_29046);
nor U32867 (N_32867,N_26999,N_28658);
or U32868 (N_32868,N_27423,N_26126);
nand U32869 (N_32869,N_25556,N_25456);
xor U32870 (N_32870,N_27242,N_26299);
or U32871 (N_32871,N_27306,N_29051);
nand U32872 (N_32872,N_26062,N_28965);
xor U32873 (N_32873,N_27710,N_26921);
nor U32874 (N_32874,N_27605,N_26348);
nand U32875 (N_32875,N_29874,N_26874);
and U32876 (N_32876,N_29888,N_25754);
xnor U32877 (N_32877,N_26427,N_26452);
nand U32878 (N_32878,N_28638,N_25477);
or U32879 (N_32879,N_25604,N_26081);
xor U32880 (N_32880,N_25450,N_26889);
nand U32881 (N_32881,N_25255,N_29505);
xnor U32882 (N_32882,N_28829,N_28285);
nand U32883 (N_32883,N_25229,N_25333);
and U32884 (N_32884,N_27807,N_27788);
xnor U32885 (N_32885,N_25280,N_27979);
nand U32886 (N_32886,N_26659,N_28302);
nand U32887 (N_32887,N_29676,N_25417);
nand U32888 (N_32888,N_28783,N_26297);
nor U32889 (N_32889,N_25116,N_27947);
nor U32890 (N_32890,N_27440,N_29561);
and U32891 (N_32891,N_27747,N_27577);
xnor U32892 (N_32892,N_28674,N_28512);
and U32893 (N_32893,N_25760,N_26818);
xnor U32894 (N_32894,N_25828,N_29979);
and U32895 (N_32895,N_28999,N_27160);
or U32896 (N_32896,N_28104,N_25108);
and U32897 (N_32897,N_28460,N_26742);
xor U32898 (N_32898,N_25303,N_27888);
xor U32899 (N_32899,N_29282,N_25333);
nor U32900 (N_32900,N_28177,N_25063);
xnor U32901 (N_32901,N_26975,N_27677);
or U32902 (N_32902,N_26581,N_28403);
xor U32903 (N_32903,N_25566,N_29903);
nand U32904 (N_32904,N_25984,N_29345);
or U32905 (N_32905,N_29503,N_27581);
or U32906 (N_32906,N_29200,N_25626);
or U32907 (N_32907,N_26888,N_25602);
xnor U32908 (N_32908,N_28350,N_28289);
or U32909 (N_32909,N_25775,N_26810);
xor U32910 (N_32910,N_28981,N_26937);
or U32911 (N_32911,N_29629,N_29469);
or U32912 (N_32912,N_26498,N_29569);
xor U32913 (N_32913,N_29704,N_28866);
or U32914 (N_32914,N_27115,N_27479);
and U32915 (N_32915,N_26733,N_25202);
or U32916 (N_32916,N_29278,N_29042);
and U32917 (N_32917,N_28278,N_25367);
nand U32918 (N_32918,N_29816,N_29643);
nor U32919 (N_32919,N_28988,N_26835);
nor U32920 (N_32920,N_26072,N_25336);
and U32921 (N_32921,N_28026,N_28418);
and U32922 (N_32922,N_29781,N_27172);
nor U32923 (N_32923,N_26423,N_26289);
and U32924 (N_32924,N_27249,N_29372);
xnor U32925 (N_32925,N_25023,N_28443);
xnor U32926 (N_32926,N_28658,N_27064);
nor U32927 (N_32927,N_26596,N_27327);
xor U32928 (N_32928,N_29896,N_25236);
or U32929 (N_32929,N_28752,N_29718);
nor U32930 (N_32930,N_27778,N_25515);
nand U32931 (N_32931,N_25720,N_26776);
xnor U32932 (N_32932,N_26913,N_27961);
nand U32933 (N_32933,N_29839,N_29356);
xor U32934 (N_32934,N_28028,N_25569);
and U32935 (N_32935,N_25071,N_26866);
nand U32936 (N_32936,N_25789,N_29456);
and U32937 (N_32937,N_29302,N_25692);
nand U32938 (N_32938,N_29365,N_29750);
and U32939 (N_32939,N_29848,N_28461);
nor U32940 (N_32940,N_27016,N_25396);
or U32941 (N_32941,N_28249,N_25089);
xor U32942 (N_32942,N_28379,N_26754);
or U32943 (N_32943,N_26422,N_28782);
nand U32944 (N_32944,N_28315,N_28747);
or U32945 (N_32945,N_26483,N_26462);
nand U32946 (N_32946,N_29156,N_28519);
or U32947 (N_32947,N_26418,N_29196);
xnor U32948 (N_32948,N_27513,N_29284);
and U32949 (N_32949,N_25231,N_26606);
nor U32950 (N_32950,N_25208,N_26295);
nand U32951 (N_32951,N_26051,N_26877);
xnor U32952 (N_32952,N_29754,N_26879);
nor U32953 (N_32953,N_27745,N_28019);
xor U32954 (N_32954,N_26893,N_29987);
nor U32955 (N_32955,N_25364,N_29538);
and U32956 (N_32956,N_29101,N_27819);
and U32957 (N_32957,N_26077,N_25509);
nor U32958 (N_32958,N_28312,N_25294);
xnor U32959 (N_32959,N_26430,N_26047);
nand U32960 (N_32960,N_26861,N_27235);
and U32961 (N_32961,N_28352,N_25019);
nand U32962 (N_32962,N_29946,N_26579);
nor U32963 (N_32963,N_29993,N_29516);
xor U32964 (N_32964,N_26809,N_29853);
xnor U32965 (N_32965,N_29644,N_28056);
xnor U32966 (N_32966,N_29078,N_26464);
xor U32967 (N_32967,N_28636,N_25807);
and U32968 (N_32968,N_26958,N_26489);
nor U32969 (N_32969,N_29527,N_29528);
nand U32970 (N_32970,N_29883,N_29344);
and U32971 (N_32971,N_27058,N_27383);
nand U32972 (N_32972,N_27532,N_28131);
and U32973 (N_32973,N_29165,N_27746);
nand U32974 (N_32974,N_28302,N_28942);
nor U32975 (N_32975,N_28524,N_29588);
nand U32976 (N_32976,N_25624,N_28634);
and U32977 (N_32977,N_25176,N_26754);
and U32978 (N_32978,N_28844,N_29194);
nand U32979 (N_32979,N_29198,N_27379);
and U32980 (N_32980,N_27286,N_29869);
xor U32981 (N_32981,N_29543,N_27660);
xor U32982 (N_32982,N_27481,N_27164);
nor U32983 (N_32983,N_28974,N_28847);
xnor U32984 (N_32984,N_26692,N_25659);
nor U32985 (N_32985,N_29582,N_28433);
xnor U32986 (N_32986,N_27931,N_29763);
nand U32987 (N_32987,N_28554,N_26339);
and U32988 (N_32988,N_28868,N_27511);
nand U32989 (N_32989,N_25888,N_26136);
nand U32990 (N_32990,N_28911,N_27194);
xor U32991 (N_32991,N_25700,N_27502);
nor U32992 (N_32992,N_27419,N_27348);
or U32993 (N_32993,N_28718,N_29547);
nand U32994 (N_32994,N_25947,N_28628);
xor U32995 (N_32995,N_28765,N_28488);
and U32996 (N_32996,N_27886,N_26755);
and U32997 (N_32997,N_29595,N_27084);
or U32998 (N_32998,N_28517,N_26148);
xor U32999 (N_32999,N_27201,N_29414);
nor U33000 (N_33000,N_28836,N_26256);
xnor U33001 (N_33001,N_28385,N_29924);
nor U33002 (N_33002,N_25096,N_29844);
nor U33003 (N_33003,N_25546,N_29089);
or U33004 (N_33004,N_25521,N_26035);
and U33005 (N_33005,N_25964,N_27214);
nor U33006 (N_33006,N_29049,N_27294);
or U33007 (N_33007,N_26872,N_25962);
nand U33008 (N_33008,N_28630,N_26834);
nor U33009 (N_33009,N_26707,N_26834);
or U33010 (N_33010,N_29788,N_26629);
or U33011 (N_33011,N_28911,N_25559);
xnor U33012 (N_33012,N_26870,N_28706);
and U33013 (N_33013,N_25282,N_25460);
or U33014 (N_33014,N_25923,N_27360);
nand U33015 (N_33015,N_27305,N_26236);
nor U33016 (N_33016,N_29513,N_26415);
nand U33017 (N_33017,N_29804,N_25811);
or U33018 (N_33018,N_26554,N_25672);
nor U33019 (N_33019,N_25118,N_25138);
nand U33020 (N_33020,N_29300,N_27406);
or U33021 (N_33021,N_29691,N_25862);
nand U33022 (N_33022,N_29880,N_28832);
or U33023 (N_33023,N_27545,N_25048);
nand U33024 (N_33024,N_29375,N_25062);
xor U33025 (N_33025,N_25755,N_26670);
or U33026 (N_33026,N_25166,N_28282);
and U33027 (N_33027,N_25976,N_29022);
nor U33028 (N_33028,N_26608,N_26096);
or U33029 (N_33029,N_25696,N_26685);
and U33030 (N_33030,N_27457,N_27964);
or U33031 (N_33031,N_29365,N_26594);
and U33032 (N_33032,N_26499,N_29227);
nor U33033 (N_33033,N_28265,N_29136);
xnor U33034 (N_33034,N_26390,N_26521);
nor U33035 (N_33035,N_27670,N_29564);
nand U33036 (N_33036,N_25084,N_26793);
nand U33037 (N_33037,N_26888,N_26625);
nand U33038 (N_33038,N_28050,N_28084);
or U33039 (N_33039,N_27847,N_27629);
nor U33040 (N_33040,N_27769,N_28633);
nand U33041 (N_33041,N_28074,N_26086);
and U33042 (N_33042,N_25592,N_29821);
or U33043 (N_33043,N_25875,N_27511);
xnor U33044 (N_33044,N_26719,N_25842);
nand U33045 (N_33045,N_25533,N_29837);
xnor U33046 (N_33046,N_26950,N_28240);
and U33047 (N_33047,N_26528,N_27520);
xor U33048 (N_33048,N_27274,N_25465);
and U33049 (N_33049,N_26547,N_27093);
xnor U33050 (N_33050,N_27594,N_25593);
or U33051 (N_33051,N_28237,N_29414);
and U33052 (N_33052,N_27553,N_28101);
nand U33053 (N_33053,N_25888,N_28555);
or U33054 (N_33054,N_26435,N_25174);
nand U33055 (N_33055,N_27610,N_28753);
nor U33056 (N_33056,N_26244,N_26016);
or U33057 (N_33057,N_25812,N_28428);
nor U33058 (N_33058,N_27863,N_29367);
or U33059 (N_33059,N_28318,N_27942);
xor U33060 (N_33060,N_26538,N_26549);
or U33061 (N_33061,N_26756,N_29558);
or U33062 (N_33062,N_29109,N_25625);
and U33063 (N_33063,N_28155,N_26350);
nor U33064 (N_33064,N_29805,N_29509);
xor U33065 (N_33065,N_25429,N_25564);
nor U33066 (N_33066,N_27029,N_26623);
nor U33067 (N_33067,N_27574,N_28859);
xor U33068 (N_33068,N_28703,N_26496);
nor U33069 (N_33069,N_29889,N_26208);
nand U33070 (N_33070,N_28493,N_27326);
xnor U33071 (N_33071,N_26492,N_27310);
nor U33072 (N_33072,N_25466,N_29803);
nor U33073 (N_33073,N_28469,N_28257);
nand U33074 (N_33074,N_28523,N_29068);
or U33075 (N_33075,N_27315,N_27430);
and U33076 (N_33076,N_29029,N_27856);
nand U33077 (N_33077,N_27770,N_25470);
or U33078 (N_33078,N_26561,N_27540);
xnor U33079 (N_33079,N_26886,N_29908);
or U33080 (N_33080,N_28482,N_25997);
or U33081 (N_33081,N_28052,N_26289);
or U33082 (N_33082,N_25527,N_27726);
and U33083 (N_33083,N_29438,N_26520);
and U33084 (N_33084,N_25819,N_28233);
nor U33085 (N_33085,N_28178,N_29642);
or U33086 (N_33086,N_26057,N_26168);
xor U33087 (N_33087,N_26134,N_28298);
nand U33088 (N_33088,N_28596,N_29646);
nand U33089 (N_33089,N_25346,N_26583);
nand U33090 (N_33090,N_25561,N_29949);
or U33091 (N_33091,N_27617,N_25101);
nor U33092 (N_33092,N_27913,N_29708);
and U33093 (N_33093,N_28423,N_25925);
or U33094 (N_33094,N_28865,N_25855);
or U33095 (N_33095,N_29271,N_27509);
nand U33096 (N_33096,N_29990,N_28332);
xor U33097 (N_33097,N_25872,N_28687);
and U33098 (N_33098,N_29329,N_28908);
and U33099 (N_33099,N_27095,N_29190);
nand U33100 (N_33100,N_25808,N_27815);
xnor U33101 (N_33101,N_29432,N_28551);
and U33102 (N_33102,N_27628,N_27102);
xnor U33103 (N_33103,N_26889,N_27357);
nand U33104 (N_33104,N_27138,N_28119);
nor U33105 (N_33105,N_29187,N_28186);
nand U33106 (N_33106,N_28707,N_25851);
or U33107 (N_33107,N_28448,N_27155);
or U33108 (N_33108,N_29312,N_26754);
xor U33109 (N_33109,N_28725,N_25861);
or U33110 (N_33110,N_28270,N_29971);
nand U33111 (N_33111,N_25116,N_26844);
and U33112 (N_33112,N_27295,N_26057);
nor U33113 (N_33113,N_28211,N_28447);
nor U33114 (N_33114,N_26326,N_28845);
xor U33115 (N_33115,N_26823,N_28402);
nand U33116 (N_33116,N_28652,N_29587);
nor U33117 (N_33117,N_26144,N_29035);
or U33118 (N_33118,N_25473,N_25945);
nand U33119 (N_33119,N_27669,N_25412);
nor U33120 (N_33120,N_25785,N_29233);
xor U33121 (N_33121,N_25516,N_25812);
xnor U33122 (N_33122,N_25250,N_27623);
and U33123 (N_33123,N_27230,N_29612);
xor U33124 (N_33124,N_27652,N_25173);
xor U33125 (N_33125,N_26078,N_29690);
or U33126 (N_33126,N_28685,N_29070);
or U33127 (N_33127,N_27130,N_29060);
xor U33128 (N_33128,N_28814,N_29433);
and U33129 (N_33129,N_28933,N_26974);
xnor U33130 (N_33130,N_29103,N_29340);
or U33131 (N_33131,N_28452,N_25348);
and U33132 (N_33132,N_28788,N_25378);
nand U33133 (N_33133,N_25017,N_25311);
or U33134 (N_33134,N_27075,N_28190);
xor U33135 (N_33135,N_27468,N_27569);
nand U33136 (N_33136,N_25911,N_26057);
nor U33137 (N_33137,N_25015,N_26582);
xnor U33138 (N_33138,N_27560,N_29939);
nor U33139 (N_33139,N_27990,N_26890);
xor U33140 (N_33140,N_28819,N_26593);
xor U33141 (N_33141,N_29401,N_26297);
nand U33142 (N_33142,N_25175,N_25864);
xor U33143 (N_33143,N_25465,N_27810);
nor U33144 (N_33144,N_27366,N_29308);
and U33145 (N_33145,N_25267,N_28912);
xnor U33146 (N_33146,N_26082,N_29128);
or U33147 (N_33147,N_27598,N_26471);
and U33148 (N_33148,N_28909,N_29391);
xnor U33149 (N_33149,N_28595,N_26891);
and U33150 (N_33150,N_26662,N_27096);
or U33151 (N_33151,N_25295,N_28426);
nand U33152 (N_33152,N_25406,N_27234);
and U33153 (N_33153,N_27698,N_29706);
xor U33154 (N_33154,N_26921,N_28872);
xor U33155 (N_33155,N_25052,N_27414);
and U33156 (N_33156,N_25567,N_25881);
or U33157 (N_33157,N_29744,N_26825);
nand U33158 (N_33158,N_27199,N_25529);
and U33159 (N_33159,N_29469,N_28326);
nor U33160 (N_33160,N_29564,N_29177);
nand U33161 (N_33161,N_29232,N_29781);
and U33162 (N_33162,N_25240,N_29568);
nor U33163 (N_33163,N_26379,N_25624);
nand U33164 (N_33164,N_25718,N_26794);
xor U33165 (N_33165,N_25791,N_26385);
or U33166 (N_33166,N_27889,N_27061);
nor U33167 (N_33167,N_28967,N_25737);
nand U33168 (N_33168,N_26577,N_26183);
or U33169 (N_33169,N_27126,N_27689);
nor U33170 (N_33170,N_27457,N_26220);
and U33171 (N_33171,N_27522,N_28936);
and U33172 (N_33172,N_26163,N_27044);
nand U33173 (N_33173,N_26880,N_27410);
and U33174 (N_33174,N_28070,N_26810);
xor U33175 (N_33175,N_25194,N_25313);
or U33176 (N_33176,N_28523,N_28097);
xor U33177 (N_33177,N_28295,N_29676);
nor U33178 (N_33178,N_25630,N_25077);
and U33179 (N_33179,N_29420,N_25128);
xor U33180 (N_33180,N_25618,N_26336);
or U33181 (N_33181,N_29989,N_25835);
or U33182 (N_33182,N_28677,N_28151);
or U33183 (N_33183,N_27365,N_26184);
and U33184 (N_33184,N_27141,N_28849);
nand U33185 (N_33185,N_28799,N_25529);
xnor U33186 (N_33186,N_26504,N_27986);
nand U33187 (N_33187,N_27866,N_28119);
xor U33188 (N_33188,N_27415,N_27984);
xnor U33189 (N_33189,N_27733,N_26100);
and U33190 (N_33190,N_28688,N_29807);
and U33191 (N_33191,N_27063,N_27052);
nand U33192 (N_33192,N_26869,N_25523);
or U33193 (N_33193,N_26346,N_25224);
nor U33194 (N_33194,N_25996,N_29831);
nor U33195 (N_33195,N_27827,N_28064);
nor U33196 (N_33196,N_26675,N_25034);
nand U33197 (N_33197,N_29876,N_29279);
nor U33198 (N_33198,N_28989,N_27419);
or U33199 (N_33199,N_28893,N_29519);
and U33200 (N_33200,N_28941,N_27027);
xor U33201 (N_33201,N_28157,N_28286);
or U33202 (N_33202,N_27437,N_26144);
nand U33203 (N_33203,N_29274,N_28350);
and U33204 (N_33204,N_28200,N_25692);
or U33205 (N_33205,N_27374,N_29579);
nand U33206 (N_33206,N_29061,N_29012);
xnor U33207 (N_33207,N_27418,N_28362);
nand U33208 (N_33208,N_27931,N_28759);
nor U33209 (N_33209,N_29709,N_29691);
xnor U33210 (N_33210,N_29406,N_25285);
or U33211 (N_33211,N_25372,N_25124);
xor U33212 (N_33212,N_28865,N_26620);
or U33213 (N_33213,N_26457,N_25116);
xnor U33214 (N_33214,N_26719,N_25762);
nor U33215 (N_33215,N_29450,N_26742);
xor U33216 (N_33216,N_27923,N_26503);
and U33217 (N_33217,N_27513,N_26113);
and U33218 (N_33218,N_27871,N_28711);
and U33219 (N_33219,N_27618,N_26525);
nor U33220 (N_33220,N_28622,N_28511);
nand U33221 (N_33221,N_29973,N_26359);
or U33222 (N_33222,N_27631,N_29086);
nand U33223 (N_33223,N_29686,N_29072);
xnor U33224 (N_33224,N_29064,N_26716);
nand U33225 (N_33225,N_27434,N_25647);
nor U33226 (N_33226,N_29047,N_28100);
nor U33227 (N_33227,N_25102,N_29765);
and U33228 (N_33228,N_27876,N_29975);
or U33229 (N_33229,N_28137,N_29517);
nand U33230 (N_33230,N_25225,N_27800);
nor U33231 (N_33231,N_25775,N_29880);
or U33232 (N_33232,N_26625,N_26813);
xor U33233 (N_33233,N_29391,N_27336);
and U33234 (N_33234,N_27636,N_25238);
or U33235 (N_33235,N_26321,N_29846);
or U33236 (N_33236,N_25285,N_25733);
and U33237 (N_33237,N_29714,N_26391);
or U33238 (N_33238,N_27494,N_28828);
and U33239 (N_33239,N_28429,N_29216);
and U33240 (N_33240,N_29511,N_26609);
and U33241 (N_33241,N_25535,N_27430);
xor U33242 (N_33242,N_25523,N_29121);
nand U33243 (N_33243,N_27580,N_27160);
and U33244 (N_33244,N_26258,N_29065);
xnor U33245 (N_33245,N_29983,N_26746);
nand U33246 (N_33246,N_26108,N_27400);
xor U33247 (N_33247,N_25211,N_28602);
nand U33248 (N_33248,N_26084,N_27984);
and U33249 (N_33249,N_28879,N_28172);
nor U33250 (N_33250,N_25458,N_25166);
nor U33251 (N_33251,N_29814,N_28373);
nor U33252 (N_33252,N_28960,N_29627);
or U33253 (N_33253,N_28998,N_25411);
nor U33254 (N_33254,N_29653,N_28592);
nor U33255 (N_33255,N_27582,N_26365);
nor U33256 (N_33256,N_29605,N_27440);
nand U33257 (N_33257,N_27669,N_26495);
or U33258 (N_33258,N_28762,N_28287);
or U33259 (N_33259,N_27053,N_26055);
xnor U33260 (N_33260,N_27867,N_28631);
and U33261 (N_33261,N_26904,N_25445);
nor U33262 (N_33262,N_28014,N_29299);
xor U33263 (N_33263,N_25625,N_29329);
or U33264 (N_33264,N_26830,N_26324);
nor U33265 (N_33265,N_27462,N_27886);
and U33266 (N_33266,N_25305,N_27245);
xor U33267 (N_33267,N_29174,N_28396);
and U33268 (N_33268,N_29074,N_25069);
nor U33269 (N_33269,N_25198,N_28521);
and U33270 (N_33270,N_26503,N_28947);
nand U33271 (N_33271,N_29345,N_29152);
and U33272 (N_33272,N_27314,N_26551);
and U33273 (N_33273,N_27041,N_29538);
xor U33274 (N_33274,N_28806,N_29010);
xnor U33275 (N_33275,N_29505,N_28486);
nand U33276 (N_33276,N_29251,N_27398);
and U33277 (N_33277,N_29472,N_28917);
xor U33278 (N_33278,N_29508,N_26224);
and U33279 (N_33279,N_25341,N_25600);
or U33280 (N_33280,N_25005,N_29039);
or U33281 (N_33281,N_29610,N_27578);
or U33282 (N_33282,N_25035,N_25036);
nor U33283 (N_33283,N_26395,N_25730);
and U33284 (N_33284,N_28370,N_26126);
or U33285 (N_33285,N_28667,N_29600);
and U33286 (N_33286,N_25693,N_29953);
nand U33287 (N_33287,N_27684,N_27694);
xnor U33288 (N_33288,N_27878,N_28736);
or U33289 (N_33289,N_29596,N_28455);
nor U33290 (N_33290,N_25648,N_26912);
or U33291 (N_33291,N_26339,N_29786);
nand U33292 (N_33292,N_29738,N_26267);
or U33293 (N_33293,N_26636,N_26002);
nor U33294 (N_33294,N_27249,N_27922);
or U33295 (N_33295,N_29001,N_27084);
and U33296 (N_33296,N_25898,N_25294);
xor U33297 (N_33297,N_28569,N_28235);
xor U33298 (N_33298,N_25043,N_29214);
or U33299 (N_33299,N_26894,N_27634);
and U33300 (N_33300,N_28267,N_26418);
or U33301 (N_33301,N_28061,N_27179);
nand U33302 (N_33302,N_28077,N_28497);
nor U33303 (N_33303,N_29826,N_26093);
xnor U33304 (N_33304,N_28035,N_26415);
xnor U33305 (N_33305,N_29331,N_29192);
nand U33306 (N_33306,N_25727,N_25525);
and U33307 (N_33307,N_29661,N_29213);
xor U33308 (N_33308,N_27930,N_28333);
xnor U33309 (N_33309,N_27917,N_27206);
nand U33310 (N_33310,N_29102,N_29879);
xnor U33311 (N_33311,N_27717,N_29872);
and U33312 (N_33312,N_29488,N_29319);
xor U33313 (N_33313,N_29324,N_28515);
xor U33314 (N_33314,N_27638,N_27687);
nor U33315 (N_33315,N_28577,N_28521);
or U33316 (N_33316,N_26469,N_27339);
nand U33317 (N_33317,N_29128,N_29762);
nor U33318 (N_33318,N_25374,N_25136);
xor U33319 (N_33319,N_29315,N_27721);
nor U33320 (N_33320,N_27427,N_25707);
or U33321 (N_33321,N_29076,N_27013);
and U33322 (N_33322,N_25940,N_27961);
nor U33323 (N_33323,N_29445,N_28946);
nand U33324 (N_33324,N_27347,N_29616);
or U33325 (N_33325,N_28561,N_25523);
nor U33326 (N_33326,N_28737,N_26448);
nand U33327 (N_33327,N_29530,N_26825);
nand U33328 (N_33328,N_28660,N_26939);
and U33329 (N_33329,N_26218,N_27509);
and U33330 (N_33330,N_26434,N_25521);
nor U33331 (N_33331,N_27415,N_25501);
xnor U33332 (N_33332,N_26670,N_28777);
and U33333 (N_33333,N_27588,N_28348);
nor U33334 (N_33334,N_28690,N_27032);
or U33335 (N_33335,N_25510,N_26459);
xnor U33336 (N_33336,N_27594,N_25842);
or U33337 (N_33337,N_25235,N_29327);
or U33338 (N_33338,N_28212,N_28679);
or U33339 (N_33339,N_27858,N_25618);
and U33340 (N_33340,N_26921,N_27459);
xnor U33341 (N_33341,N_25261,N_28848);
nand U33342 (N_33342,N_27820,N_28900);
nand U33343 (N_33343,N_29072,N_28395);
or U33344 (N_33344,N_27865,N_26236);
nor U33345 (N_33345,N_26696,N_28495);
nor U33346 (N_33346,N_28156,N_28304);
nor U33347 (N_33347,N_27345,N_26191);
and U33348 (N_33348,N_25945,N_25625);
xnor U33349 (N_33349,N_29164,N_26463);
xnor U33350 (N_33350,N_29101,N_28089);
and U33351 (N_33351,N_27852,N_25340);
xnor U33352 (N_33352,N_27703,N_26825);
xor U33353 (N_33353,N_25063,N_26338);
xor U33354 (N_33354,N_29964,N_26795);
and U33355 (N_33355,N_28829,N_29940);
xor U33356 (N_33356,N_27380,N_27274);
nor U33357 (N_33357,N_26906,N_29148);
or U33358 (N_33358,N_28555,N_29710);
or U33359 (N_33359,N_27852,N_27260);
or U33360 (N_33360,N_26170,N_26227);
or U33361 (N_33361,N_29307,N_29931);
and U33362 (N_33362,N_26488,N_27016);
nor U33363 (N_33363,N_27012,N_29116);
and U33364 (N_33364,N_26207,N_29185);
xor U33365 (N_33365,N_27278,N_26396);
xor U33366 (N_33366,N_27705,N_28854);
and U33367 (N_33367,N_28862,N_29414);
and U33368 (N_33368,N_26495,N_28199);
xnor U33369 (N_33369,N_25063,N_28876);
or U33370 (N_33370,N_28045,N_28287);
or U33371 (N_33371,N_26049,N_26682);
xnor U33372 (N_33372,N_29304,N_29079);
nor U33373 (N_33373,N_27461,N_27972);
xnor U33374 (N_33374,N_26156,N_27798);
xnor U33375 (N_33375,N_27436,N_29860);
or U33376 (N_33376,N_28333,N_28320);
and U33377 (N_33377,N_25309,N_28051);
or U33378 (N_33378,N_26355,N_27200);
and U33379 (N_33379,N_28913,N_25772);
or U33380 (N_33380,N_29968,N_29645);
nand U33381 (N_33381,N_27552,N_27408);
nand U33382 (N_33382,N_29492,N_29279);
and U33383 (N_33383,N_27370,N_27286);
or U33384 (N_33384,N_26152,N_27559);
nor U33385 (N_33385,N_29934,N_25510);
xor U33386 (N_33386,N_27324,N_25398);
xnor U33387 (N_33387,N_25932,N_27632);
or U33388 (N_33388,N_29349,N_27426);
and U33389 (N_33389,N_29073,N_29307);
nand U33390 (N_33390,N_27299,N_26952);
nor U33391 (N_33391,N_25236,N_28949);
and U33392 (N_33392,N_28464,N_28045);
or U33393 (N_33393,N_29117,N_27928);
nand U33394 (N_33394,N_27578,N_27765);
and U33395 (N_33395,N_28068,N_27959);
xnor U33396 (N_33396,N_29800,N_25940);
nand U33397 (N_33397,N_27797,N_29691);
nor U33398 (N_33398,N_29502,N_27283);
xnor U33399 (N_33399,N_28582,N_26196);
xnor U33400 (N_33400,N_25314,N_25895);
xnor U33401 (N_33401,N_27499,N_25754);
and U33402 (N_33402,N_25077,N_26626);
or U33403 (N_33403,N_29502,N_25041);
and U33404 (N_33404,N_25517,N_29492);
xor U33405 (N_33405,N_25811,N_29370);
or U33406 (N_33406,N_26814,N_25646);
xor U33407 (N_33407,N_29868,N_26719);
nor U33408 (N_33408,N_29772,N_26681);
xnor U33409 (N_33409,N_27292,N_27067);
nor U33410 (N_33410,N_28147,N_26332);
nor U33411 (N_33411,N_26399,N_28549);
nor U33412 (N_33412,N_26849,N_28905);
and U33413 (N_33413,N_25685,N_25128);
nand U33414 (N_33414,N_27358,N_27420);
or U33415 (N_33415,N_27392,N_26245);
and U33416 (N_33416,N_25420,N_29828);
nor U33417 (N_33417,N_25358,N_29354);
and U33418 (N_33418,N_27674,N_27542);
or U33419 (N_33419,N_25743,N_28848);
or U33420 (N_33420,N_26594,N_29809);
and U33421 (N_33421,N_28760,N_26723);
and U33422 (N_33422,N_29242,N_25273);
nand U33423 (N_33423,N_26912,N_26731);
xor U33424 (N_33424,N_25315,N_27335);
nor U33425 (N_33425,N_25949,N_25034);
or U33426 (N_33426,N_26202,N_25956);
nor U33427 (N_33427,N_27430,N_25630);
xnor U33428 (N_33428,N_25001,N_27640);
and U33429 (N_33429,N_28989,N_26376);
xnor U33430 (N_33430,N_27873,N_29323);
and U33431 (N_33431,N_28630,N_25155);
and U33432 (N_33432,N_25641,N_26781);
nand U33433 (N_33433,N_27301,N_27361);
or U33434 (N_33434,N_29058,N_27760);
nor U33435 (N_33435,N_29497,N_29923);
nor U33436 (N_33436,N_29693,N_28417);
and U33437 (N_33437,N_29312,N_26676);
nor U33438 (N_33438,N_26754,N_26205);
and U33439 (N_33439,N_26088,N_26981);
nor U33440 (N_33440,N_27558,N_27028);
nor U33441 (N_33441,N_26359,N_25101);
nor U33442 (N_33442,N_25961,N_29773);
or U33443 (N_33443,N_27006,N_25374);
nand U33444 (N_33444,N_26779,N_26838);
xnor U33445 (N_33445,N_27038,N_28215);
nand U33446 (N_33446,N_29902,N_26472);
nand U33447 (N_33447,N_26454,N_26947);
or U33448 (N_33448,N_29639,N_29381);
and U33449 (N_33449,N_25127,N_28621);
nand U33450 (N_33450,N_28872,N_26340);
and U33451 (N_33451,N_27286,N_28814);
or U33452 (N_33452,N_26435,N_29534);
nor U33453 (N_33453,N_29530,N_27735);
and U33454 (N_33454,N_28314,N_28918);
or U33455 (N_33455,N_26768,N_29168);
and U33456 (N_33456,N_27867,N_27987);
nor U33457 (N_33457,N_28971,N_25226);
nand U33458 (N_33458,N_29970,N_28444);
and U33459 (N_33459,N_27277,N_29081);
or U33460 (N_33460,N_29284,N_27071);
nand U33461 (N_33461,N_27422,N_26585);
and U33462 (N_33462,N_29875,N_29625);
xor U33463 (N_33463,N_29203,N_29739);
nor U33464 (N_33464,N_26993,N_27470);
and U33465 (N_33465,N_28118,N_27539);
nand U33466 (N_33466,N_26716,N_25705);
or U33467 (N_33467,N_27296,N_28663);
nand U33468 (N_33468,N_29700,N_26427);
or U33469 (N_33469,N_25140,N_29955);
nor U33470 (N_33470,N_27083,N_29999);
nand U33471 (N_33471,N_27269,N_25191);
and U33472 (N_33472,N_26781,N_29017);
nor U33473 (N_33473,N_29722,N_27925);
and U33474 (N_33474,N_29108,N_26928);
nand U33475 (N_33475,N_26213,N_28347);
nand U33476 (N_33476,N_29561,N_29491);
and U33477 (N_33477,N_26680,N_27694);
nor U33478 (N_33478,N_29241,N_27615);
nor U33479 (N_33479,N_28971,N_28830);
nand U33480 (N_33480,N_28431,N_28040);
nand U33481 (N_33481,N_26158,N_25163);
nor U33482 (N_33482,N_25689,N_26052);
or U33483 (N_33483,N_26596,N_25320);
xor U33484 (N_33484,N_28410,N_28421);
xor U33485 (N_33485,N_26794,N_28359);
and U33486 (N_33486,N_25297,N_27910);
xor U33487 (N_33487,N_29614,N_28180);
xor U33488 (N_33488,N_27890,N_26203);
and U33489 (N_33489,N_26669,N_29960);
xor U33490 (N_33490,N_29183,N_28176);
and U33491 (N_33491,N_25584,N_26442);
nand U33492 (N_33492,N_25268,N_28221);
xor U33493 (N_33493,N_28183,N_25937);
or U33494 (N_33494,N_27282,N_25046);
nand U33495 (N_33495,N_27268,N_29100);
xor U33496 (N_33496,N_28340,N_28364);
and U33497 (N_33497,N_27852,N_25217);
nand U33498 (N_33498,N_26050,N_25796);
or U33499 (N_33499,N_25814,N_26226);
nor U33500 (N_33500,N_26105,N_26563);
and U33501 (N_33501,N_25129,N_27764);
nand U33502 (N_33502,N_25130,N_29456);
and U33503 (N_33503,N_28720,N_26629);
xor U33504 (N_33504,N_28635,N_25243);
nand U33505 (N_33505,N_28642,N_25616);
nor U33506 (N_33506,N_29461,N_28230);
or U33507 (N_33507,N_25536,N_25196);
nor U33508 (N_33508,N_25885,N_25983);
or U33509 (N_33509,N_28426,N_29025);
xnor U33510 (N_33510,N_27075,N_29878);
and U33511 (N_33511,N_27524,N_25834);
and U33512 (N_33512,N_27838,N_25531);
or U33513 (N_33513,N_29788,N_28562);
xnor U33514 (N_33514,N_25119,N_27618);
nand U33515 (N_33515,N_28308,N_25003);
xnor U33516 (N_33516,N_25789,N_25601);
nor U33517 (N_33517,N_26833,N_29644);
xnor U33518 (N_33518,N_29212,N_25421);
and U33519 (N_33519,N_27672,N_27928);
nor U33520 (N_33520,N_27181,N_28135);
xor U33521 (N_33521,N_28137,N_27246);
or U33522 (N_33522,N_27751,N_28556);
or U33523 (N_33523,N_29111,N_29310);
xor U33524 (N_33524,N_26342,N_25228);
or U33525 (N_33525,N_29240,N_25642);
xor U33526 (N_33526,N_26585,N_29874);
xnor U33527 (N_33527,N_29533,N_29082);
nand U33528 (N_33528,N_25422,N_28323);
or U33529 (N_33529,N_28607,N_26873);
or U33530 (N_33530,N_26626,N_25083);
nor U33531 (N_33531,N_25439,N_29492);
nor U33532 (N_33532,N_29360,N_28363);
nor U33533 (N_33533,N_28703,N_25709);
xor U33534 (N_33534,N_26662,N_25444);
xor U33535 (N_33535,N_27277,N_28811);
and U33536 (N_33536,N_29470,N_25430);
xnor U33537 (N_33537,N_28873,N_26253);
or U33538 (N_33538,N_28855,N_28578);
nor U33539 (N_33539,N_26569,N_28576);
nand U33540 (N_33540,N_29729,N_25743);
xnor U33541 (N_33541,N_28433,N_29878);
nor U33542 (N_33542,N_25043,N_28919);
or U33543 (N_33543,N_26554,N_28906);
nor U33544 (N_33544,N_27367,N_25652);
nand U33545 (N_33545,N_28913,N_27843);
or U33546 (N_33546,N_25475,N_29936);
nand U33547 (N_33547,N_26326,N_29536);
nand U33548 (N_33548,N_25404,N_26199);
nor U33549 (N_33549,N_27692,N_27714);
and U33550 (N_33550,N_26064,N_27968);
nand U33551 (N_33551,N_28898,N_29253);
nor U33552 (N_33552,N_28472,N_27175);
and U33553 (N_33553,N_25266,N_26326);
and U33554 (N_33554,N_25203,N_29900);
nand U33555 (N_33555,N_25312,N_25392);
and U33556 (N_33556,N_29354,N_26842);
nor U33557 (N_33557,N_25044,N_27281);
and U33558 (N_33558,N_28335,N_26238);
xnor U33559 (N_33559,N_26549,N_26082);
or U33560 (N_33560,N_25572,N_26304);
xnor U33561 (N_33561,N_29170,N_28810);
or U33562 (N_33562,N_29866,N_27560);
nand U33563 (N_33563,N_26089,N_29535);
or U33564 (N_33564,N_28011,N_26252);
nor U33565 (N_33565,N_26015,N_27763);
nand U33566 (N_33566,N_26647,N_29292);
nor U33567 (N_33567,N_25146,N_26588);
nand U33568 (N_33568,N_27452,N_28729);
nand U33569 (N_33569,N_27558,N_27485);
nand U33570 (N_33570,N_26761,N_28153);
or U33571 (N_33571,N_27892,N_26720);
and U33572 (N_33572,N_25157,N_27991);
or U33573 (N_33573,N_29088,N_29614);
or U33574 (N_33574,N_27979,N_25007);
nor U33575 (N_33575,N_25644,N_26213);
or U33576 (N_33576,N_26092,N_28276);
or U33577 (N_33577,N_28821,N_28362);
or U33578 (N_33578,N_28733,N_28820);
nand U33579 (N_33579,N_29760,N_29407);
xor U33580 (N_33580,N_25687,N_26344);
or U33581 (N_33581,N_29851,N_28125);
and U33582 (N_33582,N_26158,N_26305);
and U33583 (N_33583,N_27868,N_29986);
nand U33584 (N_33584,N_29535,N_28100);
xnor U33585 (N_33585,N_26003,N_28407);
and U33586 (N_33586,N_29907,N_29403);
or U33587 (N_33587,N_25014,N_27638);
xnor U33588 (N_33588,N_28917,N_29217);
and U33589 (N_33589,N_27419,N_28093);
or U33590 (N_33590,N_26621,N_28252);
and U33591 (N_33591,N_26480,N_25739);
nor U33592 (N_33592,N_26112,N_27270);
nor U33593 (N_33593,N_26568,N_29505);
and U33594 (N_33594,N_25198,N_28063);
xnor U33595 (N_33595,N_29404,N_29186);
and U33596 (N_33596,N_29159,N_26289);
nor U33597 (N_33597,N_28618,N_29590);
xnor U33598 (N_33598,N_27727,N_25355);
nand U33599 (N_33599,N_27328,N_26729);
and U33600 (N_33600,N_25078,N_26920);
and U33601 (N_33601,N_27370,N_28797);
xor U33602 (N_33602,N_29846,N_28544);
nor U33603 (N_33603,N_27948,N_29118);
and U33604 (N_33604,N_28817,N_29807);
and U33605 (N_33605,N_28568,N_29543);
nand U33606 (N_33606,N_29343,N_28754);
or U33607 (N_33607,N_25153,N_28417);
or U33608 (N_33608,N_27085,N_28079);
xnor U33609 (N_33609,N_27791,N_29413);
nand U33610 (N_33610,N_25416,N_27284);
or U33611 (N_33611,N_25375,N_29428);
nand U33612 (N_33612,N_29022,N_29333);
or U33613 (N_33613,N_25524,N_29269);
nand U33614 (N_33614,N_26766,N_26075);
and U33615 (N_33615,N_28855,N_25825);
nor U33616 (N_33616,N_25582,N_25861);
xor U33617 (N_33617,N_25494,N_29694);
nor U33618 (N_33618,N_25597,N_29539);
and U33619 (N_33619,N_29783,N_28368);
nor U33620 (N_33620,N_28774,N_25934);
nor U33621 (N_33621,N_27264,N_29790);
and U33622 (N_33622,N_26884,N_25174);
and U33623 (N_33623,N_29941,N_25509);
xor U33624 (N_33624,N_25741,N_27727);
nand U33625 (N_33625,N_27818,N_28679);
or U33626 (N_33626,N_26580,N_26438);
nand U33627 (N_33627,N_27240,N_28030);
and U33628 (N_33628,N_27443,N_27624);
or U33629 (N_33629,N_25145,N_28542);
xor U33630 (N_33630,N_29791,N_26229);
and U33631 (N_33631,N_29081,N_29287);
nor U33632 (N_33632,N_29387,N_25529);
and U33633 (N_33633,N_28479,N_29482);
xnor U33634 (N_33634,N_27171,N_29654);
nand U33635 (N_33635,N_27212,N_29173);
nand U33636 (N_33636,N_25133,N_29336);
nand U33637 (N_33637,N_26960,N_27901);
nand U33638 (N_33638,N_27541,N_27550);
or U33639 (N_33639,N_28365,N_28759);
nand U33640 (N_33640,N_29565,N_28588);
xnor U33641 (N_33641,N_25657,N_26677);
nand U33642 (N_33642,N_29522,N_25114);
or U33643 (N_33643,N_29087,N_25972);
nand U33644 (N_33644,N_26336,N_29670);
or U33645 (N_33645,N_29857,N_26742);
xnor U33646 (N_33646,N_25811,N_28044);
or U33647 (N_33647,N_29612,N_27144);
and U33648 (N_33648,N_26503,N_25126);
nand U33649 (N_33649,N_25619,N_28534);
nand U33650 (N_33650,N_27988,N_28147);
or U33651 (N_33651,N_27734,N_29683);
nand U33652 (N_33652,N_27601,N_27353);
and U33653 (N_33653,N_27565,N_26227);
xor U33654 (N_33654,N_28400,N_26428);
and U33655 (N_33655,N_28894,N_25724);
nor U33656 (N_33656,N_29367,N_26399);
nor U33657 (N_33657,N_27920,N_25291);
and U33658 (N_33658,N_28136,N_27899);
nand U33659 (N_33659,N_25441,N_25664);
or U33660 (N_33660,N_28398,N_27423);
xnor U33661 (N_33661,N_27250,N_29630);
nand U33662 (N_33662,N_25705,N_26324);
xnor U33663 (N_33663,N_25192,N_26666);
xor U33664 (N_33664,N_29076,N_27037);
and U33665 (N_33665,N_28190,N_27692);
nand U33666 (N_33666,N_26923,N_25285);
and U33667 (N_33667,N_29172,N_27927);
and U33668 (N_33668,N_26586,N_25212);
xnor U33669 (N_33669,N_25506,N_27125);
or U33670 (N_33670,N_27818,N_25982);
xor U33671 (N_33671,N_28856,N_29863);
and U33672 (N_33672,N_29968,N_27190);
xnor U33673 (N_33673,N_28680,N_28565);
nand U33674 (N_33674,N_28708,N_27633);
nand U33675 (N_33675,N_25596,N_27927);
xor U33676 (N_33676,N_28643,N_27914);
or U33677 (N_33677,N_25706,N_28130);
nand U33678 (N_33678,N_29639,N_25391);
nand U33679 (N_33679,N_27841,N_27710);
nand U33680 (N_33680,N_27347,N_29280);
or U33681 (N_33681,N_25171,N_26976);
nor U33682 (N_33682,N_28069,N_26284);
nand U33683 (N_33683,N_29544,N_29002);
nand U33684 (N_33684,N_25055,N_26611);
nand U33685 (N_33685,N_25725,N_28136);
xnor U33686 (N_33686,N_27299,N_26277);
xor U33687 (N_33687,N_28303,N_28973);
nor U33688 (N_33688,N_25256,N_29313);
nor U33689 (N_33689,N_25119,N_25522);
xnor U33690 (N_33690,N_29619,N_29741);
and U33691 (N_33691,N_28744,N_28235);
nand U33692 (N_33692,N_29788,N_26237);
nor U33693 (N_33693,N_28544,N_29554);
xor U33694 (N_33694,N_26858,N_26784);
xor U33695 (N_33695,N_26068,N_25434);
nand U33696 (N_33696,N_25259,N_25114);
and U33697 (N_33697,N_29863,N_25969);
xor U33698 (N_33698,N_29522,N_27877);
xnor U33699 (N_33699,N_27544,N_29243);
and U33700 (N_33700,N_28125,N_25736);
or U33701 (N_33701,N_26703,N_29018);
or U33702 (N_33702,N_29130,N_29103);
nand U33703 (N_33703,N_26175,N_28849);
nand U33704 (N_33704,N_27817,N_26958);
nor U33705 (N_33705,N_29825,N_28961);
or U33706 (N_33706,N_25658,N_28791);
nand U33707 (N_33707,N_29565,N_29475);
nor U33708 (N_33708,N_26046,N_28058);
xnor U33709 (N_33709,N_27929,N_26953);
nor U33710 (N_33710,N_26177,N_25480);
nor U33711 (N_33711,N_25578,N_29907);
xor U33712 (N_33712,N_25095,N_25684);
or U33713 (N_33713,N_29088,N_25585);
nor U33714 (N_33714,N_28076,N_27338);
xnor U33715 (N_33715,N_28966,N_25019);
xnor U33716 (N_33716,N_25173,N_29298);
xnor U33717 (N_33717,N_25957,N_25116);
or U33718 (N_33718,N_26453,N_25373);
xor U33719 (N_33719,N_25488,N_25413);
nor U33720 (N_33720,N_27366,N_25026);
nor U33721 (N_33721,N_26903,N_26072);
nand U33722 (N_33722,N_29796,N_28033);
or U33723 (N_33723,N_26514,N_25353);
xor U33724 (N_33724,N_29594,N_26141);
nand U33725 (N_33725,N_26357,N_26309);
nor U33726 (N_33726,N_26065,N_29531);
xnor U33727 (N_33727,N_27988,N_27483);
xnor U33728 (N_33728,N_28848,N_25374);
or U33729 (N_33729,N_27456,N_27136);
xnor U33730 (N_33730,N_27169,N_27098);
nand U33731 (N_33731,N_27583,N_25927);
nor U33732 (N_33732,N_26756,N_25002);
and U33733 (N_33733,N_27534,N_29142);
nor U33734 (N_33734,N_28154,N_26179);
nand U33735 (N_33735,N_29755,N_26750);
nand U33736 (N_33736,N_29018,N_27012);
and U33737 (N_33737,N_25359,N_26340);
nor U33738 (N_33738,N_27400,N_25381);
nand U33739 (N_33739,N_25461,N_29664);
nor U33740 (N_33740,N_26475,N_28121);
nand U33741 (N_33741,N_26083,N_26898);
or U33742 (N_33742,N_26482,N_29543);
xnor U33743 (N_33743,N_26705,N_27425);
and U33744 (N_33744,N_26464,N_29919);
xor U33745 (N_33745,N_28477,N_25032);
and U33746 (N_33746,N_26398,N_29088);
nor U33747 (N_33747,N_28803,N_25426);
nand U33748 (N_33748,N_29465,N_26818);
xnor U33749 (N_33749,N_26527,N_27809);
xnor U33750 (N_33750,N_29437,N_29137);
xnor U33751 (N_33751,N_26969,N_26126);
nor U33752 (N_33752,N_26906,N_29134);
xor U33753 (N_33753,N_26413,N_26218);
or U33754 (N_33754,N_29196,N_25230);
nor U33755 (N_33755,N_27550,N_27769);
and U33756 (N_33756,N_26406,N_26480);
nand U33757 (N_33757,N_28303,N_25075);
xor U33758 (N_33758,N_27581,N_29360);
and U33759 (N_33759,N_25118,N_27571);
xor U33760 (N_33760,N_26935,N_28203);
nor U33761 (N_33761,N_26933,N_29118);
xnor U33762 (N_33762,N_26851,N_28255);
nand U33763 (N_33763,N_29849,N_26423);
xor U33764 (N_33764,N_27516,N_27301);
and U33765 (N_33765,N_28844,N_29597);
xnor U33766 (N_33766,N_25318,N_25980);
nand U33767 (N_33767,N_28867,N_27799);
xnor U33768 (N_33768,N_29036,N_28130);
or U33769 (N_33769,N_29826,N_25087);
nor U33770 (N_33770,N_29685,N_27935);
nor U33771 (N_33771,N_26424,N_26258);
nand U33772 (N_33772,N_28392,N_28386);
nand U33773 (N_33773,N_27599,N_26029);
nand U33774 (N_33774,N_28207,N_27493);
and U33775 (N_33775,N_28427,N_27588);
nand U33776 (N_33776,N_25237,N_26070);
or U33777 (N_33777,N_29104,N_27767);
or U33778 (N_33778,N_28012,N_28386);
nand U33779 (N_33779,N_26341,N_26528);
and U33780 (N_33780,N_25119,N_28594);
or U33781 (N_33781,N_29844,N_28338);
nor U33782 (N_33782,N_26990,N_29318);
xnor U33783 (N_33783,N_29738,N_28507);
nor U33784 (N_33784,N_26648,N_29233);
nor U33785 (N_33785,N_28382,N_25502);
and U33786 (N_33786,N_29319,N_28804);
nand U33787 (N_33787,N_26434,N_28116);
xor U33788 (N_33788,N_29272,N_29224);
nor U33789 (N_33789,N_28436,N_27298);
and U33790 (N_33790,N_25057,N_27970);
xor U33791 (N_33791,N_25952,N_29085);
nor U33792 (N_33792,N_25863,N_28438);
or U33793 (N_33793,N_28441,N_29818);
and U33794 (N_33794,N_28851,N_29777);
nand U33795 (N_33795,N_29446,N_25162);
and U33796 (N_33796,N_27452,N_27495);
nand U33797 (N_33797,N_26141,N_29162);
xnor U33798 (N_33798,N_28332,N_25826);
and U33799 (N_33799,N_29078,N_27983);
and U33800 (N_33800,N_29164,N_27764);
nor U33801 (N_33801,N_27976,N_29582);
or U33802 (N_33802,N_28809,N_27986);
nor U33803 (N_33803,N_25314,N_27119);
nand U33804 (N_33804,N_28883,N_29558);
or U33805 (N_33805,N_26305,N_26671);
and U33806 (N_33806,N_25493,N_26391);
or U33807 (N_33807,N_29201,N_29495);
and U33808 (N_33808,N_29830,N_29353);
nor U33809 (N_33809,N_26796,N_28282);
xnor U33810 (N_33810,N_27728,N_27992);
or U33811 (N_33811,N_29746,N_27723);
and U33812 (N_33812,N_29023,N_28179);
or U33813 (N_33813,N_27249,N_25721);
xor U33814 (N_33814,N_28782,N_25108);
or U33815 (N_33815,N_27102,N_25609);
and U33816 (N_33816,N_26863,N_25530);
or U33817 (N_33817,N_28984,N_28423);
or U33818 (N_33818,N_28952,N_26445);
and U33819 (N_33819,N_25792,N_26139);
xnor U33820 (N_33820,N_27407,N_25050);
xor U33821 (N_33821,N_25451,N_28145);
and U33822 (N_33822,N_26196,N_26420);
and U33823 (N_33823,N_26162,N_27661);
nand U33824 (N_33824,N_25299,N_28962);
nand U33825 (N_33825,N_29798,N_26875);
and U33826 (N_33826,N_28388,N_28421);
and U33827 (N_33827,N_28732,N_26454);
nor U33828 (N_33828,N_25722,N_25936);
nor U33829 (N_33829,N_25892,N_28585);
xnor U33830 (N_33830,N_26055,N_26267);
nand U33831 (N_33831,N_29828,N_29807);
nand U33832 (N_33832,N_26446,N_27992);
and U33833 (N_33833,N_28229,N_25915);
and U33834 (N_33834,N_27725,N_29004);
or U33835 (N_33835,N_27319,N_27366);
nor U33836 (N_33836,N_27087,N_29294);
and U33837 (N_33837,N_26980,N_28246);
or U33838 (N_33838,N_26248,N_29288);
xor U33839 (N_33839,N_25427,N_25800);
nor U33840 (N_33840,N_26953,N_29330);
xnor U33841 (N_33841,N_26049,N_27459);
xnor U33842 (N_33842,N_26929,N_25623);
and U33843 (N_33843,N_28960,N_26284);
nor U33844 (N_33844,N_27765,N_28606);
and U33845 (N_33845,N_25542,N_29312);
or U33846 (N_33846,N_25696,N_28935);
and U33847 (N_33847,N_27860,N_26369);
or U33848 (N_33848,N_25049,N_29981);
and U33849 (N_33849,N_25689,N_27866);
nand U33850 (N_33850,N_28895,N_26139);
nand U33851 (N_33851,N_26661,N_27209);
nor U33852 (N_33852,N_28443,N_26691);
xnor U33853 (N_33853,N_27005,N_26489);
nand U33854 (N_33854,N_25820,N_28347);
nor U33855 (N_33855,N_28997,N_27820);
nand U33856 (N_33856,N_29927,N_26868);
and U33857 (N_33857,N_27170,N_26023);
or U33858 (N_33858,N_28347,N_25966);
nand U33859 (N_33859,N_25789,N_28031);
nand U33860 (N_33860,N_27002,N_26685);
xor U33861 (N_33861,N_29333,N_25939);
nor U33862 (N_33862,N_26599,N_26544);
or U33863 (N_33863,N_29712,N_29882);
or U33864 (N_33864,N_26441,N_26901);
and U33865 (N_33865,N_27827,N_29313);
nand U33866 (N_33866,N_25143,N_25496);
xor U33867 (N_33867,N_28547,N_27815);
nor U33868 (N_33868,N_29028,N_25895);
and U33869 (N_33869,N_25671,N_27237);
nand U33870 (N_33870,N_26605,N_28818);
or U33871 (N_33871,N_26838,N_27010);
and U33872 (N_33872,N_26916,N_26005);
nand U33873 (N_33873,N_25723,N_29976);
xnor U33874 (N_33874,N_28367,N_28507);
xnor U33875 (N_33875,N_26046,N_27922);
or U33876 (N_33876,N_29353,N_29756);
or U33877 (N_33877,N_28470,N_27228);
nand U33878 (N_33878,N_27243,N_29484);
nand U33879 (N_33879,N_28139,N_27382);
and U33880 (N_33880,N_29062,N_29007);
nand U33881 (N_33881,N_28923,N_25375);
xnor U33882 (N_33882,N_25052,N_26489);
nor U33883 (N_33883,N_26438,N_28426);
nand U33884 (N_33884,N_27693,N_25441);
nand U33885 (N_33885,N_27608,N_26773);
or U33886 (N_33886,N_27242,N_29729);
xnor U33887 (N_33887,N_26159,N_29982);
nor U33888 (N_33888,N_25105,N_26390);
nor U33889 (N_33889,N_29121,N_28841);
or U33890 (N_33890,N_28935,N_26076);
xnor U33891 (N_33891,N_29351,N_28183);
nand U33892 (N_33892,N_25871,N_29039);
nand U33893 (N_33893,N_26916,N_28122);
nor U33894 (N_33894,N_25636,N_27953);
xnor U33895 (N_33895,N_27469,N_28524);
xor U33896 (N_33896,N_29845,N_29313);
nand U33897 (N_33897,N_28784,N_28500);
and U33898 (N_33898,N_25487,N_29717);
xor U33899 (N_33899,N_29138,N_28328);
nand U33900 (N_33900,N_26173,N_29422);
or U33901 (N_33901,N_28385,N_26100);
nand U33902 (N_33902,N_26807,N_27322);
nand U33903 (N_33903,N_26389,N_25250);
nand U33904 (N_33904,N_29233,N_27913);
nand U33905 (N_33905,N_25690,N_26730);
nand U33906 (N_33906,N_29867,N_29097);
and U33907 (N_33907,N_26469,N_25012);
nor U33908 (N_33908,N_27058,N_27587);
nor U33909 (N_33909,N_29922,N_26629);
xnor U33910 (N_33910,N_26797,N_28389);
and U33911 (N_33911,N_25547,N_26212);
nand U33912 (N_33912,N_26786,N_26393);
nor U33913 (N_33913,N_27443,N_25989);
or U33914 (N_33914,N_27962,N_28869);
and U33915 (N_33915,N_26822,N_27928);
xnor U33916 (N_33916,N_25540,N_25129);
or U33917 (N_33917,N_28589,N_25138);
and U33918 (N_33918,N_28246,N_29835);
or U33919 (N_33919,N_25674,N_25447);
and U33920 (N_33920,N_25703,N_29929);
nor U33921 (N_33921,N_25510,N_27351);
nand U33922 (N_33922,N_28206,N_29929);
nor U33923 (N_33923,N_28773,N_27563);
nand U33924 (N_33924,N_26246,N_27349);
nor U33925 (N_33925,N_29411,N_28359);
and U33926 (N_33926,N_29309,N_29956);
and U33927 (N_33927,N_29595,N_29097);
or U33928 (N_33928,N_26923,N_25101);
nand U33929 (N_33929,N_27058,N_27437);
nand U33930 (N_33930,N_27959,N_27844);
nor U33931 (N_33931,N_25659,N_25153);
nand U33932 (N_33932,N_27677,N_26943);
and U33933 (N_33933,N_28936,N_26515);
nand U33934 (N_33934,N_27749,N_27789);
xnor U33935 (N_33935,N_26881,N_26577);
xnor U33936 (N_33936,N_25088,N_25729);
or U33937 (N_33937,N_27190,N_27495);
xnor U33938 (N_33938,N_25864,N_29563);
nor U33939 (N_33939,N_28589,N_28851);
nor U33940 (N_33940,N_29106,N_27529);
and U33941 (N_33941,N_28999,N_29529);
and U33942 (N_33942,N_29473,N_29129);
xor U33943 (N_33943,N_26954,N_27475);
nor U33944 (N_33944,N_26483,N_26321);
nor U33945 (N_33945,N_29987,N_29347);
nand U33946 (N_33946,N_28256,N_25585);
xor U33947 (N_33947,N_26312,N_27183);
nor U33948 (N_33948,N_26965,N_25909);
nor U33949 (N_33949,N_27107,N_28029);
nand U33950 (N_33950,N_25098,N_27198);
and U33951 (N_33951,N_25075,N_28520);
nand U33952 (N_33952,N_26751,N_29324);
xnor U33953 (N_33953,N_25359,N_29316);
and U33954 (N_33954,N_25312,N_28454);
and U33955 (N_33955,N_29257,N_29242);
and U33956 (N_33956,N_27491,N_29380);
or U33957 (N_33957,N_26122,N_29909);
and U33958 (N_33958,N_29559,N_27214);
and U33959 (N_33959,N_29156,N_29323);
xnor U33960 (N_33960,N_26015,N_27810);
and U33961 (N_33961,N_25085,N_26510);
nand U33962 (N_33962,N_26393,N_25998);
nand U33963 (N_33963,N_29020,N_27166);
xor U33964 (N_33964,N_26683,N_25380);
nand U33965 (N_33965,N_27979,N_28659);
or U33966 (N_33966,N_27170,N_29676);
or U33967 (N_33967,N_27639,N_27090);
and U33968 (N_33968,N_29600,N_28495);
nor U33969 (N_33969,N_26149,N_27445);
or U33970 (N_33970,N_27115,N_28009);
nand U33971 (N_33971,N_25990,N_28966);
or U33972 (N_33972,N_27030,N_25789);
nor U33973 (N_33973,N_27189,N_26118);
nor U33974 (N_33974,N_26575,N_25753);
or U33975 (N_33975,N_25448,N_27205);
and U33976 (N_33976,N_26354,N_25240);
nand U33977 (N_33977,N_25244,N_28787);
and U33978 (N_33978,N_28120,N_29615);
or U33979 (N_33979,N_25407,N_28316);
nand U33980 (N_33980,N_26743,N_27980);
and U33981 (N_33981,N_26347,N_28883);
xor U33982 (N_33982,N_28148,N_27828);
and U33983 (N_33983,N_25308,N_27628);
nand U33984 (N_33984,N_26640,N_29270);
nand U33985 (N_33985,N_28150,N_25364);
and U33986 (N_33986,N_25697,N_26966);
and U33987 (N_33987,N_29505,N_29790);
nor U33988 (N_33988,N_29797,N_27044);
and U33989 (N_33989,N_28452,N_26966);
and U33990 (N_33990,N_27558,N_27146);
nand U33991 (N_33991,N_29980,N_27438);
and U33992 (N_33992,N_29178,N_29546);
nand U33993 (N_33993,N_27771,N_27537);
nor U33994 (N_33994,N_28041,N_29073);
or U33995 (N_33995,N_27193,N_25291);
xor U33996 (N_33996,N_28435,N_28968);
nor U33997 (N_33997,N_28658,N_26878);
or U33998 (N_33998,N_27373,N_26741);
and U33999 (N_33999,N_27492,N_26787);
nand U34000 (N_34000,N_28026,N_25602);
xor U34001 (N_34001,N_27394,N_28930);
nor U34002 (N_34002,N_25392,N_28090);
and U34003 (N_34003,N_26451,N_29004);
nand U34004 (N_34004,N_26435,N_28636);
nor U34005 (N_34005,N_26437,N_28904);
and U34006 (N_34006,N_26524,N_26483);
nand U34007 (N_34007,N_26798,N_25138);
xnor U34008 (N_34008,N_28764,N_29403);
nor U34009 (N_34009,N_27780,N_27473);
or U34010 (N_34010,N_26162,N_27377);
or U34011 (N_34011,N_29233,N_25124);
or U34012 (N_34012,N_29208,N_25330);
xnor U34013 (N_34013,N_27343,N_26564);
and U34014 (N_34014,N_26755,N_26288);
and U34015 (N_34015,N_29121,N_29519);
xnor U34016 (N_34016,N_26281,N_28986);
or U34017 (N_34017,N_29300,N_26309);
and U34018 (N_34018,N_25959,N_25420);
nor U34019 (N_34019,N_28198,N_25048);
nand U34020 (N_34020,N_26779,N_29343);
nor U34021 (N_34021,N_29221,N_26346);
and U34022 (N_34022,N_26357,N_28853);
xnor U34023 (N_34023,N_29377,N_29255);
and U34024 (N_34024,N_29517,N_27882);
or U34025 (N_34025,N_27738,N_29623);
nor U34026 (N_34026,N_26561,N_25595);
nor U34027 (N_34027,N_25311,N_28875);
or U34028 (N_34028,N_25857,N_26071);
nand U34029 (N_34029,N_26889,N_28857);
nand U34030 (N_34030,N_25972,N_25699);
or U34031 (N_34031,N_28789,N_25861);
or U34032 (N_34032,N_28461,N_29762);
xnor U34033 (N_34033,N_29231,N_28428);
or U34034 (N_34034,N_28194,N_29382);
and U34035 (N_34035,N_29331,N_27097);
nor U34036 (N_34036,N_25494,N_28320);
nor U34037 (N_34037,N_27113,N_27078);
nand U34038 (N_34038,N_29563,N_29949);
or U34039 (N_34039,N_26469,N_25587);
or U34040 (N_34040,N_27521,N_28913);
nand U34041 (N_34041,N_29391,N_27738);
xnor U34042 (N_34042,N_25759,N_28991);
or U34043 (N_34043,N_29305,N_28995);
nor U34044 (N_34044,N_29335,N_26707);
nor U34045 (N_34045,N_27567,N_27205);
or U34046 (N_34046,N_25195,N_25567);
and U34047 (N_34047,N_27358,N_27279);
and U34048 (N_34048,N_26631,N_25788);
and U34049 (N_34049,N_26374,N_29218);
nor U34050 (N_34050,N_26716,N_29515);
xnor U34051 (N_34051,N_27134,N_26235);
nor U34052 (N_34052,N_28161,N_26608);
xor U34053 (N_34053,N_27037,N_29455);
xor U34054 (N_34054,N_26632,N_26689);
nor U34055 (N_34055,N_28791,N_27463);
and U34056 (N_34056,N_29543,N_27401);
nor U34057 (N_34057,N_26765,N_29999);
nor U34058 (N_34058,N_26203,N_26288);
or U34059 (N_34059,N_29293,N_28470);
and U34060 (N_34060,N_27527,N_26780);
nor U34061 (N_34061,N_28614,N_29822);
or U34062 (N_34062,N_26827,N_25270);
nand U34063 (N_34063,N_28328,N_27267);
and U34064 (N_34064,N_28263,N_25525);
and U34065 (N_34065,N_27981,N_27323);
nor U34066 (N_34066,N_26383,N_26122);
or U34067 (N_34067,N_29681,N_26761);
nor U34068 (N_34068,N_29769,N_29794);
nor U34069 (N_34069,N_26638,N_26511);
nand U34070 (N_34070,N_29870,N_28011);
xnor U34071 (N_34071,N_27491,N_25034);
and U34072 (N_34072,N_27690,N_25386);
xor U34073 (N_34073,N_29050,N_26624);
xor U34074 (N_34074,N_26284,N_29904);
nand U34075 (N_34075,N_27340,N_28496);
and U34076 (N_34076,N_28475,N_25704);
xnor U34077 (N_34077,N_25499,N_25230);
and U34078 (N_34078,N_25158,N_25346);
and U34079 (N_34079,N_27529,N_28439);
nor U34080 (N_34080,N_27106,N_29971);
nor U34081 (N_34081,N_27664,N_26754);
and U34082 (N_34082,N_26153,N_28427);
nand U34083 (N_34083,N_29808,N_25868);
or U34084 (N_34084,N_26928,N_25876);
and U34085 (N_34085,N_25838,N_28908);
or U34086 (N_34086,N_26770,N_26151);
xnor U34087 (N_34087,N_29438,N_29168);
and U34088 (N_34088,N_26397,N_26896);
xnor U34089 (N_34089,N_25177,N_26115);
xor U34090 (N_34090,N_27547,N_28510);
or U34091 (N_34091,N_25835,N_29272);
nor U34092 (N_34092,N_27962,N_28556);
or U34093 (N_34093,N_25207,N_26976);
and U34094 (N_34094,N_25179,N_26688);
nand U34095 (N_34095,N_26308,N_28054);
and U34096 (N_34096,N_26346,N_25625);
or U34097 (N_34097,N_25346,N_29631);
xnor U34098 (N_34098,N_25472,N_25583);
xnor U34099 (N_34099,N_29202,N_26712);
and U34100 (N_34100,N_25816,N_27793);
nor U34101 (N_34101,N_28255,N_27420);
or U34102 (N_34102,N_29262,N_25980);
and U34103 (N_34103,N_26306,N_26814);
nor U34104 (N_34104,N_26897,N_25049);
and U34105 (N_34105,N_26253,N_26545);
nand U34106 (N_34106,N_29371,N_27767);
nor U34107 (N_34107,N_26725,N_28569);
and U34108 (N_34108,N_27623,N_27585);
nand U34109 (N_34109,N_28903,N_27640);
and U34110 (N_34110,N_29843,N_28932);
or U34111 (N_34111,N_28370,N_29100);
or U34112 (N_34112,N_25427,N_29819);
nor U34113 (N_34113,N_28946,N_25477);
nor U34114 (N_34114,N_29107,N_25297);
or U34115 (N_34115,N_27784,N_25404);
xor U34116 (N_34116,N_28740,N_27613);
nand U34117 (N_34117,N_26908,N_28385);
or U34118 (N_34118,N_29802,N_26575);
or U34119 (N_34119,N_27865,N_25887);
and U34120 (N_34120,N_25300,N_26304);
xor U34121 (N_34121,N_29237,N_29747);
and U34122 (N_34122,N_26922,N_25620);
or U34123 (N_34123,N_27909,N_28056);
xnor U34124 (N_34124,N_27055,N_25967);
or U34125 (N_34125,N_25610,N_27169);
nand U34126 (N_34126,N_26166,N_25742);
or U34127 (N_34127,N_26660,N_25833);
xor U34128 (N_34128,N_27387,N_26277);
xor U34129 (N_34129,N_27710,N_26209);
or U34130 (N_34130,N_25879,N_26591);
nor U34131 (N_34131,N_26846,N_26150);
or U34132 (N_34132,N_28614,N_27841);
xor U34133 (N_34133,N_27474,N_25872);
nand U34134 (N_34134,N_27945,N_27065);
xnor U34135 (N_34135,N_27903,N_28170);
and U34136 (N_34136,N_27459,N_27386);
or U34137 (N_34137,N_27455,N_25954);
nand U34138 (N_34138,N_25411,N_28073);
nor U34139 (N_34139,N_26296,N_29292);
or U34140 (N_34140,N_28060,N_25236);
or U34141 (N_34141,N_26731,N_28118);
or U34142 (N_34142,N_25672,N_29880);
nand U34143 (N_34143,N_29476,N_26031);
nor U34144 (N_34144,N_28099,N_27510);
and U34145 (N_34145,N_28342,N_26278);
or U34146 (N_34146,N_28190,N_27108);
and U34147 (N_34147,N_29853,N_28684);
nor U34148 (N_34148,N_27513,N_28407);
nand U34149 (N_34149,N_29586,N_29105);
and U34150 (N_34150,N_29215,N_25802);
and U34151 (N_34151,N_29753,N_28044);
nor U34152 (N_34152,N_26530,N_27255);
nand U34153 (N_34153,N_27772,N_25223);
nor U34154 (N_34154,N_27515,N_26693);
nor U34155 (N_34155,N_26749,N_29989);
nand U34156 (N_34156,N_26379,N_29923);
nand U34157 (N_34157,N_28609,N_27542);
and U34158 (N_34158,N_29192,N_27693);
nand U34159 (N_34159,N_26492,N_28135);
and U34160 (N_34160,N_29432,N_26118);
and U34161 (N_34161,N_29349,N_28772);
xnor U34162 (N_34162,N_25377,N_28850);
nor U34163 (N_34163,N_26535,N_27411);
and U34164 (N_34164,N_28266,N_26222);
nand U34165 (N_34165,N_27083,N_26415);
or U34166 (N_34166,N_29345,N_28668);
nor U34167 (N_34167,N_29658,N_29601);
xor U34168 (N_34168,N_25916,N_28525);
or U34169 (N_34169,N_29650,N_25912);
nand U34170 (N_34170,N_26420,N_25954);
nor U34171 (N_34171,N_27246,N_26130);
nor U34172 (N_34172,N_26238,N_26882);
nor U34173 (N_34173,N_28629,N_26612);
and U34174 (N_34174,N_26453,N_29836);
nand U34175 (N_34175,N_29649,N_26332);
xor U34176 (N_34176,N_29809,N_25942);
nor U34177 (N_34177,N_26160,N_26802);
and U34178 (N_34178,N_25098,N_29011);
xnor U34179 (N_34179,N_25964,N_25830);
nand U34180 (N_34180,N_27008,N_26134);
nand U34181 (N_34181,N_27366,N_27267);
nor U34182 (N_34182,N_25501,N_29254);
and U34183 (N_34183,N_28963,N_25407);
nor U34184 (N_34184,N_26440,N_28114);
nor U34185 (N_34185,N_25024,N_29797);
nand U34186 (N_34186,N_27218,N_29740);
xnor U34187 (N_34187,N_25407,N_27159);
xnor U34188 (N_34188,N_26692,N_28842);
nor U34189 (N_34189,N_28232,N_27556);
xor U34190 (N_34190,N_27030,N_25525);
xor U34191 (N_34191,N_28506,N_28462);
and U34192 (N_34192,N_29947,N_28691);
nand U34193 (N_34193,N_27868,N_28772);
or U34194 (N_34194,N_27866,N_27422);
xnor U34195 (N_34195,N_29818,N_25483);
xnor U34196 (N_34196,N_29074,N_25556);
and U34197 (N_34197,N_27515,N_29301);
nand U34198 (N_34198,N_27933,N_29284);
xnor U34199 (N_34199,N_26261,N_29542);
or U34200 (N_34200,N_25548,N_29144);
xor U34201 (N_34201,N_26396,N_27924);
nand U34202 (N_34202,N_25883,N_28259);
or U34203 (N_34203,N_29869,N_27882);
xnor U34204 (N_34204,N_29343,N_26120);
nor U34205 (N_34205,N_27882,N_26697);
and U34206 (N_34206,N_25227,N_25150);
or U34207 (N_34207,N_26574,N_29503);
and U34208 (N_34208,N_26675,N_26134);
nor U34209 (N_34209,N_29163,N_26825);
nand U34210 (N_34210,N_26189,N_28249);
and U34211 (N_34211,N_26807,N_26835);
xor U34212 (N_34212,N_26397,N_26851);
and U34213 (N_34213,N_29514,N_28186);
nand U34214 (N_34214,N_26735,N_29002);
nand U34215 (N_34215,N_25564,N_27685);
xnor U34216 (N_34216,N_27693,N_27529);
or U34217 (N_34217,N_29799,N_28883);
nor U34218 (N_34218,N_27930,N_26314);
or U34219 (N_34219,N_26998,N_27996);
and U34220 (N_34220,N_27713,N_27873);
xor U34221 (N_34221,N_25233,N_29767);
xor U34222 (N_34222,N_28217,N_25765);
xor U34223 (N_34223,N_26681,N_27940);
nor U34224 (N_34224,N_26428,N_26475);
or U34225 (N_34225,N_25699,N_27929);
or U34226 (N_34226,N_25797,N_27840);
xnor U34227 (N_34227,N_29780,N_27915);
and U34228 (N_34228,N_26917,N_28745);
or U34229 (N_34229,N_29381,N_28477);
or U34230 (N_34230,N_29239,N_27271);
and U34231 (N_34231,N_28978,N_25480);
and U34232 (N_34232,N_25643,N_28007);
xnor U34233 (N_34233,N_28207,N_26039);
or U34234 (N_34234,N_27112,N_25444);
nand U34235 (N_34235,N_26654,N_29707);
or U34236 (N_34236,N_26828,N_27416);
and U34237 (N_34237,N_29396,N_26773);
and U34238 (N_34238,N_29050,N_29496);
xnor U34239 (N_34239,N_29130,N_29147);
or U34240 (N_34240,N_25686,N_28596);
nand U34241 (N_34241,N_29271,N_25050);
xor U34242 (N_34242,N_25587,N_25851);
and U34243 (N_34243,N_28172,N_28546);
or U34244 (N_34244,N_25607,N_27993);
xor U34245 (N_34245,N_28742,N_29972);
xor U34246 (N_34246,N_26759,N_28037);
nand U34247 (N_34247,N_29224,N_25760);
nor U34248 (N_34248,N_28106,N_28129);
nand U34249 (N_34249,N_26386,N_26279);
nor U34250 (N_34250,N_28208,N_29612);
nand U34251 (N_34251,N_29682,N_27007);
nor U34252 (N_34252,N_28099,N_29291);
nand U34253 (N_34253,N_29584,N_26337);
nor U34254 (N_34254,N_26483,N_27015);
xor U34255 (N_34255,N_26686,N_28971);
nor U34256 (N_34256,N_28044,N_25831);
xnor U34257 (N_34257,N_28974,N_26932);
and U34258 (N_34258,N_26650,N_28268);
and U34259 (N_34259,N_25307,N_26705);
nor U34260 (N_34260,N_25488,N_27178);
and U34261 (N_34261,N_25390,N_26320);
nor U34262 (N_34262,N_29668,N_28450);
and U34263 (N_34263,N_27927,N_26204);
or U34264 (N_34264,N_25991,N_26246);
nand U34265 (N_34265,N_26340,N_28502);
or U34266 (N_34266,N_28002,N_25145);
nor U34267 (N_34267,N_27147,N_29270);
nand U34268 (N_34268,N_25266,N_27447);
nand U34269 (N_34269,N_28566,N_25588);
xor U34270 (N_34270,N_25333,N_27649);
nor U34271 (N_34271,N_26101,N_25300);
nand U34272 (N_34272,N_26419,N_28861);
nand U34273 (N_34273,N_26196,N_27956);
nor U34274 (N_34274,N_25302,N_26793);
nor U34275 (N_34275,N_25428,N_29251);
and U34276 (N_34276,N_26520,N_25025);
or U34277 (N_34277,N_26376,N_27836);
nand U34278 (N_34278,N_26909,N_25244);
xor U34279 (N_34279,N_28453,N_29105);
and U34280 (N_34280,N_26993,N_26864);
nand U34281 (N_34281,N_26657,N_28039);
nor U34282 (N_34282,N_26599,N_27640);
and U34283 (N_34283,N_28695,N_28800);
nand U34284 (N_34284,N_27486,N_26589);
nor U34285 (N_34285,N_27852,N_29166);
nor U34286 (N_34286,N_29174,N_26855);
and U34287 (N_34287,N_29787,N_25237);
or U34288 (N_34288,N_28191,N_26913);
and U34289 (N_34289,N_29743,N_28952);
nor U34290 (N_34290,N_27971,N_27321);
nor U34291 (N_34291,N_29906,N_28347);
or U34292 (N_34292,N_26910,N_28724);
xnor U34293 (N_34293,N_27681,N_28620);
nand U34294 (N_34294,N_28562,N_26959);
or U34295 (N_34295,N_28168,N_27223);
xor U34296 (N_34296,N_29497,N_25594);
nor U34297 (N_34297,N_25990,N_25890);
and U34298 (N_34298,N_29531,N_29659);
and U34299 (N_34299,N_29796,N_29080);
nor U34300 (N_34300,N_28718,N_26689);
nor U34301 (N_34301,N_26794,N_29982);
xor U34302 (N_34302,N_26752,N_27604);
or U34303 (N_34303,N_29341,N_27221);
xnor U34304 (N_34304,N_27716,N_29845);
or U34305 (N_34305,N_28639,N_26911);
nor U34306 (N_34306,N_29197,N_28629);
nand U34307 (N_34307,N_26348,N_26975);
or U34308 (N_34308,N_28328,N_28445);
or U34309 (N_34309,N_28767,N_27413);
nor U34310 (N_34310,N_27718,N_27698);
xnor U34311 (N_34311,N_27278,N_26803);
nor U34312 (N_34312,N_25169,N_29029);
nor U34313 (N_34313,N_26773,N_26062);
and U34314 (N_34314,N_28463,N_29505);
nor U34315 (N_34315,N_27886,N_26365);
and U34316 (N_34316,N_27439,N_26257);
xnor U34317 (N_34317,N_25798,N_26851);
or U34318 (N_34318,N_27794,N_25729);
and U34319 (N_34319,N_28215,N_27884);
or U34320 (N_34320,N_27561,N_26128);
nor U34321 (N_34321,N_26822,N_29718);
or U34322 (N_34322,N_28521,N_26302);
nor U34323 (N_34323,N_27341,N_27513);
or U34324 (N_34324,N_29643,N_28646);
or U34325 (N_34325,N_26914,N_27200);
or U34326 (N_34326,N_25639,N_25812);
xnor U34327 (N_34327,N_29949,N_28354);
nor U34328 (N_34328,N_28996,N_29356);
and U34329 (N_34329,N_28850,N_28366);
nand U34330 (N_34330,N_27941,N_29227);
and U34331 (N_34331,N_29617,N_27519);
nand U34332 (N_34332,N_25491,N_25525);
and U34333 (N_34333,N_29116,N_29594);
or U34334 (N_34334,N_27619,N_27854);
and U34335 (N_34335,N_27587,N_25031);
or U34336 (N_34336,N_26438,N_27379);
xor U34337 (N_34337,N_26619,N_27079);
nor U34338 (N_34338,N_26647,N_29664);
nor U34339 (N_34339,N_29466,N_28362);
xnor U34340 (N_34340,N_28879,N_28397);
nor U34341 (N_34341,N_25302,N_28561);
nand U34342 (N_34342,N_27271,N_29098);
nand U34343 (N_34343,N_25059,N_29484);
or U34344 (N_34344,N_29284,N_26382);
nor U34345 (N_34345,N_29621,N_29022);
and U34346 (N_34346,N_29657,N_28549);
and U34347 (N_34347,N_29390,N_29681);
or U34348 (N_34348,N_29258,N_25233);
and U34349 (N_34349,N_26620,N_27151);
nand U34350 (N_34350,N_29996,N_25963);
nand U34351 (N_34351,N_26824,N_26061);
nor U34352 (N_34352,N_25675,N_25619);
nor U34353 (N_34353,N_28510,N_29995);
or U34354 (N_34354,N_28284,N_29313);
or U34355 (N_34355,N_27136,N_28584);
xor U34356 (N_34356,N_28469,N_28901);
nor U34357 (N_34357,N_26670,N_28894);
and U34358 (N_34358,N_25479,N_28799);
or U34359 (N_34359,N_28456,N_29632);
nand U34360 (N_34360,N_28899,N_25701);
or U34361 (N_34361,N_28736,N_25913);
and U34362 (N_34362,N_27394,N_27504);
xnor U34363 (N_34363,N_27972,N_26495);
or U34364 (N_34364,N_29904,N_26423);
or U34365 (N_34365,N_26620,N_27957);
nor U34366 (N_34366,N_27517,N_29265);
nand U34367 (N_34367,N_27834,N_29259);
and U34368 (N_34368,N_28881,N_27579);
xor U34369 (N_34369,N_27109,N_27048);
nand U34370 (N_34370,N_26500,N_27024);
and U34371 (N_34371,N_25615,N_25057);
or U34372 (N_34372,N_28081,N_26201);
xor U34373 (N_34373,N_29479,N_27904);
nand U34374 (N_34374,N_26546,N_28295);
nor U34375 (N_34375,N_25962,N_25231);
or U34376 (N_34376,N_28327,N_26377);
nor U34377 (N_34377,N_27060,N_26471);
nand U34378 (N_34378,N_29115,N_26433);
nor U34379 (N_34379,N_26676,N_29432);
and U34380 (N_34380,N_27100,N_26232);
or U34381 (N_34381,N_28830,N_26254);
nor U34382 (N_34382,N_25457,N_27040);
nor U34383 (N_34383,N_27417,N_29585);
xor U34384 (N_34384,N_26539,N_28151);
and U34385 (N_34385,N_29481,N_28585);
xnor U34386 (N_34386,N_29350,N_28586);
xnor U34387 (N_34387,N_29344,N_27897);
nand U34388 (N_34388,N_27775,N_27643);
or U34389 (N_34389,N_25734,N_28373);
nand U34390 (N_34390,N_28492,N_26132);
nand U34391 (N_34391,N_25845,N_25562);
nand U34392 (N_34392,N_29848,N_25849);
xor U34393 (N_34393,N_29833,N_27825);
nand U34394 (N_34394,N_26458,N_29446);
and U34395 (N_34395,N_27683,N_27771);
nand U34396 (N_34396,N_27790,N_29363);
or U34397 (N_34397,N_25129,N_26906);
and U34398 (N_34398,N_29886,N_27623);
and U34399 (N_34399,N_29963,N_28796);
nor U34400 (N_34400,N_29049,N_28258);
nand U34401 (N_34401,N_25509,N_25301);
nand U34402 (N_34402,N_28053,N_28775);
nand U34403 (N_34403,N_28289,N_29077);
or U34404 (N_34404,N_27612,N_28429);
nand U34405 (N_34405,N_27679,N_26650);
xor U34406 (N_34406,N_27439,N_29907);
nand U34407 (N_34407,N_27307,N_27499);
nand U34408 (N_34408,N_28647,N_29611);
nand U34409 (N_34409,N_26570,N_25607);
and U34410 (N_34410,N_27157,N_25353);
or U34411 (N_34411,N_25219,N_29065);
and U34412 (N_34412,N_29487,N_28424);
xor U34413 (N_34413,N_28354,N_25464);
nand U34414 (N_34414,N_27981,N_26933);
nor U34415 (N_34415,N_27181,N_29843);
nand U34416 (N_34416,N_29263,N_26461);
xor U34417 (N_34417,N_25283,N_29409);
nor U34418 (N_34418,N_26837,N_25689);
and U34419 (N_34419,N_28929,N_28621);
nand U34420 (N_34420,N_28579,N_28397);
nand U34421 (N_34421,N_28248,N_25554);
nor U34422 (N_34422,N_28865,N_26751);
or U34423 (N_34423,N_28134,N_27601);
nand U34424 (N_34424,N_27416,N_27462);
and U34425 (N_34425,N_25725,N_28262);
nand U34426 (N_34426,N_27507,N_27265);
xnor U34427 (N_34427,N_26565,N_25906);
xnor U34428 (N_34428,N_28093,N_25281);
xor U34429 (N_34429,N_25070,N_28203);
xnor U34430 (N_34430,N_25322,N_27173);
and U34431 (N_34431,N_26361,N_25912);
xor U34432 (N_34432,N_27240,N_25812);
nor U34433 (N_34433,N_29038,N_29014);
or U34434 (N_34434,N_26426,N_27719);
and U34435 (N_34435,N_28759,N_27076);
and U34436 (N_34436,N_26429,N_26921);
nand U34437 (N_34437,N_29729,N_25696);
xnor U34438 (N_34438,N_28568,N_29674);
nor U34439 (N_34439,N_28397,N_26040);
or U34440 (N_34440,N_29688,N_26450);
nand U34441 (N_34441,N_28590,N_29424);
xor U34442 (N_34442,N_26921,N_27081);
nor U34443 (N_34443,N_26487,N_27647);
nor U34444 (N_34444,N_25732,N_28565);
nand U34445 (N_34445,N_27493,N_26678);
xnor U34446 (N_34446,N_27561,N_29939);
nor U34447 (N_34447,N_26867,N_29374);
and U34448 (N_34448,N_27082,N_28695);
nand U34449 (N_34449,N_29002,N_26035);
nor U34450 (N_34450,N_26235,N_25514);
or U34451 (N_34451,N_25378,N_26775);
nor U34452 (N_34452,N_28505,N_26652);
nand U34453 (N_34453,N_27666,N_28360);
nor U34454 (N_34454,N_26547,N_28214);
or U34455 (N_34455,N_28884,N_26168);
nand U34456 (N_34456,N_29769,N_25860);
and U34457 (N_34457,N_29241,N_26390);
or U34458 (N_34458,N_27398,N_27607);
and U34459 (N_34459,N_28009,N_29950);
xor U34460 (N_34460,N_28587,N_26118);
and U34461 (N_34461,N_28918,N_25094);
or U34462 (N_34462,N_29135,N_26796);
or U34463 (N_34463,N_28280,N_25827);
and U34464 (N_34464,N_27654,N_25550);
xor U34465 (N_34465,N_25390,N_28244);
nand U34466 (N_34466,N_26035,N_25350);
nand U34467 (N_34467,N_25117,N_26408);
nand U34468 (N_34468,N_27260,N_27657);
xor U34469 (N_34469,N_29610,N_25182);
xor U34470 (N_34470,N_28758,N_27852);
and U34471 (N_34471,N_26854,N_25592);
nand U34472 (N_34472,N_26259,N_25303);
nor U34473 (N_34473,N_27978,N_27137);
nor U34474 (N_34474,N_29942,N_29211);
nand U34475 (N_34475,N_25870,N_26306);
or U34476 (N_34476,N_29111,N_28673);
or U34477 (N_34477,N_26516,N_29221);
or U34478 (N_34478,N_28940,N_29104);
or U34479 (N_34479,N_25034,N_26751);
nor U34480 (N_34480,N_26838,N_25527);
nor U34481 (N_34481,N_28298,N_28192);
xnor U34482 (N_34482,N_29717,N_28577);
nand U34483 (N_34483,N_29992,N_29919);
xnor U34484 (N_34484,N_29830,N_29997);
nand U34485 (N_34485,N_29979,N_26715);
and U34486 (N_34486,N_27059,N_26973);
xnor U34487 (N_34487,N_26123,N_26965);
or U34488 (N_34488,N_29711,N_28217);
nand U34489 (N_34489,N_28014,N_26336);
nand U34490 (N_34490,N_29370,N_28921);
xnor U34491 (N_34491,N_25806,N_27005);
nand U34492 (N_34492,N_28184,N_26754);
nand U34493 (N_34493,N_27952,N_25249);
and U34494 (N_34494,N_26067,N_29870);
and U34495 (N_34495,N_28376,N_25547);
xnor U34496 (N_34496,N_25386,N_28121);
nand U34497 (N_34497,N_28413,N_29066);
and U34498 (N_34498,N_26917,N_25961);
nor U34499 (N_34499,N_26921,N_29247);
or U34500 (N_34500,N_28711,N_27543);
xor U34501 (N_34501,N_26123,N_25034);
and U34502 (N_34502,N_26955,N_29519);
and U34503 (N_34503,N_28575,N_28070);
nand U34504 (N_34504,N_25660,N_26660);
nand U34505 (N_34505,N_25473,N_25352);
nor U34506 (N_34506,N_29712,N_25317);
nand U34507 (N_34507,N_27591,N_25923);
nor U34508 (N_34508,N_26532,N_28396);
nand U34509 (N_34509,N_26684,N_25550);
nor U34510 (N_34510,N_26944,N_25808);
and U34511 (N_34511,N_27169,N_27854);
or U34512 (N_34512,N_27427,N_28025);
or U34513 (N_34513,N_28721,N_25366);
or U34514 (N_34514,N_25204,N_26991);
and U34515 (N_34515,N_26742,N_26757);
or U34516 (N_34516,N_25392,N_25862);
xor U34517 (N_34517,N_26793,N_28558);
nand U34518 (N_34518,N_28660,N_28917);
xnor U34519 (N_34519,N_29597,N_29642);
xor U34520 (N_34520,N_29974,N_27866);
or U34521 (N_34521,N_27485,N_28905);
and U34522 (N_34522,N_26265,N_26127);
nand U34523 (N_34523,N_26488,N_27106);
nand U34524 (N_34524,N_29932,N_28747);
and U34525 (N_34525,N_26482,N_26122);
nor U34526 (N_34526,N_25548,N_27607);
nand U34527 (N_34527,N_25470,N_25048);
nor U34528 (N_34528,N_27577,N_28330);
nand U34529 (N_34529,N_29543,N_25094);
nand U34530 (N_34530,N_25638,N_26663);
or U34531 (N_34531,N_28796,N_28897);
and U34532 (N_34532,N_29885,N_28360);
xor U34533 (N_34533,N_29479,N_29218);
xor U34534 (N_34534,N_27260,N_28031);
and U34535 (N_34535,N_26860,N_29667);
and U34536 (N_34536,N_27063,N_29703);
or U34537 (N_34537,N_29514,N_28299);
and U34538 (N_34538,N_25519,N_27364);
and U34539 (N_34539,N_26629,N_25407);
and U34540 (N_34540,N_29820,N_25869);
xor U34541 (N_34541,N_28551,N_26087);
and U34542 (N_34542,N_28053,N_29767);
xor U34543 (N_34543,N_27087,N_26760);
and U34544 (N_34544,N_27617,N_28253);
nor U34545 (N_34545,N_26937,N_27590);
nand U34546 (N_34546,N_29444,N_29456);
nor U34547 (N_34547,N_27022,N_26666);
xnor U34548 (N_34548,N_27934,N_28724);
nand U34549 (N_34549,N_29824,N_26046);
nand U34550 (N_34550,N_25916,N_27054);
nand U34551 (N_34551,N_27167,N_26498);
nand U34552 (N_34552,N_28400,N_26395);
or U34553 (N_34553,N_26491,N_28427);
nand U34554 (N_34554,N_25168,N_26791);
and U34555 (N_34555,N_29981,N_29655);
nand U34556 (N_34556,N_26486,N_27000);
or U34557 (N_34557,N_26578,N_29569);
xor U34558 (N_34558,N_29879,N_26152);
and U34559 (N_34559,N_25017,N_27615);
nor U34560 (N_34560,N_29535,N_29123);
or U34561 (N_34561,N_26192,N_28310);
nand U34562 (N_34562,N_25358,N_25909);
nand U34563 (N_34563,N_29315,N_25581);
and U34564 (N_34564,N_27273,N_26288);
xor U34565 (N_34565,N_26157,N_29233);
xor U34566 (N_34566,N_28270,N_27189);
or U34567 (N_34567,N_29027,N_28191);
or U34568 (N_34568,N_28842,N_29409);
nor U34569 (N_34569,N_29021,N_27221);
xnor U34570 (N_34570,N_29805,N_28689);
or U34571 (N_34571,N_28717,N_26674);
nor U34572 (N_34572,N_28483,N_29678);
nand U34573 (N_34573,N_27181,N_26157);
xnor U34574 (N_34574,N_26069,N_28129);
and U34575 (N_34575,N_29005,N_29057);
and U34576 (N_34576,N_27612,N_29288);
and U34577 (N_34577,N_29214,N_28067);
nand U34578 (N_34578,N_27010,N_25783);
nor U34579 (N_34579,N_27109,N_29303);
or U34580 (N_34580,N_29444,N_29602);
xnor U34581 (N_34581,N_29638,N_28349);
xnor U34582 (N_34582,N_26424,N_28673);
and U34583 (N_34583,N_27175,N_27545);
nor U34584 (N_34584,N_27689,N_29432);
xor U34585 (N_34585,N_26345,N_29858);
and U34586 (N_34586,N_27211,N_25438);
nor U34587 (N_34587,N_28252,N_29585);
xor U34588 (N_34588,N_28796,N_28575);
xor U34589 (N_34589,N_26226,N_29287);
xor U34590 (N_34590,N_26682,N_26280);
xor U34591 (N_34591,N_26684,N_28981);
nor U34592 (N_34592,N_28729,N_25900);
or U34593 (N_34593,N_28253,N_25236);
and U34594 (N_34594,N_27639,N_27024);
nand U34595 (N_34595,N_28652,N_26208);
or U34596 (N_34596,N_26350,N_28846);
xnor U34597 (N_34597,N_29560,N_29506);
or U34598 (N_34598,N_27865,N_27643);
and U34599 (N_34599,N_28416,N_28118);
or U34600 (N_34600,N_25058,N_28485);
nor U34601 (N_34601,N_29313,N_27912);
nor U34602 (N_34602,N_26966,N_29376);
or U34603 (N_34603,N_27218,N_28655);
and U34604 (N_34604,N_27949,N_26083);
and U34605 (N_34605,N_29493,N_26256);
nand U34606 (N_34606,N_29860,N_27358);
nand U34607 (N_34607,N_27702,N_26794);
nor U34608 (N_34608,N_29176,N_29857);
or U34609 (N_34609,N_27539,N_27466);
or U34610 (N_34610,N_25417,N_29270);
and U34611 (N_34611,N_25236,N_28050);
nand U34612 (N_34612,N_25267,N_28036);
nand U34613 (N_34613,N_27882,N_26996);
xor U34614 (N_34614,N_26155,N_26423);
and U34615 (N_34615,N_28757,N_26406);
and U34616 (N_34616,N_27461,N_28431);
xnor U34617 (N_34617,N_28636,N_26360);
xor U34618 (N_34618,N_28306,N_28481);
or U34619 (N_34619,N_28936,N_27321);
nand U34620 (N_34620,N_26584,N_25526);
and U34621 (N_34621,N_26110,N_28109);
and U34622 (N_34622,N_29268,N_26294);
xor U34623 (N_34623,N_28285,N_28037);
and U34624 (N_34624,N_28194,N_26968);
xor U34625 (N_34625,N_25712,N_25020);
xnor U34626 (N_34626,N_26898,N_27967);
nand U34627 (N_34627,N_27734,N_27236);
nand U34628 (N_34628,N_25092,N_26083);
xor U34629 (N_34629,N_28348,N_25456);
and U34630 (N_34630,N_26998,N_29570);
nor U34631 (N_34631,N_25154,N_27733);
and U34632 (N_34632,N_29449,N_29489);
nor U34633 (N_34633,N_26210,N_25166);
nor U34634 (N_34634,N_27219,N_25155);
and U34635 (N_34635,N_26061,N_26285);
nor U34636 (N_34636,N_25307,N_25340);
or U34637 (N_34637,N_26829,N_27423);
nor U34638 (N_34638,N_26755,N_28901);
xor U34639 (N_34639,N_26146,N_25029);
xnor U34640 (N_34640,N_25537,N_26369);
and U34641 (N_34641,N_26454,N_29927);
and U34642 (N_34642,N_26921,N_26092);
nor U34643 (N_34643,N_25763,N_28013);
or U34644 (N_34644,N_26689,N_26387);
nor U34645 (N_34645,N_27620,N_29882);
and U34646 (N_34646,N_27372,N_27510);
or U34647 (N_34647,N_26756,N_26864);
xnor U34648 (N_34648,N_28691,N_26978);
or U34649 (N_34649,N_27245,N_25004);
nor U34650 (N_34650,N_26186,N_26792);
and U34651 (N_34651,N_25263,N_28560);
or U34652 (N_34652,N_25013,N_28811);
nand U34653 (N_34653,N_29384,N_27623);
or U34654 (N_34654,N_27990,N_26760);
nor U34655 (N_34655,N_27591,N_25899);
and U34656 (N_34656,N_26726,N_25995);
and U34657 (N_34657,N_26903,N_27716);
nor U34658 (N_34658,N_28450,N_27855);
nor U34659 (N_34659,N_28684,N_28288);
and U34660 (N_34660,N_28867,N_27784);
nand U34661 (N_34661,N_25231,N_26309);
and U34662 (N_34662,N_25471,N_25283);
xnor U34663 (N_34663,N_26859,N_28553);
and U34664 (N_34664,N_25502,N_29998);
or U34665 (N_34665,N_26465,N_29687);
nor U34666 (N_34666,N_29144,N_26959);
xor U34667 (N_34667,N_28419,N_25006);
or U34668 (N_34668,N_28956,N_25777);
and U34669 (N_34669,N_25900,N_29318);
and U34670 (N_34670,N_26204,N_27089);
or U34671 (N_34671,N_27129,N_27792);
and U34672 (N_34672,N_28647,N_28071);
nand U34673 (N_34673,N_26189,N_28519);
nor U34674 (N_34674,N_28291,N_29565);
nor U34675 (N_34675,N_28437,N_29942);
nand U34676 (N_34676,N_25144,N_26208);
nand U34677 (N_34677,N_27567,N_26674);
xor U34678 (N_34678,N_26416,N_26368);
nand U34679 (N_34679,N_25229,N_29739);
nand U34680 (N_34680,N_27703,N_26071);
or U34681 (N_34681,N_28281,N_29224);
xor U34682 (N_34682,N_27400,N_25200);
or U34683 (N_34683,N_29901,N_25820);
or U34684 (N_34684,N_26961,N_28108);
or U34685 (N_34685,N_29140,N_25482);
nor U34686 (N_34686,N_29431,N_29683);
xor U34687 (N_34687,N_26911,N_27380);
nor U34688 (N_34688,N_27415,N_29494);
and U34689 (N_34689,N_27177,N_29785);
and U34690 (N_34690,N_28379,N_26382);
or U34691 (N_34691,N_27589,N_25098);
nand U34692 (N_34692,N_28084,N_27201);
and U34693 (N_34693,N_26995,N_25705);
xnor U34694 (N_34694,N_25587,N_25172);
nor U34695 (N_34695,N_29114,N_25654);
xor U34696 (N_34696,N_25039,N_27296);
and U34697 (N_34697,N_27067,N_26690);
nor U34698 (N_34698,N_27570,N_29635);
or U34699 (N_34699,N_29546,N_25439);
nand U34700 (N_34700,N_26526,N_26395);
or U34701 (N_34701,N_25120,N_26343);
nand U34702 (N_34702,N_25626,N_29487);
and U34703 (N_34703,N_29454,N_27298);
or U34704 (N_34704,N_26012,N_26781);
or U34705 (N_34705,N_29717,N_25976);
or U34706 (N_34706,N_27513,N_26386);
xnor U34707 (N_34707,N_28844,N_28218);
and U34708 (N_34708,N_27773,N_29183);
nor U34709 (N_34709,N_28082,N_29083);
or U34710 (N_34710,N_26212,N_27273);
nand U34711 (N_34711,N_25193,N_26388);
xnor U34712 (N_34712,N_28749,N_26926);
or U34713 (N_34713,N_29491,N_25971);
or U34714 (N_34714,N_25364,N_27156);
nand U34715 (N_34715,N_28527,N_27670);
nor U34716 (N_34716,N_27632,N_26802);
or U34717 (N_34717,N_29178,N_29284);
xor U34718 (N_34718,N_28986,N_28576);
and U34719 (N_34719,N_28292,N_25044);
nor U34720 (N_34720,N_27896,N_29792);
or U34721 (N_34721,N_29958,N_25250);
nor U34722 (N_34722,N_25015,N_26016);
nand U34723 (N_34723,N_26947,N_26625);
and U34724 (N_34724,N_26494,N_29230);
and U34725 (N_34725,N_26706,N_27326);
or U34726 (N_34726,N_29998,N_26795);
nand U34727 (N_34727,N_26684,N_28561);
and U34728 (N_34728,N_27121,N_29059);
nand U34729 (N_34729,N_28722,N_29656);
and U34730 (N_34730,N_25239,N_25701);
nand U34731 (N_34731,N_29764,N_28789);
and U34732 (N_34732,N_25453,N_28540);
nor U34733 (N_34733,N_29590,N_28943);
or U34734 (N_34734,N_25761,N_27267);
and U34735 (N_34735,N_26483,N_29963);
or U34736 (N_34736,N_29301,N_25300);
and U34737 (N_34737,N_26641,N_25367);
xnor U34738 (N_34738,N_27250,N_26810);
xnor U34739 (N_34739,N_26639,N_28749);
xnor U34740 (N_34740,N_27986,N_28953);
nor U34741 (N_34741,N_26682,N_29368);
nor U34742 (N_34742,N_28818,N_29997);
nand U34743 (N_34743,N_26379,N_27488);
nor U34744 (N_34744,N_26864,N_25509);
xnor U34745 (N_34745,N_28358,N_27254);
and U34746 (N_34746,N_25281,N_29061);
nand U34747 (N_34747,N_28816,N_27999);
or U34748 (N_34748,N_25696,N_25599);
xnor U34749 (N_34749,N_27905,N_27125);
xor U34750 (N_34750,N_25124,N_27348);
xor U34751 (N_34751,N_26391,N_26969);
or U34752 (N_34752,N_29707,N_25735);
and U34753 (N_34753,N_27158,N_29131);
nor U34754 (N_34754,N_29039,N_28765);
nand U34755 (N_34755,N_28234,N_25068);
nand U34756 (N_34756,N_26715,N_29840);
xnor U34757 (N_34757,N_29210,N_25794);
nand U34758 (N_34758,N_27282,N_29854);
nand U34759 (N_34759,N_25929,N_28585);
nor U34760 (N_34760,N_29099,N_27208);
nor U34761 (N_34761,N_26621,N_25270);
xor U34762 (N_34762,N_25165,N_29411);
or U34763 (N_34763,N_25690,N_25765);
nand U34764 (N_34764,N_27986,N_28484);
nor U34765 (N_34765,N_26470,N_26719);
nand U34766 (N_34766,N_26433,N_25912);
nand U34767 (N_34767,N_25642,N_25384);
and U34768 (N_34768,N_26239,N_26805);
or U34769 (N_34769,N_25284,N_27501);
xor U34770 (N_34770,N_25031,N_29685);
and U34771 (N_34771,N_25004,N_28558);
nand U34772 (N_34772,N_26403,N_28315);
and U34773 (N_34773,N_25642,N_26369);
nand U34774 (N_34774,N_25376,N_28074);
nor U34775 (N_34775,N_28155,N_28736);
xor U34776 (N_34776,N_29180,N_25514);
nand U34777 (N_34777,N_25697,N_25131);
or U34778 (N_34778,N_25792,N_29826);
nand U34779 (N_34779,N_26001,N_26943);
xnor U34780 (N_34780,N_29268,N_28334);
nor U34781 (N_34781,N_27265,N_29129);
nand U34782 (N_34782,N_27247,N_28074);
or U34783 (N_34783,N_29812,N_27298);
nand U34784 (N_34784,N_29049,N_25159);
and U34785 (N_34785,N_27102,N_28866);
xnor U34786 (N_34786,N_29193,N_28675);
and U34787 (N_34787,N_26003,N_25409);
xnor U34788 (N_34788,N_25212,N_28405);
and U34789 (N_34789,N_26937,N_25262);
and U34790 (N_34790,N_25357,N_27422);
or U34791 (N_34791,N_25376,N_26947);
or U34792 (N_34792,N_28581,N_28721);
nor U34793 (N_34793,N_25225,N_26410);
xor U34794 (N_34794,N_27121,N_26728);
nor U34795 (N_34795,N_26898,N_26037);
xor U34796 (N_34796,N_25294,N_25843);
xor U34797 (N_34797,N_27205,N_27594);
or U34798 (N_34798,N_25593,N_27682);
nand U34799 (N_34799,N_26168,N_29154);
nor U34800 (N_34800,N_25047,N_25916);
and U34801 (N_34801,N_29294,N_27768);
xnor U34802 (N_34802,N_25219,N_27039);
nand U34803 (N_34803,N_29714,N_29132);
or U34804 (N_34804,N_25821,N_28084);
or U34805 (N_34805,N_29175,N_29863);
nand U34806 (N_34806,N_29704,N_25688);
and U34807 (N_34807,N_29330,N_28727);
xor U34808 (N_34808,N_25283,N_26297);
nor U34809 (N_34809,N_26274,N_28667);
nand U34810 (N_34810,N_28875,N_29900);
xnor U34811 (N_34811,N_28394,N_28196);
xnor U34812 (N_34812,N_26937,N_26825);
xnor U34813 (N_34813,N_29616,N_26815);
or U34814 (N_34814,N_27813,N_26921);
and U34815 (N_34815,N_26092,N_29073);
or U34816 (N_34816,N_27273,N_25392);
nor U34817 (N_34817,N_25805,N_28608);
nand U34818 (N_34818,N_25895,N_25893);
and U34819 (N_34819,N_27027,N_25813);
or U34820 (N_34820,N_27753,N_27776);
or U34821 (N_34821,N_29567,N_29939);
nor U34822 (N_34822,N_25922,N_29193);
xor U34823 (N_34823,N_26413,N_25771);
or U34824 (N_34824,N_27406,N_25105);
or U34825 (N_34825,N_27688,N_29316);
and U34826 (N_34826,N_25337,N_28603);
nand U34827 (N_34827,N_29091,N_26864);
xor U34828 (N_34828,N_28128,N_28522);
nand U34829 (N_34829,N_25532,N_29993);
xnor U34830 (N_34830,N_25036,N_28112);
nand U34831 (N_34831,N_27954,N_26589);
nand U34832 (N_34832,N_26789,N_25618);
nand U34833 (N_34833,N_28604,N_28440);
nor U34834 (N_34834,N_28013,N_29731);
nand U34835 (N_34835,N_28807,N_25469);
xnor U34836 (N_34836,N_26521,N_25629);
nand U34837 (N_34837,N_27950,N_29220);
or U34838 (N_34838,N_25853,N_26700);
nand U34839 (N_34839,N_29386,N_25971);
nand U34840 (N_34840,N_29086,N_26886);
or U34841 (N_34841,N_25813,N_27394);
and U34842 (N_34842,N_29225,N_25760);
xnor U34843 (N_34843,N_26969,N_26752);
or U34844 (N_34844,N_29496,N_25142);
nand U34845 (N_34845,N_26358,N_25735);
or U34846 (N_34846,N_28531,N_28155);
xnor U34847 (N_34847,N_26190,N_28461);
nor U34848 (N_34848,N_28641,N_29149);
xnor U34849 (N_34849,N_25441,N_27710);
or U34850 (N_34850,N_29559,N_29233);
or U34851 (N_34851,N_25285,N_28415);
xnor U34852 (N_34852,N_28815,N_25957);
or U34853 (N_34853,N_29553,N_28084);
nand U34854 (N_34854,N_29342,N_28609);
and U34855 (N_34855,N_26726,N_28700);
xnor U34856 (N_34856,N_27071,N_27931);
or U34857 (N_34857,N_28720,N_28785);
nand U34858 (N_34858,N_28380,N_26414);
nor U34859 (N_34859,N_27793,N_25883);
nand U34860 (N_34860,N_27289,N_26283);
nand U34861 (N_34861,N_29452,N_28982);
and U34862 (N_34862,N_28875,N_27846);
xnor U34863 (N_34863,N_26072,N_26068);
or U34864 (N_34864,N_29605,N_28487);
or U34865 (N_34865,N_28385,N_26673);
nand U34866 (N_34866,N_26702,N_28378);
or U34867 (N_34867,N_29728,N_29503);
and U34868 (N_34868,N_29061,N_28463);
nand U34869 (N_34869,N_29985,N_25512);
or U34870 (N_34870,N_27883,N_26426);
nand U34871 (N_34871,N_29708,N_27443);
or U34872 (N_34872,N_29757,N_26381);
xor U34873 (N_34873,N_29715,N_29158);
nand U34874 (N_34874,N_27699,N_25493);
nand U34875 (N_34875,N_26911,N_25362);
or U34876 (N_34876,N_25261,N_28364);
or U34877 (N_34877,N_28189,N_28264);
nor U34878 (N_34878,N_27114,N_26937);
or U34879 (N_34879,N_28729,N_26959);
xnor U34880 (N_34880,N_29304,N_29633);
nor U34881 (N_34881,N_26152,N_27309);
or U34882 (N_34882,N_26592,N_27014);
xnor U34883 (N_34883,N_28791,N_26837);
nor U34884 (N_34884,N_27367,N_25449);
and U34885 (N_34885,N_29097,N_28080);
or U34886 (N_34886,N_26199,N_25652);
xor U34887 (N_34887,N_26124,N_28581);
nor U34888 (N_34888,N_28687,N_25109);
nand U34889 (N_34889,N_28852,N_29704);
and U34890 (N_34890,N_27506,N_25107);
xor U34891 (N_34891,N_27177,N_25839);
nand U34892 (N_34892,N_26301,N_26533);
xor U34893 (N_34893,N_27247,N_25483);
or U34894 (N_34894,N_26323,N_26885);
nand U34895 (N_34895,N_27382,N_26337);
or U34896 (N_34896,N_25019,N_25876);
nor U34897 (N_34897,N_28992,N_29890);
and U34898 (N_34898,N_25479,N_25650);
or U34899 (N_34899,N_28445,N_25334);
xnor U34900 (N_34900,N_29764,N_25359);
nor U34901 (N_34901,N_25675,N_27127);
and U34902 (N_34902,N_26197,N_28971);
nor U34903 (N_34903,N_25374,N_29501);
and U34904 (N_34904,N_27389,N_25928);
nand U34905 (N_34905,N_29733,N_25796);
and U34906 (N_34906,N_28366,N_28487);
and U34907 (N_34907,N_29393,N_27484);
nand U34908 (N_34908,N_28235,N_27012);
xor U34909 (N_34909,N_27863,N_26612);
nand U34910 (N_34910,N_25616,N_29173);
xor U34911 (N_34911,N_27776,N_28169);
nor U34912 (N_34912,N_26015,N_26384);
nor U34913 (N_34913,N_29869,N_26473);
and U34914 (N_34914,N_25482,N_25582);
or U34915 (N_34915,N_25081,N_25048);
nand U34916 (N_34916,N_29996,N_29859);
nor U34917 (N_34917,N_27637,N_25439);
nor U34918 (N_34918,N_26694,N_29230);
or U34919 (N_34919,N_28094,N_29916);
xor U34920 (N_34920,N_25562,N_26001);
xor U34921 (N_34921,N_28906,N_29712);
nor U34922 (N_34922,N_27802,N_25393);
xor U34923 (N_34923,N_26356,N_27096);
nand U34924 (N_34924,N_27896,N_28385);
or U34925 (N_34925,N_27269,N_27691);
or U34926 (N_34926,N_26948,N_25023);
xnor U34927 (N_34927,N_26187,N_28266);
xnor U34928 (N_34928,N_29953,N_25011);
or U34929 (N_34929,N_29842,N_29079);
nand U34930 (N_34930,N_26843,N_27863);
or U34931 (N_34931,N_28089,N_27500);
and U34932 (N_34932,N_25311,N_28545);
and U34933 (N_34933,N_27464,N_27764);
nand U34934 (N_34934,N_27725,N_26877);
nor U34935 (N_34935,N_26811,N_25620);
and U34936 (N_34936,N_29510,N_27258);
nor U34937 (N_34937,N_26125,N_25346);
nand U34938 (N_34938,N_27389,N_29324);
or U34939 (N_34939,N_28081,N_27642);
xnor U34940 (N_34940,N_26488,N_25457);
xor U34941 (N_34941,N_27835,N_27066);
or U34942 (N_34942,N_29480,N_29496);
nand U34943 (N_34943,N_25908,N_28550);
nand U34944 (N_34944,N_25021,N_28726);
and U34945 (N_34945,N_29966,N_28163);
xor U34946 (N_34946,N_25314,N_28861);
nand U34947 (N_34947,N_28727,N_28718);
nor U34948 (N_34948,N_28953,N_25793);
nand U34949 (N_34949,N_29522,N_26560);
nor U34950 (N_34950,N_27221,N_26903);
or U34951 (N_34951,N_26270,N_29222);
or U34952 (N_34952,N_28766,N_26984);
xnor U34953 (N_34953,N_25177,N_25829);
and U34954 (N_34954,N_29143,N_26386);
or U34955 (N_34955,N_29102,N_26887);
nand U34956 (N_34956,N_29380,N_29130);
xnor U34957 (N_34957,N_28306,N_28927);
xnor U34958 (N_34958,N_25955,N_29303);
xnor U34959 (N_34959,N_29913,N_27156);
nand U34960 (N_34960,N_28732,N_26859);
nand U34961 (N_34961,N_27223,N_27956);
or U34962 (N_34962,N_29974,N_26911);
and U34963 (N_34963,N_26105,N_28505);
or U34964 (N_34964,N_28959,N_29795);
or U34965 (N_34965,N_25312,N_25732);
and U34966 (N_34966,N_29417,N_26312);
or U34967 (N_34967,N_25115,N_26127);
xor U34968 (N_34968,N_29339,N_27426);
and U34969 (N_34969,N_28818,N_28455);
or U34970 (N_34970,N_28466,N_27074);
nor U34971 (N_34971,N_25903,N_25171);
or U34972 (N_34972,N_27326,N_25429);
or U34973 (N_34973,N_26723,N_25968);
nand U34974 (N_34974,N_27737,N_26000);
xnor U34975 (N_34975,N_29246,N_25535);
xor U34976 (N_34976,N_26655,N_28870);
xnor U34977 (N_34977,N_27125,N_29094);
nand U34978 (N_34978,N_26820,N_28984);
nor U34979 (N_34979,N_28000,N_25299);
and U34980 (N_34980,N_27725,N_27297);
and U34981 (N_34981,N_28096,N_25182);
xor U34982 (N_34982,N_29592,N_29084);
and U34983 (N_34983,N_29283,N_28112);
xnor U34984 (N_34984,N_28958,N_28625);
and U34985 (N_34985,N_27133,N_25897);
and U34986 (N_34986,N_25415,N_29373);
and U34987 (N_34987,N_26989,N_26234);
or U34988 (N_34988,N_28460,N_27339);
nor U34989 (N_34989,N_25600,N_27643);
nor U34990 (N_34990,N_28125,N_26048);
nor U34991 (N_34991,N_29590,N_27681);
xor U34992 (N_34992,N_25294,N_28654);
nor U34993 (N_34993,N_29001,N_27492);
and U34994 (N_34994,N_29463,N_29158);
or U34995 (N_34995,N_28085,N_26295);
and U34996 (N_34996,N_28052,N_28208);
xnor U34997 (N_34997,N_29483,N_29423);
nand U34998 (N_34998,N_29592,N_27060);
nor U34999 (N_34999,N_26283,N_26915);
nand U35000 (N_35000,N_31809,N_32629);
and U35001 (N_35001,N_32611,N_30928);
and U35002 (N_35002,N_33447,N_31287);
nand U35003 (N_35003,N_32441,N_31763);
xnor U35004 (N_35004,N_34292,N_30404);
xor U35005 (N_35005,N_34273,N_32677);
nor U35006 (N_35006,N_32192,N_34154);
xnor U35007 (N_35007,N_33579,N_31930);
and U35008 (N_35008,N_31300,N_34975);
nand U35009 (N_35009,N_32094,N_31887);
and U35010 (N_35010,N_34822,N_34969);
xor U35011 (N_35011,N_34918,N_34493);
and U35012 (N_35012,N_33305,N_31546);
and U35013 (N_35013,N_32656,N_32514);
nor U35014 (N_35014,N_30351,N_32168);
or U35015 (N_35015,N_30844,N_32221);
xnor U35016 (N_35016,N_31535,N_33300);
nand U35017 (N_35017,N_33753,N_33090);
nand U35018 (N_35018,N_33100,N_30623);
and U35019 (N_35019,N_33866,N_32775);
nand U35020 (N_35020,N_33429,N_32619);
or U35021 (N_35021,N_34590,N_32551);
nor U35022 (N_35022,N_30538,N_32240);
nand U35023 (N_35023,N_32031,N_31601);
or U35024 (N_35024,N_31259,N_31405);
or U35025 (N_35025,N_34520,N_33682);
and U35026 (N_35026,N_33697,N_33520);
xnor U35027 (N_35027,N_33063,N_33928);
or U35028 (N_35028,N_33835,N_31329);
nand U35029 (N_35029,N_32155,N_33119);
or U35030 (N_35030,N_31309,N_33455);
and U35031 (N_35031,N_31162,N_33553);
and U35032 (N_35032,N_32285,N_31109);
and U35033 (N_35033,N_32257,N_30205);
and U35034 (N_35034,N_32274,N_33561);
and U35035 (N_35035,N_31787,N_34882);
or U35036 (N_35036,N_31308,N_32365);
nor U35037 (N_35037,N_30174,N_30172);
nand U35038 (N_35038,N_30298,N_30143);
and U35039 (N_35039,N_30246,N_34037);
or U35040 (N_35040,N_34962,N_34106);
xor U35041 (N_35041,N_30515,N_34824);
nor U35042 (N_35042,N_33730,N_31739);
nand U35043 (N_35043,N_33062,N_31650);
or U35044 (N_35044,N_32742,N_30560);
or U35045 (N_35045,N_33482,N_30308);
nor U35046 (N_35046,N_33596,N_32975);
nor U35047 (N_35047,N_30390,N_31592);
xor U35048 (N_35048,N_33360,N_30652);
nor U35049 (N_35049,N_30954,N_34613);
nor U35050 (N_35050,N_33277,N_30929);
or U35051 (N_35051,N_30516,N_30050);
or U35052 (N_35052,N_32889,N_30433);
or U35053 (N_35053,N_33694,N_32023);
xnor U35054 (N_35054,N_32994,N_30407);
and U35055 (N_35055,N_31578,N_33160);
xor U35056 (N_35056,N_30613,N_33196);
and U35057 (N_35057,N_32260,N_33485);
xor U35058 (N_35058,N_31868,N_33871);
and U35059 (N_35059,N_34038,N_30912);
or U35060 (N_35060,N_33860,N_32186);
and U35061 (N_35061,N_33939,N_30987);
and U35062 (N_35062,N_34198,N_34617);
or U35063 (N_35063,N_34470,N_32877);
nand U35064 (N_35064,N_33911,N_31819);
xnor U35065 (N_35065,N_31937,N_34259);
or U35066 (N_35066,N_30070,N_33110);
or U35067 (N_35067,N_33782,N_33749);
or U35068 (N_35068,N_30672,N_31146);
or U35069 (N_35069,N_34475,N_33088);
nand U35070 (N_35070,N_32277,N_30425);
and U35071 (N_35071,N_30804,N_34502);
xnor U35072 (N_35072,N_34145,N_31622);
nand U35073 (N_35073,N_33388,N_31929);
and U35074 (N_35074,N_34422,N_34924);
nor U35075 (N_35075,N_31290,N_30389);
xnor U35076 (N_35076,N_32208,N_33819);
nor U35077 (N_35077,N_34076,N_32663);
xor U35078 (N_35078,N_34832,N_31494);
xnor U35079 (N_35079,N_32683,N_30013);
or U35080 (N_35080,N_33622,N_33785);
and U35081 (N_35081,N_34088,N_31397);
nor U35082 (N_35082,N_31331,N_32738);
nor U35083 (N_35083,N_31782,N_32478);
nand U35084 (N_35084,N_32512,N_34441);
nand U35085 (N_35085,N_33635,N_30925);
nand U35086 (N_35086,N_30005,N_30948);
xnor U35087 (N_35087,N_31142,N_30150);
and U35088 (N_35088,N_30221,N_30583);
nor U35089 (N_35089,N_30773,N_31894);
nand U35090 (N_35090,N_34768,N_31282);
xnor U35091 (N_35091,N_30598,N_31338);
nand U35092 (N_35092,N_30331,N_32439);
nor U35093 (N_35093,N_33272,N_32727);
and U35094 (N_35094,N_32360,N_34277);
nand U35095 (N_35095,N_33258,N_32675);
nand U35096 (N_35096,N_31200,N_34036);
nand U35097 (N_35097,N_30417,N_32386);
nand U35098 (N_35098,N_31169,N_34188);
or U35099 (N_35099,N_33283,N_31970);
xor U35100 (N_35100,N_32645,N_34801);
and U35101 (N_35101,N_33981,N_30267);
and U35102 (N_35102,N_33483,N_34724);
xnor U35103 (N_35103,N_32550,N_32247);
nor U35104 (N_35104,N_34466,N_34726);
xnor U35105 (N_35105,N_31945,N_31516);
nor U35106 (N_35106,N_32284,N_30665);
and U35107 (N_35107,N_31611,N_30119);
and U35108 (N_35108,N_32488,N_32844);
nand U35109 (N_35109,N_31833,N_32556);
nand U35110 (N_35110,N_31831,N_30203);
nand U35111 (N_35111,N_30890,N_30805);
and U35112 (N_35112,N_30363,N_31860);
and U35113 (N_35113,N_33818,N_34226);
and U35114 (N_35114,N_31942,N_30812);
nor U35115 (N_35115,N_30060,N_34405);
and U35116 (N_35116,N_34925,N_32497);
and U35117 (N_35117,N_32463,N_30158);
nor U35118 (N_35118,N_33762,N_34351);
xnor U35119 (N_35119,N_32533,N_34522);
and U35120 (N_35120,N_30814,N_32128);
nor U35121 (N_35121,N_30061,N_30816);
and U35122 (N_35122,N_30400,N_31558);
nand U35123 (N_35123,N_33612,N_31264);
nand U35124 (N_35124,N_32548,N_32602);
or U35125 (N_35125,N_32138,N_32596);
nor U35126 (N_35126,N_34847,N_33045);
and U35127 (N_35127,N_33517,N_30002);
nand U35128 (N_35128,N_33965,N_34333);
nor U35129 (N_35129,N_34451,N_34641);
xnor U35130 (N_35130,N_34045,N_34015);
nor U35131 (N_35131,N_34958,N_32188);
xnor U35132 (N_35132,N_32754,N_30091);
and U35133 (N_35133,N_34521,N_34945);
nor U35134 (N_35134,N_30513,N_30201);
xnor U35135 (N_35135,N_32074,N_30887);
or U35136 (N_35136,N_32252,N_31968);
xor U35137 (N_35137,N_32189,N_33686);
xor U35138 (N_35138,N_34258,N_34800);
xnor U35139 (N_35139,N_32909,N_33542);
and U35140 (N_35140,N_34035,N_30946);
or U35141 (N_35141,N_31055,N_33729);
or U35142 (N_35142,N_32660,N_32587);
or U35143 (N_35143,N_33324,N_30018);
xor U35144 (N_35144,N_32067,N_34872);
nand U35145 (N_35145,N_31156,N_30615);
nor U35146 (N_35146,N_32964,N_34531);
or U35147 (N_35147,N_31458,N_32396);
nor U35148 (N_35148,N_34013,N_30901);
and U35149 (N_35149,N_34647,N_33732);
and U35150 (N_35150,N_32822,N_33329);
xnor U35151 (N_35151,N_34152,N_30690);
or U35152 (N_35152,N_33214,N_34063);
or U35153 (N_35153,N_30475,N_32993);
or U35154 (N_35154,N_30995,N_32011);
nor U35155 (N_35155,N_30811,N_32271);
or U35156 (N_35156,N_34803,N_32280);
or U35157 (N_35157,N_33232,N_32137);
or U35158 (N_35158,N_31112,N_32946);
nand U35159 (N_35159,N_30693,N_31852);
nor U35160 (N_35160,N_30155,N_32412);
nand U35161 (N_35161,N_32531,N_34762);
or U35162 (N_35162,N_32345,N_33592);
nand U35163 (N_35163,N_32076,N_34902);
xor U35164 (N_35164,N_33906,N_30786);
nand U35165 (N_35165,N_34562,N_32549);
nand U35166 (N_35166,N_31450,N_33278);
nand U35167 (N_35167,N_32979,N_32697);
nor U35168 (N_35168,N_33957,N_30486);
nand U35169 (N_35169,N_33216,N_32833);
or U35170 (N_35170,N_30129,N_34221);
nor U35171 (N_35171,N_31751,N_33771);
and U35172 (N_35172,N_30863,N_31354);
and U35173 (N_35173,N_33371,N_32084);
nand U35174 (N_35174,N_34862,N_30423);
and U35175 (N_35175,N_31198,N_31054);
and U35176 (N_35176,N_31445,N_32104);
nand U35177 (N_35177,N_32323,N_32491);
and U35178 (N_35178,N_33083,N_34247);
or U35179 (N_35179,N_30998,N_32576);
or U35180 (N_35180,N_31339,N_32714);
nand U35181 (N_35181,N_32025,N_30278);
or U35182 (N_35182,N_34491,N_33608);
or U35183 (N_35183,N_31661,N_33387);
nor U35184 (N_35184,N_31472,N_34948);
nand U35185 (N_35185,N_33041,N_30955);
nand U35186 (N_35186,N_32088,N_31949);
or U35187 (N_35187,N_32187,N_34190);
nand U35188 (N_35188,N_31663,N_33850);
nand U35189 (N_35189,N_31020,N_32499);
nand U35190 (N_35190,N_30491,N_31680);
nor U35191 (N_35191,N_30067,N_32091);
nand U35192 (N_35192,N_33321,N_31413);
nor U35193 (N_35193,N_32771,N_31486);
xnor U35194 (N_35194,N_33889,N_31891);
and U35195 (N_35195,N_32781,N_33423);
nor U35196 (N_35196,N_34121,N_32246);
nor U35197 (N_35197,N_33477,N_32292);
or U35198 (N_35198,N_30364,N_34537);
nand U35199 (N_35199,N_34608,N_32899);
nand U35200 (N_35200,N_34827,N_32935);
or U35201 (N_35201,N_34812,N_30800);
or U35202 (N_35202,N_30490,N_31051);
nor U35203 (N_35203,N_30778,N_31580);
nor U35204 (N_35204,N_33863,N_33385);
xor U35205 (N_35205,N_30052,N_31188);
nor U35206 (N_35206,N_33736,N_33969);
xnor U35207 (N_35207,N_31598,N_31226);
or U35208 (N_35208,N_31237,N_30165);
or U35209 (N_35209,N_30960,N_31377);
nor U35210 (N_35210,N_31798,N_31586);
xnor U35211 (N_35211,N_34795,N_31672);
nand U35212 (N_35212,N_33728,N_30611);
nor U35213 (N_35213,N_31597,N_34289);
nor U35214 (N_35214,N_34286,N_33313);
xor U35215 (N_35215,N_31492,N_31710);
and U35216 (N_35216,N_33851,N_32959);
and U35217 (N_35217,N_32476,N_33806);
nor U35218 (N_35218,N_31743,N_31952);
nor U35219 (N_35219,N_30958,N_33737);
or U35220 (N_35220,N_32062,N_34988);
xor U35221 (N_35221,N_34379,N_31336);
and U35222 (N_35222,N_33173,N_31858);
and U35223 (N_35223,N_34715,N_33039);
nand U35224 (N_35224,N_31562,N_30612);
xor U35225 (N_35225,N_33817,N_30862);
nand U35226 (N_35226,N_30677,N_32030);
nor U35227 (N_35227,N_32853,N_33759);
and U35228 (N_35228,N_31917,N_30893);
nor U35229 (N_35229,N_30149,N_33803);
nand U35230 (N_35230,N_30350,N_34850);
or U35231 (N_35231,N_30030,N_33439);
nand U35232 (N_35232,N_33607,N_32847);
nor U35233 (N_35233,N_33954,N_34771);
or U35234 (N_35234,N_34326,N_31697);
or U35235 (N_35235,N_34275,N_32862);
and U35236 (N_35236,N_34663,N_31871);
xor U35237 (N_35237,N_32466,N_33221);
nor U35238 (N_35238,N_33653,N_33362);
and U35239 (N_35239,N_33211,N_30460);
xor U35240 (N_35240,N_33812,N_33352);
nand U35241 (N_35241,N_31322,N_30875);
xor U35242 (N_35242,N_34027,N_33980);
xor U35243 (N_35243,N_32051,N_33531);
xor U35244 (N_35244,N_31699,N_33401);
and U35245 (N_35245,N_32696,N_30401);
nand U35246 (N_35246,N_32779,N_30905);
nand U35247 (N_35247,N_33340,N_33500);
xnor U35248 (N_35248,N_34888,N_33799);
nor U35249 (N_35249,N_32881,N_32150);
or U35250 (N_35250,N_30093,N_32799);
nor U35251 (N_35251,N_33733,N_32376);
nor U35252 (N_35252,N_30430,N_31623);
nor U35253 (N_35253,N_33109,N_34581);
or U35254 (N_35254,N_33696,N_31178);
xor U35255 (N_35255,N_34923,N_30621);
xor U35256 (N_35256,N_33113,N_34806);
and U35257 (N_35257,N_30906,N_34807);
and U35258 (N_35258,N_34560,N_32393);
nand U35259 (N_35259,N_33346,N_31713);
or U35260 (N_35260,N_31490,N_33797);
nand U35261 (N_35261,N_30510,N_34165);
or U35262 (N_35262,N_32564,N_30418);
and U35263 (N_35263,N_30157,N_34965);
nand U35264 (N_35264,N_31607,N_30855);
and U35265 (N_35265,N_30802,N_34352);
nand U35266 (N_35266,N_32748,N_34587);
nor U35267 (N_35267,N_31618,N_33238);
and U35268 (N_35268,N_33882,N_33049);
xor U35269 (N_35269,N_31217,N_33183);
nor U35270 (N_35270,N_34479,N_30708);
xnor U35271 (N_35271,N_30739,N_32566);
or U35272 (N_35272,N_30818,N_30674);
and U35273 (N_35273,N_31962,N_34625);
nor U35274 (N_35274,N_32504,N_31848);
nand U35275 (N_35275,N_34687,N_34950);
or U35276 (N_35276,N_33567,N_30003);
or U35277 (N_35277,N_34779,N_34483);
nor U35278 (N_35278,N_32267,N_33804);
and U35279 (N_35279,N_31006,N_31124);
and U35280 (N_35280,N_33986,N_33073);
nor U35281 (N_35281,N_33847,N_31117);
and U35282 (N_35282,N_32012,N_33916);
and U35283 (N_35283,N_30074,N_34453);
nand U35284 (N_35284,N_32965,N_34369);
nand U35285 (N_35285,N_30085,N_32140);
nand U35286 (N_35286,N_34998,N_32015);
and U35287 (N_35287,N_33564,N_30156);
xnor U35288 (N_35288,N_34672,N_30537);
and U35289 (N_35289,N_34298,N_34769);
and U35290 (N_35290,N_33393,N_33489);
nand U35291 (N_35291,N_30329,N_34095);
or U35292 (N_35292,N_34317,N_32958);
or U35293 (N_35293,N_30324,N_33524);
nor U35294 (N_35294,N_32654,N_30294);
nand U35295 (N_35295,N_33067,N_34244);
and U35296 (N_35296,N_32179,N_30362);
nor U35297 (N_35297,N_31934,N_30315);
nor U35298 (N_35298,N_30675,N_30380);
nor U35299 (N_35299,N_34423,N_30343);
xnor U35300 (N_35300,N_34336,N_33727);
or U35301 (N_35301,N_30924,N_32956);
or U35302 (N_35302,N_30916,N_31517);
and U35303 (N_35303,N_34571,N_31368);
xor U35304 (N_35304,N_32124,N_32373);
or U35305 (N_35305,N_33287,N_34178);
nor U35306 (N_35306,N_30618,N_30581);
nor U35307 (N_35307,N_34770,N_31267);
xor U35308 (N_35308,N_31875,N_33055);
nor U35309 (N_35309,N_33478,N_32927);
xnor U35310 (N_35310,N_33501,N_30026);
or U35311 (N_35311,N_32133,N_33950);
xor U35312 (N_35312,N_32657,N_30171);
and U35313 (N_35313,N_32642,N_34424);
or U35314 (N_35314,N_32529,N_31231);
or U35315 (N_35315,N_31983,N_30597);
or U35316 (N_35316,N_34390,N_34930);
nor U35317 (N_35317,N_32195,N_34767);
or U35318 (N_35318,N_34912,N_31959);
nor U35319 (N_35319,N_32871,N_34506);
nor U35320 (N_35320,N_31495,N_30388);
xnor U35321 (N_35321,N_32756,N_32686);
or U35322 (N_35322,N_33901,N_31118);
xor U35323 (N_35323,N_30162,N_33974);
and U35324 (N_35324,N_32403,N_33035);
nand U35325 (N_35325,N_30703,N_34223);
or U35326 (N_35326,N_32778,N_32142);
and U35327 (N_35327,N_32759,N_30402);
and U35328 (N_35328,N_32008,N_31230);
and U35329 (N_35329,N_30545,N_30572);
nand U35330 (N_35330,N_33096,N_31512);
xnor U35331 (N_35331,N_30626,N_34738);
xor U35332 (N_35332,N_30034,N_32043);
xor U35333 (N_35333,N_30752,N_31053);
nand U35334 (N_35334,N_32082,N_31480);
xnor U35335 (N_35335,N_32467,N_34661);
or U35336 (N_35336,N_30188,N_34266);
nor U35337 (N_35337,N_34659,N_31366);
nor U35338 (N_35338,N_33662,N_34146);
nand U35339 (N_35339,N_32215,N_34337);
xnor U35340 (N_35340,N_31134,N_34341);
nor U35341 (N_35341,N_34429,N_31295);
or U35342 (N_35342,N_30967,N_31463);
nand U35343 (N_35343,N_30857,N_34848);
or U35344 (N_35344,N_33495,N_30250);
xnor U35345 (N_35345,N_33222,N_34340);
nand U35346 (N_35346,N_30696,N_31206);
or U35347 (N_35347,N_33141,N_33552);
nor U35348 (N_35348,N_33563,N_34355);
xnor U35349 (N_35349,N_30121,N_33359);
or U35350 (N_35350,N_32814,N_34380);
nand U35351 (N_35351,N_32745,N_30706);
and U35352 (N_35352,N_34071,N_33040);
or U35353 (N_35353,N_34682,N_32315);
and U35354 (N_35354,N_31742,N_31341);
nor U35355 (N_35355,N_32262,N_33875);
or U35356 (N_35356,N_32572,N_34311);
or U35357 (N_35357,N_31515,N_34255);
xnor U35358 (N_35358,N_34238,N_34501);
or U35359 (N_35359,N_34621,N_32859);
and U35360 (N_35360,N_31915,N_34628);
nor U35361 (N_35361,N_30130,N_31811);
xnor U35362 (N_35362,N_31089,N_34136);
nor U35363 (N_35363,N_32673,N_32495);
nor U35364 (N_35364,N_30063,N_34674);
or U35365 (N_35365,N_34471,N_34860);
xnor U35366 (N_35366,N_32109,N_32734);
or U35367 (N_35367,N_34805,N_34697);
xnor U35368 (N_35368,N_34567,N_33206);
xor U35369 (N_35369,N_34409,N_34793);
nand U35370 (N_35370,N_33503,N_31182);
xnor U35371 (N_35371,N_33493,N_31926);
nor U35372 (N_35372,N_33279,N_32122);
or U35373 (N_35373,N_32786,N_31999);
xnor U35374 (N_35374,N_30643,N_34509);
and U35375 (N_35375,N_30694,N_30872);
xnor U35376 (N_35376,N_31001,N_31242);
nor U35377 (N_35377,N_34180,N_32180);
or U35378 (N_35378,N_33118,N_30233);
and U35379 (N_35379,N_30867,N_30251);
xnor U35380 (N_35380,N_30206,N_34395);
nor U35381 (N_35381,N_31045,N_33892);
nor U35382 (N_35382,N_30064,N_30456);
nand U35383 (N_35383,N_31500,N_30489);
nor U35384 (N_35384,N_33499,N_31902);
xor U35385 (N_35385,N_34167,N_33155);
nand U35386 (N_35386,N_31931,N_31990);
and U35387 (N_35387,N_30439,N_33652);
or U35388 (N_35388,N_30951,N_32840);
nand U35389 (N_35389,N_31878,N_32668);
nand U35390 (N_35390,N_31199,N_33978);
nor U35391 (N_35391,N_30453,N_33087);
and U35392 (N_35392,N_34110,N_30768);
or U35393 (N_35393,N_30217,N_30479);
nor U35394 (N_35394,N_34069,N_32324);
or U35395 (N_35395,N_30681,N_31822);
or U35396 (N_35396,N_30019,N_32058);
xor U35397 (N_35397,N_34455,N_33722);
and U35398 (N_35398,N_31015,N_33638);
xor U35399 (N_35399,N_30219,N_30035);
and U35400 (N_35400,N_31855,N_33927);
nand U35401 (N_35401,N_31105,N_33828);
nor U35402 (N_35402,N_30228,N_32169);
nor U35403 (N_35403,N_32191,N_32235);
or U35404 (N_35404,N_34064,N_32600);
and U35405 (N_35405,N_33006,N_34338);
or U35406 (N_35406,N_31953,N_30542);
or U35407 (N_35407,N_30576,N_34143);
nor U35408 (N_35408,N_31285,N_34074);
or U35409 (N_35409,N_34439,N_31415);
or U35410 (N_35410,N_34332,N_32130);
xor U35411 (N_35411,N_33168,N_30627);
xor U35412 (N_35412,N_34974,N_32671);
or U35413 (N_35413,N_30048,N_34354);
and U35414 (N_35414,N_30579,N_30765);
or U35415 (N_35415,N_30024,N_32220);
or U35416 (N_35416,N_33302,N_34418);
or U35417 (N_35417,N_33675,N_31263);
nor U35418 (N_35418,N_30671,N_33142);
nor U35419 (N_35419,N_32326,N_31270);
xnor U35420 (N_35420,N_30330,N_31034);
and U35421 (N_35421,N_32312,N_34855);
nor U35422 (N_35422,N_30289,N_33929);
or U35423 (N_35423,N_32218,N_34607);
and U35424 (N_35424,N_30795,N_31091);
or U35425 (N_35425,N_33402,N_32527);
or U35426 (N_35426,N_34119,N_33878);
nand U35427 (N_35427,N_32793,N_32275);
nor U35428 (N_35428,N_34079,N_30841);
and U35429 (N_35429,N_34171,N_31467);
and U35430 (N_35430,N_31137,N_34891);
xor U35431 (N_35431,N_31565,N_30457);
nor U35432 (N_35432,N_30695,N_34774);
or U35433 (N_35433,N_32884,N_32562);
and U35434 (N_35434,N_30653,N_34014);
or U35435 (N_35435,N_34759,N_31273);
xor U35436 (N_35436,N_30586,N_33869);
nand U35437 (N_35437,N_34516,N_32289);
nand U35438 (N_35438,N_34139,N_33050);
nor U35439 (N_35439,N_30544,N_32349);
nor U35440 (N_35440,N_32967,N_33445);
xor U35441 (N_35441,N_30081,N_30415);
xnor U35442 (N_35442,N_31019,N_33187);
xnor U35443 (N_35443,N_30301,N_33406);
nor U35444 (N_35444,N_31132,N_30508);
xor U35445 (N_35445,N_33992,N_30610);
or U35446 (N_35446,N_33700,N_33585);
nor U35447 (N_35447,N_32182,N_32870);
nor U35448 (N_35448,N_32034,N_32579);
and U35449 (N_35449,N_34248,N_34720);
or U35450 (N_35450,N_31323,N_31664);
and U35451 (N_35451,N_32698,N_30448);
xnor U35452 (N_35452,N_34670,N_31685);
nand U35453 (N_35453,N_32395,N_30801);
and U35454 (N_35454,N_32498,N_31432);
nor U35455 (N_35455,N_33550,N_33587);
nor U35456 (N_35456,N_30183,N_31444);
xor U35457 (N_35457,N_31320,N_32295);
nor U35458 (N_35458,N_31853,N_31268);
nor U35459 (N_35459,N_32987,N_34593);
xnor U35460 (N_35460,N_32921,N_34031);
xnor U35461 (N_35461,N_33780,N_31136);
and U35462 (N_35462,N_30808,N_34569);
and U35463 (N_35463,N_30639,N_31305);
xor U35464 (N_35464,N_33516,N_33628);
nor U35465 (N_35465,N_33617,N_33166);
or U35466 (N_35466,N_31867,N_33415);
and U35467 (N_35467,N_30209,N_31176);
xnor U35468 (N_35468,N_32219,N_31197);
nand U35469 (N_35469,N_33775,N_31225);
xor U35470 (N_35470,N_33989,N_31059);
and U35471 (N_35471,N_30444,N_33243);
xor U35472 (N_35472,N_30408,N_31104);
xnor U35473 (N_35473,N_31028,N_34473);
xor U35474 (N_35474,N_31479,N_34741);
nor U35475 (N_35475,N_31684,N_32634);
nor U35476 (N_35476,N_34825,N_32607);
and U35477 (N_35477,N_34112,N_32883);
nand U35478 (N_35478,N_30136,N_34594);
and U35479 (N_35479,N_34206,N_30083);
or U35480 (N_35480,N_33123,N_32450);
nand U35481 (N_35481,N_32431,N_33072);
or U35482 (N_35482,N_32957,N_31994);
nor U35483 (N_35483,N_31964,N_30396);
nand U35484 (N_35484,N_34306,N_31534);
and U35485 (N_35485,N_30376,N_32857);
xnor U35486 (N_35486,N_30848,N_31791);
xnor U35487 (N_35487,N_34773,N_33209);
nor U35488 (N_35488,N_30838,N_32264);
nand U35489 (N_35489,N_34636,N_34241);
or U35490 (N_35490,N_33228,N_30471);
nand U35491 (N_35491,N_30909,N_34601);
nand U35492 (N_35492,N_33537,N_34689);
and U35493 (N_35493,N_30803,N_32661);
or U35494 (N_35494,N_33896,N_34443);
xor U35495 (N_35495,N_30345,N_33766);
and U35496 (N_35496,N_34230,N_31383);
nand U35497 (N_35497,N_33518,N_30414);
nor U35498 (N_35498,N_32944,N_32950);
and U35499 (N_35499,N_31049,N_33394);
nand U35500 (N_35500,N_34207,N_31437);
and U35501 (N_35501,N_31278,N_31914);
nor U35502 (N_35502,N_30266,N_33991);
or U35503 (N_35503,N_33033,N_31548);
xnor U35504 (N_35504,N_31771,N_33805);
nor U35505 (N_35505,N_30548,N_31834);
xnor U35506 (N_35506,N_32372,N_32530);
or U35507 (N_35507,N_33149,N_34400);
nor U35508 (N_35508,N_33859,N_31116);
nand U35509 (N_35509,N_34861,N_32336);
and U35510 (N_35510,N_30977,N_32282);
or U35511 (N_35511,N_32604,N_32835);
xnor U35512 (N_35512,N_33690,N_34556);
nand U35513 (N_35513,N_33641,N_32165);
and U35514 (N_35514,N_34109,N_34733);
nand U35515 (N_35515,N_34846,N_33774);
nor U35516 (N_35516,N_33430,N_31733);
or U35517 (N_35517,N_32768,N_32127);
and U35518 (N_35518,N_31038,N_30869);
nor U35519 (N_35519,N_30405,N_31951);
xnor U35520 (N_35520,N_31478,N_30562);
nor U35521 (N_35521,N_32073,N_30078);
xnor U35522 (N_35522,N_32717,N_32676);
nor U35523 (N_35523,N_34657,N_34478);
nand U35524 (N_35524,N_31152,N_34052);
nor U35525 (N_35525,N_31966,N_33404);
nor U35526 (N_35526,N_33522,N_32715);
or U35527 (N_35527,N_34267,N_30963);
nand U35528 (N_35528,N_30966,N_32653);
and U35529 (N_35529,N_33683,N_31760);
and U35530 (N_35530,N_31166,N_34877);
nor U35531 (N_35531,N_31078,N_32255);
nor U35532 (N_35532,N_30480,N_30410);
xor U35533 (N_35533,N_33855,N_31221);
nand U35534 (N_35534,N_31442,N_31399);
nand U35535 (N_35535,N_32143,N_32384);
xnor U35536 (N_35536,N_34044,N_34704);
nor U35537 (N_35537,N_30733,N_30232);
nor U35538 (N_35538,N_31777,N_32637);
nor U35539 (N_35539,N_34618,N_30886);
and U35540 (N_35540,N_32308,N_31195);
nor U35541 (N_35541,N_33605,N_31933);
or U35542 (N_35542,N_32232,N_33491);
and U35543 (N_35543,N_33207,N_30094);
xnor U35544 (N_35544,N_32093,N_32518);
nand U35545 (N_35545,N_32106,N_30441);
or U35546 (N_35546,N_34782,N_32501);
or U35547 (N_35547,N_33334,N_31021);
nor U35548 (N_35548,N_33893,N_32303);
nand U35549 (N_35549,N_34434,N_30831);
nor U35550 (N_35550,N_31901,N_32523);
nand U35551 (N_35551,N_32558,N_33203);
or U35552 (N_35552,N_34058,N_32298);
or U35553 (N_35553,N_31829,N_30651);
nand U35554 (N_35554,N_33511,N_33566);
and U35555 (N_35555,N_32214,N_34327);
nand U35556 (N_35556,N_33599,N_30455);
xnor U35557 (N_35557,N_32158,N_31508);
nand U35558 (N_35558,N_34330,N_33210);
nor U35559 (N_35559,N_34384,N_30743);
nor U35560 (N_35560,N_32054,N_30782);
or U35561 (N_35561,N_33001,N_31547);
nand U35562 (N_35562,N_31773,N_31159);
nand U35563 (N_35563,N_34917,N_34585);
nor U35564 (N_35564,N_32172,N_31716);
nand U35565 (N_35565,N_32098,N_30982);
or U35566 (N_35566,N_34224,N_31394);
and U35567 (N_35567,N_33881,N_31734);
nand U35568 (N_35568,N_32858,N_30127);
nand U35569 (N_35569,N_31541,N_30187);
xor U35570 (N_35570,N_34246,N_31671);
nand U35571 (N_35571,N_34432,N_34022);
or U35572 (N_35572,N_30667,N_32407);
or U35573 (N_35573,N_34024,N_30833);
nor U35574 (N_35574,N_30555,N_32452);
xnor U35575 (N_35575,N_31010,N_32005);
nor U35576 (N_35576,N_32595,N_33946);
and U35577 (N_35577,N_31439,N_30322);
nand U35578 (N_35578,N_34605,N_33449);
xnor U35579 (N_35579,N_30123,N_32986);
xnor U35580 (N_35580,N_31625,N_30644);
and U35581 (N_35581,N_31977,N_31276);
nand U35582 (N_35582,N_31296,N_32599);
and U35583 (N_35583,N_33140,N_32209);
nor U35584 (N_35584,N_30930,N_34300);
xnor U35585 (N_35585,N_31770,N_33384);
nor U35586 (N_35586,N_30557,N_30656);
nor U35587 (N_35587,N_30535,N_32788);
or U35588 (N_35588,N_32694,N_33372);
and U35589 (N_35589,N_30918,N_34510);
xnor U35590 (N_35590,N_33610,N_32751);
and U35591 (N_35591,N_30147,N_30997);
xor U35592 (N_35592,N_32820,N_31655);
nand U35593 (N_35593,N_32565,N_31587);
and U35594 (N_35594,N_32867,N_31865);
xor U35595 (N_35595,N_33936,N_33065);
and U35596 (N_35596,N_31647,N_34837);
or U35597 (N_35597,N_31916,N_33161);
and U35598 (N_35598,N_34213,N_34813);
nand U35599 (N_35599,N_34157,N_30584);
and U35600 (N_35600,N_30170,N_34092);
or U35601 (N_35601,N_32103,N_34904);
or U35602 (N_35602,N_34117,N_31965);
and U35603 (N_35603,N_32118,N_31509);
or U35604 (N_35604,N_31832,N_30962);
and U35605 (N_35605,N_33995,N_33422);
or U35606 (N_35606,N_32789,N_32843);
nand U35607 (N_35607,N_30277,N_31603);
and U35608 (N_35608,N_33796,N_33717);
nor U35609 (N_35609,N_34278,N_34997);
nor U35610 (N_35610,N_33658,N_33643);
nand U35611 (N_35611,N_33572,N_31065);
nor U35612 (N_35612,N_33951,N_30025);
or U35613 (N_35613,N_31788,N_33322);
and U35614 (N_35614,N_30632,N_32811);
nor U35615 (N_35615,N_34820,N_32428);
nand U35616 (N_35616,N_32545,N_31403);
and U35617 (N_35617,N_30529,N_32798);
or U35618 (N_35618,N_33114,N_32968);
or U35619 (N_35619,N_34122,N_32626);
nand U35620 (N_35620,N_31075,N_31163);
or U35621 (N_35621,N_33452,N_30932);
nor U35622 (N_35622,N_33135,N_34367);
nand U35623 (N_35623,N_30678,N_32123);
or U35624 (N_35624,N_33036,N_33470);
xor U35625 (N_35625,N_30273,N_30045);
nand U35626 (N_35626,N_30592,N_30068);
and U35627 (N_35627,N_31665,N_31843);
nor U35628 (N_35628,N_33689,N_31050);
nor U35629 (N_35629,N_31794,N_33484);
or U35630 (N_35630,N_34642,N_30032);
xor U35631 (N_35631,N_33915,N_33417);
nand U35632 (N_35632,N_34953,N_31024);
xor U35633 (N_35633,N_33188,N_31572);
nor U35634 (N_35634,N_32049,N_33464);
and U35635 (N_35635,N_34584,N_30836);
nor U35636 (N_35636,N_33538,N_31967);
and U35637 (N_35637,N_30399,N_33656);
nor U35638 (N_35638,N_34283,N_33139);
or U35639 (N_35639,N_34090,N_31525);
or U35640 (N_35640,N_31590,N_34883);
nand U35641 (N_35641,N_34508,N_32357);
xnor U35642 (N_35642,N_33331,N_33549);
xor U35643 (N_35643,N_33787,N_33163);
nand U35644 (N_35644,N_33781,N_33848);
or U35645 (N_35645,N_32666,N_32769);
xnor U35646 (N_35646,N_31094,N_31119);
nand U35647 (N_35647,N_33162,N_30777);
xor U35648 (N_35648,N_33038,N_32485);
nand U35649 (N_35649,N_33348,N_33853);
and U35650 (N_35650,N_34555,N_30866);
and U35651 (N_35651,N_33611,N_33091);
xnor U35652 (N_35652,N_33189,N_30919);
xor U35653 (N_35653,N_31944,N_31106);
nand U35654 (N_35654,N_32948,N_34301);
and U35655 (N_35655,N_30972,N_33614);
and U35656 (N_35656,N_30429,N_31140);
nor U35657 (N_35657,N_34777,N_32837);
or U35658 (N_35658,N_30870,N_32141);
xor U35659 (N_35659,N_32864,N_33868);
xnor U35660 (N_35660,N_31960,N_31514);
nand U35661 (N_35661,N_34059,N_32780);
nor U35662 (N_35662,N_33904,N_31768);
and U35663 (N_35663,N_34527,N_33897);
or U35664 (N_35664,N_31262,N_32335);
xnor U35665 (N_35665,N_34356,N_30120);
and U35666 (N_35666,N_33945,N_30917);
nor U35667 (N_35667,N_30900,N_30517);
nand U35668 (N_35668,N_32377,N_32842);
xnor U35669 (N_35669,N_32973,N_32474);
xnor U35670 (N_35670,N_31148,N_30506);
and U35671 (N_35671,N_32057,N_30447);
xnor U35672 (N_35672,N_34252,N_32250);
nand U35673 (N_35673,N_33964,N_33167);
or U35674 (N_35674,N_30772,N_34096);
nand U35675 (N_35675,N_34951,N_34640);
and U35676 (N_35676,N_34734,N_32805);
xor U35677 (N_35677,N_31074,N_34742);
xor U35678 (N_35678,N_30043,N_31984);
and U35679 (N_35679,N_30766,N_32969);
nor U35680 (N_35680,N_32823,N_34986);
nand U35681 (N_35681,N_31489,N_33646);
or U35682 (N_35682,N_33299,N_34517);
or U35683 (N_35683,N_34895,N_30409);
or U35684 (N_35684,N_33242,N_33661);
and U35685 (N_35685,N_31998,N_33958);
or U35686 (N_35686,N_31347,N_30961);
xnor U35687 (N_35687,N_33784,N_32989);
and U35688 (N_35688,N_33442,N_34312);
xor U35689 (N_35689,N_34416,N_31035);
xor U35690 (N_35690,N_34732,N_32667);
xor U35691 (N_35691,N_33138,N_31648);
xnor U35692 (N_35692,N_33600,N_32060);
or U35693 (N_35693,N_30942,N_31061);
xor U35694 (N_35694,N_30625,N_30899);
nand U35695 (N_35695,N_31315,N_33409);
and U35696 (N_35696,N_32744,N_34083);
or U35697 (N_35697,N_34546,N_31255);
or U35698 (N_35698,N_31127,N_34209);
nor U35699 (N_35699,N_31837,N_31438);
xnor U35700 (N_35700,N_34137,N_33625);
nand U35701 (N_35701,N_32424,N_31711);
xor U35702 (N_35702,N_30283,N_33874);
nand U35703 (N_35703,N_33124,N_32440);
xor U35704 (N_35704,N_30874,N_30503);
xnor U35705 (N_35705,N_30008,N_30980);
nand U35706 (N_35706,N_34179,N_31079);
xor U35707 (N_35707,N_33788,N_34616);
and U35708 (N_35708,N_30373,N_32484);
or U35709 (N_35709,N_31701,N_33327);
nand U35710 (N_35710,N_32892,N_30347);
or U35711 (N_35711,N_32194,N_33246);
xnor U35712 (N_35712,N_31576,N_32405);
and U35713 (N_35713,N_30458,N_30022);
nand U35714 (N_35714,N_31150,N_34534);
or U35715 (N_35715,N_30226,N_32617);
or U35716 (N_35716,N_34427,N_31372);
or U35717 (N_35717,N_30167,N_34919);
or U35718 (N_35718,N_33132,N_31291);
and U35719 (N_35719,N_30884,N_32087);
nand U35720 (N_35720,N_33000,N_33740);
and U35721 (N_35721,N_30182,N_30259);
and U35722 (N_35722,N_31559,N_31621);
nor U35723 (N_35723,N_32081,N_30235);
nor U35724 (N_35724,N_34968,N_31426);
nand U35725 (N_35725,N_32828,N_31669);
xor U35726 (N_35726,N_32690,N_34142);
nor U35727 (N_35727,N_32638,N_32068);
nand U35728 (N_35728,N_30968,N_31615);
xnor U35729 (N_35729,N_34245,N_31098);
and U35730 (N_35730,N_33962,N_34271);
xor U35731 (N_35731,N_30666,N_32471);
or U35732 (N_35732,N_30113,N_31180);
xnor U35733 (N_35733,N_33583,N_31398);
and U35734 (N_35734,N_30042,N_34280);
or U35735 (N_35735,N_33669,N_30454);
or U35736 (N_35736,N_32772,N_32001);
nor U35737 (N_35737,N_34655,N_34874);
nor U35738 (N_35738,N_30852,N_31897);
or U35739 (N_35739,N_32174,N_34577);
nor U35740 (N_35740,N_32996,N_31128);
or U35741 (N_35741,N_33257,N_32826);
and U35742 (N_35742,N_30263,N_30894);
nand U35743 (N_35743,N_34622,N_31212);
or U35744 (N_35744,N_33684,N_34347);
nor U35745 (N_35745,N_34626,N_33514);
or U35746 (N_35746,N_34609,N_34931);
nand U35747 (N_35747,N_31531,N_34595);
nand U35748 (N_35748,N_34991,N_33580);
nand U35749 (N_35749,N_34783,N_34790);
xor U35750 (N_35750,N_33973,N_32585);
xor U35751 (N_35751,N_32928,N_30927);
or U35752 (N_35752,N_31125,N_33688);
xor U35753 (N_35753,N_34126,N_34477);
xnor U35754 (N_35754,N_32995,N_34319);
nor U35755 (N_35755,N_31510,N_34237);
and U35756 (N_35756,N_31301,N_34032);
nand U35757 (N_35757,N_33873,N_34450);
nor U35758 (N_35758,N_32362,N_32477);
xor U35759 (N_35759,N_34937,N_32919);
nor U35760 (N_35760,N_34099,N_32674);
or U35761 (N_35761,N_31654,N_33926);
nor U35762 (N_35762,N_33862,N_34075);
xor U35763 (N_35763,N_34745,N_31780);
nor U35764 (N_35764,N_30276,N_31039);
xor U35765 (N_35765,N_30762,N_32559);
nand U35766 (N_35766,N_31851,N_33259);
xor U35767 (N_35767,N_34903,N_30813);
nand U35768 (N_35768,N_33571,N_34141);
and U35769 (N_35769,N_32069,N_33314);
and U35770 (N_35770,N_33367,N_32166);
xnor U35771 (N_35771,N_34650,N_34208);
nand U35772 (N_35772,N_33070,N_33569);
nand U35773 (N_35773,N_30440,N_34378);
xnor U35774 (N_35774,N_30799,N_30944);
and U35775 (N_35775,N_33011,N_33421);
nand U35776 (N_35776,N_31778,N_31973);
or U35777 (N_35777,N_34853,N_31205);
nor U35778 (N_35778,N_31298,N_33225);
or U35779 (N_35779,N_30125,N_34781);
and U35780 (N_35780,N_31430,N_33767);
and U35781 (N_35781,N_34987,N_34934);
and U35782 (N_35782,N_31469,N_31746);
nand U35783 (N_35783,N_31076,N_34654);
nand U35784 (N_35784,N_31067,N_34155);
nand U35785 (N_35785,N_34889,N_31849);
xor U35786 (N_35786,N_33536,N_32646);
or U35787 (N_35787,N_34552,N_31885);
and U35788 (N_35788,N_34026,N_31545);
and U35789 (N_35789,N_34183,N_31835);
or U35790 (N_35790,N_33093,N_33913);
nor U35791 (N_35791,N_33743,N_30697);
and U35792 (N_35792,N_33581,N_33654);
nor U35793 (N_35793,N_32063,N_30536);
or U35794 (N_35794,N_32460,N_33459);
nor U35795 (N_35795,N_30566,N_30820);
xnor U35796 (N_35796,N_34729,N_33190);
or U35797 (N_35797,N_30609,N_34838);
nor U35798 (N_35798,N_33558,N_34291);
nor U35799 (N_35799,N_31801,N_31154);
nor U35800 (N_35800,N_30207,N_33525);
xnor U35801 (N_35801,N_31738,N_32406);
nor U35802 (N_35802,N_30071,N_31097);
xnor U35803 (N_35803,N_33560,N_30481);
xnor U35804 (N_35804,N_30445,N_34410);
or U35805 (N_35805,N_34977,N_33453);
nor U35806 (N_35806,N_33846,N_34474);
or U35807 (N_35807,N_31676,N_33005);
nor U35808 (N_35808,N_32390,N_33551);
and U35809 (N_35809,N_33023,N_32249);
nor U35810 (N_35810,N_33342,N_30514);
xor U35811 (N_35811,N_32893,N_32687);
and U35812 (N_35812,N_32574,N_34756);
nor U35813 (N_35813,N_32044,N_30984);
xnor U35814 (N_35814,N_34468,N_34973);
and U35815 (N_35815,N_32342,N_31170);
nand U35816 (N_35816,N_34750,N_30255);
nor U35817 (N_35817,N_31260,N_34376);
xnor U35818 (N_35818,N_30789,N_33909);
nand U35819 (N_35819,N_30341,N_30138);
nand U35820 (N_35820,N_31507,N_30846);
nand U35821 (N_35821,N_30553,N_31956);
nor U35822 (N_35822,N_30431,N_31864);
and U35823 (N_35823,N_31284,N_32906);
and U35824 (N_35824,N_33618,N_34442);
nand U35825 (N_35825,N_32055,N_33251);
xor U35826 (N_35826,N_33064,N_31209);
nor U35827 (N_35827,N_30339,N_31732);
xnor U35828 (N_35828,N_34886,N_32286);
xor U35829 (N_35829,N_31484,N_33673);
nor U35830 (N_35830,N_34368,N_33648);
and U35831 (N_35831,N_32914,N_33793);
nand U35832 (N_35832,N_33679,N_30477);
nor U35833 (N_35833,N_31012,N_34030);
nand U35834 (N_35834,N_34412,N_31412);
or U35835 (N_35835,N_32749,N_32560);
nand U35836 (N_35836,N_31606,N_33263);
or U35837 (N_35837,N_30282,N_33018);
nand U35838 (N_35838,N_33007,N_33009);
xnor U35839 (N_35839,N_32258,N_32366);
and U35840 (N_35840,N_34028,N_32391);
nor U35841 (N_35841,N_30406,N_32041);
nor U35842 (N_35842,N_32577,N_31431);
and U35843 (N_35843,N_32263,N_31526);
and U35844 (N_35844,N_32378,N_30629);
or U35845 (N_35845,N_30482,N_30356);
and U35846 (N_35846,N_33266,N_33121);
xnor U35847 (N_35847,N_32006,N_34749);
nor U35848 (N_35848,N_30334,N_30595);
nor U35849 (N_35849,N_34614,N_32831);
or U35850 (N_35850,N_31186,N_34668);
nor U35851 (N_35851,N_31869,N_32184);
or U35852 (N_35852,N_30647,N_32695);
or U35853 (N_35853,N_32953,N_30923);
nor U35854 (N_35854,N_31544,N_32534);
xnor U35855 (N_35855,N_33171,N_31083);
xnor U35856 (N_35856,N_33588,N_32680);
or U35857 (N_35857,N_33956,N_34707);
xor U35858 (N_35858,N_33202,N_31992);
and U35859 (N_35859,N_30975,N_31850);
or U35860 (N_35860,N_31758,N_32614);
or U35861 (N_35861,N_34538,N_33837);
nor U35862 (N_35862,N_33107,N_32999);
xor U35863 (N_35863,N_33541,N_32977);
and U35864 (N_35864,N_32454,N_30214);
or U35865 (N_35865,N_32434,N_30574);
nand U35866 (N_35866,N_30220,N_30781);
or U35867 (N_35867,N_32146,N_30096);
nand U35868 (N_35868,N_33144,N_34694);
or U35869 (N_35869,N_34664,N_34403);
nor U35870 (N_35870,N_31972,N_34195);
or U35871 (N_35871,N_33521,N_31256);
or U35872 (N_35872,N_30314,N_34936);
nand U35873 (N_35873,N_32776,N_31138);
nand U35874 (N_35874,N_33735,N_33507);
nor U35875 (N_35875,N_32433,N_32261);
xor U35876 (N_35876,N_34511,N_34431);
and U35877 (N_35877,N_33667,N_30175);
nand U35878 (N_35878,N_34242,N_33834);
nand U35879 (N_35879,N_33076,N_31637);
and U35880 (N_35880,N_32568,N_31179);
xor U35881 (N_35881,N_34495,N_31304);
and U35882 (N_35882,N_34576,N_30943);
and U35883 (N_35883,N_32065,N_31923);
nor U35884 (N_35884,N_30225,N_32139);
nand U35885 (N_35885,N_30507,N_34070);
or U35886 (N_35886,N_30131,N_30252);
nor U35887 (N_35887,N_33220,N_30497);
xor U35888 (N_35888,N_31696,N_34780);
xor U35889 (N_35889,N_32723,N_32852);
nand U35890 (N_35890,N_34809,N_30936);
xor U35891 (N_35891,N_34541,N_31954);
nand U35892 (N_35892,N_33042,N_32866);
and U35893 (N_35893,N_33758,N_34764);
or U35894 (N_35894,N_34865,N_30009);
nand U35895 (N_35895,N_33555,N_30224);
nor U35896 (N_35896,N_34163,N_30741);
xnor U35897 (N_35897,N_34498,N_34128);
or U35898 (N_35898,N_32204,N_30312);
nor U35899 (N_35899,N_33169,N_33702);
nand U35900 (N_35900,N_34718,N_32856);
nor U35901 (N_35901,N_33923,N_30145);
xor U35902 (N_35902,N_32511,N_31149);
xor U35903 (N_35903,N_32582,N_31406);
or U35904 (N_35904,N_32506,N_34019);
xor U35905 (N_35905,N_31202,N_30578);
xor U35906 (N_35906,N_31017,N_30934);
nor U35907 (N_35907,N_31360,N_32597);
and U35908 (N_35908,N_32713,N_34249);
nand U35909 (N_35909,N_32105,N_30725);
nor U35910 (N_35910,N_30950,N_33052);
xnor U35911 (N_35911,N_31496,N_33726);
xor U35912 (N_35912,N_30066,N_31555);
and U35913 (N_35913,N_32797,N_34138);
nand U35914 (N_35914,N_30683,N_30850);
or U35915 (N_35915,N_32089,N_32932);
xor U35916 (N_35916,N_33089,N_30729);
or U35917 (N_35917,N_34671,N_33508);
nand U35918 (N_35918,N_31319,N_34867);
and U35919 (N_35919,N_33836,N_34835);
or U35920 (N_35920,N_32245,N_31838);
nand U35921 (N_35921,N_32251,N_30754);
nor U35922 (N_35922,N_34573,N_31612);
and U35923 (N_35923,N_33292,N_30160);
nor U35924 (N_35924,N_30198,N_32299);
or U35925 (N_35925,N_31673,N_33990);
nand U35926 (N_35926,N_32291,N_30749);
nand U35927 (N_35927,N_34503,N_33347);
and U35928 (N_35928,N_31131,N_32760);
xnor U35929 (N_35929,N_30292,N_32669);
or U35930 (N_35930,N_33910,N_31073);
and U35931 (N_35931,N_31946,N_30518);
and U35932 (N_35932,N_34307,N_33380);
or U35933 (N_35933,N_31543,N_34274);
or U35934 (N_35934,N_34104,N_33357);
nor U35935 (N_35935,N_31451,N_30437);
xor U35936 (N_35936,N_31971,N_32625);
xor U35937 (N_35937,N_34459,N_30346);
or U35938 (N_35938,N_33456,N_33420);
nor U35939 (N_35939,N_34727,N_32019);
nand U35940 (N_35940,N_33856,N_34467);
or U35941 (N_35941,N_30858,N_30039);
or U35942 (N_35942,N_31704,N_30367);
xor U35943 (N_35943,N_30511,N_30981);
and U35944 (N_35944,N_33761,N_34197);
or U35945 (N_35945,N_31975,N_33366);
nand U35946 (N_35946,N_30432,N_32636);
nand U35947 (N_35947,N_33952,N_33752);
nor U35948 (N_35948,N_30474,N_32763);
nor U35949 (N_35949,N_33506,N_30306);
or U35950 (N_35950,N_34387,N_33003);
and U35951 (N_35951,N_32332,N_34651);
nand U35952 (N_35952,N_31830,N_30040);
xnor U35953 (N_35953,N_30546,N_34884);
nor U35954 (N_35954,N_33941,N_30607);
nor U35955 (N_35955,N_32500,N_34740);
or U35956 (N_35956,N_31101,N_30939);
and U35957 (N_35957,N_32070,N_34564);
and U35958 (N_35958,N_30759,N_32254);
nor U35959 (N_35959,N_34158,N_31058);
nor U35960 (N_35960,N_30730,N_30360);
or U35961 (N_35961,N_33573,N_30015);
or U35962 (N_35962,N_32538,N_34878);
nand U35963 (N_35963,N_34359,N_30381);
and U35964 (N_35964,N_34012,N_33085);
or U35965 (N_35965,N_34653,N_30153);
xnor U35966 (N_35966,N_34392,N_33562);
nand U35967 (N_35967,N_32469,N_32418);
nor U35968 (N_35968,N_31337,N_33333);
nor U35969 (N_35969,N_34488,N_32924);
or U35970 (N_35970,N_30088,N_30342);
xnor U35971 (N_35971,N_31561,N_34879);
or U35972 (N_35972,N_32701,N_33884);
nand U35973 (N_35973,N_32190,N_31289);
nor U35974 (N_35974,N_31783,N_31371);
nor U35975 (N_35975,N_34677,N_32681);
or U35976 (N_35976,N_32615,N_34675);
and U35977 (N_35977,N_32907,N_30427);
nand U35978 (N_35978,N_32203,N_33261);
nor U35979 (N_35979,N_31769,N_33823);
or U35980 (N_35980,N_34120,N_34219);
and U35981 (N_35981,N_32288,N_31882);
and U35982 (N_35982,N_34688,N_34251);
nand U35983 (N_35983,N_32300,N_32111);
and U35984 (N_35984,N_30673,N_30271);
and U35985 (N_35985,N_33756,N_31139);
or U35986 (N_35986,N_34118,N_33708);
xnor U35987 (N_35987,N_34565,N_31980);
nor U35988 (N_35988,N_30797,N_30422);
and U35989 (N_35989,N_30974,N_34232);
and U35990 (N_35990,N_32022,N_31044);
xor U35991 (N_35991,N_30057,N_34842);
and U35992 (N_35992,N_32561,N_32480);
nor U35993 (N_35993,N_32461,N_32972);
nand U35994 (N_35994,N_34563,N_32939);
and U35995 (N_35995,N_31351,N_31477);
nand U35996 (N_35996,N_30663,N_34559);
xnor U35997 (N_35997,N_32120,N_34182);
xor U35998 (N_35998,N_34956,N_32790);
nand U35999 (N_35999,N_31529,N_31485);
or U36000 (N_36000,N_30883,N_31947);
nand U36001 (N_36001,N_34898,N_32268);
xnor U36002 (N_36002,N_30118,N_31632);
nor U36003 (N_36003,N_33053,N_30649);
xor U36004 (N_36004,N_32117,N_34788);
xor U36005 (N_36005,N_34203,N_30122);
and U36006 (N_36006,N_31581,N_31803);
and U36007 (N_36007,N_31861,N_33463);
or U36008 (N_36008,N_33794,N_32845);
and U36009 (N_36009,N_30531,N_32624);
nor U36010 (N_36010,N_34134,N_31005);
nand U36011 (N_36011,N_30323,N_33575);
or U36012 (N_36012,N_30828,N_33350);
nand U36013 (N_36013,N_31184,N_30585);
nor U36014 (N_36014,N_30940,N_33325);
xor U36015 (N_36015,N_30567,N_32721);
xor U36016 (N_36016,N_32173,N_30161);
nand U36017 (N_36017,N_31257,N_30616);
and U36018 (N_36018,N_34706,N_30021);
nor U36019 (N_36019,N_33437,N_32635);
nor U36020 (N_36020,N_30670,N_31626);
or U36021 (N_36021,N_34604,N_33349);
and U36022 (N_36022,N_34010,N_34873);
nand U36023 (N_36023,N_33373,N_30680);
or U36024 (N_36024,N_33280,N_30420);
and U36025 (N_36025,N_30717,N_34797);
xor U36026 (N_36026,N_34419,N_30898);
nor U36027 (N_36027,N_33105,N_32544);
nor U36028 (N_36028,N_32731,N_33999);
or U36029 (N_36029,N_34928,N_32515);
and U36030 (N_36030,N_31542,N_33917);
nand U36031 (N_36031,N_33934,N_31857);
and U36032 (N_36032,N_34635,N_30029);
and U36033 (N_36033,N_31391,N_32328);
or U36034 (N_36034,N_33742,N_32783);
or U36035 (N_36035,N_32708,N_34446);
or U36036 (N_36036,N_33754,N_31636);
xnor U36037 (N_36037,N_30714,N_33117);
and U36038 (N_36038,N_32473,N_34539);
xor U36039 (N_36039,N_33376,N_33170);
and U36040 (N_36040,N_33026,N_30395);
or U36041 (N_36041,N_32175,N_34196);
and U36042 (N_36042,N_30104,N_33791);
nand U36043 (N_36043,N_31157,N_32492);
nand U36044 (N_36044,N_32703,N_30640);
nor U36045 (N_36045,N_31359,N_34428);
and U36046 (N_36046,N_34582,N_34736);
nand U36047 (N_36047,N_34843,N_30891);
or U36048 (N_36048,N_34739,N_31468);
xor U36049 (N_36049,N_34250,N_34362);
nand U36050 (N_36050,N_32092,N_30196);
nor U36051 (N_36051,N_33016,N_31246);
xor U36052 (N_36052,N_31056,N_34002);
and U36053 (N_36053,N_31227,N_33330);
nand U36054 (N_36054,N_34217,N_34366);
nand U36055 (N_36055,N_34485,N_30757);
nor U36056 (N_36056,N_34492,N_32389);
nand U36057 (N_36057,N_30727,N_32586);
and U36058 (N_36058,N_31293,N_30541);
xnor U36059 (N_36059,N_30272,N_34034);
and U36060 (N_36060,N_33998,N_31845);
xnor U36061 (N_36061,N_30261,N_34082);
nand U36062 (N_36062,N_32319,N_32621);
nand U36063 (N_36063,N_32567,N_34528);
nand U36064 (N_36064,N_31731,N_34114);
or U36065 (N_36065,N_33712,N_31682);
xor U36066 (N_36066,N_34060,N_30715);
nor U36067 (N_36067,N_31382,N_33125);
xor U36068 (N_36068,N_30829,N_32368);
and U36069 (N_36069,N_31985,N_30307);
nor U36070 (N_36070,N_32096,N_30319);
nor U36071 (N_36071,N_30732,N_34892);
nand U36072 (N_36072,N_33122,N_33577);
nand U36073 (N_36073,N_31454,N_32293);
xnor U36074 (N_36074,N_30462,N_31963);
nand U36075 (N_36075,N_32606,N_34826);
and U36076 (N_36076,N_34957,N_33890);
and U36077 (N_36077,N_32042,N_32990);
xor U36078 (N_36078,N_32154,N_32101);
or U36079 (N_36079,N_30107,N_31499);
and U36080 (N_36080,N_33887,N_30117);
nor U36081 (N_36081,N_30163,N_34284);
and U36082 (N_36082,N_30809,N_33037);
or U36083 (N_36083,N_34303,N_33391);
and U36084 (N_36084,N_31328,N_34802);
and U36085 (N_36085,N_30181,N_30533);
and U36086 (N_36086,N_30080,N_34684);
nor U36087 (N_36087,N_30965,N_33274);
and U36088 (N_36088,N_30184,N_32281);
nor U36089 (N_36089,N_30140,N_34444);
and U36090 (N_36090,N_34187,N_30704);
xor U36091 (N_36091,N_33158,N_31108);
and U36092 (N_36092,N_32974,N_30473);
or U36093 (N_36093,N_33902,N_30240);
nor U36094 (N_36094,N_33311,N_33413);
or U36095 (N_36095,N_32388,N_32157);
xnor U36096 (N_36096,N_33195,N_32021);
xor U36097 (N_36097,N_31556,N_34067);
nor U36098 (N_36098,N_31880,N_32346);
or U36099 (N_36099,N_31080,N_32453);
nor U36100 (N_36100,N_31554,N_30498);
xnor U36101 (N_36101,N_30229,N_34893);
xnor U36102 (N_36102,N_31380,N_34947);
nand U36103 (N_36103,N_34816,N_34871);
and U36104 (N_36104,N_34433,N_31103);
or U36105 (N_36105,N_32729,N_32356);
and U36106 (N_36106,N_31678,N_33800);
xor U36107 (N_36107,N_33268,N_34540);
xnor U36108 (N_36108,N_33498,N_30817);
or U36109 (N_36109,N_32631,N_33019);
and U36110 (N_36110,N_33010,N_31806);
nor U36111 (N_36111,N_34910,N_34097);
and U36112 (N_36112,N_31588,N_32265);
and U36113 (N_36113,N_30202,N_33770);
nand U36114 (N_36114,N_30738,N_32526);
and U36115 (N_36115,N_33888,N_33748);
nor U36116 (N_36116,N_31340,N_33594);
nand U36117 (N_36117,N_34920,N_31120);
nand U36118 (N_36118,N_32546,N_31717);
nand U36119 (N_36119,N_32547,N_30231);
nor U36120 (N_36120,N_33031,N_34696);
or U36121 (N_36121,N_31317,N_31691);
nor U36122 (N_36122,N_31286,N_33075);
and U36123 (N_36123,N_34547,N_31033);
xnor U36124 (N_36124,N_31793,N_33290);
xnor U36125 (N_36125,N_33948,N_30105);
or U36126 (N_36126,N_31404,N_34482);
and U36127 (N_36127,N_34775,N_31436);
or U36128 (N_36128,N_32524,N_33411);
nand U36129 (N_36129,N_31123,N_31272);
or U36130 (N_36130,N_33460,N_32410);
nor U36131 (N_36131,N_34523,N_32949);
and U36132 (N_36132,N_31658,N_32479);
nor U36133 (N_36133,N_31823,N_30459);
nor U36134 (N_36134,N_31909,N_33604);
or U36135 (N_36135,N_34132,N_30239);
xnor U36136 (N_36136,N_30352,N_32449);
nand U36137 (N_36137,N_32211,N_34906);
nand U36138 (N_36138,N_31240,N_30398);
nand U36139 (N_36139,N_30526,N_33938);
xor U36140 (N_36140,N_31306,N_32229);
xnor U36141 (N_36141,N_32520,N_31715);
xor U36142 (N_36142,N_34227,N_33068);
nand U36143 (N_36143,N_30007,N_33319);
or U36144 (N_36144,N_31330,N_30500);
xnor U36145 (N_36145,N_33301,N_32750);
xor U36146 (N_36146,N_33809,N_30745);
nand U36147 (N_36147,N_33370,N_31841);
and U36148 (N_36148,N_34375,N_31524);
xnor U36149 (N_36149,N_32131,N_34220);
nand U36150 (N_36150,N_33985,N_30173);
or U36151 (N_36151,N_30810,N_30606);
xnor U36152 (N_36152,N_32608,N_31043);
xor U36153 (N_36153,N_30839,N_32413);
nor U36154 (N_36154,N_33354,N_33883);
nor U36155 (N_36155,N_32854,N_32732);
nor U36156 (N_36156,N_33230,N_33972);
or U36157 (N_36157,N_33143,N_32705);
or U36158 (N_36158,N_32046,N_31313);
nor U36159 (N_36159,N_33412,N_31303);
or U36160 (N_36160,N_31847,N_33179);
nor U36161 (N_36161,N_30821,N_32112);
and U36162 (N_36162,N_32033,N_34798);
and U36163 (N_36163,N_34819,N_31173);
or U36164 (N_36164,N_33602,N_33526);
or U36165 (N_36165,N_33701,N_32409);
or U36166 (N_36166,N_34691,N_30877);
nor U36167 (N_36167,N_31688,N_32355);
nand U36168 (N_36168,N_32962,N_30089);
and U36169 (N_36169,N_30638,N_33159);
or U36170 (N_36170,N_32659,N_30617);
nand U36171 (N_36171,N_31595,N_31473);
and U36172 (N_36172,N_33227,N_34343);
nor U36173 (N_36173,N_31827,N_30788);
and U36174 (N_36174,N_34334,N_33197);
nand U36175 (N_36175,N_34103,N_30487);
and U36176 (N_36176,N_32829,N_33598);
nand U36177 (N_36177,N_31002,N_32080);
or U36178 (N_36178,N_31644,N_30659);
nand U36179 (N_36179,N_32662,N_30840);
nor U36180 (N_36180,N_33315,N_32719);
xor U36181 (N_36181,N_33996,N_33903);
nor U36182 (N_36182,N_34413,N_33647);
nand U36183 (N_36183,N_31344,N_34730);
and U36184 (N_36184,N_34320,N_33381);
nor U36185 (N_36185,N_34864,N_30783);
nand U36186 (N_36186,N_31023,N_32850);
and U36187 (N_36187,N_31957,N_30442);
nand U36188 (N_36188,N_32808,N_34404);
or U36189 (N_36189,N_34915,N_33734);
xor U36190 (N_36190,N_30134,N_32437);
and U36191 (N_36191,N_34606,N_33446);
or U36192 (N_36192,N_34890,N_33443);
and U36193 (N_36193,N_33472,N_33584);
nor U36194 (N_36194,N_32314,N_33200);
nor U36195 (N_36195,N_31527,N_30100);
xnor U36196 (N_36196,N_30769,N_32102);
and U36197 (N_36197,N_33677,N_34192);
or U36198 (N_36198,N_30570,N_31409);
nor U36199 (N_36199,N_30186,N_32200);
xnor U36200 (N_36200,N_31642,N_32392);
nor U36201 (N_36201,N_33918,N_34656);
or U36202 (N_36202,N_32622,N_32053);
and U36203 (N_36203,N_32317,N_34844);
nor U36204 (N_36204,N_31087,N_33687);
and U36205 (N_36205,N_31774,N_30636);
nand U36206 (N_36206,N_30028,N_30952);
nor U36207 (N_36207,N_33937,N_32752);
xor U36208 (N_36208,N_32197,N_31940);
or U36209 (N_36209,N_31121,N_32978);
nor U36210 (N_36210,N_34437,N_33432);
xor U36211 (N_36211,N_32724,N_33126);
xnor U36212 (N_36212,N_32316,N_32446);
xnor U36213 (N_36213,N_30552,N_34549);
nor U36214 (N_36214,N_34705,N_33488);
nor U36215 (N_36215,N_34228,N_32100);
xor U36216 (N_36216,N_31522,N_30520);
or U36217 (N_36217,N_34637,N_34345);
nand U36218 (N_36218,N_33497,N_34325);
and U36219 (N_36219,N_31551,N_32443);
or U36220 (N_36220,N_30599,N_34299);
nor U36221 (N_36221,N_33795,N_34009);
and U36222 (N_36222,N_33164,N_34944);
and U36223 (N_36223,N_33764,N_31574);
nor U36224 (N_36224,N_33260,N_33642);
xnor U36225 (N_36225,N_31175,N_34766);
nor U36226 (N_36226,N_34632,N_30059);
nand U36227 (N_36227,N_32216,N_30502);
and U36228 (N_36228,N_32040,N_32110);
nor U36229 (N_36229,N_32554,N_31395);
or U36230 (N_36230,N_30871,N_30868);
nor U36231 (N_36231,N_31820,N_34065);
xor U36232 (N_36232,N_34728,N_34981);
xnor U36233 (N_36233,N_32481,N_30337);
nand U36234 (N_36234,N_33328,N_34050);
xnor U36235 (N_36235,N_33867,N_33403);
nand U36236 (N_36236,N_30244,N_34630);
and U36237 (N_36237,N_30177,N_33877);
xnor U36238 (N_36238,N_32746,N_33601);
and U36239 (N_36239,N_33845,N_33691);
xor U36240 (N_36240,N_30731,N_31805);
nor U36241 (N_36241,N_33291,N_31418);
nand U36242 (N_36242,N_33627,N_30358);
nand U36243 (N_36243,N_33308,N_34162);
or U36244 (N_36244,N_34212,N_32341);
nor U36245 (N_36245,N_34868,N_32399);
xnor U36246 (N_36246,N_33490,N_32610);
nand U36247 (N_36247,N_30976,N_30124);
nand U36248 (N_36248,N_32758,N_32970);
xor U36249 (N_36249,N_33223,N_34814);
or U36250 (N_36250,N_34721,N_32311);
nand U36251 (N_36251,N_31591,N_34818);
xnor U36252 (N_36252,N_30856,N_32234);
or U36253 (N_36253,N_30815,N_30979);
nor U36254 (N_36254,N_30558,N_34507);
xor U36255 (N_36255,N_31905,N_30949);
nor U36256 (N_36256,N_30403,N_33059);
nand U36257 (N_36257,N_32874,N_30655);
xor U36258 (N_36258,N_34166,N_34662);
nand U36259 (N_36259,N_31281,N_31384);
nand U36260 (N_36260,N_33634,N_34669);
nor U36261 (N_36261,N_30600,N_32163);
nand U36262 (N_36262,N_30904,N_33870);
nand U36263 (N_36263,N_31222,N_33802);
nor U36264 (N_36264,N_30746,N_32900);
and U36265 (N_36265,N_31211,N_30387);
or U36266 (N_36266,N_32891,N_30534);
nand U36267 (N_36267,N_33323,N_33418);
xnor U36268 (N_36268,N_33811,N_31705);
and U36269 (N_36269,N_31025,N_32097);
or U36270 (N_36270,N_34678,N_30532);
xnor U36271 (N_36271,N_33256,N_30310);
nor U36272 (N_36272,N_33826,N_32306);
or U36273 (N_36273,N_31610,N_31349);
and U36274 (N_36274,N_34056,N_32066);
or U36275 (N_36275,N_32802,N_33184);
nand U36276 (N_36276,N_34543,N_30328);
nand U36277 (N_36277,N_30210,N_32382);
nand U36278 (N_36278,N_31772,N_33613);
or U36279 (N_36279,N_31594,N_33265);
nor U36280 (N_36280,N_30467,N_32923);
or U36281 (N_36281,N_34023,N_30859);
and U36282 (N_36282,N_30547,N_33177);
or U36283 (N_36283,N_33609,N_31487);
xnor U36284 (N_36284,N_32736,N_30412);
xor U36285 (N_36285,N_33198,N_32095);
and U36286 (N_36286,N_34875,N_32039);
nor U36287 (N_36287,N_33949,N_34186);
and U36288 (N_36288,N_32493,N_34685);
and U36289 (N_36289,N_33540,N_34315);
nand U36290 (N_36290,N_32313,N_31725);
nor U36291 (N_36291,N_31192,N_31709);
nand U36292 (N_36292,N_31297,N_32930);
xor U36293 (N_36293,N_32014,N_32457);
nand U36294 (N_36294,N_32371,N_32904);
nor U36295 (N_36295,N_31752,N_30097);
and U36296 (N_36296,N_31719,N_32702);
nand U36297 (N_36297,N_32358,N_32830);
nor U36298 (N_36298,N_33841,N_34612);
xor U36299 (N_36299,N_32880,N_34193);
xor U36300 (N_36300,N_30075,N_33426);
or U36301 (N_36301,N_31265,N_31722);
and U36302 (N_36302,N_32327,N_32872);
nor U36303 (N_36303,N_33015,N_31981);
xor U36304 (N_36304,N_31571,N_31269);
nor U36305 (N_36305,N_31870,N_32026);
xor U36306 (N_36306,N_30956,N_34978);
nand U36307 (N_36307,N_30996,N_30713);
nand U36308 (N_36308,N_33487,N_33718);
nand U36309 (N_36309,N_34236,N_34305);
and U36310 (N_36310,N_34580,N_33544);
xor U36311 (N_36311,N_34216,N_32050);
or U36312 (N_36312,N_33739,N_31638);
nand U36313 (N_36313,N_31877,N_30494);
and U36314 (N_36314,N_33919,N_33907);
xnor U36315 (N_36315,N_32077,N_32451);
nand U36316 (N_36316,N_30286,N_31617);
nand U36317 (N_36317,N_32640,N_31779);
and U36318 (N_36318,N_33699,N_33034);
or U36319 (N_36319,N_30556,N_34761);
xor U36320 (N_36320,N_33709,N_30264);
nand U36321 (N_36321,N_34261,N_32849);
and U36322 (N_36322,N_30705,N_31447);
xnor U36323 (N_36323,N_32483,N_33481);
nand U36324 (N_36324,N_31031,N_33790);
nand U36325 (N_36325,N_31077,N_32107);
nand U36326 (N_36326,N_33768,N_33082);
or U36327 (N_36327,N_31627,N_34200);
nand U36328 (N_36328,N_31086,N_31634);
xnor U36329 (N_36329,N_30238,N_34205);
xor U36330 (N_36330,N_32777,N_32882);
nand U36331 (N_36331,N_30926,N_34716);
and U36332 (N_36332,N_30044,N_33399);
nand U36333 (N_36333,N_31987,N_34673);
xor U36334 (N_36334,N_33778,N_33905);
or U36335 (N_36335,N_33310,N_34939);
nand U36336 (N_36336,N_33275,N_30661);
or U36337 (N_36337,N_34566,N_30397);
and U36338 (N_36338,N_32773,N_33760);
xnor U36339 (N_36339,N_30132,N_33080);
and U36340 (N_36340,N_34339,N_34792);
nand U36341 (N_36341,N_32573,N_34151);
nand U36342 (N_36342,N_34000,N_33205);
and U36343 (N_36343,N_32224,N_30760);
xor U36344 (N_36344,N_33547,N_30305);
nor U36345 (N_36345,N_32510,N_33344);
nor U36346 (N_36346,N_32135,N_30662);
or U36347 (N_36347,N_31706,N_33137);
or U36348 (N_36348,N_33645,N_30284);
nand U36349 (N_36349,N_30216,N_34859);
and U36350 (N_36350,N_30451,N_31641);
and U36351 (N_36351,N_30710,N_34222);
or U36352 (N_36352,N_32836,N_32832);
nor U36353 (N_36353,N_32156,N_31693);
or U36354 (N_36354,N_33217,N_31932);
and U36355 (N_36355,N_32159,N_31193);
nor U36356 (N_36356,N_31069,N_34053);
and U36357 (N_36357,N_34620,N_30230);
and U36358 (N_36358,N_34276,N_30847);
nor U36359 (N_36359,N_30637,N_32416);
or U36360 (N_36360,N_34093,N_32387);
nand U36361 (N_36361,N_34578,N_32553);
and U36362 (N_36362,N_33970,N_33473);
nor U36363 (N_36363,N_33382,N_33102);
xnor U36364 (N_36364,N_30748,N_32149);
nor U36365 (N_36365,N_34496,N_34703);
and U36366 (N_36366,N_33231,N_31251);
or U36367 (N_36367,N_30098,N_32037);
nand U36368 (N_36368,N_34399,N_33480);
xnor U36369 (N_36369,N_33273,N_33725);
xnor U36370 (N_36370,N_34817,N_33084);
xnor U36371 (N_36371,N_30472,N_34257);
or U36372 (N_36372,N_34735,N_31311);
xor U36373 (N_36373,N_30291,N_32253);
xnor U36374 (N_36374,N_31608,N_30527);
nor U36375 (N_36375,N_30992,N_34057);
nand U36376 (N_36376,N_31666,N_34281);
or U36377 (N_36377,N_33711,N_31645);
nand U36378 (N_36378,N_31381,N_30826);
xor U36379 (N_36379,N_30372,N_31821);
nand U36380 (N_36380,N_32810,N_32709);
or U36381 (N_36381,N_30164,N_33116);
xnor U36382 (N_36382,N_33419,N_30237);
nor U36383 (N_36383,N_33204,N_32541);
and U36384 (N_36384,N_31046,N_33825);
and U36385 (N_36385,N_33326,N_33636);
or U36386 (N_36386,N_32508,N_32183);
nor U36387 (N_36387,N_31969,N_34869);
nand U36388 (N_36388,N_33505,N_31776);
and U36389 (N_36389,N_31016,N_34435);
or U36390 (N_36390,N_33469,N_31407);
xnor U36391 (N_36391,N_34199,N_32816);
xor U36392 (N_36392,N_32010,N_31790);
nor U36393 (N_36393,N_32593,N_34040);
xnor U36394 (N_36394,N_30072,N_33621);
or U36395 (N_36395,N_34184,N_31164);
xnor U36396 (N_36396,N_30758,N_33844);
nor U36397 (N_36397,N_30280,N_30249);
nor U36398 (N_36398,N_32770,N_32244);
nand U36399 (N_36399,N_32943,N_33289);
nand U36400 (N_36400,N_33629,N_34445);
or U36401 (N_36401,N_32207,N_31537);
nand U36402 (N_36402,N_31893,N_31388);
nor U36403 (N_36403,N_33839,N_31493);
xor U36404 (N_36404,N_30099,N_32241);
or U36405 (N_36405,N_31792,N_34845);
or U36406 (N_36406,N_33961,N_30645);
nand U36407 (N_36407,N_31239,N_31670);
nand U36408 (N_36408,N_32320,N_31208);
or U36409 (N_36409,N_33513,N_33448);
and U36410 (N_36410,N_33115,N_33245);
nand U36411 (N_36411,N_31234,N_32321);
nor U36412 (N_36412,N_31629,N_31828);
nand U36413 (N_36413,N_34415,N_33465);
xnor U36414 (N_36414,N_33002,N_32961);
and U36415 (N_36415,N_31812,N_34452);
and U36416 (N_36416,N_30834,N_30234);
xnor U36417 (N_36417,N_33953,N_31913);
or U36418 (N_36418,N_31440,N_34262);
nor U36419 (N_36419,N_30391,N_33968);
nor U36420 (N_36420,N_33715,N_31071);
xnor U36421 (N_36421,N_34302,N_32394);
or U36422 (N_36422,N_31153,N_34029);
nand U36423 (N_36423,N_30204,N_31252);
nand U36424 (N_36424,N_34692,N_31989);
nand U36425 (N_36425,N_32623,N_30669);
xor U36426 (N_36426,N_31037,N_30853);
nand U36427 (N_36427,N_31357,N_34996);
xor U36428 (N_36428,N_34194,N_30168);
and U36429 (N_36429,N_33539,N_34645);
nand U36430 (N_36430,N_31032,N_33975);
nor U36431 (N_36431,N_32448,N_34486);
nor U36432 (N_36432,N_31151,N_32897);
nor U36433 (N_36433,N_33389,N_33976);
or U36434 (N_36434,N_31389,N_30496);
or U36435 (N_36435,N_34394,N_34346);
and U36436 (N_36436,N_30349,N_32649);
nor U36437 (N_36437,N_34148,N_33281);
nor U36438 (N_36438,N_30485,N_32304);
and U36439 (N_36439,N_34078,N_30483);
or U36440 (N_36440,N_34646,N_31674);
and U36441 (N_36441,N_32706,N_30499);
nand U36442 (N_36442,N_32027,N_31007);
nand U36443 (N_36443,N_30523,N_31470);
nand U36444 (N_36444,N_32223,N_31008);
or U36445 (N_36445,N_33681,N_31280);
nor U36446 (N_36446,N_34708,N_31775);
nor U36447 (N_36447,N_31243,N_31068);
xor U36448 (N_36448,N_34020,N_32425);
or U36449 (N_36449,N_31889,N_30126);
nand U36450 (N_36450,N_34597,N_31191);
and U36451 (N_36451,N_33267,N_30199);
and U36452 (N_36452,N_34087,N_33997);
or U36453 (N_36453,N_32879,N_33462);
or U36454 (N_36454,N_30849,N_30550);
or U36455 (N_36455,N_34297,N_30790);
and U36456 (N_36456,N_30603,N_33182);
nand U36457 (N_36457,N_32230,N_32279);
or U36458 (N_36458,N_33651,N_33128);
and U36459 (N_36459,N_32509,N_33475);
or U36460 (N_36460,N_32238,N_31130);
nand U36461 (N_36461,N_33942,N_34811);
nand U36462 (N_36462,N_31539,N_31047);
nor U36463 (N_36463,N_34420,N_33297);
and U36464 (N_36464,N_33237,N_33644);
or U36465 (N_36465,N_34382,N_31464);
nand U36466 (N_36466,N_30056,N_31147);
and U36467 (N_36467,N_32947,N_31411);
and U36468 (N_36468,N_30296,N_30191);
nand U36469 (N_36469,N_30017,N_34967);
and U36470 (N_36470,N_31321,N_30726);
and U36471 (N_36471,N_30501,N_30933);
and U36472 (N_36472,N_33920,N_32834);
and U36473 (N_36473,N_31795,N_32269);
or U36474 (N_36474,N_30587,N_30784);
or U36475 (N_36475,N_30055,N_31345);
xnor U36476 (N_36476,N_32824,N_31609);
nand U36477 (N_36477,N_32813,N_32915);
nand U36478 (N_36478,N_32578,N_31271);
and U36479 (N_36479,N_31364,N_33374);
and U36480 (N_36480,N_31907,N_30953);
or U36481 (N_36481,N_33494,N_34111);
nor U36482 (N_36482,N_31813,N_34006);
or U36483 (N_36483,N_31919,N_31528);
or U36484 (N_36484,N_34698,N_31333);
or U36485 (N_36485,N_30465,N_34554);
nor U36486 (N_36486,N_33156,N_31424);
nor U36487 (N_36487,N_30313,N_33071);
nand U36488 (N_36488,N_31628,N_34839);
or U36489 (N_36489,N_30151,N_30058);
nand U36490 (N_36490,N_30464,N_32898);
xnor U36491 (N_36491,N_31040,N_34254);
and U36492 (N_36492,N_32916,N_31392);
or U36493 (N_36493,N_33512,N_33398);
and U36494 (N_36494,N_33578,N_32651);
and U36495 (N_36495,N_32278,N_32791);
nand U36496 (N_36496,N_30378,N_30691);
and U36497 (N_36497,N_31113,N_34049);
and U36498 (N_36498,N_33249,N_32419);
nor U36499 (N_36499,N_34897,N_32000);
xor U36500 (N_36500,N_34282,N_32784);
nand U36501 (N_36501,N_33304,N_32997);
xor U36502 (N_36502,N_33680,N_33534);
or U36503 (N_36503,N_31633,N_34046);
nor U36504 (N_36504,N_30614,N_31219);
or U36505 (N_36505,N_33886,N_31720);
nand U36506 (N_36506,N_32555,N_30993);
nor U36507 (N_36507,N_31566,N_30660);
or U36508 (N_36508,N_32767,N_31564);
nand U36509 (N_36509,N_34623,N_31950);
nand U36510 (N_36510,N_30888,N_31457);
xnor U36511 (N_36511,N_31201,N_31765);
nand U36512 (N_36512,N_33375,N_33944);
nor U36513 (N_36513,N_31908,N_30624);
or U36514 (N_36514,N_31220,N_33765);
and U36515 (N_36515,N_32426,N_33390);
and U36516 (N_36516,N_31244,N_33769);
or U36517 (N_36517,N_32632,N_31703);
or U36518 (N_36518,N_33548,N_32196);
or U36519 (N_36519,N_34310,N_30046);
nor U36520 (N_36520,N_33358,N_30428);
or U36521 (N_36521,N_30519,N_34500);
nor U36522 (N_36522,N_31976,N_30227);
nor U36523 (N_36523,N_34018,N_33486);
and U36524 (N_36524,N_33930,N_33630);
and U36525 (N_36525,N_30837,N_32085);
or U36526 (N_36526,N_34411,N_31979);
and U36527 (N_36527,N_34927,N_31635);
nand U36528 (N_36528,N_33816,N_32601);
nor U36529 (N_36529,N_31030,N_32658);
xor U36530 (N_36530,N_30135,N_30994);
xor U36531 (N_36531,N_32886,N_31228);
xnor U36532 (N_36532,N_31567,N_31476);
or U36533 (N_36533,N_34841,N_33515);
nor U36534 (N_36534,N_30685,N_34786);
nand U36535 (N_36535,N_32688,N_33705);
or U36536 (N_36536,N_33444,N_32167);
nor U36537 (N_36537,N_30524,N_32691);
and U36538 (N_36538,N_32908,N_34239);
xor U36539 (N_36539,N_34526,N_33914);
xnor U36540 (N_36540,N_33857,N_31759);
or U36541 (N_36541,N_31854,N_31299);
and U36542 (N_36542,N_34408,N_32270);
and U36543 (N_36543,N_31310,N_32333);
nor U36544 (N_36544,N_32612,N_31659);
or U36545 (N_36545,N_31346,N_33885);
xnor U36546 (N_36546,N_31604,N_30889);
nand U36547 (N_36547,N_34021,N_34983);
nor U36548 (N_36548,N_34922,N_33043);
or U36549 (N_36549,N_30320,N_31840);
nand U36550 (N_36550,N_31708,N_32787);
or U36551 (N_36551,N_34264,N_31552);
or U36552 (N_36552,N_30369,N_33235);
and U36553 (N_36553,N_30290,N_32225);
and U36554 (N_36554,N_34169,N_31158);
nor U36555 (N_36555,N_32468,N_31238);
nor U36556 (N_36556,N_32665,N_32296);
nor U36557 (N_36557,N_30701,N_31401);
nor U36558 (N_36558,N_32936,N_34125);
or U36559 (N_36559,N_31000,N_30365);
nand U36560 (N_36560,N_30822,N_33741);
and U36561 (N_36561,N_34880,N_30971);
and U36562 (N_36562,N_32806,N_34982);
nor U36563 (N_36563,N_33603,N_33721);
nor U36564 (N_36564,N_30604,N_34066);
xor U36565 (N_36565,N_33527,N_30419);
xor U36566 (N_36566,N_30522,N_31266);
and U36567 (N_36567,N_34440,N_33650);
nor U36568 (N_36568,N_32353,N_30630);
nor U36569 (N_36569,N_33032,N_32400);
nand U36570 (N_36570,N_32210,N_31356);
nor U36571 (N_36571,N_33530,N_34572);
xnor U36572 (N_36572,N_32134,N_34385);
or U36573 (N_36573,N_34438,N_33424);
xnor U36574 (N_36574,N_34365,N_30385);
xor U36575 (N_36575,N_33678,N_33066);
and U36576 (N_36576,N_31099,N_33695);
nor U36577 (N_36577,N_31041,N_32693);
and U36578 (N_36578,N_30737,N_32905);
nand U36579 (N_36579,N_31474,N_34100);
and U36580 (N_36580,N_31093,N_33606);
nand U36581 (N_36581,N_31141,N_34701);
and U36582 (N_36582,N_31579,N_32730);
xor U36583 (N_36583,N_34426,N_30041);
and U36584 (N_36584,N_33664,N_34202);
xnor U36585 (N_36585,N_31013,N_31160);
xnor U36586 (N_36586,N_34921,N_32177);
nor U36587 (N_36587,N_31808,N_30077);
or U36588 (N_36588,N_34611,N_31428);
nor U36589 (N_36589,N_31824,N_30922);
nand U36590 (N_36590,N_30416,N_32710);
and U36591 (N_36591,N_34489,N_30133);
and U36592 (N_36592,N_33303,N_31859);
and U36593 (N_36593,N_30495,N_30509);
or U36594 (N_36594,N_32873,N_34648);
and U36595 (N_36595,N_34381,N_32815);
xor U36596 (N_36596,N_33738,N_30895);
or U36597 (N_36597,N_30258,N_34808);
or U36598 (N_36598,N_34108,N_31557);
and U36599 (N_36599,N_32507,N_32672);
xnor U36600 (N_36600,N_32740,N_34529);
nand U36601 (N_36601,N_31235,N_31570);
or U36602 (N_36602,N_33434,N_33316);
and U36603 (N_36603,N_31064,N_30086);
nor U36604 (N_36604,N_33020,N_33095);
xnor U36605 (N_36605,N_34107,N_31996);
nand U36606 (N_36606,N_30438,N_33108);
xor U36607 (N_36607,N_34374,N_33746);
xnor U36608 (N_36608,N_31014,N_33288);
or U36609 (N_36609,N_30069,N_32064);
and U36610 (N_36610,N_34723,N_30742);
or U36611 (N_36611,N_30382,N_31167);
xnor U36612 (N_36612,N_32934,N_30361);
xnor U36613 (N_36613,N_34831,N_33379);
nor U36614 (N_36614,N_31003,N_30590);
nand U36615 (N_36615,N_30751,N_34823);
and U36616 (N_36616,N_33894,N_31504);
and U36617 (N_36617,N_33922,N_31955);
nand U36618 (N_36618,N_31254,N_30880);
nor U36619 (N_36619,N_31318,N_33427);
or U36620 (N_36620,N_31102,N_34525);
nand U36621 (N_36621,N_30357,N_34398);
or U36622 (N_36622,N_33451,N_33668);
or U36623 (N_36623,N_33813,N_34331);
nand U36624 (N_36624,N_32911,N_33474);
nor U36625 (N_36625,N_32144,N_30370);
and U36626 (N_36626,N_30379,N_30353);
or U36627 (N_36627,N_31314,N_30152);
nand U36628 (N_36628,N_31928,N_31911);
nand U36629 (N_36629,N_33755,N_32417);
xnor U36630 (N_36630,N_30049,N_32804);
and U36631 (N_36631,N_30807,N_33960);
or U36632 (N_36632,N_32861,N_34908);
nand U36633 (N_36633,N_30915,N_34344);
nor U36634 (N_36634,N_31677,N_32910);
or U36635 (N_36635,N_31207,N_34073);
nand U36636 (N_36636,N_33264,N_34627);
or U36637 (N_36637,N_30470,N_33341);
and U36638 (N_36638,N_34116,N_34229);
nand U36639 (N_36639,N_31185,N_33051);
xnor U36640 (N_36640,N_30108,N_32287);
nor U36641 (N_36641,N_31194,N_32181);
or U36642 (N_36642,N_32351,N_31585);
xor U36643 (N_36643,N_31129,N_31506);
nand U36644 (N_36644,N_34709,N_31518);
or U36645 (N_36645,N_30303,N_32592);
or U36646 (N_36646,N_31082,N_31724);
nand U36647 (N_36647,N_32305,N_31241);
nand U36648 (N_36648,N_31694,N_30668);
or U36649 (N_36649,N_31325,N_30492);
nor U36650 (N_36650,N_32735,N_34113);
xnor U36651 (N_36651,N_32113,N_31090);
or U36652 (N_36652,N_31755,N_33519);
nor U36653 (N_36653,N_30728,N_32933);
nor U36654 (N_36654,N_34711,N_30299);
and U36655 (N_36655,N_32017,N_34955);
xnor U36656 (N_36656,N_32535,N_33935);
nand U36657 (N_36657,N_32618,N_30327);
or U36658 (N_36658,N_30192,N_31643);
or U36659 (N_36659,N_32415,N_31740);
and U36660 (N_36660,N_30154,N_32682);
or U36661 (N_36661,N_33597,N_33963);
xor U36662 (N_36662,N_30476,N_30141);
or U36663 (N_36663,N_33854,N_30892);
and U36664 (N_36664,N_30180,N_34047);
nand U36665 (N_36665,N_33130,N_30027);
xor U36666 (N_36666,N_34314,N_30521);
and U36667 (N_36667,N_33181,N_33576);
and U36668 (N_36668,N_34717,N_31786);
and U36669 (N_36669,N_30166,N_31434);
and U36670 (N_36670,N_34062,N_31938);
and U36671 (N_36671,N_33241,N_34772);
xor U36672 (N_36672,N_33988,N_31283);
or U36673 (N_36673,N_33027,N_33967);
nand U36674 (N_36674,N_30602,N_33719);
nor U36675 (N_36675,N_33492,N_30628);
nor U36676 (N_36676,N_32340,N_31247);
nor U36677 (N_36677,N_30798,N_34901);
nand U36678 (N_36678,N_34476,N_31726);
nand U36679 (N_36679,N_34061,N_34102);
nand U36680 (N_36680,N_30038,N_32380);
and U36681 (N_36681,N_32951,N_31660);
nor U36682 (N_36682,N_31575,N_31253);
nor U36683 (N_36683,N_32212,N_34757);
or U36684 (N_36684,N_31892,N_31471);
xor U36685 (N_36685,N_30700,N_32796);
and U36686 (N_36686,N_32517,N_30771);
xnor U36687 (N_36687,N_30721,N_30014);
nor U36688 (N_36688,N_31560,N_30011);
xor U36689 (N_36689,N_33175,N_31807);
nor U36690 (N_36690,N_30092,N_31441);
nand U36691 (N_36691,N_34260,N_30344);
xnor U36692 (N_36692,N_31423,N_30791);
and U36693 (N_36693,N_34681,N_31408);
and U36694 (N_36694,N_32354,N_32379);
or U36695 (N_36695,N_31721,N_30594);
nand U36696 (N_36696,N_31723,N_33626);
xor U36697 (N_36697,N_33133,N_33450);
nand U36698 (N_36698,N_31497,N_32540);
nand U36699 (N_36699,N_34004,N_34436);
xor U36700 (N_36700,N_33165,N_33186);
nor U36701 (N_36701,N_33254,N_34414);
nor U36702 (N_36702,N_33410,N_30450);
or U36703 (N_36703,N_32032,N_33178);
xnor U36704 (N_36704,N_31375,N_32359);
and U36705 (N_36705,N_32397,N_34589);
and U36706 (N_36706,N_32290,N_33111);
and U36707 (N_36707,N_31600,N_30937);
or U36708 (N_36708,N_31115,N_32931);
and U36709 (N_36709,N_30260,N_31135);
nor U36710 (N_36710,N_30641,N_32981);
xnor U36711 (N_36711,N_31936,N_33056);
and U36712 (N_36712,N_34971,N_34810);
nor U36713 (N_36713,N_32352,N_34497);
and U36714 (N_36714,N_34940,N_34725);
nor U36715 (N_36715,N_30864,N_31275);
xor U36716 (N_36716,N_33891,N_30761);
and U36717 (N_36717,N_33745,N_30208);
and U36718 (N_36718,N_31762,N_30287);
nand U36719 (N_36719,N_32699,N_31872);
xnor U36720 (N_36720,N_33747,N_34834);
xor U36721 (N_36721,N_31839,N_32528);
nor U36722 (N_36722,N_32537,N_34799);
or U36723 (N_36723,N_30193,N_30114);
nand U36724 (N_36724,N_30340,N_34665);
and U36725 (N_36725,N_31532,N_31475);
xnor U36726 (N_36726,N_30368,N_32348);
or U36727 (N_36727,N_30336,N_30332);
xor U36728 (N_36728,N_34174,N_30564);
xor U36729 (N_36729,N_30551,N_33821);
xnor U36730 (N_36730,N_34900,N_30222);
and U36731 (N_36731,N_34051,N_32894);
and U36732 (N_36732,N_30990,N_30128);
nand U36733 (N_36733,N_33048,N_34017);
nor U36734 (N_36734,N_33510,N_31896);
nand U36735 (N_36735,N_34615,N_31011);
xnor U36736 (N_36736,N_30698,N_34610);
and U36737 (N_36737,N_32361,N_32960);
and U36738 (N_36738,N_34089,N_34758);
nor U36739 (N_36739,N_31753,N_33193);
nor U36740 (N_36740,N_31172,N_31096);
or U36741 (N_36741,N_32383,N_30004);
nand U36742 (N_36742,N_32639,N_34885);
nand U36743 (N_36743,N_33899,N_33355);
and U36744 (N_36744,N_33081,N_32912);
nor U36745 (N_36745,N_34042,N_31288);
nand U36746 (N_36746,N_33054,N_33830);
xor U36747 (N_36747,N_33565,N_33751);
xnor U36748 (N_36748,N_32803,N_33586);
and U36749 (N_36749,N_32002,N_30010);
nand U36750 (N_36750,N_32442,N_30304);
nor U36751 (N_36751,N_30112,N_31084);
xnor U36752 (N_36752,N_32865,N_30964);
xnor U36753 (N_36753,N_31616,N_31335);
and U36754 (N_36754,N_32536,N_33345);
or U36755 (N_36755,N_30383,N_34214);
or U36756 (N_36756,N_30257,N_34481);
nand U36757 (N_36757,N_34349,N_31417);
xor U36758 (N_36758,N_34909,N_30111);
nand U36759 (N_36759,N_30986,N_33101);
nor U36760 (N_36760,N_30218,N_32998);
xor U36761 (N_36761,N_33931,N_33858);
xnor U36762 (N_36762,N_34397,N_34358);
xnor U36763 (N_36763,N_31991,N_31419);
nand U36764 (N_36764,N_31446,N_30689);
nor U36765 (N_36765,N_30443,N_31757);
xor U36766 (N_36766,N_34457,N_30907);
nand U36767 (N_36767,N_30274,N_33639);
nand U36768 (N_36768,N_33152,N_31085);
or U36769 (N_36769,N_33820,N_33570);
and U36770 (N_36770,N_31605,N_34407);
or U36771 (N_36771,N_33104,N_34005);
or U36772 (N_36772,N_31904,N_32647);
nor U36773 (N_36773,N_32785,N_31324);
nand U36774 (N_36774,N_30830,N_31502);
xor U36775 (N_36775,N_34778,N_30824);
nor U36776 (N_36776,N_32171,N_30335);
and U36777 (N_36777,N_33368,N_30139);
nor U36778 (N_36778,N_32059,N_33286);
xnor U36779 (N_36779,N_31613,N_32941);
or U36780 (N_36780,N_31181,N_32364);
nand U36781 (N_36781,N_32334,N_33724);
and U36782 (N_36782,N_32239,N_33441);
xnor U36783 (N_36783,N_34253,N_33619);
and U36784 (N_36784,N_30747,N_33092);
or U36785 (N_36785,N_34693,N_30780);
and U36786 (N_36786,N_34941,N_32035);
nor U36787 (N_36787,N_30559,N_30109);
nor U36788 (N_36788,N_34043,N_30082);
xor U36789 (N_36789,N_34173,N_32583);
nor U36790 (N_36790,N_32937,N_34619);
xor U36791 (N_36791,N_30605,N_30776);
xor U36792 (N_36792,N_32148,N_34077);
and U36793 (N_36793,N_30144,N_34504);
nor U36794 (N_36794,N_32711,N_33849);
or U36795 (N_36795,N_32525,N_32521);
xor U36796 (N_36796,N_32226,N_34796);
and U36797 (N_36797,N_33876,N_34176);
or U36798 (N_36798,N_34098,N_32185);
nand U36799 (N_36799,N_34600,N_32028);
xor U36800 (N_36800,N_33842,N_33792);
nor U36801 (N_36801,N_32620,N_30016);
or U36802 (N_36802,N_31747,N_34719);
or U36803 (N_36803,N_34949,N_32231);
and U36804 (N_36804,N_31165,N_33706);
nand U36805 (N_36805,N_32444,N_33763);
nor U36806 (N_36806,N_31883,N_30991);
nand U36807 (N_36807,N_33479,N_31203);
and U36808 (N_36808,N_33396,N_34634);
nand U36809 (N_36809,N_30941,N_32048);
nand U36810 (N_36810,N_34448,N_33336);
nor U36811 (N_36811,N_33017,N_31327);
nor U36812 (N_36812,N_33397,N_30561);
and U36813 (N_36813,N_34575,N_30317);
nor U36814 (N_36814,N_32971,N_34048);
xnor U36815 (N_36815,N_33993,N_32741);
xor U36816 (N_36816,N_34318,N_32633);
or U36817 (N_36817,N_33192,N_30065);
xnor U36818 (N_36818,N_33364,N_32016);
nand U36819 (N_36819,N_30881,N_30195);
or U36820 (N_36820,N_34377,N_34287);
nand U36821 (N_36821,N_34929,N_31692);
nand U36822 (N_36822,N_30248,N_30293);
nand U36823 (N_36823,N_30935,N_33276);
and U36824 (N_36824,N_31649,N_31110);
nor U36825 (N_36825,N_30709,N_33435);
xnor U36826 (N_36826,N_34185,N_34386);
xor U36827 (N_36827,N_30806,N_30931);
and U36828 (N_36828,N_30571,N_34954);
nand U36829 (N_36829,N_33832,N_33332);
nor U36830 (N_36830,N_31429,N_30692);
and U36831 (N_36831,N_34713,N_30563);
nor U36832 (N_36832,N_34373,N_32432);
xor U36833 (N_36833,N_34321,N_33236);
and U36834 (N_36834,N_32940,N_32641);
nor U36835 (N_36835,N_34976,N_34084);
nand U36836 (N_36836,N_31223,N_32496);
nand U36837 (N_36837,N_30775,N_34553);
xor U36838 (N_36838,N_31453,N_31422);
nand U36839 (N_36839,N_31218,N_31455);
and U36840 (N_36840,N_32075,N_31261);
nor U36841 (N_36841,N_30865,N_34515);
nand U36842 (N_36842,N_34680,N_31114);
xnor U36843 (N_36843,N_32920,N_34086);
nand U36844 (N_36844,N_30311,N_30102);
and U36845 (N_36845,N_30101,N_31569);
nand U36846 (N_36846,N_32575,N_34933);
nand U36847 (N_36847,N_31631,N_30648);
and U36848 (N_36848,N_34211,N_34753);
and U36849 (N_36849,N_30095,N_33337);
or U36850 (N_36850,N_34309,N_31277);
or U36851 (N_36851,N_32079,N_30735);
and U36852 (N_36852,N_32992,N_33339);
nor U36853 (N_36853,N_34308,N_32227);
nand U36854 (N_36854,N_32519,N_32072);
or U36855 (N_36855,N_33671,N_34907);
or U36856 (N_36856,N_34935,N_34938);
or U36857 (N_36857,N_32679,N_34041);
nand U36858 (N_36858,N_33865,N_32807);
nor U36859 (N_36859,N_34744,N_30620);
and U36860 (N_36860,N_32447,N_32330);
xnor U36861 (N_36861,N_34535,N_32009);
nor U36862 (N_36862,N_31941,N_34763);
xor U36863 (N_36863,N_33827,N_34960);
xor U36864 (N_36864,N_34127,N_31997);
or U36865 (N_36865,N_34544,N_31060);
nor U36866 (N_36866,N_30371,N_33649);
or U36867 (N_36867,N_33244,N_31004);
nand U36868 (N_36868,N_31761,N_33777);
and U36869 (N_36869,N_30384,N_33589);
nand U36870 (N_36870,N_33633,N_33250);
or U36871 (N_36871,N_34551,N_34999);
or U36872 (N_36872,N_33710,N_30265);
and U36873 (N_36873,N_33425,N_33145);
xor U36874 (N_36874,N_30854,N_32408);
and U36875 (N_36875,N_32007,N_32809);
nor U36876 (N_36876,N_32494,N_34905);
nand U36877 (N_36877,N_31009,N_33431);
and U36878 (N_36878,N_30176,N_31505);
nor U36879 (N_36879,N_33012,N_30269);
nor U36880 (N_36880,N_32164,N_30302);
nor U36881 (N_36881,N_33436,N_34995);
nand U36882 (N_36882,N_31844,N_33229);
nand U36883 (N_36883,N_30938,N_33545);
or U36884 (N_36884,N_30446,N_34091);
xnor U36885 (N_36885,N_31133,N_32765);
and U36886 (N_36886,N_34829,N_33959);
nor U36887 (N_36887,N_30983,N_30582);
xor U36888 (N_36888,N_32024,N_34952);
and U36889 (N_36889,N_33185,N_31177);
nor U36890 (N_36890,N_31307,N_34536);
xnor U36891 (N_36891,N_33282,N_32704);
or U36892 (N_36892,N_30411,N_33131);
nand U36893 (N_36893,N_30194,N_31568);
nand U36894 (N_36894,N_31018,N_30989);
and U36895 (N_36895,N_31036,N_30723);
and U36896 (N_36896,N_32465,N_31802);
or U36897 (N_36897,N_30885,N_30722);
xnor U36898 (N_36898,N_33247,N_30236);
and U36899 (N_36899,N_31886,N_34961);
xnor U36900 (N_36900,N_31920,N_31921);
or U36901 (N_36901,N_32584,N_31842);
and U36902 (N_36902,N_34514,N_33335);
xnor U36903 (N_36903,N_31702,N_31718);
nand U36904 (N_36904,N_33433,N_34524);
or U36905 (N_36905,N_33977,N_30608);
nor U36906 (N_36906,N_32984,N_30142);
nor U36907 (N_36907,N_30873,N_30253);
and U36908 (N_36908,N_33377,N_32136);
nor U36909 (N_36909,N_32099,N_31350);
xor U36910 (N_36910,N_31355,N_33623);
nor U36911 (N_36911,N_31922,N_33454);
nor U36912 (N_36912,N_33069,N_34755);
nor U36913 (N_36913,N_30920,N_31161);
and U36914 (N_36914,N_31448,N_34461);
nor U36915 (N_36915,N_32516,N_33191);
xnor U36916 (N_36916,N_30785,N_32887);
nor U36917 (N_36917,N_31895,N_34464);
xor U36918 (N_36918,N_34153,N_30006);
or U36919 (N_36919,N_32581,N_33129);
xnor U36920 (N_36920,N_31374,N_33843);
and U36921 (N_36921,N_32206,N_31646);
nand U36922 (N_36922,N_31675,N_31995);
or U36923 (N_36923,N_34294,N_33383);
nor U36924 (N_36924,N_34743,N_32522);
and U36925 (N_36925,N_34295,N_31656);
and U36926 (N_36926,N_34599,N_31679);
xnor U36927 (N_36927,N_33707,N_33676);
nand U36928 (N_36928,N_34293,N_30268);
and U36929 (N_36929,N_32988,N_30596);
nand U36930 (N_36930,N_30338,N_33317);
xnor U36931 (N_36931,N_30851,N_33808);
nor U36932 (N_36932,N_31052,N_30794);
and U36933 (N_36933,N_31348,N_31312);
nor U36934 (N_36934,N_32652,N_31521);
nor U36935 (N_36935,N_31189,N_31249);
and U36936 (N_36936,N_34462,N_33252);
nor U36937 (N_36937,N_33172,N_34913);
or U36938 (N_36938,N_34972,N_34747);
or U36939 (N_36939,N_32664,N_31744);
nand U36940 (N_36940,N_32628,N_32248);
xor U36941 (N_36941,N_31784,N_34794);
nor U36942 (N_36942,N_30711,N_33933);
and U36943 (N_36943,N_34984,N_33079);
nor U36944 (N_36944,N_34639,N_30642);
nand U36945 (N_36945,N_32202,N_33640);
nand U36946 (N_36946,N_33692,N_30588);
and U36947 (N_36947,N_30861,N_31986);
and U36948 (N_36948,N_34370,N_34963);
or U36949 (N_36949,N_34712,N_33532);
or U36950 (N_36950,N_31589,N_34055);
and U36951 (N_36951,N_30079,N_34406);
and U36952 (N_36952,N_33546,N_33306);
xor U36953 (N_36953,N_32013,N_34513);
nor U36954 (N_36954,N_32435,N_31029);
or U36955 (N_36955,N_30375,N_30463);
nand U36956 (N_36956,N_34383,N_31196);
nor U36957 (N_36957,N_30959,N_32370);
and U36958 (N_36958,N_32543,N_33496);
xor U36959 (N_36959,N_32486,N_33004);
or U36960 (N_36960,N_34602,N_33030);
and U36961 (N_36961,N_34268,N_31924);
nor U36962 (N_36962,N_31379,N_33098);
xor U36963 (N_36963,N_33924,N_34290);
xor U36964 (N_36964,N_33386,N_34172);
and U36965 (N_36965,N_32233,N_34993);
nand U36966 (N_36966,N_34456,N_32472);
xor U36967 (N_36967,N_31224,N_32414);
xnor U36968 (N_36968,N_31026,N_33509);
nand U36969 (N_36969,N_34943,N_30051);
nand U36970 (N_36970,N_31695,N_33966);
or U36971 (N_36971,N_31390,N_32283);
xnor U36972 (N_36972,N_32256,N_32337);
and U36973 (N_36973,N_30908,N_32222);
xor U36974 (N_36974,N_32489,N_32728);
xnor U36975 (N_36975,N_31236,N_34054);
xor U36976 (N_36976,N_31657,N_32718);
and U36977 (N_36977,N_34542,N_32170);
and U36978 (N_36978,N_31961,N_30452);
xor U36979 (N_36979,N_30275,N_31683);
or U36980 (N_36980,N_30718,N_32003);
nand U36981 (N_36981,N_32588,N_34391);
nor U36982 (N_36982,N_33468,N_30658);
nor U36983 (N_36983,N_33982,N_30756);
nor U36984 (N_36984,N_34649,N_34329);
xnor U36985 (N_36985,N_33293,N_32863);
or U36986 (N_36986,N_32052,N_33014);
nand U36987 (N_36987,N_30321,N_31190);
or U36988 (N_36988,N_31250,N_31396);
or U36989 (N_36989,N_31846,N_34360);
xnor U36990 (N_36990,N_34469,N_31690);
nor U36991 (N_36991,N_32198,N_34990);
or U36992 (N_36992,N_31573,N_31584);
nor U36993 (N_36993,N_32381,N_31856);
xnor U36994 (N_36994,N_31826,N_31814);
nor U36995 (N_36995,N_32272,N_32821);
and U36996 (N_36996,N_30377,N_32963);
or U36997 (N_36997,N_31421,N_31022);
nand U36998 (N_36998,N_34256,N_34992);
nor U36999 (N_36999,N_34272,N_30466);
or U37000 (N_37000,N_31459,N_34629);
nand U37001 (N_37001,N_32818,N_32162);
xnor U37002 (N_37002,N_31898,N_33665);
xnor U37003 (N_37003,N_34449,N_31700);
xor U37004 (N_37004,N_32552,N_30033);
xnor U37005 (N_37005,N_31063,N_32228);
or U37006 (N_37006,N_34243,N_33637);
xnor U37007 (N_37007,N_32331,N_34353);
nand U37008 (N_37008,N_30860,N_34699);
nor U37009 (N_37009,N_31766,N_31072);
nor U37010 (N_37010,N_34876,N_34215);
nor U37011 (N_37011,N_34690,N_30243);
or U37012 (N_37012,N_32684,N_30957);
nand U37013 (N_37013,N_32427,N_33458);
nor U37014 (N_37014,N_34624,N_31491);
and U37015 (N_37015,N_33219,N_32018);
nand U37016 (N_37016,N_30062,N_32318);
xnor U37017 (N_37017,N_34210,N_33025);
and U37018 (N_37018,N_32061,N_31326);
xnor U37019 (N_37019,N_30348,N_30211);
or U37020 (N_37020,N_33814,N_32955);
or U37021 (N_37021,N_31274,N_34454);
or U37022 (N_37022,N_31754,N_32609);
nand U37023 (N_37023,N_32753,N_31736);
xor U37024 (N_37024,N_31582,N_33461);
xnor U37025 (N_37025,N_30436,N_33568);
nor U37026 (N_37026,N_30985,N_34760);
and U37027 (N_37027,N_31466,N_33833);
and U37028 (N_37028,N_30724,N_33103);
nor U37029 (N_37029,N_31799,N_30945);
xnor U37030 (N_37030,N_31343,N_33786);
and U37031 (N_37031,N_33971,N_33294);
xor U37032 (N_37032,N_31974,N_31764);
and U37033 (N_37033,N_34714,N_31062);
nor U37034 (N_37034,N_30750,N_33880);
xnor U37035 (N_37035,N_32153,N_32505);
nand U37036 (N_37036,N_32764,N_30719);
nand U37037 (N_37037,N_30913,N_33467);
or U37038 (N_37038,N_34288,N_33838);
nor U37039 (N_37039,N_32503,N_32090);
or U37040 (N_37040,N_34430,N_32817);
nor U37041 (N_37041,N_30426,N_33476);
nor U37042 (N_37042,N_34324,N_34072);
nand U37043 (N_37043,N_32888,N_31210);
nand U37044 (N_37044,N_30684,N_32650);
nand U37045 (N_37045,N_33127,N_31639);
or U37046 (N_37046,N_32430,N_31088);
xor U37047 (N_37047,N_31910,N_32176);
xnor U37048 (N_37048,N_33194,N_34124);
nand U37049 (N_37049,N_30676,N_30577);
and U37050 (N_37050,N_33057,N_31369);
nor U37051 (N_37051,N_33361,N_30484);
nand U37052 (N_37052,N_32712,N_34676);
nand U37053 (N_37053,N_32643,N_31100);
nor U37054 (N_37054,N_33659,N_31342);
nor U37055 (N_37055,N_31614,N_30634);
or U37056 (N_37056,N_32917,N_34533);
or U37057 (N_37057,N_33233,N_34851);
nor U37058 (N_37058,N_32329,N_33044);
and U37059 (N_37059,N_34700,N_33798);
or U37060 (N_37060,N_34322,N_30779);
nand U37061 (N_37061,N_33556,N_32047);
nor U37062 (N_37062,N_31066,N_31836);
nor U37063 (N_37063,N_34658,N_33523);
or U37064 (N_37064,N_32121,N_33407);
nand U37065 (N_37065,N_33595,N_34916);
nor U37066 (N_37066,N_33099,N_34472);
nor U37067 (N_37067,N_33815,N_30879);
or U37068 (N_37068,N_32436,N_31767);
or U37069 (N_37069,N_31536,N_30413);
nor U37070 (N_37070,N_33060,N_31818);
or U37071 (N_37071,N_32325,N_32502);
nand U37072 (N_37072,N_34361,N_31903);
nor U37073 (N_37073,N_32985,N_32369);
or U37074 (N_37074,N_32056,N_33554);
or U37075 (N_37075,N_30910,N_34003);
nor U37076 (N_37076,N_31890,N_33147);
nand U37077 (N_37077,N_32307,N_32178);
nand U37078 (N_37078,N_30000,N_30528);
nor U37079 (N_37079,N_34371,N_33086);
or U37080 (N_37080,N_32761,N_30896);
nor U37081 (N_37081,N_31988,N_33772);
or U37082 (N_37082,N_32860,N_34530);
xor U37083 (N_37083,N_30734,N_32801);
and U37084 (N_37084,N_33208,N_31662);
nand U37085 (N_37085,N_34866,N_34545);
or U37086 (N_37086,N_34789,N_32670);
and U37087 (N_37087,N_30770,N_31365);
and U37088 (N_37088,N_34568,N_33295);
nand U37089 (N_37089,N_33106,N_33408);
nand U37090 (N_37090,N_30753,N_32242);
nor U37091 (N_37091,N_32363,N_31741);
or U37092 (N_37092,N_30593,N_31168);
xor U37093 (N_37093,N_33174,N_30435);
and U37094 (N_37094,N_33912,N_33632);
nand U37095 (N_37095,N_32827,N_31294);
nand U37096 (N_37096,N_32145,N_30116);
nand U37097 (N_37097,N_32213,N_33061);
nor U37098 (N_37098,N_32375,N_32570);
or U37099 (N_37099,N_30573,N_33685);
or U37100 (N_37100,N_31816,N_30281);
and U37101 (N_37101,N_32792,N_30295);
nand U37102 (N_37102,N_33698,N_32743);
nand U37103 (N_37103,N_34025,N_31461);
nor U37104 (N_37104,N_34133,N_30169);
nand U37105 (N_37105,N_34505,N_32627);
nor U37106 (N_37106,N_30279,N_32737);
nand U37107 (N_37107,N_32429,N_34421);
nand U37108 (N_37108,N_31433,N_32890);
xnor U37109 (N_37109,N_30589,N_30707);
or U37110 (N_37110,N_34218,N_31681);
nand U37111 (N_37111,N_30424,N_34296);
or U37112 (N_37112,N_30223,N_31425);
xor U37113 (N_37113,N_32420,N_31107);
and U37114 (N_37114,N_32782,N_34150);
or U37115 (N_37115,N_31796,N_33400);
nand U37116 (N_37116,N_31993,N_33136);
nand U37117 (N_37117,N_30300,N_34702);
or U37118 (N_37118,N_34304,N_32848);
nand U37119 (N_37119,N_33351,N_32237);
xnor U37120 (N_37120,N_30073,N_34235);
or U37121 (N_37121,N_32590,N_34081);
xor U37122 (N_37122,N_32774,N_30654);
or U37123 (N_37123,N_32678,N_33180);
nor U37124 (N_37124,N_32344,N_30488);
nor U37125 (N_37125,N_34348,N_34966);
or U37126 (N_37126,N_31596,N_30921);
xnor U37127 (N_37127,N_33773,N_34586);
or U37128 (N_37128,N_31667,N_34458);
or U37129 (N_37129,N_34570,N_34487);
and U37130 (N_37130,N_32276,N_34490);
nand U37131 (N_37131,N_31729,N_33270);
nand U37132 (N_37132,N_33074,N_33405);
nand U37133 (N_37133,N_32132,N_33047);
nor U37134 (N_37134,N_34550,N_31081);
and U37135 (N_37135,N_32603,N_34519);
and U37136 (N_37136,N_34094,N_33776);
nor U37137 (N_37137,N_31686,N_31145);
and U37138 (N_37138,N_33097,N_33312);
or U37139 (N_37139,N_32869,N_32855);
nand U37140 (N_37140,N_30973,N_32812);
or U37141 (N_37141,N_34402,N_34683);
nor U37142 (N_37142,N_32655,N_30633);
nand U37143 (N_37143,N_33008,N_31248);
and U37144 (N_37144,N_31027,N_32125);
nand U37145 (N_37145,N_31513,N_31482);
and U37146 (N_37146,N_31884,N_33615);
and U37147 (N_37147,N_32841,N_31873);
xnor U37148 (N_37148,N_34666,N_30947);
nand U37149 (N_37149,N_31906,N_34068);
or U37150 (N_37150,N_34784,N_33979);
xor U37151 (N_37151,N_33024,N_33810);
xnor U37152 (N_37152,N_33457,N_31416);
or U37153 (N_37153,N_34911,N_32825);
nor U37154 (N_37154,N_33226,N_31730);
nand U37155 (N_37155,N_30575,N_30212);
xnor U37156 (N_37156,N_30755,N_34849);
nand U37157 (N_37157,N_30540,N_34484);
nand U37158 (N_37158,N_33861,N_30549);
or U37159 (N_37159,N_33218,N_33021);
or U37160 (N_37160,N_32569,N_32438);
nand U37161 (N_37161,N_34785,N_31737);
nand U37162 (N_37162,N_30421,N_33872);
nand U37163 (N_37163,N_34870,N_32071);
xnor U37164 (N_37164,N_31781,N_33318);
nand U37165 (N_37165,N_30179,N_32922);
nor U37166 (N_37166,N_33343,N_34460);
nand U37167 (N_37167,N_32459,N_31863);
and U37168 (N_37168,N_32115,N_30569);
or U37169 (N_37169,N_30053,N_33983);
or U37170 (N_37170,N_34695,N_30819);
or U37171 (N_37171,N_30988,N_32878);
and U37172 (N_37172,N_32794,N_34791);
and U37173 (N_37173,N_30505,N_30355);
xnor U37174 (N_37174,N_32991,N_31602);
nand U37175 (N_37175,N_34033,N_31620);
nor U37176 (N_37176,N_31549,N_32199);
nor U37177 (N_37177,N_30631,N_30469);
nand U37178 (N_37178,N_34357,N_31874);
and U37179 (N_37179,N_32613,N_34776);
and U37180 (N_37180,N_30178,N_30316);
nand U37181 (N_37181,N_32402,N_34899);
and U37182 (N_37182,N_31229,N_33824);
or U37183 (N_37183,N_31410,N_33864);
or U37184 (N_37184,N_31599,N_31748);
and U37185 (N_37185,N_33471,N_32594);
or U37186 (N_37186,N_31258,N_30635);
or U37187 (N_37187,N_30978,N_32302);
or U37188 (N_37188,N_33353,N_32901);
nor U37189 (N_37189,N_33672,N_33879);
xnor U37190 (N_37190,N_31939,N_30020);
nand U37191 (N_37191,N_31370,N_30318);
nor U37192 (N_37192,N_31712,N_30878);
nor U37193 (N_37193,N_34932,N_32876);
and U37194 (N_37194,N_34852,N_33271);
nor U37195 (N_37195,N_33801,N_32129);
nor U37196 (N_37196,N_33590,N_32692);
and U37197 (N_37197,N_32589,N_31978);
nor U37198 (N_37198,N_31174,N_30619);
nor U37199 (N_37199,N_30493,N_31918);
nand U37200 (N_37200,N_33925,N_32700);
or U37201 (N_37201,N_31519,N_30087);
xnor U37202 (N_37202,N_31825,N_32644);
nand U37203 (N_37203,N_32896,N_34748);
nor U37204 (N_37204,N_32532,N_33807);
xor U37205 (N_37205,N_33591,N_32310);
and U37206 (N_37206,N_31042,N_32322);
nor U37207 (N_37207,N_30468,N_31530);
and U37208 (N_37208,N_32918,N_31789);
xnor U37209 (N_37209,N_34233,N_30037);
xnor U37210 (N_37210,N_31948,N_34887);
and U37211 (N_37211,N_33955,N_30682);
or U37212 (N_37212,N_34135,N_33504);
or U37213 (N_37213,N_33239,N_34787);
and U37214 (N_37214,N_30823,N_31817);
nand U37215 (N_37215,N_34129,N_30159);
nor U37216 (N_37216,N_34363,N_34765);
nor U37217 (N_37217,N_31443,N_31362);
xnor U37218 (N_37218,N_34579,N_32747);
or U37219 (N_37219,N_31334,N_34105);
or U37220 (N_37220,N_33720,N_34316);
nor U37221 (N_37221,N_34225,N_31750);
nand U37222 (N_37222,N_31653,N_33723);
nand U37223 (N_37223,N_31462,N_33120);
and U37224 (N_37224,N_32404,N_31577);
or U37225 (N_37225,N_33284,N_34011);
and U37226 (N_37226,N_30146,N_34447);
and U37227 (N_37227,N_30882,N_33704);
or U37228 (N_37228,N_33146,N_34313);
and U37229 (N_37229,N_30543,N_34364);
or U37230 (N_37230,N_30792,N_31899);
nor U37231 (N_37231,N_30326,N_32648);
nor U37232 (N_37232,N_31804,N_31958);
xnor U37233 (N_37233,N_33713,N_33154);
and U37234 (N_37234,N_31460,N_32309);
nand U37235 (N_37235,N_32580,N_32725);
and U37236 (N_37236,N_32273,N_32689);
nand U37237 (N_37237,N_33987,N_34964);
or U37238 (N_37238,N_31797,N_34463);
and U37239 (N_37239,N_31233,N_32976);
nand U37240 (N_37240,N_30796,N_30242);
xnor U37241 (N_37241,N_32895,N_30842);
or U37242 (N_37242,N_31687,N_33528);
and U37243 (N_37243,N_33157,N_33285);
and U37244 (N_37244,N_34115,N_30679);
or U37245 (N_37245,N_30366,N_32243);
xnor U37246 (N_37246,N_30622,N_33543);
and U37247 (N_37247,N_31481,N_32083);
nand U37248 (N_37248,N_30999,N_33134);
nand U37249 (N_37249,N_31376,N_32464);
nor U37250 (N_37250,N_33670,N_30720);
xnor U37251 (N_37251,N_34149,N_31553);
nor U37252 (N_37252,N_30688,N_32401);
and U37253 (N_37253,N_31593,N_34231);
and U37254 (N_37254,N_32201,N_30530);
nand U37255 (N_37255,N_34830,N_32707);
xor U37256 (N_37256,N_34856,N_31879);
and U37257 (N_37257,N_33094,N_32903);
nor U37258 (N_37258,N_30646,N_32445);
and U37259 (N_37259,N_33502,N_32942);
nor U37260 (N_37260,N_32217,N_33416);
nand U37261 (N_37261,N_34638,N_30047);
or U37262 (N_37262,N_31279,N_32236);
nand U37263 (N_37263,N_34591,N_33655);
or U37264 (N_37264,N_31302,N_31501);
nor U37265 (N_37265,N_31143,N_32297);
and U37266 (N_37266,N_31155,N_34557);
nand U37267 (N_37267,N_32722,N_33438);
nand U37268 (N_37268,N_33624,N_32755);
xnor U37269 (N_37269,N_34660,N_30825);
nor U37270 (N_37270,N_32036,N_30189);
nor U37271 (N_37271,N_33932,N_33559);
nand U37272 (N_37272,N_34857,N_32966);
and U37273 (N_37273,N_32160,N_32925);
nand U37274 (N_37274,N_31452,N_33365);
nand U37275 (N_37275,N_30554,N_33369);
or U37276 (N_37276,N_34833,N_33829);
and U37277 (N_37277,N_33940,N_34279);
nor U37278 (N_37278,N_31361,N_34558);
nor U37279 (N_37279,N_31465,N_32301);
nand U37280 (N_37280,N_31171,N_31386);
nor U37281 (N_37281,N_32462,N_33148);
nor U37282 (N_37282,N_32423,N_31092);
xnor U37283 (N_37283,N_30148,N_32913);
or U37284 (N_37284,N_34836,N_30568);
or U37285 (N_37285,N_34175,N_30716);
and U37286 (N_37286,N_30354,N_33557);
xor U37287 (N_37287,N_31668,N_30736);
xnor U37288 (N_37288,N_33153,N_32795);
nand U37289 (N_37289,N_34147,N_32954);
nand U37290 (N_37290,N_33750,N_31483);
xor U37291 (N_37291,N_30374,N_34854);
xnor U37292 (N_37292,N_33716,N_33255);
and U37293 (N_37293,N_34881,N_32339);
xor U37294 (N_37294,N_32126,N_32343);
xnor U37295 (N_37295,N_30309,N_33240);
xor U37296 (N_37296,N_33631,N_31749);
nor U37297 (N_37297,N_32938,N_34170);
xnor U37298 (N_37298,N_31095,N_32838);
nor U37299 (N_37299,N_31214,N_32490);
xor U37300 (N_37300,N_34263,N_30190);
nor U37301 (N_37301,N_32605,N_30393);
and U37302 (N_37302,N_30793,N_32020);
nor U37303 (N_37303,N_31122,N_31048);
and U37304 (N_37304,N_34189,N_33112);
xnor U37305 (N_37305,N_31111,N_33898);
xor U37306 (N_37306,N_30767,N_30386);
or U37307 (N_37307,N_32557,N_30394);
and U37308 (N_37308,N_32542,N_34265);
nand U37309 (N_37309,N_33077,N_32766);
nand U37310 (N_37310,N_32259,N_30740);
or U37311 (N_37311,N_34389,N_31785);
xor U37312 (N_37312,N_31745,N_34144);
nor U37313 (N_37313,N_33296,N_33212);
nand U37314 (N_37314,N_34942,N_34754);
nor U37315 (N_37315,N_33248,N_30036);
or U37316 (N_37316,N_30001,N_33994);
xnor U37317 (N_37317,N_34994,N_32851);
or U37318 (N_37318,N_34140,N_30539);
xnor U37319 (N_37319,N_30787,N_30601);
nor U37320 (N_37320,N_30969,N_31538);
and U37321 (N_37321,N_34342,N_32616);
xnor U37322 (N_37322,N_32147,N_31367);
or U37323 (N_37323,N_32482,N_30215);
xor U37324 (N_37324,N_32367,N_32108);
nor U37325 (N_37325,N_32398,N_30580);
nand U37326 (N_37326,N_30333,N_30197);
nand U37327 (N_37327,N_34388,N_30200);
or U37328 (N_37328,N_31245,N_33363);
nor U37329 (N_37329,N_31232,N_33657);
nand U37330 (N_37330,N_32470,N_34372);
and U37331 (N_37331,N_31810,N_31435);
xor U37332 (N_37332,N_32374,N_32598);
nor U37333 (N_37333,N_31385,N_34518);
and U37334 (N_37334,N_32716,N_31387);
nand U37335 (N_37335,N_34161,N_33028);
and U37336 (N_37336,N_31378,N_34731);
nor U37337 (N_37337,N_33414,N_31353);
xnor U37338 (N_37338,N_34679,N_32839);
nor U37339 (N_37339,N_31540,N_34592);
nand U37340 (N_37340,N_30702,N_31070);
and U37341 (N_37341,N_31533,N_33199);
nor U37342 (N_37342,N_32004,N_34270);
nand U37343 (N_37343,N_30525,N_31927);
nand U37344 (N_37344,N_30664,N_31689);
and U37345 (N_37345,N_31456,N_30262);
nor U37346 (N_37346,N_34465,N_33150);
nand U37347 (N_37347,N_34234,N_33620);
or U37348 (N_37348,N_30245,N_32726);
nor U37349 (N_37349,N_34751,N_30241);
nor U37350 (N_37350,N_33947,N_30031);
nor U37351 (N_37351,N_30914,N_30023);
or U37352 (N_37352,N_31698,N_32982);
xnor U37353 (N_37353,N_34007,N_32739);
nor U37354 (N_37354,N_31144,N_34970);
nor U37355 (N_37355,N_33831,N_32456);
xor U37356 (N_37356,N_31815,N_30827);
nor U37357 (N_37357,N_33663,N_31624);
xnor U37358 (N_37358,N_30285,N_33783);
nand U37359 (N_37359,N_34085,N_30137);
nand U37360 (N_37360,N_30054,N_30970);
or U37361 (N_37361,N_30084,N_30712);
nand U37362 (N_37362,N_34985,N_33309);
xor U37363 (N_37363,N_32455,N_32421);
nor U37364 (N_37364,N_34168,N_32385);
xor U37365 (N_37365,N_33320,N_32151);
xor U37366 (N_37366,N_31204,N_34746);
and U37367 (N_37367,N_33779,N_30012);
nand U37368 (N_37368,N_33269,N_31400);
xor U37369 (N_37369,N_33466,N_30254);
nand U37370 (N_37370,N_34979,N_33029);
and U37371 (N_37371,N_33593,N_32114);
nor U37372 (N_37372,N_33529,N_34980);
nor U37373 (N_37373,N_32630,N_31488);
nand U37374 (N_37374,N_34016,N_30911);
xnor U37375 (N_37375,N_34240,N_34177);
and U37376 (N_37376,N_33895,N_30110);
or U37377 (N_37377,N_31363,N_31583);
or U37378 (N_37378,N_34858,N_31057);
and U37379 (N_37379,N_34946,N_30247);
xor U37380 (N_37380,N_31866,N_32294);
xnor U37381 (N_37381,N_33533,N_33298);
nand U37382 (N_37382,N_32193,N_32819);
nand U37383 (N_37383,N_34840,N_30657);
and U37384 (N_37384,N_34548,N_34425);
nor U37385 (N_37385,N_32563,N_33262);
or U37386 (N_37386,N_34828,N_31427);
nand U37387 (N_37387,N_32902,N_31216);
xnor U37388 (N_37388,N_34583,N_34532);
nand U37389 (N_37389,N_32458,N_33234);
nand U37390 (N_37390,N_32926,N_32945);
xor U37391 (N_37391,N_34164,N_30090);
nor U37392 (N_37392,N_33022,N_33840);
nand U37393 (N_37393,N_33943,N_31420);
xor U37394 (N_37394,N_33822,N_30103);
nor U37395 (N_37395,N_33307,N_33378);
nand U37396 (N_37396,N_30650,N_31943);
nor U37397 (N_37397,N_33215,N_30774);
nor U37398 (N_37398,N_33338,N_33253);
nand U37399 (N_37399,N_33703,N_34156);
nand U37400 (N_37400,N_33440,N_32868);
nor U37401 (N_37401,N_31187,N_34494);
nor U37402 (N_37402,N_33535,N_30297);
nor U37403 (N_37403,N_31735,N_33660);
xor U37404 (N_37404,N_31619,N_30744);
nor U37405 (N_37405,N_33714,N_33428);
xnor U37406 (N_37406,N_34926,N_33213);
nor U37407 (N_37407,N_34328,N_30686);
xnor U37408 (N_37408,N_33666,N_33616);
nor U37409 (N_37409,N_33078,N_31630);
or U37410 (N_37410,N_32571,N_31550);
nand U37411 (N_37411,N_30449,N_30512);
nor U37412 (N_37412,N_34894,N_30325);
nor U37413 (N_37413,N_34131,N_34080);
nor U37414 (N_37414,N_31714,N_32846);
xor U37415 (N_37415,N_33908,N_30832);
or U37416 (N_37416,N_32757,N_31756);
nor U37417 (N_37417,N_34574,N_33058);
and U37418 (N_37418,N_34204,N_31414);
xnor U37419 (N_37419,N_32983,N_33046);
nor U37420 (N_37420,N_32338,N_34417);
nand U37421 (N_37421,N_34914,N_34393);
nand U37422 (N_37422,N_32513,N_32733);
nand U37423 (N_37423,N_33574,N_31183);
nor U37424 (N_37424,N_32885,N_31888);
nor U37425 (N_37425,N_30835,N_30897);
xnor U37426 (N_37426,N_33921,N_34896);
or U37427 (N_37427,N_31358,N_34101);
or U37428 (N_37428,N_32086,N_30902);
or U37429 (N_37429,N_30843,N_33176);
nand U37430 (N_37430,N_34644,N_33693);
xnor U37431 (N_37431,N_31498,N_34191);
and U37432 (N_37432,N_34396,N_34959);
xnor U37433 (N_37433,N_30461,N_32029);
nand U37434 (N_37434,N_30392,N_33224);
or U37435 (N_37435,N_32266,N_31876);
and U37436 (N_37436,N_30764,N_32929);
nor U37437 (N_37437,N_31982,N_34989);
nand U37438 (N_37438,N_34512,N_30478);
nor U37439 (N_37439,N_32347,N_30076);
nor U37440 (N_37440,N_31523,N_34123);
nand U37441 (N_37441,N_31912,N_32422);
nand U37442 (N_37442,N_30115,N_34863);
nor U37443 (N_37443,N_34159,N_32038);
or U37444 (N_37444,N_30565,N_32952);
xor U37445 (N_37445,N_30845,N_34480);
and U37446 (N_37446,N_34643,N_32205);
or U37447 (N_37447,N_30687,N_30270);
nand U37448 (N_37448,N_34596,N_34710);
nand U37449 (N_37449,N_32411,N_32487);
nand U37450 (N_37450,N_32152,N_33392);
nand U37451 (N_37451,N_31332,N_34598);
or U37452 (N_37452,N_30106,N_33395);
or U37453 (N_37453,N_31563,N_31935);
nor U37454 (N_37454,N_33201,N_34499);
or U37455 (N_37455,N_34603,N_32350);
nand U37456 (N_37456,N_34752,N_34130);
nor U37457 (N_37457,N_32685,N_34633);
and U37458 (N_37458,N_34269,N_31126);
xor U37459 (N_37459,N_30185,N_32762);
nand U37460 (N_37460,N_31707,N_34631);
and U37461 (N_37461,N_32980,N_33789);
nand U37462 (N_37462,N_31727,N_31652);
nor U37463 (N_37463,N_31373,N_30591);
nor U37464 (N_37464,N_31213,N_32800);
or U37465 (N_37465,N_30213,N_32475);
xnor U37466 (N_37466,N_34737,N_31862);
and U37467 (N_37467,N_33731,N_32720);
nor U37468 (N_37468,N_32539,N_31449);
or U37469 (N_37469,N_34350,N_32591);
or U37470 (N_37470,N_33984,N_34335);
xnor U37471 (N_37471,N_30876,N_34181);
xor U37472 (N_37472,N_33757,N_30903);
nand U37473 (N_37473,N_32875,N_31511);
nand U37474 (N_37474,N_30504,N_33582);
nand U37475 (N_37475,N_34588,N_31800);
and U37476 (N_37476,N_31520,N_34039);
xnor U37477 (N_37477,N_30434,N_31292);
xnor U37478 (N_37478,N_32161,N_31881);
nand U37479 (N_37479,N_32116,N_31215);
and U37480 (N_37480,N_31393,N_33356);
nor U37481 (N_37481,N_30699,N_34686);
xor U37482 (N_37482,N_30256,N_34160);
xnor U37483 (N_37483,N_34804,N_31402);
and U37484 (N_37484,N_34401,N_34008);
nand U37485 (N_37485,N_34201,N_31900);
nor U37486 (N_37486,N_34001,N_33013);
and U37487 (N_37487,N_34561,N_33900);
and U37488 (N_37488,N_33852,N_33151);
nand U37489 (N_37489,N_31316,N_32078);
or U37490 (N_37490,N_34323,N_33674);
nand U37491 (N_37491,N_31640,N_31651);
and U37492 (N_37492,N_30763,N_31728);
nor U37493 (N_37493,N_34815,N_32045);
nor U37494 (N_37494,N_34652,N_30288);
or U37495 (N_37495,N_31503,N_34667);
nor U37496 (N_37496,N_30359,N_34285);
nand U37497 (N_37497,N_32119,N_31352);
nor U37498 (N_37498,N_31925,N_33744);
or U37499 (N_37499,N_34722,N_34821);
and U37500 (N_37500,N_34266,N_32903);
nand U37501 (N_37501,N_33342,N_32821);
nand U37502 (N_37502,N_30160,N_30215);
or U37503 (N_37503,N_31000,N_33270);
nor U37504 (N_37504,N_33137,N_34343);
xor U37505 (N_37505,N_33207,N_33220);
and U37506 (N_37506,N_33856,N_31526);
nand U37507 (N_37507,N_31824,N_34244);
or U37508 (N_37508,N_34419,N_31418);
nor U37509 (N_37509,N_33759,N_34166);
and U37510 (N_37510,N_32116,N_31835);
nor U37511 (N_37511,N_33673,N_31363);
xor U37512 (N_37512,N_32591,N_34528);
or U37513 (N_37513,N_34635,N_30178);
nand U37514 (N_37514,N_33632,N_30104);
and U37515 (N_37515,N_33189,N_31093);
nor U37516 (N_37516,N_34728,N_34444);
nor U37517 (N_37517,N_34164,N_30953);
xor U37518 (N_37518,N_30070,N_33671);
nor U37519 (N_37519,N_34366,N_31831);
nor U37520 (N_37520,N_32881,N_31505);
xnor U37521 (N_37521,N_30161,N_31507);
and U37522 (N_37522,N_32800,N_32428);
xor U37523 (N_37523,N_34516,N_32183);
xnor U37524 (N_37524,N_30261,N_31852);
or U37525 (N_37525,N_31449,N_33631);
and U37526 (N_37526,N_30717,N_31008);
or U37527 (N_37527,N_33030,N_31755);
and U37528 (N_37528,N_30897,N_32924);
and U37529 (N_37529,N_30777,N_31615);
xor U37530 (N_37530,N_33063,N_31131);
nand U37531 (N_37531,N_34867,N_30793);
or U37532 (N_37532,N_32656,N_30797);
xor U37533 (N_37533,N_31967,N_31379);
xor U37534 (N_37534,N_33899,N_33829);
or U37535 (N_37535,N_34218,N_31528);
xnor U37536 (N_37536,N_33796,N_31117);
or U37537 (N_37537,N_34982,N_32328);
nand U37538 (N_37538,N_33073,N_33074);
and U37539 (N_37539,N_30883,N_34812);
or U37540 (N_37540,N_32309,N_32131);
or U37541 (N_37541,N_31720,N_32827);
nor U37542 (N_37542,N_31940,N_34648);
nor U37543 (N_37543,N_33239,N_30469);
nand U37544 (N_37544,N_31026,N_33692);
or U37545 (N_37545,N_33458,N_32350);
nand U37546 (N_37546,N_33184,N_31211);
and U37547 (N_37547,N_32422,N_31039);
nand U37548 (N_37548,N_32616,N_30244);
and U37549 (N_37549,N_31364,N_30463);
nor U37550 (N_37550,N_34228,N_32248);
and U37551 (N_37551,N_32994,N_34364);
xnor U37552 (N_37552,N_32521,N_33426);
nor U37553 (N_37553,N_34346,N_30701);
xor U37554 (N_37554,N_32075,N_30729);
and U37555 (N_37555,N_30161,N_31359);
xnor U37556 (N_37556,N_32031,N_32410);
or U37557 (N_37557,N_32691,N_34475);
xor U37558 (N_37558,N_32795,N_32553);
nor U37559 (N_37559,N_30724,N_30333);
nand U37560 (N_37560,N_30921,N_30715);
and U37561 (N_37561,N_32717,N_30884);
xnor U37562 (N_37562,N_33709,N_34141);
xor U37563 (N_37563,N_31319,N_34969);
xnor U37564 (N_37564,N_34296,N_34242);
nand U37565 (N_37565,N_34007,N_33147);
nand U37566 (N_37566,N_34910,N_30045);
nor U37567 (N_37567,N_34556,N_34852);
nor U37568 (N_37568,N_32388,N_30821);
nor U37569 (N_37569,N_34199,N_30531);
or U37570 (N_37570,N_31558,N_34742);
nor U37571 (N_37571,N_34930,N_31765);
or U37572 (N_37572,N_33076,N_32442);
and U37573 (N_37573,N_30882,N_32123);
nand U37574 (N_37574,N_30509,N_34958);
nand U37575 (N_37575,N_33979,N_31399);
nor U37576 (N_37576,N_34188,N_33310);
nor U37577 (N_37577,N_31395,N_33276);
and U37578 (N_37578,N_32711,N_32219);
xor U37579 (N_37579,N_32747,N_34730);
xor U37580 (N_37580,N_30664,N_34251);
nand U37581 (N_37581,N_33462,N_34466);
nor U37582 (N_37582,N_32548,N_32582);
nor U37583 (N_37583,N_34140,N_33655);
nor U37584 (N_37584,N_32311,N_30904);
and U37585 (N_37585,N_34849,N_34188);
or U37586 (N_37586,N_33890,N_31883);
and U37587 (N_37587,N_32959,N_33752);
nor U37588 (N_37588,N_32506,N_34060);
and U37589 (N_37589,N_32149,N_30336);
xnor U37590 (N_37590,N_31016,N_31248);
nor U37591 (N_37591,N_32181,N_34817);
or U37592 (N_37592,N_30679,N_32749);
xnor U37593 (N_37593,N_31718,N_32875);
nand U37594 (N_37594,N_33711,N_30094);
nand U37595 (N_37595,N_32129,N_34608);
or U37596 (N_37596,N_30968,N_30958);
and U37597 (N_37597,N_34554,N_30212);
nand U37598 (N_37598,N_33748,N_31544);
nor U37599 (N_37599,N_31793,N_30123);
and U37600 (N_37600,N_34712,N_31257);
or U37601 (N_37601,N_32356,N_32774);
and U37602 (N_37602,N_33992,N_32218);
and U37603 (N_37603,N_31637,N_34997);
and U37604 (N_37604,N_33013,N_33379);
and U37605 (N_37605,N_30886,N_30375);
nor U37606 (N_37606,N_32772,N_30871);
xnor U37607 (N_37607,N_31854,N_32343);
xor U37608 (N_37608,N_33820,N_34227);
or U37609 (N_37609,N_34139,N_32125);
or U37610 (N_37610,N_31397,N_32683);
and U37611 (N_37611,N_30107,N_32540);
nand U37612 (N_37612,N_30187,N_30005);
or U37613 (N_37613,N_30844,N_33690);
or U37614 (N_37614,N_32306,N_30529);
or U37615 (N_37615,N_32182,N_34631);
xor U37616 (N_37616,N_30399,N_34354);
nor U37617 (N_37617,N_33152,N_33005);
nor U37618 (N_37618,N_34296,N_31520);
xor U37619 (N_37619,N_31888,N_30871);
xnor U37620 (N_37620,N_32942,N_33334);
or U37621 (N_37621,N_30677,N_30743);
nand U37622 (N_37622,N_32457,N_30972);
xnor U37623 (N_37623,N_32421,N_34927);
nand U37624 (N_37624,N_33972,N_32079);
nand U37625 (N_37625,N_33519,N_31958);
xor U37626 (N_37626,N_33776,N_32501);
xnor U37627 (N_37627,N_34052,N_33266);
nor U37628 (N_37628,N_34205,N_34640);
and U37629 (N_37629,N_30285,N_33560);
nor U37630 (N_37630,N_32230,N_34408);
xnor U37631 (N_37631,N_32496,N_31656);
nor U37632 (N_37632,N_32942,N_31790);
and U37633 (N_37633,N_31671,N_32630);
nand U37634 (N_37634,N_30204,N_30876);
or U37635 (N_37635,N_30225,N_31973);
xor U37636 (N_37636,N_30005,N_31116);
or U37637 (N_37637,N_34599,N_31760);
and U37638 (N_37638,N_30640,N_32089);
xor U37639 (N_37639,N_30865,N_30626);
nand U37640 (N_37640,N_32480,N_33318);
nor U37641 (N_37641,N_33244,N_31758);
nand U37642 (N_37642,N_32820,N_32226);
and U37643 (N_37643,N_30894,N_30847);
xor U37644 (N_37644,N_32406,N_33469);
nor U37645 (N_37645,N_32408,N_34169);
or U37646 (N_37646,N_31744,N_34390);
nor U37647 (N_37647,N_33462,N_31707);
nor U37648 (N_37648,N_32453,N_33644);
nor U37649 (N_37649,N_31039,N_32174);
and U37650 (N_37650,N_30565,N_32705);
or U37651 (N_37651,N_32972,N_34996);
nand U37652 (N_37652,N_34838,N_33505);
or U37653 (N_37653,N_30685,N_33738);
nand U37654 (N_37654,N_32822,N_32630);
and U37655 (N_37655,N_30251,N_30823);
and U37656 (N_37656,N_34966,N_30451);
and U37657 (N_37657,N_30800,N_30532);
and U37658 (N_37658,N_33363,N_32708);
and U37659 (N_37659,N_34358,N_31976);
and U37660 (N_37660,N_30279,N_33351);
or U37661 (N_37661,N_30822,N_33476);
xnor U37662 (N_37662,N_30990,N_33484);
and U37663 (N_37663,N_33110,N_32320);
xnor U37664 (N_37664,N_30299,N_33773);
nor U37665 (N_37665,N_32056,N_31797);
nor U37666 (N_37666,N_31993,N_34140);
or U37667 (N_37667,N_32266,N_31262);
or U37668 (N_37668,N_33807,N_31809);
and U37669 (N_37669,N_31202,N_34947);
or U37670 (N_37670,N_33854,N_32830);
xor U37671 (N_37671,N_30267,N_34883);
or U37672 (N_37672,N_33157,N_32538);
and U37673 (N_37673,N_32665,N_32986);
or U37674 (N_37674,N_32694,N_30223);
xnor U37675 (N_37675,N_31682,N_32596);
and U37676 (N_37676,N_32344,N_31832);
nand U37677 (N_37677,N_34781,N_33476);
nand U37678 (N_37678,N_33790,N_34474);
nor U37679 (N_37679,N_34257,N_34762);
xor U37680 (N_37680,N_31971,N_32759);
nand U37681 (N_37681,N_32236,N_31199);
xnor U37682 (N_37682,N_34987,N_34048);
and U37683 (N_37683,N_34404,N_33667);
nor U37684 (N_37684,N_32819,N_34911);
xor U37685 (N_37685,N_30914,N_33794);
nor U37686 (N_37686,N_34316,N_31529);
nand U37687 (N_37687,N_33179,N_34842);
and U37688 (N_37688,N_30046,N_30390);
or U37689 (N_37689,N_31344,N_32339);
and U37690 (N_37690,N_34707,N_33800);
nand U37691 (N_37691,N_34339,N_32814);
xnor U37692 (N_37692,N_34877,N_31923);
nand U37693 (N_37693,N_33116,N_34465);
or U37694 (N_37694,N_33843,N_30511);
nand U37695 (N_37695,N_33624,N_34995);
and U37696 (N_37696,N_30647,N_32552);
nand U37697 (N_37697,N_31647,N_32603);
nor U37698 (N_37698,N_32571,N_30451);
nor U37699 (N_37699,N_32157,N_31355);
or U37700 (N_37700,N_33830,N_34674);
and U37701 (N_37701,N_33713,N_31652);
or U37702 (N_37702,N_34235,N_30721);
xnor U37703 (N_37703,N_34957,N_34567);
xnor U37704 (N_37704,N_34668,N_33306);
xor U37705 (N_37705,N_33043,N_32734);
nand U37706 (N_37706,N_32337,N_31190);
nand U37707 (N_37707,N_30975,N_30014);
and U37708 (N_37708,N_30102,N_30462);
or U37709 (N_37709,N_30651,N_31967);
xor U37710 (N_37710,N_33816,N_31076);
and U37711 (N_37711,N_31338,N_30072);
and U37712 (N_37712,N_31239,N_31841);
nor U37713 (N_37713,N_31353,N_32830);
nor U37714 (N_37714,N_32605,N_33539);
and U37715 (N_37715,N_33053,N_33595);
xnor U37716 (N_37716,N_30675,N_30668);
xnor U37717 (N_37717,N_31378,N_34610);
nor U37718 (N_37718,N_30863,N_31521);
or U37719 (N_37719,N_32103,N_31850);
or U37720 (N_37720,N_30377,N_32534);
or U37721 (N_37721,N_32241,N_34776);
nand U37722 (N_37722,N_32136,N_34083);
nand U37723 (N_37723,N_32465,N_32085);
xor U37724 (N_37724,N_30351,N_30834);
xor U37725 (N_37725,N_31735,N_31746);
and U37726 (N_37726,N_31733,N_34021);
or U37727 (N_37727,N_33300,N_34934);
and U37728 (N_37728,N_34089,N_31125);
and U37729 (N_37729,N_34860,N_32593);
or U37730 (N_37730,N_31349,N_30790);
and U37731 (N_37731,N_30369,N_32195);
or U37732 (N_37732,N_34030,N_33566);
and U37733 (N_37733,N_33129,N_33806);
nand U37734 (N_37734,N_30103,N_30519);
and U37735 (N_37735,N_31882,N_33921);
nor U37736 (N_37736,N_30929,N_34117);
and U37737 (N_37737,N_33717,N_33325);
xor U37738 (N_37738,N_34278,N_32093);
nor U37739 (N_37739,N_34139,N_30106);
or U37740 (N_37740,N_33386,N_30440);
nor U37741 (N_37741,N_30732,N_34712);
nand U37742 (N_37742,N_30430,N_32081);
and U37743 (N_37743,N_30161,N_31058);
nor U37744 (N_37744,N_34150,N_31410);
or U37745 (N_37745,N_32238,N_34644);
xnor U37746 (N_37746,N_33917,N_34462);
nor U37747 (N_37747,N_33313,N_31994);
or U37748 (N_37748,N_33160,N_32231);
and U37749 (N_37749,N_30622,N_32712);
xnor U37750 (N_37750,N_31377,N_30063);
nand U37751 (N_37751,N_32203,N_32555);
nand U37752 (N_37752,N_33514,N_31977);
xnor U37753 (N_37753,N_33210,N_32356);
and U37754 (N_37754,N_33941,N_33241);
nor U37755 (N_37755,N_34714,N_30639);
nand U37756 (N_37756,N_34644,N_32894);
xnor U37757 (N_37757,N_31156,N_34099);
and U37758 (N_37758,N_30691,N_33138);
and U37759 (N_37759,N_32768,N_34884);
nand U37760 (N_37760,N_33627,N_32408);
and U37761 (N_37761,N_30292,N_34361);
or U37762 (N_37762,N_30508,N_32259);
nand U37763 (N_37763,N_33029,N_30398);
xnor U37764 (N_37764,N_31719,N_30402);
xor U37765 (N_37765,N_31248,N_34347);
nor U37766 (N_37766,N_30401,N_34447);
or U37767 (N_37767,N_30684,N_32500);
xnor U37768 (N_37768,N_33289,N_33639);
nor U37769 (N_37769,N_32551,N_30763);
or U37770 (N_37770,N_30149,N_33247);
or U37771 (N_37771,N_31573,N_30147);
and U37772 (N_37772,N_32245,N_32967);
nand U37773 (N_37773,N_31965,N_30585);
nor U37774 (N_37774,N_32513,N_33835);
nor U37775 (N_37775,N_30726,N_34090);
or U37776 (N_37776,N_31293,N_32102);
nand U37777 (N_37777,N_32299,N_30738);
nand U37778 (N_37778,N_32899,N_34151);
and U37779 (N_37779,N_30077,N_33194);
xnor U37780 (N_37780,N_33808,N_33823);
nand U37781 (N_37781,N_31377,N_33398);
xnor U37782 (N_37782,N_31008,N_32295);
nor U37783 (N_37783,N_34166,N_31783);
or U37784 (N_37784,N_30649,N_31249);
or U37785 (N_37785,N_33931,N_34844);
nor U37786 (N_37786,N_30362,N_31780);
or U37787 (N_37787,N_30111,N_32430);
nor U37788 (N_37788,N_31277,N_31805);
nand U37789 (N_37789,N_34482,N_30545);
or U37790 (N_37790,N_30680,N_32452);
or U37791 (N_37791,N_31841,N_34056);
or U37792 (N_37792,N_30663,N_33885);
or U37793 (N_37793,N_31943,N_31469);
nor U37794 (N_37794,N_34583,N_32710);
or U37795 (N_37795,N_30979,N_32451);
nand U37796 (N_37796,N_33708,N_32149);
or U37797 (N_37797,N_33007,N_31497);
or U37798 (N_37798,N_31583,N_31956);
nor U37799 (N_37799,N_32882,N_30498);
and U37800 (N_37800,N_34831,N_33857);
nand U37801 (N_37801,N_33483,N_31687);
nand U37802 (N_37802,N_31957,N_33838);
or U37803 (N_37803,N_34069,N_30454);
xor U37804 (N_37804,N_32229,N_32033);
and U37805 (N_37805,N_30592,N_31092);
or U37806 (N_37806,N_34568,N_32474);
nand U37807 (N_37807,N_31669,N_30453);
nor U37808 (N_37808,N_32197,N_33002);
or U37809 (N_37809,N_33814,N_34004);
nand U37810 (N_37810,N_31605,N_34838);
and U37811 (N_37811,N_31345,N_30967);
nor U37812 (N_37812,N_34394,N_30611);
or U37813 (N_37813,N_30960,N_31094);
nand U37814 (N_37814,N_30442,N_34523);
and U37815 (N_37815,N_30489,N_30921);
and U37816 (N_37816,N_31778,N_30509);
xnor U37817 (N_37817,N_30460,N_30406);
or U37818 (N_37818,N_33926,N_34436);
or U37819 (N_37819,N_32121,N_30143);
nor U37820 (N_37820,N_34652,N_34056);
nor U37821 (N_37821,N_32274,N_33050);
nor U37822 (N_37822,N_34500,N_32581);
or U37823 (N_37823,N_32596,N_30676);
nor U37824 (N_37824,N_31695,N_32696);
xnor U37825 (N_37825,N_34213,N_31484);
and U37826 (N_37826,N_30170,N_33549);
nand U37827 (N_37827,N_31324,N_33752);
nor U37828 (N_37828,N_34419,N_31156);
nor U37829 (N_37829,N_30038,N_32624);
nor U37830 (N_37830,N_30059,N_30234);
nand U37831 (N_37831,N_33775,N_34072);
xnor U37832 (N_37832,N_33642,N_31471);
nand U37833 (N_37833,N_32204,N_31930);
nand U37834 (N_37834,N_30408,N_32144);
nand U37835 (N_37835,N_32464,N_30765);
nor U37836 (N_37836,N_34473,N_31835);
xor U37837 (N_37837,N_33555,N_32849);
xnor U37838 (N_37838,N_34781,N_34207);
and U37839 (N_37839,N_31365,N_32240);
nor U37840 (N_37840,N_33881,N_34338);
nor U37841 (N_37841,N_31674,N_30605);
xnor U37842 (N_37842,N_31561,N_31709);
and U37843 (N_37843,N_33160,N_32425);
nand U37844 (N_37844,N_34610,N_33086);
and U37845 (N_37845,N_33644,N_32561);
nand U37846 (N_37846,N_30382,N_30808);
and U37847 (N_37847,N_33695,N_30692);
and U37848 (N_37848,N_32419,N_34649);
and U37849 (N_37849,N_31699,N_33009);
nand U37850 (N_37850,N_33516,N_33842);
xor U37851 (N_37851,N_31579,N_34371);
and U37852 (N_37852,N_30014,N_32958);
nand U37853 (N_37853,N_31928,N_30785);
nor U37854 (N_37854,N_31286,N_30226);
nor U37855 (N_37855,N_32559,N_34727);
and U37856 (N_37856,N_32133,N_33315);
nor U37857 (N_37857,N_30018,N_30973);
or U37858 (N_37858,N_32671,N_30834);
or U37859 (N_37859,N_30120,N_31522);
nor U37860 (N_37860,N_33389,N_31881);
and U37861 (N_37861,N_30303,N_33207);
nor U37862 (N_37862,N_31970,N_32198);
or U37863 (N_37863,N_34856,N_30602);
nor U37864 (N_37864,N_32774,N_33235);
and U37865 (N_37865,N_32603,N_32984);
and U37866 (N_37866,N_32505,N_33658);
or U37867 (N_37867,N_33706,N_33926);
or U37868 (N_37868,N_34291,N_30872);
and U37869 (N_37869,N_34866,N_34096);
or U37870 (N_37870,N_34791,N_33667);
nand U37871 (N_37871,N_32377,N_34673);
or U37872 (N_37872,N_33969,N_31597);
xnor U37873 (N_37873,N_31073,N_34093);
or U37874 (N_37874,N_30189,N_33727);
or U37875 (N_37875,N_31439,N_30482);
xor U37876 (N_37876,N_33603,N_34872);
xor U37877 (N_37877,N_31240,N_31462);
and U37878 (N_37878,N_32476,N_31010);
nand U37879 (N_37879,N_32117,N_31774);
and U37880 (N_37880,N_32617,N_32339);
xor U37881 (N_37881,N_33649,N_33478);
and U37882 (N_37882,N_30784,N_33214);
and U37883 (N_37883,N_34464,N_34977);
xor U37884 (N_37884,N_34270,N_33959);
nand U37885 (N_37885,N_33852,N_32446);
nand U37886 (N_37886,N_33635,N_30827);
nor U37887 (N_37887,N_31401,N_33131);
xnor U37888 (N_37888,N_31557,N_31051);
and U37889 (N_37889,N_31498,N_33914);
or U37890 (N_37890,N_33555,N_30921);
xnor U37891 (N_37891,N_33230,N_30266);
xnor U37892 (N_37892,N_30555,N_34679);
xor U37893 (N_37893,N_32151,N_33940);
and U37894 (N_37894,N_30679,N_30770);
xor U37895 (N_37895,N_33023,N_32031);
xor U37896 (N_37896,N_30392,N_32928);
xnor U37897 (N_37897,N_30504,N_30253);
nor U37898 (N_37898,N_34069,N_34881);
nor U37899 (N_37899,N_32439,N_30237);
nand U37900 (N_37900,N_31103,N_32428);
xnor U37901 (N_37901,N_31165,N_34617);
and U37902 (N_37902,N_30695,N_31721);
nor U37903 (N_37903,N_30102,N_32660);
and U37904 (N_37904,N_33713,N_34198);
nand U37905 (N_37905,N_31885,N_34087);
and U37906 (N_37906,N_33439,N_32464);
nor U37907 (N_37907,N_30046,N_31463);
or U37908 (N_37908,N_32266,N_33911);
nand U37909 (N_37909,N_30033,N_31683);
or U37910 (N_37910,N_30120,N_33981);
or U37911 (N_37911,N_30627,N_30425);
nor U37912 (N_37912,N_34719,N_33364);
nor U37913 (N_37913,N_34816,N_32344);
xnor U37914 (N_37914,N_31592,N_34319);
or U37915 (N_37915,N_34900,N_30511);
and U37916 (N_37916,N_30406,N_30738);
nand U37917 (N_37917,N_34313,N_34746);
and U37918 (N_37918,N_34536,N_32454);
and U37919 (N_37919,N_30628,N_34314);
nor U37920 (N_37920,N_30240,N_33500);
and U37921 (N_37921,N_32199,N_32315);
or U37922 (N_37922,N_34712,N_32080);
xnor U37923 (N_37923,N_31034,N_31851);
xor U37924 (N_37924,N_32434,N_34483);
or U37925 (N_37925,N_34854,N_31493);
or U37926 (N_37926,N_34064,N_34856);
or U37927 (N_37927,N_32158,N_32604);
nand U37928 (N_37928,N_30224,N_33049);
and U37929 (N_37929,N_34002,N_33766);
or U37930 (N_37930,N_33968,N_34027);
xor U37931 (N_37931,N_30047,N_31753);
or U37932 (N_37932,N_31853,N_34037);
nor U37933 (N_37933,N_33363,N_34055);
and U37934 (N_37934,N_31444,N_32168);
and U37935 (N_37935,N_34220,N_34084);
xnor U37936 (N_37936,N_32513,N_31847);
or U37937 (N_37937,N_33453,N_32761);
or U37938 (N_37938,N_31391,N_30946);
nand U37939 (N_37939,N_33083,N_30731);
nand U37940 (N_37940,N_30811,N_33070);
xnor U37941 (N_37941,N_31552,N_33601);
nand U37942 (N_37942,N_32133,N_31902);
nor U37943 (N_37943,N_31064,N_31875);
or U37944 (N_37944,N_32291,N_34150);
nor U37945 (N_37945,N_32436,N_33047);
xor U37946 (N_37946,N_33716,N_33887);
or U37947 (N_37947,N_32515,N_32445);
and U37948 (N_37948,N_33245,N_34429);
and U37949 (N_37949,N_31228,N_34431);
or U37950 (N_37950,N_33049,N_32398);
nand U37951 (N_37951,N_31219,N_31159);
xnor U37952 (N_37952,N_31383,N_34134);
nor U37953 (N_37953,N_34142,N_30026);
and U37954 (N_37954,N_33756,N_31830);
nor U37955 (N_37955,N_31118,N_31117);
nand U37956 (N_37956,N_32177,N_30046);
nand U37957 (N_37957,N_31623,N_32897);
nand U37958 (N_37958,N_31832,N_32899);
and U37959 (N_37959,N_33156,N_31776);
nand U37960 (N_37960,N_33109,N_32801);
or U37961 (N_37961,N_32426,N_31705);
xor U37962 (N_37962,N_32102,N_30650);
and U37963 (N_37963,N_32646,N_32537);
and U37964 (N_37964,N_30772,N_30739);
nor U37965 (N_37965,N_32585,N_32976);
nor U37966 (N_37966,N_32196,N_31915);
nand U37967 (N_37967,N_32695,N_34928);
or U37968 (N_37968,N_31166,N_34435);
and U37969 (N_37969,N_34029,N_34360);
and U37970 (N_37970,N_31162,N_34859);
or U37971 (N_37971,N_30064,N_31886);
or U37972 (N_37972,N_32604,N_31185);
nand U37973 (N_37973,N_30581,N_32937);
xnor U37974 (N_37974,N_31723,N_31044);
nor U37975 (N_37975,N_30010,N_34059);
xor U37976 (N_37976,N_34107,N_33196);
nand U37977 (N_37977,N_31192,N_34137);
and U37978 (N_37978,N_30609,N_30004);
nor U37979 (N_37979,N_34294,N_31237);
and U37980 (N_37980,N_31761,N_31932);
nand U37981 (N_37981,N_31527,N_33117);
xnor U37982 (N_37982,N_33119,N_34556);
nand U37983 (N_37983,N_32486,N_34491);
nor U37984 (N_37984,N_31744,N_33220);
nand U37985 (N_37985,N_30319,N_31304);
and U37986 (N_37986,N_30312,N_31726);
or U37987 (N_37987,N_34173,N_32365);
or U37988 (N_37988,N_31702,N_32503);
nor U37989 (N_37989,N_30799,N_31514);
xor U37990 (N_37990,N_32693,N_33987);
nor U37991 (N_37991,N_30298,N_30919);
xor U37992 (N_37992,N_33059,N_32288);
or U37993 (N_37993,N_30928,N_33129);
xnor U37994 (N_37994,N_32777,N_32011);
or U37995 (N_37995,N_34296,N_33411);
xor U37996 (N_37996,N_32576,N_34384);
xor U37997 (N_37997,N_34628,N_30510);
nor U37998 (N_37998,N_32806,N_30383);
nand U37999 (N_37999,N_32716,N_33509);
xor U38000 (N_38000,N_30868,N_33127);
nor U38001 (N_38001,N_32195,N_34297);
nand U38002 (N_38002,N_32779,N_30480);
and U38003 (N_38003,N_34081,N_32160);
or U38004 (N_38004,N_32204,N_33957);
or U38005 (N_38005,N_30474,N_33137);
nor U38006 (N_38006,N_33774,N_34486);
nand U38007 (N_38007,N_33931,N_30430);
nor U38008 (N_38008,N_33171,N_31964);
nor U38009 (N_38009,N_30463,N_30896);
xor U38010 (N_38010,N_30878,N_30640);
and U38011 (N_38011,N_34162,N_31037);
xnor U38012 (N_38012,N_31926,N_33845);
xor U38013 (N_38013,N_30472,N_30852);
nor U38014 (N_38014,N_32826,N_34575);
xnor U38015 (N_38015,N_32368,N_31247);
and U38016 (N_38016,N_32231,N_33192);
and U38017 (N_38017,N_33145,N_32441);
xor U38018 (N_38018,N_30715,N_30162);
xnor U38019 (N_38019,N_30907,N_31601);
nand U38020 (N_38020,N_32443,N_30774);
and U38021 (N_38021,N_30643,N_32113);
nand U38022 (N_38022,N_31205,N_31524);
and U38023 (N_38023,N_34294,N_31790);
nand U38024 (N_38024,N_34853,N_34923);
or U38025 (N_38025,N_31018,N_32920);
nand U38026 (N_38026,N_30668,N_31957);
and U38027 (N_38027,N_32777,N_31908);
or U38028 (N_38028,N_34827,N_34948);
and U38029 (N_38029,N_32724,N_34520);
nand U38030 (N_38030,N_31313,N_34076);
nand U38031 (N_38031,N_30585,N_31896);
xnor U38032 (N_38032,N_32191,N_33473);
nor U38033 (N_38033,N_31023,N_31326);
nor U38034 (N_38034,N_31275,N_31216);
or U38035 (N_38035,N_34249,N_34505);
xor U38036 (N_38036,N_32724,N_34609);
nand U38037 (N_38037,N_34328,N_34626);
xor U38038 (N_38038,N_33342,N_32162);
nand U38039 (N_38039,N_33963,N_34963);
nand U38040 (N_38040,N_34268,N_34733);
nand U38041 (N_38041,N_33767,N_31574);
or U38042 (N_38042,N_30204,N_32754);
or U38043 (N_38043,N_32043,N_33205);
nor U38044 (N_38044,N_34421,N_30140);
nor U38045 (N_38045,N_30682,N_33129);
nor U38046 (N_38046,N_30180,N_33674);
xnor U38047 (N_38047,N_31758,N_32888);
or U38048 (N_38048,N_31235,N_33384);
xor U38049 (N_38049,N_33709,N_32786);
nor U38050 (N_38050,N_31988,N_31630);
and U38051 (N_38051,N_33044,N_34374);
nor U38052 (N_38052,N_33101,N_31805);
xor U38053 (N_38053,N_31692,N_32838);
xnor U38054 (N_38054,N_31884,N_32743);
and U38055 (N_38055,N_32657,N_32953);
and U38056 (N_38056,N_30652,N_31324);
nor U38057 (N_38057,N_32664,N_33709);
and U38058 (N_38058,N_31163,N_32969);
nor U38059 (N_38059,N_32869,N_33688);
or U38060 (N_38060,N_33214,N_34128);
nand U38061 (N_38061,N_32266,N_34899);
nor U38062 (N_38062,N_30255,N_31084);
xor U38063 (N_38063,N_33910,N_32868);
and U38064 (N_38064,N_30657,N_34609);
and U38065 (N_38065,N_30908,N_34327);
and U38066 (N_38066,N_32829,N_33592);
or U38067 (N_38067,N_33369,N_34499);
or U38068 (N_38068,N_34852,N_34517);
and U38069 (N_38069,N_32200,N_33746);
nor U38070 (N_38070,N_33810,N_33272);
and U38071 (N_38071,N_32484,N_30704);
nand U38072 (N_38072,N_32525,N_33145);
nand U38073 (N_38073,N_34410,N_33577);
xor U38074 (N_38074,N_30309,N_31245);
or U38075 (N_38075,N_31548,N_32250);
nor U38076 (N_38076,N_31825,N_33290);
and U38077 (N_38077,N_30568,N_32590);
nand U38078 (N_38078,N_31459,N_34622);
or U38079 (N_38079,N_31369,N_34424);
or U38080 (N_38080,N_30240,N_30916);
or U38081 (N_38081,N_30316,N_32430);
and U38082 (N_38082,N_33312,N_32051);
nand U38083 (N_38083,N_33068,N_34204);
nand U38084 (N_38084,N_32902,N_33293);
and U38085 (N_38085,N_34053,N_33305);
nor U38086 (N_38086,N_33384,N_31202);
and U38087 (N_38087,N_34340,N_32738);
nand U38088 (N_38088,N_33041,N_32843);
nor U38089 (N_38089,N_30020,N_30925);
nor U38090 (N_38090,N_34414,N_34850);
or U38091 (N_38091,N_32905,N_33865);
and U38092 (N_38092,N_32301,N_30326);
nand U38093 (N_38093,N_34743,N_33062);
and U38094 (N_38094,N_33101,N_34123);
xor U38095 (N_38095,N_33176,N_32282);
and U38096 (N_38096,N_30216,N_30909);
nand U38097 (N_38097,N_33370,N_30310);
nor U38098 (N_38098,N_32510,N_30402);
nor U38099 (N_38099,N_33906,N_30495);
nor U38100 (N_38100,N_33013,N_34524);
and U38101 (N_38101,N_30884,N_34609);
xnor U38102 (N_38102,N_32717,N_30226);
xor U38103 (N_38103,N_30235,N_30922);
nand U38104 (N_38104,N_34878,N_30541);
nor U38105 (N_38105,N_30000,N_33124);
and U38106 (N_38106,N_34526,N_34039);
nor U38107 (N_38107,N_30730,N_33970);
or U38108 (N_38108,N_34540,N_30163);
or U38109 (N_38109,N_31955,N_30078);
nand U38110 (N_38110,N_31550,N_30408);
or U38111 (N_38111,N_34915,N_34261);
nor U38112 (N_38112,N_32112,N_31992);
nand U38113 (N_38113,N_34471,N_33711);
nor U38114 (N_38114,N_31774,N_33531);
and U38115 (N_38115,N_33095,N_32593);
and U38116 (N_38116,N_33109,N_33997);
or U38117 (N_38117,N_33573,N_32512);
nand U38118 (N_38118,N_34211,N_33355);
or U38119 (N_38119,N_30541,N_30477);
nor U38120 (N_38120,N_30141,N_30995);
xor U38121 (N_38121,N_31391,N_33201);
or U38122 (N_38122,N_34638,N_30632);
xnor U38123 (N_38123,N_30235,N_32405);
and U38124 (N_38124,N_32880,N_32437);
nand U38125 (N_38125,N_30315,N_34041);
nor U38126 (N_38126,N_32718,N_32148);
and U38127 (N_38127,N_32592,N_34900);
nor U38128 (N_38128,N_32858,N_32719);
and U38129 (N_38129,N_31958,N_30821);
or U38130 (N_38130,N_30870,N_32730);
nand U38131 (N_38131,N_32503,N_31903);
or U38132 (N_38132,N_31504,N_33626);
nor U38133 (N_38133,N_30099,N_31058);
nor U38134 (N_38134,N_34862,N_33670);
and U38135 (N_38135,N_31484,N_34089);
nand U38136 (N_38136,N_32151,N_30298);
nand U38137 (N_38137,N_30827,N_33620);
nand U38138 (N_38138,N_33244,N_31279);
xor U38139 (N_38139,N_30472,N_33178);
or U38140 (N_38140,N_33858,N_34082);
nand U38141 (N_38141,N_34985,N_30834);
xnor U38142 (N_38142,N_31802,N_30306);
and U38143 (N_38143,N_30207,N_34551);
xor U38144 (N_38144,N_32314,N_31411);
nor U38145 (N_38145,N_32042,N_32708);
or U38146 (N_38146,N_30228,N_33044);
or U38147 (N_38147,N_34389,N_34439);
and U38148 (N_38148,N_32168,N_34248);
xnor U38149 (N_38149,N_34662,N_30763);
nand U38150 (N_38150,N_30302,N_31233);
nor U38151 (N_38151,N_30000,N_34147);
xnor U38152 (N_38152,N_34977,N_31196);
xnor U38153 (N_38153,N_33325,N_31869);
or U38154 (N_38154,N_31610,N_34655);
nor U38155 (N_38155,N_32600,N_31494);
and U38156 (N_38156,N_33531,N_34071);
and U38157 (N_38157,N_32932,N_32456);
nor U38158 (N_38158,N_31432,N_33045);
and U38159 (N_38159,N_32600,N_31252);
xor U38160 (N_38160,N_31674,N_32885);
nor U38161 (N_38161,N_30301,N_34594);
nor U38162 (N_38162,N_30074,N_33103);
nand U38163 (N_38163,N_32449,N_32243);
xnor U38164 (N_38164,N_32323,N_34075);
xor U38165 (N_38165,N_31259,N_34056);
and U38166 (N_38166,N_30079,N_31740);
nand U38167 (N_38167,N_34726,N_34537);
nand U38168 (N_38168,N_31591,N_30607);
nor U38169 (N_38169,N_30740,N_30948);
or U38170 (N_38170,N_33364,N_31361);
nor U38171 (N_38171,N_34656,N_34767);
nand U38172 (N_38172,N_34991,N_31290);
and U38173 (N_38173,N_33911,N_31697);
xnor U38174 (N_38174,N_33520,N_33101);
xnor U38175 (N_38175,N_31200,N_30602);
or U38176 (N_38176,N_31536,N_33097);
nand U38177 (N_38177,N_31105,N_34085);
nor U38178 (N_38178,N_30416,N_34541);
and U38179 (N_38179,N_34399,N_32635);
and U38180 (N_38180,N_31096,N_32678);
xor U38181 (N_38181,N_34603,N_33534);
xnor U38182 (N_38182,N_34400,N_33859);
xnor U38183 (N_38183,N_33957,N_31877);
nand U38184 (N_38184,N_34774,N_34084);
nand U38185 (N_38185,N_34661,N_31651);
nor U38186 (N_38186,N_30884,N_31904);
xor U38187 (N_38187,N_32713,N_34428);
or U38188 (N_38188,N_33152,N_32367);
or U38189 (N_38189,N_33360,N_34534);
nand U38190 (N_38190,N_33000,N_33298);
nor U38191 (N_38191,N_34054,N_31672);
nor U38192 (N_38192,N_33343,N_32162);
nor U38193 (N_38193,N_33133,N_33783);
and U38194 (N_38194,N_31716,N_31134);
xnor U38195 (N_38195,N_33136,N_30747);
nor U38196 (N_38196,N_32988,N_30812);
and U38197 (N_38197,N_31778,N_30661);
nor U38198 (N_38198,N_31562,N_31133);
xnor U38199 (N_38199,N_33924,N_32270);
and U38200 (N_38200,N_30185,N_31586);
or U38201 (N_38201,N_32117,N_31555);
xor U38202 (N_38202,N_30517,N_30762);
nand U38203 (N_38203,N_30962,N_33349);
or U38204 (N_38204,N_34300,N_34516);
nor U38205 (N_38205,N_31970,N_33562);
xor U38206 (N_38206,N_33917,N_32419);
and U38207 (N_38207,N_31447,N_34784);
xnor U38208 (N_38208,N_30042,N_30251);
nor U38209 (N_38209,N_30717,N_33600);
xnor U38210 (N_38210,N_32341,N_32331);
and U38211 (N_38211,N_31672,N_32063);
nor U38212 (N_38212,N_33464,N_34940);
and U38213 (N_38213,N_33062,N_34390);
xnor U38214 (N_38214,N_34721,N_34396);
nor U38215 (N_38215,N_32333,N_31906);
or U38216 (N_38216,N_30042,N_33137);
xnor U38217 (N_38217,N_33288,N_34428);
xnor U38218 (N_38218,N_30176,N_32298);
xor U38219 (N_38219,N_31399,N_33522);
nand U38220 (N_38220,N_31047,N_31441);
or U38221 (N_38221,N_31008,N_30312);
or U38222 (N_38222,N_31177,N_33157);
xor U38223 (N_38223,N_32817,N_33373);
nor U38224 (N_38224,N_30463,N_30684);
or U38225 (N_38225,N_30245,N_31584);
xnor U38226 (N_38226,N_30278,N_34928);
or U38227 (N_38227,N_32178,N_34320);
nand U38228 (N_38228,N_34917,N_30893);
nand U38229 (N_38229,N_34381,N_30891);
xor U38230 (N_38230,N_30900,N_32315);
nor U38231 (N_38231,N_34653,N_34280);
and U38232 (N_38232,N_31388,N_34405);
or U38233 (N_38233,N_31547,N_31034);
xor U38234 (N_38234,N_32955,N_32293);
nor U38235 (N_38235,N_31632,N_33246);
nand U38236 (N_38236,N_32822,N_32178);
nand U38237 (N_38237,N_33342,N_33517);
or U38238 (N_38238,N_33923,N_32018);
nor U38239 (N_38239,N_34402,N_33202);
nand U38240 (N_38240,N_34912,N_30146);
xor U38241 (N_38241,N_30455,N_30336);
nor U38242 (N_38242,N_30774,N_34827);
nand U38243 (N_38243,N_31833,N_34473);
nor U38244 (N_38244,N_34978,N_34381);
and U38245 (N_38245,N_33116,N_31806);
nand U38246 (N_38246,N_33201,N_34907);
nor U38247 (N_38247,N_32363,N_30994);
xor U38248 (N_38248,N_32565,N_34356);
and U38249 (N_38249,N_32804,N_30801);
nor U38250 (N_38250,N_33346,N_33844);
xor U38251 (N_38251,N_32061,N_32986);
xnor U38252 (N_38252,N_31658,N_33824);
or U38253 (N_38253,N_32921,N_31253);
xor U38254 (N_38254,N_33902,N_31319);
and U38255 (N_38255,N_33936,N_30905);
nand U38256 (N_38256,N_34605,N_30113);
nor U38257 (N_38257,N_34151,N_31038);
or U38258 (N_38258,N_31246,N_30467);
and U38259 (N_38259,N_34543,N_30145);
xor U38260 (N_38260,N_32641,N_33562);
xnor U38261 (N_38261,N_31295,N_31800);
and U38262 (N_38262,N_32207,N_34873);
nand U38263 (N_38263,N_30878,N_30847);
and U38264 (N_38264,N_30673,N_33526);
or U38265 (N_38265,N_32189,N_30255);
xor U38266 (N_38266,N_33170,N_34065);
and U38267 (N_38267,N_31721,N_33438);
or U38268 (N_38268,N_33532,N_32389);
nand U38269 (N_38269,N_32183,N_34915);
nor U38270 (N_38270,N_33347,N_30089);
nand U38271 (N_38271,N_31452,N_31112);
xnor U38272 (N_38272,N_33269,N_32410);
nor U38273 (N_38273,N_32065,N_32080);
xor U38274 (N_38274,N_33794,N_34293);
and U38275 (N_38275,N_33882,N_32110);
xnor U38276 (N_38276,N_32477,N_33551);
nand U38277 (N_38277,N_34300,N_34475);
or U38278 (N_38278,N_30537,N_33909);
nand U38279 (N_38279,N_31624,N_34330);
and U38280 (N_38280,N_33641,N_33091);
and U38281 (N_38281,N_33657,N_34562);
xnor U38282 (N_38282,N_32165,N_31830);
xnor U38283 (N_38283,N_30488,N_32783);
and U38284 (N_38284,N_32830,N_32436);
nand U38285 (N_38285,N_33655,N_33383);
nand U38286 (N_38286,N_30041,N_31056);
nor U38287 (N_38287,N_32893,N_31031);
nand U38288 (N_38288,N_30015,N_33645);
xor U38289 (N_38289,N_30947,N_32115);
nand U38290 (N_38290,N_31830,N_31449);
or U38291 (N_38291,N_32215,N_34620);
or U38292 (N_38292,N_30426,N_31832);
nand U38293 (N_38293,N_31680,N_30928);
or U38294 (N_38294,N_30563,N_30631);
nor U38295 (N_38295,N_32295,N_34263);
and U38296 (N_38296,N_33625,N_34621);
or U38297 (N_38297,N_32786,N_31955);
xor U38298 (N_38298,N_30520,N_31458);
or U38299 (N_38299,N_34483,N_34009);
xor U38300 (N_38300,N_34200,N_31671);
xnor U38301 (N_38301,N_34466,N_30223);
nand U38302 (N_38302,N_34311,N_33786);
and U38303 (N_38303,N_32300,N_30455);
xnor U38304 (N_38304,N_34484,N_34523);
nor U38305 (N_38305,N_32771,N_31038);
nand U38306 (N_38306,N_34290,N_33537);
nor U38307 (N_38307,N_33765,N_31785);
nand U38308 (N_38308,N_33738,N_33498);
nor U38309 (N_38309,N_34535,N_31146);
nor U38310 (N_38310,N_34072,N_34229);
and U38311 (N_38311,N_33999,N_31553);
nand U38312 (N_38312,N_32662,N_32871);
nor U38313 (N_38313,N_33505,N_32292);
xnor U38314 (N_38314,N_32615,N_32322);
and U38315 (N_38315,N_30611,N_33735);
nor U38316 (N_38316,N_33702,N_30955);
xnor U38317 (N_38317,N_32476,N_33524);
xnor U38318 (N_38318,N_31523,N_31856);
xor U38319 (N_38319,N_34734,N_33333);
or U38320 (N_38320,N_34233,N_31404);
and U38321 (N_38321,N_32530,N_34091);
nor U38322 (N_38322,N_31853,N_31579);
nand U38323 (N_38323,N_31310,N_32959);
nor U38324 (N_38324,N_33864,N_32532);
nand U38325 (N_38325,N_31565,N_30162);
nand U38326 (N_38326,N_33623,N_31801);
or U38327 (N_38327,N_30200,N_31000);
nand U38328 (N_38328,N_31503,N_31222);
nand U38329 (N_38329,N_34295,N_34091);
nand U38330 (N_38330,N_31926,N_31251);
and U38331 (N_38331,N_33574,N_32544);
or U38332 (N_38332,N_31630,N_32390);
xor U38333 (N_38333,N_32669,N_31438);
xor U38334 (N_38334,N_30546,N_32260);
nand U38335 (N_38335,N_33459,N_32178);
nor U38336 (N_38336,N_31593,N_34508);
nor U38337 (N_38337,N_34027,N_34230);
nand U38338 (N_38338,N_31284,N_33669);
xor U38339 (N_38339,N_32489,N_32933);
nor U38340 (N_38340,N_30203,N_30932);
nand U38341 (N_38341,N_30738,N_31581);
xor U38342 (N_38342,N_31862,N_34055);
xor U38343 (N_38343,N_33200,N_33215);
nor U38344 (N_38344,N_30930,N_32409);
nand U38345 (N_38345,N_34484,N_34508);
nand U38346 (N_38346,N_34290,N_32505);
xor U38347 (N_38347,N_30873,N_34737);
and U38348 (N_38348,N_33389,N_33927);
nor U38349 (N_38349,N_32327,N_32139);
or U38350 (N_38350,N_34633,N_33384);
and U38351 (N_38351,N_32830,N_31305);
nand U38352 (N_38352,N_34591,N_33092);
nand U38353 (N_38353,N_30458,N_30510);
and U38354 (N_38354,N_30102,N_30147);
nor U38355 (N_38355,N_34577,N_32340);
nand U38356 (N_38356,N_34356,N_33292);
and U38357 (N_38357,N_31201,N_31290);
nand U38358 (N_38358,N_30229,N_34185);
and U38359 (N_38359,N_32223,N_34760);
nand U38360 (N_38360,N_32288,N_32682);
xnor U38361 (N_38361,N_33036,N_31190);
nand U38362 (N_38362,N_31971,N_32160);
xnor U38363 (N_38363,N_33086,N_34693);
nand U38364 (N_38364,N_30094,N_30665);
and U38365 (N_38365,N_34248,N_32659);
nor U38366 (N_38366,N_30931,N_34430);
nor U38367 (N_38367,N_30527,N_33297);
nand U38368 (N_38368,N_34030,N_30498);
and U38369 (N_38369,N_34181,N_30104);
and U38370 (N_38370,N_33919,N_34815);
nand U38371 (N_38371,N_31938,N_31335);
nand U38372 (N_38372,N_31277,N_32547);
xnor U38373 (N_38373,N_30539,N_34325);
nand U38374 (N_38374,N_33326,N_31014);
nand U38375 (N_38375,N_31039,N_31264);
and U38376 (N_38376,N_30466,N_30162);
nor U38377 (N_38377,N_34544,N_30016);
nor U38378 (N_38378,N_32653,N_31582);
and U38379 (N_38379,N_30104,N_34308);
xnor U38380 (N_38380,N_30960,N_31304);
xor U38381 (N_38381,N_33371,N_33291);
nand U38382 (N_38382,N_32043,N_31503);
and U38383 (N_38383,N_33361,N_32107);
nand U38384 (N_38384,N_34517,N_34606);
nor U38385 (N_38385,N_34324,N_34443);
and U38386 (N_38386,N_34111,N_34298);
and U38387 (N_38387,N_33107,N_31565);
nand U38388 (N_38388,N_32387,N_32930);
nand U38389 (N_38389,N_33734,N_31050);
and U38390 (N_38390,N_30098,N_34651);
and U38391 (N_38391,N_30456,N_30641);
or U38392 (N_38392,N_32282,N_33636);
or U38393 (N_38393,N_31138,N_34495);
xor U38394 (N_38394,N_33304,N_30003);
xnor U38395 (N_38395,N_32792,N_33206);
and U38396 (N_38396,N_30348,N_32631);
xnor U38397 (N_38397,N_30827,N_32325);
or U38398 (N_38398,N_32334,N_33301);
and U38399 (N_38399,N_33613,N_31647);
and U38400 (N_38400,N_31096,N_31965);
nor U38401 (N_38401,N_32280,N_34142);
or U38402 (N_38402,N_33915,N_30107);
nand U38403 (N_38403,N_30193,N_34378);
and U38404 (N_38404,N_33174,N_30992);
nor U38405 (N_38405,N_31201,N_30281);
or U38406 (N_38406,N_34875,N_30048);
xor U38407 (N_38407,N_33927,N_30713);
nand U38408 (N_38408,N_30733,N_34692);
and U38409 (N_38409,N_32127,N_30885);
nor U38410 (N_38410,N_32938,N_32208);
nand U38411 (N_38411,N_33416,N_33118);
nand U38412 (N_38412,N_32193,N_30001);
xnor U38413 (N_38413,N_31001,N_31367);
nor U38414 (N_38414,N_34317,N_30756);
nand U38415 (N_38415,N_30397,N_30316);
or U38416 (N_38416,N_31945,N_33166);
xor U38417 (N_38417,N_33128,N_33665);
nor U38418 (N_38418,N_34639,N_34948);
and U38419 (N_38419,N_34030,N_33124);
nor U38420 (N_38420,N_34851,N_32776);
nor U38421 (N_38421,N_30519,N_30864);
nor U38422 (N_38422,N_34804,N_34992);
nor U38423 (N_38423,N_30323,N_30091);
or U38424 (N_38424,N_33995,N_33889);
or U38425 (N_38425,N_30873,N_31350);
nor U38426 (N_38426,N_34089,N_31012);
xnor U38427 (N_38427,N_34240,N_34734);
and U38428 (N_38428,N_31898,N_33321);
nor U38429 (N_38429,N_32041,N_33432);
or U38430 (N_38430,N_33541,N_31753);
nand U38431 (N_38431,N_31886,N_30759);
or U38432 (N_38432,N_32105,N_31869);
xnor U38433 (N_38433,N_33798,N_31581);
xor U38434 (N_38434,N_31761,N_31183);
nor U38435 (N_38435,N_33133,N_31111);
nand U38436 (N_38436,N_33942,N_30949);
nand U38437 (N_38437,N_32409,N_34709);
xnor U38438 (N_38438,N_33674,N_30943);
nor U38439 (N_38439,N_33083,N_34091);
or U38440 (N_38440,N_33641,N_33023);
and U38441 (N_38441,N_31987,N_33960);
nand U38442 (N_38442,N_33041,N_30641);
nor U38443 (N_38443,N_34010,N_34732);
nand U38444 (N_38444,N_32745,N_30464);
nand U38445 (N_38445,N_34482,N_31568);
nand U38446 (N_38446,N_30470,N_32376);
or U38447 (N_38447,N_33735,N_30188);
xor U38448 (N_38448,N_34406,N_30994);
or U38449 (N_38449,N_30162,N_32952);
and U38450 (N_38450,N_32474,N_30137);
or U38451 (N_38451,N_32786,N_32781);
nand U38452 (N_38452,N_34454,N_31305);
or U38453 (N_38453,N_34093,N_34292);
nor U38454 (N_38454,N_30906,N_33093);
nand U38455 (N_38455,N_34177,N_34484);
xnor U38456 (N_38456,N_32076,N_31038);
nand U38457 (N_38457,N_32589,N_32659);
nand U38458 (N_38458,N_30250,N_33033);
nor U38459 (N_38459,N_31183,N_33715);
xor U38460 (N_38460,N_30017,N_30613);
nand U38461 (N_38461,N_34659,N_32841);
xor U38462 (N_38462,N_34312,N_32758);
nand U38463 (N_38463,N_30119,N_31560);
nor U38464 (N_38464,N_30895,N_31120);
nand U38465 (N_38465,N_30063,N_34807);
or U38466 (N_38466,N_30639,N_31754);
nand U38467 (N_38467,N_30074,N_31022);
nand U38468 (N_38468,N_33262,N_31762);
or U38469 (N_38469,N_33432,N_32152);
nor U38470 (N_38470,N_34569,N_33667);
nor U38471 (N_38471,N_30513,N_34307);
or U38472 (N_38472,N_32173,N_33606);
or U38473 (N_38473,N_31616,N_33315);
xnor U38474 (N_38474,N_32468,N_31710);
xnor U38475 (N_38475,N_33701,N_34672);
nor U38476 (N_38476,N_32748,N_34147);
xnor U38477 (N_38477,N_32925,N_32151);
nor U38478 (N_38478,N_32791,N_33312);
nor U38479 (N_38479,N_31129,N_31253);
nand U38480 (N_38480,N_34758,N_30187);
nand U38481 (N_38481,N_30966,N_30075);
nor U38482 (N_38482,N_30893,N_34798);
nand U38483 (N_38483,N_30403,N_33812);
or U38484 (N_38484,N_30023,N_31203);
xor U38485 (N_38485,N_31357,N_33015);
nand U38486 (N_38486,N_31061,N_31419);
and U38487 (N_38487,N_32384,N_34302);
nand U38488 (N_38488,N_32287,N_30871);
and U38489 (N_38489,N_31978,N_32207);
xor U38490 (N_38490,N_33782,N_31374);
or U38491 (N_38491,N_30284,N_34455);
or U38492 (N_38492,N_34240,N_34519);
nor U38493 (N_38493,N_34336,N_32337);
xnor U38494 (N_38494,N_34075,N_34542);
nor U38495 (N_38495,N_31239,N_34097);
nor U38496 (N_38496,N_33312,N_31695);
and U38497 (N_38497,N_34299,N_30099);
nor U38498 (N_38498,N_33237,N_33469);
nand U38499 (N_38499,N_30596,N_30678);
or U38500 (N_38500,N_34422,N_33251);
xor U38501 (N_38501,N_34302,N_30203);
nor U38502 (N_38502,N_32848,N_31658);
nand U38503 (N_38503,N_31464,N_30191);
nand U38504 (N_38504,N_32423,N_30206);
and U38505 (N_38505,N_33640,N_33014);
nand U38506 (N_38506,N_33001,N_31335);
xor U38507 (N_38507,N_33510,N_31006);
or U38508 (N_38508,N_31016,N_30096);
nand U38509 (N_38509,N_33137,N_33393);
xor U38510 (N_38510,N_31798,N_30294);
and U38511 (N_38511,N_30688,N_30587);
nor U38512 (N_38512,N_30641,N_33611);
and U38513 (N_38513,N_34302,N_31126);
nor U38514 (N_38514,N_31959,N_34852);
nand U38515 (N_38515,N_33009,N_31624);
and U38516 (N_38516,N_31617,N_32162);
and U38517 (N_38517,N_34199,N_33984);
or U38518 (N_38518,N_30453,N_33027);
xor U38519 (N_38519,N_34797,N_34128);
or U38520 (N_38520,N_34366,N_32814);
or U38521 (N_38521,N_33643,N_30059);
nand U38522 (N_38522,N_33402,N_34541);
nor U38523 (N_38523,N_33687,N_32453);
nor U38524 (N_38524,N_30664,N_34074);
and U38525 (N_38525,N_33674,N_31256);
nor U38526 (N_38526,N_30825,N_32697);
nand U38527 (N_38527,N_33122,N_34388);
xnor U38528 (N_38528,N_33375,N_30926);
and U38529 (N_38529,N_34611,N_31392);
or U38530 (N_38530,N_33990,N_30692);
nand U38531 (N_38531,N_31422,N_30863);
nand U38532 (N_38532,N_34479,N_31612);
xnor U38533 (N_38533,N_32940,N_32076);
nand U38534 (N_38534,N_34237,N_32987);
or U38535 (N_38535,N_32406,N_32861);
nand U38536 (N_38536,N_33936,N_33040);
and U38537 (N_38537,N_33693,N_33735);
xor U38538 (N_38538,N_32316,N_32032);
and U38539 (N_38539,N_32193,N_34089);
xnor U38540 (N_38540,N_33632,N_31065);
nor U38541 (N_38541,N_33734,N_31025);
or U38542 (N_38542,N_30691,N_34687);
xor U38543 (N_38543,N_33349,N_30646);
xor U38544 (N_38544,N_31796,N_32667);
nand U38545 (N_38545,N_32856,N_31509);
xnor U38546 (N_38546,N_32376,N_30260);
xor U38547 (N_38547,N_31089,N_30002);
nand U38548 (N_38548,N_33581,N_32258);
nor U38549 (N_38549,N_30473,N_33044);
nor U38550 (N_38550,N_32404,N_34026);
and U38551 (N_38551,N_32694,N_32415);
and U38552 (N_38552,N_32050,N_31819);
nand U38553 (N_38553,N_34934,N_31290);
nor U38554 (N_38554,N_30990,N_33722);
nor U38555 (N_38555,N_34022,N_30668);
or U38556 (N_38556,N_31191,N_34798);
nand U38557 (N_38557,N_33612,N_31689);
nor U38558 (N_38558,N_32408,N_32032);
or U38559 (N_38559,N_31743,N_31375);
or U38560 (N_38560,N_31592,N_30719);
nor U38561 (N_38561,N_33671,N_32719);
or U38562 (N_38562,N_30333,N_33556);
nor U38563 (N_38563,N_33821,N_32865);
nand U38564 (N_38564,N_33204,N_34757);
xor U38565 (N_38565,N_31005,N_30934);
or U38566 (N_38566,N_33815,N_31601);
nor U38567 (N_38567,N_32399,N_30413);
or U38568 (N_38568,N_30343,N_34116);
nand U38569 (N_38569,N_32613,N_34050);
nand U38570 (N_38570,N_31827,N_33602);
and U38571 (N_38571,N_30748,N_32140);
nand U38572 (N_38572,N_30115,N_34648);
nand U38573 (N_38573,N_30232,N_34577);
nand U38574 (N_38574,N_31214,N_30203);
and U38575 (N_38575,N_34180,N_30843);
xnor U38576 (N_38576,N_32711,N_33317);
xor U38577 (N_38577,N_34669,N_33283);
xor U38578 (N_38578,N_34925,N_31499);
and U38579 (N_38579,N_34905,N_33762);
nand U38580 (N_38580,N_32420,N_32707);
and U38581 (N_38581,N_33425,N_31412);
nand U38582 (N_38582,N_32479,N_32849);
xor U38583 (N_38583,N_34026,N_33302);
xor U38584 (N_38584,N_33806,N_30125);
nand U38585 (N_38585,N_34934,N_31256);
xor U38586 (N_38586,N_34178,N_31456);
xnor U38587 (N_38587,N_34762,N_34898);
nor U38588 (N_38588,N_34436,N_33903);
nand U38589 (N_38589,N_33183,N_33434);
and U38590 (N_38590,N_31094,N_31250);
xor U38591 (N_38591,N_33576,N_31852);
or U38592 (N_38592,N_34660,N_33759);
nor U38593 (N_38593,N_33738,N_32261);
xor U38594 (N_38594,N_31742,N_30693);
xnor U38595 (N_38595,N_33576,N_34718);
nand U38596 (N_38596,N_31853,N_32243);
nand U38597 (N_38597,N_33575,N_33430);
or U38598 (N_38598,N_33093,N_34318);
or U38599 (N_38599,N_30903,N_33195);
nor U38600 (N_38600,N_33092,N_31684);
and U38601 (N_38601,N_34075,N_33859);
and U38602 (N_38602,N_33165,N_32809);
xnor U38603 (N_38603,N_30673,N_31296);
xnor U38604 (N_38604,N_34960,N_34582);
and U38605 (N_38605,N_34464,N_34889);
and U38606 (N_38606,N_30689,N_31552);
xor U38607 (N_38607,N_32750,N_31986);
or U38608 (N_38608,N_33678,N_31153);
or U38609 (N_38609,N_32645,N_34825);
and U38610 (N_38610,N_32441,N_30480);
or U38611 (N_38611,N_31750,N_30726);
or U38612 (N_38612,N_31805,N_34817);
and U38613 (N_38613,N_34091,N_31983);
nand U38614 (N_38614,N_34258,N_33681);
or U38615 (N_38615,N_31623,N_30330);
and U38616 (N_38616,N_33259,N_31619);
nand U38617 (N_38617,N_33346,N_32024);
and U38618 (N_38618,N_32922,N_30063);
and U38619 (N_38619,N_34724,N_30647);
xor U38620 (N_38620,N_33970,N_31089);
or U38621 (N_38621,N_30498,N_34779);
nor U38622 (N_38622,N_34178,N_31660);
or U38623 (N_38623,N_32456,N_33361);
or U38624 (N_38624,N_34804,N_30608);
nor U38625 (N_38625,N_34299,N_32021);
nand U38626 (N_38626,N_34780,N_34471);
or U38627 (N_38627,N_30092,N_30774);
and U38628 (N_38628,N_34974,N_34199);
and U38629 (N_38629,N_30650,N_30460);
nand U38630 (N_38630,N_34202,N_34272);
and U38631 (N_38631,N_32856,N_33079);
or U38632 (N_38632,N_34159,N_32811);
nand U38633 (N_38633,N_30771,N_30761);
nand U38634 (N_38634,N_33781,N_30038);
nor U38635 (N_38635,N_32044,N_32375);
or U38636 (N_38636,N_33354,N_30913);
xnor U38637 (N_38637,N_32840,N_32776);
or U38638 (N_38638,N_32653,N_32854);
nor U38639 (N_38639,N_33572,N_31002);
nor U38640 (N_38640,N_31400,N_31034);
xnor U38641 (N_38641,N_34703,N_32279);
nand U38642 (N_38642,N_33845,N_32252);
and U38643 (N_38643,N_31126,N_31908);
nor U38644 (N_38644,N_31699,N_32954);
or U38645 (N_38645,N_34136,N_32726);
or U38646 (N_38646,N_31299,N_34948);
or U38647 (N_38647,N_34275,N_33934);
xnor U38648 (N_38648,N_31935,N_32912);
nand U38649 (N_38649,N_31100,N_34919);
and U38650 (N_38650,N_34400,N_32232);
and U38651 (N_38651,N_31118,N_34927);
nand U38652 (N_38652,N_33066,N_34457);
xor U38653 (N_38653,N_30106,N_30168);
and U38654 (N_38654,N_32542,N_33380);
xor U38655 (N_38655,N_31883,N_34454);
or U38656 (N_38656,N_32669,N_31211);
xnor U38657 (N_38657,N_34199,N_34133);
xor U38658 (N_38658,N_31155,N_32106);
xnor U38659 (N_38659,N_34035,N_30071);
and U38660 (N_38660,N_33416,N_32944);
xor U38661 (N_38661,N_33122,N_34781);
nand U38662 (N_38662,N_31906,N_31665);
or U38663 (N_38663,N_32307,N_33391);
nor U38664 (N_38664,N_31703,N_31418);
xor U38665 (N_38665,N_33483,N_33817);
nor U38666 (N_38666,N_34808,N_30466);
nand U38667 (N_38667,N_30221,N_30011);
nor U38668 (N_38668,N_31445,N_30672);
or U38669 (N_38669,N_30983,N_31472);
and U38670 (N_38670,N_32180,N_34975);
xor U38671 (N_38671,N_31563,N_33555);
or U38672 (N_38672,N_34407,N_30138);
xor U38673 (N_38673,N_30422,N_34288);
and U38674 (N_38674,N_31060,N_30644);
or U38675 (N_38675,N_30411,N_31649);
or U38676 (N_38676,N_32053,N_33321);
xor U38677 (N_38677,N_30254,N_34782);
or U38678 (N_38678,N_33646,N_34350);
nand U38679 (N_38679,N_34028,N_32540);
xnor U38680 (N_38680,N_32890,N_32009);
and U38681 (N_38681,N_32096,N_34454);
nand U38682 (N_38682,N_34768,N_31518);
and U38683 (N_38683,N_32901,N_30098);
nand U38684 (N_38684,N_34455,N_33512);
xnor U38685 (N_38685,N_30519,N_33499);
nor U38686 (N_38686,N_30918,N_33105);
or U38687 (N_38687,N_31379,N_34025);
and U38688 (N_38688,N_30047,N_31009);
or U38689 (N_38689,N_30229,N_34944);
xor U38690 (N_38690,N_30580,N_34779);
xor U38691 (N_38691,N_32112,N_33186);
or U38692 (N_38692,N_33923,N_34865);
xor U38693 (N_38693,N_31531,N_34523);
nand U38694 (N_38694,N_34404,N_32893);
or U38695 (N_38695,N_32721,N_30604);
and U38696 (N_38696,N_31809,N_34173);
or U38697 (N_38697,N_32063,N_33155);
xor U38698 (N_38698,N_33117,N_33578);
and U38699 (N_38699,N_33284,N_32646);
xor U38700 (N_38700,N_32174,N_32627);
xnor U38701 (N_38701,N_31272,N_32733);
nand U38702 (N_38702,N_31402,N_32895);
and U38703 (N_38703,N_31792,N_34463);
xor U38704 (N_38704,N_33103,N_32755);
nand U38705 (N_38705,N_33054,N_33475);
xor U38706 (N_38706,N_33280,N_31092);
nand U38707 (N_38707,N_33844,N_30062);
and U38708 (N_38708,N_32097,N_31837);
and U38709 (N_38709,N_34549,N_31031);
xnor U38710 (N_38710,N_32352,N_33639);
nand U38711 (N_38711,N_31844,N_31020);
and U38712 (N_38712,N_33061,N_33995);
and U38713 (N_38713,N_33006,N_31089);
or U38714 (N_38714,N_31278,N_33381);
xor U38715 (N_38715,N_32726,N_34353);
and U38716 (N_38716,N_33314,N_34959);
nor U38717 (N_38717,N_34645,N_31022);
xnor U38718 (N_38718,N_31792,N_34226);
nor U38719 (N_38719,N_34837,N_32889);
or U38720 (N_38720,N_30965,N_30109);
xor U38721 (N_38721,N_34247,N_32023);
nor U38722 (N_38722,N_34452,N_32934);
nor U38723 (N_38723,N_32540,N_34791);
nand U38724 (N_38724,N_31706,N_32399);
and U38725 (N_38725,N_32213,N_30743);
and U38726 (N_38726,N_30766,N_34002);
nor U38727 (N_38727,N_32486,N_32022);
xor U38728 (N_38728,N_33829,N_31380);
nor U38729 (N_38729,N_33959,N_33809);
nor U38730 (N_38730,N_31036,N_32443);
and U38731 (N_38731,N_34759,N_31348);
xnor U38732 (N_38732,N_31194,N_30993);
or U38733 (N_38733,N_30460,N_34052);
and U38734 (N_38734,N_34401,N_30028);
and U38735 (N_38735,N_34791,N_33666);
nand U38736 (N_38736,N_34829,N_31821);
and U38737 (N_38737,N_33031,N_34667);
xor U38738 (N_38738,N_32608,N_30854);
and U38739 (N_38739,N_31399,N_34346);
and U38740 (N_38740,N_30224,N_30528);
nand U38741 (N_38741,N_34573,N_34292);
nand U38742 (N_38742,N_33649,N_32824);
xor U38743 (N_38743,N_32539,N_31273);
xor U38744 (N_38744,N_32349,N_31309);
xor U38745 (N_38745,N_31768,N_31916);
nand U38746 (N_38746,N_30768,N_34577);
or U38747 (N_38747,N_34526,N_33684);
xnor U38748 (N_38748,N_31196,N_31861);
nor U38749 (N_38749,N_33640,N_33424);
and U38750 (N_38750,N_30361,N_33772);
nand U38751 (N_38751,N_30918,N_32096);
xnor U38752 (N_38752,N_33050,N_32971);
and U38753 (N_38753,N_34716,N_32687);
or U38754 (N_38754,N_31587,N_34510);
nor U38755 (N_38755,N_34519,N_32035);
nand U38756 (N_38756,N_31177,N_32713);
and U38757 (N_38757,N_34804,N_32185);
nor U38758 (N_38758,N_34260,N_32447);
xnor U38759 (N_38759,N_31429,N_33827);
or U38760 (N_38760,N_31777,N_32724);
nand U38761 (N_38761,N_33088,N_31750);
xnor U38762 (N_38762,N_31525,N_31331);
xor U38763 (N_38763,N_31170,N_33345);
nand U38764 (N_38764,N_34809,N_31628);
nand U38765 (N_38765,N_32405,N_34007);
nand U38766 (N_38766,N_33757,N_31233);
or U38767 (N_38767,N_34801,N_34410);
nor U38768 (N_38768,N_34767,N_30914);
or U38769 (N_38769,N_34401,N_33881);
nand U38770 (N_38770,N_33628,N_33752);
nor U38771 (N_38771,N_34718,N_34120);
and U38772 (N_38772,N_32049,N_31002);
and U38773 (N_38773,N_30861,N_30628);
nand U38774 (N_38774,N_31987,N_33885);
nor U38775 (N_38775,N_32665,N_31090);
nand U38776 (N_38776,N_33524,N_30335);
nand U38777 (N_38777,N_34867,N_30646);
or U38778 (N_38778,N_32339,N_32449);
nand U38779 (N_38779,N_34116,N_30417);
xnor U38780 (N_38780,N_31707,N_30923);
and U38781 (N_38781,N_33023,N_33361);
and U38782 (N_38782,N_30364,N_33975);
nor U38783 (N_38783,N_32990,N_30331);
xor U38784 (N_38784,N_33467,N_34397);
nand U38785 (N_38785,N_31683,N_33357);
nor U38786 (N_38786,N_30458,N_32026);
and U38787 (N_38787,N_34438,N_30878);
nor U38788 (N_38788,N_31910,N_34799);
nor U38789 (N_38789,N_32214,N_34256);
nand U38790 (N_38790,N_33089,N_34576);
nand U38791 (N_38791,N_30932,N_31589);
nand U38792 (N_38792,N_33409,N_32532);
xor U38793 (N_38793,N_33141,N_32590);
nor U38794 (N_38794,N_33733,N_30644);
nor U38795 (N_38795,N_31278,N_31460);
nand U38796 (N_38796,N_30845,N_34063);
or U38797 (N_38797,N_34683,N_34828);
nand U38798 (N_38798,N_33286,N_33488);
nand U38799 (N_38799,N_34503,N_30088);
nor U38800 (N_38800,N_30303,N_32244);
nor U38801 (N_38801,N_31716,N_34020);
xnor U38802 (N_38802,N_32076,N_33538);
nor U38803 (N_38803,N_30027,N_34855);
nand U38804 (N_38804,N_33954,N_30004);
and U38805 (N_38805,N_32887,N_34681);
or U38806 (N_38806,N_33027,N_31788);
nand U38807 (N_38807,N_31440,N_32401);
nor U38808 (N_38808,N_33199,N_30635);
xor U38809 (N_38809,N_30397,N_30969);
or U38810 (N_38810,N_34773,N_31323);
xor U38811 (N_38811,N_34583,N_34543);
nor U38812 (N_38812,N_31275,N_31187);
or U38813 (N_38813,N_34913,N_30068);
and U38814 (N_38814,N_33014,N_30866);
xnor U38815 (N_38815,N_33048,N_32547);
xor U38816 (N_38816,N_31523,N_34005);
xnor U38817 (N_38817,N_32649,N_31586);
nor U38818 (N_38818,N_30807,N_32547);
xnor U38819 (N_38819,N_34237,N_31168);
nand U38820 (N_38820,N_31585,N_32779);
nand U38821 (N_38821,N_30988,N_30520);
and U38822 (N_38822,N_31890,N_30786);
nand U38823 (N_38823,N_33873,N_31686);
nand U38824 (N_38824,N_33929,N_34486);
nand U38825 (N_38825,N_31075,N_31519);
or U38826 (N_38826,N_34288,N_31758);
nor U38827 (N_38827,N_32130,N_34326);
or U38828 (N_38828,N_34922,N_34352);
and U38829 (N_38829,N_30382,N_32990);
or U38830 (N_38830,N_34836,N_31782);
or U38831 (N_38831,N_31501,N_34474);
xnor U38832 (N_38832,N_31802,N_33375);
nand U38833 (N_38833,N_33464,N_34729);
nor U38834 (N_38834,N_30650,N_33296);
xnor U38835 (N_38835,N_34191,N_34254);
xnor U38836 (N_38836,N_32040,N_32693);
or U38837 (N_38837,N_30753,N_31760);
xnor U38838 (N_38838,N_30701,N_32119);
and U38839 (N_38839,N_30172,N_32908);
or U38840 (N_38840,N_33436,N_30375);
or U38841 (N_38841,N_30030,N_33613);
or U38842 (N_38842,N_34310,N_31443);
nand U38843 (N_38843,N_32158,N_34426);
nor U38844 (N_38844,N_32766,N_31356);
xor U38845 (N_38845,N_31064,N_31083);
and U38846 (N_38846,N_30442,N_31738);
xnor U38847 (N_38847,N_32302,N_33817);
and U38848 (N_38848,N_33643,N_31880);
or U38849 (N_38849,N_33847,N_32126);
and U38850 (N_38850,N_33740,N_33096);
or U38851 (N_38851,N_31791,N_32650);
nand U38852 (N_38852,N_31534,N_34239);
nand U38853 (N_38853,N_30974,N_32228);
xor U38854 (N_38854,N_32002,N_32103);
nand U38855 (N_38855,N_32440,N_33387);
and U38856 (N_38856,N_30354,N_31559);
nor U38857 (N_38857,N_30257,N_31577);
xnor U38858 (N_38858,N_31753,N_31148);
xnor U38859 (N_38859,N_30053,N_32978);
xnor U38860 (N_38860,N_31400,N_32935);
xnor U38861 (N_38861,N_33646,N_32284);
or U38862 (N_38862,N_30323,N_33128);
nand U38863 (N_38863,N_32335,N_30011);
nor U38864 (N_38864,N_34291,N_30645);
and U38865 (N_38865,N_32278,N_32189);
nor U38866 (N_38866,N_31677,N_31711);
or U38867 (N_38867,N_34760,N_31189);
nor U38868 (N_38868,N_33530,N_33905);
and U38869 (N_38869,N_32176,N_33066);
xor U38870 (N_38870,N_34753,N_33874);
xor U38871 (N_38871,N_33244,N_34022);
nor U38872 (N_38872,N_32597,N_33160);
nand U38873 (N_38873,N_34262,N_34432);
nor U38874 (N_38874,N_31084,N_32437);
xor U38875 (N_38875,N_34340,N_31184);
xnor U38876 (N_38876,N_34105,N_31395);
nand U38877 (N_38877,N_32682,N_33201);
nor U38878 (N_38878,N_34906,N_30792);
or U38879 (N_38879,N_34474,N_30161);
nor U38880 (N_38880,N_34859,N_32514);
or U38881 (N_38881,N_32127,N_31383);
and U38882 (N_38882,N_31512,N_33577);
and U38883 (N_38883,N_33266,N_32397);
xor U38884 (N_38884,N_33562,N_33089);
xor U38885 (N_38885,N_31874,N_34863);
xor U38886 (N_38886,N_30308,N_34308);
nand U38887 (N_38887,N_31717,N_30268);
or U38888 (N_38888,N_33594,N_31076);
and U38889 (N_38889,N_32430,N_33782);
nor U38890 (N_38890,N_31272,N_31923);
or U38891 (N_38891,N_30894,N_34654);
xnor U38892 (N_38892,N_32650,N_33624);
xor U38893 (N_38893,N_34240,N_30865);
and U38894 (N_38894,N_31944,N_30334);
xor U38895 (N_38895,N_31848,N_33494);
or U38896 (N_38896,N_34544,N_30468);
nor U38897 (N_38897,N_32358,N_31219);
nor U38898 (N_38898,N_32714,N_34267);
xnor U38899 (N_38899,N_34831,N_30644);
xor U38900 (N_38900,N_32973,N_31867);
and U38901 (N_38901,N_31002,N_30796);
or U38902 (N_38902,N_32679,N_31891);
nand U38903 (N_38903,N_31926,N_32512);
or U38904 (N_38904,N_32132,N_31050);
nand U38905 (N_38905,N_31923,N_30306);
nand U38906 (N_38906,N_32719,N_33339);
or U38907 (N_38907,N_32361,N_34435);
nor U38908 (N_38908,N_32882,N_34499);
and U38909 (N_38909,N_31537,N_34728);
nand U38910 (N_38910,N_32752,N_32222);
and U38911 (N_38911,N_32884,N_33271);
nand U38912 (N_38912,N_30634,N_31966);
or U38913 (N_38913,N_32360,N_32075);
nand U38914 (N_38914,N_33443,N_30703);
xor U38915 (N_38915,N_31420,N_34855);
and U38916 (N_38916,N_32495,N_33955);
and U38917 (N_38917,N_31575,N_32673);
and U38918 (N_38918,N_31688,N_33507);
xnor U38919 (N_38919,N_31316,N_31825);
nor U38920 (N_38920,N_31154,N_32909);
nand U38921 (N_38921,N_30771,N_30812);
and U38922 (N_38922,N_31624,N_32041);
nand U38923 (N_38923,N_31504,N_33065);
or U38924 (N_38924,N_32714,N_32911);
nand U38925 (N_38925,N_30807,N_31183);
or U38926 (N_38926,N_34172,N_34362);
nand U38927 (N_38927,N_33124,N_30050);
nor U38928 (N_38928,N_34135,N_32109);
and U38929 (N_38929,N_32747,N_34131);
xnor U38930 (N_38930,N_33602,N_30421);
xor U38931 (N_38931,N_31195,N_30200);
xor U38932 (N_38932,N_32892,N_32181);
nor U38933 (N_38933,N_33320,N_31667);
or U38934 (N_38934,N_30174,N_34366);
xor U38935 (N_38935,N_32174,N_33547);
nor U38936 (N_38936,N_30099,N_34635);
nor U38937 (N_38937,N_32876,N_33567);
nor U38938 (N_38938,N_31030,N_30027);
xnor U38939 (N_38939,N_33846,N_31966);
nand U38940 (N_38940,N_34183,N_34398);
nor U38941 (N_38941,N_34144,N_33049);
nor U38942 (N_38942,N_31720,N_31729);
or U38943 (N_38943,N_34641,N_31641);
or U38944 (N_38944,N_31500,N_31789);
and U38945 (N_38945,N_32952,N_34961);
nor U38946 (N_38946,N_31823,N_34530);
or U38947 (N_38947,N_34125,N_33643);
xnor U38948 (N_38948,N_34070,N_33314);
nand U38949 (N_38949,N_32123,N_30701);
nand U38950 (N_38950,N_30959,N_34851);
xnor U38951 (N_38951,N_34813,N_31149);
nand U38952 (N_38952,N_34136,N_30770);
nor U38953 (N_38953,N_34486,N_33410);
and U38954 (N_38954,N_30699,N_32621);
or U38955 (N_38955,N_30924,N_34832);
nor U38956 (N_38956,N_34808,N_34965);
nand U38957 (N_38957,N_33462,N_31953);
xor U38958 (N_38958,N_33963,N_33043);
xor U38959 (N_38959,N_30118,N_32478);
and U38960 (N_38960,N_32448,N_33291);
and U38961 (N_38961,N_31157,N_31281);
nand U38962 (N_38962,N_32981,N_31650);
nand U38963 (N_38963,N_33411,N_31789);
xor U38964 (N_38964,N_30074,N_34635);
xor U38965 (N_38965,N_33193,N_32980);
or U38966 (N_38966,N_31557,N_30006);
nand U38967 (N_38967,N_32377,N_33211);
or U38968 (N_38968,N_31715,N_32182);
xnor U38969 (N_38969,N_33982,N_34423);
and U38970 (N_38970,N_33461,N_31548);
nor U38971 (N_38971,N_31336,N_33678);
or U38972 (N_38972,N_34466,N_31916);
nand U38973 (N_38973,N_32351,N_33332);
nor U38974 (N_38974,N_30492,N_32711);
nand U38975 (N_38975,N_33046,N_32273);
nand U38976 (N_38976,N_30806,N_32290);
and U38977 (N_38977,N_34181,N_30484);
nand U38978 (N_38978,N_31115,N_30604);
nand U38979 (N_38979,N_34250,N_30593);
nor U38980 (N_38980,N_32532,N_34650);
and U38981 (N_38981,N_31664,N_34843);
xnor U38982 (N_38982,N_33675,N_31739);
xor U38983 (N_38983,N_31731,N_34872);
nor U38984 (N_38984,N_30135,N_30095);
nand U38985 (N_38985,N_31639,N_34831);
and U38986 (N_38986,N_34153,N_33664);
or U38987 (N_38987,N_30573,N_30705);
or U38988 (N_38988,N_33840,N_33952);
and U38989 (N_38989,N_30725,N_33245);
xnor U38990 (N_38990,N_33300,N_30844);
or U38991 (N_38991,N_34267,N_31023);
nand U38992 (N_38992,N_30415,N_32554);
nor U38993 (N_38993,N_32149,N_34063);
xnor U38994 (N_38994,N_34173,N_31034);
xor U38995 (N_38995,N_32344,N_33070);
nand U38996 (N_38996,N_31553,N_33243);
and U38997 (N_38997,N_32637,N_34532);
nor U38998 (N_38998,N_34518,N_30189);
and U38999 (N_38999,N_33679,N_31073);
nand U39000 (N_39000,N_32247,N_33406);
nand U39001 (N_39001,N_33060,N_34372);
xnor U39002 (N_39002,N_33230,N_30734);
and U39003 (N_39003,N_31061,N_34144);
xnor U39004 (N_39004,N_32740,N_32866);
nor U39005 (N_39005,N_34151,N_32093);
or U39006 (N_39006,N_30699,N_31495);
and U39007 (N_39007,N_33248,N_34488);
and U39008 (N_39008,N_33055,N_30243);
and U39009 (N_39009,N_33604,N_31606);
nor U39010 (N_39010,N_30076,N_31309);
nor U39011 (N_39011,N_31340,N_32894);
nand U39012 (N_39012,N_32487,N_32203);
nand U39013 (N_39013,N_31461,N_30732);
and U39014 (N_39014,N_32303,N_33978);
and U39015 (N_39015,N_30718,N_32008);
and U39016 (N_39016,N_32727,N_30278);
and U39017 (N_39017,N_30050,N_31228);
nand U39018 (N_39018,N_32422,N_31227);
nand U39019 (N_39019,N_33399,N_30010);
and U39020 (N_39020,N_30368,N_33547);
xor U39021 (N_39021,N_30570,N_32869);
nand U39022 (N_39022,N_32087,N_32345);
nand U39023 (N_39023,N_32802,N_31544);
xor U39024 (N_39024,N_31581,N_33598);
nand U39025 (N_39025,N_31358,N_30203);
or U39026 (N_39026,N_30634,N_32598);
nor U39027 (N_39027,N_32287,N_34219);
and U39028 (N_39028,N_30532,N_31521);
nor U39029 (N_39029,N_30611,N_32173);
xnor U39030 (N_39030,N_34675,N_31655);
nand U39031 (N_39031,N_33357,N_34237);
or U39032 (N_39032,N_30441,N_33925);
or U39033 (N_39033,N_33393,N_31372);
nor U39034 (N_39034,N_32338,N_31928);
nand U39035 (N_39035,N_32948,N_31904);
nor U39036 (N_39036,N_31176,N_30236);
or U39037 (N_39037,N_30073,N_32773);
nand U39038 (N_39038,N_33645,N_32671);
or U39039 (N_39039,N_30574,N_33255);
and U39040 (N_39040,N_34328,N_33762);
nand U39041 (N_39041,N_33466,N_33914);
nand U39042 (N_39042,N_34738,N_32851);
xnor U39043 (N_39043,N_34613,N_31221);
nand U39044 (N_39044,N_34960,N_34414);
and U39045 (N_39045,N_31087,N_32871);
or U39046 (N_39046,N_30553,N_33790);
xor U39047 (N_39047,N_30728,N_31635);
and U39048 (N_39048,N_33358,N_34572);
nor U39049 (N_39049,N_30880,N_32311);
nand U39050 (N_39050,N_33015,N_32059);
and U39051 (N_39051,N_33193,N_33519);
and U39052 (N_39052,N_33804,N_32755);
xnor U39053 (N_39053,N_32020,N_34017);
nor U39054 (N_39054,N_30106,N_32773);
xnor U39055 (N_39055,N_34590,N_30694);
nand U39056 (N_39056,N_34363,N_31363);
nand U39057 (N_39057,N_31030,N_32416);
or U39058 (N_39058,N_31726,N_31375);
nand U39059 (N_39059,N_33574,N_34218);
and U39060 (N_39060,N_34084,N_31292);
and U39061 (N_39061,N_30821,N_31920);
nand U39062 (N_39062,N_32853,N_32767);
nand U39063 (N_39063,N_30564,N_30776);
xor U39064 (N_39064,N_31959,N_32168);
or U39065 (N_39065,N_31562,N_34700);
or U39066 (N_39066,N_31985,N_32912);
nand U39067 (N_39067,N_30857,N_33040);
nand U39068 (N_39068,N_31617,N_31445);
or U39069 (N_39069,N_30368,N_34868);
and U39070 (N_39070,N_31634,N_30803);
xnor U39071 (N_39071,N_32934,N_34553);
nand U39072 (N_39072,N_33217,N_34106);
or U39073 (N_39073,N_30225,N_33690);
and U39074 (N_39074,N_32791,N_33027);
and U39075 (N_39075,N_31891,N_33295);
and U39076 (N_39076,N_32699,N_32031);
xor U39077 (N_39077,N_32759,N_30802);
xor U39078 (N_39078,N_32756,N_33155);
or U39079 (N_39079,N_33685,N_33188);
or U39080 (N_39080,N_34080,N_31366);
nand U39081 (N_39081,N_30253,N_33380);
xor U39082 (N_39082,N_33200,N_34286);
nand U39083 (N_39083,N_30404,N_32884);
xor U39084 (N_39084,N_31125,N_34467);
and U39085 (N_39085,N_31886,N_31469);
or U39086 (N_39086,N_31555,N_30588);
nor U39087 (N_39087,N_34610,N_31317);
and U39088 (N_39088,N_33607,N_34934);
or U39089 (N_39089,N_32490,N_31252);
xnor U39090 (N_39090,N_30641,N_33323);
or U39091 (N_39091,N_31073,N_32290);
xnor U39092 (N_39092,N_30107,N_34799);
nand U39093 (N_39093,N_30215,N_33222);
nand U39094 (N_39094,N_31643,N_30173);
nor U39095 (N_39095,N_31099,N_30450);
nand U39096 (N_39096,N_30579,N_33062);
and U39097 (N_39097,N_33554,N_34760);
nand U39098 (N_39098,N_34683,N_34414);
nor U39099 (N_39099,N_34901,N_32926);
nor U39100 (N_39100,N_30305,N_34791);
nand U39101 (N_39101,N_34370,N_32490);
nor U39102 (N_39102,N_34774,N_33277);
nand U39103 (N_39103,N_32097,N_34899);
nor U39104 (N_39104,N_30885,N_34629);
nor U39105 (N_39105,N_31226,N_30817);
nand U39106 (N_39106,N_32938,N_32783);
nand U39107 (N_39107,N_31808,N_31140);
and U39108 (N_39108,N_31342,N_30742);
xnor U39109 (N_39109,N_32107,N_31171);
and U39110 (N_39110,N_33272,N_34221);
or U39111 (N_39111,N_30079,N_33133);
or U39112 (N_39112,N_34309,N_33017);
nor U39113 (N_39113,N_33773,N_32714);
and U39114 (N_39114,N_32285,N_33910);
and U39115 (N_39115,N_32408,N_30430);
or U39116 (N_39116,N_31645,N_34530);
nand U39117 (N_39117,N_32758,N_31323);
nor U39118 (N_39118,N_34692,N_31003);
or U39119 (N_39119,N_34132,N_32575);
xor U39120 (N_39120,N_32071,N_34844);
xnor U39121 (N_39121,N_30600,N_30734);
or U39122 (N_39122,N_34389,N_30396);
nor U39123 (N_39123,N_31237,N_32647);
xnor U39124 (N_39124,N_30715,N_30764);
or U39125 (N_39125,N_32828,N_30233);
xor U39126 (N_39126,N_33618,N_31116);
xnor U39127 (N_39127,N_30312,N_31038);
nand U39128 (N_39128,N_30871,N_33171);
nor U39129 (N_39129,N_31827,N_33763);
and U39130 (N_39130,N_34262,N_32021);
or U39131 (N_39131,N_34406,N_34863);
and U39132 (N_39132,N_33408,N_30339);
nor U39133 (N_39133,N_34480,N_34081);
xnor U39134 (N_39134,N_30904,N_31380);
nor U39135 (N_39135,N_31439,N_33310);
nor U39136 (N_39136,N_30857,N_32857);
nor U39137 (N_39137,N_32241,N_34413);
and U39138 (N_39138,N_30270,N_30539);
xor U39139 (N_39139,N_30682,N_33949);
or U39140 (N_39140,N_31862,N_30715);
nor U39141 (N_39141,N_34515,N_33569);
and U39142 (N_39142,N_30439,N_33601);
xor U39143 (N_39143,N_32167,N_34029);
xor U39144 (N_39144,N_34976,N_34640);
nor U39145 (N_39145,N_30458,N_33137);
nand U39146 (N_39146,N_33885,N_32253);
or U39147 (N_39147,N_33004,N_30260);
or U39148 (N_39148,N_32164,N_34450);
nand U39149 (N_39149,N_34694,N_34980);
and U39150 (N_39150,N_30445,N_30072);
and U39151 (N_39151,N_34518,N_34859);
nand U39152 (N_39152,N_32368,N_30225);
nand U39153 (N_39153,N_34914,N_32905);
nand U39154 (N_39154,N_31801,N_33640);
nand U39155 (N_39155,N_32421,N_33484);
xor U39156 (N_39156,N_31959,N_30732);
nand U39157 (N_39157,N_31663,N_32789);
nand U39158 (N_39158,N_32893,N_30549);
nand U39159 (N_39159,N_33564,N_30168);
nor U39160 (N_39160,N_33205,N_31323);
and U39161 (N_39161,N_34714,N_30129);
xor U39162 (N_39162,N_34458,N_33884);
and U39163 (N_39163,N_31668,N_30288);
nor U39164 (N_39164,N_32377,N_30242);
nand U39165 (N_39165,N_32639,N_33576);
nor U39166 (N_39166,N_30698,N_33119);
xor U39167 (N_39167,N_31627,N_31074);
nand U39168 (N_39168,N_33880,N_31521);
xnor U39169 (N_39169,N_31673,N_34620);
or U39170 (N_39170,N_31951,N_33628);
or U39171 (N_39171,N_34778,N_31645);
nor U39172 (N_39172,N_34856,N_34838);
or U39173 (N_39173,N_30558,N_34014);
and U39174 (N_39174,N_34151,N_34823);
xor U39175 (N_39175,N_31190,N_32155);
nand U39176 (N_39176,N_34075,N_31574);
xor U39177 (N_39177,N_32680,N_31682);
or U39178 (N_39178,N_32106,N_31029);
nor U39179 (N_39179,N_34120,N_30498);
or U39180 (N_39180,N_33703,N_33476);
and U39181 (N_39181,N_34244,N_34438);
xor U39182 (N_39182,N_30801,N_31295);
nand U39183 (N_39183,N_33719,N_33587);
and U39184 (N_39184,N_30352,N_32551);
nor U39185 (N_39185,N_34073,N_33675);
xor U39186 (N_39186,N_33910,N_31782);
or U39187 (N_39187,N_34391,N_30483);
nor U39188 (N_39188,N_31994,N_32518);
xor U39189 (N_39189,N_31898,N_30428);
or U39190 (N_39190,N_30782,N_30088);
xor U39191 (N_39191,N_32285,N_34592);
nand U39192 (N_39192,N_31390,N_33182);
nand U39193 (N_39193,N_30035,N_30144);
nand U39194 (N_39194,N_30536,N_33275);
xor U39195 (N_39195,N_33662,N_31751);
xnor U39196 (N_39196,N_34116,N_30306);
nor U39197 (N_39197,N_33233,N_33424);
nand U39198 (N_39198,N_31059,N_32098);
and U39199 (N_39199,N_32993,N_34251);
nor U39200 (N_39200,N_30679,N_34047);
and U39201 (N_39201,N_33591,N_30132);
or U39202 (N_39202,N_30597,N_32876);
or U39203 (N_39203,N_31405,N_34009);
or U39204 (N_39204,N_33375,N_32321);
nand U39205 (N_39205,N_34323,N_30376);
nor U39206 (N_39206,N_30471,N_34494);
xor U39207 (N_39207,N_31964,N_30458);
nand U39208 (N_39208,N_34932,N_30931);
nand U39209 (N_39209,N_34044,N_31715);
nor U39210 (N_39210,N_32208,N_33939);
xnor U39211 (N_39211,N_32426,N_31765);
xnor U39212 (N_39212,N_31626,N_32732);
nand U39213 (N_39213,N_30779,N_33208);
xor U39214 (N_39214,N_32312,N_33544);
nand U39215 (N_39215,N_30892,N_34277);
nand U39216 (N_39216,N_34775,N_31518);
nor U39217 (N_39217,N_34911,N_33994);
and U39218 (N_39218,N_32249,N_34406);
nor U39219 (N_39219,N_31793,N_33842);
or U39220 (N_39220,N_34576,N_34274);
or U39221 (N_39221,N_34487,N_33021);
xor U39222 (N_39222,N_31177,N_30237);
and U39223 (N_39223,N_33468,N_33051);
xor U39224 (N_39224,N_34953,N_30100);
or U39225 (N_39225,N_34423,N_33791);
nand U39226 (N_39226,N_34057,N_31586);
and U39227 (N_39227,N_32603,N_32107);
xor U39228 (N_39228,N_32060,N_32677);
nand U39229 (N_39229,N_30272,N_34083);
nand U39230 (N_39230,N_31144,N_33275);
xnor U39231 (N_39231,N_31032,N_30825);
or U39232 (N_39232,N_34008,N_31968);
nand U39233 (N_39233,N_31490,N_34418);
nor U39234 (N_39234,N_30625,N_31369);
nand U39235 (N_39235,N_34840,N_31180);
nor U39236 (N_39236,N_31855,N_34481);
nand U39237 (N_39237,N_30471,N_31750);
or U39238 (N_39238,N_33968,N_34832);
nand U39239 (N_39239,N_32859,N_31906);
or U39240 (N_39240,N_31898,N_32404);
nand U39241 (N_39241,N_34142,N_34638);
xor U39242 (N_39242,N_32121,N_33378);
and U39243 (N_39243,N_33550,N_34788);
or U39244 (N_39244,N_31619,N_33677);
nor U39245 (N_39245,N_30687,N_33717);
or U39246 (N_39246,N_31396,N_33055);
or U39247 (N_39247,N_33395,N_33446);
nor U39248 (N_39248,N_30504,N_32219);
xnor U39249 (N_39249,N_32190,N_34364);
or U39250 (N_39250,N_32189,N_33506);
nand U39251 (N_39251,N_31849,N_30485);
or U39252 (N_39252,N_31331,N_33133);
and U39253 (N_39253,N_31141,N_34844);
nor U39254 (N_39254,N_32964,N_31055);
and U39255 (N_39255,N_33378,N_31652);
or U39256 (N_39256,N_32867,N_31687);
and U39257 (N_39257,N_32050,N_33288);
or U39258 (N_39258,N_32664,N_30913);
nor U39259 (N_39259,N_34843,N_31999);
or U39260 (N_39260,N_30843,N_30389);
and U39261 (N_39261,N_30333,N_33084);
xnor U39262 (N_39262,N_32603,N_32383);
nor U39263 (N_39263,N_33571,N_30804);
or U39264 (N_39264,N_30812,N_32935);
and U39265 (N_39265,N_31467,N_31683);
nor U39266 (N_39266,N_32958,N_34193);
nand U39267 (N_39267,N_32602,N_31586);
and U39268 (N_39268,N_32530,N_32043);
and U39269 (N_39269,N_31348,N_32865);
or U39270 (N_39270,N_33709,N_30565);
or U39271 (N_39271,N_33049,N_30958);
nand U39272 (N_39272,N_32876,N_31213);
xor U39273 (N_39273,N_31157,N_30468);
or U39274 (N_39274,N_34281,N_33847);
nand U39275 (N_39275,N_34728,N_30706);
nor U39276 (N_39276,N_34947,N_31357);
nand U39277 (N_39277,N_32863,N_31611);
nand U39278 (N_39278,N_32976,N_31110);
nor U39279 (N_39279,N_30337,N_33409);
xnor U39280 (N_39280,N_34289,N_33333);
or U39281 (N_39281,N_33309,N_33186);
and U39282 (N_39282,N_34018,N_32051);
and U39283 (N_39283,N_34764,N_32550);
or U39284 (N_39284,N_31902,N_34052);
nand U39285 (N_39285,N_30325,N_32366);
or U39286 (N_39286,N_30896,N_31084);
nand U39287 (N_39287,N_34252,N_31036);
and U39288 (N_39288,N_30227,N_32613);
nand U39289 (N_39289,N_30389,N_30860);
nand U39290 (N_39290,N_32348,N_34945);
nand U39291 (N_39291,N_34234,N_31519);
and U39292 (N_39292,N_32362,N_33263);
and U39293 (N_39293,N_34330,N_33144);
and U39294 (N_39294,N_34237,N_30901);
xnor U39295 (N_39295,N_30987,N_34193);
nand U39296 (N_39296,N_32536,N_33251);
nor U39297 (N_39297,N_31703,N_30325);
or U39298 (N_39298,N_33665,N_31302);
xor U39299 (N_39299,N_32667,N_34606);
nor U39300 (N_39300,N_32008,N_32433);
nor U39301 (N_39301,N_34117,N_31542);
nor U39302 (N_39302,N_34298,N_30564);
and U39303 (N_39303,N_30160,N_33442);
or U39304 (N_39304,N_34124,N_33817);
xor U39305 (N_39305,N_30359,N_34621);
nor U39306 (N_39306,N_30687,N_30747);
and U39307 (N_39307,N_34565,N_30059);
nor U39308 (N_39308,N_32817,N_32597);
or U39309 (N_39309,N_34764,N_33216);
nand U39310 (N_39310,N_32095,N_33992);
xor U39311 (N_39311,N_31344,N_31418);
and U39312 (N_39312,N_32113,N_31937);
xnor U39313 (N_39313,N_30243,N_31765);
nor U39314 (N_39314,N_31822,N_30073);
xnor U39315 (N_39315,N_31956,N_32871);
and U39316 (N_39316,N_33048,N_31553);
nor U39317 (N_39317,N_33956,N_30813);
xor U39318 (N_39318,N_31170,N_32591);
nand U39319 (N_39319,N_31184,N_31063);
nand U39320 (N_39320,N_34831,N_30090);
xor U39321 (N_39321,N_31378,N_33018);
nor U39322 (N_39322,N_31830,N_31517);
nor U39323 (N_39323,N_33606,N_31832);
nand U39324 (N_39324,N_31849,N_31781);
and U39325 (N_39325,N_32314,N_32177);
or U39326 (N_39326,N_30896,N_31405);
nand U39327 (N_39327,N_31477,N_30230);
nand U39328 (N_39328,N_32792,N_34563);
nand U39329 (N_39329,N_31048,N_33754);
nand U39330 (N_39330,N_32406,N_32590);
xor U39331 (N_39331,N_34654,N_32350);
nand U39332 (N_39332,N_34579,N_33321);
and U39333 (N_39333,N_33426,N_30309);
and U39334 (N_39334,N_33432,N_33606);
xor U39335 (N_39335,N_31908,N_34250);
and U39336 (N_39336,N_31701,N_30830);
or U39337 (N_39337,N_34003,N_31703);
xnor U39338 (N_39338,N_31180,N_31748);
or U39339 (N_39339,N_32118,N_31102);
nor U39340 (N_39340,N_33468,N_33728);
xor U39341 (N_39341,N_30401,N_30935);
xnor U39342 (N_39342,N_30125,N_34673);
or U39343 (N_39343,N_32497,N_30106);
nor U39344 (N_39344,N_30658,N_32085);
and U39345 (N_39345,N_33549,N_34332);
xor U39346 (N_39346,N_34181,N_31304);
nand U39347 (N_39347,N_32093,N_30697);
or U39348 (N_39348,N_32578,N_30645);
nand U39349 (N_39349,N_31059,N_34728);
or U39350 (N_39350,N_31695,N_34416);
or U39351 (N_39351,N_33117,N_31689);
xnor U39352 (N_39352,N_34031,N_34051);
nand U39353 (N_39353,N_32545,N_30826);
xnor U39354 (N_39354,N_34884,N_33114);
xor U39355 (N_39355,N_32219,N_33802);
or U39356 (N_39356,N_31014,N_33591);
or U39357 (N_39357,N_31934,N_30772);
nand U39358 (N_39358,N_34251,N_31488);
xor U39359 (N_39359,N_30202,N_30707);
and U39360 (N_39360,N_33477,N_31276);
nand U39361 (N_39361,N_32719,N_32737);
nor U39362 (N_39362,N_34539,N_34715);
nor U39363 (N_39363,N_32412,N_32166);
and U39364 (N_39364,N_34858,N_34789);
nand U39365 (N_39365,N_30545,N_32689);
nand U39366 (N_39366,N_31017,N_32807);
and U39367 (N_39367,N_33118,N_30954);
and U39368 (N_39368,N_30317,N_31615);
nand U39369 (N_39369,N_32081,N_31426);
nand U39370 (N_39370,N_31707,N_33403);
nand U39371 (N_39371,N_30202,N_31567);
xnor U39372 (N_39372,N_32986,N_34461);
nand U39373 (N_39373,N_31418,N_32721);
nand U39374 (N_39374,N_32016,N_34863);
nand U39375 (N_39375,N_30777,N_31943);
xor U39376 (N_39376,N_31955,N_32721);
nor U39377 (N_39377,N_31945,N_34875);
nand U39378 (N_39378,N_34446,N_32132);
nand U39379 (N_39379,N_32650,N_31154);
nand U39380 (N_39380,N_34846,N_30951);
and U39381 (N_39381,N_30860,N_30222);
or U39382 (N_39382,N_33873,N_33895);
nor U39383 (N_39383,N_33469,N_32409);
xnor U39384 (N_39384,N_30452,N_34162);
nor U39385 (N_39385,N_32871,N_34260);
xnor U39386 (N_39386,N_30466,N_30081);
or U39387 (N_39387,N_32987,N_31813);
nand U39388 (N_39388,N_31181,N_31994);
nand U39389 (N_39389,N_31988,N_30493);
and U39390 (N_39390,N_34233,N_34010);
xnor U39391 (N_39391,N_33941,N_30189);
and U39392 (N_39392,N_34809,N_31120);
or U39393 (N_39393,N_33683,N_34606);
and U39394 (N_39394,N_33793,N_33720);
or U39395 (N_39395,N_31169,N_30967);
or U39396 (N_39396,N_34207,N_33452);
xor U39397 (N_39397,N_34125,N_30363);
xor U39398 (N_39398,N_32664,N_30864);
nor U39399 (N_39399,N_30064,N_34172);
xnor U39400 (N_39400,N_31741,N_32201);
or U39401 (N_39401,N_32050,N_31009);
nand U39402 (N_39402,N_31285,N_34369);
nand U39403 (N_39403,N_32336,N_33669);
and U39404 (N_39404,N_32349,N_31688);
nor U39405 (N_39405,N_33243,N_34897);
or U39406 (N_39406,N_31962,N_33122);
nand U39407 (N_39407,N_33273,N_30490);
nor U39408 (N_39408,N_30784,N_34170);
nor U39409 (N_39409,N_34569,N_33234);
nor U39410 (N_39410,N_31360,N_33373);
or U39411 (N_39411,N_32099,N_33684);
or U39412 (N_39412,N_34934,N_31664);
nand U39413 (N_39413,N_30540,N_30408);
or U39414 (N_39414,N_34711,N_33503);
xnor U39415 (N_39415,N_31128,N_30795);
nand U39416 (N_39416,N_30642,N_34103);
or U39417 (N_39417,N_30394,N_32193);
and U39418 (N_39418,N_31266,N_30827);
nand U39419 (N_39419,N_31157,N_34823);
nor U39420 (N_39420,N_31621,N_30443);
and U39421 (N_39421,N_33120,N_34346);
nand U39422 (N_39422,N_30013,N_34428);
or U39423 (N_39423,N_32365,N_31903);
and U39424 (N_39424,N_30716,N_30421);
xnor U39425 (N_39425,N_32622,N_33236);
nand U39426 (N_39426,N_34871,N_34386);
nand U39427 (N_39427,N_33404,N_33541);
nand U39428 (N_39428,N_33730,N_32066);
and U39429 (N_39429,N_34599,N_34384);
xor U39430 (N_39430,N_30287,N_32775);
xor U39431 (N_39431,N_33524,N_32226);
nor U39432 (N_39432,N_32931,N_30778);
nand U39433 (N_39433,N_34623,N_30914);
nand U39434 (N_39434,N_31474,N_31582);
nor U39435 (N_39435,N_32936,N_33473);
or U39436 (N_39436,N_33153,N_30823);
and U39437 (N_39437,N_33845,N_31931);
xor U39438 (N_39438,N_31739,N_30366);
or U39439 (N_39439,N_34220,N_34596);
xor U39440 (N_39440,N_30637,N_30816);
xnor U39441 (N_39441,N_31471,N_33757);
nand U39442 (N_39442,N_31755,N_30507);
or U39443 (N_39443,N_30175,N_32548);
nor U39444 (N_39444,N_33645,N_30431);
nand U39445 (N_39445,N_31203,N_32973);
nor U39446 (N_39446,N_30045,N_30038);
xor U39447 (N_39447,N_33188,N_32561);
xnor U39448 (N_39448,N_34595,N_34013);
nand U39449 (N_39449,N_34407,N_31847);
and U39450 (N_39450,N_33190,N_32650);
and U39451 (N_39451,N_30680,N_33742);
and U39452 (N_39452,N_30054,N_30011);
xnor U39453 (N_39453,N_33221,N_34530);
and U39454 (N_39454,N_32554,N_33919);
xnor U39455 (N_39455,N_32169,N_31254);
xor U39456 (N_39456,N_31089,N_32114);
nand U39457 (N_39457,N_34528,N_31118);
nor U39458 (N_39458,N_34042,N_31184);
or U39459 (N_39459,N_30603,N_33339);
xnor U39460 (N_39460,N_32173,N_32421);
and U39461 (N_39461,N_30960,N_30231);
and U39462 (N_39462,N_31475,N_33588);
and U39463 (N_39463,N_34758,N_30907);
and U39464 (N_39464,N_32693,N_33986);
nor U39465 (N_39465,N_31777,N_30433);
nor U39466 (N_39466,N_31379,N_33483);
xor U39467 (N_39467,N_30709,N_32328);
nand U39468 (N_39468,N_32569,N_30252);
xnor U39469 (N_39469,N_34883,N_34731);
or U39470 (N_39470,N_34912,N_33146);
or U39471 (N_39471,N_34232,N_31042);
nand U39472 (N_39472,N_30007,N_32495);
nor U39473 (N_39473,N_30259,N_30023);
xnor U39474 (N_39474,N_31873,N_31115);
xnor U39475 (N_39475,N_32223,N_30590);
xnor U39476 (N_39476,N_33761,N_33512);
and U39477 (N_39477,N_34545,N_33360);
xor U39478 (N_39478,N_34698,N_31565);
or U39479 (N_39479,N_30916,N_34588);
nand U39480 (N_39480,N_34091,N_32380);
or U39481 (N_39481,N_31453,N_34786);
nand U39482 (N_39482,N_34736,N_31740);
xor U39483 (N_39483,N_32080,N_32919);
xor U39484 (N_39484,N_30625,N_32873);
and U39485 (N_39485,N_34491,N_32446);
nand U39486 (N_39486,N_30946,N_32968);
xnor U39487 (N_39487,N_34020,N_30266);
and U39488 (N_39488,N_34556,N_33518);
nand U39489 (N_39489,N_30405,N_30784);
nand U39490 (N_39490,N_30006,N_32559);
nand U39491 (N_39491,N_30167,N_31708);
nor U39492 (N_39492,N_31860,N_30454);
nor U39493 (N_39493,N_32933,N_34771);
or U39494 (N_39494,N_31451,N_32070);
xor U39495 (N_39495,N_34810,N_31419);
or U39496 (N_39496,N_32436,N_30332);
xnor U39497 (N_39497,N_30466,N_33437);
nor U39498 (N_39498,N_30941,N_34632);
nand U39499 (N_39499,N_33632,N_32421);
or U39500 (N_39500,N_30204,N_32906);
and U39501 (N_39501,N_31052,N_31952);
nor U39502 (N_39502,N_34663,N_32652);
xnor U39503 (N_39503,N_30459,N_31571);
and U39504 (N_39504,N_31347,N_32041);
nor U39505 (N_39505,N_31635,N_34421);
and U39506 (N_39506,N_34163,N_31886);
nand U39507 (N_39507,N_31810,N_30639);
nand U39508 (N_39508,N_31987,N_30543);
xor U39509 (N_39509,N_31034,N_33803);
nor U39510 (N_39510,N_34271,N_33243);
nand U39511 (N_39511,N_34099,N_30311);
nor U39512 (N_39512,N_33585,N_32830);
xor U39513 (N_39513,N_30848,N_30471);
or U39514 (N_39514,N_34680,N_31616);
xnor U39515 (N_39515,N_33805,N_33744);
and U39516 (N_39516,N_31734,N_33779);
nor U39517 (N_39517,N_32204,N_32196);
xor U39518 (N_39518,N_34034,N_32085);
nand U39519 (N_39519,N_30858,N_31954);
or U39520 (N_39520,N_32559,N_33800);
nand U39521 (N_39521,N_34586,N_32393);
and U39522 (N_39522,N_33489,N_31608);
or U39523 (N_39523,N_34791,N_30717);
nor U39524 (N_39524,N_30137,N_34795);
nor U39525 (N_39525,N_30762,N_34217);
nor U39526 (N_39526,N_32300,N_33254);
or U39527 (N_39527,N_34148,N_34390);
nor U39528 (N_39528,N_34071,N_31820);
nor U39529 (N_39529,N_33834,N_30155);
nor U39530 (N_39530,N_30068,N_32693);
or U39531 (N_39531,N_31847,N_33686);
and U39532 (N_39532,N_34613,N_30929);
or U39533 (N_39533,N_33490,N_31837);
or U39534 (N_39534,N_34651,N_34095);
nand U39535 (N_39535,N_30155,N_30085);
xor U39536 (N_39536,N_34051,N_30928);
xor U39537 (N_39537,N_30106,N_34837);
and U39538 (N_39538,N_32417,N_34475);
and U39539 (N_39539,N_31100,N_34427);
and U39540 (N_39540,N_30191,N_31314);
and U39541 (N_39541,N_33108,N_30442);
and U39542 (N_39542,N_32737,N_31135);
or U39543 (N_39543,N_30916,N_31452);
nor U39544 (N_39544,N_31654,N_31676);
and U39545 (N_39545,N_33353,N_33124);
nand U39546 (N_39546,N_31417,N_34317);
nor U39547 (N_39547,N_34388,N_33961);
nand U39548 (N_39548,N_34895,N_30537);
xnor U39549 (N_39549,N_31588,N_30478);
nor U39550 (N_39550,N_33725,N_33351);
or U39551 (N_39551,N_34639,N_31359);
nand U39552 (N_39552,N_34150,N_33282);
xnor U39553 (N_39553,N_32955,N_30257);
xnor U39554 (N_39554,N_32576,N_31971);
nand U39555 (N_39555,N_33953,N_33033);
nand U39556 (N_39556,N_32926,N_34033);
or U39557 (N_39557,N_31656,N_31024);
nor U39558 (N_39558,N_33650,N_32887);
or U39559 (N_39559,N_33292,N_33348);
or U39560 (N_39560,N_34330,N_32485);
or U39561 (N_39561,N_33309,N_31767);
xnor U39562 (N_39562,N_33197,N_30088);
or U39563 (N_39563,N_34524,N_31856);
xnor U39564 (N_39564,N_31549,N_30600);
xor U39565 (N_39565,N_33454,N_32682);
nand U39566 (N_39566,N_32509,N_34896);
or U39567 (N_39567,N_34925,N_32898);
nand U39568 (N_39568,N_31684,N_34708);
nand U39569 (N_39569,N_32326,N_32964);
nor U39570 (N_39570,N_31842,N_31769);
or U39571 (N_39571,N_33752,N_31345);
or U39572 (N_39572,N_34462,N_31022);
and U39573 (N_39573,N_34519,N_34942);
or U39574 (N_39574,N_33481,N_31551);
or U39575 (N_39575,N_33126,N_34521);
nor U39576 (N_39576,N_30023,N_31306);
nand U39577 (N_39577,N_33954,N_31274);
or U39578 (N_39578,N_33388,N_30993);
and U39579 (N_39579,N_33970,N_31011);
nand U39580 (N_39580,N_30720,N_31703);
xor U39581 (N_39581,N_32791,N_31204);
nand U39582 (N_39582,N_33270,N_30915);
xor U39583 (N_39583,N_30809,N_32299);
or U39584 (N_39584,N_31680,N_30276);
nand U39585 (N_39585,N_32583,N_34640);
and U39586 (N_39586,N_33401,N_32440);
xor U39587 (N_39587,N_32024,N_34439);
nand U39588 (N_39588,N_34439,N_32221);
and U39589 (N_39589,N_33523,N_33524);
xor U39590 (N_39590,N_30018,N_32231);
xnor U39591 (N_39591,N_30078,N_31403);
and U39592 (N_39592,N_30375,N_34618);
xor U39593 (N_39593,N_34871,N_32090);
xor U39594 (N_39594,N_30183,N_30149);
or U39595 (N_39595,N_34026,N_32691);
and U39596 (N_39596,N_33446,N_31599);
nor U39597 (N_39597,N_34930,N_33689);
or U39598 (N_39598,N_31997,N_32349);
xnor U39599 (N_39599,N_30202,N_30089);
or U39600 (N_39600,N_32144,N_30801);
and U39601 (N_39601,N_30730,N_34067);
nand U39602 (N_39602,N_33013,N_30895);
nand U39603 (N_39603,N_34740,N_30287);
or U39604 (N_39604,N_33015,N_32865);
or U39605 (N_39605,N_33661,N_33128);
nand U39606 (N_39606,N_30564,N_31898);
nor U39607 (N_39607,N_33657,N_33586);
and U39608 (N_39608,N_32453,N_34412);
xnor U39609 (N_39609,N_31877,N_34576);
or U39610 (N_39610,N_31740,N_33340);
nand U39611 (N_39611,N_33441,N_34156);
nand U39612 (N_39612,N_34335,N_33085);
nor U39613 (N_39613,N_34954,N_30268);
nor U39614 (N_39614,N_30995,N_33457);
or U39615 (N_39615,N_31689,N_30258);
and U39616 (N_39616,N_32807,N_33317);
xnor U39617 (N_39617,N_31506,N_32336);
nor U39618 (N_39618,N_32983,N_32524);
or U39619 (N_39619,N_32782,N_30961);
xor U39620 (N_39620,N_31298,N_31206);
nand U39621 (N_39621,N_31515,N_34866);
nand U39622 (N_39622,N_33529,N_30953);
or U39623 (N_39623,N_34629,N_34265);
or U39624 (N_39624,N_34374,N_34079);
or U39625 (N_39625,N_32934,N_32487);
and U39626 (N_39626,N_32632,N_32030);
xnor U39627 (N_39627,N_32508,N_31768);
nand U39628 (N_39628,N_31912,N_34105);
or U39629 (N_39629,N_34691,N_33346);
nand U39630 (N_39630,N_31498,N_33611);
nor U39631 (N_39631,N_33739,N_30500);
and U39632 (N_39632,N_31400,N_32839);
or U39633 (N_39633,N_34220,N_31596);
nand U39634 (N_39634,N_32850,N_33209);
and U39635 (N_39635,N_30649,N_30366);
or U39636 (N_39636,N_33556,N_34787);
xnor U39637 (N_39637,N_32963,N_31056);
or U39638 (N_39638,N_32915,N_34281);
xnor U39639 (N_39639,N_31929,N_31597);
or U39640 (N_39640,N_32331,N_32618);
or U39641 (N_39641,N_33548,N_34183);
nand U39642 (N_39642,N_31147,N_31687);
xnor U39643 (N_39643,N_32588,N_30690);
nand U39644 (N_39644,N_33109,N_31996);
nor U39645 (N_39645,N_31329,N_32378);
nor U39646 (N_39646,N_33123,N_32575);
or U39647 (N_39647,N_34726,N_34921);
xnor U39648 (N_39648,N_33177,N_31303);
or U39649 (N_39649,N_34288,N_30540);
nor U39650 (N_39650,N_32331,N_31166);
and U39651 (N_39651,N_33049,N_32547);
or U39652 (N_39652,N_31120,N_32137);
nor U39653 (N_39653,N_30641,N_33694);
or U39654 (N_39654,N_30300,N_31627);
nor U39655 (N_39655,N_31004,N_31253);
or U39656 (N_39656,N_31444,N_34116);
xnor U39657 (N_39657,N_33169,N_30465);
or U39658 (N_39658,N_33812,N_32103);
or U39659 (N_39659,N_32264,N_32042);
nor U39660 (N_39660,N_31779,N_32120);
and U39661 (N_39661,N_33068,N_30801);
xor U39662 (N_39662,N_34365,N_31192);
nand U39663 (N_39663,N_30509,N_34398);
nor U39664 (N_39664,N_33142,N_31722);
nor U39665 (N_39665,N_34944,N_30779);
nor U39666 (N_39666,N_33770,N_33010);
or U39667 (N_39667,N_31172,N_31568);
or U39668 (N_39668,N_30870,N_30194);
nor U39669 (N_39669,N_32758,N_34260);
or U39670 (N_39670,N_32599,N_34266);
xor U39671 (N_39671,N_32115,N_34532);
and U39672 (N_39672,N_32856,N_31612);
nand U39673 (N_39673,N_32468,N_32453);
or U39674 (N_39674,N_34307,N_32928);
nand U39675 (N_39675,N_31259,N_30112);
xnor U39676 (N_39676,N_34140,N_30992);
xor U39677 (N_39677,N_34271,N_33559);
and U39678 (N_39678,N_32352,N_33914);
nand U39679 (N_39679,N_33952,N_32578);
and U39680 (N_39680,N_32238,N_30427);
nand U39681 (N_39681,N_32795,N_30179);
and U39682 (N_39682,N_31671,N_30447);
and U39683 (N_39683,N_34515,N_33048);
nand U39684 (N_39684,N_32031,N_34468);
nand U39685 (N_39685,N_32776,N_31828);
xnor U39686 (N_39686,N_30740,N_33898);
and U39687 (N_39687,N_32652,N_34713);
xor U39688 (N_39688,N_34949,N_34857);
nor U39689 (N_39689,N_34228,N_34953);
nor U39690 (N_39690,N_34966,N_33746);
and U39691 (N_39691,N_32977,N_30482);
nor U39692 (N_39692,N_32897,N_30122);
nand U39693 (N_39693,N_32138,N_32643);
nand U39694 (N_39694,N_34125,N_33485);
nor U39695 (N_39695,N_32419,N_33463);
and U39696 (N_39696,N_31645,N_31348);
nor U39697 (N_39697,N_34699,N_32271);
or U39698 (N_39698,N_32056,N_33082);
xnor U39699 (N_39699,N_32467,N_34688);
xor U39700 (N_39700,N_34014,N_31856);
nand U39701 (N_39701,N_34254,N_30386);
xnor U39702 (N_39702,N_30237,N_30056);
or U39703 (N_39703,N_33745,N_32875);
xor U39704 (N_39704,N_31004,N_31121);
or U39705 (N_39705,N_34204,N_32108);
nor U39706 (N_39706,N_32570,N_30023);
xor U39707 (N_39707,N_30335,N_33481);
and U39708 (N_39708,N_33604,N_30353);
or U39709 (N_39709,N_32276,N_33148);
and U39710 (N_39710,N_34359,N_30378);
nor U39711 (N_39711,N_30825,N_31137);
and U39712 (N_39712,N_31235,N_33413);
and U39713 (N_39713,N_32918,N_30682);
nand U39714 (N_39714,N_33052,N_32407);
or U39715 (N_39715,N_34957,N_30866);
or U39716 (N_39716,N_32500,N_33157);
nand U39717 (N_39717,N_32245,N_30385);
xor U39718 (N_39718,N_33856,N_30584);
nor U39719 (N_39719,N_33255,N_31001);
nor U39720 (N_39720,N_30974,N_30418);
or U39721 (N_39721,N_33647,N_34161);
and U39722 (N_39722,N_32587,N_33088);
nand U39723 (N_39723,N_34939,N_30135);
or U39724 (N_39724,N_34826,N_32034);
nor U39725 (N_39725,N_32747,N_34675);
and U39726 (N_39726,N_32265,N_32895);
xnor U39727 (N_39727,N_33260,N_30299);
xor U39728 (N_39728,N_32566,N_31369);
nand U39729 (N_39729,N_33750,N_32345);
nand U39730 (N_39730,N_32746,N_34459);
xnor U39731 (N_39731,N_33470,N_33759);
or U39732 (N_39732,N_31628,N_30035);
and U39733 (N_39733,N_34536,N_34927);
nor U39734 (N_39734,N_33570,N_30503);
and U39735 (N_39735,N_34613,N_33951);
nand U39736 (N_39736,N_31715,N_30976);
xnor U39737 (N_39737,N_33311,N_32223);
nor U39738 (N_39738,N_34411,N_30283);
xor U39739 (N_39739,N_30624,N_32958);
xor U39740 (N_39740,N_30428,N_30691);
xnor U39741 (N_39741,N_31798,N_30338);
nand U39742 (N_39742,N_33067,N_33661);
xor U39743 (N_39743,N_34319,N_31694);
nor U39744 (N_39744,N_33038,N_31526);
nor U39745 (N_39745,N_30390,N_31883);
nor U39746 (N_39746,N_30201,N_31808);
or U39747 (N_39747,N_34158,N_30255);
xnor U39748 (N_39748,N_32632,N_33147);
nor U39749 (N_39749,N_30468,N_31984);
nor U39750 (N_39750,N_33099,N_32550);
nor U39751 (N_39751,N_34195,N_31368);
nand U39752 (N_39752,N_33090,N_33338);
nor U39753 (N_39753,N_32320,N_30990);
nor U39754 (N_39754,N_34566,N_32042);
nand U39755 (N_39755,N_33608,N_32538);
nand U39756 (N_39756,N_32605,N_34738);
or U39757 (N_39757,N_34511,N_31181);
nor U39758 (N_39758,N_32056,N_32836);
or U39759 (N_39759,N_31138,N_32901);
or U39760 (N_39760,N_31286,N_31838);
xnor U39761 (N_39761,N_31246,N_34441);
nor U39762 (N_39762,N_30931,N_30510);
nand U39763 (N_39763,N_34295,N_33096);
and U39764 (N_39764,N_34542,N_33974);
or U39765 (N_39765,N_31494,N_31486);
xor U39766 (N_39766,N_32928,N_31404);
nor U39767 (N_39767,N_34939,N_31497);
or U39768 (N_39768,N_30601,N_34675);
nand U39769 (N_39769,N_32271,N_30931);
nand U39770 (N_39770,N_34672,N_32717);
nor U39771 (N_39771,N_34533,N_34167);
nor U39772 (N_39772,N_34573,N_31684);
nand U39773 (N_39773,N_32307,N_34056);
or U39774 (N_39774,N_30164,N_33329);
and U39775 (N_39775,N_31762,N_31060);
nor U39776 (N_39776,N_31164,N_34437);
and U39777 (N_39777,N_33516,N_34020);
xnor U39778 (N_39778,N_31006,N_34337);
and U39779 (N_39779,N_33548,N_32822);
nand U39780 (N_39780,N_31546,N_33774);
or U39781 (N_39781,N_34754,N_30820);
nand U39782 (N_39782,N_32204,N_34302);
and U39783 (N_39783,N_31754,N_33667);
and U39784 (N_39784,N_30778,N_30022);
nor U39785 (N_39785,N_33644,N_31868);
nand U39786 (N_39786,N_33156,N_31749);
or U39787 (N_39787,N_33866,N_31881);
or U39788 (N_39788,N_31999,N_33479);
or U39789 (N_39789,N_32806,N_33090);
and U39790 (N_39790,N_33392,N_32217);
or U39791 (N_39791,N_32512,N_33502);
nor U39792 (N_39792,N_30132,N_34779);
xor U39793 (N_39793,N_32008,N_32124);
or U39794 (N_39794,N_34896,N_30103);
and U39795 (N_39795,N_34858,N_32410);
nand U39796 (N_39796,N_32522,N_31787);
nand U39797 (N_39797,N_31583,N_33830);
and U39798 (N_39798,N_33007,N_33076);
and U39799 (N_39799,N_33678,N_34767);
and U39800 (N_39800,N_30495,N_30645);
nand U39801 (N_39801,N_34385,N_33647);
nand U39802 (N_39802,N_30494,N_31334);
nor U39803 (N_39803,N_32709,N_30422);
and U39804 (N_39804,N_31171,N_32455);
and U39805 (N_39805,N_30545,N_31685);
or U39806 (N_39806,N_32884,N_32344);
nand U39807 (N_39807,N_33027,N_34535);
and U39808 (N_39808,N_33111,N_33795);
nand U39809 (N_39809,N_34097,N_31059);
or U39810 (N_39810,N_30849,N_31144);
nor U39811 (N_39811,N_30043,N_32166);
and U39812 (N_39812,N_32024,N_32535);
nand U39813 (N_39813,N_32464,N_34916);
xnor U39814 (N_39814,N_33646,N_30929);
nand U39815 (N_39815,N_32229,N_30527);
or U39816 (N_39816,N_31379,N_31241);
or U39817 (N_39817,N_32536,N_32395);
and U39818 (N_39818,N_32564,N_32011);
nor U39819 (N_39819,N_31808,N_33872);
nand U39820 (N_39820,N_30227,N_32894);
or U39821 (N_39821,N_30987,N_31949);
nor U39822 (N_39822,N_30107,N_34125);
xor U39823 (N_39823,N_33847,N_32281);
and U39824 (N_39824,N_34992,N_30520);
nand U39825 (N_39825,N_32169,N_34219);
nor U39826 (N_39826,N_31505,N_34688);
nand U39827 (N_39827,N_32634,N_32019);
nor U39828 (N_39828,N_31319,N_32334);
nor U39829 (N_39829,N_31411,N_33437);
nand U39830 (N_39830,N_32616,N_32828);
and U39831 (N_39831,N_32034,N_32921);
nor U39832 (N_39832,N_33788,N_33142);
xnor U39833 (N_39833,N_33047,N_30401);
nor U39834 (N_39834,N_30750,N_31485);
nand U39835 (N_39835,N_31044,N_30904);
and U39836 (N_39836,N_30824,N_31852);
nand U39837 (N_39837,N_30504,N_30684);
or U39838 (N_39838,N_32227,N_33584);
and U39839 (N_39839,N_32500,N_31795);
or U39840 (N_39840,N_33318,N_34653);
xnor U39841 (N_39841,N_30144,N_32027);
nor U39842 (N_39842,N_33327,N_31083);
nor U39843 (N_39843,N_32410,N_32015);
and U39844 (N_39844,N_34010,N_30447);
nand U39845 (N_39845,N_30413,N_33972);
nand U39846 (N_39846,N_32336,N_30207);
or U39847 (N_39847,N_34036,N_31549);
nand U39848 (N_39848,N_34431,N_33753);
or U39849 (N_39849,N_33001,N_30769);
nand U39850 (N_39850,N_34494,N_33983);
xnor U39851 (N_39851,N_33725,N_34769);
or U39852 (N_39852,N_30675,N_33843);
xnor U39853 (N_39853,N_32978,N_34970);
nand U39854 (N_39854,N_34905,N_31253);
xnor U39855 (N_39855,N_33169,N_34120);
nand U39856 (N_39856,N_34226,N_34506);
nor U39857 (N_39857,N_32207,N_30500);
nor U39858 (N_39858,N_30054,N_30119);
or U39859 (N_39859,N_32373,N_30471);
nand U39860 (N_39860,N_32900,N_33138);
and U39861 (N_39861,N_32234,N_32955);
nor U39862 (N_39862,N_32999,N_32217);
nor U39863 (N_39863,N_31851,N_32441);
or U39864 (N_39864,N_31252,N_31520);
nand U39865 (N_39865,N_30241,N_32480);
or U39866 (N_39866,N_34745,N_32896);
and U39867 (N_39867,N_32005,N_31954);
nand U39868 (N_39868,N_30982,N_32507);
nor U39869 (N_39869,N_31272,N_33221);
nand U39870 (N_39870,N_33803,N_34240);
nor U39871 (N_39871,N_33941,N_31644);
xor U39872 (N_39872,N_33148,N_32704);
xor U39873 (N_39873,N_33789,N_33547);
nand U39874 (N_39874,N_32967,N_32122);
xor U39875 (N_39875,N_30696,N_34830);
xor U39876 (N_39876,N_30554,N_33992);
nor U39877 (N_39877,N_34360,N_33715);
nor U39878 (N_39878,N_34071,N_30327);
or U39879 (N_39879,N_31718,N_31936);
xor U39880 (N_39880,N_32596,N_34574);
nor U39881 (N_39881,N_34184,N_31652);
and U39882 (N_39882,N_31974,N_33626);
or U39883 (N_39883,N_33085,N_31093);
nand U39884 (N_39884,N_32266,N_30913);
and U39885 (N_39885,N_30232,N_32050);
nand U39886 (N_39886,N_30499,N_34145);
or U39887 (N_39887,N_31162,N_34173);
xor U39888 (N_39888,N_30413,N_33496);
or U39889 (N_39889,N_32024,N_32190);
xor U39890 (N_39890,N_32627,N_31318);
xnor U39891 (N_39891,N_34007,N_34120);
or U39892 (N_39892,N_34078,N_34837);
nand U39893 (N_39893,N_33992,N_31834);
nand U39894 (N_39894,N_32294,N_30888);
and U39895 (N_39895,N_33741,N_34658);
nor U39896 (N_39896,N_33350,N_30069);
and U39897 (N_39897,N_33717,N_30027);
nor U39898 (N_39898,N_32926,N_33861);
and U39899 (N_39899,N_32553,N_33718);
or U39900 (N_39900,N_33101,N_34170);
xor U39901 (N_39901,N_31557,N_32900);
and U39902 (N_39902,N_34833,N_32435);
or U39903 (N_39903,N_30637,N_31046);
nor U39904 (N_39904,N_30451,N_34570);
and U39905 (N_39905,N_30261,N_31973);
nand U39906 (N_39906,N_34498,N_32658);
nor U39907 (N_39907,N_30850,N_34026);
nor U39908 (N_39908,N_31494,N_34035);
or U39909 (N_39909,N_31441,N_32553);
or U39910 (N_39910,N_30110,N_34568);
xor U39911 (N_39911,N_33739,N_30305);
and U39912 (N_39912,N_33823,N_32279);
and U39913 (N_39913,N_34206,N_34475);
and U39914 (N_39914,N_32523,N_31969);
xor U39915 (N_39915,N_33803,N_32879);
and U39916 (N_39916,N_32821,N_33126);
xnor U39917 (N_39917,N_33164,N_32251);
nand U39918 (N_39918,N_31945,N_30790);
and U39919 (N_39919,N_31782,N_33325);
and U39920 (N_39920,N_30004,N_30330);
nor U39921 (N_39921,N_31303,N_32619);
xor U39922 (N_39922,N_34023,N_31925);
or U39923 (N_39923,N_32246,N_30028);
or U39924 (N_39924,N_31500,N_30638);
or U39925 (N_39925,N_32598,N_32911);
nand U39926 (N_39926,N_32426,N_30118);
or U39927 (N_39927,N_34284,N_30043);
and U39928 (N_39928,N_32385,N_32607);
or U39929 (N_39929,N_31605,N_33611);
or U39930 (N_39930,N_31297,N_32409);
nand U39931 (N_39931,N_30977,N_30799);
or U39932 (N_39932,N_31096,N_31658);
and U39933 (N_39933,N_34803,N_30873);
nor U39934 (N_39934,N_32975,N_30087);
nand U39935 (N_39935,N_31627,N_30991);
nor U39936 (N_39936,N_33204,N_30601);
and U39937 (N_39937,N_30005,N_32379);
nand U39938 (N_39938,N_31792,N_31244);
xnor U39939 (N_39939,N_34300,N_32778);
or U39940 (N_39940,N_34182,N_34493);
and U39941 (N_39941,N_32760,N_32248);
or U39942 (N_39942,N_32778,N_33981);
nand U39943 (N_39943,N_30039,N_32582);
xor U39944 (N_39944,N_31417,N_32055);
xor U39945 (N_39945,N_34525,N_31261);
nor U39946 (N_39946,N_34008,N_32448);
xnor U39947 (N_39947,N_33132,N_32349);
nor U39948 (N_39948,N_34540,N_32242);
xnor U39949 (N_39949,N_30490,N_34700);
or U39950 (N_39950,N_32040,N_32365);
xnor U39951 (N_39951,N_34622,N_34518);
and U39952 (N_39952,N_30962,N_30707);
nor U39953 (N_39953,N_34324,N_34225);
xor U39954 (N_39954,N_30538,N_34315);
or U39955 (N_39955,N_30038,N_30555);
or U39956 (N_39956,N_30586,N_31129);
and U39957 (N_39957,N_34034,N_31720);
or U39958 (N_39958,N_30621,N_34754);
and U39959 (N_39959,N_31071,N_30871);
nor U39960 (N_39960,N_30450,N_30245);
xnor U39961 (N_39961,N_30287,N_32466);
xnor U39962 (N_39962,N_33468,N_34594);
nor U39963 (N_39963,N_33284,N_34900);
or U39964 (N_39964,N_30684,N_34231);
or U39965 (N_39965,N_34086,N_30746);
nand U39966 (N_39966,N_30592,N_30962);
nor U39967 (N_39967,N_34891,N_32596);
xor U39968 (N_39968,N_32427,N_34218);
nand U39969 (N_39969,N_34452,N_31137);
nor U39970 (N_39970,N_32577,N_30988);
or U39971 (N_39971,N_34344,N_30433);
nor U39972 (N_39972,N_33543,N_31893);
or U39973 (N_39973,N_30130,N_33123);
xor U39974 (N_39974,N_30002,N_32278);
xnor U39975 (N_39975,N_30860,N_33958);
xnor U39976 (N_39976,N_34722,N_31089);
or U39977 (N_39977,N_31276,N_30374);
xnor U39978 (N_39978,N_31562,N_32505);
xnor U39979 (N_39979,N_33349,N_33063);
or U39980 (N_39980,N_32169,N_33936);
and U39981 (N_39981,N_33493,N_34025);
xnor U39982 (N_39982,N_30614,N_30825);
xor U39983 (N_39983,N_31040,N_30963);
or U39984 (N_39984,N_34110,N_33247);
and U39985 (N_39985,N_30366,N_32244);
or U39986 (N_39986,N_32522,N_32847);
xor U39987 (N_39987,N_34605,N_34995);
nand U39988 (N_39988,N_33212,N_31303);
nand U39989 (N_39989,N_33743,N_34369);
nand U39990 (N_39990,N_30478,N_32216);
or U39991 (N_39991,N_30655,N_32497);
and U39992 (N_39992,N_31343,N_33433);
or U39993 (N_39993,N_33971,N_32671);
nand U39994 (N_39994,N_33895,N_33995);
xnor U39995 (N_39995,N_34442,N_34466);
nand U39996 (N_39996,N_30767,N_30788);
nor U39997 (N_39997,N_34600,N_34669);
xor U39998 (N_39998,N_33273,N_33748);
nor U39999 (N_39999,N_34917,N_32700);
nor U40000 (N_40000,N_37723,N_35909);
nor U40001 (N_40001,N_37921,N_36856);
xnor U40002 (N_40002,N_38275,N_37024);
nor U40003 (N_40003,N_37357,N_36992);
or U40004 (N_40004,N_39039,N_39281);
nor U40005 (N_40005,N_39772,N_38580);
nand U40006 (N_40006,N_35529,N_39589);
xor U40007 (N_40007,N_39502,N_39321);
and U40008 (N_40008,N_38908,N_35277);
nand U40009 (N_40009,N_36884,N_35645);
xor U40010 (N_40010,N_35172,N_36976);
and U40011 (N_40011,N_39179,N_35553);
xor U40012 (N_40012,N_37827,N_36215);
nand U40013 (N_40013,N_35445,N_39542);
nor U40014 (N_40014,N_37695,N_38759);
or U40015 (N_40015,N_35632,N_38902);
xor U40016 (N_40016,N_38661,N_36205);
or U40017 (N_40017,N_37093,N_36096);
and U40018 (N_40018,N_35948,N_37547);
nand U40019 (N_40019,N_37198,N_35256);
xor U40020 (N_40020,N_37822,N_36592);
or U40021 (N_40021,N_35204,N_39245);
xor U40022 (N_40022,N_35524,N_37929);
nand U40023 (N_40023,N_36582,N_36858);
nand U40024 (N_40024,N_38567,N_36488);
xor U40025 (N_40025,N_37499,N_39976);
nand U40026 (N_40026,N_35362,N_39751);
xnor U40027 (N_40027,N_39251,N_39145);
nor U40028 (N_40028,N_35346,N_39747);
nor U40029 (N_40029,N_35535,N_39963);
or U40030 (N_40030,N_36366,N_35706);
nand U40031 (N_40031,N_38290,N_37472);
nor U40032 (N_40032,N_38937,N_38488);
nand U40033 (N_40033,N_37603,N_36612);
nor U40034 (N_40034,N_36514,N_37879);
nand U40035 (N_40035,N_37164,N_36193);
nand U40036 (N_40036,N_38552,N_36028);
nor U40037 (N_40037,N_38927,N_38970);
nor U40038 (N_40038,N_37758,N_36532);
xnor U40039 (N_40039,N_37911,N_37835);
nand U40040 (N_40040,N_36484,N_38781);
and U40041 (N_40041,N_37548,N_38144);
nand U40042 (N_40042,N_38260,N_37288);
and U40043 (N_40043,N_35967,N_37173);
xor U40044 (N_40044,N_37149,N_36122);
xnor U40045 (N_40045,N_35578,N_35726);
nor U40046 (N_40046,N_37229,N_39022);
or U40047 (N_40047,N_35890,N_38160);
nor U40048 (N_40048,N_36168,N_38663);
or U40049 (N_40049,N_38324,N_35205);
nor U40050 (N_40050,N_35418,N_35989);
and U40051 (N_40051,N_37242,N_36460);
xnor U40052 (N_40052,N_38001,N_38996);
and U40053 (N_40053,N_35298,N_35244);
xnor U40054 (N_40054,N_37171,N_37840);
nand U40055 (N_40055,N_36424,N_36436);
nor U40056 (N_40056,N_36453,N_37832);
and U40057 (N_40057,N_39010,N_35474);
and U40058 (N_40058,N_38120,N_38691);
or U40059 (N_40059,N_37086,N_35022);
xor U40060 (N_40060,N_35426,N_35801);
and U40061 (N_40061,N_38504,N_38683);
and U40062 (N_40062,N_35634,N_35109);
nor U40063 (N_40063,N_36165,N_39773);
and U40064 (N_40064,N_35211,N_39319);
or U40065 (N_40065,N_39551,N_35379);
nand U40066 (N_40066,N_38130,N_38039);
xor U40067 (N_40067,N_39209,N_37128);
and U40068 (N_40068,N_38490,N_37477);
nor U40069 (N_40069,N_36570,N_37251);
or U40070 (N_40070,N_39725,N_38826);
nor U40071 (N_40071,N_39811,N_36386);
xor U40072 (N_40072,N_38242,N_36253);
nor U40073 (N_40073,N_35284,N_36023);
or U40074 (N_40074,N_38869,N_35302);
xor U40075 (N_40075,N_39442,N_36075);
nor U40076 (N_40076,N_37290,N_38430);
nand U40077 (N_40077,N_35233,N_37215);
nand U40078 (N_40078,N_35491,N_39930);
or U40079 (N_40079,N_39396,N_39866);
nand U40080 (N_40080,N_36316,N_35365);
or U40081 (N_40081,N_37464,N_38117);
and U40082 (N_40082,N_38388,N_36723);
or U40083 (N_40083,N_39633,N_36815);
or U40084 (N_40084,N_39878,N_37436);
or U40085 (N_40085,N_35138,N_39398);
nand U40086 (N_40086,N_36093,N_39750);
nor U40087 (N_40087,N_36236,N_37543);
nor U40088 (N_40088,N_38443,N_37742);
xnor U40089 (N_40089,N_39112,N_35325);
or U40090 (N_40090,N_35950,N_39777);
or U40091 (N_40091,N_36701,N_36050);
and U40092 (N_40092,N_37442,N_36523);
nand U40093 (N_40093,N_38178,N_39832);
xor U40094 (N_40094,N_38100,N_37587);
and U40095 (N_40095,N_36382,N_36969);
nor U40096 (N_40096,N_39186,N_35031);
nor U40097 (N_40097,N_36932,N_36194);
xnor U40098 (N_40098,N_35131,N_39044);
nor U40099 (N_40099,N_38159,N_38833);
xor U40100 (N_40100,N_36005,N_37344);
or U40101 (N_40101,N_37939,N_38838);
nand U40102 (N_40102,N_38960,N_39820);
nand U40103 (N_40103,N_38135,N_37932);
nor U40104 (N_40104,N_36014,N_38403);
xor U40105 (N_40105,N_37381,N_37775);
and U40106 (N_40106,N_39916,N_36825);
nor U40107 (N_40107,N_39220,N_39570);
or U40108 (N_40108,N_36358,N_37841);
xnor U40109 (N_40109,N_37618,N_35758);
nor U40110 (N_40110,N_38813,N_35868);
xnor U40111 (N_40111,N_35020,N_37426);
xor U40112 (N_40112,N_38727,N_35943);
nor U40113 (N_40113,N_39320,N_39051);
nand U40114 (N_40114,N_38844,N_39523);
and U40115 (N_40115,N_38456,N_35595);
and U40116 (N_40116,N_39060,N_35877);
xor U40117 (N_40117,N_39835,N_38731);
nor U40118 (N_40118,N_39505,N_35518);
or U40119 (N_40119,N_38498,N_39488);
and U40120 (N_40120,N_38177,N_39315);
xor U40121 (N_40121,N_38419,N_37162);
xnor U40122 (N_40122,N_36718,N_38478);
nand U40123 (N_40123,N_38469,N_37201);
or U40124 (N_40124,N_35384,N_36148);
xnor U40125 (N_40125,N_38263,N_35644);
xor U40126 (N_40126,N_37525,N_38939);
nand U40127 (N_40127,N_38817,N_39225);
nand U40128 (N_40128,N_35755,N_35123);
and U40129 (N_40129,N_37757,N_36384);
or U40130 (N_40130,N_39983,N_38816);
xor U40131 (N_40131,N_37546,N_38695);
or U40132 (N_40132,N_39541,N_36729);
and U40133 (N_40133,N_36266,N_37561);
or U40134 (N_40134,N_39250,N_36027);
and U40135 (N_40135,N_39170,N_35319);
or U40136 (N_40136,N_35923,N_37038);
nand U40137 (N_40137,N_38630,N_39533);
or U40138 (N_40138,N_39036,N_37174);
nand U40139 (N_40139,N_38739,N_35729);
nor U40140 (N_40140,N_35059,N_38107);
or U40141 (N_40141,N_38044,N_35704);
nor U40142 (N_40142,N_35028,N_35224);
nand U40143 (N_40143,N_35519,N_37953);
and U40144 (N_40144,N_36016,N_39338);
and U40145 (N_40145,N_38397,N_35276);
xnor U40146 (N_40146,N_37247,N_36954);
nand U40147 (N_40147,N_37334,N_36130);
xor U40148 (N_40148,N_35452,N_38672);
nor U40149 (N_40149,N_36048,N_39719);
nand U40150 (N_40150,N_36774,N_37973);
or U40151 (N_40151,N_37816,N_36784);
and U40152 (N_40152,N_38035,N_35293);
nand U40153 (N_40153,N_39588,N_35710);
nor U40154 (N_40154,N_36792,N_39681);
nor U40155 (N_40155,N_38602,N_35235);
nor U40156 (N_40156,N_39208,N_36750);
nand U40157 (N_40157,N_37387,N_35778);
nor U40158 (N_40158,N_36051,N_38866);
and U40159 (N_40159,N_39810,N_38934);
nand U40160 (N_40160,N_39642,N_36281);
nand U40161 (N_40161,N_35451,N_39525);
nor U40162 (N_40162,N_35528,N_36212);
nor U40163 (N_40163,N_35148,N_38936);
nor U40164 (N_40164,N_39363,N_39974);
xnor U40165 (N_40165,N_38392,N_39439);
nor U40166 (N_40166,N_39047,N_35843);
and U40167 (N_40167,N_36150,N_36272);
xnor U40168 (N_40168,N_35825,N_39775);
nor U40169 (N_40169,N_36035,N_35157);
nand U40170 (N_40170,N_39114,N_35613);
nor U40171 (N_40171,N_36249,N_39723);
xor U40172 (N_40172,N_39796,N_38226);
xor U40173 (N_40173,N_39211,N_39556);
nor U40174 (N_40174,N_38991,N_39131);
nand U40175 (N_40175,N_36221,N_37943);
or U40176 (N_40176,N_36605,N_35116);
xor U40177 (N_40177,N_35337,N_37813);
nand U40178 (N_40178,N_37498,N_36095);
nand U40179 (N_40179,N_37506,N_39380);
or U40180 (N_40180,N_38550,N_39507);
nand U40181 (N_40181,N_39021,N_37398);
nor U40182 (N_40182,N_35942,N_35567);
xnor U40183 (N_40183,N_35894,N_37443);
or U40184 (N_40184,N_39711,N_37428);
or U40185 (N_40185,N_38264,N_35620);
and U40186 (N_40186,N_38283,N_36434);
nor U40187 (N_40187,N_37274,N_37884);
xnor U40188 (N_40188,N_39361,N_37747);
nand U40189 (N_40189,N_35096,N_37914);
xnor U40190 (N_40190,N_36588,N_35262);
nand U40191 (N_40191,N_36099,N_38616);
or U40192 (N_40192,N_36581,N_36039);
xor U40193 (N_40193,N_36388,N_38357);
and U40194 (N_40194,N_38441,N_35464);
and U40195 (N_40195,N_36821,N_36720);
nor U40196 (N_40196,N_36673,N_38969);
or U40197 (N_40197,N_38855,N_36848);
nand U40198 (N_40198,N_38423,N_35124);
nand U40199 (N_40199,N_38832,N_39953);
or U40200 (N_40200,N_38500,N_38646);
or U40201 (N_40201,N_35514,N_39168);
nor U40202 (N_40202,N_38598,N_38581);
nor U40203 (N_40203,N_35132,N_37692);
and U40204 (N_40204,N_35380,N_38474);
or U40205 (N_40205,N_38089,N_37704);
and U40206 (N_40206,N_35169,N_37016);
or U40207 (N_40207,N_38576,N_38401);
xnor U40208 (N_40208,N_39341,N_38992);
nor U40209 (N_40209,N_35347,N_39142);
xnor U40210 (N_40210,N_36807,N_38561);
or U40211 (N_40211,N_35711,N_38217);
or U40212 (N_40212,N_38626,N_36136);
nor U40213 (N_40213,N_38252,N_38479);
nor U40214 (N_40214,N_39804,N_35676);
and U40215 (N_40215,N_35505,N_36875);
nand U40216 (N_40216,N_38148,N_35822);
nand U40217 (N_40217,N_38657,N_37330);
nand U40218 (N_40218,N_39371,N_39115);
and U40219 (N_40219,N_35984,N_36070);
nor U40220 (N_40220,N_36461,N_36563);
or U40221 (N_40221,N_36579,N_37262);
or U40222 (N_40222,N_39276,N_39692);
and U40223 (N_40223,N_37266,N_39237);
and U40224 (N_40224,N_38468,N_39936);
or U40225 (N_40225,N_38231,N_36534);
and U40226 (N_40226,N_35087,N_35078);
or U40227 (N_40227,N_37748,N_36731);
or U40228 (N_40228,N_35777,N_35062);
nand U40229 (N_40229,N_37053,N_38734);
and U40230 (N_40230,N_37912,N_38076);
and U40231 (N_40231,N_39076,N_35639);
or U40232 (N_40232,N_38821,N_36738);
nand U40233 (N_40233,N_37018,N_37135);
or U40234 (N_40234,N_35428,N_37046);
xnor U40235 (N_40235,N_35623,N_35986);
nor U40236 (N_40236,N_37388,N_38282);
nand U40237 (N_40237,N_38358,N_37806);
or U40238 (N_40238,N_38890,N_39040);
nor U40239 (N_40239,N_37651,N_36827);
nand U40240 (N_40240,N_36061,N_36066);
or U40241 (N_40241,N_39347,N_35137);
xor U40242 (N_40242,N_35378,N_35376);
xnor U40243 (N_40243,N_37314,N_38095);
nor U40244 (N_40244,N_36322,N_35831);
or U40245 (N_40245,N_39616,N_35545);
xnor U40246 (N_40246,N_35876,N_37390);
xnor U40247 (N_40247,N_36739,N_35306);
nand U40248 (N_40248,N_37446,N_38942);
or U40249 (N_40249,N_37803,N_39028);
nor U40250 (N_40250,N_37085,N_38235);
and U40251 (N_40251,N_39275,N_37938);
or U40252 (N_40252,N_36567,N_38917);
nor U40253 (N_40253,N_35811,N_38415);
xor U40254 (N_40254,N_36258,N_37975);
nor U40255 (N_40255,N_39912,N_35775);
nor U40256 (N_40256,N_35725,N_37203);
nor U40257 (N_40257,N_38863,N_37719);
xor U40258 (N_40258,N_36776,N_39664);
xor U40259 (N_40259,N_39892,N_37327);
or U40260 (N_40260,N_36345,N_39924);
or U40261 (N_40261,N_37819,N_37836);
nor U40262 (N_40262,N_39676,N_35867);
nand U40263 (N_40263,N_35506,N_38523);
and U40264 (N_40264,N_38239,N_35992);
and U40265 (N_40265,N_39537,N_38472);
xnor U40266 (N_40266,N_38615,N_39137);
and U40267 (N_40267,N_35566,N_39941);
nand U40268 (N_40268,N_39235,N_39867);
nand U40269 (N_40269,N_35902,N_37602);
nand U40270 (N_40270,N_36472,N_37319);
nor U40271 (N_40271,N_37647,N_35438);
nand U40272 (N_40272,N_37689,N_37453);
xnor U40273 (N_40273,N_38245,N_37966);
nand U40274 (N_40274,N_38475,N_38434);
xor U40275 (N_40275,N_39718,N_37555);
and U40276 (N_40276,N_38929,N_38604);
or U40277 (N_40277,N_39543,N_39012);
nand U40278 (N_40278,N_38671,N_39094);
xor U40279 (N_40279,N_36317,N_35227);
or U40280 (N_40280,N_39492,N_36965);
nor U40281 (N_40281,N_39253,N_36564);
xnor U40282 (N_40282,N_35317,N_35118);
and U40283 (N_40283,N_37040,N_35274);
xor U40284 (N_40284,N_38447,N_35812);
xnor U40285 (N_40285,N_37562,N_36115);
xor U40286 (N_40286,N_37361,N_35421);
xor U40287 (N_40287,N_36762,N_39068);
nand U40288 (N_40288,N_39070,N_37339);
and U40289 (N_40289,N_36600,N_36397);
or U40290 (N_40290,N_39462,N_38648);
and U40291 (N_40291,N_39101,N_35593);
and U40292 (N_40292,N_35795,N_35653);
or U40293 (N_40293,N_38020,N_36730);
nand U40294 (N_40294,N_38097,N_39998);
or U40295 (N_40295,N_35178,N_35579);
and U40296 (N_40296,N_37280,N_38494);
and U40297 (N_40297,N_38225,N_39697);
and U40298 (N_40298,N_36601,N_37877);
and U40299 (N_40299,N_35839,N_37125);
nand U40300 (N_40300,N_39727,N_37277);
or U40301 (N_40301,N_35463,N_36758);
xnor U40302 (N_40302,N_36407,N_37531);
xnor U40303 (N_40303,N_35181,N_39746);
nand U40304 (N_40304,N_35727,N_39149);
xor U40305 (N_40305,N_39814,N_39509);
nor U40306 (N_40306,N_37631,N_39590);
xnor U40307 (N_40307,N_39860,N_35918);
nor U40308 (N_40308,N_37788,N_36062);
xor U40309 (N_40309,N_35366,N_36209);
nand U40310 (N_40310,N_39298,N_39368);
nor U40311 (N_40311,N_38935,N_38795);
nor U40312 (N_40312,N_35817,N_36896);
or U40313 (N_40313,N_37480,N_39739);
and U40314 (N_40314,N_37050,N_39215);
xor U40315 (N_40315,N_35335,N_37530);
nand U40316 (N_40316,N_36192,N_38753);
or U40317 (N_40317,N_36157,N_37590);
nand U40318 (N_40318,N_35794,N_39914);
nor U40319 (N_40319,N_36337,N_37102);
xor U40320 (N_40320,N_37485,N_38512);
nor U40321 (N_40321,N_39701,N_37569);
and U40322 (N_40322,N_36552,N_38063);
and U40323 (N_40323,N_39348,N_36142);
nor U40324 (N_40324,N_36808,N_38293);
nor U40325 (N_40325,N_38328,N_39444);
xnor U40326 (N_40326,N_39248,N_36371);
xnor U40327 (N_40327,N_39651,N_37897);
nor U40328 (N_40328,N_39562,N_35196);
xnor U40329 (N_40329,N_37131,N_39325);
nor U40330 (N_40330,N_35643,N_38574);
or U40331 (N_40331,N_35760,N_35815);
xor U40332 (N_40332,N_36981,N_37764);
xnor U40333 (N_40333,N_38516,N_38954);
xor U40334 (N_40334,N_36110,N_39636);
nor U40335 (N_40335,N_36970,N_37513);
nor U40336 (N_40336,N_37267,N_37500);
nand U40337 (N_40337,N_36753,N_38705);
or U40338 (N_40338,N_36541,N_38366);
xor U40339 (N_40339,N_38674,N_39143);
nor U40340 (N_40340,N_35879,N_37154);
and U40341 (N_40341,N_39576,N_38306);
nand U40342 (N_40342,N_39201,N_38059);
or U40343 (N_40343,N_39546,N_39567);
and U40344 (N_40344,N_39313,N_35935);
nand U40345 (N_40345,N_37739,N_36707);
xor U40346 (N_40346,N_39083,N_37430);
and U40347 (N_40347,N_35003,N_37456);
nor U40348 (N_40348,N_36084,N_36603);
nand U40349 (N_40349,N_36880,N_37249);
and U40350 (N_40350,N_39691,N_38215);
nor U40351 (N_40351,N_39432,N_38182);
nor U40352 (N_40352,N_35025,N_37657);
or U40353 (N_40353,N_35300,N_39715);
nor U40354 (N_40354,N_37915,N_38706);
and U40355 (N_40355,N_37101,N_37654);
nand U40356 (N_40356,N_35265,N_39180);
or U40357 (N_40357,N_38741,N_37948);
xnor U40358 (N_40358,N_38414,N_38973);
and U40359 (N_40359,N_36917,N_35083);
or U40360 (N_40360,N_38887,N_38880);
nand U40361 (N_40361,N_38670,N_35446);
or U40362 (N_40362,N_39957,N_39932);
or U40363 (N_40363,N_39359,N_37650);
xnor U40364 (N_40364,N_39929,N_39880);
xnor U40365 (N_40365,N_38334,N_36100);
nor U40366 (N_40366,N_38905,N_39034);
nand U40367 (N_40367,N_35997,N_35521);
xor U40368 (N_40368,N_37260,N_38008);
xnor U40369 (N_40369,N_37861,N_39939);
nor U40370 (N_40370,N_37801,N_37312);
nand U40371 (N_40371,N_36539,N_37400);
and U40372 (N_40372,N_36881,N_36224);
nor U40373 (N_40373,N_35896,N_38590);
nor U40374 (N_40374,N_36922,N_37575);
nor U40375 (N_40375,N_36370,N_36405);
or U40376 (N_40376,N_39285,N_35938);
and U40377 (N_40377,N_39879,N_36616);
xnor U40378 (N_40378,N_38575,N_38014);
and U40379 (N_40379,N_38372,N_37325);
nor U40380 (N_40380,N_36107,N_38399);
nand U40381 (N_40381,N_36659,N_35226);
xnor U40382 (N_40382,N_35947,N_37054);
or U40383 (N_40383,N_37843,N_38825);
or U40384 (N_40384,N_39203,N_35499);
or U40385 (N_40385,N_38104,N_36556);
or U40386 (N_40386,N_38061,N_37702);
xnor U40387 (N_40387,N_35416,N_36331);
xnor U40388 (N_40388,N_37521,N_35323);
or U40389 (N_40389,N_36147,N_39877);
and U40390 (N_40390,N_37963,N_37550);
xnor U40391 (N_40391,N_38466,N_36483);
and U40392 (N_40392,N_35228,N_35952);
xor U40393 (N_40393,N_35720,N_36744);
or U40394 (N_40394,N_37039,N_35170);
or U40395 (N_40395,N_36938,N_39874);
or U40396 (N_40396,N_36132,N_36949);
nand U40397 (N_40397,N_38452,N_35674);
nand U40398 (N_40398,N_35372,N_36485);
nand U40399 (N_40399,N_36172,N_37217);
and U40400 (N_40400,N_35949,N_35468);
xor U40401 (N_40401,N_35910,N_38187);
or U40402 (N_40402,N_37675,N_37823);
nor U40403 (N_40403,N_36412,N_38493);
and U40404 (N_40404,N_37165,N_36933);
xnor U40405 (N_40405,N_36913,N_36839);
nand U40406 (N_40406,N_35987,N_35539);
and U40407 (N_40407,N_37828,N_38322);
or U40408 (N_40408,N_35016,N_36230);
xnor U40409 (N_40409,N_39569,N_37553);
xnor U40410 (N_40410,N_35012,N_37401);
nand U40411 (N_40411,N_35456,N_38158);
xor U40412 (N_40412,N_35991,N_35677);
nor U40413 (N_40413,N_36843,N_37415);
and U40414 (N_40414,N_35483,N_37954);
and U40415 (N_40415,N_35312,N_38715);
xnor U40416 (N_40416,N_36112,N_37504);
and U40417 (N_40417,N_37981,N_39062);
nand U40418 (N_40418,N_35387,N_36072);
or U40419 (N_40419,N_37126,N_38726);
or U40420 (N_40420,N_37540,N_39106);
nand U40421 (N_40421,N_38628,N_36270);
xor U40422 (N_40422,N_35916,N_36809);
nor U40423 (N_40423,N_36983,N_38595);
and U40424 (N_40424,N_37871,N_37526);
nor U40425 (N_40425,N_37382,N_37920);
and U40426 (N_40426,N_39922,N_38644);
or U40427 (N_40427,N_36754,N_39210);
or U40428 (N_40428,N_37536,N_39061);
xnor U40429 (N_40429,N_36324,N_39284);
xor U40430 (N_40430,N_35127,N_36625);
and U40431 (N_40431,N_38304,N_37449);
or U40432 (N_40432,N_38658,N_36114);
nand U40433 (N_40433,N_36479,N_37123);
xor U40434 (N_40434,N_37141,N_38482);
nand U40435 (N_40435,N_35749,N_37609);
and U40436 (N_40436,N_36262,N_37652);
xor U40437 (N_40437,N_35609,N_39863);
and U40438 (N_40438,N_38820,N_39489);
or U40439 (N_40439,N_38874,N_38766);
and U40440 (N_40440,N_36246,N_39601);
xnor U40441 (N_40441,N_38128,N_38547);
nand U40442 (N_40442,N_36134,N_39103);
nand U40443 (N_40443,N_37916,N_36285);
and U40444 (N_40444,N_35957,N_38471);
nand U40445 (N_40445,N_39408,N_38704);
nand U40446 (N_40446,N_36446,N_38974);
nand U40447 (N_40447,N_36926,N_36389);
nor U40448 (N_40448,N_37490,N_36013);
xor U40449 (N_40449,N_38463,N_37892);
xnor U40450 (N_40450,N_37202,N_35614);
nor U40451 (N_40451,N_35305,N_35963);
nand U40452 (N_40452,N_39286,N_37471);
or U40453 (N_40453,N_38112,N_35391);
nand U40454 (N_40454,N_39078,N_35834);
and U40455 (N_40455,N_39845,N_35819);
or U40456 (N_40456,N_38300,N_38241);
nor U40457 (N_40457,N_37077,N_35906);
nor U40458 (N_40458,N_37311,N_38621);
nand U40459 (N_40459,N_37391,N_36861);
or U40460 (N_40460,N_36895,N_35734);
or U40461 (N_40461,N_39053,N_38331);
and U40462 (N_40462,N_37493,N_38899);
nand U40463 (N_40463,N_36174,N_35102);
xor U40464 (N_40464,N_35513,N_37476);
xor U40465 (N_40465,N_35691,N_35163);
nor U40466 (N_40466,N_38732,N_37419);
or U40467 (N_40467,N_39228,N_37354);
xnor U40468 (N_40468,N_36458,N_37061);
and U40469 (N_40469,N_39423,N_38513);
xnor U40470 (N_40470,N_35556,N_36457);
xnor U40471 (N_40471,N_39352,N_35719);
xor U40472 (N_40472,N_36801,N_37643);
and U40473 (N_40473,N_36392,N_38639);
nand U40474 (N_40474,N_36678,N_35282);
nand U40475 (N_40475,N_37514,N_39227);
xor U40476 (N_40476,N_35125,N_35253);
xor U40477 (N_40477,N_37495,N_37027);
and U40478 (N_40478,N_39872,N_36629);
xnor U40479 (N_40479,N_37740,N_39650);
or U40480 (N_40480,N_38713,N_36214);
nor U40481 (N_40481,N_38794,N_38889);
and U40482 (N_40482,N_35437,N_39096);
or U40483 (N_40483,N_39230,N_36996);
or U40484 (N_40484,N_36300,N_39638);
xnor U40485 (N_40485,N_36845,N_36440);
xnor U40486 (N_40486,N_39198,N_35238);
nor U40487 (N_40487,N_39896,N_37263);
and U40488 (N_40488,N_35517,N_37935);
and U40489 (N_40489,N_39294,N_35806);
or U40490 (N_40490,N_39148,N_35339);
and U40491 (N_40491,N_39175,N_35728);
or U40492 (N_40492,N_35304,N_39519);
or U40493 (N_40493,N_39274,N_38216);
and U40494 (N_40494,N_36007,N_37629);
xnor U40495 (N_40495,N_38022,N_39770);
nand U40496 (N_40496,N_38873,N_38707);
and U40497 (N_40497,N_38611,N_37238);
xor U40498 (N_40498,N_37397,N_35884);
and U40499 (N_40499,N_36773,N_39241);
and U40500 (N_40500,N_36906,N_35833);
xor U40501 (N_40501,N_38417,N_37900);
nand U40502 (N_40502,N_38383,N_36709);
or U40503 (N_40503,N_36368,N_38023);
xor U40504 (N_40504,N_36203,N_39379);
or U40505 (N_40505,N_35219,N_36053);
nand U40506 (N_40506,N_38398,N_39194);
nand U40507 (N_40507,N_38975,N_39736);
nand U40508 (N_40508,N_37922,N_38932);
nand U40509 (N_40509,N_35368,N_39960);
or U40510 (N_40510,N_37990,N_38218);
and U40511 (N_40511,N_38859,N_36610);
or U40512 (N_40512,N_36507,N_37055);
or U40513 (N_40513,N_37451,N_35097);
or U40514 (N_40514,N_35352,N_39048);
or U40515 (N_40515,N_37684,N_35142);
and U40516 (N_40516,N_39921,N_36771);
and U40517 (N_40517,N_37292,N_39434);
and U40518 (N_40518,N_35269,N_35095);
and U40519 (N_40519,N_38315,N_38316);
nor U40520 (N_40520,N_36671,N_38277);
or U40521 (N_40521,N_37231,N_37600);
or U40522 (N_40522,N_38738,N_36494);
xnor U40523 (N_40523,N_37193,N_39803);
xnor U40524 (N_40524,N_37291,N_37160);
or U40525 (N_40525,N_38752,N_36664);
and U40526 (N_40526,N_36390,N_37411);
and U40527 (N_40527,N_39837,N_36269);
and U40528 (N_40528,N_37974,N_37621);
and U40529 (N_40529,N_35073,N_35479);
nand U40530 (N_40530,N_35326,N_39580);
xnor U40531 (N_40531,N_37904,N_36538);
or U40532 (N_40532,N_36010,N_37244);
or U40533 (N_40533,N_36682,N_38000);
or U40534 (N_40534,N_35334,N_39031);
nor U40535 (N_40535,N_36662,N_35694);
nand U40536 (N_40536,N_35254,N_38990);
xnor U40537 (N_40537,N_37091,N_38108);
nor U40538 (N_40538,N_36463,N_36078);
xor U40539 (N_40539,N_39173,N_37581);
or U40540 (N_40540,N_35841,N_36660);
and U40541 (N_40541,N_38074,N_35576);
or U40542 (N_40542,N_38754,N_35946);
or U40543 (N_40543,N_36726,N_35864);
xor U40544 (N_40544,N_37967,N_37044);
nor U40545 (N_40545,N_35121,N_38485);
nand U40546 (N_40546,N_37591,N_38094);
or U40547 (N_40547,N_38768,N_38229);
or U40548 (N_40548,N_35531,N_35607);
and U40549 (N_40549,N_36443,N_39670);
and U40550 (N_40550,N_36737,N_35444);
nor U40551 (N_40551,N_38110,N_36639);
xnor U40552 (N_40552,N_36973,N_36356);
nand U40553 (N_40553,N_35069,N_37095);
or U40554 (N_40554,N_39392,N_35592);
xor U40555 (N_40555,N_36781,N_37004);
or U40556 (N_40556,N_36456,N_39610);
xor U40557 (N_40557,N_35060,N_37824);
nor U40558 (N_40558,N_38017,N_36763);
or U40559 (N_40559,N_36886,N_39608);
nor U40560 (N_40560,N_35686,N_37894);
or U40561 (N_40561,N_36591,N_37750);
or U40562 (N_40562,N_38530,N_36780);
nor U40563 (N_40563,N_37956,N_36242);
and U40564 (N_40564,N_35321,N_36942);
nand U40565 (N_40565,N_38814,N_38151);
nor U40566 (N_40566,N_36474,N_37011);
nor U40567 (N_40567,N_37985,N_39122);
nand U40568 (N_40568,N_37902,N_37118);
or U40569 (N_40569,N_37888,N_36898);
xor U40570 (N_40570,N_36788,N_37106);
or U40571 (N_40571,N_37958,N_35907);
and U40572 (N_40572,N_35920,N_38026);
nor U40573 (N_40573,N_37554,N_35005);
or U40574 (N_40574,N_38435,N_36510);
nor U40575 (N_40575,N_35435,N_37982);
or U40576 (N_40576,N_37414,N_38649);
nand U40577 (N_40577,N_37649,N_36001);
nand U40578 (N_40578,N_38004,N_36513);
nand U40579 (N_40579,N_36802,N_38308);
nand U40580 (N_40580,N_37984,N_36073);
xnor U40581 (N_40581,N_37971,N_39102);
or U40582 (N_40582,N_38154,N_37003);
xor U40583 (N_40583,N_35144,N_39920);
nand U40584 (N_40584,N_39428,N_37056);
xnor U40585 (N_40585,N_36057,N_38634);
nor U40586 (N_40586,N_36951,N_38665);
xor U40587 (N_40587,N_36467,N_37403);
xnor U40588 (N_40588,N_38594,N_35332);
xor U40589 (N_40589,N_35252,N_36298);
or U40590 (N_40590,N_35849,N_37439);
and U40591 (N_40591,N_38786,N_37028);
xnor U40592 (N_40592,N_38565,N_38223);
and U40593 (N_40593,N_36844,N_37728);
xnor U40594 (N_40594,N_36840,N_39020);
or U40595 (N_40595,N_36622,N_38473);
nand U40596 (N_40596,N_38164,N_35548);
nor U40597 (N_40597,N_35600,N_37763);
and U40598 (N_40598,N_36188,N_37298);
or U40599 (N_40599,N_39885,N_36022);
nor U40600 (N_40600,N_36235,N_37156);
and U40601 (N_40601,N_35612,N_36841);
nand U40602 (N_40602,N_39130,N_39729);
nand U40603 (N_40603,N_38756,N_37299);
nor U40604 (N_40604,N_35616,N_37596);
or U40605 (N_40605,N_38395,N_38746);
xnor U40606 (N_40606,N_36223,N_39309);
or U40607 (N_40607,N_37735,N_37437);
nor U40608 (N_40608,N_35465,N_36451);
and U40609 (N_40609,N_37103,N_37712);
and U40610 (N_40610,N_39037,N_35936);
xor U40611 (N_40611,N_35515,N_37573);
nand U40612 (N_40612,N_35275,N_38486);
nor U40613 (N_40613,N_35603,N_36459);
or U40614 (N_40614,N_39190,N_35861);
nand U40615 (N_40615,N_38484,N_36422);
or U40616 (N_40616,N_36716,N_39630);
or U40617 (N_40617,N_38172,N_38262);
and U40618 (N_40618,N_38278,N_35742);
or U40619 (N_40619,N_36857,N_37852);
or U40620 (N_40620,N_35808,N_35079);
nor U40621 (N_40621,N_39536,N_38933);
nor U40622 (N_40622,N_37286,N_38122);
and U40623 (N_40623,N_39495,N_39862);
nor U40624 (N_40624,N_39574,N_37194);
nor U40625 (N_40625,N_37754,N_39433);
or U40626 (N_40626,N_38963,N_38281);
xor U40627 (N_40627,N_37374,N_35045);
or U40628 (N_40628,N_36522,N_39358);
xor U40629 (N_40629,N_37020,N_37834);
xor U40630 (N_40630,N_39264,N_38961);
and U40631 (N_40631,N_38583,N_37508);
and U40632 (N_40632,N_35941,N_36817);
xnor U40633 (N_40633,N_38904,N_37876);
nand U40634 (N_40634,N_38194,N_38666);
or U40635 (N_40635,N_37110,N_35375);
xnor U40636 (N_40636,N_36111,N_36243);
or U40637 (N_40637,N_39985,N_36077);
and U40638 (N_40638,N_35540,N_35192);
nand U40639 (N_40639,N_36959,N_39594);
or U40640 (N_40640,N_37371,N_36068);
or U40641 (N_40641,N_38142,N_35359);
nand U40642 (N_40642,N_38668,N_39377);
nor U40643 (N_40643,N_39654,N_35286);
nor U40644 (N_40644,N_35635,N_37632);
nor U40645 (N_40645,N_39579,N_35744);
nand U40646 (N_40646,N_39282,N_39015);
nor U40647 (N_40647,N_39024,N_36182);
nor U40648 (N_40648,N_38232,N_38455);
or U40649 (N_40649,N_38424,N_38072);
or U40650 (N_40650,N_35712,N_37870);
or U40651 (N_40651,N_36128,N_38519);
and U40652 (N_40652,N_38643,N_37356);
or U40653 (N_40653,N_39655,N_38841);
or U40654 (N_40654,N_37706,N_37640);
xor U40655 (N_40655,N_35713,N_36064);
xnor U40656 (N_40656,N_36184,N_37161);
and U40657 (N_40657,N_39003,N_36376);
xnor U40658 (N_40658,N_37962,N_39113);
nand U40659 (N_40659,N_37404,N_38957);
nor U40660 (N_40660,N_35313,N_39217);
or U40661 (N_40661,N_37599,N_37365);
or U40662 (N_40662,N_36395,N_36225);
and U40663 (N_40663,N_35164,N_39612);
or U40664 (N_40664,N_39384,N_36206);
nand U40665 (N_40665,N_38579,N_38845);
and U40666 (N_40666,N_37905,N_35046);
nand U40667 (N_40667,N_38735,N_37968);
or U40668 (N_40668,N_35182,N_38408);
nand U40669 (N_40669,N_37794,N_39997);
and U40670 (N_40670,N_38425,N_37349);
or U40671 (N_40671,N_36086,N_37753);
and U40672 (N_40672,N_36469,N_37478);
xnor U40673 (N_40673,N_38551,N_38679);
or U40674 (N_40674,N_36185,N_36200);
nand U40675 (N_40675,N_39204,N_36432);
xor U40676 (N_40676,N_35968,N_38296);
xor U40677 (N_40677,N_38137,N_38327);
nand U40678 (N_40678,N_35011,N_38313);
nand U40679 (N_40679,N_36340,N_38355);
nand U40680 (N_40680,N_37475,N_37423);
or U40681 (N_40681,N_36597,N_35122);
or U40682 (N_40682,N_35648,N_38722);
and U40683 (N_40683,N_36287,N_35000);
xnor U40684 (N_40684,N_38714,N_35889);
xor U40685 (N_40685,N_35975,N_35068);
nand U40686 (N_40686,N_36850,N_35824);
xnor U40687 (N_40687,N_38188,N_37283);
or U40688 (N_40688,N_36167,N_38828);
xnor U40689 (N_40689,N_36855,N_39069);
nor U40690 (N_40690,N_39337,N_39430);
xnor U40691 (N_40691,N_35433,N_35194);
or U40692 (N_40692,N_38013,N_38654);
nand U40693 (N_40693,N_35113,N_39369);
or U40694 (N_40694,N_39722,N_39171);
or U40695 (N_40695,N_38601,N_35774);
and U40696 (N_40696,N_39386,N_35427);
xor U40697 (N_40697,N_38553,N_39511);
nor U40698 (N_40698,N_35225,N_38351);
or U40699 (N_40699,N_35919,N_39534);
nor U40700 (N_40700,N_38462,N_39893);
and U40701 (N_40701,N_38389,N_36890);
nor U40702 (N_40702,N_37996,N_36198);
nor U40703 (N_40703,N_36336,N_38692);
or U40704 (N_40704,N_37729,N_39197);
xnor U40705 (N_40705,N_38546,N_39455);
or U40706 (N_40706,N_37137,N_35084);
xnor U40707 (N_40707,N_39496,N_39402);
nor U40708 (N_40708,N_35114,N_38767);
and U40709 (N_40709,N_36863,N_37383);
nand U40710 (N_40710,N_38511,N_37771);
nor U40711 (N_40711,N_39512,N_39571);
nor U40712 (N_40712,N_37316,N_35061);
xnor U40713 (N_40713,N_37326,N_36296);
and U40714 (N_40714,N_38367,N_38165);
or U40715 (N_40715,N_37470,N_35858);
nand U40716 (N_40716,N_37792,N_35569);
xor U40717 (N_40717,N_36191,N_37969);
or U40718 (N_40718,N_35422,N_36162);
or U40719 (N_40719,N_38949,N_35747);
nor U40720 (N_40720,N_35240,N_36279);
nor U40721 (N_40721,N_35027,N_38209);
xnor U40722 (N_40722,N_38977,N_39159);
nand U40723 (N_40723,N_39678,N_38180);
xor U40724 (N_40724,N_38019,N_36691);
nor U40725 (N_40725,N_35598,N_35088);
or U40726 (N_40726,N_39855,N_38045);
or U40727 (N_40727,N_39458,N_38125);
and U40728 (N_40728,N_38374,N_38418);
nor U40729 (N_40729,N_38856,N_36751);
xor U40730 (N_40730,N_35126,N_38048);
or U40731 (N_40731,N_35038,N_36181);
nand U40732 (N_40732,N_38088,N_37462);
or U40733 (N_40733,N_38129,N_35051);
or U40734 (N_40734,N_38637,N_38799);
xor U40735 (N_40735,N_35489,N_35561);
nor U40736 (N_40736,N_37300,N_39672);
nor U40737 (N_40737,N_39838,N_39800);
and U40738 (N_40738,N_39460,N_37447);
xnor U40739 (N_40739,N_39331,N_36775);
xor U40740 (N_40740,N_39119,N_36529);
and U40741 (N_40741,N_35041,N_39817);
nand U40742 (N_40742,N_36511,N_38109);
or U40743 (N_40743,N_38132,N_37474);
or U40744 (N_40744,N_38321,N_36420);
nand U40745 (N_40745,N_37114,N_39129);
xor U40746 (N_40746,N_39644,N_37875);
xor U40747 (N_40747,N_38685,N_35408);
or U40748 (N_40748,N_35656,N_39859);
or U40749 (N_40749,N_39793,N_39289);
xnor U40750 (N_40750,N_38748,N_38539);
and U40751 (N_40751,N_36273,N_35261);
or U40752 (N_40752,N_39954,N_35763);
xnor U40753 (N_40753,N_36994,N_36849);
nand U40754 (N_40754,N_37496,N_37176);
and U40755 (N_40755,N_35383,N_35692);
nor U40756 (N_40756,N_39768,N_35572);
nand U40757 (N_40757,N_38150,N_39740);
and U40758 (N_40758,N_38382,N_36935);
or U40759 (N_40759,N_36733,N_38477);
nor U40760 (N_40760,N_35779,N_38168);
nand U40761 (N_40761,N_36292,N_35733);
nand U40762 (N_40762,N_37463,N_38481);
xor U40763 (N_40763,N_36972,N_39214);
xor U40764 (N_40764,N_37432,N_36454);
or U40765 (N_40765,N_36462,N_38699);
and U40766 (N_40766,N_36929,N_35092);
or U40767 (N_40767,N_35743,N_37682);
xor U40768 (N_40768,N_36621,N_37369);
xor U40769 (N_40769,N_37205,N_38694);
xnor U40770 (N_40770,N_38272,N_39771);
nor U40771 (N_40771,N_37925,N_36799);
or U40772 (N_40772,N_37279,N_39032);
xor U40773 (N_40773,N_36585,N_39394);
or U40774 (N_40774,N_36025,N_38764);
nor U40775 (N_40775,N_39187,N_36826);
nor U40776 (N_40776,N_35296,N_36465);
or U40777 (N_40777,N_35671,N_38921);
or U40778 (N_40778,N_39503,N_37170);
nor U40779 (N_40779,N_38564,N_37034);
and U40780 (N_40780,N_37207,N_38370);
xor U40781 (N_40781,N_36559,N_36641);
nor U40782 (N_40782,N_36989,N_35845);
nand U40783 (N_40783,N_39595,N_36160);
xor U40784 (N_40784,N_36765,N_37927);
nor U40785 (N_40785,N_38725,N_38200);
and U40786 (N_40786,N_36766,N_36090);
nand U40787 (N_40787,N_35409,N_36527);
nor U40788 (N_40788,N_39157,N_39884);
and U40789 (N_40789,N_39497,N_39937);
or U40790 (N_40790,N_36476,N_39744);
xor U40791 (N_40791,N_37509,N_38751);
xor U40792 (N_40792,N_38876,N_38910);
nand U40793 (N_40793,N_35338,N_39351);
nand U40794 (N_40794,N_38720,N_38185);
nand U40795 (N_40795,N_36904,N_38656);
nor U40796 (N_40796,N_35241,N_39623);
xnor U40797 (N_40797,N_36144,N_36265);
or U40798 (N_40798,N_35621,N_36648);
xor U40799 (N_40799,N_35432,N_39055);
nor U40800 (N_40800,N_38912,N_35933);
nand U40801 (N_40801,N_39889,N_37810);
or U40802 (N_40802,N_39244,N_36294);
or U40803 (N_40803,N_35057,N_38460);
nor U40804 (N_40804,N_36712,N_37994);
xor U40805 (N_40805,N_38445,N_35467);
and U40806 (N_40806,N_38761,N_37821);
nand U40807 (N_40807,N_36819,N_35101);
nand U40808 (N_40808,N_39558,N_35995);
and U40809 (N_40809,N_39150,N_36752);
or U40810 (N_40810,N_37697,N_38633);
xor U40811 (N_40811,N_36596,N_39684);
nor U40812 (N_40812,N_37180,N_35972);
nor U40813 (N_40813,N_39592,N_37988);
or U40814 (N_40814,N_36519,N_39990);
xnor U40815 (N_40815,N_38809,N_36832);
xnor U40816 (N_40816,N_37272,N_38797);
nor U40817 (N_40817,N_37063,N_36990);
nor U40818 (N_40818,N_35956,N_39011);
nor U40819 (N_40819,N_35979,N_37059);
nor U40820 (N_40820,N_35583,N_39084);
nor U40821 (N_40821,N_36778,N_38846);
or U40822 (N_40822,N_38589,N_38559);
and U40823 (N_40823,N_38058,N_39152);
or U40824 (N_40824,N_38793,N_39902);
or U40825 (N_40825,N_36217,N_39378);
or U40826 (N_40826,N_36692,N_37333);
nor U40827 (N_40827,N_35039,N_38870);
nand U40828 (N_40828,N_37057,N_36525);
or U40829 (N_40829,N_39812,N_35998);
nor U40830 (N_40830,N_37132,N_39030);
nand U40831 (N_40831,N_35990,N_35201);
nor U40832 (N_40832,N_36478,N_39846);
nand U40833 (N_40833,N_39952,N_35415);
nor U40834 (N_40834,N_37276,N_35052);
xnor U40835 (N_40835,N_35209,N_39549);
xor U40836 (N_40836,N_37048,N_37389);
or U40837 (N_40837,N_36042,N_37946);
or U40838 (N_40838,N_38353,N_38919);
xor U40839 (N_40839,N_35065,N_38033);
nor U40840 (N_40840,N_37566,N_39781);
or U40841 (N_40841,N_37660,N_39093);
or U40842 (N_40842,N_35484,N_39680);
nand U40843 (N_40843,N_38007,N_39544);
and U40844 (N_40844,N_38854,N_38755);
nor U40845 (N_40845,N_37332,N_35093);
or U40846 (N_40846,N_39927,N_38962);
nor U40847 (N_40847,N_39501,N_35602);
xor U40848 (N_40848,N_39014,N_39410);
and U40849 (N_40849,N_36343,N_36643);
and U40850 (N_40850,N_38861,N_39045);
and U40851 (N_40851,N_36924,N_39792);
nand U40852 (N_40852,N_36916,N_36824);
or U40853 (N_40853,N_35457,N_39586);
xor U40854 (N_40854,N_35570,N_36862);
or U40855 (N_40855,N_37235,N_37551);
nor U40856 (N_40856,N_35899,N_37166);
nand U40857 (N_40857,N_37363,N_37673);
nand U40858 (N_40858,N_35898,N_39707);
and U40859 (N_40859,N_37151,N_35850);
or U40860 (N_40860,N_39913,N_37179);
or U40861 (N_40861,N_38368,N_36967);
and U40862 (N_40862,N_38562,N_36327);
xor U40863 (N_40863,N_39184,N_36810);
or U40864 (N_40864,N_36486,N_35200);
nor U40865 (N_40865,N_36728,N_37646);
nand U40866 (N_40866,N_39456,N_37705);
and U40867 (N_40867,N_37329,N_38742);
xor U40868 (N_40868,N_38900,N_37930);
and U40869 (N_40869,N_35199,N_39661);
xnor U40870 (N_40870,N_36491,N_39585);
nand U40871 (N_40871,N_39295,N_37549);
nand U40872 (N_40872,N_36814,N_39385);
nor U40873 (N_40873,N_38448,N_39308);
and U40874 (N_40874,N_37152,N_39299);
xor U40875 (N_40875,N_35492,N_38709);
nand U40876 (N_40876,N_35577,N_39881);
nand U40877 (N_40877,N_35345,N_37105);
nand U40878 (N_40878,N_37289,N_35701);
or U40879 (N_40879,N_39584,N_36030);
xor U40880 (N_40880,N_39287,N_38537);
or U40881 (N_40881,N_38470,N_39323);
and U40882 (N_40882,N_39268,N_35476);
and U40883 (N_40883,N_37109,N_38204);
xnor U40884 (N_40884,N_37505,N_39322);
nor U40885 (N_40885,N_36238,N_38227);
xor U40886 (N_40886,N_37658,N_37294);
nand U40887 (N_40887,N_39986,N_38320);
and U40888 (N_40888,N_39424,N_37987);
and U40889 (N_40889,N_39970,N_39605);
or U40890 (N_40890,N_36124,N_37773);
or U40891 (N_40891,N_38749,N_39307);
or U40892 (N_40892,N_38057,N_38918);
nand U40893 (N_40893,N_38708,N_36414);
xor U40894 (N_40894,N_36897,N_35555);
nor U40895 (N_40895,N_36747,N_35954);
or U40896 (N_40896,N_35827,N_38003);
xnor U40897 (N_40897,N_37814,N_35960);
and U40898 (N_40898,N_39335,N_35367);
or U40899 (N_40899,N_37804,N_35872);
xnor U40900 (N_40900,N_36497,N_39857);
and U40901 (N_40901,N_38769,N_36798);
nand U40902 (N_40902,N_37343,N_38771);
nor U40903 (N_40903,N_35912,N_38680);
xnor U40904 (N_40904,N_39842,N_35411);
nor U40905 (N_40905,N_39640,N_38212);
and U40906 (N_40906,N_37701,N_36735);
or U40907 (N_40907,N_39823,N_38385);
and U40908 (N_40908,N_37515,N_36681);
xor U40909 (N_40909,N_35560,N_39764);
xor U40910 (N_40910,N_38234,N_36237);
nand U40911 (N_40911,N_38804,N_36315);
and U40912 (N_40912,N_36123,N_35697);
or U40913 (N_40913,N_38659,N_38916);
nand U40914 (N_40914,N_39151,N_35324);
and U40915 (N_40915,N_38386,N_37090);
or U40916 (N_40916,N_36958,N_39370);
and U40917 (N_40917,N_38400,N_38687);
or U40918 (N_40918,N_35111,N_37409);
and U40919 (N_40919,N_37785,N_38319);
nor U40920 (N_40920,N_38603,N_38875);
and U40921 (N_40921,N_35229,N_39353);
and U40922 (N_40922,N_39782,N_35526);
and U40923 (N_40923,N_37623,N_39917);
nand U40924 (N_40924,N_36190,N_39972);
and U40925 (N_40925,N_35322,N_38570);
and U40926 (N_40926,N_36964,N_39095);
and U40927 (N_40927,N_36447,N_36787);
or U40928 (N_40928,N_39484,N_39390);
nor U40929 (N_40929,N_39035,N_39191);
nand U40930 (N_40930,N_39128,N_35354);
and U40931 (N_40931,N_36952,N_37225);
and U40932 (N_40932,N_36568,N_39461);
nand U40933 (N_40933,N_35294,N_35373);
nand U40934 (N_40934,N_35067,N_36919);
or U40935 (N_40935,N_35147,N_37459);
nand U40936 (N_40936,N_35502,N_37172);
nor U40937 (N_40937,N_35082,N_36722);
xnor U40938 (N_40938,N_37212,N_39959);
nand U40939 (N_40939,N_37630,N_37481);
xor U40940 (N_40940,N_35363,N_38220);
xor U40941 (N_40941,N_36900,N_35404);
nand U40942 (N_40942,N_35611,N_39445);
nand U40943 (N_40943,N_39822,N_36657);
nor U40944 (N_40944,N_36323,N_39848);
nand U40945 (N_40945,N_38276,N_35667);
nand U40946 (N_40946,N_39138,N_38199);
and U40947 (N_40947,N_35564,N_36431);
nor U40948 (N_40948,N_39758,N_39864);
nand U40949 (N_40949,N_39625,N_37214);
xnor U40950 (N_40950,N_35552,N_39238);
xor U40951 (N_40951,N_39328,N_36433);
nand U40952 (N_40952,N_39710,N_37593);
or U40953 (N_40953,N_37620,N_35789);
and U40954 (N_40954,N_38054,N_38036);
nor U40955 (N_40955,N_39659,N_37659);
nor U40956 (N_40956,N_35958,N_36620);
or U40957 (N_40957,N_36795,N_36984);
nor U40958 (N_40958,N_37527,N_35962);
xor U40959 (N_40959,N_37845,N_36721);
or U40960 (N_40960,N_37157,N_36851);
and U40961 (N_40961,N_37139,N_39968);
nor U40962 (N_40962,N_39975,N_38084);
nand U40963 (N_40963,N_38777,N_37560);
nor U40964 (N_40964,N_37317,N_37239);
or U40965 (N_40965,N_38224,N_36686);
xnor U40966 (N_40966,N_37951,N_38760);
xor U40967 (N_40967,N_38426,N_36126);
nor U40968 (N_40968,N_36398,N_36569);
nand U40969 (N_40969,N_36346,N_37450);
and U40970 (N_40970,N_39329,N_37142);
nand U40971 (N_40971,N_38138,N_39695);
xnor U40972 (N_40972,N_35678,N_39259);
nand U40973 (N_40973,N_39925,N_36882);
and U40974 (N_40974,N_36286,N_37309);
xor U40975 (N_40975,N_35307,N_38114);
or U40976 (N_40976,N_39945,N_37080);
xor U40977 (N_40977,N_36151,N_35848);
nand U40978 (N_40978,N_38597,N_37092);
nand U40979 (N_40979,N_39529,N_36668);
or U40980 (N_40980,N_38787,N_35273);
xnor U40981 (N_40981,N_36961,N_38624);
nand U40982 (N_40982,N_37633,N_36357);
nor U40983 (N_40983,N_39033,N_37192);
nor U40984 (N_40984,N_35940,N_37178);
xor U40985 (N_40985,N_38213,N_39947);
nand U40986 (N_40986,N_37108,N_39992);
nor U40987 (N_40987,N_36646,N_39624);
nand U40988 (N_40988,N_36351,N_38196);
nand U40989 (N_40989,N_39107,N_35143);
nor U40990 (N_40990,N_36868,N_36377);
nand U40991 (N_40991,N_35769,N_35072);
nand U40992 (N_40992,N_39383,N_39573);
nand U40993 (N_40993,N_35724,N_35066);
and U40994 (N_40994,N_38294,N_35330);
nand U40995 (N_40995,N_39448,N_35349);
nor U40996 (N_40996,N_35482,N_38179);
nor U40997 (N_40997,N_38733,N_38631);
or U40998 (N_40998,N_36557,N_37538);
xnor U40999 (N_40999,N_36234,N_39098);
or U41000 (N_41000,N_39403,N_38066);
nor U41001 (N_41001,N_39969,N_35626);
nand U41002 (N_41002,N_36767,N_39716);
nand U41003 (N_41003,N_36638,N_37837);
xnor U41004 (N_41004,N_38614,N_39405);
xnor U41005 (N_41005,N_35389,N_38106);
xor U41006 (N_41006,N_35737,N_39923);
nor U41007 (N_41007,N_39450,N_37029);
nor U41008 (N_41008,N_39306,N_39786);
nor U41009 (N_41009,N_38420,N_37433);
nand U41010 (N_41010,N_36437,N_36618);
nand U41011 (N_41011,N_37770,N_36777);
xnor U41012 (N_41012,N_37907,N_38641);
xor U41013 (N_41013,N_37957,N_35485);
or U41014 (N_41014,N_38850,N_35856);
nand U41015 (N_41015,N_35781,N_36700);
nand U41016 (N_41016,N_36831,N_39553);
and U41017 (N_41017,N_38857,N_36158);
and U41018 (N_41018,N_39841,N_37078);
nand U41019 (N_41019,N_39265,N_37908);
and U41020 (N_41020,N_39221,N_36250);
and U41021 (N_41021,N_39717,N_37574);
nand U41022 (N_41022,N_37303,N_37711);
nand U41023 (N_41023,N_35390,N_39813);
nor U41024 (N_41024,N_36106,N_35165);
nand U41025 (N_41025,N_36741,N_39077);
and U41026 (N_41026,N_35184,N_35646);
or U41027 (N_41027,N_36704,N_35327);
or U41028 (N_41028,N_38155,N_39155);
or U41029 (N_41029,N_36516,N_37259);
and U41030 (N_41030,N_39234,N_36080);
and U41031 (N_41031,N_36820,N_37315);
xor U41032 (N_41032,N_38343,N_39714);
and U41033 (N_41033,N_39938,N_36993);
and U41034 (N_41034,N_38077,N_37568);
nand U41035 (N_41035,N_38789,N_38717);
and U41036 (N_41036,N_37256,N_38627);
nand U41037 (N_41037,N_37860,N_37863);
and U41038 (N_41038,N_36477,N_37341);
xor U41039 (N_41039,N_37671,N_36416);
and U41040 (N_41040,N_37557,N_37385);
or U41041 (N_41041,N_36226,N_39267);
and U41042 (N_41042,N_35177,N_39981);
nor U41043 (N_41043,N_38849,N_35797);
nand U41044 (N_41044,N_38642,N_39632);
or U41045 (N_41045,N_39412,N_37146);
xnor U41046 (N_41046,N_37216,N_35601);
or U41047 (N_41047,N_36883,N_38566);
nor U41048 (N_41048,N_38521,N_39088);
nand U41049 (N_41049,N_36891,N_38901);
or U41050 (N_41050,N_36426,N_37934);
xnor U41051 (N_41051,N_39449,N_36804);
xor U41052 (N_41052,N_35786,N_36944);
xnor U41053 (N_41053,N_39473,N_37779);
nor U41054 (N_41054,N_38303,N_38119);
nand U41055 (N_41055,N_37351,N_39491);
nor U41056 (N_41056,N_36833,N_38736);
nor U41057 (N_41057,N_39480,N_37532);
nand U41058 (N_41058,N_35764,N_38848);
or U41059 (N_41059,N_39174,N_39219);
nand U41060 (N_41060,N_36120,N_37222);
xor U41061 (N_41061,N_35403,N_39646);
nor U41062 (N_41062,N_35892,N_39391);
or U41063 (N_41063,N_36402,N_38071);
xor U41064 (N_41064,N_39134,N_39406);
or U41065 (N_41065,N_37664,N_37370);
or U41066 (N_41066,N_39946,N_37978);
nor U41067 (N_41067,N_37594,N_35799);
nand U41068 (N_41068,N_38503,N_35973);
or U41069 (N_41069,N_36312,N_37218);
xnor U41070 (N_41070,N_37878,N_38405);
nor U41071 (N_41071,N_39243,N_35236);
and U41072 (N_41072,N_38544,N_37147);
and U41073 (N_41073,N_36445,N_36571);
nor U41074 (N_41074,N_39357,N_36687);
or U41075 (N_41075,N_36760,N_37961);
nor U41076 (N_41076,N_37282,N_37190);
nand U41077 (N_41077,N_35766,N_38291);
nand U41078 (N_41078,N_38533,N_39561);
and U41079 (N_41079,N_35374,N_39066);
and U41080 (N_41080,N_39100,N_37189);
or U41081 (N_41081,N_37305,N_36791);
nor U41082 (N_41082,N_39825,N_38465);
or U41083 (N_41083,N_35193,N_35796);
xor U41084 (N_41084,N_37082,N_36308);
or U41085 (N_41085,N_38333,N_39609);
nor U41086 (N_41086,N_39454,N_38162);
nand U41087 (N_41087,N_39421,N_39706);
or U41088 (N_41088,N_37168,N_35882);
and U41089 (N_41089,N_38881,N_35006);
nand U41090 (N_41090,N_35112,N_36876);
nor U41091 (N_41091,N_38431,N_38652);
and U41092 (N_41092,N_37887,N_37607);
nor U41093 (N_41093,N_38214,N_39619);
nand U41094 (N_41094,N_39355,N_35268);
and U41095 (N_41095,N_35336,N_35927);
and U41096 (N_41096,N_36632,N_36874);
nand U41097 (N_41097,N_37420,N_36056);
and U41098 (N_41098,N_38175,N_35466);
xnor U41099 (N_41099,N_37928,N_36732);
xnor U41100 (N_41100,N_38043,N_37100);
and U41101 (N_41101,N_37393,N_35119);
nand U41102 (N_41102,N_37895,N_36372);
nor U41103 (N_41103,N_38819,N_37228);
or U41104 (N_41104,N_35441,N_39897);
nor U41105 (N_41105,N_36748,N_36580);
or U41106 (N_41106,N_35168,N_38047);
or U41107 (N_41107,N_36101,N_39002);
nand U41108 (N_41108,N_35255,N_36962);
nand U41109 (N_41109,N_38173,N_39934);
or U41110 (N_41110,N_39833,N_36669);
and U41111 (N_41111,N_39749,N_37539);
nor U41112 (N_41112,N_36031,N_38085);
nor U41113 (N_41113,N_37232,N_35089);
nor U41114 (N_41114,N_38198,N_35930);
nand U41115 (N_41115,N_36943,N_39388);
xnor U41116 (N_41116,N_38555,N_37489);
xor U41117 (N_41117,N_37933,N_39490);
nor U41118 (N_41118,N_39895,N_35429);
or U41119 (N_41119,N_38763,N_35928);
nor U41120 (N_41120,N_37552,N_37233);
and U41121 (N_41121,N_37230,N_35104);
nand U41122 (N_41122,N_37831,N_35974);
or U41123 (N_41123,N_39345,N_35606);
and U41124 (N_41124,N_36127,N_39013);
xor U41125 (N_41125,N_37812,N_38785);
or U41126 (N_41126,N_36468,N_39780);
or U41127 (N_41127,N_35377,N_37350);
and U41128 (N_41128,N_36574,N_35443);
xnor U41129 (N_41129,N_39776,N_36187);
and U41130 (N_41130,N_38806,N_38723);
nand U41131 (N_41131,N_38573,N_39260);
or U41132 (N_41132,N_38971,N_37191);
nor U41133 (N_41133,N_39816,N_35477);
xnor U41134 (N_41134,N_36466,N_37893);
nand U41135 (N_41135,N_37265,N_35187);
xnor U41136 (N_41136,N_36229,N_37601);
xor U41137 (N_41137,N_36725,N_38998);
or U41138 (N_41138,N_37503,N_37873);
nor U41139 (N_41139,N_36176,N_36378);
or U41140 (N_41140,N_36490,N_35018);
or U41141 (N_41141,N_37913,N_39526);
or U41142 (N_41142,N_39508,N_36021);
nor U41143 (N_41143,N_36734,N_36259);
nor U41144 (N_41144,N_39851,N_38163);
nand U41145 (N_41145,N_37661,N_38702);
xor U41146 (N_41146,N_36594,N_36442);
xor U41147 (N_41147,N_39297,N_38131);
or U41148 (N_41148,N_35695,N_36506);
nand U41149 (N_41149,N_36565,N_37624);
nor U41150 (N_41150,N_38042,N_38943);
xor U41151 (N_41151,N_38548,N_35160);
or U41152 (N_41152,N_38457,N_37441);
nor U41153 (N_41153,N_35944,N_35859);
or U41154 (N_41154,N_38247,N_35537);
and U41155 (N_41155,N_36789,N_37345);
xnor U41156 (N_41156,N_39425,N_35853);
or U41157 (N_41157,N_39105,N_36998);
and U41158 (N_41158,N_35887,N_35015);
nor U41159 (N_41159,N_38698,N_38255);
xor U41160 (N_41160,N_35735,N_39797);
nor U41161 (N_41161,N_36689,N_38815);
and U41162 (N_41162,N_36040,N_36313);
nor U41163 (N_41163,N_37615,N_38524);
nor U41164 (N_41164,N_37465,N_35911);
or U41165 (N_41165,N_36985,N_39702);
and U41166 (N_41166,N_38563,N_38149);
and U41167 (N_41167,N_35915,N_37275);
or U41168 (N_41168,N_38166,N_37936);
and U41169 (N_41169,N_35242,N_37577);
nand U41170 (N_41170,N_36991,N_36369);
and U41171 (N_41171,N_37768,N_35913);
and U41172 (N_41172,N_38677,N_39283);
nor U41173 (N_41173,N_36724,N_35804);
nor U41174 (N_41174,N_37580,N_37297);
nor U41175 (N_41175,N_35655,N_39468);
nand U41176 (N_41176,N_35610,N_38858);
or U41177 (N_41177,N_36306,N_38356);
xnor U41178 (N_41178,N_35310,N_37529);
nand U41179 (N_41179,N_35295,N_35840);
nor U41180 (N_41180,N_36854,N_35328);
and U41181 (N_41181,N_36846,N_35257);
or U41182 (N_41182,N_38696,N_36133);
or U41183 (N_41183,N_39477,N_35605);
or U41184 (N_41184,N_36499,N_35527);
nor U41185 (N_41185,N_36103,N_36493);
nor U41186 (N_41186,N_37392,N_37145);
nor U41187 (N_41187,N_38442,N_37182);
nand U41188 (N_41188,N_37234,N_36655);
and U41189 (N_41189,N_39891,N_35202);
and U41190 (N_41190,N_35830,N_38233);
nor U41191 (N_41191,N_35687,N_38103);
and U41192 (N_41192,N_39242,N_37584);
nand U41193 (N_41193,N_39596,N_39222);
nand U41194 (N_41194,N_35821,N_36694);
xnor U41195 (N_41195,N_38711,N_35033);
and U41196 (N_41196,N_39809,N_37417);
nor U41197 (N_41197,N_37867,N_38978);
xor U41198 (N_41198,N_36940,N_36542);
nand U41199 (N_41199,N_37842,N_38230);
or U41200 (N_41200,N_36052,N_35454);
and U41201 (N_41201,N_39853,N_36383);
xnor U41202 (N_41202,N_36873,N_38206);
nand U41203 (N_41203,N_38349,N_37236);
nor U41204 (N_41204,N_36693,N_36367);
nor U41205 (N_41205,N_35580,N_35188);
nor U41206 (N_41206,N_35267,N_39806);
nor U41207 (N_41207,N_37995,N_39550);
or U41208 (N_41208,N_35448,N_38489);
nand U41209 (N_41209,N_39757,N_39162);
or U41210 (N_41210,N_36869,N_35047);
and U41211 (N_41211,N_37782,N_35718);
nand U41212 (N_41212,N_37181,N_38396);
and U41213 (N_41213,N_38676,N_37278);
nor U41214 (N_41214,N_36770,N_36301);
nor U41215 (N_41215,N_35120,N_38323);
or U41216 (N_41216,N_38450,N_36352);
xnor U41217 (N_41217,N_37534,N_37188);
and U41218 (N_41218,N_37336,N_38690);
or U41219 (N_41219,N_38078,N_35013);
nand U41220 (N_41220,N_35551,N_36149);
xor U41221 (N_41221,N_39269,N_39029);
nor U41222 (N_41222,N_38113,N_39404);
nor U41223 (N_41223,N_37579,N_35647);
and U41224 (N_41224,N_36606,N_39581);
nor U41225 (N_41225,N_38843,N_38169);
nor U41226 (N_41226,N_37111,N_39252);
nand U41227 (N_41227,N_37983,N_38986);
and U41228 (N_41228,N_35054,N_39476);
nor U41229 (N_41229,N_36019,N_39389);
xor U41230 (N_41230,N_35546,N_37542);
xor U41231 (N_41231,N_38377,N_36438);
xor U41232 (N_41232,N_39136,N_37896);
or U41233 (N_41233,N_36393,N_35563);
or U41234 (N_41234,N_38831,N_38222);
or U41235 (N_41235,N_37710,N_35554);
xor U41236 (N_41236,N_39539,N_39144);
and U41237 (N_41237,N_38593,N_37076);
nand U41238 (N_41238,N_37113,N_35628);
nand U41239 (N_41239,N_38632,N_35504);
nor U41240 (N_41240,N_39399,N_37784);
or U41241 (N_41241,N_38947,N_37776);
nor U41242 (N_41242,N_38348,N_37583);
nor U41243 (N_41243,N_35007,N_35624);
or U41244 (N_41244,N_39538,N_38556);
and U41245 (N_41245,N_38989,N_39856);
and U41246 (N_41246,N_39041,N_36094);
xnor U41247 (N_41247,N_37062,N_37502);
xor U41248 (N_41248,N_37722,N_39409);
and U41249 (N_41249,N_38507,N_35396);
xnor U41250 (N_41250,N_35773,N_39397);
nor U41251 (N_41251,N_35081,N_35965);
xor U41252 (N_41252,N_36330,N_38373);
nand U41253 (N_41253,N_39001,N_35115);
nand U41254 (N_41254,N_36244,N_36471);
and U41255 (N_41255,N_39593,N_39652);
and U41256 (N_41256,N_39614,N_37375);
nand U41257 (N_41257,N_38952,N_35208);
nor U41258 (N_41258,N_37285,N_35883);
xor U41259 (N_41259,N_37384,N_36871);
nand U41260 (N_41260,N_36889,N_35792);
and U41261 (N_41261,N_35604,N_39498);
nor U41262 (N_41262,N_35581,N_36956);
or U41263 (N_41263,N_39311,N_37199);
and U41264 (N_41264,N_38105,N_38360);
and U41265 (N_41265,N_36289,N_36492);
and U41266 (N_41266,N_35922,N_37467);
nor U41267 (N_41267,N_35652,N_39984);
and U41268 (N_41268,N_39724,N_35800);
or U41269 (N_41269,N_35076,N_39240);
and U41270 (N_41270,N_39081,N_37049);
xor U41271 (N_41271,N_39063,N_37537);
xor U41272 (N_41272,N_37293,N_35098);
nand U41273 (N_41273,N_37976,N_39346);
or U41274 (N_41274,N_37257,N_39979);
xor U41275 (N_41275,N_37041,N_36859);
or U41276 (N_41276,N_36960,N_37738);
or U41277 (N_41277,N_36903,N_38682);
and U41278 (N_41278,N_36509,N_39705);
or U41279 (N_41279,N_37084,N_38006);
and U41280 (N_41280,N_36806,N_37117);
nor U41281 (N_41281,N_37700,N_35931);
or U41282 (N_41282,N_38146,N_38852);
and U41283 (N_41283,N_38492,N_37075);
or U41284 (N_41284,N_37663,N_39446);
or U41285 (N_41285,N_39270,N_38959);
or U41286 (N_41286,N_38651,N_39365);
or U41287 (N_41287,N_38812,N_35239);
nand U41288 (N_41288,N_36002,N_38824);
xnor U41289 (N_41289,N_37899,N_38380);
and U41290 (N_41290,N_35009,N_37901);
or U41291 (N_41291,N_35679,N_35750);
xnor U41292 (N_41292,N_37528,N_37605);
and U41293 (N_41293,N_36925,N_38807);
nand U41294 (N_41294,N_36887,N_35130);
or U41295 (N_41295,N_38369,N_39882);
nor U41296 (N_41296,N_37774,N_37395);
xnor U41297 (N_41297,N_36228,N_35231);
or U41298 (N_41298,N_39935,N_36945);
and U41299 (N_41299,N_37986,N_37497);
and U41300 (N_41300,N_37227,N_39904);
nand U41301 (N_41301,N_36645,N_38096);
nor U41302 (N_41302,N_35034,N_38688);
or U41303 (N_41303,N_39453,N_35246);
nand U41304 (N_41304,N_37372,N_38599);
nor U41305 (N_41305,N_39317,N_39074);
and U41306 (N_41306,N_35036,N_37786);
xnor U41307 (N_41307,N_36375,N_37725);
nand U41308 (N_41308,N_35615,N_36615);
nor U41309 (N_41309,N_37992,N_38903);
and U41310 (N_41310,N_38152,N_36299);
and U41311 (N_41311,N_35732,N_35937);
nor U41312 (N_41312,N_37469,N_35398);
xor U41313 (N_41313,N_35353,N_37999);
xor U41314 (N_41314,N_35281,N_37849);
nor U41315 (N_41315,N_35303,N_36982);
nand U41316 (N_41316,N_38860,N_37931);
or U41317 (N_41317,N_35810,N_36575);
nand U41318 (N_41318,N_39247,N_38650);
or U41319 (N_41319,N_36547,N_35029);
and U41320 (N_41320,N_39685,N_36524);
and U41321 (N_41321,N_37677,N_36449);
and U41322 (N_41322,N_36923,N_37368);
xor U41323 (N_41323,N_36348,N_36349);
xor U41324 (N_41324,N_36609,N_36783);
nand U41325 (N_41325,N_37853,N_37253);
or U41326 (N_41326,N_39218,N_39948);
nor U41327 (N_41327,N_39564,N_38285);
and U41328 (N_41328,N_37073,N_37026);
and U41329 (N_41329,N_38134,N_38123);
and U41330 (N_41330,N_36549,N_35271);
nand U41331 (N_41331,N_35869,N_35174);
and U41332 (N_41332,N_36572,N_36360);
nand U41333 (N_41333,N_35617,N_36888);
nand U41334 (N_41334,N_38346,N_35220);
and U41335 (N_41335,N_36866,N_36498);
and U41336 (N_41336,N_38508,N_35381);
nor U41337 (N_41337,N_38016,N_38347);
nand U41338 (N_41338,N_37653,N_35721);
nor U41339 (N_41339,N_36811,N_37337);
or U41340 (N_41340,N_35180,N_38143);
or U41341 (N_41341,N_38757,N_37006);
xor U41342 (N_41342,N_39258,N_35410);
nor U41343 (N_41343,N_37858,N_37952);
nor U41344 (N_41344,N_38412,N_35550);
and U41345 (N_41345,N_38983,N_36800);
nor U41346 (N_41346,N_39109,N_35993);
and U41347 (N_41347,N_39154,N_39127);
nor U41348 (N_41348,N_35230,N_36311);
xnor U41349 (N_41349,N_38842,N_39006);
and U41350 (N_41350,N_36614,N_39133);
nand U41351 (N_41351,N_38520,N_39513);
nand U41352 (N_41352,N_35450,N_37558);
nor U41353 (N_41353,N_36761,N_39905);
or U41354 (N_41354,N_36170,N_39815);
and U41355 (N_41355,N_35575,N_38948);
nor U41356 (N_41356,N_36785,N_39943);
and U41357 (N_41357,N_36189,N_35133);
nor U41358 (N_41358,N_36496,N_39799);
nand U41359 (N_41359,N_36628,N_38280);
or U41360 (N_41360,N_39622,N_39836);
nand U41361 (N_41361,N_35042,N_37820);
or U41362 (N_41362,N_37667,N_37331);
nor U41363 (N_41363,N_38040,N_39419);
xor U41364 (N_41364,N_38145,N_39689);
nand U41365 (N_41365,N_39086,N_37636);
nand U41366 (N_41366,N_39795,N_39522);
and U41367 (N_41367,N_38219,N_38925);
nor U41368 (N_41368,N_36087,N_38099);
nor U41369 (N_41369,N_36521,N_38273);
nand U41370 (N_41370,N_38124,N_38891);
or U41371 (N_41371,N_35442,N_39950);
nor U41372 (N_41372,N_37859,N_36038);
or U41373 (N_41373,N_36475,N_38897);
xor U41374 (N_41374,N_39915,N_38938);
xor U41375 (N_41375,N_37195,N_39530);
or U41376 (N_41376,N_35495,N_37405);
xor U41377 (N_41377,N_38596,N_35021);
nor U41378 (N_41378,N_36248,N_35260);
xnor U41379 (N_41379,N_38496,N_35714);
nor U41380 (N_41380,N_39146,N_39634);
xnor U41381 (N_41381,N_39918,N_37585);
and U41382 (N_41382,N_39944,N_37743);
or U41383 (N_41383,N_37413,N_37487);
nand U41384 (N_41384,N_38776,N_37204);
nand U41385 (N_41385,N_37094,N_36155);
and U41386 (N_41386,N_36018,N_35110);
and U41387 (N_41387,N_35161,N_37868);
nand U41388 (N_41388,N_35393,N_38413);
xor U41389 (N_41389,N_39831,N_36779);
xor U41390 (N_41390,N_36842,N_36218);
or U41391 (N_41391,N_35213,N_38712);
nor U41392 (N_41392,N_38086,N_39987);
nand U41393 (N_41393,N_37183,N_37761);
nand U41394 (N_41394,N_35961,N_39649);
nand U41395 (N_41395,N_36586,N_36104);
xor U41396 (N_41396,N_37522,N_36284);
nor U41397 (N_41397,N_37817,N_38823);
nand U41398 (N_41398,N_39506,N_39698);
nand U41399 (N_41399,N_36354,N_38068);
or U41400 (N_41400,N_35480,N_36560);
xor U41401 (N_41401,N_36860,N_38083);
nor U41402 (N_41402,N_37572,N_37130);
or U41403 (N_41403,N_37066,N_36540);
and U41404 (N_41404,N_39532,N_35953);
nor U41405 (N_41405,N_38052,N_37438);
nor U41406 (N_41406,N_37058,N_37769);
nand U41407 (N_41407,N_37980,N_39965);
nand U41408 (N_41408,N_37556,N_39801);
and U41409 (N_41409,N_36257,N_37377);
or U41410 (N_41410,N_37524,N_38337);
nor U41411 (N_41411,N_39756,N_35412);
or U41412 (N_41412,N_35195,N_36361);
or U41413 (N_41413,N_38228,N_39290);
nand U41414 (N_41414,N_39687,N_35846);
and U41415 (N_41415,N_36867,N_36239);
nor U41416 (N_41416,N_39472,N_37254);
xor U41417 (N_41417,N_39177,N_39464);
nor U41418 (N_41418,N_39075,N_36667);
nand U41419 (N_41419,N_38529,N_35863);
xnor U41420 (N_41420,N_39535,N_39414);
and U41421 (N_41421,N_39054,N_35820);
xnor U41422 (N_41422,N_36677,N_36032);
nand U41423 (N_41423,N_35873,N_35536);
nor U41424 (N_41424,N_35980,N_37150);
or U41425 (N_41425,N_39667,N_38506);
or U41426 (N_41426,N_39886,N_37854);
or U41427 (N_41427,N_39199,N_38636);
nand U41428 (N_41428,N_37883,N_38697);
and U41429 (N_41429,N_36410,N_35243);
and U41430 (N_41430,N_36109,N_37482);
or U41431 (N_41431,N_37838,N_38464);
nor U41432 (N_41432,N_39395,N_35530);
and U41433 (N_41433,N_38087,N_35430);
and U41434 (N_41434,N_36046,N_37269);
or U41435 (N_41435,N_39504,N_37793);
or U41436 (N_41436,N_39202,N_37811);
or U41437 (N_41437,N_37271,N_36054);
or U41438 (N_41438,N_35885,N_35776);
and U41439 (N_41439,N_35129,N_36675);
nand U41440 (N_41440,N_39677,N_36803);
nand U41441 (N_41441,N_37127,N_35891);
xnor U41442 (N_41442,N_38192,N_36768);
or U41443 (N_41443,N_39254,N_37408);
nor U41444 (N_41444,N_36905,N_37458);
or U41445 (N_41445,N_37136,N_38922);
nor U41446 (N_41446,N_39951,N_36291);
and U41447 (N_41447,N_39049,N_39333);
nor U41448 (N_41448,N_39362,N_38140);
xnor U41449 (N_41449,N_35136,N_36464);
nand U41450 (N_41450,N_37308,N_39195);
nor U41451 (N_41451,N_36813,N_39852);
and U41452 (N_41452,N_39273,N_39583);
nand U41453 (N_41453,N_36997,N_39766);
or U41454 (N_41454,N_37668,N_36635);
and U41455 (N_41455,N_37533,N_38525);
and U41456 (N_41456,N_38851,N_39887);
xnor U41457 (N_41457,N_35070,N_38988);
nor U41458 (N_41458,N_36353,N_37067);
nor U41459 (N_41459,N_35173,N_39545);
or U41460 (N_41460,N_36688,N_35473);
nor U41461 (N_41461,N_36399,N_38354);
nor U41462 (N_41462,N_38645,N_35486);
nor U41463 (N_41463,N_37213,N_39515);
nand U41464 (N_41464,N_35921,N_37167);
or U41465 (N_41465,N_36044,N_36373);
nand U41466 (N_41466,N_37635,N_36578);
nor U41467 (N_41467,N_35030,N_38788);
or U41468 (N_41468,N_38193,N_38190);
xor U41469 (N_41469,N_36364,N_35002);
or U41470 (N_41470,N_39336,N_36980);
and U41471 (N_41471,N_39840,N_39475);
nand U41472 (N_41472,N_38681,N_39602);
or U41473 (N_41473,N_37622,N_35386);
or U41474 (N_41474,N_37119,N_38541);
or U41475 (N_41475,N_38311,N_39212);
or U41476 (N_41476,N_35394,N_37945);
nor U41477 (N_41477,N_37295,N_36877);
xor U41478 (N_41478,N_39870,N_35685);
nor U41479 (N_41479,N_37898,N_36255);
nor U41480 (N_41480,N_39147,N_37306);
or U41481 (N_41481,N_39755,N_39785);
nor U41482 (N_41482,N_37720,N_39118);
xnor U41483 (N_41483,N_37805,N_36141);
and U41484 (N_41484,N_36537,N_38700);
and U41485 (N_41485,N_35469,N_36227);
or U41486 (N_41486,N_35279,N_36823);
and U41487 (N_41487,N_35657,N_37000);
and U41488 (N_41488,N_39999,N_36222);
or U41489 (N_41489,N_37122,N_38987);
and U41490 (N_41490,N_39334,N_36271);
or U41491 (N_41491,N_37891,N_39193);
nand U41492 (N_41492,N_37950,N_37638);
nand U41493 (N_41493,N_37626,N_36166);
or U41494 (N_41494,N_37846,N_39660);
xor U41495 (N_41495,N_35382,N_38662);
xor U41496 (N_41496,N_36082,N_38835);
and U41497 (N_41497,N_38361,N_39568);
xnor U41498 (N_41498,N_37427,N_39808);
or U41499 (N_41499,N_37906,N_36329);
nand U41500 (N_41500,N_35315,N_36508);
nor U41501 (N_41501,N_38801,N_36975);
and U41502 (N_41502,N_36213,N_37360);
and U41503 (N_41503,N_35672,N_37851);
xnor U41504 (N_41504,N_38830,N_39340);
nor U41505 (N_41505,N_38002,N_39683);
nand U41506 (N_41506,N_36595,N_36531);
nand U41507 (N_41507,N_37425,N_37466);
nand U41508 (N_41508,N_39375,N_35717);
nand U41509 (N_41509,N_35829,N_38612);
xor U41510 (N_41510,N_38740,N_37592);
xor U41511 (N_41511,N_35434,N_36647);
nor U41512 (N_41512,N_37744,N_36830);
nor U41513 (N_41513,N_36297,N_35053);
or U41514 (N_41514,N_38678,N_37991);
and U41515 (N_41515,N_37047,N_37941);
nor U41516 (N_41516,N_39213,N_35090);
or U41517 (N_41517,N_36481,N_39310);
nor U41518 (N_41518,N_38803,N_38606);
and U41519 (N_41519,N_39271,N_37116);
and U41520 (N_41520,N_39807,N_39582);
xor U41521 (N_41521,N_36715,N_36562);
or U41522 (N_41522,N_37072,N_38330);
and U41523 (N_41523,N_37972,N_36865);
nand U41524 (N_41524,N_38339,N_38557);
or U41525 (N_41525,N_38913,N_37096);
nor U41526 (N_41526,N_37604,N_36838);
nand U41527 (N_41527,N_35976,N_36034);
nand U41528 (N_41528,N_36576,N_37847);
or U41529 (N_41529,N_35017,N_39611);
or U41530 (N_41530,N_39141,N_36129);
and U41531 (N_41531,N_39111,N_35730);
and U41532 (N_41532,N_39778,N_36714);
nand U41533 (N_41533,N_38778,N_35512);
nand U41534 (N_41534,N_36335,N_37359);
xor U41535 (N_41535,N_37155,N_37516);
or U41536 (N_41536,N_39700,N_37013);
and U41537 (N_41537,N_37479,N_35329);
and U41538 (N_41538,N_36719,N_37177);
nor U41539 (N_41539,N_38288,N_38030);
and U41540 (N_41540,N_35475,N_39296);
and U41541 (N_41541,N_38065,N_37678);
xnor U41542 (N_41542,N_39120,N_36121);
nand U41543 (N_41543,N_39657,N_35050);
and U41544 (N_41544,N_39977,N_39524);
and U41545 (N_41545,N_39429,N_37030);
nand U41546 (N_41546,N_39216,N_37009);
xor U41547 (N_41547,N_35152,N_37313);
and U41548 (N_41548,N_37429,N_36197);
nand U41549 (N_41549,N_35914,N_38005);
xnor U41550 (N_41550,N_39312,N_39058);
or U41551 (N_41551,N_35008,N_37713);
xor U41552 (N_41552,N_35314,N_38364);
or U41553 (N_41553,N_38161,N_38994);
nand U41554 (N_41554,N_39418,N_36651);
nand U41555 (N_41555,N_35414,N_38056);
nand U41556 (N_41556,N_37455,N_38183);
nor U41557 (N_41557,N_38027,N_36977);
or U41558 (N_41558,N_38893,N_39621);
nand U41559 (N_41559,N_36344,N_39451);
or U41560 (N_41560,N_36554,N_37140);
nor U41561 (N_41561,N_39376,N_35908);
nand U41562 (N_41562,N_35245,N_39783);
or U41563 (N_41563,N_38625,N_39482);
and U41564 (N_41564,N_39183,N_38037);
nand U41565 (N_41565,N_36333,N_39767);
nand U41566 (N_41566,N_37937,N_37809);
or U41567 (N_41567,N_39065,N_39139);
nand U41568 (N_41568,N_35637,N_36543);
nand U41569 (N_41569,N_37310,N_37578);
nand U41570 (N_41570,N_37518,N_39528);
nor U41571 (N_41571,N_36047,N_35525);
xnor U41572 (N_41572,N_39278,N_38394);
nand U41573 (N_41573,N_36968,N_36757);
nand U41574 (N_41574,N_36482,N_35917);
or U41575 (N_41575,N_36986,N_39487);
nor U41576 (N_41576,N_39861,N_37488);
nand U41577 (N_41577,N_37752,N_36374);
nand U41578 (N_41578,N_39988,N_37460);
and U41579 (N_41579,N_39366,N_35107);
xnor U41580 (N_41580,N_38461,N_37918);
and U41581 (N_41581,N_38940,N_35590);
or U41582 (N_41582,N_39903,N_35419);
xnor U41583 (N_41583,N_35557,N_39279);
and U41584 (N_41584,N_35793,N_38867);
xor U41585 (N_41585,N_35842,N_39958);
or U41586 (N_41586,N_37696,N_39046);
or U41587 (N_41587,N_37143,N_36139);
xor U41588 (N_41588,N_35985,N_39026);
or U41589 (N_41589,N_36544,N_36927);
nand U41590 (N_41590,N_35597,N_38174);
xor U41591 (N_41591,N_35496,N_37866);
xnor U41592 (N_41592,N_36713,N_35049);
or U41593 (N_41593,N_35431,N_35080);
nand U41594 (N_41594,N_38139,N_39262);
and U41595 (N_41595,N_39089,N_36418);
nor U41596 (N_41596,N_37184,N_38176);
and U41597 (N_41597,N_35934,N_37535);
nor U41598 (N_41598,N_37864,N_39639);
or U41599 (N_41599,N_37098,N_36178);
nor U41600 (N_41600,N_36703,N_38411);
or U41601 (N_41601,N_35582,N_36604);
or U41602 (N_41602,N_37917,N_38883);
nand U41603 (N_41603,N_39578,N_37353);
xnor U41604 (N_41604,N_36450,N_37586);
and U41605 (N_41605,N_38721,N_39607);
xor U41606 (N_41606,N_37511,N_37571);
nor U41607 (N_41607,N_37412,N_39900);
and U41608 (N_41608,N_35272,N_37565);
nor U41609 (N_41609,N_37598,N_39627);
nand U41610 (N_41610,N_39431,N_38404);
or U41611 (N_41611,N_35895,N_38907);
nor U41612 (N_41612,N_35627,N_35731);
or U41613 (N_41613,N_39470,N_39126);
nor U41614 (N_41614,N_36899,N_38497);
and U41615 (N_41615,N_35897,N_38944);
nand U41616 (N_41616,N_36974,N_35689);
nand U41617 (N_41617,N_38578,N_36118);
and U41618 (N_41618,N_37270,N_39779);
or U41619 (N_41619,N_36650,N_38522);
nand U41620 (N_41620,N_35746,N_36794);
and U41621 (N_41621,N_36901,N_37919);
or U41622 (N_41622,N_35696,N_35105);
xnor U41623 (N_41623,N_35287,N_39819);
xnor U41624 (N_41624,N_35739,N_35401);
nand U41625 (N_41625,N_35459,N_35077);
or U41626 (N_41626,N_38997,N_35439);
nor U41627 (N_41627,N_39413,N_35436);
nand U41628 (N_41628,N_37709,N_37616);
nand U41629 (N_41629,N_38345,N_35903);
and U41630 (N_41630,N_38538,N_38931);
nand U41631 (N_41631,N_38197,N_38780);
nand U41632 (N_41632,N_37942,N_38446);
xnor U41633 (N_41633,N_36836,N_35650);
or U41634 (N_41634,N_35333,N_38428);
or U41635 (N_41635,N_37492,N_36024);
and U41636 (N_41636,N_36231,N_35702);
nor U41637 (N_41637,N_35176,N_35585);
xor U41638 (N_41638,N_37258,N_35881);
nor U41639 (N_41639,N_39056,N_36870);
nor U41640 (N_41640,N_39693,N_36517);
and U41641 (N_41641,N_37264,N_35516);
xnor U41642 (N_41642,N_35424,N_35782);
nand U41643 (N_41643,N_36470,N_36947);
or U41644 (N_41644,N_38387,N_35955);
nor U41645 (N_41645,N_36558,N_36401);
nor U41646 (N_41646,N_39457,N_38136);
and U41647 (N_41647,N_35828,N_37909);
xnor U41648 (N_41648,N_35844,N_36314);
nand U41649 (N_41649,N_39721,N_35740);
nor U41650 (N_41650,N_38911,N_38619);
and U41651 (N_41651,N_38010,N_39387);
and U41652 (N_41652,N_37717,N_36153);
and U41653 (N_41653,N_38329,N_35185);
and U41654 (N_41654,N_36834,N_38309);
nand U41655 (N_41655,N_39350,N_35970);
and U41656 (N_41656,N_37848,N_36545);
or U41657 (N_41657,N_38079,N_37669);
or U41658 (N_41658,N_35638,N_35668);
nor U41659 (N_41659,N_38946,N_38956);
or U41660 (N_41660,N_39478,N_36146);
or U41661 (N_41661,N_36918,N_36864);
or U41662 (N_41662,N_35153,N_35523);
or U41663 (N_41663,N_35447,N_38600);
nand U41664 (N_41664,N_38067,N_39961);
or U41665 (N_41665,N_36936,N_36501);
or U41666 (N_41666,N_35532,N_37133);
xor U41667 (N_41667,N_37186,N_38127);
or U41668 (N_41668,N_35458,N_38864);
nand U41669 (N_41669,N_37158,N_39666);
nor U41670 (N_41670,N_39600,N_36334);
xnor U41671 (N_41671,N_38585,N_35832);
and U41672 (N_41672,N_38673,N_39301);
nor U41673 (N_41673,N_35715,N_35014);
nand U41674 (N_41674,N_39057,N_38549);
nand U41675 (N_41675,N_35149,N_36699);
nor U41676 (N_41676,N_39300,N_37874);
xnor U41677 (N_41677,N_35978,N_37570);
or U41678 (N_41678,N_35688,N_37815);
nand U41679 (N_41679,N_39291,N_35166);
nor U41680 (N_41680,N_38926,N_36280);
or U41681 (N_41681,N_36036,N_38834);
xor U41682 (N_41682,N_36071,N_37210);
nand U41683 (N_41683,N_39563,N_36342);
or U41684 (N_41684,N_38818,N_35488);
and U41685 (N_41685,N_38582,N_36059);
nand U41686 (N_41686,N_39552,N_36736);
xor U41687 (N_41687,N_36404,N_35522);
xnor U41688 (N_41688,N_38459,N_36448);
xnor U41689 (N_41689,N_36408,N_35886);
or U41690 (N_41690,N_36480,N_37352);
nor U41691 (N_41691,N_39466,N_35223);
xnor U41692 (N_41692,N_36041,N_38909);
nor U41693 (N_41693,N_35703,N_38393);
nor U41694 (N_41694,N_38102,N_39232);
xnor U41695 (N_41695,N_35640,N_37708);
nor U41696 (N_41696,N_36630,N_37856);
nand U41697 (N_41697,N_35826,N_35805);
or U41698 (N_41698,N_35470,N_35056);
nand U41699 (N_41699,N_39117,N_38018);
xor U41700 (N_41700,N_38980,N_36816);
xnor U41701 (N_41701,N_37628,N_38993);
and U41702 (N_41702,N_36953,N_36081);
or U41703 (N_41703,N_39577,N_36293);
and U41704 (N_41704,N_39629,N_36307);
nand U41705 (N_41705,N_36339,N_35478);
nor U41706 (N_41706,N_35722,N_36156);
or U41707 (N_41707,N_36261,N_37666);
and U41708 (N_41708,N_35771,N_39829);
nor U41709 (N_41709,N_36138,N_38314);
or U41710 (N_41710,N_38332,N_35619);
nor U41711 (N_41711,N_38265,N_39085);
and U41712 (N_41712,N_35503,N_35212);
xor U41713 (N_41713,N_35259,N_39277);
nor U41714 (N_41714,N_36355,N_35270);
or U41715 (N_41715,N_36853,N_36435);
nand U41716 (N_41716,N_36535,N_37608);
xor U41717 (N_41717,N_38951,N_39899);
or U41718 (N_41718,N_39082,N_38307);
nor U41719 (N_41719,N_37138,N_37022);
nor U41720 (N_41720,N_37993,N_38350);
nand U41721 (N_41721,N_39520,N_36619);
nand U41722 (N_41722,N_38502,N_39092);
nor U41723 (N_41723,N_38896,N_36455);
xnor U41724 (N_41724,N_35344,N_38587);
nor U41725 (N_41725,N_39784,N_36102);
and U41726 (N_41726,N_35865,N_36894);
or U41727 (N_41727,N_39302,N_36067);
xor U41728 (N_41728,N_39761,N_39931);
or U41729 (N_41729,N_38865,N_38029);
xnor U41730 (N_41730,N_36742,N_35071);
xnor U41731 (N_41731,N_36233,N_37486);
nand U41732 (N_41732,N_36793,N_38483);
xor U41733 (N_41733,N_35971,N_37394);
nand U41734 (N_41734,N_38133,N_39071);
and U41735 (N_41735,N_36636,N_37087);
and U41736 (N_41736,N_35154,N_35234);
nor U41737 (N_41737,N_39443,N_35651);
and U41738 (N_41738,N_38729,N_39158);
xor U41739 (N_41739,N_38773,N_39080);
or U41740 (N_41740,N_39991,N_37307);
or U41741 (N_41741,N_39849,N_35364);
or U41742 (N_41742,N_39663,N_35290);
nor U41743 (N_41743,N_35405,N_37960);
nand U41744 (N_41744,N_36452,N_37444);
nand U41745 (N_41745,N_37924,N_36837);
and U41746 (N_41746,N_36219,N_36444);
nor U41747 (N_41747,N_39467,N_36391);
xnor U41748 (N_41748,N_38610,N_39971);
nand U41749 (N_41749,N_39865,N_38545);
nand U41750 (N_41750,N_38237,N_37376);
and U41751 (N_41751,N_37687,N_38436);
and U41752 (N_41752,N_36379,N_37949);
nor U41753 (N_41753,N_35103,N_36204);
nor U41754 (N_41754,N_35852,N_37889);
nor U41755 (N_41755,N_38221,N_38743);
nand U41756 (N_41756,N_37340,N_36011);
and U41757 (N_41757,N_37716,N_38157);
and U41758 (N_41758,N_39613,N_39440);
or U41759 (N_41759,N_38069,N_36359);
and U41760 (N_41760,N_37402,N_37544);
or U41761 (N_41761,N_35449,N_35880);
xnor U41762 (N_41762,N_37680,N_35085);
xnor U41763 (N_41763,N_35608,N_39828);
or U41764 (N_41764,N_37001,N_38126);
and U41765 (N_41765,N_35589,N_35994);
xor U41766 (N_41766,N_37910,N_37796);
xnor U41767 (N_41767,N_39381,N_37865);
xnor U41768 (N_41768,N_38862,N_37807);
nor U41769 (N_41769,N_39559,N_38325);
nand U41770 (N_41770,N_35558,N_35186);
or U41771 (N_41771,N_39898,N_38728);
or U41772 (N_41772,N_39617,N_35044);
and U41773 (N_41773,N_39907,N_36561);
xnor U41774 (N_41774,N_37787,N_37074);
xnor U41775 (N_41775,N_36955,N_35289);
nand U41776 (N_41776,N_37698,N_38526);
and U41777 (N_41777,N_36930,N_37031);
nor U41778 (N_41778,N_36288,N_35297);
nand U41779 (N_41779,N_37691,N_39631);
and U41780 (N_41780,N_35399,N_38402);
nand U41781 (N_41781,N_35893,N_37541);
nor U41782 (N_41782,N_39565,N_39263);
nand U41783 (N_41783,N_36999,N_35171);
xor U41784 (N_41784,N_36587,N_35263);
nor U41785 (N_41785,N_36143,N_38737);
and U41786 (N_41786,N_38558,N_39486);
xor U41787 (N_41787,N_37685,N_36533);
or U41788 (N_41788,N_35183,N_39426);
xor U41789 (N_41789,N_35361,N_38745);
or U41790 (N_41790,N_38156,N_38259);
nand U41791 (N_41791,N_35649,N_35024);
nor U41792 (N_41792,N_37281,N_38758);
and U41793 (N_41793,N_37644,N_36161);
xor U41794 (N_41794,N_39339,N_35351);
and U41795 (N_41795,N_37798,N_38352);
or U41796 (N_41796,N_38208,N_38882);
or U41797 (N_41797,N_39788,N_39587);
xnor U41798 (N_41798,N_36008,N_35417);
nand U41799 (N_41799,N_37435,N_37163);
nand U41800 (N_41800,N_37989,N_38249);
or U41801 (N_41801,N_39821,N_37196);
and U41802 (N_41802,N_36852,N_37749);
xnor U41803 (N_41803,N_39826,N_38542);
nor U41804 (N_41804,N_36043,N_38432);
or U41805 (N_41805,N_36746,N_36350);
xnor U41806 (N_41806,N_35586,N_37211);
and U41807 (N_41807,N_37612,N_36631);
or U41808 (N_41808,N_36302,N_39266);
xor U41809 (N_41809,N_35139,N_37576);
nor U41810 (N_41810,N_36268,N_37002);
or U41811 (N_41811,N_35772,N_35770);
nor U41812 (N_41812,N_36995,N_39189);
and U41813 (N_41813,N_39733,N_38167);
or U41814 (N_41814,N_39344,N_35063);
and U41815 (N_41815,N_35159,N_39223);
or U41816 (N_41816,N_37328,N_36009);
and U41817 (N_41817,N_37833,N_37089);
nor U41818 (N_41818,N_35809,N_35541);
xnor U41819 (N_41819,N_37619,N_35507);
and U41820 (N_41820,N_39647,N_38049);
nand U41821 (N_41821,N_36818,N_35534);
xor U41822 (N_41822,N_36911,N_39087);
xor U41823 (N_41823,N_37564,N_38534);
or U41824 (N_41824,N_36941,N_38655);
nand U41825 (N_41825,N_38021,N_39906);
nand U41826 (N_41826,N_39735,N_38958);
nor U41827 (N_41827,N_39305,N_38453);
and U41828 (N_41828,N_36037,N_35878);
or U41829 (N_41829,N_37639,N_37434);
or U41830 (N_41830,N_36518,N_37944);
nand U41831 (N_41831,N_36241,N_38379);
nor U41832 (N_41832,N_38341,N_36309);
or U41833 (N_41833,N_38684,N_39407);
and U41834 (N_41834,N_37734,N_38605);
and U41835 (N_41835,N_36674,N_37112);
or U41836 (N_41836,N_37032,N_39008);
xor U41837 (N_41837,N_38266,N_36318);
or U41838 (N_41838,N_38572,N_37320);
and U41839 (N_41839,N_35355,N_37606);
and U41840 (N_41840,N_37765,N_35641);
nand U41841 (N_41841,N_36415,N_36033);
and U41842 (N_41842,N_37407,N_38041);
nor U41843 (N_41843,N_38923,N_37025);
and U41844 (N_41844,N_37261,N_39762);
or U41845 (N_41845,N_38892,N_37338);
or U41846 (N_41846,N_38046,N_37862);
nand U41847 (N_41847,N_35248,N_37380);
nor U41848 (N_41848,N_39973,N_38476);
xor U41849 (N_41849,N_38064,N_38279);
nor U41850 (N_41850,N_35542,N_37241);
nor U41851 (N_41851,N_39643,N_38879);
and U41852 (N_41852,N_38770,N_37731);
nor U41853 (N_41853,N_37964,N_35498);
nand U41854 (N_41854,N_38532,N_38568);
or U41855 (N_41855,N_36245,N_37642);
or U41856 (N_41856,N_36413,N_37121);
or U41857 (N_41857,N_38438,N_36661);
xnor U41858 (N_41858,N_38618,N_38847);
nand U41859 (N_41859,N_38384,N_36872);
nand U41860 (N_41860,N_39517,N_36536);
nand U41861 (N_41861,N_38837,N_36277);
nor U41862 (N_41862,N_37070,N_36878);
nor U41863 (N_41863,N_37517,N_36004);
nor U41864 (N_41864,N_38540,N_36247);
nor U41865 (N_41865,N_36573,N_39956);
nor U41866 (N_41866,N_39869,N_39401);
nor U41867 (N_41867,N_37613,N_38121);
nor U41868 (N_41868,N_35266,N_39774);
or U41869 (N_41869,N_36546,N_38338);
and U41870 (N_41870,N_38966,N_39521);
xor U41871 (N_41871,N_37890,N_36551);
and U41872 (N_41872,N_38689,N_35490);
xor U41873 (N_41873,N_35500,N_35681);
nand U41874 (N_41874,N_35664,N_38359);
xnor U41875 (N_41875,N_38774,N_38302);
and U41876 (N_41876,N_35074,N_37418);
nand U41877 (N_41877,N_35316,N_35203);
and U41878 (N_41878,N_38635,N_39481);
or U41879 (N_41879,N_38261,N_36504);
xor U41880 (N_41880,N_38081,N_39847);
nor U41881 (N_41881,N_39598,N_38790);
nand U41882 (N_41882,N_36417,N_35753);
xnor U41883 (N_41883,N_35197,N_35348);
or U41884 (N_41884,N_37348,N_36000);
nor U41885 (N_41885,N_35100,N_35925);
and U41886 (N_41886,N_36786,N_39890);
xnor U41887 (N_41887,N_38181,N_38487);
xor U41888 (N_41888,N_35756,N_38667);
xnor U41889 (N_41889,N_37036,N_37268);
or U41890 (N_41890,N_37637,N_37494);
xor U41891 (N_41891,N_39790,N_36325);
xor U41892 (N_41892,N_35320,N_38772);
nand U41893 (N_41893,N_37772,N_37431);
or U41894 (N_41894,N_39493,N_39172);
nand U41895 (N_41895,N_36963,N_35754);
nand U41896 (N_41896,N_37223,N_35035);
and U41897 (N_41897,N_39121,N_36216);
nor U41898 (N_41898,N_36380,N_38591);
xor U41899 (N_41899,N_35091,N_36252);
xnor U41900 (N_41900,N_36290,N_37886);
and U41901 (N_41901,N_39000,N_35283);
and U41902 (N_41902,N_38390,N_39469);
nand U41903 (N_41903,N_38467,N_37169);
and U41904 (N_41904,N_35699,N_37015);
nor U41905 (N_41905,N_35981,N_35900);
or U41906 (N_41906,N_39514,N_39949);
nor U41907 (N_41907,N_36642,N_38295);
and U41908 (N_41908,N_36201,N_36637);
nor U41909 (N_41909,N_36338,N_37224);
nor U41910 (N_41910,N_39280,N_37733);
nand U41911 (N_41911,N_36079,N_35761);
nand U41912 (N_41912,N_37060,N_38669);
nor U41913 (N_41913,N_39665,N_39435);
and U41914 (N_41914,N_38964,N_38914);
or U41915 (N_41915,N_35250,N_39025);
nand U41916 (N_41916,N_38050,N_39554);
or U41917 (N_41917,N_36666,N_37284);
nor U41918 (N_41918,N_38340,N_38499);
nand U41919 (N_41919,N_36015,N_36698);
nand U41920 (N_41920,N_37491,N_36154);
nand U41921 (N_41921,N_36577,N_37209);
or U41922 (N_41922,N_39233,N_39728);
nand U41923 (N_41923,N_37693,N_36633);
nand U41924 (N_41924,N_39955,N_35357);
and U41925 (N_41925,N_38878,N_36611);
nor U41926 (N_41926,N_35851,N_36987);
nand U41927 (N_41927,N_38808,N_36063);
xnor U41928 (N_41928,N_35866,N_35547);
nand U41929 (N_41929,N_39686,N_39436);
and U41930 (N_41930,N_39688,N_36029);
nor U41931 (N_41931,N_39181,N_39249);
xnor U41932 (N_41932,N_39185,N_36914);
and U41933 (N_41933,N_38409,N_38093);
or U41934 (N_41934,N_37756,N_37033);
xor U41935 (N_41935,N_39641,N_36649);
or U41936 (N_41936,N_35625,N_37627);
and U41937 (N_41937,N_38191,N_35487);
or U41938 (N_41938,N_35217,N_36749);
and U41939 (N_41939,N_38429,N_35215);
xnor U41940 (N_41940,N_37947,N_35629);
and U41941 (N_41941,N_35206,N_35340);
nand U41942 (N_41942,N_35533,N_37715);
nor U41943 (N_41943,N_36745,N_38840);
xnor U41944 (N_41944,N_37979,N_38976);
xnor U41945 (N_41945,N_36400,N_38701);
and U41946 (N_41946,N_36274,N_35959);
nand U41947 (N_41947,N_39246,N_37208);
nor U41948 (N_41948,N_36885,N_39980);
nor U41949 (N_41949,N_39023,N_39548);
xnor U41950 (N_41950,N_37721,N_38062);
xnor U41951 (N_41951,N_38298,N_35010);
xnor U41952 (N_41952,N_39875,N_39090);
nand U41953 (N_41953,N_39962,N_38898);
nand U41954 (N_41954,N_35982,N_35951);
xor U41955 (N_41955,N_39557,N_37457);
and U41956 (N_41956,N_36711,N_39690);
and U41957 (N_41957,N_39566,N_39004);
or U41958 (N_41958,N_37694,N_35128);
nor U41959 (N_41959,N_39738,N_37672);
nor U41960 (N_41960,N_38116,N_37839);
nand U41961 (N_41961,N_38421,N_38184);
and U41962 (N_41962,N_38440,N_39161);
and U41963 (N_41963,N_36512,N_36263);
xnor U41964 (N_41964,N_36304,N_39909);
xor U41965 (N_41965,N_39911,N_35803);
nand U41966 (N_41966,N_39982,N_35784);
and U41967 (N_41967,N_38617,N_38791);
and U41968 (N_41968,N_35040,N_36341);
xnor U41969 (N_41969,N_37248,N_35251);
xor U41970 (N_41970,N_38070,N_35871);
and U41971 (N_41971,N_38528,N_39272);
xor U41972 (N_41972,N_39942,N_39009);
nand U41973 (N_41973,N_36589,N_39261);
xor U41974 (N_41974,N_37243,N_36829);
xnor U41975 (N_41975,N_36140,N_39839);
nor U41976 (N_41976,N_38073,N_37830);
nand U41977 (N_41977,N_39753,N_36232);
nand U41978 (N_41978,N_39769,N_37012);
xnor U41979 (N_41979,N_36583,N_38253);
or U41980 (N_41980,N_39603,N_37791);
nand U41981 (N_41981,N_36950,N_36772);
or U41982 (N_41982,N_37448,N_39742);
nand U41983 (N_41983,N_37855,N_38082);
nand U41984 (N_41984,N_36303,N_37219);
nand U41985 (N_41985,N_36909,N_35440);
nor U41986 (N_41986,N_36717,N_35568);
and U41987 (N_41987,N_35179,N_36708);
and U41988 (N_41988,N_39160,N_37923);
nor U41989 (N_41989,N_38894,N_39016);
nor U41990 (N_41990,N_39416,N_38141);
and U41991 (N_41991,N_35599,N_39675);
nor U41992 (N_41992,N_38211,N_36598);
nor U41993 (N_41993,N_39658,N_35221);
and U41994 (N_41994,N_36186,N_39167);
nand U41995 (N_41995,N_35765,N_39703);
and U41996 (N_41996,N_37755,N_39479);
nor U41997 (N_41997,N_36797,N_38101);
nor U41998 (N_41998,N_37364,N_38930);
and U41999 (N_41999,N_36326,N_36988);
nand U42000 (N_42000,N_37246,N_36305);
nor U42001 (N_42001,N_35622,N_38984);
xor U42002 (N_42002,N_39606,N_39737);
and U42003 (N_42003,N_37869,N_35633);
nor U42004 (N_42004,N_35983,N_35023);
or U42005 (N_42005,N_39648,N_38719);
or U42006 (N_42006,N_37081,N_38371);
nand U42007 (N_42007,N_36634,N_38535);
xnor U42008 (N_42008,N_38613,N_35587);
or U42009 (N_42009,N_36171,N_35790);
xor U42010 (N_42010,N_38827,N_37965);
nand U42011 (N_42011,N_39064,N_36503);
xnor U42012 (N_42012,N_36550,N_37762);
xor U42013 (N_42013,N_39850,N_39373);
nand U42014 (N_42014,N_35214,N_38495);
and U42015 (N_42015,N_36362,N_37373);
or U42016 (N_42016,N_36164,N_35939);
nor U42017 (N_42017,N_37780,N_39873);
xor U42018 (N_42018,N_37124,N_38906);
and U42019 (N_42019,N_38297,N_38407);
nor U42020 (N_42020,N_36879,N_35690);
nand U42021 (N_42021,N_36421,N_39140);
nor U42022 (N_42022,N_35309,N_35594);
nor U42023 (N_42023,N_36644,N_38999);
xnor U42024 (N_42024,N_38028,N_37881);
nor U42025 (N_42025,N_35232,N_39292);
nor U42026 (N_42026,N_36394,N_36089);
or U42027 (N_42027,N_39597,N_39635);
and U42028 (N_42028,N_38972,N_37625);
or U42029 (N_42029,N_37882,N_35343);
xor U42030 (N_42030,N_38686,N_37422);
and U42031 (N_42031,N_36812,N_36428);
nor U42032 (N_42032,N_36653,N_39669);
xor U42033 (N_42033,N_35150,N_35932);
nand U42034 (N_42034,N_39731,N_36210);
and U42035 (N_42035,N_35631,N_36108);
and U42036 (N_42036,N_38888,N_39910);
nand U42037 (N_42037,N_39079,N_37042);
or U42038 (N_42038,N_39132,N_38955);
xor U42039 (N_42039,N_39050,N_35762);
nand U42040 (N_42040,N_35094,N_38363);
xor U42041 (N_42041,N_35680,N_35460);
xor U42042 (N_42042,N_39518,N_38945);
or U42043 (N_42043,N_38718,N_38299);
nand U42044 (N_42044,N_37718,N_37043);
and U42045 (N_42045,N_38515,N_36211);
and U42046 (N_42046,N_37378,N_36473);
nor U42047 (N_42047,N_38240,N_38895);
xnor U42048 (N_42048,N_38501,N_35285);
nor U42049 (N_42049,N_37781,N_39928);
nand U42050 (N_42050,N_36640,N_38375);
and U42051 (N_42051,N_38810,N_35508);
and U42052 (N_42052,N_35787,N_35299);
xnor U42053 (N_42053,N_35562,N_37484);
and U42054 (N_42054,N_37071,N_35905);
and U42055 (N_42055,N_39073,N_36495);
or U42056 (N_42056,N_35904,N_39994);
xnor U42057 (N_42057,N_36003,N_38871);
nand U42058 (N_42058,N_38638,N_36602);
nand U42059 (N_42059,N_35663,N_38560);
nor U42060 (N_42060,N_35596,N_36553);
or U42061 (N_42061,N_35813,N_35210);
nor U42062 (N_42062,N_38378,N_39933);
xnor U42063 (N_42063,N_36074,N_39067);
and U42064 (N_42064,N_36283,N_39239);
nor U42065 (N_42065,N_37144,N_35988);
and U42066 (N_42066,N_35684,N_37926);
xnor U42067 (N_42067,N_35658,N_37690);
or U42068 (N_42068,N_37115,N_35783);
nand U42069 (N_42069,N_37589,N_37252);
and U42070 (N_42070,N_38075,N_35135);
nand U42071 (N_42071,N_39547,N_36764);
and U42072 (N_42072,N_39257,N_37641);
or U42073 (N_42073,N_36979,N_39153);
nand U42074 (N_42074,N_39712,N_39485);
nor U42075 (N_42075,N_37237,N_38588);
nor U42076 (N_42076,N_39354,N_35388);
or U42077 (N_42077,N_39360,N_35341);
or U42078 (N_42078,N_35662,N_36179);
and U42079 (N_42079,N_39483,N_35977);
nand U42080 (N_42080,N_37129,N_38009);
and U42081 (N_42081,N_39531,N_39091);
or U42082 (N_42082,N_37674,N_37545);
and U42083 (N_42083,N_35705,N_38269);
or U42084 (N_42084,N_35207,N_38433);
and U42085 (N_42085,N_37099,N_39382);
and U42086 (N_42086,N_39420,N_37454);
and U42087 (N_42087,N_35075,N_37826);
and U42088 (N_42088,N_39104,N_38664);
nor U42089 (N_42089,N_37582,N_38491);
nor U42090 (N_42090,N_38995,N_39901);
nand U42091 (N_42091,N_35472,N_37240);
and U42092 (N_42092,N_37079,N_36097);
xnor U42093 (N_42093,N_36085,N_35654);
and U42094 (N_42094,N_36928,N_39844);
nand U42095 (N_42095,N_35510,N_35058);
nor U42096 (N_42096,N_38744,N_37421);
nor U42097 (N_42097,N_35420,N_36264);
nor U42098 (N_42098,N_38251,N_36690);
nand U42099 (N_42099,N_38985,N_38829);
xnor U42100 (N_42100,N_36425,N_37783);
nand U42101 (N_42101,N_37656,N_37379);
or U42102 (N_42102,N_38267,N_36624);
nand U42103 (N_42103,N_35823,N_36835);
nand U42104 (N_42104,N_35591,N_38115);
and U42105 (N_42105,N_39205,N_36528);
nor U42106 (N_42106,N_36240,N_35342);
nand U42107 (N_42107,N_38839,N_39441);
nand U42108 (N_42108,N_39123,N_38257);
nand U42109 (N_42109,N_39318,N_39192);
or U42110 (N_42110,N_39745,N_38015);
nand U42111 (N_42111,N_35237,N_39059);
and U42112 (N_42112,N_35630,N_36566);
nand U42113 (N_42113,N_38335,N_37665);
nand U42114 (N_42114,N_39255,N_37134);
nor U42115 (N_42115,N_37318,N_36695);
nor U42116 (N_42116,N_39393,N_36177);
and U42117 (N_42117,N_36710,N_36427);
nor U42118 (N_42118,N_39967,N_36697);
or U42119 (N_42119,N_36939,N_39671);
and U42120 (N_42120,N_38640,N_38802);
xor U42121 (N_42121,N_35278,N_39332);
and U42122 (N_42122,N_39324,N_36769);
or U42123 (N_42123,N_39471,N_35425);
and U42124 (N_42124,N_35835,N_35838);
xor U42125 (N_42125,N_39052,N_35291);
nand U42126 (N_42126,N_38250,N_38730);
nand U42127 (N_42127,N_35738,N_35642);
nand U42128 (N_42128,N_38592,N_38210);
or U42129 (N_42129,N_35501,N_35693);
and U42130 (N_42130,N_38376,N_35675);
or U42131 (N_42131,N_37019,N_36915);
xnor U42132 (N_42132,N_39732,N_39135);
or U42133 (N_42133,N_39883,N_36658);
nor U42134 (N_42134,N_36515,N_39668);
and U42135 (N_42135,N_39818,N_37778);
or U42136 (N_42136,N_35026,N_39696);
and U42137 (N_42137,N_39176,N_36320);
nand U42138 (N_42138,N_37335,N_39871);
nand U42139 (N_42139,N_37064,N_39726);
and U42140 (N_42140,N_38365,N_38505);
xnor U42141 (N_42141,N_38189,N_38362);
nor U42142 (N_42142,N_35099,N_36026);
xor U42143 (N_42143,N_38782,N_37410);
nor U42144 (N_42144,N_39099,N_38647);
or U42145 (N_42145,N_35926,N_35249);
xnor U42146 (N_42146,N_39734,N_35400);
or U42147 (N_42147,N_38024,N_36608);
nand U42148 (N_42148,N_35588,N_35407);
xnor U42149 (N_42149,N_39293,N_35798);
nand U42150 (N_42150,N_38254,N_36092);
or U42151 (N_42151,N_36091,N_35032);
xnor U42152 (N_42152,N_38805,N_35573);
or U42153 (N_42153,N_38238,N_35791);
or U42154 (N_42154,N_39108,N_38207);
xor U42155 (N_42155,N_38422,N_39494);
or U42156 (N_42156,N_36135,N_38536);
or U42157 (N_42157,N_35966,N_36656);
and U42158 (N_42158,N_36113,N_38586);
nand U42159 (N_42159,N_38872,N_38480);
or U42160 (N_42160,N_37304,N_39926);
and U42161 (N_42161,N_36083,N_36385);
and U42162 (N_42162,N_38244,N_37037);
nor U42163 (N_42163,N_36702,N_37342);
and U42164 (N_42164,N_39288,N_39626);
and U42165 (N_42165,N_38981,N_39628);
and U42166 (N_42166,N_39989,N_39437);
nor U42167 (N_42167,N_39802,N_37301);
or U42168 (N_42168,N_39752,N_39575);
or U42169 (N_42169,N_38391,N_36419);
and U42170 (N_42170,N_38941,N_38025);
xor U42171 (N_42171,N_35494,N_37679);
xnor U42172 (N_42172,N_38518,N_38693);
xor U42173 (N_42173,N_39682,N_37751);
xor U42174 (N_42174,N_37367,N_35055);
and U42175 (N_42175,N_35043,N_36049);
nand U42176 (N_42176,N_35709,N_36396);
or U42177 (N_42177,N_37302,N_38554);
or U42178 (N_42178,N_39125,N_38195);
nand U42179 (N_42179,N_37736,N_39038);
or U42180 (N_42180,N_39694,N_37023);
xnor U42181 (N_42181,N_39919,N_35356);
and U42182 (N_42182,N_36966,N_39572);
xor U42183 (N_42183,N_39018,N_36555);
xnor U42184 (N_42184,N_35996,N_36822);
nand U42185 (N_42185,N_39007,N_39868);
nand U42186 (N_42186,N_37445,N_36548);
nand U42187 (N_42187,N_35218,N_39798);
or U42188 (N_42188,N_37746,N_35360);
xnor U42189 (N_42189,N_35175,N_38514);
nor U42190 (N_42190,N_37008,N_35673);
or U42191 (N_42191,N_37399,N_35768);
and U42192 (N_42192,N_39599,N_35331);
or U42193 (N_42193,N_35862,N_35802);
nand U42194 (N_42194,N_38868,N_39043);
nand U42195 (N_42195,N_37510,N_36119);
nand U42196 (N_42196,N_39754,N_38256);
or U42197 (N_42197,N_37676,N_39555);
xor U42198 (N_42198,N_37148,N_35870);
or U42199 (N_42199,N_39615,N_35392);
xor U42200 (N_42200,N_37977,N_35453);
nand U42201 (N_42201,N_39229,N_38031);
xnor U42202 (N_42202,N_39116,N_39182);
nand U42203 (N_42203,N_36254,N_39188);
nand U42204 (N_42204,N_37767,N_39372);
nand U42205 (N_42205,N_37808,N_35301);
and U42206 (N_42206,N_38703,N_37732);
xnor U42207 (N_42207,N_39164,N_39858);
or U42208 (N_42208,N_37358,N_35520);
and U42209 (N_42209,N_36931,N_35371);
and U42210 (N_42210,N_39438,N_36705);
nor U42211 (N_42211,N_35670,N_39206);
xor U42212 (N_42212,N_39499,N_36409);
xor U42213 (N_42213,N_38312,N_39748);
nand U42214 (N_42214,N_39200,N_38444);
nand U42215 (N_42215,N_36183,N_36098);
or U42216 (N_42216,N_35191,N_37255);
xor U42217 (N_42217,N_35292,N_38620);
or U42218 (N_42218,N_36105,N_36590);
nor U42219 (N_42219,N_39207,N_39704);
nor U42220 (N_42220,N_38243,N_39995);
nand U42221 (N_42221,N_36782,N_38950);
nor U42222 (N_42222,N_38454,N_36159);
or U42223 (N_42223,N_39330,N_36680);
nand U42224 (N_42224,N_37745,N_37010);
or U42225 (N_42225,N_35816,N_38051);
and U42226 (N_42226,N_35462,N_35001);
or U42227 (N_42227,N_37424,N_38527);
nor U42228 (N_42228,N_38784,N_35659);
and U42229 (N_42229,N_39888,N_36652);
xor U42230 (N_42230,N_37802,N_36670);
or U42231 (N_42231,N_36365,N_39854);
xor U42232 (N_42232,N_35924,N_39516);
xnor U42233 (N_42233,N_37970,N_37688);
or U42234 (N_42234,N_38623,N_38629);
or U42235 (N_42235,N_36759,N_36796);
nand U42236 (N_42236,N_37366,N_35155);
or U42237 (N_42237,N_37714,N_35222);
nand U42238 (N_42238,N_39527,N_37885);
nand U42239 (N_42239,N_37355,N_39400);
nand U42240 (N_42240,N_38928,N_36683);
and U42241 (N_42241,N_38248,N_35757);
nor U42242 (N_42242,N_36321,N_36441);
and U42243 (N_42243,N_39673,N_36006);
nand U42244 (N_42244,N_35481,N_38968);
xor U42245 (N_42245,N_35471,N_36593);
or U42246 (N_42246,N_36607,N_35019);
nand U42247 (N_42247,N_38967,N_36076);
xnor U42248 (N_42248,N_35723,N_37187);
or U42249 (N_42249,N_37523,N_39165);
nor U42250 (N_42250,N_37051,N_36500);
or U42251 (N_42251,N_36672,N_36599);
xor U42252 (N_42252,N_38750,N_35752);
nand U42253 (N_42253,N_38783,N_36295);
xor U42254 (N_42254,N_37287,N_37396);
nor U42255 (N_42255,N_37940,N_39604);
or U42256 (N_42256,N_37007,N_36060);
nor U42257 (N_42257,N_37468,N_37880);
and U42258 (N_42258,N_38090,N_35141);
nor U42259 (N_42259,N_36256,N_35929);
nor U42260 (N_42260,N_35669,N_37461);
or U42261 (N_42261,N_36828,N_39843);
nand U42262 (N_42262,N_37097,N_38012);
xor U42263 (N_42263,N_36684,N_35751);
or U42264 (N_42264,N_36489,N_35759);
xor U42265 (N_42265,N_38765,N_38543);
nand U42266 (N_42266,N_35788,N_38326);
and U42267 (N_42267,N_35189,N_38531);
nor U42268 (N_42268,N_38577,N_38800);
nand U42269 (N_42269,N_35964,N_37473);
or U42270 (N_42270,N_38416,N_39447);
or U42271 (N_42271,N_36934,N_38205);
or U42272 (N_42272,N_38822,N_39662);
or U42273 (N_42273,N_39894,N_35707);
and U42274 (N_42274,N_36805,N_37005);
nor U42275 (N_42275,N_39465,N_39637);
or U42276 (N_42276,N_38080,N_36627);
nor U42277 (N_42277,N_39540,N_37346);
xnor U42278 (N_42278,N_38289,N_35660);
or U42279 (N_42279,N_38318,N_39653);
nor U42280 (N_42280,N_38437,N_35780);
nand U42281 (N_42281,N_37520,N_39834);
xnor U42282 (N_42282,N_39824,N_38886);
or U42283 (N_42283,N_37200,N_36202);
nand U42284 (N_42284,N_38982,N_37800);
nand U42285 (N_42285,N_37107,N_35106);
and U42286 (N_42286,N_36069,N_38877);
nand U42287 (N_42287,N_39741,N_37324);
nand U42288 (N_42288,N_36180,N_36196);
nor U42289 (N_42289,N_37611,N_37567);
xnor U42290 (N_42290,N_36487,N_35198);
xnor U42291 (N_42291,N_39474,N_39794);
and U42292 (N_42292,N_36740,N_38118);
nand U42293 (N_42293,N_38011,N_36020);
nand U42294 (N_42294,N_37017,N_35461);
or U42295 (N_42295,N_37362,N_37068);
or U42296 (N_42296,N_38836,N_36116);
nor U42297 (N_42297,N_38796,N_35854);
xor U42298 (N_42298,N_38920,N_37120);
or U42299 (N_42299,N_36978,N_36502);
and U42300 (N_42300,N_37440,N_36526);
and U42301 (N_42301,N_37483,N_39178);
and U42302 (N_42302,N_39830,N_35190);
or U42303 (N_42303,N_37321,N_38607);
or U42304 (N_42304,N_36946,N_39699);
xor U42305 (N_42305,N_39422,N_37727);
and U42306 (N_42306,N_35493,N_36921);
or U42307 (N_42307,N_36065,N_39027);
and U42308 (N_42308,N_38202,N_37959);
and U42309 (N_42309,N_37686,N_38038);
xor U42310 (N_42310,N_37045,N_37296);
or U42311 (N_42311,N_38427,N_39978);
xnor U42312 (N_42312,N_36260,N_35455);
nand U42313 (N_42313,N_36756,N_37175);
nand U42314 (N_42314,N_35162,N_39618);
nor U42315 (N_42315,N_35402,N_36743);
and U42316 (N_42316,N_37844,N_37617);
nor U42317 (N_42317,N_37563,N_35574);
nand U42318 (N_42318,N_39805,N_37724);
nor U42319 (N_42319,N_39017,N_38410);
nor U42320 (N_42320,N_35350,N_36012);
nand U42321 (N_42321,N_36430,N_37512);
nor U42322 (N_42322,N_35741,N_37730);
nand U42323 (N_42323,N_39316,N_39256);
or U42324 (N_42324,N_35134,N_35543);
nand U42325 (N_42325,N_38092,N_38716);
nand U42326 (N_42326,N_39760,N_35086);
or U42327 (N_42327,N_36169,N_35901);
or U42328 (N_42328,N_38762,N_36617);
or U42329 (N_42329,N_37777,N_39427);
and U42330 (N_42330,N_38236,N_38798);
and U42331 (N_42331,N_38965,N_35146);
xor U42332 (N_42332,N_37273,N_35860);
nand U42333 (N_42333,N_36276,N_39303);
or U42334 (N_42334,N_39415,N_39713);
xnor U42335 (N_42335,N_38653,N_37797);
and U42336 (N_42336,N_38439,N_37507);
nor U42337 (N_42337,N_38336,N_37052);
or U42338 (N_42338,N_36696,N_36937);
xor U42339 (N_42339,N_37829,N_39656);
xnor U42340 (N_42340,N_36058,N_36267);
xnor U42341 (N_42341,N_35048,N_35666);
nor U42342 (N_42342,N_35369,N_39964);
nor U42343 (N_42343,N_35511,N_38034);
and U42344 (N_42344,N_38305,N_37206);
or U42345 (N_42345,N_36220,N_36332);
and U42346 (N_42346,N_39620,N_39730);
nand U42347 (N_42347,N_38203,N_36282);
or U42348 (N_42348,N_38301,N_38091);
and U42349 (N_42349,N_35716,N_35140);
or U42350 (N_42350,N_37857,N_36907);
nand U42351 (N_42351,N_38779,N_35288);
or U42352 (N_42352,N_39720,N_36195);
nor U42353 (N_42353,N_39304,N_39763);
and U42354 (N_42354,N_39674,N_39765);
or U42355 (N_42355,N_35167,N_35549);
nor U42356 (N_42356,N_35358,N_39759);
xnor U42357 (N_42357,N_39042,N_39709);
xnor U42358 (N_42358,N_36310,N_38675);
nand U42359 (N_42359,N_38608,N_38111);
nor U42360 (N_42360,N_39827,N_37955);
or U42361 (N_42361,N_35708,N_36017);
or U42362 (N_42362,N_39966,N_35836);
or U42363 (N_42363,N_38287,N_36626);
xor U42364 (N_42364,N_37153,N_37595);
and U42365 (N_42365,N_36055,N_37825);
nor U42366 (N_42366,N_35969,N_37069);
xor U42367 (N_42367,N_37850,N_39019);
nor U42368 (N_42368,N_39993,N_38147);
or U42369 (N_42369,N_37648,N_38811);
nor U42370 (N_42370,N_36676,N_36381);
or U42371 (N_42371,N_39196,N_39326);
and U42372 (N_42372,N_37662,N_37021);
and U42373 (N_42373,N_36948,N_37799);
and U42374 (N_42374,N_35875,N_35814);
nor U42375 (N_42375,N_36902,N_36175);
and U42376 (N_42376,N_37452,N_35571);
nor U42377 (N_42377,N_36584,N_39743);
nor U42378 (N_42378,N_38406,N_35888);
and U42379 (N_42379,N_37872,N_37670);
and U42380 (N_42380,N_35158,N_37245);
nand U42381 (N_42381,N_38571,N_38724);
nand U42382 (N_42382,N_37220,N_36663);
xnor U42383 (N_42383,N_39374,N_39560);
xnor U42384 (N_42384,N_37737,N_38286);
or U42385 (N_42385,N_36319,N_37065);
and U42386 (N_42386,N_37681,N_39876);
or U42387 (N_42387,N_37588,N_38953);
and U42388 (N_42388,N_35037,N_37104);
nand U42389 (N_42389,N_36613,N_35748);
and U42390 (N_42390,N_39708,N_35785);
and U42391 (N_42391,N_39789,N_35700);
nand U42392 (N_42392,N_36727,N_38344);
or U42393 (N_42393,N_35311,N_35818);
nand U42394 (N_42394,N_37789,N_39156);
nor U42395 (N_42395,N_38201,N_35736);
nor U42396 (N_42396,N_39349,N_35509);
nand U42397 (N_42397,N_35538,N_38381);
or U42398 (N_42398,N_36520,N_38053);
and U42399 (N_42399,N_36971,N_36411);
or U42400 (N_42400,N_36137,N_38509);
or U42401 (N_42401,N_38451,N_38317);
nand U42402 (N_42402,N_35151,N_36910);
xnor U42403 (N_42403,N_39169,N_38660);
nand U42404 (N_42404,N_36623,N_37501);
and U42405 (N_42405,N_37655,N_37707);
xor U42406 (N_42406,N_36207,N_39411);
and U42407 (N_42407,N_35847,N_35559);
or U42408 (N_42408,N_39787,N_39996);
xor U42409 (N_42409,N_36117,N_38153);
and U42410 (N_42410,N_37221,N_37014);
xnor U42411 (N_42411,N_35636,N_36275);
nor U42412 (N_42412,N_35395,N_36439);
xnor U42413 (N_42413,N_37760,N_39343);
xor U42414 (N_42414,N_37790,N_37559);
xor U42415 (N_42415,N_38274,N_36847);
or U42416 (N_42416,N_35216,N_35413);
or U42417 (N_42417,N_35665,N_35258);
xor U42418 (N_42418,N_39231,N_38569);
or U42419 (N_42419,N_37634,N_36251);
and U42420 (N_42420,N_36328,N_35698);
xor U42421 (N_42421,N_36088,N_36665);
or U42422 (N_42422,N_38979,N_38885);
xor U42423 (N_42423,N_38098,N_36685);
nand U42424 (N_42424,N_39591,N_38284);
nand U42425 (N_42425,N_39327,N_38924);
and U42426 (N_42426,N_35683,N_36429);
xnor U42427 (N_42427,N_37903,N_39236);
and U42428 (N_42428,N_36957,N_39417);
xor U42429 (N_42429,N_36131,N_35264);
or U42430 (N_42430,N_39459,N_38186);
or U42431 (N_42431,N_38246,N_36892);
and U42432 (N_42432,N_38792,N_38258);
nor U42433 (N_42433,N_37795,N_35117);
or U42434 (N_42434,N_38170,N_36145);
nand U42435 (N_42435,N_36199,N_39645);
nand U42436 (N_42436,N_38710,N_35807);
nor U42437 (N_42437,N_35318,N_35565);
or U42438 (N_42438,N_37699,N_37610);
nor U42439 (N_42439,N_37226,N_36755);
and U42440 (N_42440,N_37998,N_37416);
xor U42441 (N_42441,N_37997,N_38775);
nor U42442 (N_42442,N_38609,N_39224);
xnor U42443 (N_42443,N_37197,N_37726);
nor U42444 (N_42444,N_38171,N_36125);
and U42445 (N_42445,N_37322,N_35857);
or U42446 (N_42446,N_36347,N_36912);
or U42447 (N_42447,N_35945,N_39452);
nor U42448 (N_42448,N_35855,N_39342);
or U42449 (N_42449,N_38884,N_35497);
nor U42450 (N_42450,N_39364,N_38458);
and U42451 (N_42451,N_38517,N_36406);
xnor U42452 (N_42452,N_37185,N_36893);
and U42453 (N_42453,N_35280,N_35999);
xnor U42454 (N_42454,N_39314,N_38060);
nand U42455 (N_42455,N_37406,N_36363);
xor U42456 (N_42456,N_35156,N_39940);
and U42457 (N_42457,N_37035,N_37597);
and U42458 (N_42458,N_39679,N_38032);
or U42459 (N_42459,N_35618,N_37683);
nand U42460 (N_42460,N_38271,N_36152);
or U42461 (N_42461,N_35682,N_35837);
xnor U42462 (N_42462,N_36908,N_39791);
and U42463 (N_42463,N_36505,N_37614);
nand U42464 (N_42464,N_36387,N_36530);
nand U42465 (N_42465,N_39005,N_35004);
and U42466 (N_42466,N_35874,N_36045);
nor U42467 (N_42467,N_36920,N_37088);
nor U42468 (N_42468,N_38449,N_35308);
xor U42469 (N_42469,N_37347,N_38055);
nor U42470 (N_42470,N_37645,N_35397);
nand U42471 (N_42471,N_36163,N_39463);
nor U42472 (N_42472,N_38342,N_39124);
nand U42473 (N_42473,N_39163,N_35385);
nor U42474 (N_42474,N_36173,N_38510);
nand U42475 (N_42475,N_37759,N_37386);
and U42476 (N_42476,N_38310,N_35584);
and U42477 (N_42477,N_35423,N_35406);
nor U42478 (N_42478,N_39510,N_38268);
nor U42479 (N_42479,N_37323,N_39110);
and U42480 (N_42480,N_35745,N_36403);
and U42481 (N_42481,N_35370,N_39097);
nor U42482 (N_42482,N_38915,N_36208);
xnor U42483 (N_42483,N_37519,N_35767);
nand U42484 (N_42484,N_36790,N_37741);
xnor U42485 (N_42485,N_38853,N_39166);
and U42486 (N_42486,N_39367,N_39356);
nor U42487 (N_42487,N_37250,N_38270);
or U42488 (N_42488,N_38292,N_35108);
xnor U42489 (N_42489,N_36679,N_39072);
nor U42490 (N_42490,N_36278,N_37083);
nor U42491 (N_42491,N_36706,N_39226);
xnor U42492 (N_42492,N_37766,N_37818);
and U42493 (N_42493,N_39908,N_37703);
or U42494 (N_42494,N_39500,N_35544);
nand U42495 (N_42495,N_36654,N_38747);
nor U42496 (N_42496,N_35247,N_38584);
and U42497 (N_42497,N_38622,N_36423);
or U42498 (N_42498,N_35064,N_35661);
nor U42499 (N_42499,N_37159,N_35145);
xor U42500 (N_42500,N_39016,N_36260);
or U42501 (N_42501,N_39333,N_38238);
and U42502 (N_42502,N_36210,N_38592);
or U42503 (N_42503,N_39061,N_36905);
and U42504 (N_42504,N_39538,N_37345);
nand U42505 (N_42505,N_37550,N_38813);
or U42506 (N_42506,N_36293,N_38451);
or U42507 (N_42507,N_37593,N_39061);
xnor U42508 (N_42508,N_35337,N_39297);
or U42509 (N_42509,N_36858,N_39460);
nand U42510 (N_42510,N_38449,N_35916);
nand U42511 (N_42511,N_36562,N_36613);
and U42512 (N_42512,N_35623,N_39714);
or U42513 (N_42513,N_38314,N_35280);
nand U42514 (N_42514,N_35509,N_35909);
or U42515 (N_42515,N_36005,N_37544);
or U42516 (N_42516,N_38238,N_36332);
nand U42517 (N_42517,N_37115,N_37183);
or U42518 (N_42518,N_35873,N_38145);
nor U42519 (N_42519,N_36802,N_37323);
and U42520 (N_42520,N_37337,N_38747);
xnor U42521 (N_42521,N_38300,N_37165);
or U42522 (N_42522,N_37611,N_38415);
nor U42523 (N_42523,N_35542,N_36898);
nor U42524 (N_42524,N_39438,N_36137);
xor U42525 (N_42525,N_39438,N_39473);
and U42526 (N_42526,N_35209,N_36737);
nand U42527 (N_42527,N_35244,N_35877);
and U42528 (N_42528,N_38195,N_36437);
xor U42529 (N_42529,N_39316,N_37442);
and U42530 (N_42530,N_38238,N_38421);
xor U42531 (N_42531,N_39143,N_38630);
nor U42532 (N_42532,N_36257,N_36949);
nand U42533 (N_42533,N_37406,N_37713);
or U42534 (N_42534,N_39223,N_38106);
and U42535 (N_42535,N_39608,N_39317);
or U42536 (N_42536,N_38345,N_36633);
nand U42537 (N_42537,N_36868,N_39520);
or U42538 (N_42538,N_39107,N_35883);
nor U42539 (N_42539,N_35272,N_38013);
or U42540 (N_42540,N_36882,N_38860);
nor U42541 (N_42541,N_37964,N_36320);
nand U42542 (N_42542,N_39847,N_36421);
and U42543 (N_42543,N_39878,N_38163);
nor U42544 (N_42544,N_38850,N_37280);
and U42545 (N_42545,N_35047,N_39757);
xor U42546 (N_42546,N_37003,N_39785);
nand U42547 (N_42547,N_39486,N_36211);
nor U42548 (N_42548,N_37594,N_37712);
nor U42549 (N_42549,N_35737,N_38566);
xor U42550 (N_42550,N_36007,N_39556);
and U42551 (N_42551,N_36661,N_35973);
nand U42552 (N_42552,N_35090,N_36218);
nand U42553 (N_42553,N_38603,N_39669);
nor U42554 (N_42554,N_39683,N_35333);
xor U42555 (N_42555,N_38030,N_35532);
and U42556 (N_42556,N_36577,N_37493);
and U42557 (N_42557,N_38746,N_38439);
or U42558 (N_42558,N_37680,N_39462);
xnor U42559 (N_42559,N_35650,N_38998);
or U42560 (N_42560,N_39725,N_37983);
nor U42561 (N_42561,N_37533,N_36285);
and U42562 (N_42562,N_39884,N_39970);
or U42563 (N_42563,N_38820,N_37914);
and U42564 (N_42564,N_38522,N_36028);
or U42565 (N_42565,N_37533,N_39861);
nand U42566 (N_42566,N_35039,N_35036);
or U42567 (N_42567,N_39986,N_36909);
nor U42568 (N_42568,N_35101,N_37964);
and U42569 (N_42569,N_35624,N_39169);
nand U42570 (N_42570,N_39312,N_38967);
nor U42571 (N_42571,N_39052,N_36016);
nand U42572 (N_42572,N_39094,N_39978);
nand U42573 (N_42573,N_36164,N_38385);
xnor U42574 (N_42574,N_39347,N_38515);
and U42575 (N_42575,N_36921,N_36479);
or U42576 (N_42576,N_39179,N_36540);
nand U42577 (N_42577,N_39270,N_35674);
nand U42578 (N_42578,N_39545,N_37742);
or U42579 (N_42579,N_39467,N_39771);
xnor U42580 (N_42580,N_38558,N_39952);
nor U42581 (N_42581,N_35748,N_37775);
xnor U42582 (N_42582,N_35100,N_36049);
nand U42583 (N_42583,N_37377,N_39849);
or U42584 (N_42584,N_36711,N_36375);
xor U42585 (N_42585,N_39621,N_35281);
or U42586 (N_42586,N_38882,N_37575);
nand U42587 (N_42587,N_39562,N_37549);
xnor U42588 (N_42588,N_38558,N_36916);
or U42589 (N_42589,N_35757,N_37078);
nor U42590 (N_42590,N_37372,N_37283);
and U42591 (N_42591,N_35928,N_39686);
nand U42592 (N_42592,N_36116,N_37466);
nand U42593 (N_42593,N_38061,N_37359);
xor U42594 (N_42594,N_37504,N_35788);
nand U42595 (N_42595,N_38088,N_37741);
xnor U42596 (N_42596,N_36587,N_38177);
nand U42597 (N_42597,N_36328,N_39122);
or U42598 (N_42598,N_35794,N_39031);
nor U42599 (N_42599,N_38306,N_37754);
nor U42600 (N_42600,N_38474,N_39886);
or U42601 (N_42601,N_39616,N_37913);
nor U42602 (N_42602,N_36849,N_38566);
nor U42603 (N_42603,N_39168,N_39733);
nand U42604 (N_42604,N_38327,N_37552);
and U42605 (N_42605,N_36209,N_37844);
and U42606 (N_42606,N_37322,N_35679);
nand U42607 (N_42607,N_35638,N_37254);
or U42608 (N_42608,N_38533,N_36535);
nand U42609 (N_42609,N_38743,N_38092);
or U42610 (N_42610,N_36396,N_35531);
xor U42611 (N_42611,N_38281,N_35336);
or U42612 (N_42612,N_36352,N_35436);
xnor U42613 (N_42613,N_35781,N_36302);
nand U42614 (N_42614,N_36428,N_36609);
xor U42615 (N_42615,N_35629,N_38754);
or U42616 (N_42616,N_37087,N_37261);
and U42617 (N_42617,N_35187,N_36475);
xor U42618 (N_42618,N_39306,N_35727);
nand U42619 (N_42619,N_39004,N_38228);
or U42620 (N_42620,N_35183,N_38087);
nor U42621 (N_42621,N_38028,N_37684);
nand U42622 (N_42622,N_35555,N_35240);
nor U42623 (N_42623,N_36990,N_36763);
nor U42624 (N_42624,N_39780,N_38945);
and U42625 (N_42625,N_36795,N_36229);
nor U42626 (N_42626,N_37470,N_38024);
xnor U42627 (N_42627,N_38965,N_37998);
or U42628 (N_42628,N_39512,N_38633);
xor U42629 (N_42629,N_38693,N_36113);
nand U42630 (N_42630,N_35548,N_37376);
nand U42631 (N_42631,N_36065,N_36093);
nor U42632 (N_42632,N_35842,N_36706);
nor U42633 (N_42633,N_38853,N_39480);
xor U42634 (N_42634,N_36410,N_37847);
nand U42635 (N_42635,N_35313,N_35099);
nor U42636 (N_42636,N_38532,N_36415);
nand U42637 (N_42637,N_36260,N_35030);
and U42638 (N_42638,N_37782,N_39692);
nand U42639 (N_42639,N_39862,N_38488);
nand U42640 (N_42640,N_35986,N_36476);
nand U42641 (N_42641,N_37583,N_37705);
nand U42642 (N_42642,N_38306,N_38922);
nand U42643 (N_42643,N_39263,N_38892);
xnor U42644 (N_42644,N_37162,N_38686);
xor U42645 (N_42645,N_38193,N_38301);
and U42646 (N_42646,N_36317,N_35927);
and U42647 (N_42647,N_37872,N_35820);
nor U42648 (N_42648,N_36253,N_36887);
nor U42649 (N_42649,N_35471,N_37515);
or U42650 (N_42650,N_35436,N_36881);
nand U42651 (N_42651,N_35299,N_37844);
and U42652 (N_42652,N_35243,N_37075);
xnor U42653 (N_42653,N_35135,N_36667);
nor U42654 (N_42654,N_39248,N_38549);
nand U42655 (N_42655,N_37214,N_35921);
xnor U42656 (N_42656,N_35614,N_36435);
or U42657 (N_42657,N_39277,N_39596);
xnor U42658 (N_42658,N_36728,N_35258);
nor U42659 (N_42659,N_37955,N_39794);
nor U42660 (N_42660,N_36453,N_37072);
and U42661 (N_42661,N_37483,N_37721);
and U42662 (N_42662,N_35800,N_37941);
nand U42663 (N_42663,N_35063,N_39157);
nand U42664 (N_42664,N_39359,N_38138);
xor U42665 (N_42665,N_35553,N_39173);
or U42666 (N_42666,N_37753,N_39124);
xor U42667 (N_42667,N_38216,N_39501);
nor U42668 (N_42668,N_38958,N_39921);
nor U42669 (N_42669,N_36974,N_39446);
and U42670 (N_42670,N_37101,N_37261);
and U42671 (N_42671,N_37888,N_36376);
nand U42672 (N_42672,N_38229,N_35033);
nor U42673 (N_42673,N_37137,N_38650);
xor U42674 (N_42674,N_35795,N_35278);
nor U42675 (N_42675,N_35295,N_35046);
nand U42676 (N_42676,N_37857,N_36511);
xor U42677 (N_42677,N_35786,N_38481);
xnor U42678 (N_42678,N_36487,N_38201);
nand U42679 (N_42679,N_39195,N_37725);
nor U42680 (N_42680,N_35918,N_35316);
nor U42681 (N_42681,N_38015,N_38901);
and U42682 (N_42682,N_37801,N_36649);
nand U42683 (N_42683,N_37532,N_38303);
or U42684 (N_42684,N_38773,N_38248);
or U42685 (N_42685,N_36620,N_38790);
xor U42686 (N_42686,N_35628,N_38612);
and U42687 (N_42687,N_37659,N_36968);
nand U42688 (N_42688,N_35975,N_37348);
or U42689 (N_42689,N_39445,N_38384);
nand U42690 (N_42690,N_36825,N_37806);
and U42691 (N_42691,N_36105,N_37071);
or U42692 (N_42692,N_37689,N_38580);
and U42693 (N_42693,N_35747,N_38113);
nor U42694 (N_42694,N_39871,N_38152);
nand U42695 (N_42695,N_38431,N_36403);
xor U42696 (N_42696,N_37827,N_39714);
or U42697 (N_42697,N_35817,N_35669);
xor U42698 (N_42698,N_35964,N_39458);
and U42699 (N_42699,N_36598,N_36919);
or U42700 (N_42700,N_37267,N_38003);
nor U42701 (N_42701,N_39103,N_35023);
xnor U42702 (N_42702,N_35174,N_37439);
and U42703 (N_42703,N_37594,N_37959);
or U42704 (N_42704,N_35478,N_37768);
or U42705 (N_42705,N_38601,N_35259);
xor U42706 (N_42706,N_37613,N_37188);
and U42707 (N_42707,N_36288,N_39954);
xnor U42708 (N_42708,N_38727,N_38748);
nand U42709 (N_42709,N_39174,N_35061);
and U42710 (N_42710,N_37823,N_35573);
and U42711 (N_42711,N_35122,N_36267);
and U42712 (N_42712,N_37770,N_38302);
and U42713 (N_42713,N_35718,N_36212);
and U42714 (N_42714,N_35248,N_37469);
xor U42715 (N_42715,N_38038,N_38477);
or U42716 (N_42716,N_38878,N_36107);
nand U42717 (N_42717,N_36546,N_38194);
nor U42718 (N_42718,N_35915,N_35079);
nor U42719 (N_42719,N_36931,N_39407);
nor U42720 (N_42720,N_37381,N_38146);
and U42721 (N_42721,N_38864,N_38964);
nand U42722 (N_42722,N_39566,N_35045);
xnor U42723 (N_42723,N_38536,N_36196);
xor U42724 (N_42724,N_36496,N_35963);
and U42725 (N_42725,N_35312,N_39307);
xor U42726 (N_42726,N_36770,N_39686);
nor U42727 (N_42727,N_35701,N_39497);
nand U42728 (N_42728,N_36519,N_36690);
or U42729 (N_42729,N_39101,N_39123);
nor U42730 (N_42730,N_37247,N_37091);
and U42731 (N_42731,N_35384,N_37201);
nand U42732 (N_42732,N_35175,N_38415);
nor U42733 (N_42733,N_36429,N_37432);
nand U42734 (N_42734,N_38483,N_39004);
nor U42735 (N_42735,N_38095,N_35677);
nand U42736 (N_42736,N_39926,N_38722);
and U42737 (N_42737,N_36458,N_38000);
nand U42738 (N_42738,N_35075,N_39808);
and U42739 (N_42739,N_36847,N_35428);
and U42740 (N_42740,N_36616,N_36654);
xor U42741 (N_42741,N_39799,N_36250);
and U42742 (N_42742,N_37703,N_39627);
and U42743 (N_42743,N_36644,N_38090);
or U42744 (N_42744,N_36465,N_37089);
or U42745 (N_42745,N_39199,N_36518);
or U42746 (N_42746,N_35884,N_39037);
nand U42747 (N_42747,N_39006,N_35211);
and U42748 (N_42748,N_39743,N_35775);
and U42749 (N_42749,N_36880,N_36067);
nor U42750 (N_42750,N_35793,N_39747);
nor U42751 (N_42751,N_38693,N_35981);
nand U42752 (N_42752,N_39064,N_35897);
nand U42753 (N_42753,N_38632,N_38261);
nor U42754 (N_42754,N_35298,N_35124);
nand U42755 (N_42755,N_35553,N_39694);
or U42756 (N_42756,N_36155,N_37709);
xnor U42757 (N_42757,N_36267,N_35643);
nor U42758 (N_42758,N_36715,N_35222);
or U42759 (N_42759,N_39094,N_37097);
and U42760 (N_42760,N_38893,N_36124);
or U42761 (N_42761,N_39151,N_35756);
xor U42762 (N_42762,N_37460,N_38244);
nor U42763 (N_42763,N_35305,N_37453);
and U42764 (N_42764,N_39819,N_39790);
xor U42765 (N_42765,N_38661,N_38103);
nor U42766 (N_42766,N_39060,N_36973);
nor U42767 (N_42767,N_38719,N_35130);
nand U42768 (N_42768,N_36161,N_37064);
and U42769 (N_42769,N_38184,N_38198);
nor U42770 (N_42770,N_36487,N_37454);
and U42771 (N_42771,N_39347,N_38550);
xnor U42772 (N_42772,N_37538,N_37670);
xnor U42773 (N_42773,N_38390,N_37690);
and U42774 (N_42774,N_37023,N_36114);
and U42775 (N_42775,N_37194,N_36234);
xnor U42776 (N_42776,N_38445,N_37475);
nor U42777 (N_42777,N_36893,N_39161);
or U42778 (N_42778,N_37101,N_36525);
nor U42779 (N_42779,N_38509,N_35618);
nand U42780 (N_42780,N_38325,N_37082);
nor U42781 (N_42781,N_35079,N_36337);
nor U42782 (N_42782,N_35457,N_35651);
and U42783 (N_42783,N_35197,N_35064);
nand U42784 (N_42784,N_37452,N_35912);
nor U42785 (N_42785,N_35087,N_39507);
nand U42786 (N_42786,N_39506,N_38794);
or U42787 (N_42787,N_36783,N_36821);
nand U42788 (N_42788,N_37856,N_35141);
or U42789 (N_42789,N_39655,N_39113);
and U42790 (N_42790,N_35009,N_38434);
xor U42791 (N_42791,N_38617,N_39460);
xor U42792 (N_42792,N_35104,N_39486);
nor U42793 (N_42793,N_36316,N_38449);
nor U42794 (N_42794,N_37066,N_36057);
nand U42795 (N_42795,N_39094,N_35253);
xnor U42796 (N_42796,N_35821,N_35742);
nand U42797 (N_42797,N_39692,N_39736);
or U42798 (N_42798,N_35148,N_38238);
nor U42799 (N_42799,N_38256,N_39808);
nand U42800 (N_42800,N_36600,N_36474);
xor U42801 (N_42801,N_36831,N_39205);
xnor U42802 (N_42802,N_36183,N_36513);
nor U42803 (N_42803,N_37571,N_35850);
or U42804 (N_42804,N_39619,N_38159);
nand U42805 (N_42805,N_36004,N_38582);
xor U42806 (N_42806,N_38752,N_39459);
xor U42807 (N_42807,N_38058,N_38988);
xnor U42808 (N_42808,N_39247,N_38664);
nor U42809 (N_42809,N_36214,N_37497);
nor U42810 (N_42810,N_35240,N_39874);
nand U42811 (N_42811,N_38814,N_35328);
nor U42812 (N_42812,N_36866,N_38263);
nand U42813 (N_42813,N_39932,N_38092);
and U42814 (N_42814,N_37096,N_35478);
nand U42815 (N_42815,N_39819,N_37201);
nor U42816 (N_42816,N_35597,N_38939);
nand U42817 (N_42817,N_38855,N_37841);
or U42818 (N_42818,N_38092,N_35687);
xnor U42819 (N_42819,N_36118,N_37408);
or U42820 (N_42820,N_39175,N_36861);
and U42821 (N_42821,N_36304,N_39186);
xnor U42822 (N_42822,N_36981,N_35045);
xor U42823 (N_42823,N_35231,N_36084);
nor U42824 (N_42824,N_37548,N_35242);
and U42825 (N_42825,N_39731,N_35317);
and U42826 (N_42826,N_38301,N_39171);
or U42827 (N_42827,N_37746,N_38199);
nand U42828 (N_42828,N_36587,N_39287);
nand U42829 (N_42829,N_39516,N_35471);
nor U42830 (N_42830,N_36472,N_37106);
nand U42831 (N_42831,N_37788,N_36636);
nor U42832 (N_42832,N_39190,N_39611);
nand U42833 (N_42833,N_38330,N_38846);
and U42834 (N_42834,N_37990,N_36898);
xor U42835 (N_42835,N_38095,N_37783);
and U42836 (N_42836,N_38124,N_38667);
nor U42837 (N_42837,N_38742,N_37278);
nor U42838 (N_42838,N_36426,N_35120);
or U42839 (N_42839,N_38975,N_38295);
and U42840 (N_42840,N_35328,N_35635);
xnor U42841 (N_42841,N_38209,N_39667);
or U42842 (N_42842,N_36660,N_39511);
or U42843 (N_42843,N_37730,N_36200);
xnor U42844 (N_42844,N_35956,N_36857);
or U42845 (N_42845,N_38263,N_38099);
nand U42846 (N_42846,N_38593,N_37846);
nand U42847 (N_42847,N_36945,N_35614);
nor U42848 (N_42848,N_35339,N_36895);
xnor U42849 (N_42849,N_39736,N_37338);
and U42850 (N_42850,N_35690,N_38238);
nor U42851 (N_42851,N_35583,N_39637);
or U42852 (N_42852,N_38574,N_39082);
xor U42853 (N_42853,N_37491,N_36526);
xnor U42854 (N_42854,N_39331,N_36321);
or U42855 (N_42855,N_36146,N_35190);
nand U42856 (N_42856,N_39028,N_35303);
nor U42857 (N_42857,N_36583,N_38756);
or U42858 (N_42858,N_36862,N_37702);
and U42859 (N_42859,N_36174,N_36733);
or U42860 (N_42860,N_38014,N_37549);
nand U42861 (N_42861,N_37679,N_37087);
nand U42862 (N_42862,N_35351,N_39927);
and U42863 (N_42863,N_35925,N_39798);
nor U42864 (N_42864,N_38956,N_37752);
or U42865 (N_42865,N_36092,N_38042);
or U42866 (N_42866,N_35635,N_35335);
nor U42867 (N_42867,N_38358,N_39193);
xor U42868 (N_42868,N_35765,N_39444);
xnor U42869 (N_42869,N_36258,N_36106);
or U42870 (N_42870,N_39229,N_35990);
and U42871 (N_42871,N_39072,N_36492);
or U42872 (N_42872,N_35939,N_35221);
or U42873 (N_42873,N_35384,N_38755);
and U42874 (N_42874,N_36780,N_36225);
or U42875 (N_42875,N_37046,N_37203);
and U42876 (N_42876,N_39670,N_35875);
xnor U42877 (N_42877,N_35023,N_37975);
nor U42878 (N_42878,N_38575,N_37724);
nand U42879 (N_42879,N_36554,N_37013);
xnor U42880 (N_42880,N_35283,N_35042);
nor U42881 (N_42881,N_37667,N_39569);
xor U42882 (N_42882,N_36975,N_36778);
and U42883 (N_42883,N_38657,N_38488);
xnor U42884 (N_42884,N_35820,N_39523);
or U42885 (N_42885,N_36642,N_36158);
nor U42886 (N_42886,N_36193,N_35215);
and U42887 (N_42887,N_38943,N_39078);
nand U42888 (N_42888,N_36925,N_38035);
nand U42889 (N_42889,N_39647,N_36051);
nand U42890 (N_42890,N_36541,N_39893);
and U42891 (N_42891,N_38779,N_36944);
or U42892 (N_42892,N_36950,N_35237);
and U42893 (N_42893,N_39605,N_35685);
and U42894 (N_42894,N_35916,N_37995);
and U42895 (N_42895,N_37708,N_36221);
xnor U42896 (N_42896,N_39591,N_35877);
nor U42897 (N_42897,N_35899,N_35587);
nor U42898 (N_42898,N_37580,N_38983);
xnor U42899 (N_42899,N_37695,N_37448);
nor U42900 (N_42900,N_37913,N_38364);
xor U42901 (N_42901,N_38998,N_38248);
and U42902 (N_42902,N_38600,N_39650);
nand U42903 (N_42903,N_37984,N_37699);
xor U42904 (N_42904,N_36746,N_38722);
xor U42905 (N_42905,N_35880,N_36805);
nor U42906 (N_42906,N_35211,N_35856);
and U42907 (N_42907,N_36097,N_39843);
and U42908 (N_42908,N_36957,N_35570);
and U42909 (N_42909,N_39992,N_38534);
nand U42910 (N_42910,N_35312,N_39929);
or U42911 (N_42911,N_35844,N_36015);
or U42912 (N_42912,N_39014,N_38552);
or U42913 (N_42913,N_35508,N_39386);
nor U42914 (N_42914,N_39828,N_39125);
nor U42915 (N_42915,N_35470,N_36635);
nand U42916 (N_42916,N_39948,N_38265);
and U42917 (N_42917,N_38066,N_35642);
nor U42918 (N_42918,N_37707,N_36859);
nand U42919 (N_42919,N_38425,N_36865);
nand U42920 (N_42920,N_39226,N_36223);
and U42921 (N_42921,N_37029,N_37654);
nor U42922 (N_42922,N_38265,N_39653);
and U42923 (N_42923,N_37770,N_35171);
and U42924 (N_42924,N_39633,N_38694);
or U42925 (N_42925,N_35014,N_36011);
nand U42926 (N_42926,N_36281,N_37763);
xnor U42927 (N_42927,N_36079,N_36908);
nand U42928 (N_42928,N_36054,N_35943);
nor U42929 (N_42929,N_39454,N_37692);
xnor U42930 (N_42930,N_37799,N_35144);
or U42931 (N_42931,N_36598,N_39034);
or U42932 (N_42932,N_35523,N_37155);
or U42933 (N_42933,N_37836,N_39640);
nand U42934 (N_42934,N_36192,N_35879);
nand U42935 (N_42935,N_39428,N_36265);
or U42936 (N_42936,N_39968,N_36508);
and U42937 (N_42937,N_35862,N_39494);
or U42938 (N_42938,N_36879,N_38419);
or U42939 (N_42939,N_39318,N_39401);
xor U42940 (N_42940,N_39337,N_36999);
xor U42941 (N_42941,N_36660,N_38195);
xor U42942 (N_42942,N_39967,N_35154);
and U42943 (N_42943,N_38018,N_37583);
nand U42944 (N_42944,N_39112,N_39654);
xor U42945 (N_42945,N_35506,N_38417);
and U42946 (N_42946,N_38377,N_35375);
or U42947 (N_42947,N_39331,N_36718);
and U42948 (N_42948,N_35688,N_39675);
xor U42949 (N_42949,N_39698,N_35221);
and U42950 (N_42950,N_38946,N_37671);
and U42951 (N_42951,N_38536,N_39935);
and U42952 (N_42952,N_35672,N_36580);
nor U42953 (N_42953,N_37067,N_38203);
and U42954 (N_42954,N_38670,N_37986);
nor U42955 (N_42955,N_38945,N_37089);
or U42956 (N_42956,N_37871,N_36704);
or U42957 (N_42957,N_36873,N_36070);
or U42958 (N_42958,N_36069,N_35330);
or U42959 (N_42959,N_37117,N_36349);
nor U42960 (N_42960,N_38178,N_37228);
and U42961 (N_42961,N_36622,N_39597);
nand U42962 (N_42962,N_38202,N_38442);
and U42963 (N_42963,N_36393,N_39118);
nand U42964 (N_42964,N_39030,N_35453);
and U42965 (N_42965,N_39498,N_39167);
nor U42966 (N_42966,N_37015,N_37243);
xor U42967 (N_42967,N_39628,N_35941);
nor U42968 (N_42968,N_37234,N_37873);
nor U42969 (N_42969,N_37118,N_38366);
or U42970 (N_42970,N_39248,N_37098);
xor U42971 (N_42971,N_36635,N_38139);
and U42972 (N_42972,N_38994,N_37019);
and U42973 (N_42973,N_39356,N_39631);
and U42974 (N_42974,N_37911,N_35003);
xnor U42975 (N_42975,N_38000,N_36503);
nand U42976 (N_42976,N_36032,N_39718);
nand U42977 (N_42977,N_37525,N_39011);
nor U42978 (N_42978,N_37464,N_36211);
nand U42979 (N_42979,N_39694,N_37728);
or U42980 (N_42980,N_39069,N_35136);
nand U42981 (N_42981,N_37716,N_36908);
nor U42982 (N_42982,N_39492,N_38949);
and U42983 (N_42983,N_36870,N_38007);
xnor U42984 (N_42984,N_37432,N_39162);
and U42985 (N_42985,N_36091,N_36415);
xor U42986 (N_42986,N_38747,N_36817);
and U42987 (N_42987,N_39100,N_36199);
nand U42988 (N_42988,N_36558,N_39220);
and U42989 (N_42989,N_38729,N_36479);
and U42990 (N_42990,N_38253,N_38680);
and U42991 (N_42991,N_39039,N_38347);
nand U42992 (N_42992,N_36514,N_37642);
nand U42993 (N_42993,N_36684,N_38046);
nor U42994 (N_42994,N_38777,N_35339);
xor U42995 (N_42995,N_38546,N_39906);
xnor U42996 (N_42996,N_35608,N_37887);
nor U42997 (N_42997,N_35959,N_39573);
nor U42998 (N_42998,N_35485,N_39944);
nor U42999 (N_42999,N_39965,N_36530);
nand U43000 (N_43000,N_36449,N_36593);
xnor U43001 (N_43001,N_35171,N_37438);
nor U43002 (N_43002,N_39153,N_36205);
nand U43003 (N_43003,N_38743,N_36087);
nor U43004 (N_43004,N_39922,N_38098);
or U43005 (N_43005,N_39150,N_39434);
nand U43006 (N_43006,N_37509,N_36584);
nor U43007 (N_43007,N_39440,N_38647);
or U43008 (N_43008,N_39761,N_35881);
nor U43009 (N_43009,N_39002,N_36609);
or U43010 (N_43010,N_36096,N_36664);
or U43011 (N_43011,N_35725,N_39104);
nor U43012 (N_43012,N_35624,N_36799);
nor U43013 (N_43013,N_37866,N_36374);
xor U43014 (N_43014,N_35910,N_35378);
and U43015 (N_43015,N_35184,N_37968);
nor U43016 (N_43016,N_35379,N_37818);
or U43017 (N_43017,N_36679,N_36331);
or U43018 (N_43018,N_35344,N_38110);
or U43019 (N_43019,N_35043,N_38399);
nand U43020 (N_43020,N_38881,N_35109);
xor U43021 (N_43021,N_38791,N_39550);
and U43022 (N_43022,N_35174,N_37512);
xnor U43023 (N_43023,N_38442,N_38464);
and U43024 (N_43024,N_37492,N_35732);
nand U43025 (N_43025,N_35126,N_36118);
and U43026 (N_43026,N_39051,N_38667);
or U43027 (N_43027,N_39881,N_38312);
nand U43028 (N_43028,N_35743,N_35545);
nor U43029 (N_43029,N_35988,N_37913);
nor U43030 (N_43030,N_38888,N_36126);
nor U43031 (N_43031,N_37936,N_38862);
nor U43032 (N_43032,N_37466,N_37622);
xnor U43033 (N_43033,N_36681,N_39995);
nand U43034 (N_43034,N_36811,N_37282);
and U43035 (N_43035,N_37361,N_35602);
and U43036 (N_43036,N_37619,N_38494);
and U43037 (N_43037,N_35888,N_36078);
nor U43038 (N_43038,N_39742,N_35876);
xor U43039 (N_43039,N_35214,N_39837);
nor U43040 (N_43040,N_35618,N_36096);
or U43041 (N_43041,N_36750,N_35717);
nand U43042 (N_43042,N_36622,N_37392);
xor U43043 (N_43043,N_35869,N_36039);
nand U43044 (N_43044,N_39378,N_36294);
nand U43045 (N_43045,N_38844,N_38768);
and U43046 (N_43046,N_37858,N_36280);
nor U43047 (N_43047,N_38217,N_35173);
nand U43048 (N_43048,N_38730,N_35469);
nor U43049 (N_43049,N_37366,N_39467);
nand U43050 (N_43050,N_38452,N_35013);
or U43051 (N_43051,N_37750,N_37938);
xor U43052 (N_43052,N_36963,N_36198);
nand U43053 (N_43053,N_35735,N_37067);
and U43054 (N_43054,N_36397,N_36368);
nand U43055 (N_43055,N_38699,N_36844);
nand U43056 (N_43056,N_37620,N_38057);
nand U43057 (N_43057,N_37717,N_37872);
xor U43058 (N_43058,N_38293,N_35802);
and U43059 (N_43059,N_35790,N_38048);
nor U43060 (N_43060,N_35071,N_37114);
xor U43061 (N_43061,N_38927,N_37266);
or U43062 (N_43062,N_37036,N_35907);
nor U43063 (N_43063,N_35437,N_35621);
nor U43064 (N_43064,N_39503,N_35664);
xor U43065 (N_43065,N_39611,N_36961);
xnor U43066 (N_43066,N_37410,N_36923);
nor U43067 (N_43067,N_38148,N_36565);
or U43068 (N_43068,N_37952,N_39407);
xor U43069 (N_43069,N_35970,N_35506);
and U43070 (N_43070,N_36231,N_39657);
nor U43071 (N_43071,N_35919,N_35472);
nor U43072 (N_43072,N_35582,N_38043);
nand U43073 (N_43073,N_35281,N_37818);
and U43074 (N_43074,N_38620,N_37113);
and U43075 (N_43075,N_38525,N_38927);
nor U43076 (N_43076,N_37867,N_39648);
nor U43077 (N_43077,N_38681,N_35817);
or U43078 (N_43078,N_38731,N_35243);
nand U43079 (N_43079,N_39306,N_36637);
xnor U43080 (N_43080,N_36119,N_36936);
xor U43081 (N_43081,N_37734,N_37499);
nor U43082 (N_43082,N_38298,N_36872);
and U43083 (N_43083,N_35712,N_37347);
nand U43084 (N_43084,N_37636,N_36163);
nor U43085 (N_43085,N_38552,N_37261);
xor U43086 (N_43086,N_35816,N_39696);
nor U43087 (N_43087,N_39806,N_39343);
or U43088 (N_43088,N_36597,N_37792);
xor U43089 (N_43089,N_39216,N_37837);
nor U43090 (N_43090,N_37069,N_36176);
nand U43091 (N_43091,N_38332,N_38865);
xnor U43092 (N_43092,N_35174,N_36302);
nand U43093 (N_43093,N_35694,N_39448);
xor U43094 (N_43094,N_38500,N_35280);
xnor U43095 (N_43095,N_38386,N_36925);
nand U43096 (N_43096,N_37156,N_38567);
and U43097 (N_43097,N_38347,N_38056);
nand U43098 (N_43098,N_37258,N_36628);
xor U43099 (N_43099,N_37320,N_37965);
nor U43100 (N_43100,N_36726,N_38760);
and U43101 (N_43101,N_36763,N_37144);
nor U43102 (N_43102,N_37601,N_36221);
xor U43103 (N_43103,N_38959,N_39199);
or U43104 (N_43104,N_38479,N_38555);
xor U43105 (N_43105,N_35104,N_38349);
xor U43106 (N_43106,N_38595,N_36673);
nand U43107 (N_43107,N_39585,N_37553);
or U43108 (N_43108,N_35328,N_38150);
and U43109 (N_43109,N_36456,N_38498);
or U43110 (N_43110,N_36646,N_38448);
nand U43111 (N_43111,N_38172,N_39192);
and U43112 (N_43112,N_35832,N_39224);
nand U43113 (N_43113,N_39288,N_37525);
nor U43114 (N_43114,N_38629,N_38911);
nand U43115 (N_43115,N_37853,N_35278);
nor U43116 (N_43116,N_36839,N_38898);
xor U43117 (N_43117,N_35914,N_37852);
and U43118 (N_43118,N_39082,N_39935);
nor U43119 (N_43119,N_38701,N_37837);
or U43120 (N_43120,N_39352,N_39975);
xnor U43121 (N_43121,N_36817,N_39200);
and U43122 (N_43122,N_37092,N_39709);
nand U43123 (N_43123,N_39205,N_38629);
and U43124 (N_43124,N_35430,N_39691);
or U43125 (N_43125,N_35342,N_36863);
nand U43126 (N_43126,N_37414,N_37680);
and U43127 (N_43127,N_36277,N_39476);
nand U43128 (N_43128,N_38707,N_39845);
xor U43129 (N_43129,N_35936,N_35615);
or U43130 (N_43130,N_36011,N_36440);
xnor U43131 (N_43131,N_39152,N_38420);
and U43132 (N_43132,N_35879,N_38339);
or U43133 (N_43133,N_38984,N_38288);
or U43134 (N_43134,N_36606,N_39755);
nor U43135 (N_43135,N_36968,N_36068);
or U43136 (N_43136,N_39116,N_35653);
or U43137 (N_43137,N_35290,N_35244);
and U43138 (N_43138,N_35056,N_39217);
nand U43139 (N_43139,N_37333,N_35369);
and U43140 (N_43140,N_39765,N_39785);
nor U43141 (N_43141,N_37272,N_36407);
nor U43142 (N_43142,N_39020,N_38512);
or U43143 (N_43143,N_36395,N_38459);
or U43144 (N_43144,N_37820,N_35431);
xor U43145 (N_43145,N_37160,N_36988);
and U43146 (N_43146,N_38595,N_36988);
nand U43147 (N_43147,N_36830,N_36404);
nand U43148 (N_43148,N_36138,N_37912);
nand U43149 (N_43149,N_39977,N_38565);
or U43150 (N_43150,N_36359,N_36835);
xor U43151 (N_43151,N_35361,N_39144);
and U43152 (N_43152,N_38208,N_35366);
nand U43153 (N_43153,N_36753,N_37335);
nand U43154 (N_43154,N_39695,N_36675);
and U43155 (N_43155,N_38141,N_38626);
nand U43156 (N_43156,N_37605,N_39524);
xnor U43157 (N_43157,N_37320,N_37312);
nor U43158 (N_43158,N_39732,N_36698);
or U43159 (N_43159,N_36401,N_35152);
or U43160 (N_43160,N_35281,N_35773);
xnor U43161 (N_43161,N_37352,N_35957);
or U43162 (N_43162,N_37985,N_36500);
xnor U43163 (N_43163,N_37383,N_39236);
xnor U43164 (N_43164,N_39523,N_38445);
nand U43165 (N_43165,N_35001,N_38752);
and U43166 (N_43166,N_37588,N_39039);
nor U43167 (N_43167,N_38166,N_39960);
nor U43168 (N_43168,N_35017,N_38449);
nor U43169 (N_43169,N_39541,N_37180);
and U43170 (N_43170,N_35648,N_35465);
or U43171 (N_43171,N_35746,N_36742);
or U43172 (N_43172,N_35424,N_36655);
nand U43173 (N_43173,N_35651,N_38672);
xnor U43174 (N_43174,N_39675,N_39242);
and U43175 (N_43175,N_36112,N_36679);
and U43176 (N_43176,N_36590,N_36949);
nor U43177 (N_43177,N_37131,N_39561);
xor U43178 (N_43178,N_36089,N_37836);
nor U43179 (N_43179,N_37786,N_37773);
and U43180 (N_43180,N_37859,N_37315);
nand U43181 (N_43181,N_35632,N_38105);
or U43182 (N_43182,N_35337,N_38056);
nor U43183 (N_43183,N_39073,N_36052);
or U43184 (N_43184,N_38635,N_39963);
nor U43185 (N_43185,N_36803,N_38796);
and U43186 (N_43186,N_38483,N_39263);
nand U43187 (N_43187,N_37116,N_39731);
xnor U43188 (N_43188,N_36769,N_39851);
and U43189 (N_43189,N_39199,N_36870);
or U43190 (N_43190,N_39472,N_37170);
xor U43191 (N_43191,N_38014,N_37769);
nand U43192 (N_43192,N_35990,N_38979);
or U43193 (N_43193,N_38706,N_39370);
or U43194 (N_43194,N_37354,N_35448);
nor U43195 (N_43195,N_35641,N_37924);
and U43196 (N_43196,N_38242,N_37840);
nand U43197 (N_43197,N_35056,N_39900);
xor U43198 (N_43198,N_39761,N_35554);
and U43199 (N_43199,N_38454,N_38056);
xor U43200 (N_43200,N_39649,N_36705);
or U43201 (N_43201,N_37672,N_39153);
nand U43202 (N_43202,N_37328,N_35390);
or U43203 (N_43203,N_38482,N_38945);
nor U43204 (N_43204,N_39523,N_36448);
nand U43205 (N_43205,N_35460,N_36897);
nand U43206 (N_43206,N_39850,N_39337);
and U43207 (N_43207,N_38990,N_37178);
nor U43208 (N_43208,N_37201,N_38847);
xor U43209 (N_43209,N_39646,N_36363);
nor U43210 (N_43210,N_35245,N_37868);
and U43211 (N_43211,N_38895,N_37367);
nand U43212 (N_43212,N_37836,N_38019);
and U43213 (N_43213,N_39753,N_38756);
and U43214 (N_43214,N_39243,N_39953);
nand U43215 (N_43215,N_35826,N_35337);
or U43216 (N_43216,N_35513,N_39616);
and U43217 (N_43217,N_37856,N_39006);
nand U43218 (N_43218,N_39222,N_39409);
or U43219 (N_43219,N_38209,N_38458);
or U43220 (N_43220,N_39465,N_36245);
and U43221 (N_43221,N_38396,N_38995);
xnor U43222 (N_43222,N_35880,N_37598);
nand U43223 (N_43223,N_38793,N_39688);
and U43224 (N_43224,N_36083,N_39812);
and U43225 (N_43225,N_38209,N_35536);
nor U43226 (N_43226,N_35002,N_35596);
and U43227 (N_43227,N_38958,N_35162);
or U43228 (N_43228,N_35365,N_39570);
or U43229 (N_43229,N_39614,N_38414);
or U43230 (N_43230,N_36324,N_37868);
xor U43231 (N_43231,N_38508,N_35505);
nor U43232 (N_43232,N_37977,N_39205);
or U43233 (N_43233,N_35086,N_36711);
xor U43234 (N_43234,N_38906,N_39639);
or U43235 (N_43235,N_39551,N_36668);
xor U43236 (N_43236,N_37863,N_37361);
nand U43237 (N_43237,N_39126,N_36899);
xnor U43238 (N_43238,N_37922,N_36276);
nor U43239 (N_43239,N_36289,N_38148);
and U43240 (N_43240,N_35650,N_39596);
xnor U43241 (N_43241,N_38733,N_37399);
nor U43242 (N_43242,N_38250,N_36270);
or U43243 (N_43243,N_36447,N_37096);
or U43244 (N_43244,N_36302,N_36327);
and U43245 (N_43245,N_38536,N_39094);
nand U43246 (N_43246,N_36048,N_37975);
nand U43247 (N_43247,N_35422,N_38305);
xor U43248 (N_43248,N_38042,N_39268);
nand U43249 (N_43249,N_37805,N_36153);
and U43250 (N_43250,N_37770,N_36061);
nand U43251 (N_43251,N_35240,N_39570);
xor U43252 (N_43252,N_35841,N_39448);
nand U43253 (N_43253,N_36407,N_35331);
xnor U43254 (N_43254,N_37288,N_37618);
nand U43255 (N_43255,N_37604,N_39581);
xor U43256 (N_43256,N_37655,N_39756);
and U43257 (N_43257,N_37026,N_39357);
nor U43258 (N_43258,N_39632,N_38633);
or U43259 (N_43259,N_35360,N_35608);
and U43260 (N_43260,N_36942,N_36355);
nor U43261 (N_43261,N_35207,N_36117);
and U43262 (N_43262,N_39030,N_38766);
nor U43263 (N_43263,N_36831,N_35361);
or U43264 (N_43264,N_35605,N_37868);
nand U43265 (N_43265,N_39429,N_38406);
or U43266 (N_43266,N_35639,N_38699);
nand U43267 (N_43267,N_35067,N_38464);
xor U43268 (N_43268,N_36436,N_38968);
nand U43269 (N_43269,N_37590,N_35052);
nor U43270 (N_43270,N_38732,N_38555);
nand U43271 (N_43271,N_37456,N_38762);
nand U43272 (N_43272,N_36225,N_38747);
nor U43273 (N_43273,N_39101,N_37194);
and U43274 (N_43274,N_37270,N_37768);
nor U43275 (N_43275,N_38880,N_38500);
xor U43276 (N_43276,N_36171,N_35981);
or U43277 (N_43277,N_39287,N_37738);
xor U43278 (N_43278,N_36199,N_39982);
xnor U43279 (N_43279,N_37926,N_37470);
nor U43280 (N_43280,N_35761,N_39761);
nand U43281 (N_43281,N_36882,N_39401);
or U43282 (N_43282,N_39805,N_37968);
and U43283 (N_43283,N_38440,N_35434);
and U43284 (N_43284,N_37004,N_39406);
nor U43285 (N_43285,N_38555,N_37691);
nand U43286 (N_43286,N_36621,N_35720);
nor U43287 (N_43287,N_37546,N_38180);
xor U43288 (N_43288,N_37797,N_35045);
nand U43289 (N_43289,N_35006,N_37536);
and U43290 (N_43290,N_36148,N_35420);
or U43291 (N_43291,N_35120,N_36232);
xnor U43292 (N_43292,N_36055,N_35266);
nand U43293 (N_43293,N_39927,N_37796);
xor U43294 (N_43294,N_35729,N_36919);
or U43295 (N_43295,N_36344,N_38222);
nor U43296 (N_43296,N_36068,N_37470);
nor U43297 (N_43297,N_36725,N_38988);
nor U43298 (N_43298,N_37206,N_39017);
nand U43299 (N_43299,N_36814,N_36415);
xor U43300 (N_43300,N_39617,N_38019);
nand U43301 (N_43301,N_38190,N_39967);
nor U43302 (N_43302,N_38735,N_39749);
nand U43303 (N_43303,N_38260,N_39663);
xor U43304 (N_43304,N_39522,N_39059);
and U43305 (N_43305,N_36662,N_35738);
or U43306 (N_43306,N_39978,N_38335);
or U43307 (N_43307,N_35060,N_38075);
and U43308 (N_43308,N_35783,N_37202);
xnor U43309 (N_43309,N_38145,N_38701);
or U43310 (N_43310,N_38597,N_36470);
nand U43311 (N_43311,N_39950,N_38358);
and U43312 (N_43312,N_36586,N_37651);
or U43313 (N_43313,N_39420,N_39653);
or U43314 (N_43314,N_35297,N_35634);
xnor U43315 (N_43315,N_38143,N_38310);
or U43316 (N_43316,N_39267,N_39717);
xor U43317 (N_43317,N_39276,N_39797);
nand U43318 (N_43318,N_37924,N_35620);
xnor U43319 (N_43319,N_39476,N_35833);
nor U43320 (N_43320,N_36659,N_36811);
nand U43321 (N_43321,N_37857,N_37575);
or U43322 (N_43322,N_37452,N_38595);
xor U43323 (N_43323,N_35621,N_39137);
xor U43324 (N_43324,N_39549,N_35828);
and U43325 (N_43325,N_36347,N_38927);
nand U43326 (N_43326,N_39364,N_36665);
nand U43327 (N_43327,N_39093,N_38666);
nor U43328 (N_43328,N_35599,N_37317);
or U43329 (N_43329,N_37069,N_39619);
or U43330 (N_43330,N_39519,N_39993);
or U43331 (N_43331,N_39189,N_36005);
nor U43332 (N_43332,N_37030,N_38394);
xor U43333 (N_43333,N_35769,N_39448);
nor U43334 (N_43334,N_38980,N_38981);
xor U43335 (N_43335,N_37141,N_38246);
nor U43336 (N_43336,N_38040,N_35898);
or U43337 (N_43337,N_36106,N_37095);
xnor U43338 (N_43338,N_38696,N_39491);
nand U43339 (N_43339,N_37301,N_35398);
nor U43340 (N_43340,N_36346,N_36936);
or U43341 (N_43341,N_37164,N_39339);
nor U43342 (N_43342,N_35088,N_39786);
and U43343 (N_43343,N_35679,N_35132);
or U43344 (N_43344,N_37942,N_36733);
nand U43345 (N_43345,N_36806,N_39269);
nor U43346 (N_43346,N_38131,N_39461);
and U43347 (N_43347,N_36267,N_35361);
nand U43348 (N_43348,N_37450,N_37024);
or U43349 (N_43349,N_36653,N_37635);
nand U43350 (N_43350,N_38899,N_38949);
and U43351 (N_43351,N_36403,N_35878);
xor U43352 (N_43352,N_39109,N_35616);
and U43353 (N_43353,N_36781,N_35883);
or U43354 (N_43354,N_37553,N_39875);
nand U43355 (N_43355,N_35338,N_38187);
or U43356 (N_43356,N_39045,N_37307);
and U43357 (N_43357,N_38420,N_38247);
or U43358 (N_43358,N_36059,N_35144);
nand U43359 (N_43359,N_37583,N_36901);
xnor U43360 (N_43360,N_37043,N_36324);
or U43361 (N_43361,N_35081,N_36861);
nand U43362 (N_43362,N_39501,N_35276);
xor U43363 (N_43363,N_35162,N_36652);
and U43364 (N_43364,N_38649,N_39411);
and U43365 (N_43365,N_38091,N_38024);
and U43366 (N_43366,N_39141,N_37414);
nand U43367 (N_43367,N_36150,N_38143);
xnor U43368 (N_43368,N_38502,N_39652);
and U43369 (N_43369,N_38193,N_35918);
and U43370 (N_43370,N_36083,N_39383);
and U43371 (N_43371,N_36295,N_37030);
and U43372 (N_43372,N_37389,N_35836);
and U43373 (N_43373,N_37219,N_35230);
nor U43374 (N_43374,N_38955,N_37947);
xnor U43375 (N_43375,N_39259,N_36135);
and U43376 (N_43376,N_39235,N_35575);
xor U43377 (N_43377,N_35724,N_35385);
nor U43378 (N_43378,N_36023,N_35281);
nand U43379 (N_43379,N_38792,N_39122);
and U43380 (N_43380,N_38701,N_35090);
and U43381 (N_43381,N_39665,N_37997);
and U43382 (N_43382,N_35473,N_36263);
nor U43383 (N_43383,N_36788,N_37778);
nand U43384 (N_43384,N_38036,N_39132);
xnor U43385 (N_43385,N_37541,N_37602);
or U43386 (N_43386,N_35887,N_35950);
nor U43387 (N_43387,N_37666,N_38281);
or U43388 (N_43388,N_36066,N_35618);
and U43389 (N_43389,N_37898,N_39484);
nor U43390 (N_43390,N_38747,N_35020);
nand U43391 (N_43391,N_39451,N_36006);
xor U43392 (N_43392,N_38490,N_36497);
nand U43393 (N_43393,N_37871,N_35701);
and U43394 (N_43394,N_36110,N_38550);
xnor U43395 (N_43395,N_37210,N_38167);
nor U43396 (N_43396,N_35328,N_37163);
nand U43397 (N_43397,N_37522,N_36804);
nand U43398 (N_43398,N_36164,N_36293);
or U43399 (N_43399,N_35515,N_35192);
nor U43400 (N_43400,N_36134,N_37822);
or U43401 (N_43401,N_35389,N_35894);
nand U43402 (N_43402,N_35517,N_39427);
or U43403 (N_43403,N_38040,N_35448);
xnor U43404 (N_43404,N_36806,N_36245);
or U43405 (N_43405,N_35530,N_36175);
nand U43406 (N_43406,N_36500,N_35474);
xnor U43407 (N_43407,N_35004,N_36263);
and U43408 (N_43408,N_39576,N_35069);
nand U43409 (N_43409,N_39983,N_35196);
and U43410 (N_43410,N_35418,N_35860);
and U43411 (N_43411,N_37896,N_36910);
and U43412 (N_43412,N_36722,N_36313);
or U43413 (N_43413,N_36548,N_39970);
and U43414 (N_43414,N_39273,N_38874);
xnor U43415 (N_43415,N_35309,N_39924);
nor U43416 (N_43416,N_35552,N_37142);
or U43417 (N_43417,N_39192,N_36145);
or U43418 (N_43418,N_35428,N_35761);
nand U43419 (N_43419,N_39502,N_39636);
nor U43420 (N_43420,N_36420,N_35943);
nor U43421 (N_43421,N_35953,N_36830);
xnor U43422 (N_43422,N_36449,N_38275);
nand U43423 (N_43423,N_35801,N_38303);
and U43424 (N_43424,N_36388,N_37087);
nor U43425 (N_43425,N_35042,N_37612);
and U43426 (N_43426,N_36650,N_38560);
xor U43427 (N_43427,N_39163,N_39756);
and U43428 (N_43428,N_36386,N_36754);
xor U43429 (N_43429,N_37619,N_36897);
xnor U43430 (N_43430,N_37021,N_37053);
and U43431 (N_43431,N_37286,N_35229);
nand U43432 (N_43432,N_37044,N_38361);
xnor U43433 (N_43433,N_38699,N_39581);
and U43434 (N_43434,N_39834,N_36252);
xor U43435 (N_43435,N_35784,N_36291);
nand U43436 (N_43436,N_39576,N_37951);
and U43437 (N_43437,N_39014,N_36926);
nor U43438 (N_43438,N_36068,N_35630);
xnor U43439 (N_43439,N_36916,N_39856);
and U43440 (N_43440,N_37464,N_35459);
nand U43441 (N_43441,N_39514,N_37639);
nand U43442 (N_43442,N_38427,N_36279);
and U43443 (N_43443,N_38150,N_37914);
xor U43444 (N_43444,N_38584,N_39812);
and U43445 (N_43445,N_39543,N_35416);
nand U43446 (N_43446,N_39639,N_38096);
or U43447 (N_43447,N_37892,N_35803);
xor U43448 (N_43448,N_37230,N_37396);
nand U43449 (N_43449,N_38224,N_39370);
or U43450 (N_43450,N_37078,N_35383);
nand U43451 (N_43451,N_36019,N_39065);
or U43452 (N_43452,N_38602,N_37443);
and U43453 (N_43453,N_39245,N_35683);
nor U43454 (N_43454,N_35726,N_36892);
and U43455 (N_43455,N_38183,N_39829);
xnor U43456 (N_43456,N_38529,N_38050);
or U43457 (N_43457,N_36865,N_36063);
xor U43458 (N_43458,N_39112,N_38703);
nor U43459 (N_43459,N_37258,N_38007);
or U43460 (N_43460,N_35452,N_38481);
and U43461 (N_43461,N_39451,N_39254);
xor U43462 (N_43462,N_38004,N_37987);
nor U43463 (N_43463,N_35400,N_37301);
xor U43464 (N_43464,N_36779,N_39231);
nand U43465 (N_43465,N_36694,N_39949);
nand U43466 (N_43466,N_36573,N_37931);
or U43467 (N_43467,N_38170,N_35971);
and U43468 (N_43468,N_37656,N_36937);
or U43469 (N_43469,N_39945,N_39491);
nor U43470 (N_43470,N_35819,N_37135);
nand U43471 (N_43471,N_38116,N_36235);
nand U43472 (N_43472,N_38997,N_36836);
or U43473 (N_43473,N_37612,N_38509);
nand U43474 (N_43474,N_37000,N_38519);
xnor U43475 (N_43475,N_36716,N_37048);
nand U43476 (N_43476,N_36601,N_39008);
xnor U43477 (N_43477,N_38846,N_37811);
nor U43478 (N_43478,N_37754,N_35940);
xnor U43479 (N_43479,N_38369,N_39030);
xor U43480 (N_43480,N_36105,N_35393);
xnor U43481 (N_43481,N_39191,N_37494);
and U43482 (N_43482,N_37912,N_36838);
nor U43483 (N_43483,N_36056,N_38008);
xor U43484 (N_43484,N_38403,N_39412);
or U43485 (N_43485,N_35361,N_39268);
or U43486 (N_43486,N_35307,N_35513);
nor U43487 (N_43487,N_37224,N_39580);
nor U43488 (N_43488,N_36312,N_39523);
and U43489 (N_43489,N_39284,N_39365);
xnor U43490 (N_43490,N_38589,N_37363);
xnor U43491 (N_43491,N_39754,N_35142);
xor U43492 (N_43492,N_36617,N_39061);
or U43493 (N_43493,N_38381,N_36501);
xor U43494 (N_43494,N_36619,N_36447);
xnor U43495 (N_43495,N_37995,N_39367);
xnor U43496 (N_43496,N_39547,N_37921);
and U43497 (N_43497,N_36825,N_38770);
nor U43498 (N_43498,N_35606,N_35690);
xnor U43499 (N_43499,N_38321,N_35693);
xor U43500 (N_43500,N_35181,N_37121);
nor U43501 (N_43501,N_37747,N_35401);
xor U43502 (N_43502,N_35706,N_35998);
xnor U43503 (N_43503,N_39605,N_35916);
nor U43504 (N_43504,N_38019,N_38127);
nand U43505 (N_43505,N_36412,N_37004);
nand U43506 (N_43506,N_37533,N_39796);
xnor U43507 (N_43507,N_38816,N_36421);
xnor U43508 (N_43508,N_39872,N_36819);
nor U43509 (N_43509,N_36826,N_36305);
nand U43510 (N_43510,N_38406,N_37503);
and U43511 (N_43511,N_35756,N_36526);
and U43512 (N_43512,N_36945,N_37213);
and U43513 (N_43513,N_36892,N_39823);
nand U43514 (N_43514,N_36643,N_36084);
or U43515 (N_43515,N_37181,N_35520);
nor U43516 (N_43516,N_39734,N_38071);
and U43517 (N_43517,N_37539,N_38997);
nor U43518 (N_43518,N_37633,N_35445);
nand U43519 (N_43519,N_39320,N_35643);
xor U43520 (N_43520,N_35657,N_38676);
nor U43521 (N_43521,N_36045,N_37848);
nor U43522 (N_43522,N_38402,N_37703);
nand U43523 (N_43523,N_35355,N_37903);
nand U43524 (N_43524,N_39504,N_37529);
nor U43525 (N_43525,N_37996,N_37229);
or U43526 (N_43526,N_36129,N_38265);
or U43527 (N_43527,N_36891,N_38015);
nor U43528 (N_43528,N_37467,N_35868);
xor U43529 (N_43529,N_35968,N_38578);
and U43530 (N_43530,N_36444,N_35119);
or U43531 (N_43531,N_37145,N_35648);
nor U43532 (N_43532,N_38866,N_38493);
nand U43533 (N_43533,N_38492,N_38160);
and U43534 (N_43534,N_37270,N_38406);
xor U43535 (N_43535,N_35458,N_39272);
nor U43536 (N_43536,N_37159,N_38270);
xor U43537 (N_43537,N_37570,N_36833);
and U43538 (N_43538,N_35521,N_37847);
or U43539 (N_43539,N_36478,N_39425);
and U43540 (N_43540,N_39970,N_39123);
or U43541 (N_43541,N_35847,N_38771);
nand U43542 (N_43542,N_39679,N_38149);
and U43543 (N_43543,N_37007,N_35082);
or U43544 (N_43544,N_35215,N_36843);
and U43545 (N_43545,N_36569,N_35756);
nand U43546 (N_43546,N_36778,N_35351);
nor U43547 (N_43547,N_35146,N_36965);
xor U43548 (N_43548,N_37962,N_35286);
or U43549 (N_43549,N_37179,N_36654);
xnor U43550 (N_43550,N_35562,N_35786);
nor U43551 (N_43551,N_37316,N_38772);
xor U43552 (N_43552,N_37919,N_36232);
xor U43553 (N_43553,N_39325,N_38538);
nor U43554 (N_43554,N_36338,N_35570);
and U43555 (N_43555,N_35960,N_37433);
and U43556 (N_43556,N_39611,N_36944);
and U43557 (N_43557,N_38246,N_38906);
or U43558 (N_43558,N_36944,N_39436);
or U43559 (N_43559,N_37380,N_36165);
nand U43560 (N_43560,N_39823,N_36548);
nor U43561 (N_43561,N_37554,N_35506);
or U43562 (N_43562,N_35029,N_39227);
xor U43563 (N_43563,N_38707,N_38046);
and U43564 (N_43564,N_39728,N_36283);
nand U43565 (N_43565,N_38290,N_35249);
and U43566 (N_43566,N_37961,N_36142);
nand U43567 (N_43567,N_38629,N_37039);
nor U43568 (N_43568,N_39326,N_39043);
and U43569 (N_43569,N_38799,N_36646);
or U43570 (N_43570,N_35679,N_36027);
nand U43571 (N_43571,N_37310,N_39715);
nand U43572 (N_43572,N_35473,N_36079);
nor U43573 (N_43573,N_38640,N_35032);
and U43574 (N_43574,N_35131,N_39301);
and U43575 (N_43575,N_35765,N_35425);
and U43576 (N_43576,N_36803,N_37114);
nor U43577 (N_43577,N_36774,N_37498);
or U43578 (N_43578,N_36714,N_35411);
nand U43579 (N_43579,N_39771,N_36705);
nor U43580 (N_43580,N_36870,N_38485);
and U43581 (N_43581,N_35307,N_36557);
nor U43582 (N_43582,N_35763,N_39331);
or U43583 (N_43583,N_35618,N_38463);
nor U43584 (N_43584,N_39379,N_39606);
or U43585 (N_43585,N_35439,N_38247);
nor U43586 (N_43586,N_35935,N_35304);
and U43587 (N_43587,N_35235,N_38674);
or U43588 (N_43588,N_39695,N_36600);
nor U43589 (N_43589,N_35910,N_37902);
or U43590 (N_43590,N_35778,N_36320);
nor U43591 (N_43591,N_36851,N_36481);
or U43592 (N_43592,N_38308,N_35578);
or U43593 (N_43593,N_38728,N_37455);
and U43594 (N_43594,N_35162,N_38218);
nand U43595 (N_43595,N_37620,N_38717);
nor U43596 (N_43596,N_39652,N_37923);
nor U43597 (N_43597,N_36307,N_35552);
or U43598 (N_43598,N_38625,N_39366);
xor U43599 (N_43599,N_36760,N_39758);
nor U43600 (N_43600,N_35227,N_39212);
and U43601 (N_43601,N_39779,N_37910);
or U43602 (N_43602,N_38289,N_36080);
nor U43603 (N_43603,N_38419,N_38083);
nand U43604 (N_43604,N_37666,N_36136);
nor U43605 (N_43605,N_39216,N_39791);
nor U43606 (N_43606,N_39798,N_39091);
nor U43607 (N_43607,N_38424,N_35712);
nor U43608 (N_43608,N_38965,N_36150);
or U43609 (N_43609,N_35949,N_36866);
and U43610 (N_43610,N_38641,N_39538);
and U43611 (N_43611,N_38603,N_37232);
and U43612 (N_43612,N_38217,N_35518);
xnor U43613 (N_43613,N_39941,N_39839);
nor U43614 (N_43614,N_35047,N_37484);
nor U43615 (N_43615,N_36140,N_37763);
nor U43616 (N_43616,N_39153,N_39258);
and U43617 (N_43617,N_36226,N_35765);
nand U43618 (N_43618,N_37269,N_39860);
or U43619 (N_43619,N_36914,N_36842);
xor U43620 (N_43620,N_38741,N_36812);
xor U43621 (N_43621,N_35888,N_37005);
and U43622 (N_43622,N_35981,N_39680);
or U43623 (N_43623,N_38552,N_37922);
or U43624 (N_43624,N_39205,N_38565);
and U43625 (N_43625,N_38464,N_38982);
nor U43626 (N_43626,N_37607,N_39968);
and U43627 (N_43627,N_39960,N_37092);
nand U43628 (N_43628,N_37543,N_35298);
and U43629 (N_43629,N_39686,N_36389);
nor U43630 (N_43630,N_35864,N_35473);
nand U43631 (N_43631,N_35642,N_35121);
or U43632 (N_43632,N_37963,N_39502);
or U43633 (N_43633,N_37081,N_37759);
or U43634 (N_43634,N_35450,N_35066);
nand U43635 (N_43635,N_36960,N_39997);
or U43636 (N_43636,N_36379,N_36203);
xor U43637 (N_43637,N_37610,N_35358);
nand U43638 (N_43638,N_39188,N_36774);
nor U43639 (N_43639,N_38965,N_38392);
xnor U43640 (N_43640,N_36472,N_36875);
xnor U43641 (N_43641,N_39555,N_38323);
nand U43642 (N_43642,N_36925,N_39932);
and U43643 (N_43643,N_38742,N_39764);
nor U43644 (N_43644,N_36462,N_38517);
nor U43645 (N_43645,N_35709,N_36349);
xnor U43646 (N_43646,N_35702,N_39847);
nor U43647 (N_43647,N_37309,N_35040);
nor U43648 (N_43648,N_37296,N_37341);
or U43649 (N_43649,N_35243,N_37294);
nor U43650 (N_43650,N_38044,N_38692);
xnor U43651 (N_43651,N_39716,N_35162);
nand U43652 (N_43652,N_35131,N_39467);
nand U43653 (N_43653,N_35432,N_36165);
and U43654 (N_43654,N_37595,N_36955);
and U43655 (N_43655,N_38538,N_35541);
nor U43656 (N_43656,N_38936,N_35354);
or U43657 (N_43657,N_39964,N_35337);
and U43658 (N_43658,N_38744,N_39927);
and U43659 (N_43659,N_38269,N_35174);
or U43660 (N_43660,N_37511,N_37689);
xor U43661 (N_43661,N_37795,N_36322);
or U43662 (N_43662,N_39748,N_38123);
xnor U43663 (N_43663,N_35129,N_38435);
or U43664 (N_43664,N_39930,N_35893);
or U43665 (N_43665,N_35981,N_37833);
xnor U43666 (N_43666,N_37430,N_37660);
and U43667 (N_43667,N_36142,N_36842);
and U43668 (N_43668,N_36446,N_39512);
and U43669 (N_43669,N_36666,N_36523);
and U43670 (N_43670,N_37395,N_39489);
nor U43671 (N_43671,N_37861,N_35946);
nand U43672 (N_43672,N_39332,N_39139);
xor U43673 (N_43673,N_37234,N_36643);
or U43674 (N_43674,N_39306,N_36473);
or U43675 (N_43675,N_35453,N_38180);
or U43676 (N_43676,N_36210,N_37087);
xnor U43677 (N_43677,N_36139,N_37090);
xnor U43678 (N_43678,N_35179,N_36322);
nand U43679 (N_43679,N_36369,N_38684);
nor U43680 (N_43680,N_36079,N_39724);
and U43681 (N_43681,N_36889,N_35755);
nand U43682 (N_43682,N_35673,N_37471);
and U43683 (N_43683,N_39409,N_37482);
or U43684 (N_43684,N_38041,N_37029);
nor U43685 (N_43685,N_35676,N_35123);
and U43686 (N_43686,N_37396,N_38921);
and U43687 (N_43687,N_39099,N_37325);
xor U43688 (N_43688,N_37022,N_38416);
nand U43689 (N_43689,N_38384,N_37800);
or U43690 (N_43690,N_39258,N_39550);
nand U43691 (N_43691,N_35516,N_37745);
and U43692 (N_43692,N_39209,N_37039);
nor U43693 (N_43693,N_36644,N_39346);
xor U43694 (N_43694,N_37689,N_35159);
and U43695 (N_43695,N_38250,N_39144);
and U43696 (N_43696,N_38636,N_37437);
nor U43697 (N_43697,N_35419,N_36025);
and U43698 (N_43698,N_38330,N_39499);
nand U43699 (N_43699,N_35189,N_35284);
or U43700 (N_43700,N_37083,N_39649);
nor U43701 (N_43701,N_39217,N_36278);
xor U43702 (N_43702,N_39189,N_36134);
nand U43703 (N_43703,N_39459,N_38513);
nand U43704 (N_43704,N_37819,N_39566);
xor U43705 (N_43705,N_37553,N_39197);
nand U43706 (N_43706,N_38158,N_36384);
and U43707 (N_43707,N_38398,N_39945);
nand U43708 (N_43708,N_39116,N_38200);
xnor U43709 (N_43709,N_39850,N_38261);
nor U43710 (N_43710,N_39828,N_35469);
or U43711 (N_43711,N_38117,N_38467);
xor U43712 (N_43712,N_36910,N_35240);
or U43713 (N_43713,N_36763,N_35232);
or U43714 (N_43714,N_35046,N_36516);
nor U43715 (N_43715,N_36772,N_38366);
and U43716 (N_43716,N_37341,N_38365);
nand U43717 (N_43717,N_35227,N_35151);
nor U43718 (N_43718,N_39248,N_35778);
nor U43719 (N_43719,N_39501,N_36717);
or U43720 (N_43720,N_39878,N_39275);
and U43721 (N_43721,N_39460,N_38978);
nor U43722 (N_43722,N_37680,N_35271);
nand U43723 (N_43723,N_35519,N_39365);
and U43724 (N_43724,N_39506,N_35512);
xnor U43725 (N_43725,N_35695,N_35658);
nand U43726 (N_43726,N_38284,N_39545);
or U43727 (N_43727,N_39186,N_38771);
nand U43728 (N_43728,N_39980,N_36682);
nor U43729 (N_43729,N_35625,N_36477);
xnor U43730 (N_43730,N_35640,N_37162);
or U43731 (N_43731,N_35018,N_39288);
and U43732 (N_43732,N_35662,N_37569);
nand U43733 (N_43733,N_38877,N_39317);
and U43734 (N_43734,N_36606,N_36504);
nor U43735 (N_43735,N_37185,N_38589);
nand U43736 (N_43736,N_38325,N_39968);
or U43737 (N_43737,N_35511,N_37806);
or U43738 (N_43738,N_38817,N_36050);
nand U43739 (N_43739,N_36079,N_38043);
nor U43740 (N_43740,N_39486,N_35248);
or U43741 (N_43741,N_37271,N_38984);
nand U43742 (N_43742,N_36373,N_39424);
nand U43743 (N_43743,N_39232,N_35634);
nor U43744 (N_43744,N_38245,N_38862);
and U43745 (N_43745,N_37150,N_38102);
nand U43746 (N_43746,N_36235,N_36776);
and U43747 (N_43747,N_35957,N_35930);
xnor U43748 (N_43748,N_37497,N_36518);
nand U43749 (N_43749,N_38974,N_38349);
nor U43750 (N_43750,N_36554,N_38850);
nand U43751 (N_43751,N_36403,N_39986);
and U43752 (N_43752,N_35078,N_37897);
xnor U43753 (N_43753,N_39056,N_39853);
nand U43754 (N_43754,N_37459,N_38762);
xor U43755 (N_43755,N_35272,N_35720);
and U43756 (N_43756,N_38195,N_39865);
nor U43757 (N_43757,N_37988,N_36677);
nand U43758 (N_43758,N_37055,N_36892);
and U43759 (N_43759,N_37795,N_35864);
xor U43760 (N_43760,N_36354,N_38210);
and U43761 (N_43761,N_39839,N_35939);
nor U43762 (N_43762,N_39366,N_36186);
or U43763 (N_43763,N_35131,N_38711);
and U43764 (N_43764,N_35527,N_36098);
xor U43765 (N_43765,N_37285,N_39870);
nor U43766 (N_43766,N_35190,N_35499);
nor U43767 (N_43767,N_37654,N_39934);
and U43768 (N_43768,N_39510,N_37481);
or U43769 (N_43769,N_39140,N_38044);
nor U43770 (N_43770,N_35754,N_39062);
nor U43771 (N_43771,N_39857,N_38532);
nand U43772 (N_43772,N_38980,N_35865);
and U43773 (N_43773,N_39184,N_38334);
nor U43774 (N_43774,N_37605,N_39074);
nor U43775 (N_43775,N_36626,N_36330);
nand U43776 (N_43776,N_35289,N_35670);
xnor U43777 (N_43777,N_39358,N_35996);
xor U43778 (N_43778,N_36907,N_36436);
xnor U43779 (N_43779,N_36344,N_39134);
nand U43780 (N_43780,N_39711,N_37086);
nor U43781 (N_43781,N_37199,N_36441);
nand U43782 (N_43782,N_35738,N_35736);
nand U43783 (N_43783,N_38188,N_39756);
and U43784 (N_43784,N_39251,N_37691);
nand U43785 (N_43785,N_36515,N_35199);
nand U43786 (N_43786,N_37018,N_37626);
nand U43787 (N_43787,N_39545,N_38086);
nand U43788 (N_43788,N_36157,N_37122);
nand U43789 (N_43789,N_37693,N_35229);
nand U43790 (N_43790,N_38977,N_35695);
nor U43791 (N_43791,N_36066,N_38636);
xnor U43792 (N_43792,N_35364,N_35338);
nand U43793 (N_43793,N_38148,N_35258);
and U43794 (N_43794,N_39960,N_39240);
or U43795 (N_43795,N_35872,N_37277);
nor U43796 (N_43796,N_38332,N_35962);
xor U43797 (N_43797,N_37689,N_35549);
and U43798 (N_43798,N_39423,N_36188);
and U43799 (N_43799,N_37586,N_38504);
and U43800 (N_43800,N_36564,N_36254);
or U43801 (N_43801,N_39899,N_37572);
or U43802 (N_43802,N_35992,N_38163);
and U43803 (N_43803,N_37069,N_35999);
or U43804 (N_43804,N_39388,N_37628);
xnor U43805 (N_43805,N_38946,N_39746);
nor U43806 (N_43806,N_35468,N_35727);
and U43807 (N_43807,N_39573,N_37992);
xnor U43808 (N_43808,N_38495,N_37845);
nand U43809 (N_43809,N_36457,N_39087);
and U43810 (N_43810,N_38265,N_37801);
or U43811 (N_43811,N_39457,N_39919);
and U43812 (N_43812,N_38891,N_38474);
nor U43813 (N_43813,N_38875,N_39661);
nand U43814 (N_43814,N_39674,N_36721);
or U43815 (N_43815,N_36279,N_39615);
and U43816 (N_43816,N_38870,N_38733);
xnor U43817 (N_43817,N_39128,N_39106);
or U43818 (N_43818,N_37315,N_38560);
xnor U43819 (N_43819,N_38493,N_38328);
or U43820 (N_43820,N_35294,N_35005);
nand U43821 (N_43821,N_38576,N_35382);
xor U43822 (N_43822,N_35712,N_37173);
xor U43823 (N_43823,N_37687,N_37652);
and U43824 (N_43824,N_35269,N_38973);
or U43825 (N_43825,N_38449,N_38796);
nor U43826 (N_43826,N_36758,N_39116);
or U43827 (N_43827,N_35987,N_38253);
nor U43828 (N_43828,N_35886,N_38391);
and U43829 (N_43829,N_38777,N_38986);
xor U43830 (N_43830,N_35399,N_38487);
and U43831 (N_43831,N_35867,N_37293);
and U43832 (N_43832,N_35651,N_37106);
nand U43833 (N_43833,N_36188,N_39820);
or U43834 (N_43834,N_35746,N_38023);
nand U43835 (N_43835,N_36180,N_37527);
nor U43836 (N_43836,N_37645,N_38081);
or U43837 (N_43837,N_39968,N_36087);
xor U43838 (N_43838,N_38576,N_35325);
or U43839 (N_43839,N_36515,N_38971);
and U43840 (N_43840,N_38392,N_39233);
xor U43841 (N_43841,N_36773,N_37296);
nand U43842 (N_43842,N_39772,N_35752);
and U43843 (N_43843,N_35982,N_36104);
nand U43844 (N_43844,N_38768,N_38436);
xnor U43845 (N_43845,N_36149,N_38279);
nand U43846 (N_43846,N_39672,N_35629);
or U43847 (N_43847,N_35752,N_35379);
xor U43848 (N_43848,N_39272,N_38439);
and U43849 (N_43849,N_39941,N_39730);
or U43850 (N_43850,N_36508,N_39695);
nor U43851 (N_43851,N_39419,N_36236);
nand U43852 (N_43852,N_38503,N_37595);
nand U43853 (N_43853,N_37781,N_36975);
and U43854 (N_43854,N_39296,N_36609);
and U43855 (N_43855,N_38449,N_36030);
and U43856 (N_43856,N_37023,N_36818);
nor U43857 (N_43857,N_38123,N_36237);
nor U43858 (N_43858,N_36822,N_39613);
and U43859 (N_43859,N_37787,N_36857);
or U43860 (N_43860,N_36599,N_37418);
and U43861 (N_43861,N_38073,N_39036);
nand U43862 (N_43862,N_35394,N_39068);
nand U43863 (N_43863,N_37692,N_37214);
xor U43864 (N_43864,N_35794,N_38032);
nor U43865 (N_43865,N_37418,N_35510);
nand U43866 (N_43866,N_35804,N_37550);
xnor U43867 (N_43867,N_37200,N_37334);
or U43868 (N_43868,N_39608,N_36022);
xnor U43869 (N_43869,N_39819,N_36714);
or U43870 (N_43870,N_38542,N_35459);
or U43871 (N_43871,N_36830,N_38252);
nor U43872 (N_43872,N_38248,N_36844);
nand U43873 (N_43873,N_35772,N_35513);
nor U43874 (N_43874,N_35252,N_38403);
nor U43875 (N_43875,N_37199,N_35430);
nor U43876 (N_43876,N_39739,N_36460);
nor U43877 (N_43877,N_35915,N_37630);
nand U43878 (N_43878,N_38295,N_39316);
xnor U43879 (N_43879,N_37338,N_38680);
and U43880 (N_43880,N_39405,N_39792);
and U43881 (N_43881,N_35783,N_36601);
or U43882 (N_43882,N_36628,N_35697);
or U43883 (N_43883,N_37611,N_39261);
nor U43884 (N_43884,N_37202,N_38661);
nand U43885 (N_43885,N_39072,N_35642);
and U43886 (N_43886,N_36721,N_38062);
nand U43887 (N_43887,N_35344,N_36900);
nor U43888 (N_43888,N_36196,N_35695);
xor U43889 (N_43889,N_38959,N_35455);
and U43890 (N_43890,N_39479,N_38277);
and U43891 (N_43891,N_37727,N_39039);
nor U43892 (N_43892,N_35739,N_35640);
and U43893 (N_43893,N_36152,N_36627);
nand U43894 (N_43894,N_35052,N_35936);
and U43895 (N_43895,N_35769,N_37064);
or U43896 (N_43896,N_39294,N_39402);
or U43897 (N_43897,N_35723,N_35573);
xor U43898 (N_43898,N_36114,N_35697);
nor U43899 (N_43899,N_36410,N_39561);
and U43900 (N_43900,N_39361,N_36228);
nand U43901 (N_43901,N_36940,N_37516);
and U43902 (N_43902,N_35878,N_37162);
xor U43903 (N_43903,N_39556,N_36385);
and U43904 (N_43904,N_39262,N_36013);
or U43905 (N_43905,N_39386,N_37625);
and U43906 (N_43906,N_37832,N_39385);
nand U43907 (N_43907,N_38231,N_36459);
xor U43908 (N_43908,N_35626,N_37077);
xor U43909 (N_43909,N_36717,N_38338);
or U43910 (N_43910,N_35949,N_36965);
xor U43911 (N_43911,N_35048,N_35841);
or U43912 (N_43912,N_39390,N_38792);
and U43913 (N_43913,N_36391,N_37288);
xnor U43914 (N_43914,N_37236,N_36665);
nor U43915 (N_43915,N_35691,N_38718);
nand U43916 (N_43916,N_35526,N_38985);
or U43917 (N_43917,N_35595,N_37893);
and U43918 (N_43918,N_35512,N_37703);
or U43919 (N_43919,N_38810,N_39780);
xnor U43920 (N_43920,N_39667,N_38944);
nor U43921 (N_43921,N_39905,N_36837);
and U43922 (N_43922,N_38247,N_37915);
xnor U43923 (N_43923,N_35696,N_35984);
xor U43924 (N_43924,N_38603,N_35997);
or U43925 (N_43925,N_37136,N_38687);
xor U43926 (N_43926,N_35307,N_35793);
nor U43927 (N_43927,N_38280,N_38748);
nand U43928 (N_43928,N_36021,N_35956);
and U43929 (N_43929,N_35011,N_39110);
or U43930 (N_43930,N_39792,N_37032);
nor U43931 (N_43931,N_38745,N_35468);
xnor U43932 (N_43932,N_35375,N_38460);
or U43933 (N_43933,N_38858,N_39597);
nand U43934 (N_43934,N_39158,N_37923);
xnor U43935 (N_43935,N_37024,N_38836);
xor U43936 (N_43936,N_38216,N_35153);
nand U43937 (N_43937,N_37346,N_39744);
nor U43938 (N_43938,N_37144,N_37661);
and U43939 (N_43939,N_39306,N_38453);
or U43940 (N_43940,N_36255,N_37159);
and U43941 (N_43941,N_38523,N_38090);
or U43942 (N_43942,N_36821,N_37650);
and U43943 (N_43943,N_39386,N_39479);
nor U43944 (N_43944,N_38452,N_39691);
or U43945 (N_43945,N_37499,N_39589);
nand U43946 (N_43946,N_36052,N_36139);
and U43947 (N_43947,N_37575,N_36986);
and U43948 (N_43948,N_38260,N_38213);
nor U43949 (N_43949,N_39117,N_37367);
xnor U43950 (N_43950,N_35405,N_35612);
xnor U43951 (N_43951,N_36235,N_36072);
xnor U43952 (N_43952,N_35869,N_35626);
and U43953 (N_43953,N_37858,N_38675);
and U43954 (N_43954,N_36656,N_36363);
and U43955 (N_43955,N_37004,N_36638);
or U43956 (N_43956,N_35926,N_37122);
nand U43957 (N_43957,N_36157,N_38756);
nand U43958 (N_43958,N_37074,N_39434);
xnor U43959 (N_43959,N_39193,N_36636);
or U43960 (N_43960,N_35277,N_35972);
xor U43961 (N_43961,N_37652,N_39692);
nor U43962 (N_43962,N_37243,N_39598);
nand U43963 (N_43963,N_38624,N_39614);
nand U43964 (N_43964,N_39568,N_37152);
nor U43965 (N_43965,N_37791,N_39228);
and U43966 (N_43966,N_37997,N_37144);
or U43967 (N_43967,N_37052,N_35033);
and U43968 (N_43968,N_35487,N_37625);
xor U43969 (N_43969,N_37090,N_38169);
xor U43970 (N_43970,N_39085,N_37075);
or U43971 (N_43971,N_36323,N_35073);
and U43972 (N_43972,N_35262,N_35433);
xnor U43973 (N_43973,N_39548,N_37510);
nor U43974 (N_43974,N_37752,N_38145);
xor U43975 (N_43975,N_38139,N_35073);
or U43976 (N_43976,N_39860,N_37117);
nor U43977 (N_43977,N_39529,N_36289);
and U43978 (N_43978,N_39565,N_39631);
xnor U43979 (N_43979,N_38678,N_37144);
and U43980 (N_43980,N_37296,N_39627);
xor U43981 (N_43981,N_38197,N_35676);
nand U43982 (N_43982,N_36737,N_36285);
nor U43983 (N_43983,N_39188,N_35799);
and U43984 (N_43984,N_36144,N_38702);
and U43985 (N_43985,N_37118,N_38443);
and U43986 (N_43986,N_39216,N_35302);
xnor U43987 (N_43987,N_39017,N_35075);
nor U43988 (N_43988,N_39717,N_35021);
or U43989 (N_43989,N_35051,N_35252);
and U43990 (N_43990,N_35533,N_38949);
nor U43991 (N_43991,N_35057,N_35592);
xor U43992 (N_43992,N_36175,N_36077);
xor U43993 (N_43993,N_35162,N_37932);
nand U43994 (N_43994,N_37057,N_39408);
and U43995 (N_43995,N_39173,N_37118);
nor U43996 (N_43996,N_36678,N_36466);
or U43997 (N_43997,N_35944,N_38731);
nor U43998 (N_43998,N_35824,N_35244);
nand U43999 (N_43999,N_35549,N_39960);
nand U44000 (N_44000,N_36627,N_37637);
nor U44001 (N_44001,N_36834,N_36001);
and U44002 (N_44002,N_36938,N_38159);
or U44003 (N_44003,N_39718,N_37524);
or U44004 (N_44004,N_39458,N_37149);
or U44005 (N_44005,N_38489,N_35004);
xnor U44006 (N_44006,N_35588,N_39117);
or U44007 (N_44007,N_35692,N_38821);
nor U44008 (N_44008,N_39648,N_39548);
xnor U44009 (N_44009,N_36256,N_36647);
nor U44010 (N_44010,N_37425,N_37680);
nor U44011 (N_44011,N_37042,N_38261);
or U44012 (N_44012,N_39857,N_36735);
nand U44013 (N_44013,N_35430,N_39045);
xnor U44014 (N_44014,N_35575,N_38354);
nand U44015 (N_44015,N_36722,N_37786);
or U44016 (N_44016,N_35758,N_37960);
nor U44017 (N_44017,N_36897,N_36652);
or U44018 (N_44018,N_35687,N_38818);
and U44019 (N_44019,N_37107,N_39729);
and U44020 (N_44020,N_35537,N_37499);
and U44021 (N_44021,N_39167,N_39320);
or U44022 (N_44022,N_37408,N_39176);
or U44023 (N_44023,N_39684,N_39045);
and U44024 (N_44024,N_36171,N_35736);
or U44025 (N_44025,N_39345,N_39003);
nand U44026 (N_44026,N_36175,N_37406);
nor U44027 (N_44027,N_36123,N_39129);
xor U44028 (N_44028,N_36078,N_38774);
or U44029 (N_44029,N_37713,N_39593);
xor U44030 (N_44030,N_37670,N_37926);
or U44031 (N_44031,N_36077,N_37998);
or U44032 (N_44032,N_39536,N_38974);
xor U44033 (N_44033,N_35100,N_39793);
or U44034 (N_44034,N_37130,N_38586);
and U44035 (N_44035,N_37145,N_37594);
or U44036 (N_44036,N_37129,N_35714);
nor U44037 (N_44037,N_35343,N_38536);
nor U44038 (N_44038,N_36469,N_39901);
xor U44039 (N_44039,N_35293,N_36774);
nand U44040 (N_44040,N_35947,N_37955);
xor U44041 (N_44041,N_36197,N_36493);
and U44042 (N_44042,N_39308,N_37592);
nor U44043 (N_44043,N_35410,N_38106);
nor U44044 (N_44044,N_39900,N_37774);
and U44045 (N_44045,N_39181,N_37829);
xnor U44046 (N_44046,N_37746,N_36591);
nand U44047 (N_44047,N_37153,N_36231);
xnor U44048 (N_44048,N_35380,N_36306);
or U44049 (N_44049,N_36215,N_36787);
and U44050 (N_44050,N_38117,N_38833);
and U44051 (N_44051,N_35687,N_37829);
or U44052 (N_44052,N_36014,N_39370);
xnor U44053 (N_44053,N_38122,N_35367);
nand U44054 (N_44054,N_36525,N_36307);
nor U44055 (N_44055,N_39944,N_39410);
xnor U44056 (N_44056,N_37915,N_38280);
nand U44057 (N_44057,N_39408,N_39071);
nor U44058 (N_44058,N_38510,N_38446);
and U44059 (N_44059,N_36849,N_39255);
nand U44060 (N_44060,N_35551,N_36389);
nand U44061 (N_44061,N_36042,N_37666);
xor U44062 (N_44062,N_37050,N_37522);
nor U44063 (N_44063,N_36093,N_35494);
xnor U44064 (N_44064,N_38617,N_38588);
and U44065 (N_44065,N_37381,N_36357);
xnor U44066 (N_44066,N_37235,N_38074);
and U44067 (N_44067,N_36327,N_39322);
xnor U44068 (N_44068,N_37334,N_38557);
nand U44069 (N_44069,N_38697,N_38822);
nor U44070 (N_44070,N_39850,N_35609);
xor U44071 (N_44071,N_37519,N_38937);
xnor U44072 (N_44072,N_39357,N_39129);
or U44073 (N_44073,N_36172,N_38964);
and U44074 (N_44074,N_36567,N_37885);
and U44075 (N_44075,N_38918,N_39007);
nand U44076 (N_44076,N_37354,N_37441);
nand U44077 (N_44077,N_36610,N_35751);
and U44078 (N_44078,N_39807,N_38164);
or U44079 (N_44079,N_36501,N_38340);
nand U44080 (N_44080,N_39715,N_36272);
nor U44081 (N_44081,N_38480,N_36940);
xnor U44082 (N_44082,N_35927,N_37743);
nand U44083 (N_44083,N_38814,N_35706);
nor U44084 (N_44084,N_38620,N_37455);
or U44085 (N_44085,N_36210,N_39657);
and U44086 (N_44086,N_39747,N_39233);
nor U44087 (N_44087,N_38855,N_36235);
nor U44088 (N_44088,N_39468,N_37295);
xnor U44089 (N_44089,N_37427,N_37730);
or U44090 (N_44090,N_38871,N_37012);
or U44091 (N_44091,N_39953,N_38343);
nor U44092 (N_44092,N_39620,N_39905);
nand U44093 (N_44093,N_36805,N_38432);
or U44094 (N_44094,N_39517,N_35804);
xor U44095 (N_44095,N_37151,N_38523);
and U44096 (N_44096,N_36815,N_38522);
xor U44097 (N_44097,N_38443,N_35308);
or U44098 (N_44098,N_38513,N_36263);
nor U44099 (N_44099,N_38085,N_35832);
and U44100 (N_44100,N_35837,N_36151);
nand U44101 (N_44101,N_38493,N_35445);
nand U44102 (N_44102,N_38513,N_38724);
nor U44103 (N_44103,N_38339,N_37811);
or U44104 (N_44104,N_37014,N_36535);
and U44105 (N_44105,N_37731,N_35609);
xor U44106 (N_44106,N_35881,N_36386);
or U44107 (N_44107,N_39588,N_36977);
or U44108 (N_44108,N_36892,N_37788);
xor U44109 (N_44109,N_39950,N_37487);
nand U44110 (N_44110,N_37683,N_37868);
or U44111 (N_44111,N_37777,N_37180);
xnor U44112 (N_44112,N_39132,N_37341);
xor U44113 (N_44113,N_35206,N_38679);
or U44114 (N_44114,N_36212,N_36739);
or U44115 (N_44115,N_36950,N_38283);
or U44116 (N_44116,N_36750,N_36063);
xor U44117 (N_44117,N_36885,N_35534);
and U44118 (N_44118,N_37537,N_39658);
xor U44119 (N_44119,N_39218,N_38983);
nand U44120 (N_44120,N_37674,N_35214);
or U44121 (N_44121,N_37194,N_39860);
nor U44122 (N_44122,N_37622,N_35848);
and U44123 (N_44123,N_38924,N_36179);
nand U44124 (N_44124,N_38298,N_39389);
or U44125 (N_44125,N_36197,N_38040);
nor U44126 (N_44126,N_35677,N_35260);
xor U44127 (N_44127,N_36949,N_37045);
or U44128 (N_44128,N_38823,N_37231);
nor U44129 (N_44129,N_36864,N_39131);
or U44130 (N_44130,N_36042,N_35579);
or U44131 (N_44131,N_39803,N_39873);
or U44132 (N_44132,N_35965,N_36527);
and U44133 (N_44133,N_36640,N_38068);
nor U44134 (N_44134,N_36051,N_38519);
and U44135 (N_44135,N_37745,N_39842);
nor U44136 (N_44136,N_36748,N_35542);
and U44137 (N_44137,N_35000,N_39639);
xnor U44138 (N_44138,N_36663,N_37471);
and U44139 (N_44139,N_37458,N_38748);
or U44140 (N_44140,N_39859,N_35164);
and U44141 (N_44141,N_39392,N_35842);
or U44142 (N_44142,N_37851,N_35805);
nand U44143 (N_44143,N_38926,N_35918);
nand U44144 (N_44144,N_39419,N_36601);
nand U44145 (N_44145,N_39499,N_38625);
or U44146 (N_44146,N_39187,N_37228);
nand U44147 (N_44147,N_35071,N_39269);
or U44148 (N_44148,N_37328,N_38527);
xor U44149 (N_44149,N_36734,N_35698);
nor U44150 (N_44150,N_36201,N_39517);
and U44151 (N_44151,N_35173,N_36947);
nor U44152 (N_44152,N_38697,N_37164);
or U44153 (N_44153,N_35052,N_37149);
and U44154 (N_44154,N_35717,N_39502);
nor U44155 (N_44155,N_35598,N_35076);
or U44156 (N_44156,N_36527,N_37287);
and U44157 (N_44157,N_37043,N_37186);
and U44158 (N_44158,N_36270,N_37329);
xor U44159 (N_44159,N_36518,N_38389);
or U44160 (N_44160,N_36990,N_39009);
or U44161 (N_44161,N_36747,N_37196);
xor U44162 (N_44162,N_38531,N_36071);
nand U44163 (N_44163,N_36383,N_39795);
nand U44164 (N_44164,N_36205,N_39922);
or U44165 (N_44165,N_38406,N_39825);
and U44166 (N_44166,N_36442,N_38118);
nand U44167 (N_44167,N_37137,N_37573);
nor U44168 (N_44168,N_38090,N_37922);
nor U44169 (N_44169,N_36766,N_35306);
nand U44170 (N_44170,N_36109,N_39565);
xnor U44171 (N_44171,N_35570,N_35166);
nor U44172 (N_44172,N_38137,N_36514);
or U44173 (N_44173,N_35354,N_36382);
and U44174 (N_44174,N_39328,N_39875);
or U44175 (N_44175,N_39774,N_37793);
nor U44176 (N_44176,N_39751,N_38172);
or U44177 (N_44177,N_38235,N_37579);
xnor U44178 (N_44178,N_39006,N_38310);
and U44179 (N_44179,N_37648,N_35609);
and U44180 (N_44180,N_37495,N_36995);
nor U44181 (N_44181,N_38534,N_36644);
nor U44182 (N_44182,N_39606,N_36684);
or U44183 (N_44183,N_39909,N_38131);
or U44184 (N_44184,N_35066,N_39778);
nor U44185 (N_44185,N_39197,N_39478);
nor U44186 (N_44186,N_38628,N_39848);
nand U44187 (N_44187,N_35447,N_39013);
nor U44188 (N_44188,N_37043,N_35970);
and U44189 (N_44189,N_39066,N_38270);
nor U44190 (N_44190,N_39391,N_36709);
nand U44191 (N_44191,N_36782,N_38040);
nand U44192 (N_44192,N_37189,N_36063);
and U44193 (N_44193,N_39568,N_35492);
and U44194 (N_44194,N_37923,N_36491);
xor U44195 (N_44195,N_36266,N_35416);
nor U44196 (N_44196,N_37210,N_39331);
or U44197 (N_44197,N_39713,N_35071);
and U44198 (N_44198,N_37394,N_37138);
or U44199 (N_44199,N_38471,N_38835);
nand U44200 (N_44200,N_38878,N_35710);
nand U44201 (N_44201,N_39052,N_35303);
xor U44202 (N_44202,N_39663,N_38189);
nand U44203 (N_44203,N_38593,N_39712);
or U44204 (N_44204,N_37538,N_38219);
or U44205 (N_44205,N_35779,N_36285);
and U44206 (N_44206,N_38002,N_39455);
and U44207 (N_44207,N_36845,N_35548);
nand U44208 (N_44208,N_38040,N_37622);
or U44209 (N_44209,N_38186,N_38202);
nor U44210 (N_44210,N_39026,N_36689);
nor U44211 (N_44211,N_38235,N_39834);
and U44212 (N_44212,N_38877,N_39056);
or U44213 (N_44213,N_38822,N_39291);
and U44214 (N_44214,N_35470,N_35404);
nand U44215 (N_44215,N_37258,N_38228);
or U44216 (N_44216,N_35802,N_38512);
and U44217 (N_44217,N_37940,N_37469);
nor U44218 (N_44218,N_37737,N_36601);
nor U44219 (N_44219,N_39652,N_37919);
or U44220 (N_44220,N_38406,N_38103);
and U44221 (N_44221,N_37198,N_39825);
nor U44222 (N_44222,N_38928,N_36842);
nand U44223 (N_44223,N_37416,N_35231);
xor U44224 (N_44224,N_37262,N_39704);
xnor U44225 (N_44225,N_39964,N_37297);
or U44226 (N_44226,N_39151,N_35355);
xnor U44227 (N_44227,N_36755,N_35102);
and U44228 (N_44228,N_39083,N_37862);
nand U44229 (N_44229,N_39581,N_37736);
nand U44230 (N_44230,N_37923,N_36219);
and U44231 (N_44231,N_36506,N_35350);
nor U44232 (N_44232,N_39767,N_35672);
or U44233 (N_44233,N_36780,N_35084);
nand U44234 (N_44234,N_37463,N_38015);
and U44235 (N_44235,N_38034,N_37628);
nand U44236 (N_44236,N_36986,N_38126);
nand U44237 (N_44237,N_37763,N_37618);
nand U44238 (N_44238,N_39626,N_37305);
or U44239 (N_44239,N_39606,N_39718);
or U44240 (N_44240,N_38398,N_36082);
and U44241 (N_44241,N_35322,N_36129);
and U44242 (N_44242,N_39368,N_38672);
and U44243 (N_44243,N_37278,N_36559);
xor U44244 (N_44244,N_39029,N_35601);
and U44245 (N_44245,N_38484,N_37832);
xor U44246 (N_44246,N_39812,N_37370);
and U44247 (N_44247,N_36893,N_39423);
and U44248 (N_44248,N_39791,N_36352);
or U44249 (N_44249,N_37594,N_35485);
nand U44250 (N_44250,N_39688,N_37808);
xor U44251 (N_44251,N_37813,N_35079);
or U44252 (N_44252,N_36328,N_39893);
nand U44253 (N_44253,N_37659,N_35901);
or U44254 (N_44254,N_35624,N_35945);
nand U44255 (N_44255,N_35365,N_38742);
nand U44256 (N_44256,N_39540,N_35445);
nand U44257 (N_44257,N_39730,N_36442);
nor U44258 (N_44258,N_36571,N_37676);
nand U44259 (N_44259,N_37501,N_38089);
xor U44260 (N_44260,N_39459,N_36703);
nor U44261 (N_44261,N_39019,N_36034);
nand U44262 (N_44262,N_36979,N_35774);
and U44263 (N_44263,N_36936,N_36342);
nor U44264 (N_44264,N_35742,N_39916);
nand U44265 (N_44265,N_38337,N_38370);
or U44266 (N_44266,N_35213,N_36394);
xor U44267 (N_44267,N_36700,N_36994);
nand U44268 (N_44268,N_39210,N_36206);
xor U44269 (N_44269,N_39232,N_35832);
and U44270 (N_44270,N_35371,N_35343);
and U44271 (N_44271,N_38917,N_39149);
or U44272 (N_44272,N_36941,N_38623);
and U44273 (N_44273,N_38770,N_35788);
xnor U44274 (N_44274,N_35251,N_37551);
and U44275 (N_44275,N_35681,N_35841);
xor U44276 (N_44276,N_36879,N_38574);
and U44277 (N_44277,N_35295,N_35577);
nor U44278 (N_44278,N_39474,N_35190);
or U44279 (N_44279,N_35305,N_36861);
nand U44280 (N_44280,N_37262,N_35461);
xor U44281 (N_44281,N_37379,N_36251);
nand U44282 (N_44282,N_38443,N_39980);
nand U44283 (N_44283,N_37015,N_35733);
nor U44284 (N_44284,N_39248,N_36769);
or U44285 (N_44285,N_36120,N_37868);
nand U44286 (N_44286,N_37856,N_35109);
nor U44287 (N_44287,N_35992,N_36041);
and U44288 (N_44288,N_39164,N_35634);
nand U44289 (N_44289,N_36332,N_35358);
nand U44290 (N_44290,N_36680,N_39650);
nand U44291 (N_44291,N_39699,N_36057);
nand U44292 (N_44292,N_38961,N_36781);
and U44293 (N_44293,N_36103,N_37538);
xor U44294 (N_44294,N_36742,N_37030);
or U44295 (N_44295,N_38435,N_38497);
nand U44296 (N_44296,N_36353,N_39364);
nor U44297 (N_44297,N_39524,N_37312);
nand U44298 (N_44298,N_39809,N_36336);
xnor U44299 (N_44299,N_35386,N_38285);
or U44300 (N_44300,N_35962,N_39797);
nor U44301 (N_44301,N_36777,N_36211);
and U44302 (N_44302,N_39795,N_36839);
and U44303 (N_44303,N_38764,N_35634);
nor U44304 (N_44304,N_35456,N_38666);
xor U44305 (N_44305,N_39123,N_36254);
nor U44306 (N_44306,N_37335,N_38435);
or U44307 (N_44307,N_36490,N_39099);
xnor U44308 (N_44308,N_36410,N_38225);
nor U44309 (N_44309,N_36658,N_37417);
nor U44310 (N_44310,N_37277,N_35484);
nor U44311 (N_44311,N_36333,N_37255);
and U44312 (N_44312,N_35008,N_36309);
nor U44313 (N_44313,N_37520,N_37650);
and U44314 (N_44314,N_35901,N_38634);
and U44315 (N_44315,N_38350,N_35997);
or U44316 (N_44316,N_35305,N_39520);
and U44317 (N_44317,N_38025,N_39952);
or U44318 (N_44318,N_35421,N_35240);
and U44319 (N_44319,N_38551,N_35782);
and U44320 (N_44320,N_35765,N_35078);
or U44321 (N_44321,N_36072,N_37795);
nand U44322 (N_44322,N_37615,N_37120);
nor U44323 (N_44323,N_37398,N_39643);
or U44324 (N_44324,N_38769,N_39329);
or U44325 (N_44325,N_36415,N_35136);
xor U44326 (N_44326,N_36689,N_35205);
nand U44327 (N_44327,N_39670,N_37454);
xnor U44328 (N_44328,N_35526,N_38459);
xor U44329 (N_44329,N_39718,N_35279);
nand U44330 (N_44330,N_37461,N_39508);
nand U44331 (N_44331,N_35048,N_36667);
or U44332 (N_44332,N_39747,N_36262);
xnor U44333 (N_44333,N_36922,N_37238);
nor U44334 (N_44334,N_36775,N_35867);
nand U44335 (N_44335,N_36955,N_36326);
or U44336 (N_44336,N_37830,N_37325);
or U44337 (N_44337,N_35185,N_37207);
nand U44338 (N_44338,N_35447,N_36579);
xor U44339 (N_44339,N_38042,N_39733);
or U44340 (N_44340,N_36445,N_36172);
xnor U44341 (N_44341,N_39760,N_35554);
xnor U44342 (N_44342,N_36649,N_36857);
nor U44343 (N_44343,N_37801,N_37552);
nor U44344 (N_44344,N_38572,N_38562);
and U44345 (N_44345,N_37626,N_38182);
nand U44346 (N_44346,N_36289,N_39085);
nand U44347 (N_44347,N_35294,N_37776);
nand U44348 (N_44348,N_38612,N_37601);
xor U44349 (N_44349,N_36394,N_35311);
and U44350 (N_44350,N_38094,N_36761);
or U44351 (N_44351,N_37181,N_37661);
nor U44352 (N_44352,N_38888,N_38096);
or U44353 (N_44353,N_38201,N_38961);
nor U44354 (N_44354,N_37552,N_37149);
nand U44355 (N_44355,N_36327,N_36628);
and U44356 (N_44356,N_35699,N_36077);
or U44357 (N_44357,N_37389,N_38596);
nand U44358 (N_44358,N_36475,N_39526);
xor U44359 (N_44359,N_39145,N_39053);
and U44360 (N_44360,N_39683,N_35257);
nor U44361 (N_44361,N_37269,N_38223);
nand U44362 (N_44362,N_37118,N_37140);
or U44363 (N_44363,N_37287,N_38546);
and U44364 (N_44364,N_38849,N_38552);
nor U44365 (N_44365,N_37035,N_37762);
nand U44366 (N_44366,N_39485,N_36167);
or U44367 (N_44367,N_38813,N_36896);
xor U44368 (N_44368,N_39180,N_37805);
xnor U44369 (N_44369,N_38064,N_36697);
xnor U44370 (N_44370,N_38527,N_39916);
and U44371 (N_44371,N_38116,N_38739);
nand U44372 (N_44372,N_35666,N_36524);
nor U44373 (N_44373,N_38242,N_39062);
nor U44374 (N_44374,N_38861,N_37389);
nor U44375 (N_44375,N_36287,N_38904);
nor U44376 (N_44376,N_37007,N_36793);
and U44377 (N_44377,N_36104,N_39783);
nor U44378 (N_44378,N_37716,N_37827);
or U44379 (N_44379,N_37880,N_36171);
xnor U44380 (N_44380,N_38956,N_36331);
or U44381 (N_44381,N_36402,N_38813);
xnor U44382 (N_44382,N_38854,N_37118);
xor U44383 (N_44383,N_37586,N_39002);
nor U44384 (N_44384,N_37362,N_38297);
and U44385 (N_44385,N_37880,N_39945);
or U44386 (N_44386,N_37391,N_36560);
or U44387 (N_44387,N_36665,N_36617);
and U44388 (N_44388,N_38578,N_38288);
xor U44389 (N_44389,N_38620,N_36280);
xnor U44390 (N_44390,N_39993,N_36140);
xnor U44391 (N_44391,N_38311,N_36415);
xnor U44392 (N_44392,N_39771,N_36948);
and U44393 (N_44393,N_38063,N_35672);
or U44394 (N_44394,N_38590,N_36698);
nand U44395 (N_44395,N_37154,N_37853);
and U44396 (N_44396,N_37731,N_35195);
and U44397 (N_44397,N_39357,N_39493);
xor U44398 (N_44398,N_35537,N_36453);
or U44399 (N_44399,N_37716,N_36176);
nor U44400 (N_44400,N_36518,N_38059);
and U44401 (N_44401,N_36338,N_39008);
and U44402 (N_44402,N_36508,N_39781);
and U44403 (N_44403,N_37002,N_39068);
nor U44404 (N_44404,N_39776,N_39453);
nand U44405 (N_44405,N_35768,N_35412);
nand U44406 (N_44406,N_35892,N_39478);
nor U44407 (N_44407,N_39754,N_36247);
and U44408 (N_44408,N_37090,N_37987);
or U44409 (N_44409,N_37624,N_38577);
xnor U44410 (N_44410,N_38926,N_35203);
xor U44411 (N_44411,N_36642,N_38081);
nor U44412 (N_44412,N_35550,N_39622);
xnor U44413 (N_44413,N_37225,N_35593);
and U44414 (N_44414,N_36855,N_36035);
nor U44415 (N_44415,N_36558,N_37654);
nor U44416 (N_44416,N_37024,N_38522);
or U44417 (N_44417,N_37915,N_37867);
xor U44418 (N_44418,N_39481,N_36886);
xor U44419 (N_44419,N_38406,N_36951);
xnor U44420 (N_44420,N_36975,N_36080);
nor U44421 (N_44421,N_38884,N_35151);
nor U44422 (N_44422,N_36369,N_36004);
and U44423 (N_44423,N_39070,N_38874);
and U44424 (N_44424,N_36192,N_38362);
xor U44425 (N_44425,N_36689,N_39087);
nand U44426 (N_44426,N_36110,N_37122);
or U44427 (N_44427,N_35736,N_36546);
and U44428 (N_44428,N_37880,N_35551);
nor U44429 (N_44429,N_35171,N_37219);
and U44430 (N_44430,N_37879,N_35572);
xnor U44431 (N_44431,N_38973,N_35454);
and U44432 (N_44432,N_38533,N_38556);
nand U44433 (N_44433,N_38476,N_38482);
nand U44434 (N_44434,N_35477,N_35040);
nand U44435 (N_44435,N_35234,N_35382);
nor U44436 (N_44436,N_37210,N_39192);
or U44437 (N_44437,N_38538,N_35338);
or U44438 (N_44438,N_39860,N_36859);
and U44439 (N_44439,N_39392,N_36730);
xor U44440 (N_44440,N_37025,N_39470);
nor U44441 (N_44441,N_39663,N_36293);
and U44442 (N_44442,N_37714,N_39918);
or U44443 (N_44443,N_38989,N_37863);
and U44444 (N_44444,N_37749,N_35845);
or U44445 (N_44445,N_35682,N_37176);
xor U44446 (N_44446,N_38502,N_38740);
nand U44447 (N_44447,N_37578,N_36179);
nor U44448 (N_44448,N_37441,N_36608);
or U44449 (N_44449,N_38682,N_36107);
xnor U44450 (N_44450,N_38618,N_38890);
and U44451 (N_44451,N_38305,N_36438);
or U44452 (N_44452,N_35945,N_39873);
and U44453 (N_44453,N_36355,N_38062);
or U44454 (N_44454,N_37952,N_35612);
nor U44455 (N_44455,N_38468,N_37945);
or U44456 (N_44456,N_37178,N_39375);
and U44457 (N_44457,N_36750,N_35875);
or U44458 (N_44458,N_36924,N_36530);
and U44459 (N_44459,N_37823,N_37812);
nand U44460 (N_44460,N_38554,N_35778);
or U44461 (N_44461,N_37751,N_37052);
and U44462 (N_44462,N_35992,N_35629);
xor U44463 (N_44463,N_35155,N_36145);
nand U44464 (N_44464,N_36579,N_37327);
or U44465 (N_44465,N_38004,N_39229);
nor U44466 (N_44466,N_37269,N_36100);
and U44467 (N_44467,N_36132,N_37516);
nor U44468 (N_44468,N_35884,N_36081);
and U44469 (N_44469,N_38546,N_37054);
nand U44470 (N_44470,N_37461,N_39166);
nand U44471 (N_44471,N_37603,N_39685);
or U44472 (N_44472,N_36768,N_37278);
xnor U44473 (N_44473,N_38398,N_38068);
nand U44474 (N_44474,N_37433,N_39780);
or U44475 (N_44475,N_38337,N_37569);
or U44476 (N_44476,N_35926,N_37906);
nand U44477 (N_44477,N_36966,N_37804);
and U44478 (N_44478,N_39989,N_35187);
xor U44479 (N_44479,N_38280,N_35292);
xor U44480 (N_44480,N_36966,N_35306);
and U44481 (N_44481,N_38503,N_39461);
and U44482 (N_44482,N_36435,N_36687);
and U44483 (N_44483,N_39901,N_39152);
nor U44484 (N_44484,N_39460,N_36643);
nor U44485 (N_44485,N_35084,N_38373);
and U44486 (N_44486,N_37953,N_36076);
nor U44487 (N_44487,N_38129,N_35413);
xor U44488 (N_44488,N_36205,N_38462);
and U44489 (N_44489,N_39664,N_37508);
or U44490 (N_44490,N_36668,N_39354);
or U44491 (N_44491,N_39825,N_36996);
nand U44492 (N_44492,N_37387,N_37731);
and U44493 (N_44493,N_37753,N_36223);
nand U44494 (N_44494,N_37582,N_37590);
nor U44495 (N_44495,N_35789,N_39432);
or U44496 (N_44496,N_35763,N_38309);
nor U44497 (N_44497,N_36343,N_35865);
or U44498 (N_44498,N_38645,N_39514);
nor U44499 (N_44499,N_36748,N_36450);
xnor U44500 (N_44500,N_38429,N_38244);
xnor U44501 (N_44501,N_35316,N_36979);
or U44502 (N_44502,N_35168,N_36912);
nand U44503 (N_44503,N_39715,N_36633);
and U44504 (N_44504,N_36879,N_36707);
or U44505 (N_44505,N_35614,N_36794);
or U44506 (N_44506,N_35068,N_35646);
nand U44507 (N_44507,N_37013,N_36338);
or U44508 (N_44508,N_36221,N_38315);
nor U44509 (N_44509,N_38302,N_39021);
or U44510 (N_44510,N_39383,N_38496);
nor U44511 (N_44511,N_37632,N_39091);
and U44512 (N_44512,N_36386,N_37216);
nand U44513 (N_44513,N_38306,N_35846);
nand U44514 (N_44514,N_39532,N_37128);
nor U44515 (N_44515,N_35014,N_37879);
nand U44516 (N_44516,N_36365,N_36756);
and U44517 (N_44517,N_35218,N_39016);
nand U44518 (N_44518,N_39468,N_37283);
or U44519 (N_44519,N_39981,N_36092);
and U44520 (N_44520,N_38798,N_38712);
nor U44521 (N_44521,N_36955,N_37455);
xnor U44522 (N_44522,N_36650,N_36460);
and U44523 (N_44523,N_39463,N_36370);
nand U44524 (N_44524,N_37378,N_39767);
nor U44525 (N_44525,N_39423,N_37599);
nor U44526 (N_44526,N_36816,N_36955);
nor U44527 (N_44527,N_36394,N_36436);
nand U44528 (N_44528,N_37241,N_38650);
nand U44529 (N_44529,N_37520,N_36589);
nand U44530 (N_44530,N_38334,N_35087);
xnor U44531 (N_44531,N_35039,N_35255);
and U44532 (N_44532,N_39737,N_37148);
nand U44533 (N_44533,N_37741,N_38883);
or U44534 (N_44534,N_36213,N_39435);
or U44535 (N_44535,N_37805,N_37699);
xor U44536 (N_44536,N_38088,N_37558);
nand U44537 (N_44537,N_38880,N_38735);
nand U44538 (N_44538,N_35793,N_36150);
xnor U44539 (N_44539,N_39640,N_38371);
nor U44540 (N_44540,N_37604,N_37354);
xor U44541 (N_44541,N_35975,N_38171);
nand U44542 (N_44542,N_35349,N_39504);
xnor U44543 (N_44543,N_38354,N_35517);
nand U44544 (N_44544,N_36775,N_39006);
or U44545 (N_44545,N_38617,N_39168);
and U44546 (N_44546,N_39406,N_35951);
or U44547 (N_44547,N_35906,N_37772);
xnor U44548 (N_44548,N_37088,N_37441);
xnor U44549 (N_44549,N_39862,N_38234);
and U44550 (N_44550,N_39240,N_36893);
nand U44551 (N_44551,N_36544,N_38101);
and U44552 (N_44552,N_38326,N_38288);
or U44553 (N_44553,N_39856,N_35091);
nand U44554 (N_44554,N_36961,N_36145);
nor U44555 (N_44555,N_38161,N_39740);
nand U44556 (N_44556,N_38339,N_36350);
and U44557 (N_44557,N_38635,N_36982);
and U44558 (N_44558,N_39059,N_36743);
nor U44559 (N_44559,N_36385,N_39569);
nand U44560 (N_44560,N_39558,N_39799);
nor U44561 (N_44561,N_37495,N_37981);
and U44562 (N_44562,N_37165,N_36223);
nand U44563 (N_44563,N_35121,N_37606);
nor U44564 (N_44564,N_39156,N_37746);
nand U44565 (N_44565,N_35900,N_36386);
or U44566 (N_44566,N_39559,N_38946);
nor U44567 (N_44567,N_38534,N_38992);
xor U44568 (N_44568,N_38670,N_38005);
nand U44569 (N_44569,N_39534,N_38000);
or U44570 (N_44570,N_38816,N_39712);
nor U44571 (N_44571,N_37667,N_38375);
nor U44572 (N_44572,N_39407,N_36943);
and U44573 (N_44573,N_38236,N_39105);
or U44574 (N_44574,N_35718,N_35658);
xnor U44575 (N_44575,N_35759,N_35980);
and U44576 (N_44576,N_37605,N_35887);
nand U44577 (N_44577,N_35010,N_36753);
xor U44578 (N_44578,N_39538,N_37908);
nand U44579 (N_44579,N_38419,N_39363);
and U44580 (N_44580,N_36197,N_35164);
nor U44581 (N_44581,N_37481,N_36826);
and U44582 (N_44582,N_38787,N_35620);
xor U44583 (N_44583,N_35125,N_36537);
nand U44584 (N_44584,N_35327,N_35356);
or U44585 (N_44585,N_39670,N_39462);
nor U44586 (N_44586,N_36225,N_37211);
nand U44587 (N_44587,N_36615,N_35263);
and U44588 (N_44588,N_36569,N_38689);
nor U44589 (N_44589,N_36971,N_38690);
nand U44590 (N_44590,N_39901,N_36433);
or U44591 (N_44591,N_35014,N_39176);
or U44592 (N_44592,N_38356,N_37806);
and U44593 (N_44593,N_37797,N_37091);
and U44594 (N_44594,N_36134,N_36794);
or U44595 (N_44595,N_39750,N_39248);
nand U44596 (N_44596,N_39739,N_38458);
xor U44597 (N_44597,N_37657,N_39287);
nor U44598 (N_44598,N_37499,N_37707);
xnor U44599 (N_44599,N_36431,N_36085);
xnor U44600 (N_44600,N_35027,N_39073);
nor U44601 (N_44601,N_36493,N_35374);
nor U44602 (N_44602,N_36167,N_38186);
nand U44603 (N_44603,N_37602,N_38261);
nor U44604 (N_44604,N_36545,N_39722);
or U44605 (N_44605,N_37417,N_39574);
nand U44606 (N_44606,N_35065,N_35823);
nor U44607 (N_44607,N_35873,N_35481);
nor U44608 (N_44608,N_35140,N_38700);
nor U44609 (N_44609,N_38290,N_39217);
nor U44610 (N_44610,N_36195,N_39741);
nor U44611 (N_44611,N_37595,N_35805);
xnor U44612 (N_44612,N_37817,N_35178);
or U44613 (N_44613,N_37389,N_37652);
xnor U44614 (N_44614,N_37521,N_38731);
or U44615 (N_44615,N_36518,N_39132);
xnor U44616 (N_44616,N_37203,N_35125);
or U44617 (N_44617,N_39756,N_37830);
and U44618 (N_44618,N_37466,N_37989);
or U44619 (N_44619,N_39451,N_35410);
nor U44620 (N_44620,N_37150,N_35931);
and U44621 (N_44621,N_37243,N_38013);
and U44622 (N_44622,N_37948,N_35711);
nand U44623 (N_44623,N_37164,N_38775);
xnor U44624 (N_44624,N_36065,N_39640);
nor U44625 (N_44625,N_38473,N_39318);
nor U44626 (N_44626,N_38897,N_35966);
or U44627 (N_44627,N_39877,N_37266);
and U44628 (N_44628,N_39120,N_35070);
xnor U44629 (N_44629,N_38986,N_37321);
nor U44630 (N_44630,N_36237,N_36995);
xor U44631 (N_44631,N_38768,N_39762);
and U44632 (N_44632,N_39651,N_37485);
nand U44633 (N_44633,N_37315,N_35780);
nor U44634 (N_44634,N_35305,N_36873);
nor U44635 (N_44635,N_38069,N_36025);
or U44636 (N_44636,N_38505,N_35824);
and U44637 (N_44637,N_37153,N_37889);
nand U44638 (N_44638,N_36180,N_37670);
or U44639 (N_44639,N_35483,N_35464);
nand U44640 (N_44640,N_35527,N_36746);
and U44641 (N_44641,N_37545,N_39149);
nand U44642 (N_44642,N_37276,N_37408);
and U44643 (N_44643,N_37914,N_37533);
nor U44644 (N_44644,N_39255,N_38515);
nor U44645 (N_44645,N_37459,N_37199);
xor U44646 (N_44646,N_38302,N_36989);
xor U44647 (N_44647,N_36210,N_39503);
and U44648 (N_44648,N_37963,N_39590);
nor U44649 (N_44649,N_37875,N_37758);
or U44650 (N_44650,N_35657,N_38008);
nor U44651 (N_44651,N_36565,N_38482);
or U44652 (N_44652,N_35919,N_38943);
xor U44653 (N_44653,N_36220,N_36552);
and U44654 (N_44654,N_38951,N_38604);
xnor U44655 (N_44655,N_37437,N_37646);
or U44656 (N_44656,N_37904,N_35653);
xnor U44657 (N_44657,N_37685,N_38172);
nand U44658 (N_44658,N_37855,N_38076);
nor U44659 (N_44659,N_37503,N_36665);
xnor U44660 (N_44660,N_36974,N_38022);
nand U44661 (N_44661,N_38888,N_39740);
nor U44662 (N_44662,N_36531,N_36821);
nand U44663 (N_44663,N_36137,N_36314);
nand U44664 (N_44664,N_36329,N_35038);
nand U44665 (N_44665,N_38229,N_39831);
or U44666 (N_44666,N_35954,N_35695);
and U44667 (N_44667,N_37132,N_39351);
nand U44668 (N_44668,N_37859,N_36895);
nand U44669 (N_44669,N_39252,N_35539);
nand U44670 (N_44670,N_36769,N_36479);
or U44671 (N_44671,N_35127,N_37518);
nor U44672 (N_44672,N_35054,N_37764);
nor U44673 (N_44673,N_38444,N_38686);
nor U44674 (N_44674,N_39360,N_35335);
xnor U44675 (N_44675,N_35352,N_37041);
nor U44676 (N_44676,N_35755,N_39977);
and U44677 (N_44677,N_39235,N_35810);
nand U44678 (N_44678,N_38908,N_38834);
xor U44679 (N_44679,N_39026,N_35863);
or U44680 (N_44680,N_35881,N_36507);
nand U44681 (N_44681,N_35760,N_39474);
nor U44682 (N_44682,N_35377,N_35958);
or U44683 (N_44683,N_35820,N_37776);
or U44684 (N_44684,N_39037,N_36873);
and U44685 (N_44685,N_36662,N_36001);
nand U44686 (N_44686,N_37902,N_35627);
nand U44687 (N_44687,N_36890,N_37199);
nand U44688 (N_44688,N_38321,N_37984);
nand U44689 (N_44689,N_36417,N_38056);
nor U44690 (N_44690,N_35379,N_36338);
and U44691 (N_44691,N_37469,N_38550);
nor U44692 (N_44692,N_37198,N_35482);
or U44693 (N_44693,N_39031,N_35399);
nor U44694 (N_44694,N_38365,N_35633);
nand U44695 (N_44695,N_36829,N_35861);
and U44696 (N_44696,N_35594,N_36997);
xor U44697 (N_44697,N_38219,N_38626);
nand U44698 (N_44698,N_38984,N_35078);
xor U44699 (N_44699,N_37582,N_35146);
or U44700 (N_44700,N_37133,N_36549);
xor U44701 (N_44701,N_37114,N_38489);
and U44702 (N_44702,N_37845,N_37227);
or U44703 (N_44703,N_37624,N_36576);
xnor U44704 (N_44704,N_35982,N_37162);
or U44705 (N_44705,N_36069,N_38035);
or U44706 (N_44706,N_35427,N_38509);
nand U44707 (N_44707,N_36808,N_36791);
nand U44708 (N_44708,N_36223,N_38091);
nor U44709 (N_44709,N_35053,N_38789);
and U44710 (N_44710,N_35780,N_36848);
nor U44711 (N_44711,N_37681,N_35590);
nor U44712 (N_44712,N_38770,N_39828);
nand U44713 (N_44713,N_35637,N_36899);
nor U44714 (N_44714,N_35726,N_36713);
or U44715 (N_44715,N_35563,N_35425);
xnor U44716 (N_44716,N_39161,N_39273);
and U44717 (N_44717,N_37152,N_37953);
xnor U44718 (N_44718,N_35116,N_39165);
nand U44719 (N_44719,N_35574,N_39741);
or U44720 (N_44720,N_37553,N_37108);
or U44721 (N_44721,N_35594,N_39537);
nand U44722 (N_44722,N_38457,N_36294);
nor U44723 (N_44723,N_39034,N_37387);
and U44724 (N_44724,N_37953,N_39077);
or U44725 (N_44725,N_39274,N_39334);
xnor U44726 (N_44726,N_36265,N_37458);
or U44727 (N_44727,N_35438,N_36632);
nand U44728 (N_44728,N_37601,N_38516);
nand U44729 (N_44729,N_37156,N_35088);
nor U44730 (N_44730,N_38739,N_38554);
or U44731 (N_44731,N_37629,N_37236);
or U44732 (N_44732,N_38210,N_39522);
nor U44733 (N_44733,N_38321,N_35201);
nand U44734 (N_44734,N_35030,N_38539);
xnor U44735 (N_44735,N_36249,N_39687);
nor U44736 (N_44736,N_39929,N_39911);
or U44737 (N_44737,N_38407,N_36933);
or U44738 (N_44738,N_35014,N_36745);
nor U44739 (N_44739,N_39586,N_35422);
xor U44740 (N_44740,N_38638,N_36695);
nand U44741 (N_44741,N_38527,N_36433);
nand U44742 (N_44742,N_35545,N_36347);
or U44743 (N_44743,N_35037,N_38042);
and U44744 (N_44744,N_35225,N_36828);
and U44745 (N_44745,N_35222,N_37718);
and U44746 (N_44746,N_39864,N_39382);
xnor U44747 (N_44747,N_39797,N_36444);
nor U44748 (N_44748,N_39687,N_39450);
or U44749 (N_44749,N_37961,N_35435);
and U44750 (N_44750,N_35105,N_38450);
nor U44751 (N_44751,N_39563,N_37052);
nor U44752 (N_44752,N_39396,N_38635);
or U44753 (N_44753,N_36508,N_38771);
nand U44754 (N_44754,N_37787,N_35484);
or U44755 (N_44755,N_37655,N_36275);
xor U44756 (N_44756,N_38931,N_39220);
or U44757 (N_44757,N_38434,N_39177);
nor U44758 (N_44758,N_36634,N_39174);
and U44759 (N_44759,N_37976,N_39304);
and U44760 (N_44760,N_35606,N_37094);
and U44761 (N_44761,N_39527,N_36125);
nand U44762 (N_44762,N_38824,N_38614);
or U44763 (N_44763,N_35412,N_36881);
xor U44764 (N_44764,N_38218,N_37363);
nor U44765 (N_44765,N_38333,N_35152);
and U44766 (N_44766,N_38163,N_39016);
nor U44767 (N_44767,N_36865,N_36778);
nand U44768 (N_44768,N_36914,N_39106);
or U44769 (N_44769,N_35074,N_39771);
nand U44770 (N_44770,N_37324,N_39560);
and U44771 (N_44771,N_38657,N_37803);
and U44772 (N_44772,N_37917,N_39017);
xor U44773 (N_44773,N_35903,N_38775);
or U44774 (N_44774,N_38829,N_36085);
nand U44775 (N_44775,N_37795,N_39271);
xor U44776 (N_44776,N_35361,N_35326);
nand U44777 (N_44777,N_38069,N_39667);
nor U44778 (N_44778,N_35560,N_36956);
xnor U44779 (N_44779,N_38158,N_35621);
xnor U44780 (N_44780,N_38821,N_35806);
nor U44781 (N_44781,N_39349,N_39162);
nor U44782 (N_44782,N_38513,N_37137);
nand U44783 (N_44783,N_36251,N_35846);
or U44784 (N_44784,N_35408,N_35820);
xnor U44785 (N_44785,N_38343,N_36236);
nor U44786 (N_44786,N_36510,N_36692);
nand U44787 (N_44787,N_37057,N_38665);
nand U44788 (N_44788,N_39777,N_37572);
and U44789 (N_44789,N_36898,N_36231);
xnor U44790 (N_44790,N_38600,N_36910);
or U44791 (N_44791,N_38431,N_37539);
xor U44792 (N_44792,N_39999,N_39732);
nor U44793 (N_44793,N_35965,N_37796);
and U44794 (N_44794,N_37952,N_35014);
or U44795 (N_44795,N_39944,N_36117);
or U44796 (N_44796,N_35971,N_39283);
nand U44797 (N_44797,N_35184,N_39953);
or U44798 (N_44798,N_37717,N_37741);
and U44799 (N_44799,N_35194,N_39952);
xnor U44800 (N_44800,N_37242,N_37170);
xnor U44801 (N_44801,N_37471,N_37294);
nor U44802 (N_44802,N_35004,N_38199);
or U44803 (N_44803,N_36789,N_39253);
and U44804 (N_44804,N_37524,N_39990);
or U44805 (N_44805,N_36347,N_35895);
xor U44806 (N_44806,N_35686,N_37932);
nor U44807 (N_44807,N_36611,N_38139);
and U44808 (N_44808,N_37619,N_35120);
and U44809 (N_44809,N_37582,N_35789);
xor U44810 (N_44810,N_38798,N_36213);
nand U44811 (N_44811,N_38851,N_36997);
nand U44812 (N_44812,N_38357,N_39791);
or U44813 (N_44813,N_35379,N_38959);
xor U44814 (N_44814,N_37826,N_35698);
nand U44815 (N_44815,N_39364,N_39909);
nand U44816 (N_44816,N_37382,N_38235);
or U44817 (N_44817,N_35050,N_37918);
and U44818 (N_44818,N_35523,N_38388);
nand U44819 (N_44819,N_35608,N_35525);
xor U44820 (N_44820,N_38979,N_39915);
or U44821 (N_44821,N_36294,N_38388);
nand U44822 (N_44822,N_39727,N_37235);
nor U44823 (N_44823,N_38198,N_36115);
and U44824 (N_44824,N_38535,N_37135);
and U44825 (N_44825,N_39526,N_37967);
nand U44826 (N_44826,N_36449,N_37124);
nor U44827 (N_44827,N_38109,N_37283);
nor U44828 (N_44828,N_38492,N_38226);
and U44829 (N_44829,N_39173,N_39736);
nor U44830 (N_44830,N_37562,N_39052);
and U44831 (N_44831,N_38370,N_37756);
or U44832 (N_44832,N_39074,N_37394);
nor U44833 (N_44833,N_39174,N_36312);
or U44834 (N_44834,N_39569,N_35758);
nand U44835 (N_44835,N_36439,N_36824);
nand U44836 (N_44836,N_38214,N_39039);
nor U44837 (N_44837,N_38632,N_35646);
and U44838 (N_44838,N_39833,N_38186);
xor U44839 (N_44839,N_35567,N_35596);
nor U44840 (N_44840,N_37761,N_37986);
xor U44841 (N_44841,N_37629,N_38787);
xnor U44842 (N_44842,N_37591,N_35417);
xor U44843 (N_44843,N_37341,N_36114);
nor U44844 (N_44844,N_38228,N_39532);
or U44845 (N_44845,N_38653,N_36534);
nand U44846 (N_44846,N_35508,N_35297);
nand U44847 (N_44847,N_36224,N_39375);
xnor U44848 (N_44848,N_39784,N_38961);
nor U44849 (N_44849,N_35472,N_36200);
and U44850 (N_44850,N_37068,N_38924);
xor U44851 (N_44851,N_38383,N_38858);
or U44852 (N_44852,N_38062,N_38791);
nand U44853 (N_44853,N_37361,N_36901);
nor U44854 (N_44854,N_35728,N_35966);
nand U44855 (N_44855,N_35777,N_36029);
nand U44856 (N_44856,N_35444,N_35341);
and U44857 (N_44857,N_37196,N_38377);
xor U44858 (N_44858,N_39344,N_39166);
xnor U44859 (N_44859,N_38658,N_38100);
xor U44860 (N_44860,N_39084,N_38365);
or U44861 (N_44861,N_35448,N_36333);
and U44862 (N_44862,N_39472,N_36938);
xnor U44863 (N_44863,N_36756,N_37252);
and U44864 (N_44864,N_38503,N_38688);
nor U44865 (N_44865,N_37699,N_38390);
nand U44866 (N_44866,N_36577,N_38357);
or U44867 (N_44867,N_39807,N_35141);
nor U44868 (N_44868,N_36339,N_38690);
or U44869 (N_44869,N_38737,N_37698);
nor U44870 (N_44870,N_37482,N_39092);
and U44871 (N_44871,N_37698,N_36485);
nor U44872 (N_44872,N_37074,N_37394);
or U44873 (N_44873,N_38941,N_36580);
and U44874 (N_44874,N_36206,N_35142);
and U44875 (N_44875,N_35923,N_36094);
or U44876 (N_44876,N_39926,N_38764);
and U44877 (N_44877,N_38866,N_35453);
nor U44878 (N_44878,N_37593,N_35873);
nor U44879 (N_44879,N_35787,N_39185);
or U44880 (N_44880,N_38294,N_39427);
nand U44881 (N_44881,N_35284,N_36648);
and U44882 (N_44882,N_39488,N_38452);
nand U44883 (N_44883,N_38195,N_35563);
xnor U44884 (N_44884,N_35638,N_37949);
or U44885 (N_44885,N_37089,N_36013);
and U44886 (N_44886,N_37856,N_35359);
and U44887 (N_44887,N_36349,N_39533);
and U44888 (N_44888,N_38959,N_36954);
xor U44889 (N_44889,N_39602,N_35368);
or U44890 (N_44890,N_35719,N_36924);
nand U44891 (N_44891,N_36101,N_36491);
and U44892 (N_44892,N_35051,N_37937);
xor U44893 (N_44893,N_37542,N_36108);
nand U44894 (N_44894,N_38057,N_36102);
and U44895 (N_44895,N_37764,N_39155);
or U44896 (N_44896,N_36500,N_36383);
xnor U44897 (N_44897,N_39169,N_36452);
nor U44898 (N_44898,N_38531,N_37961);
or U44899 (N_44899,N_39107,N_36532);
or U44900 (N_44900,N_38532,N_37836);
xnor U44901 (N_44901,N_38991,N_37351);
nor U44902 (N_44902,N_36853,N_37547);
xnor U44903 (N_44903,N_39341,N_39058);
or U44904 (N_44904,N_35878,N_39393);
or U44905 (N_44905,N_39580,N_38458);
nand U44906 (N_44906,N_35938,N_39042);
nor U44907 (N_44907,N_35812,N_36013);
or U44908 (N_44908,N_35867,N_38153);
and U44909 (N_44909,N_37365,N_39395);
or U44910 (N_44910,N_37790,N_35103);
nand U44911 (N_44911,N_39969,N_37177);
nor U44912 (N_44912,N_39149,N_39264);
nor U44913 (N_44913,N_35236,N_38244);
nand U44914 (N_44914,N_38179,N_39391);
nor U44915 (N_44915,N_35779,N_35232);
xor U44916 (N_44916,N_37435,N_38998);
and U44917 (N_44917,N_36539,N_36397);
nor U44918 (N_44918,N_35724,N_36009);
nand U44919 (N_44919,N_35086,N_35180);
and U44920 (N_44920,N_38635,N_36582);
nand U44921 (N_44921,N_38173,N_38484);
xnor U44922 (N_44922,N_38112,N_35766);
xor U44923 (N_44923,N_35910,N_36686);
nand U44924 (N_44924,N_37656,N_35548);
and U44925 (N_44925,N_36532,N_38111);
or U44926 (N_44926,N_35228,N_39998);
or U44927 (N_44927,N_38339,N_35817);
or U44928 (N_44928,N_36510,N_36553);
nor U44929 (N_44929,N_38206,N_39719);
and U44930 (N_44930,N_39630,N_39785);
xnor U44931 (N_44931,N_36981,N_35496);
nand U44932 (N_44932,N_39140,N_37474);
or U44933 (N_44933,N_39546,N_37239);
xor U44934 (N_44934,N_36274,N_39721);
and U44935 (N_44935,N_38729,N_36284);
nand U44936 (N_44936,N_37794,N_36567);
xor U44937 (N_44937,N_35835,N_36163);
or U44938 (N_44938,N_37719,N_38484);
xnor U44939 (N_44939,N_35554,N_37155);
xnor U44940 (N_44940,N_36981,N_39421);
and U44941 (N_44941,N_37064,N_37025);
nor U44942 (N_44942,N_39231,N_38457);
nand U44943 (N_44943,N_38988,N_38232);
nand U44944 (N_44944,N_39371,N_36713);
nor U44945 (N_44945,N_35988,N_35791);
nor U44946 (N_44946,N_38889,N_36896);
nor U44947 (N_44947,N_38494,N_39046);
nand U44948 (N_44948,N_36972,N_37436);
xnor U44949 (N_44949,N_36300,N_38016);
or U44950 (N_44950,N_38723,N_36386);
nor U44951 (N_44951,N_37266,N_39590);
nor U44952 (N_44952,N_39558,N_36038);
nor U44953 (N_44953,N_37187,N_35442);
nor U44954 (N_44954,N_36565,N_36184);
and U44955 (N_44955,N_36897,N_38432);
nand U44956 (N_44956,N_35066,N_37832);
or U44957 (N_44957,N_37555,N_38510);
or U44958 (N_44958,N_38374,N_36989);
or U44959 (N_44959,N_36464,N_35366);
nand U44960 (N_44960,N_37360,N_35198);
xnor U44961 (N_44961,N_39762,N_37358);
or U44962 (N_44962,N_36366,N_36223);
nor U44963 (N_44963,N_37686,N_35551);
xor U44964 (N_44964,N_38824,N_35730);
nand U44965 (N_44965,N_36187,N_38070);
xnor U44966 (N_44966,N_37109,N_36004);
xor U44967 (N_44967,N_38149,N_38872);
and U44968 (N_44968,N_37838,N_38585);
and U44969 (N_44969,N_37998,N_39328);
xnor U44970 (N_44970,N_39835,N_38104);
xor U44971 (N_44971,N_36821,N_39506);
nand U44972 (N_44972,N_39800,N_35723);
nand U44973 (N_44973,N_38104,N_39431);
xor U44974 (N_44974,N_37088,N_35831);
nand U44975 (N_44975,N_37355,N_38457);
xnor U44976 (N_44976,N_38847,N_36177);
nor U44977 (N_44977,N_38450,N_36961);
xnor U44978 (N_44978,N_36218,N_39288);
or U44979 (N_44979,N_38246,N_37192);
or U44980 (N_44980,N_38442,N_37414);
xor U44981 (N_44981,N_37633,N_37794);
nor U44982 (N_44982,N_35028,N_38474);
and U44983 (N_44983,N_35165,N_37810);
nand U44984 (N_44984,N_36231,N_38878);
and U44985 (N_44985,N_35975,N_35551);
and U44986 (N_44986,N_37080,N_36024);
xnor U44987 (N_44987,N_35607,N_37089);
or U44988 (N_44988,N_36215,N_36807);
and U44989 (N_44989,N_38186,N_39801);
nor U44990 (N_44990,N_36582,N_39649);
and U44991 (N_44991,N_35455,N_37480);
or U44992 (N_44992,N_39186,N_39523);
nand U44993 (N_44993,N_39650,N_37188);
nor U44994 (N_44994,N_37184,N_36169);
or U44995 (N_44995,N_35166,N_38483);
nand U44996 (N_44996,N_37418,N_35526);
xnor U44997 (N_44997,N_37346,N_38183);
xor U44998 (N_44998,N_37709,N_38045);
or U44999 (N_44999,N_37322,N_36224);
or U45000 (N_45000,N_41433,N_44496);
and U45001 (N_45001,N_42361,N_42861);
or U45002 (N_45002,N_41550,N_40743);
or U45003 (N_45003,N_43766,N_44489);
or U45004 (N_45004,N_44666,N_42642);
or U45005 (N_45005,N_43130,N_42452);
nor U45006 (N_45006,N_41650,N_41792);
xnor U45007 (N_45007,N_41221,N_40197);
nor U45008 (N_45008,N_42946,N_43344);
nor U45009 (N_45009,N_41220,N_43887);
xor U45010 (N_45010,N_41463,N_44890);
nand U45011 (N_45011,N_44031,N_40703);
or U45012 (N_45012,N_42271,N_43245);
nand U45013 (N_45013,N_40740,N_43394);
xor U45014 (N_45014,N_41021,N_41479);
and U45015 (N_45015,N_44994,N_42535);
nand U45016 (N_45016,N_41873,N_44225);
or U45017 (N_45017,N_41342,N_42560);
or U45018 (N_45018,N_43131,N_41471);
nor U45019 (N_45019,N_40512,N_40771);
or U45020 (N_45020,N_44485,N_41632);
nor U45021 (N_45021,N_44852,N_44613);
or U45022 (N_45022,N_40144,N_41834);
or U45023 (N_45023,N_43443,N_44174);
nor U45024 (N_45024,N_44744,N_42230);
or U45025 (N_45025,N_40358,N_43060);
nand U45026 (N_45026,N_41399,N_40220);
nand U45027 (N_45027,N_42791,N_42103);
nor U45028 (N_45028,N_42729,N_44332);
nand U45029 (N_45029,N_42493,N_40010);
xor U45030 (N_45030,N_41435,N_42462);
xor U45031 (N_45031,N_40023,N_41974);
xor U45032 (N_45032,N_41907,N_41567);
xnor U45033 (N_45033,N_43108,N_42239);
nor U45034 (N_45034,N_41752,N_40605);
nor U45035 (N_45035,N_41276,N_40606);
nor U45036 (N_45036,N_41770,N_41110);
and U45037 (N_45037,N_43189,N_44090);
nor U45038 (N_45038,N_40819,N_40151);
nor U45039 (N_45039,N_42099,N_40398);
and U45040 (N_45040,N_40631,N_42305);
or U45041 (N_45041,N_41505,N_40071);
xnor U45042 (N_45042,N_43603,N_42682);
and U45043 (N_45043,N_42996,N_41185);
xnor U45044 (N_45044,N_40239,N_42189);
nand U45045 (N_45045,N_42685,N_44961);
or U45046 (N_45046,N_41558,N_40135);
or U45047 (N_45047,N_41118,N_41261);
nand U45048 (N_45048,N_40416,N_42628);
nand U45049 (N_45049,N_42436,N_42908);
xor U45050 (N_45050,N_40537,N_40850);
and U45051 (N_45051,N_43611,N_44635);
or U45052 (N_45052,N_41100,N_41436);
xnor U45053 (N_45053,N_44384,N_43963);
and U45054 (N_45054,N_42592,N_43264);
or U45055 (N_45055,N_42926,N_43505);
and U45056 (N_45056,N_43370,N_44997);
nand U45057 (N_45057,N_42767,N_41078);
nand U45058 (N_45058,N_40190,N_41379);
nor U45059 (N_45059,N_41251,N_44142);
xor U45060 (N_45060,N_44520,N_44980);
nor U45061 (N_45061,N_41778,N_42526);
or U45062 (N_45062,N_42033,N_43573);
or U45063 (N_45063,N_41538,N_42384);
nand U45064 (N_45064,N_40293,N_40435);
or U45065 (N_45065,N_43374,N_43751);
or U45066 (N_45066,N_43989,N_42427);
and U45067 (N_45067,N_43973,N_40422);
and U45068 (N_45068,N_41853,N_43786);
nor U45069 (N_45069,N_43492,N_43268);
nand U45070 (N_45070,N_44071,N_40470);
nor U45071 (N_45071,N_43087,N_40581);
nand U45072 (N_45072,N_44558,N_44220);
nand U45073 (N_45073,N_44781,N_43064);
nand U45074 (N_45074,N_43898,N_42837);
nor U45075 (N_45075,N_41204,N_42575);
or U45076 (N_45076,N_42788,N_41697);
and U45077 (N_45077,N_43544,N_43826);
nand U45078 (N_45078,N_40322,N_40074);
nand U45079 (N_45079,N_43210,N_42419);
and U45080 (N_45080,N_44417,N_40951);
xor U45081 (N_45081,N_44521,N_41037);
or U45082 (N_45082,N_43650,N_41941);
and U45083 (N_45083,N_41687,N_43450);
nor U45084 (N_45084,N_44081,N_40112);
xor U45085 (N_45085,N_41267,N_42985);
nand U45086 (N_45086,N_40738,N_43322);
or U45087 (N_45087,N_44568,N_43534);
xor U45088 (N_45088,N_44293,N_41361);
or U45089 (N_45089,N_43749,N_41010);
and U45090 (N_45090,N_40718,N_41564);
and U45091 (N_45091,N_44894,N_42613);
xor U45092 (N_45092,N_40615,N_42794);
and U45093 (N_45093,N_44300,N_43678);
and U45094 (N_45094,N_41408,N_40733);
xor U45095 (N_45095,N_41540,N_41349);
xor U45096 (N_45096,N_44963,N_42118);
nand U45097 (N_45097,N_41732,N_43366);
and U45098 (N_45098,N_41786,N_41020);
xor U45099 (N_45099,N_43148,N_40042);
or U45100 (N_45100,N_44414,N_43985);
nor U45101 (N_45101,N_44787,N_41248);
xnor U45102 (N_45102,N_42517,N_44574);
nand U45103 (N_45103,N_41059,N_43696);
xnor U45104 (N_45104,N_43385,N_41457);
nand U45105 (N_45105,N_42223,N_40651);
or U45106 (N_45106,N_40421,N_41655);
and U45107 (N_45107,N_40305,N_43454);
xnor U45108 (N_45108,N_42124,N_41129);
and U45109 (N_45109,N_42913,N_42536);
xnor U45110 (N_45110,N_43888,N_40759);
or U45111 (N_45111,N_44572,N_40570);
or U45112 (N_45112,N_43354,N_42078);
xor U45113 (N_45113,N_43185,N_42705);
nand U45114 (N_45114,N_44340,N_40063);
xnor U45115 (N_45115,N_43251,N_41278);
xor U45116 (N_45116,N_43035,N_41948);
or U45117 (N_45117,N_41288,N_44383);
and U45118 (N_45118,N_42978,N_44027);
xor U45119 (N_45119,N_43029,N_42081);
and U45120 (N_45120,N_42332,N_44625);
or U45121 (N_45121,N_44688,N_40451);
nand U45122 (N_45122,N_41289,N_41430);
xnor U45123 (N_45123,N_43367,N_41231);
or U45124 (N_45124,N_41054,N_44169);
xor U45125 (N_45125,N_41504,N_42066);
nor U45126 (N_45126,N_43875,N_41242);
or U45127 (N_45127,N_44830,N_40404);
xor U45128 (N_45128,N_43904,N_40812);
or U45129 (N_45129,N_44874,N_40228);
nand U45130 (N_45130,N_43353,N_44887);
nand U45131 (N_45131,N_40194,N_41742);
or U45132 (N_45132,N_43209,N_42145);
xnor U45133 (N_45133,N_43738,N_43926);
xnor U45134 (N_45134,N_40287,N_43164);
nand U45135 (N_45135,N_43843,N_42654);
nand U45136 (N_45136,N_41958,N_44735);
nor U45137 (N_45137,N_40386,N_42465);
nand U45138 (N_45138,N_43255,N_42894);
nand U45139 (N_45139,N_40900,N_41704);
and U45140 (N_45140,N_40060,N_43677);
xor U45141 (N_45141,N_41817,N_41145);
and U45142 (N_45142,N_41382,N_44705);
xor U45143 (N_45143,N_42382,N_41611);
and U45144 (N_45144,N_42021,N_43760);
nand U45145 (N_45145,N_42292,N_42525);
or U45146 (N_45146,N_41336,N_43540);
xor U45147 (N_45147,N_40321,N_42570);
nor U45148 (N_45148,N_42780,N_43566);
nand U45149 (N_45149,N_43393,N_44038);
nand U45150 (N_45150,N_41138,N_42012);
and U45151 (N_45151,N_40656,N_44540);
and U45152 (N_45152,N_40936,N_41956);
nand U45153 (N_45153,N_43339,N_44942);
xor U45154 (N_45154,N_40028,N_41648);
or U45155 (N_45155,N_44073,N_44776);
nor U45156 (N_45156,N_43277,N_43978);
and U45157 (N_45157,N_41940,N_43088);
and U45158 (N_45158,N_41406,N_43300);
and U45159 (N_45159,N_42387,N_40344);
nand U45160 (N_45160,N_44179,N_44708);
nand U45161 (N_45161,N_44999,N_40476);
and U45162 (N_45162,N_44684,N_41761);
or U45163 (N_45163,N_40585,N_40173);
and U45164 (N_45164,N_40254,N_41726);
nor U45165 (N_45165,N_42298,N_41158);
and U45166 (N_45166,N_43921,N_43024);
xor U45167 (N_45167,N_40623,N_41884);
and U45168 (N_45168,N_44117,N_44310);
nor U45169 (N_45169,N_40439,N_42067);
or U45170 (N_45170,N_42331,N_43023);
nor U45171 (N_45171,N_44096,N_43192);
or U45172 (N_45172,N_40977,N_41023);
xnor U45173 (N_45173,N_43880,N_43476);
nor U45174 (N_45174,N_41685,N_43818);
nor U45175 (N_45175,N_42824,N_43578);
xor U45176 (N_45176,N_42619,N_41901);
nor U45177 (N_45177,N_41529,N_41394);
or U45178 (N_45178,N_42070,N_42456);
or U45179 (N_45179,N_44850,N_40635);
xnor U45180 (N_45180,N_40885,N_41556);
xor U45181 (N_45181,N_43698,N_44262);
and U45182 (N_45182,N_40230,N_44514);
xor U45183 (N_45183,N_43780,N_42610);
nand U45184 (N_45184,N_41089,N_41425);
nand U45185 (N_45185,N_44104,N_42337);
nor U45186 (N_45186,N_43408,N_42359);
and U45187 (N_45187,N_44659,N_42637);
nor U45188 (N_45188,N_40877,N_41772);
nor U45189 (N_45189,N_43866,N_43181);
nand U45190 (N_45190,N_40887,N_40918);
or U45191 (N_45191,N_42074,N_44392);
or U45192 (N_45192,N_43250,N_42825);
and U45193 (N_45193,N_41448,N_42144);
xor U45194 (N_45194,N_42235,N_42333);
xnor U45195 (N_45195,N_44740,N_40990);
or U45196 (N_45196,N_44566,N_42704);
or U45197 (N_45197,N_43554,N_42414);
nor U45198 (N_45198,N_43533,N_43585);
or U45199 (N_45199,N_41085,N_42415);
or U45200 (N_45200,N_41308,N_42141);
xor U45201 (N_45201,N_40572,N_41048);
nor U45202 (N_45202,N_40500,N_42163);
nand U45203 (N_45203,N_42111,N_42950);
nand U45204 (N_45204,N_44903,N_41109);
nor U45205 (N_45205,N_43934,N_41052);
xnor U45206 (N_45206,N_40523,N_41597);
and U45207 (N_45207,N_42403,N_41216);
and U45208 (N_45208,N_44115,N_40210);
nand U45209 (N_45209,N_41861,N_40111);
nand U45210 (N_45210,N_41115,N_43036);
xor U45211 (N_45211,N_42718,N_42968);
xnor U45212 (N_45212,N_44032,N_41372);
nand U45213 (N_45213,N_41870,N_40515);
and U45214 (N_45214,N_43691,N_44188);
nand U45215 (N_45215,N_42905,N_43247);
or U45216 (N_45216,N_43062,N_41994);
xnor U45217 (N_45217,N_44814,N_44686);
or U45218 (N_45218,N_42725,N_43178);
and U45219 (N_45219,N_41709,N_42170);
nand U45220 (N_45220,N_43183,N_41700);
or U45221 (N_45221,N_43073,N_42813);
and U45222 (N_45222,N_44407,N_42851);
nor U45223 (N_45223,N_44416,N_43371);
nor U45224 (N_45224,N_40353,N_43357);
nor U45225 (N_45225,N_40896,N_44916);
and U45226 (N_45226,N_40625,N_40616);
nand U45227 (N_45227,N_43886,N_41081);
xnor U45228 (N_45228,N_42938,N_42994);
or U45229 (N_45229,N_43695,N_42107);
nor U45230 (N_45230,N_43195,N_41928);
xnor U45231 (N_45231,N_43772,N_43383);
and U45232 (N_45232,N_43937,N_41389);
xor U45233 (N_45233,N_40622,N_42951);
and U45234 (N_45234,N_42155,N_43712);
and U45235 (N_45235,N_43262,N_42552);
and U45236 (N_45236,N_43365,N_43136);
nor U45237 (N_45237,N_41624,N_40637);
and U45238 (N_45238,N_40310,N_40876);
xor U45239 (N_45239,N_43984,N_40155);
nand U45240 (N_45240,N_44009,N_43083);
and U45241 (N_45241,N_40148,N_42339);
nor U45242 (N_45242,N_41850,N_42133);
or U45243 (N_45243,N_44856,N_44316);
or U45244 (N_45244,N_42374,N_40872);
and U45245 (N_45245,N_40780,N_44432);
xnor U45246 (N_45246,N_40846,N_41264);
or U45247 (N_45247,N_43707,N_40005);
and U45248 (N_45248,N_43474,N_42161);
xnor U45249 (N_45249,N_40880,N_40630);
and U45250 (N_45250,N_42097,N_44336);
xnor U45251 (N_45251,N_43304,N_43722);
or U45252 (N_45252,N_43467,N_41771);
and U45253 (N_45253,N_42551,N_42715);
or U45254 (N_45254,N_43123,N_44844);
nor U45255 (N_45255,N_43539,N_44891);
or U45256 (N_45256,N_43170,N_40289);
or U45257 (N_45257,N_44294,N_43422);
nor U45258 (N_45258,N_43610,N_42931);
and U45259 (N_45259,N_40970,N_42940);
or U45260 (N_45260,N_44733,N_41461);
xor U45261 (N_45261,N_40187,N_41661);
nand U45262 (N_45262,N_40215,N_42770);
nand U45263 (N_45263,N_43555,N_43078);
or U45264 (N_45264,N_41219,N_43961);
or U45265 (N_45265,N_41729,N_43413);
xnor U45266 (N_45266,N_41006,N_44638);
nand U45267 (N_45267,N_43473,N_43097);
xor U45268 (N_45268,N_40768,N_40399);
xor U45269 (N_45269,N_42591,N_43105);
nand U45270 (N_45270,N_40108,N_42381);
and U45271 (N_45271,N_44137,N_44256);
and U45272 (N_45272,N_44996,N_44642);
and U45273 (N_45273,N_41015,N_43574);
nor U45274 (N_45274,N_40307,N_41071);
and U45275 (N_45275,N_42231,N_41593);
and U45276 (N_45276,N_41469,N_40776);
xnor U45277 (N_45277,N_44986,N_41583);
xnor U45278 (N_45278,N_40450,N_41523);
and U45279 (N_45279,N_43661,N_40696);
nor U45280 (N_45280,N_42598,N_44691);
or U45281 (N_45281,N_44778,N_42280);
nor U45282 (N_45282,N_44350,N_41723);
or U45283 (N_45283,N_44650,N_44736);
or U45284 (N_45284,N_41534,N_43463);
xor U45285 (N_45285,N_41617,N_42405);
nor U45286 (N_45286,N_41183,N_43620);
and U45287 (N_45287,N_41801,N_44077);
xnor U45288 (N_45288,N_44656,N_44399);
nand U45289 (N_45289,N_43403,N_40529);
nand U45290 (N_45290,N_43602,N_42909);
or U45291 (N_45291,N_40950,N_42420);
xor U45292 (N_45292,N_41487,N_40916);
nor U45293 (N_45293,N_42354,N_42018);
xor U45294 (N_45294,N_43718,N_41165);
and U45295 (N_45295,N_42944,N_43863);
or U45296 (N_45296,N_44984,N_40649);
nand U45297 (N_45297,N_40502,N_44085);
nor U45298 (N_45298,N_44330,N_41311);
nor U45299 (N_45299,N_41470,N_40666);
nor U45300 (N_45300,N_40947,N_43957);
and U45301 (N_45301,N_44957,N_44357);
nand U45302 (N_45302,N_43177,N_44059);
nand U45303 (N_45303,N_40415,N_41547);
nand U45304 (N_45304,N_40946,N_42564);
and U45305 (N_45305,N_44567,N_41944);
xor U45306 (N_45306,N_40047,N_43966);
nor U45307 (N_45307,N_40789,N_41123);
or U45308 (N_45308,N_42808,N_44352);
nor U45309 (N_45309,N_41630,N_43828);
xor U45310 (N_45310,N_44526,N_43321);
nor U45311 (N_45311,N_41124,N_40737);
nor U45312 (N_45312,N_43905,N_43616);
and U45313 (N_45313,N_40482,N_44189);
or U45314 (N_45314,N_43580,N_44442);
and U45315 (N_45315,N_40778,N_42444);
or U45316 (N_45316,N_41882,N_44762);
or U45317 (N_45317,N_42793,N_42411);
or U45318 (N_45318,N_44221,N_40143);
and U45319 (N_45319,N_41472,N_43015);
and U45320 (N_45320,N_42627,N_44079);
nand U45321 (N_45321,N_43221,N_40160);
xnor U45322 (N_45322,N_44093,N_43857);
xor U45323 (N_45323,N_40553,N_44973);
or U45324 (N_45324,N_43793,N_44466);
xor U45325 (N_45325,N_41991,N_41580);
xnor U45326 (N_45326,N_44657,N_43225);
xnor U45327 (N_45327,N_42751,N_41409);
nor U45328 (N_45328,N_41266,N_40756);
nand U45329 (N_45329,N_43519,N_42407);
xor U45330 (N_45330,N_41888,N_40243);
or U45331 (N_45331,N_43945,N_44579);
nand U45332 (N_45332,N_41933,N_44014);
nor U45333 (N_45333,N_43672,N_43731);
nand U45334 (N_45334,N_40096,N_40362);
xor U45335 (N_45335,N_40985,N_43276);
nand U45336 (N_45336,N_41075,N_42678);
nor U45337 (N_45337,N_44562,N_41068);
nand U45338 (N_45338,N_42283,N_44155);
or U45339 (N_45339,N_43508,N_43597);
nand U45340 (N_45340,N_41776,N_41365);
nor U45341 (N_45341,N_43615,N_40464);
and U45342 (N_45342,N_42860,N_41635);
or U45343 (N_45343,N_42928,N_44868);
xor U45344 (N_45344,N_43488,N_42364);
or U45345 (N_45345,N_44478,N_42774);
nand U45346 (N_45346,N_41511,N_40280);
and U45347 (N_45347,N_40397,N_41539);
nor U45348 (N_45348,N_41516,N_41329);
or U45349 (N_45349,N_40146,N_43831);
and U45350 (N_45350,N_41682,N_44841);
xor U45351 (N_45351,N_42421,N_44730);
and U45352 (N_45352,N_42798,N_44196);
and U45353 (N_45353,N_42779,N_44569);
and U45354 (N_45354,N_42984,N_40767);
xor U45355 (N_45355,N_44931,N_43726);
nor U45356 (N_45356,N_43536,N_44696);
xor U45357 (N_45357,N_42220,N_40027);
nor U45358 (N_45358,N_40881,N_41164);
nor U45359 (N_45359,N_41209,N_41669);
or U45360 (N_45360,N_42504,N_42334);
nand U45361 (N_45361,N_44611,N_40820);
nand U45362 (N_45362,N_42497,N_44582);
xor U45363 (N_45363,N_43171,N_40853);
nand U45364 (N_45364,N_42912,N_42540);
xor U45365 (N_45365,N_44285,N_40021);
nand U45366 (N_45366,N_44929,N_40483);
nor U45367 (N_45367,N_42939,N_44813);
or U45368 (N_45368,N_44265,N_41891);
nand U45369 (N_45369,N_44333,N_41681);
nor U45370 (N_45370,N_43281,N_40433);
nand U45371 (N_45371,N_40949,N_43667);
xor U45372 (N_45372,N_43338,N_40290);
nor U45373 (N_45373,N_41375,N_43323);
nor U45374 (N_45374,N_44449,N_43058);
nor U45375 (N_45375,N_43736,N_41855);
or U45376 (N_45376,N_41633,N_41887);
or U45377 (N_45377,N_42109,N_43889);
nor U45378 (N_45378,N_42040,N_43636);
xor U45379 (N_45379,N_41005,N_44492);
and U45380 (N_45380,N_44967,N_41473);
or U45381 (N_45381,N_42043,N_42703);
or U45382 (N_45382,N_44018,N_43920);
nor U45383 (N_45383,N_43457,N_42963);
or U45384 (N_45384,N_44677,N_41293);
or U45385 (N_45385,N_40029,N_44893);
nor U45386 (N_45386,N_44643,N_42446);
xnor U45387 (N_45387,N_44128,N_40061);
and U45388 (N_45388,N_44818,N_43758);
nand U45389 (N_45389,N_44321,N_43071);
nor U45390 (N_45390,N_43638,N_41555);
or U45391 (N_45391,N_41922,N_43743);
xnor U45392 (N_45392,N_44063,N_43201);
or U45393 (N_45393,N_40497,N_42904);
nor U45394 (N_45394,N_43019,N_43750);
nand U45395 (N_45395,N_41274,N_43759);
nand U45396 (N_45396,N_43535,N_41820);
xor U45397 (N_45397,N_42884,N_40177);
and U45398 (N_45398,N_44319,N_43571);
or U45399 (N_45399,N_42643,N_42889);
nand U45400 (N_45400,N_41309,N_41481);
nor U45401 (N_45401,N_41476,N_44879);
nor U45402 (N_45402,N_42676,N_40810);
xnor U45403 (N_45403,N_44726,N_44950);
xnor U45404 (N_45404,N_43941,N_41995);
or U45405 (N_45405,N_41520,N_44683);
or U45406 (N_45406,N_44325,N_44535);
nand U45407 (N_45407,N_42122,N_41356);
or U45408 (N_45408,N_44051,N_44109);
or U45409 (N_45409,N_42819,N_40323);
and U45410 (N_45410,N_41376,N_41854);
or U45411 (N_45411,N_44555,N_43767);
nor U45412 (N_45412,N_40418,N_43595);
nor U45413 (N_45413,N_40627,N_40647);
or U45414 (N_45414,N_41727,N_44045);
nor U45415 (N_45415,N_43755,N_42069);
nand U45416 (N_45416,N_40982,N_43784);
nand U45417 (N_45417,N_42172,N_43121);
nand U45418 (N_45418,N_41639,N_44193);
xor U45419 (N_45419,N_42936,N_40834);
nor U45420 (N_45420,N_40890,N_44054);
and U45421 (N_45421,N_42186,N_42661);
nand U45422 (N_45422,N_42869,N_41782);
nand U45423 (N_45423,N_43982,N_43607);
and U45424 (N_45424,N_40368,N_43272);
or U45425 (N_45425,N_43047,N_44720);
or U45426 (N_45426,N_40527,N_40869);
or U45427 (N_45427,N_40691,N_40829);
or U45428 (N_45428,N_43319,N_42631);
nor U45429 (N_45429,N_44075,N_43909);
nand U45430 (N_45430,N_44528,N_40349);
or U45431 (N_45431,N_40840,N_40717);
or U45432 (N_45432,N_43378,N_41571);
nor U45433 (N_45433,N_43987,N_44923);
or U45434 (N_45434,N_42972,N_40463);
nor U45435 (N_45435,N_40679,N_42677);
nand U45436 (N_45436,N_42802,N_41252);
xor U45437 (N_45437,N_41514,N_40965);
and U45438 (N_45438,N_41077,N_42867);
nor U45439 (N_45439,N_41692,N_42815);
xor U45440 (N_45440,N_42449,N_44329);
nand U45441 (N_45441,N_41728,N_43512);
nor U45442 (N_45442,N_42692,N_40413);
nor U45443 (N_45443,N_42579,N_44775);
or U45444 (N_45444,N_43452,N_42686);
and U45445 (N_45445,N_43693,N_40076);
and U45446 (N_45446,N_44175,N_40870);
or U45447 (N_45447,N_41544,N_40602);
nand U45448 (N_45448,N_41125,N_41413);
or U45449 (N_45449,N_44172,N_44920);
or U45450 (N_45450,N_41318,N_42893);
nand U45451 (N_45451,N_44364,N_42136);
xnor U45452 (N_45452,N_43377,N_41284);
and U45453 (N_45453,N_42666,N_40457);
xor U45454 (N_45454,N_40424,N_44822);
or U45455 (N_45455,N_41024,N_43783);
nand U45456 (N_45456,N_44639,N_41838);
xor U45457 (N_45457,N_40882,N_44181);
or U45458 (N_45458,N_40090,N_41238);
nand U45459 (N_45459,N_44224,N_44064);
nor U45460 (N_45460,N_44171,N_40892);
or U45461 (N_45461,N_41208,N_44545);
and U45462 (N_45462,N_42370,N_40967);
or U45463 (N_45463,N_42521,N_40403);
nor U45464 (N_45464,N_43350,N_42473);
nor U45465 (N_45465,N_43199,N_42247);
and U45466 (N_45466,N_42031,N_40849);
nand U45467 (N_45467,N_43407,N_43082);
or U45468 (N_45468,N_43910,N_40038);
xnor U45469 (N_45469,N_41103,N_42982);
xnor U45470 (N_45470,N_41152,N_41032);
nand U45471 (N_45471,N_40569,N_41184);
xnor U45472 (N_45472,N_44888,N_43263);
nand U45473 (N_45473,N_44785,N_43665);
and U45474 (N_45474,N_40964,N_41401);
nand U45475 (N_45475,N_43115,N_42395);
and U45476 (N_45476,N_41065,N_43127);
nor U45477 (N_45477,N_42638,N_42844);
nand U45478 (N_45478,N_42655,N_44043);
xor U45479 (N_45479,N_43846,N_44264);
and U45480 (N_45480,N_42303,N_41025);
nand U45481 (N_45481,N_42702,N_42367);
xnor U45482 (N_45482,N_44112,N_41173);
and U45483 (N_45483,N_44886,N_42020);
nand U45484 (N_45484,N_42533,N_43771);
and U45485 (N_45485,N_41362,N_41805);
xor U45486 (N_45486,N_44266,N_42828);
or U45487 (N_45487,N_44501,N_43441);
nand U45488 (N_45488,N_42149,N_43625);
nand U45489 (N_45489,N_44989,N_40188);
or U45490 (N_45490,N_43617,N_44118);
xor U45491 (N_45491,N_42262,N_42014);
or U45492 (N_45492,N_44490,N_43404);
xor U45493 (N_45493,N_44147,N_43447);
nor U45494 (N_45494,N_41892,N_43477);
nand U45495 (N_45495,N_44421,N_43798);
xnor U45496 (N_45496,N_41591,N_42123);
nand U45497 (N_45497,N_42320,N_44606);
nand U45498 (N_45498,N_44025,N_41438);
xnor U45499 (N_45499,N_42611,N_41918);
and U45500 (N_45500,N_43343,N_40514);
and U45501 (N_45501,N_41146,N_42087);
xor U45502 (N_45502,N_40822,N_43194);
and U45503 (N_45503,N_43762,N_41910);
xnor U45504 (N_45504,N_41257,N_42903);
xnor U45505 (N_45505,N_42487,N_40779);
xor U45506 (N_45506,N_43290,N_44202);
nand U45507 (N_45507,N_42875,N_40884);
xnor U45508 (N_45508,N_42746,N_41450);
nor U45509 (N_45509,N_41588,N_43933);
nor U45510 (N_45510,N_42625,N_42921);
xor U45511 (N_45511,N_44324,N_42958);
xnor U45512 (N_45512,N_44896,N_41715);
or U45513 (N_45513,N_44998,N_44295);
nor U45514 (N_45514,N_40231,N_41136);
nand U45515 (N_45515,N_41637,N_43837);
nor U45516 (N_45516,N_43236,N_40879);
or U45517 (N_45517,N_42915,N_43384);
xor U45518 (N_45518,N_41133,N_41354);
nor U45519 (N_45519,N_40419,N_40494);
nor U45520 (N_45520,N_42577,N_43315);
nand U45521 (N_45521,N_44612,N_44159);
or U45522 (N_45522,N_41875,N_42690);
nand U45523 (N_45523,N_44645,N_42817);
nand U45524 (N_45524,N_41105,N_42171);
nor U45525 (N_45525,N_43745,N_43336);
nand U45526 (N_45526,N_44792,N_40499);
nand U45527 (N_45527,N_43425,N_44486);
xor U45528 (N_45528,N_41116,N_40377);
nand U45529 (N_45529,N_40980,N_41768);
xnor U45530 (N_45530,N_44382,N_41708);
nand U45531 (N_45531,N_43552,N_43705);
nor U45532 (N_45532,N_40645,N_43458);
xor U45533 (N_45533,N_43618,N_42539);
or U45534 (N_45534,N_40122,N_40831);
and U45535 (N_45535,N_42046,N_44919);
nor U45536 (N_45536,N_41047,N_44668);
or U45537 (N_45537,N_41960,N_41939);
nand U45538 (N_45538,N_43017,N_43327);
nor U45539 (N_45539,N_41169,N_42233);
nand U45540 (N_45540,N_41587,N_41652);
and U45541 (N_45541,N_43306,N_43753);
or U45542 (N_45542,N_43232,N_44828);
nor U45543 (N_45543,N_43868,N_43946);
nand U45544 (N_45544,N_42358,N_43411);
xor U45545 (N_45545,N_43174,N_41364);
nand U45546 (N_45546,N_43680,N_44446);
or U45547 (N_45547,N_43094,N_40815);
nand U45548 (N_45548,N_41783,N_40342);
or U45549 (N_45549,N_42312,N_43902);
xnor U45550 (N_45550,N_41082,N_44010);
or U45551 (N_45551,N_40923,N_42723);
nand U45552 (N_45552,N_44679,N_42532);
and U45553 (N_45553,N_42763,N_42326);
and U45554 (N_45554,N_40086,N_43563);
xnor U45555 (N_45555,N_42134,N_42064);
and U45556 (N_45556,N_43862,N_43802);
xnor U45557 (N_45557,N_44626,N_44049);
nand U45558 (N_45558,N_41959,N_42084);
nor U45559 (N_45559,N_43288,N_43165);
nor U45560 (N_45560,N_40491,N_44764);
nand U45561 (N_45561,N_43175,N_42534);
xor U45562 (N_45562,N_41878,N_44124);
or U45563 (N_45563,N_43216,N_44050);
or U45564 (N_45564,N_40065,N_40522);
and U45565 (N_45565,N_42392,N_43844);
nand U45566 (N_45566,N_41346,N_41625);
xnor U45567 (N_45567,N_42448,N_42582);
or U45568 (N_45568,N_42041,N_43522);
or U45569 (N_45569,N_40784,N_41104);
xor U45570 (N_45570,N_44680,N_40095);
nand U45571 (N_45571,N_44816,N_43806);
or U45572 (N_45572,N_41283,N_41390);
xor U45573 (N_45573,N_40898,N_41695);
or U45574 (N_45574,N_41607,N_44274);
nor U45575 (N_45575,N_40244,N_44937);
or U45576 (N_45576,N_40018,N_42783);
nand U45577 (N_45577,N_42167,N_41460);
nand U45578 (N_45578,N_44634,N_41097);
and U45579 (N_45579,N_44769,N_40013);
nand U45580 (N_45580,N_40862,N_43710);
nand U45581 (N_45581,N_42300,N_41494);
nor U45582 (N_45582,N_42091,N_41810);
xnor U45583 (N_45583,N_43820,N_42659);
nand U45584 (N_45584,N_40531,N_44284);
nand U45585 (N_45585,N_40678,N_43335);
nand U45586 (N_45586,N_43503,N_41760);
and U45587 (N_45587,N_40919,N_40994);
and U45588 (N_45588,N_41812,N_41620);
xnor U45589 (N_45589,N_41902,N_44902);
nor U45590 (N_45590,N_44729,N_43593);
and U45591 (N_45591,N_43674,N_44773);
or U45592 (N_45592,N_43347,N_42471);
or U45593 (N_45593,N_42797,N_44445);
xnor U45594 (N_45594,N_40628,N_42035);
and U45595 (N_45595,N_41112,N_42218);
nor U45596 (N_45596,N_41355,N_40278);
nand U45597 (N_45597,N_41900,N_44586);
nor U45598 (N_45598,N_44098,N_42455);
and U45599 (N_45599,N_40997,N_43805);
xor U45600 (N_45600,N_43151,N_42775);
and U45601 (N_45601,N_43879,N_42507);
xor U45602 (N_45602,N_40566,N_40246);
nor U45603 (N_45603,N_43790,N_40655);
xor U45604 (N_45604,N_42732,N_42836);
nand U45605 (N_45605,N_42036,N_41860);
and U45606 (N_45606,N_42485,N_42311);
xnor U45607 (N_45607,N_42265,N_42174);
and U45608 (N_45608,N_44301,N_44621);
nor U45609 (N_45609,N_41176,N_44737);
or U45610 (N_45610,N_44065,N_42826);
and U45611 (N_45611,N_44798,N_41061);
or U45612 (N_45612,N_44186,N_41862);
or U45613 (N_45613,N_44056,N_43715);
nand U45614 (N_45614,N_42618,N_43436);
or U45615 (N_45615,N_43230,N_42841);
or U45616 (N_45616,N_41358,N_41130);
or U45617 (N_45617,N_40772,N_42325);
and U45618 (N_45618,N_40447,N_41612);
xor U45619 (N_45619,N_42656,N_40611);
and U45620 (N_45620,N_41106,N_41911);
nand U45621 (N_45621,N_41977,N_40408);
nor U45622 (N_45622,N_41432,N_42308);
nor U45623 (N_45623,N_40312,N_43479);
and U45624 (N_45624,N_40719,N_43764);
or U45625 (N_45625,N_41707,N_42740);
and U45626 (N_45626,N_43605,N_44123);
xor U45627 (N_45627,N_40448,N_42773);
and U45628 (N_45628,N_44543,N_42697);
or U45629 (N_45629,N_41192,N_40367);
xor U45630 (N_45630,N_43683,N_42322);
nand U45631 (N_45631,N_44722,N_43316);
xnor U45632 (N_45632,N_44460,N_43011);
and U45633 (N_45633,N_42263,N_42304);
nand U45634 (N_45634,N_42648,N_44685);
xor U45635 (N_45635,N_40348,N_40875);
or U45636 (N_45636,N_42918,N_41066);
and U45637 (N_45637,N_43243,N_40178);
or U45638 (N_45638,N_43911,N_44309);
or U45639 (N_45639,N_42886,N_42424);
nor U45640 (N_45640,N_43841,N_43079);
nand U45641 (N_45641,N_43046,N_41965);
or U45642 (N_45642,N_42106,N_43007);
nor U45643 (N_45643,N_44819,N_41644);
nand U45644 (N_45644,N_40978,N_44883);
nand U45645 (N_45645,N_42645,N_42741);
xnor U45646 (N_45646,N_40401,N_43424);
nand U45647 (N_45647,N_42556,N_41144);
xnor U45648 (N_45648,N_43003,N_42809);
or U45649 (N_45649,N_42193,N_44156);
nor U45650 (N_45650,N_42042,N_41162);
and U45651 (N_45651,N_42285,N_44461);
nand U45652 (N_45652,N_40986,N_40817);
or U45653 (N_45653,N_42396,N_42512);
xor U45654 (N_45654,N_43103,N_41636);
and U45655 (N_45655,N_42660,N_43777);
nor U45656 (N_45656,N_44036,N_44267);
or U45657 (N_45657,N_42518,N_43013);
nand U45658 (N_45658,N_44431,N_42249);
xnor U45659 (N_45659,N_40864,N_43590);
or U45660 (N_45660,N_41987,N_43794);
and U45661 (N_45661,N_44662,N_40436);
nand U45662 (N_45662,N_44546,N_44724);
nor U45663 (N_45663,N_44561,N_44949);
xnor U45664 (N_45664,N_40031,N_44088);
and U45665 (N_45665,N_43624,N_41828);
xor U45666 (N_45666,N_42513,N_43543);
nand U45667 (N_45667,N_44279,N_44342);
xnor U45668 (N_45668,N_42906,N_40886);
xnor U45669 (N_45669,N_43313,N_42350);
and U45670 (N_45670,N_43830,N_44004);
and U45671 (N_45671,N_44616,N_40402);
xor U45672 (N_45672,N_42199,N_44959);
nor U45673 (N_45673,N_40993,N_43270);
nor U45674 (N_45674,N_43730,N_42017);
or U45675 (N_45675,N_41369,N_42412);
xor U45676 (N_45676,N_42256,N_44347);
and U45677 (N_45677,N_43485,N_41297);
nand U45678 (N_45678,N_40049,N_40676);
and U45679 (N_45679,N_43768,N_44055);
or U45680 (N_45680,N_40059,N_41378);
xnor U45681 (N_45681,N_41087,N_42609);
xor U45682 (N_45682,N_44020,N_44375);
and U45683 (N_45683,N_42529,N_41452);
and U45684 (N_45684,N_43329,N_44272);
and U45685 (N_45685,N_40709,N_41203);
or U45686 (N_45686,N_41733,N_42795);
and U45687 (N_45687,N_44952,N_42191);
nand U45688 (N_45688,N_44714,N_44801);
nand U45689 (N_45689,N_41485,N_42182);
nor U45690 (N_45690,N_41975,N_44557);
and U45691 (N_45691,N_43967,N_40331);
nor U45692 (N_45692,N_44103,N_44201);
xor U45693 (N_45693,N_41576,N_43648);
and U45694 (N_45694,N_42187,N_40109);
or U45695 (N_45695,N_43807,N_43733);
and U45696 (N_45696,N_44302,N_41629);
nor U45697 (N_45697,N_41777,N_44857);
and U45698 (N_45698,N_40934,N_43302);
or U45699 (N_45699,N_43386,N_42130);
and U45700 (N_45700,N_40078,N_42417);
xor U45701 (N_45701,N_40609,N_40601);
or U45702 (N_45702,N_41499,N_44212);
or U45703 (N_45703,N_42491,N_43913);
nor U45704 (N_45704,N_43445,N_42620);
and U45705 (N_45705,N_43697,N_44651);
nand U45706 (N_45706,N_43095,N_43619);
xor U45707 (N_45707,N_42833,N_41043);
and U45708 (N_45708,N_44983,N_43871);
xnor U45709 (N_45709,N_44971,N_42954);
xor U45710 (N_45710,N_41058,N_44608);
or U45711 (N_45711,N_42297,N_44870);
nor U45712 (N_45712,N_44244,N_40443);
or U45713 (N_45713,N_40124,N_44248);
or U45714 (N_45714,N_40009,N_41525);
or U45715 (N_45715,N_41483,N_42830);
nor U45716 (N_45716,N_44593,N_42110);
nand U45717 (N_45717,N_41645,N_41254);
nor U45718 (N_45718,N_44675,N_40034);
nand U45719 (N_45719,N_43781,N_41656);
and U45720 (N_45720,N_40237,N_40462);
nor U45721 (N_45721,N_42624,N_41224);
or U45722 (N_45722,N_42183,N_43813);
nor U45723 (N_45723,N_40101,N_43341);
xnor U45724 (N_45724,N_44068,N_43207);
xor U45725 (N_45725,N_41200,N_40167);
nor U45726 (N_45726,N_41790,N_44556);
or U45727 (N_45727,N_43145,N_41028);
xor U45728 (N_45728,N_42397,N_40658);
xnor U45729 (N_45729,N_42037,N_43246);
nand U45730 (N_45730,N_40579,N_40972);
nor U45731 (N_45731,N_43654,N_40513);
xnor U45732 (N_45732,N_41102,N_41763);
and U45733 (N_45733,N_43581,N_40675);
or U45734 (N_45734,N_40674,N_41148);
and U45735 (N_45735,N_41170,N_40684);
and U45736 (N_45736,N_41962,N_40070);
xnor U45737 (N_45737,N_41823,N_42398);
xor U45738 (N_45738,N_41559,N_44618);
and U45739 (N_45739,N_43352,N_42158);
nand U45740 (N_45740,N_43222,N_40521);
nand U45741 (N_45741,N_41793,N_43356);
or U45742 (N_45742,N_42789,N_40981);
xnor U45743 (N_45743,N_40088,N_44078);
nand U45744 (N_45744,N_43873,N_44367);
xor U45745 (N_45745,N_41013,N_43051);
nand U45746 (N_45746,N_42438,N_42098);
nand U45747 (N_45747,N_41134,N_40412);
nor U45748 (N_45748,N_41055,N_42747);
nand U45749 (N_45749,N_41604,N_44653);
or U45750 (N_45750,N_41521,N_40176);
nand U45751 (N_45751,N_44779,N_42463);
xor U45752 (N_45752,N_41440,N_43054);
nor U45753 (N_45753,N_43675,N_40548);
xor U45754 (N_45754,N_41424,N_41477);
and U45755 (N_45755,N_43196,N_42034);
or U45756 (N_45756,N_44110,N_44303);
and U45757 (N_45757,N_42148,N_42727);
and U45758 (N_45758,N_42131,N_42689);
xnor U45759 (N_45759,N_40075,N_41292);
or U45760 (N_45760,N_41541,N_40438);
xor U45761 (N_45761,N_43634,N_42927);
nor U45762 (N_45762,N_40156,N_42243);
or U45763 (N_45763,N_40329,N_43184);
nor U45764 (N_45764,N_43072,N_41923);
and U45765 (N_45765,N_41359,N_43342);
nor U45766 (N_45766,N_41475,N_41937);
xor U45767 (N_45767,N_42899,N_42022);
nor U45768 (N_45768,N_44158,N_40827);
nor U45769 (N_45769,N_40264,N_43464);
xor U45770 (N_45770,N_42188,N_41608);
and U45771 (N_45771,N_40098,N_43048);
xor U45772 (N_45772,N_44796,N_40056);
nand U45773 (N_45773,N_41551,N_43415);
or U45774 (N_45774,N_41259,N_43213);
nor U45775 (N_45775,N_42301,N_42855);
or U45776 (N_45776,N_44213,N_40325);
or U45777 (N_45777,N_44559,N_42500);
nand U45778 (N_45778,N_42739,N_41147);
xnor U45779 (N_45779,N_43594,N_41301);
xor U45780 (N_45780,N_41039,N_44988);
or U45781 (N_45781,N_40479,N_44150);
nand U45782 (N_45782,N_41531,N_43260);
or U45783 (N_45783,N_42399,N_44426);
nor U45784 (N_45784,N_42542,N_42484);
xor U45785 (N_45785,N_43851,N_44019);
or U45786 (N_45786,N_43685,N_41280);
nand U45787 (N_45787,N_40945,N_44922);
and U45788 (N_45788,N_42644,N_42390);
nand U45789 (N_45789,N_42088,N_40055);
xnor U45790 (N_45790,N_44908,N_44881);
and U45791 (N_45791,N_40301,N_43291);
or U45792 (N_45792,N_42596,N_44312);
or U45793 (N_45793,N_44397,N_44795);
xor U45794 (N_45794,N_43681,N_40240);
and U45795 (N_45795,N_43486,N_43139);
and U45796 (N_45796,N_43421,N_41779);
or U45797 (N_45797,N_42910,N_43002);
or U45798 (N_45798,N_44195,N_42437);
nor U45799 (N_45799,N_42987,N_41310);
nand U45800 (N_45800,N_41969,N_42089);
and U45801 (N_45801,N_43298,N_40927);
xor U45802 (N_45802,N_41557,N_44283);
and U45803 (N_45803,N_40754,N_41654);
xor U45804 (N_45804,N_41275,N_42967);
nand U45805 (N_45805,N_41294,N_41827);
or U45806 (N_45806,N_44260,N_42733);
and U45807 (N_45807,N_40119,N_41212);
nand U45808 (N_45808,N_44905,N_42356);
or U45809 (N_45809,N_43975,N_40942);
and U45810 (N_45810,N_40409,N_44425);
nor U45811 (N_45811,N_43500,N_41874);
or U45812 (N_45812,N_40341,N_40261);
or U45813 (N_45813,N_40066,N_44784);
or U45814 (N_45814,N_43405,N_43545);
and U45815 (N_45815,N_43435,N_42948);
nand U45816 (N_45816,N_44146,N_42784);
or U45817 (N_45817,N_43754,N_43387);
and U45818 (N_45818,N_43514,N_40456);
xor U45819 (N_45819,N_44275,N_40216);
and U45820 (N_45820,N_42215,N_43076);
and U45821 (N_45821,N_42606,N_44519);
nor U45822 (N_45822,N_41712,N_40791);
nand U45823 (N_45823,N_43525,N_43576);
and U45824 (N_45824,N_40706,N_44829);
xor U45825 (N_45825,N_41377,N_44331);
nor U45826 (N_45826,N_42766,N_44995);
xnor U45827 (N_45827,N_43676,N_41398);
nor U45828 (N_45828,N_43430,N_44026);
xor U45829 (N_45829,N_41766,N_42251);
or U45830 (N_45830,N_43475,N_43114);
nand U45831 (N_45831,N_43694,N_40828);
xor U45832 (N_45832,N_41495,N_43493);
and U45833 (N_45833,N_41851,N_44126);
and U45834 (N_45834,N_40437,N_44754);
nor U45835 (N_45835,N_44900,N_43655);
xor U45836 (N_45836,N_40902,N_40123);
nor U45837 (N_45837,N_44571,N_43312);
or U45838 (N_45838,N_44947,N_41373);
and U45839 (N_45839,N_44390,N_42472);
xnor U45840 (N_45840,N_41713,N_41554);
or U45841 (N_45841,N_41228,N_42388);
nor U45842 (N_45842,N_40247,N_44405);
nor U45843 (N_45843,N_40998,N_44057);
or U45844 (N_45844,N_43117,N_41459);
and U45845 (N_45845,N_42630,N_40039);
or U45846 (N_45846,N_40306,N_44777);
and U45847 (N_45847,N_43397,N_41665);
nor U45848 (N_45848,N_40384,N_42428);
nor U45849 (N_45849,N_40851,N_40901);
nor U45850 (N_45850,N_42641,N_42827);
nor U45851 (N_45851,N_40894,N_42765);
xnor U45852 (N_45852,N_42016,N_41848);
or U45853 (N_45853,N_41434,N_44437);
nand U45854 (N_45854,N_42688,N_41135);
xnor U45855 (N_45855,N_40449,N_40608);
and U45856 (N_45856,N_40542,N_44763);
nand U45857 (N_45857,N_42468,N_44005);
or U45858 (N_45858,N_42962,N_42621);
or U45859 (N_45859,N_41721,N_43030);
nor U45860 (N_45860,N_44505,N_43284);
nand U45861 (N_45861,N_41972,N_42947);
nor U45862 (N_45862,N_40343,N_41175);
and U45863 (N_45863,N_43041,N_43652);
nand U45864 (N_45864,N_40895,N_42663);
nor U45865 (N_45865,N_42672,N_41041);
and U45866 (N_45866,N_40337,N_44024);
nand U45867 (N_45867,N_43231,N_44204);
nand U45868 (N_45868,N_41754,N_42885);
nand U45869 (N_45869,N_41099,N_40369);
xor U45870 (N_45870,N_41016,N_43922);
nor U45871 (N_45871,N_42707,N_42082);
and U45872 (N_45872,N_41676,N_41150);
nor U45873 (N_45873,N_41683,N_40432);
or U45874 (N_45874,N_43240,N_43042);
and U45875 (N_45875,N_40378,N_43116);
xor U45876 (N_45876,N_42053,N_43627);
or U45877 (N_45877,N_41879,N_43267);
nand U45878 (N_45878,N_40712,N_44719);
and U45879 (N_45879,N_43138,N_44832);
xor U45880 (N_45880,N_40186,N_43557);
and U45881 (N_45881,N_43622,N_40001);
or U45882 (N_45882,N_44360,N_43656);
and U45883 (N_45883,N_44231,N_42615);
nor U45884 (N_45884,N_41716,N_42864);
nor U45885 (N_45885,N_40465,N_40252);
xor U45886 (N_45886,N_40407,N_41009);
or U45887 (N_45887,N_43916,N_40166);
nand U45888 (N_45888,N_40366,N_40988);
nor U45889 (N_45889,N_43609,N_44839);
or U45890 (N_45890,N_44749,N_42208);
nor U45891 (N_45891,N_44847,N_41631);
nand U45892 (N_45892,N_40202,N_40619);
xor U45893 (N_45893,N_43701,N_44892);
and U45894 (N_45894,N_43163,N_43269);
nor U45895 (N_45895,N_42811,N_43487);
and U45896 (N_45896,N_40273,N_40295);
nor U45897 (N_45897,N_41904,N_42699);
xor U45898 (N_45898,N_40161,N_41331);
xnor U45899 (N_45899,N_44094,N_43739);
and U45900 (N_45900,N_44344,N_41569);
xor U45901 (N_45901,N_41664,N_42294);
and U45902 (N_45902,N_41549,N_41229);
or U45903 (N_45903,N_42492,N_41968);
nand U45904 (N_45904,N_44958,N_42015);
nor U45905 (N_45905,N_43811,N_43349);
nand U45906 (N_45906,N_40888,N_40257);
xnor U45907 (N_45907,N_42681,N_42983);
and U45908 (N_45908,N_42995,N_42476);
and U45909 (N_45909,N_41287,N_42440);
and U45910 (N_45910,N_41451,N_43962);
xor U45911 (N_45911,N_41423,N_42470);
nand U45912 (N_45912,N_40414,N_44371);
or U45913 (N_45913,N_40236,N_44578);
xnor U45914 (N_45914,N_42458,N_44921);
nand U45915 (N_45915,N_41641,N_43090);
xnor U45916 (N_45916,N_40434,N_40928);
nor U45917 (N_45917,N_44910,N_40267);
xor U45918 (N_45918,N_41386,N_42709);
nand U45919 (N_45919,N_43822,N_43583);
or U45920 (N_45920,N_43690,N_44060);
and U45921 (N_45921,N_41205,N_41935);
nor U45922 (N_45922,N_40040,N_43204);
xnor U45923 (N_45923,N_40125,N_44956);
xnor U45924 (N_45924,N_40961,N_41675);
and U45925 (N_45925,N_44356,N_42990);
xor U45926 (N_45926,N_41600,N_44865);
or U45927 (N_45927,N_44452,N_41127);
or U45928 (N_45928,N_44817,N_40092);
or U45929 (N_45929,N_43198,N_43156);
and U45930 (N_45930,N_42778,N_41101);
or U45931 (N_45931,N_40550,N_41575);
xnor U45932 (N_45932,N_40175,N_40140);
xnor U45933 (N_45933,N_41367,N_40480);
xor U45934 (N_45934,N_44121,N_44809);
nor U45935 (N_45935,N_40984,N_41739);
nand U45936 (N_45936,N_41755,N_43621);
nor U45937 (N_45937,N_42157,N_43208);
and U45938 (N_45938,N_40516,N_40245);
xor U45939 (N_45939,N_40372,N_43568);
nand U45940 (N_45940,N_40485,N_40493);
nor U45941 (N_45941,N_41429,N_40002);
and U45942 (N_45942,N_40258,N_44235);
xor U45943 (N_45943,N_40910,N_40577);
nand U45944 (N_45944,N_43993,N_43663);
nand U45945 (N_45945,N_44338,N_44339);
nand U45946 (N_45946,N_42969,N_42971);
and U45947 (N_45947,N_44187,N_41328);
nor U45948 (N_45948,N_40596,N_40748);
nor U45949 (N_45949,N_43285,N_41223);
and U45950 (N_45950,N_43577,N_43044);
nand U45951 (N_45951,N_40734,N_42101);
nand U45952 (N_45952,N_44022,N_40790);
and U45953 (N_45953,N_44884,N_41711);
or U45954 (N_45954,N_40459,N_44824);
and U45955 (N_45955,N_42095,N_43040);
and U45956 (N_45956,N_42999,N_43645);
nor U45957 (N_45957,N_41412,N_44499);
xor U45958 (N_45958,N_42759,N_42464);
nor U45959 (N_45959,N_40241,N_42006);
and U45960 (N_45960,N_44439,N_44002);
nand U45961 (N_45961,N_40142,N_41063);
nand U45962 (N_45962,N_44738,N_43840);
or U45963 (N_45963,N_42344,N_40996);
or U45964 (N_45964,N_41191,N_43708);
or U45965 (N_45965,N_43935,N_42068);
or U45966 (N_45966,N_43586,N_40340);
nor U45967 (N_45967,N_43340,N_44468);
xnor U45968 (N_45968,N_42714,N_42557);
nand U45969 (N_45969,N_40162,N_42584);
nor U45970 (N_45970,N_40181,N_44182);
nand U45971 (N_45971,N_43037,N_44909);
or U45972 (N_45972,N_40503,N_41273);
nor U45973 (N_45973,N_43289,N_40586);
and U45974 (N_45974,N_42519,N_44767);
nand U45975 (N_45975,N_41478,N_41794);
or U45976 (N_45976,N_44658,N_43122);
xor U45977 (N_45977,N_40564,N_40583);
or U45978 (N_45978,N_43410,N_44508);
nor U45979 (N_45979,N_42180,N_44935);
or U45980 (N_45980,N_44768,N_43389);
and U45981 (N_45981,N_42207,N_40387);
nor U45982 (N_45982,N_41674,N_43598);
nor U45983 (N_45983,N_42252,N_44928);
xor U45984 (N_45984,N_41693,N_41258);
xor U45985 (N_45985,N_42974,N_42916);
nor U45986 (N_45986,N_42616,N_43426);
xor U45987 (N_45987,N_43834,N_44966);
nor U45988 (N_45988,N_41366,N_42576);
and U45989 (N_45989,N_44239,N_44372);
or U45990 (N_45990,N_40963,N_43747);
nor U45991 (N_45991,N_43110,N_43877);
or U45992 (N_45992,N_44924,N_41889);
nor U45993 (N_45993,N_42156,N_44273);
xnor U45994 (N_45994,N_40660,N_40426);
and U45995 (N_45995,N_41090,N_41022);
xnor U45996 (N_45996,N_42907,N_40116);
nor U45997 (N_45997,N_44450,N_41662);
nor U45998 (N_45998,N_41912,N_41804);
and U45999 (N_45999,N_43244,N_42874);
nor U46000 (N_46000,N_43469,N_41323);
or U46001 (N_46001,N_41315,N_40471);
or U46002 (N_46002,N_43432,N_43490);
or U46003 (N_46003,N_40613,N_40782);
nand U46004 (N_46004,N_40201,N_40841);
xnor U46005 (N_46005,N_44756,N_44747);
nand U46006 (N_46006,N_43000,N_43434);
nor U46007 (N_46007,N_41214,N_43004);
xor U46008 (N_46008,N_44620,N_42804);
or U46009 (N_46009,N_40868,N_40104);
nor U46010 (N_46010,N_42961,N_42562);
and U46011 (N_46011,N_42175,N_42195);
and U46012 (N_46012,N_43257,N_43632);
nor U46013 (N_46013,N_42425,N_44759);
xnor U46014 (N_46014,N_40073,N_43107);
xor U46015 (N_46015,N_40711,N_41508);
nor U46016 (N_46016,N_41268,N_40195);
nor U46017 (N_46017,N_43358,N_43368);
and U46018 (N_46018,N_43200,N_44046);
or U46019 (N_46019,N_43553,N_40466);
xnor U46020 (N_46020,N_41579,N_44134);
or U46021 (N_46021,N_42386,N_40939);
and U46022 (N_46022,N_42531,N_40327);
nor U46023 (N_46023,N_41824,N_44532);
nand U46024 (N_46024,N_43451,N_42801);
nand U46025 (N_46025,N_40727,N_44378);
nor U46026 (N_46026,N_40180,N_40147);
nor U46027 (N_46027,N_41552,N_42602);
and U46028 (N_46028,N_40496,N_40788);
and U46029 (N_46029,N_44934,N_43020);
nand U46030 (N_46030,N_41789,N_42650);
nand U46031 (N_46031,N_43006,N_44307);
and U46032 (N_46032,N_44534,N_44974);
and U46033 (N_46033,N_44793,N_41237);
nor U46034 (N_46034,N_40509,N_40232);
and U46035 (N_46035,N_41069,N_40960);
nand U46036 (N_46036,N_43970,N_43033);
or U46037 (N_46037,N_43713,N_40989);
xnor U46038 (N_46038,N_44531,N_43591);
and U46039 (N_46039,N_42258,N_43546);
nand U46040 (N_46040,N_40957,N_44652);
and U46041 (N_46041,N_40057,N_40339);
xnor U46042 (N_46042,N_43642,N_44389);
xnor U46043 (N_46043,N_44825,N_42376);
nor U46044 (N_46044,N_42684,N_40922);
xor U46045 (N_46045,N_43028,N_43125);
or U46046 (N_46046,N_42164,N_41642);
nor U46047 (N_46047,N_42888,N_44484);
xor U46048 (N_46048,N_43517,N_42168);
nand U46049 (N_46049,N_41730,N_42716);
xor U46050 (N_46050,N_44628,N_44194);
xnor U46051 (N_46051,N_42639,N_41829);
nor U46052 (N_46052,N_44385,N_42822);
xor U46053 (N_46053,N_40486,N_42451);
and U46054 (N_46054,N_40847,N_40821);
or U46055 (N_46055,N_43400,N_43495);
nor U46056 (N_46056,N_41658,N_44717);
and U46057 (N_46057,N_44475,N_42330);
nor U46058 (N_46058,N_41781,N_44622);
xor U46059 (N_46059,N_42422,N_44913);
or U46060 (N_46060,N_43320,N_41119);
nor U46061 (N_46061,N_40643,N_40539);
nand U46062 (N_46062,N_41159,N_43526);
nand U46063 (N_46063,N_43684,N_44087);
or U46064 (N_46064,N_44515,N_44834);
nand U46065 (N_46065,N_42501,N_42777);
xnor U46066 (N_46066,N_40604,N_42203);
xor U46067 (N_46067,N_40836,N_41166);
or U46068 (N_46068,N_40006,N_40765);
and U46069 (N_46069,N_42083,N_41137);
or U46070 (N_46070,N_40417,N_42900);
nand U46071 (N_46071,N_40599,N_42937);
xnor U46072 (N_46072,N_42329,N_40848);
nand U46073 (N_46073,N_44457,N_41230);
xor U46074 (N_46074,N_40871,N_43134);
or U46075 (N_46075,N_41898,N_43080);
or U46076 (N_46076,N_40924,N_41671);
xnor U46077 (N_46077,N_41813,N_44143);
xnor U46078 (N_46078,N_40224,N_44000);
or U46079 (N_46079,N_44003,N_43954);
xor U46080 (N_46080,N_42079,N_42205);
xnor U46081 (N_46081,N_42508,N_40110);
or U46082 (N_46082,N_43092,N_40319);
nor U46083 (N_46083,N_42051,N_41843);
nor U46084 (N_46084,N_43810,N_44734);
nor U46085 (N_46085,N_40453,N_44600);
nand U46086 (N_46086,N_42838,N_40968);
xnor U46087 (N_46087,N_43720,N_43588);
and U46088 (N_46088,N_42351,N_41333);
nor U46089 (N_46089,N_44393,N_42402);
nor U46090 (N_46090,N_41725,N_44589);
xor U46091 (N_46091,N_44216,N_41598);
nand U46092 (N_46092,N_40490,N_41491);
nand U46093 (N_46093,N_42761,N_40547);
nand U46094 (N_46094,N_42286,N_43729);
nand U46095 (N_46095,N_40149,N_40781);
and U46096 (N_46096,N_43334,N_42004);
or U46097 (N_46097,N_41592,N_42045);
nor U46098 (N_46098,N_44786,N_41395);
or U46099 (N_46099,N_41809,N_40856);
or U46100 (N_46100,N_41610,N_44218);
nor U46101 (N_46101,N_40907,N_43649);
xnor U46102 (N_46102,N_42050,N_43907);
and U46103 (N_46103,N_44978,N_42701);
or U46104 (N_46104,N_42538,N_43668);
nor U46105 (N_46105,N_43431,N_44398);
nor U46106 (N_46106,N_41180,N_42856);
nand U46107 (N_46107,N_40801,N_43782);
and U46108 (N_46108,N_40222,N_41869);
and U46109 (N_46109,N_43948,N_43748);
and U46110 (N_46110,N_42138,N_44516);
nor U46111 (N_46111,N_41553,N_41249);
nand U46112 (N_46112,N_43112,N_41663);
xnor U46113 (N_46113,N_42748,N_42883);
or U46114 (N_46114,N_44451,N_43742);
nand U46115 (N_46115,N_44082,N_42302);
and U46116 (N_46116,N_42897,N_41585);
and U46117 (N_46117,N_41256,N_42226);
and U46118 (N_46118,N_44671,N_40750);
nor U46119 (N_46119,N_40955,N_44259);
and U46120 (N_46120,N_41437,N_43995);
nor U46121 (N_46121,N_40391,N_42891);
xor U46122 (N_46122,N_43765,N_43965);
xnor U46123 (N_46123,N_40576,N_44208);
nor U46124 (N_46124,N_41053,N_43345);
nor U46125 (N_46125,N_43647,N_44670);
nand U46126 (N_46126,N_40250,N_40285);
and U46127 (N_46127,N_44525,N_42445);
nor U46128 (N_46128,N_43773,N_44880);
nor U46129 (N_46129,N_40082,N_40165);
xor U46130 (N_46130,N_42139,N_40941);
xnor U46131 (N_46131,N_43662,N_41806);
xnor U46132 (N_46132,N_40089,N_40371);
nor U46133 (N_46133,N_42044,N_43314);
nor U46134 (N_46134,N_41347,N_40823);
xor U46135 (N_46135,N_44084,N_44507);
and U46136 (N_46136,N_44710,N_41177);
xnor U46137 (N_46137,N_40300,N_44413);
nor U46138 (N_46138,N_42027,N_41619);
xor U46139 (N_46139,N_40535,N_44472);
or U46140 (N_46140,N_42687,N_43892);
xnor U46141 (N_46141,N_42803,N_42352);
nor U46142 (N_46142,N_40760,N_42353);
and U46143 (N_46143,N_41684,N_43305);
nand U46144 (N_46144,N_40705,N_44660);
xnor U46145 (N_46145,N_42981,N_41154);
xor U46146 (N_46146,N_43325,N_41961);
xnor U46147 (N_46147,N_40083,N_44138);
xnor U46148 (N_46148,N_43734,N_40944);
xor U46149 (N_46149,N_44227,N_44553);
xnor U46150 (N_46150,N_41188,N_44821);
xor U46151 (N_46151,N_41757,N_41758);
nand U46152 (N_46152,N_42585,N_40671);
and U46153 (N_46153,N_43774,N_44320);
xor U46154 (N_46154,N_40118,N_40087);
and U46155 (N_46155,N_40603,N_40363);
nand U46156 (N_46156,N_44376,N_42986);
nor U46157 (N_46157,N_44241,N_44304);
or U46158 (N_46158,N_41453,N_41380);
nor U46159 (N_46159,N_44474,N_41201);
and U46160 (N_46160,N_41528,N_40704);
nor U46161 (N_46161,N_41883,N_40565);
and U46162 (N_46162,N_43038,N_40292);
nand U46163 (N_46163,N_43381,N_43237);
nand U46164 (N_46164,N_44810,N_41240);
or U46165 (N_46165,N_42176,N_40953);
nand U46166 (N_46166,N_43412,N_44315);
nand U46167 (N_46167,N_41833,N_41383);
nor U46168 (N_46168,N_41677,N_40610);
xnor U46169 (N_46169,N_42120,N_44549);
and U46170 (N_46170,N_43956,N_40221);
and U46171 (N_46171,N_41038,N_44723);
or U46172 (N_46172,N_41673,N_42039);
and U46173 (N_46173,N_43986,N_44076);
nand U46174 (N_46174,N_42558,N_43286);
and U46175 (N_46175,N_40646,N_42010);
or U46176 (N_46176,N_40724,N_42917);
or U46177 (N_46177,N_43809,N_41422);
and U46178 (N_46178,N_43666,N_42055);
and U46179 (N_46179,N_40809,N_42433);
nand U46180 (N_46180,N_40992,N_41927);
and U46181 (N_46181,N_42475,N_40269);
or U46182 (N_46182,N_40824,N_43440);
nor U46183 (N_46183,N_43193,N_44926);
nand U46184 (N_46184,N_43936,N_44168);
nand U46185 (N_46185,N_40816,N_40019);
nand U46186 (N_46186,N_41193,N_40835);
nand U46187 (N_46187,N_42975,N_41374);
nor U46188 (N_46188,N_44915,N_43484);
and U46189 (N_46189,N_40481,N_43481);
nand U46190 (N_46190,N_43520,N_44497);
nor U46191 (N_46191,N_41640,N_41160);
xnor U46192 (N_46192,N_42237,N_41111);
xor U46193 (N_46193,N_41260,N_41060);
nor U46194 (N_46194,N_41027,N_40904);
xor U46195 (N_46195,N_42509,N_41524);
or U46196 (N_46196,N_43714,N_42142);
nor U46197 (N_46197,N_41182,N_40345);
and U46198 (N_46198,N_42001,N_41092);
and U46199 (N_46199,N_42442,N_42340);
and U46200 (N_46200,N_40722,N_43162);
and U46201 (N_46201,N_41718,N_41526);
and U46202 (N_46202,N_41747,N_43865);
and U46203 (N_46203,N_44592,N_43238);
nand U46204 (N_46204,N_42469,N_41822);
xnor U46205 (N_46205,N_42368,N_44648);
and U46206 (N_46206,N_44197,N_41225);
or U46207 (N_46207,N_43548,N_44854);
nor U46208 (N_46208,N_44707,N_42264);
nand U46209 (N_46209,N_43912,N_40133);
nand U46210 (N_46210,N_44139,N_43884);
xor U46211 (N_46211,N_40207,N_40917);
or U46212 (N_46212,N_43099,N_42026);
nor U46213 (N_46213,N_41474,N_40484);
nor U46214 (N_46214,N_42930,N_44113);
nand U46215 (N_46215,N_43929,N_41818);
nor U46216 (N_46216,N_41121,N_40844);
and U46217 (N_46217,N_43567,N_44510);
xnor U46218 (N_46218,N_40891,N_40276);
xor U46219 (N_46219,N_44323,N_43001);
xor U46220 (N_46220,N_43915,N_44594);
nand U46221 (N_46221,N_44842,N_43098);
or U46222 (N_46222,N_42919,N_42622);
nand U46223 (N_46223,N_43455,N_43853);
nand U46224 (N_46224,N_41872,N_44552);
and U46225 (N_46225,N_40153,N_40590);
nor U46226 (N_46226,N_44791,N_40315);
and U46227 (N_46227,N_41269,N_42090);
nand U46228 (N_46228,N_41626,N_40452);
and U46229 (N_46229,N_40354,N_44930);
and U46230 (N_46230,N_41003,N_44591);
nor U46231 (N_46231,N_40429,N_44430);
nand U46232 (N_46232,N_43086,N_40843);
nand U46233 (N_46233,N_42310,N_42092);
nand U46234 (N_46234,N_43296,N_43161);
nand U46235 (N_46235,N_41402,N_42965);
xnor U46236 (N_46236,N_44408,N_43128);
xor U46237 (N_46237,N_40455,N_40909);
nor U46238 (N_46238,N_43372,N_44203);
or U46239 (N_46239,N_43241,N_40388);
nor U46240 (N_46240,N_43234,N_40333);
and U46241 (N_46241,N_40383,N_41327);
and U46242 (N_46242,N_40373,N_42104);
or U46243 (N_46243,N_44580,N_41536);
xnor U46244 (N_46244,N_40562,N_44441);
xnor U46245 (N_46245,N_41679,N_42670);
xnor U46246 (N_46246,N_43497,N_43604);
and U46247 (N_46247,N_44932,N_43769);
xor U46248 (N_46248,N_42275,N_42846);
or U46249 (N_46249,N_40730,N_44386);
nor U46250 (N_46250,N_42850,N_40507);
and U46251 (N_46251,N_40731,N_41603);
and U46252 (N_46252,N_41098,N_42214);
nand U46253 (N_46253,N_43817,N_42317);
nor U46254 (N_46254,N_41131,N_44361);
nand U46255 (N_46255,N_41431,N_44447);
nor U46256 (N_46256,N_41686,N_40931);
or U46257 (N_46257,N_44992,N_41441);
nand U46258 (N_46258,N_44037,N_40017);
and U46259 (N_46259,N_40938,N_40011);
and U46260 (N_46260,N_41012,N_42169);
and U46261 (N_46261,N_43757,N_44962);
xor U46262 (N_46262,N_44365,N_40238);
nor U46263 (N_46263,N_42745,N_40549);
or U46264 (N_46264,N_41953,N_42375);
and U46265 (N_46265,N_44477,N_44454);
or U46266 (N_46266,N_41298,N_40430);
and U46267 (N_46267,N_42295,N_40695);
or U46268 (N_46268,N_40253,N_43643);
xnor U46269 (N_46269,N_44436,N_44268);
nor U46270 (N_46270,N_40126,N_40392);
or U46271 (N_46271,N_40227,N_44029);
xor U46272 (N_46272,N_40016,N_40282);
and U46273 (N_46273,N_44095,N_44925);
and U46274 (N_46274,N_42960,N_44427);
nor U46275 (N_46275,N_40652,N_44665);
and U46276 (N_46276,N_44089,N_43510);
nor U46277 (N_46277,N_42708,N_40357);
nand U46278 (N_46278,N_44422,N_44180);
nand U46279 (N_46279,N_41865,N_40802);
nand U46280 (N_46280,N_43091,N_43994);
xor U46281 (N_46281,N_43135,N_40266);
nor U46282 (N_46282,N_44654,N_43214);
xor U46283 (N_46283,N_41073,N_42496);
or U46284 (N_46284,N_44576,N_41317);
nand U46285 (N_46285,N_42712,N_40304);
nand U46286 (N_46286,N_44305,N_44907);
nand U46287 (N_46287,N_41442,N_41084);
nor U46288 (N_46288,N_43188,N_42132);
xnor U46289 (N_46289,N_44990,N_44409);
nand U46290 (N_46290,N_41896,N_42902);
nand U46291 (N_46291,N_42197,N_43053);
xnor U46292 (N_46292,N_43483,N_44165);
xnor U46293 (N_46293,N_41886,N_44129);
and U46294 (N_46294,N_40411,N_42515);
and U46295 (N_46295,N_40067,N_42113);
nor U46296 (N_46296,N_41142,N_42075);
nand U46297 (N_46297,N_43960,N_44864);
nand U46298 (N_46298,N_43971,N_44242);
nand U46299 (N_46299,N_40270,N_41970);
and U46300 (N_46300,N_44419,N_44721);
and U46301 (N_46301,N_42502,N_42772);
nand U46302 (N_46302,N_40163,N_43075);
and U46303 (N_46303,N_44918,N_41720);
and U46304 (N_46304,N_42313,N_41983);
nor U46305 (N_46305,N_42482,N_41057);
and U46306 (N_46306,N_44649,N_41070);
xor U46307 (N_46307,N_40935,N_42952);
and U46308 (N_46308,N_40742,N_42296);
or U46309 (N_46309,N_44166,N_43513);
and U46310 (N_46310,N_40262,N_41706);
nor U46311 (N_46311,N_42434,N_40969);
xnor U46312 (N_46312,N_44602,N_44415);
and U46313 (N_46313,N_40131,N_42876);
and U46314 (N_46314,N_42369,N_44455);
and U46315 (N_46315,N_43703,N_43812);
xor U46316 (N_46316,N_40205,N_43233);
nor U46317 (N_46317,N_41917,N_42595);
xor U46318 (N_46318,N_42077,N_43453);
nand U46319 (N_46319,N_42914,N_42640);
and U46320 (N_46320,N_44509,N_42178);
or U46321 (N_46321,N_40966,N_43599);
or U46322 (N_46322,N_42032,N_42194);
nand U46323 (N_46323,N_40015,N_40905);
and U46324 (N_46324,N_42213,N_41067);
xor U46325 (N_46325,N_42603,N_40991);
nand U46326 (N_46326,N_44053,N_44228);
or U46327 (N_46327,N_44191,N_40192);
nand U46328 (N_46328,N_42834,N_43575);
or U46329 (N_46329,N_43297,N_40582);
or U46330 (N_46330,N_42413,N_44506);
xor U46331 (N_46331,N_40735,N_44939);
nand U46332 (N_46332,N_40857,N_41954);
and U46333 (N_46333,N_40680,N_42589);
nand U46334 (N_46334,N_40617,N_43670);
nor U46335 (N_46335,N_41480,N_40620);
and U46336 (N_46336,N_41740,N_44690);
nand U46337 (N_46337,N_41226,N_41319);
nand U46338 (N_46338,N_40477,N_43317);
nand U46339 (N_46339,N_40571,N_42270);
nor U46340 (N_46340,N_44848,N_41957);
nor U46341 (N_46341,N_44107,N_44177);
nor U46342 (N_46342,N_41407,N_40068);
and U46343 (N_46343,N_44153,N_44570);
nand U46344 (N_46344,N_43274,N_44674);
or U46345 (N_46345,N_43157,N_41234);
or U46346 (N_46346,N_40248,N_41798);
or U46347 (N_46347,N_43644,N_44379);
and U46348 (N_46348,N_41190,N_41774);
xnor U46349 (N_46349,N_43223,N_44236);
or U46350 (N_46350,N_43756,N_41750);
and U46351 (N_46351,N_43847,N_42726);
and U46352 (N_46352,N_42719,N_44845);
nor U46353 (N_46353,N_43359,N_43498);
and U46354 (N_46354,N_43878,N_42102);
nor U46355 (N_46355,N_43254,N_43084);
nand U46356 (N_46356,N_42796,N_43499);
nor U46357 (N_46357,N_40081,N_40271);
xnor U46358 (N_46358,N_43919,N_40764);
and U46359 (N_46359,N_43999,N_43955);
and U46360 (N_46360,N_41179,N_42966);
and U46361 (N_46361,N_44099,N_43056);
nand U46362 (N_46362,N_42269,N_42184);
and U46363 (N_46363,N_44624,N_44483);
or U46364 (N_46364,N_43998,N_42105);
xnor U46365 (N_46365,N_42842,N_43180);
nor U46366 (N_46366,N_42166,N_40664);
and U46367 (N_46367,N_40958,N_43399);
and U46368 (N_46368,N_44529,N_41796);
or U46369 (N_46369,N_44640,N_42970);
nand U46370 (N_46370,N_40382,N_43996);
xor U46371 (N_46371,N_41743,N_43858);
or U46372 (N_46372,N_42201,N_44289);
and U46373 (N_46373,N_44253,N_41515);
xnor U46374 (N_46374,N_41353,N_42453);
xnor U46375 (N_46375,N_41949,N_43081);
and U46376 (N_46376,N_44355,N_43203);
nor U46377 (N_46377,N_41599,N_44554);
nand U46378 (N_46378,N_42866,N_40137);
nor U46379 (N_46379,N_40692,N_40159);
or U46380 (N_46380,N_40785,N_43992);
nor U46381 (N_46381,N_42911,N_42435);
nand U46382 (N_46382,N_43529,N_43176);
or U46383 (N_46383,N_42429,N_40889);
nor U46384 (N_46384,N_44806,N_42486);
xnor U46385 (N_46385,N_42522,N_42200);
and U46386 (N_46386,N_40741,N_43444);
xor U46387 (N_46387,N_42657,N_41488);
nor U46388 (N_46388,N_44190,N_43049);
nor U46389 (N_46389,N_43318,N_42898);
and U46390 (N_46390,N_40640,N_42059);
nand U46391 (N_46391,N_43235,N_41837);
xnor U46392 (N_46392,N_41320,N_41351);
nor U46393 (N_46393,N_43763,N_42206);
nor U46394 (N_46394,N_43328,N_43396);
nand U46395 (N_46395,N_44826,N_44851);
nor U46396 (N_46396,N_40182,N_41890);
nor U46397 (N_46397,N_44314,N_42115);
nand U46398 (N_46398,N_42593,N_42675);
xnor U46399 (N_46399,N_44577,N_42561);
xor U46400 (N_46400,N_44536,N_41932);
nand U46401 (N_46401,N_40314,N_42307);
nor U46402 (N_46402,N_43428,N_41384);
or U46403 (N_46403,N_43137,N_42165);
nand U46404 (N_46404,N_43409,N_40179);
or U46405 (N_46405,N_43089,N_43901);
nand U46406 (N_46406,N_44164,N_43043);
or U46407 (N_46407,N_43282,N_40929);
xor U46408 (N_46408,N_40203,N_44258);
xor U46409 (N_46409,N_41018,N_41044);
or U46410 (N_46410,N_42776,N_43900);
nor U46411 (N_46411,N_44713,N_41218);
nor U46412 (N_46412,N_43132,N_42959);
nand U46413 (N_46413,N_42288,N_40288);
nand U46414 (N_46414,N_41751,N_44160);
and U46415 (N_46415,N_41596,N_41532);
and U46416 (N_46416,N_40263,N_44811);
nor U46417 (N_46417,N_43931,N_43468);
xnor U46418 (N_46418,N_44831,N_44070);
or U46419 (N_46419,N_40260,N_40792);
and U46420 (N_46420,N_43824,N_42599);
and U46421 (N_46421,N_40469,N_40543);
nor U46422 (N_46422,N_44581,N_42680);
and U46423 (N_46423,N_41447,N_40976);
nand U46424 (N_46424,N_43728,N_43789);
nor U46425 (N_46425,N_42404,N_42807);
nand U46426 (N_46426,N_43628,N_44282);
nor U46427 (N_46427,N_40644,N_40568);
nor U46428 (N_46428,N_40591,N_40012);
nand U46429 (N_46429,N_40117,N_43106);
and U46430 (N_46430,N_42942,N_42241);
and U46431 (N_46431,N_41500,N_44341);
nor U46432 (N_46432,N_40053,N_42261);
and U46433 (N_46433,N_40035,N_42008);
nor U46434 (N_46434,N_42379,N_40551);
or U46435 (N_46435,N_44617,N_43398);
nor U46436 (N_46436,N_40952,N_40621);
nand U46437 (N_46437,N_42782,N_43252);
or U46438 (N_46438,N_43059,N_44230);
nor U46439 (N_46439,N_43600,N_44780);
and U46440 (N_46440,N_40690,N_42278);
and U46441 (N_46441,N_41908,N_41731);
nand U46442 (N_46442,N_41019,N_42617);
nand U46443 (N_46443,N_42342,N_42769);
xor U46444 (N_46444,N_44459,N_40100);
or U46445 (N_46445,N_41363,N_43679);
nor U46446 (N_46446,N_42764,N_43217);
nor U46447 (N_46447,N_40317,N_40229);
or U46448 (N_46448,N_43009,N_40489);
xor U46449 (N_46449,N_43211,N_44564);
nand U46450 (N_46450,N_40311,N_40554);
nor U46451 (N_46451,N_41627,N_40555);
xnor U46452 (N_46452,N_41307,N_44269);
or U46453 (N_46453,N_40234,N_43401);
xor U46454 (N_46454,N_41852,N_40379);
nor U46455 (N_46455,N_44938,N_40518);
or U46456 (N_46456,N_42706,N_42162);
nand U46457 (N_46457,N_41561,N_43541);
or U46458 (N_46458,N_40653,N_44185);
or U46459 (N_46459,N_42348,N_43979);
or U46460 (N_46460,N_42494,N_43925);
and U46461 (N_46461,N_42100,N_42664);
nand U46462 (N_46462,N_44548,N_41046);
or U46463 (N_46463,N_44827,N_41986);
xor U46464 (N_46464,N_42393,N_43256);
xor U46465 (N_46465,N_43872,N_41811);
or U46466 (N_46466,N_41513,N_42409);
nand U46467 (N_46467,N_40128,N_43799);
xnor U46468 (N_46468,N_40072,N_43932);
and U46469 (N_46469,N_43355,N_44587);
nand U46470 (N_46470,N_40689,N_41368);
and U46471 (N_46471,N_44987,N_42478);
and U46472 (N_46472,N_44746,N_40360);
nor U46473 (N_46473,N_41079,N_43027);
nor U46474 (N_46474,N_42632,N_40185);
or U46475 (N_46475,N_43012,N_41493);
nand U46476 (N_46476,N_43168,N_41788);
nand U46477 (N_46477,N_44458,N_40225);
nand U46478 (N_46478,N_40025,N_44802);
xor U46479 (N_46479,N_44276,N_43547);
nor U46480 (N_46480,N_40506,N_42210);
or U46481 (N_46481,N_42988,N_40198);
and U46482 (N_46482,N_40141,N_44960);
and U46483 (N_46483,N_44731,N_44039);
or U46484 (N_46484,N_43930,N_40024);
nor U46485 (N_46485,N_40930,N_41565);
and U46486 (N_46486,N_41050,N_42371);
xor U46487 (N_46487,N_43700,N_42291);
nand U46488 (N_46488,N_42222,N_43149);
nor U46489 (N_46489,N_44211,N_42720);
nor U46490 (N_46490,N_41456,N_41428);
nand U46491 (N_46491,N_44500,N_44597);
nor U46492 (N_46492,N_44774,N_44524);
xnor U46493 (N_46493,N_43331,N_44807);
xnor U46494 (N_46494,N_42372,N_44257);
or U46495 (N_46495,N_44152,N_40654);
nor U46496 (N_46496,N_42259,N_43118);
xor U46497 (N_46497,N_43741,N_42196);
or U46498 (N_46498,N_43564,N_44034);
xnor U46499 (N_46499,N_43630,N_40526);
xnor U46500 (N_46500,N_43261,N_43348);
and U46501 (N_46501,N_40758,N_43022);
xnor U46502 (N_46502,N_41816,N_41239);
xor U46503 (N_46503,N_41647,N_44605);
or U46504 (N_46504,N_44667,N_41094);
nor U46505 (N_46505,N_40867,N_44092);
and U46506 (N_46506,N_41643,N_40461);
and U46507 (N_46507,N_40858,N_43660);
and U46508 (N_46508,N_43803,N_42805);
or U46509 (N_46509,N_40334,N_40158);
and U46510 (N_46510,N_44979,N_40318);
nand U46511 (N_46511,N_42378,N_43923);
xor U46512 (N_46512,N_40766,N_44823);
and U46513 (N_46513,N_41030,N_41455);
or U46514 (N_46514,N_42441,N_40138);
or U46515 (N_46515,N_44678,N_40164);
nand U46516 (N_46516,N_43885,N_44476);
nor U46517 (N_46517,N_44585,N_42002);
xor U46518 (N_46518,N_40775,N_41187);
nor U46519 (N_46519,N_41590,N_44251);
and U46520 (N_46520,N_41930,N_42728);
and U46521 (N_46521,N_44977,N_43537);
xnor U46522 (N_46522,N_42750,N_40355);
xnor U46523 (N_46523,N_41830,N_40385);
nand U46524 (N_46524,N_44933,N_42072);
xor U46525 (N_46525,N_44429,N_43776);
and U46526 (N_46526,N_41967,N_44630);
or U46527 (N_46527,N_43959,N_42713);
and U46528 (N_46528,N_44317,N_42383);
or U46529 (N_46529,N_42923,N_44805);
and U46530 (N_46530,N_44229,N_41735);
nand U46531 (N_46531,N_40657,N_43894);
xnor U46532 (N_46532,N_44711,N_43990);
nor U46533 (N_46533,N_42696,N_42646);
nor U46534 (N_46534,N_41210,N_43068);
nand U46535 (N_46535,N_41181,N_43018);
nand U46536 (N_46536,N_44790,N_40763);
nor U46537 (N_46537,N_42048,N_43133);
nor U46538 (N_46538,N_44699,N_42736);
nand U46539 (N_46539,N_40532,N_41748);
nor U46540 (N_46540,N_42253,N_43026);
xnor U46541 (N_46541,N_44904,N_43893);
xnor U46542 (N_46542,N_42119,N_40710);
and U46543 (N_46543,N_41360,N_44491);
xnor U46544 (N_46544,N_41344,N_43562);
nor U46545 (N_46545,N_41357,N_44252);
or U46546 (N_46546,N_44270,N_44017);
and U46547 (N_46547,N_43657,N_42454);
and U46548 (N_46548,N_44964,N_43606);
and U46549 (N_46549,N_42527,N_43864);
nor U46550 (N_46550,N_42550,N_40080);
xor U46551 (N_46551,N_40093,N_44575);
or U46552 (N_46552,N_43524,N_44940);
nor U46553 (N_46553,N_44406,N_41272);
and U46554 (N_46554,N_41688,N_42000);
nor U46555 (N_46555,N_41194,N_40533);
or U46556 (N_46556,N_41535,N_42495);
nand U46557 (N_46557,N_44623,N_43154);
xor U46558 (N_46558,N_40428,N_41143);
xnor U46559 (N_46559,N_44993,N_42683);
nor U46560 (N_46560,N_41831,N_44632);
xnor U46561 (N_46561,N_44048,N_40694);
nor U46562 (N_46562,N_44975,N_40094);
nor U46563 (N_46563,N_40468,N_42279);
or U46564 (N_46564,N_42964,N_41577);
or U46565 (N_46565,N_43120,N_42980);
or U46566 (N_46566,N_40999,N_41836);
nand U46567 (N_46567,N_44808,N_40612);
nor U46568 (N_46568,N_42929,N_41397);
nand U46569 (N_46569,N_42933,N_40114);
and U46570 (N_46570,N_43721,N_43491);
and U46571 (N_46571,N_44794,N_43518);
nor U46572 (N_46572,N_44106,N_43478);
and U46573 (N_46573,N_43658,N_42128);
nand U46574 (N_46574,N_42086,N_43153);
nand U46575 (N_46575,N_43727,N_40440);
xnor U46576 (N_46576,N_42389,N_40517);
xor U46577 (N_46577,N_43770,N_42439);
and U46578 (N_46578,N_44838,N_42242);
xnor U46579 (N_46579,N_43687,N_40932);
nor U46580 (N_46580,N_42572,N_43190);
xor U46581 (N_46581,N_40598,N_41609);
nor U46582 (N_46582,N_42679,N_42992);
and U46583 (N_46583,N_42147,N_41074);
nor U46584 (N_46584,N_44343,N_44402);
or U46585 (N_46585,N_44673,N_44732);
nand U46586 (N_46586,N_42013,N_43055);
xor U46587 (N_46587,N_41404,N_43502);
or U46588 (N_46588,N_40152,N_43969);
and U46589 (N_46589,N_40661,N_41616);
nor U46590 (N_46590,N_43823,N_42316);
nand U46591 (N_46591,N_41724,N_44288);
or U46592 (N_46592,N_40033,N_40510);
and U46593 (N_46593,N_40183,N_43166);
and U46594 (N_46594,N_44609,N_42257);
and U46595 (N_46595,N_42229,N_41859);
and U46596 (N_46596,N_40046,N_43206);
and U46597 (N_46597,N_41417,N_40588);
nand U46598 (N_46598,N_44245,N_41343);
nor U46599 (N_46599,N_42065,N_40749);
and U46600 (N_46600,N_42760,N_41916);
xor U46601 (N_46601,N_43311,N_41113);
xnor U46602 (N_46602,N_42054,N_44403);
xor U46603 (N_46603,N_44697,N_42814);
and U46604 (N_46604,N_41876,N_44373);
and U46605 (N_46605,N_43845,N_40519);
and U46606 (N_46606,N_41035,N_43867);
nand U46607 (N_46607,N_41168,N_42151);
nor U46608 (N_46608,N_41672,N_42159);
or U46609 (N_46609,N_41929,N_42461);
nand U46610 (N_46610,N_44423,N_44418);
and U46611 (N_46611,N_40487,N_41017);
nor U46612 (N_46612,N_44885,N_41243);
or U46613 (N_46613,N_40723,N_40524);
and U46614 (N_46614,N_41391,N_43939);
xor U46615 (N_46615,N_41841,N_40973);
xor U46616 (N_46616,N_42049,N_41849);
or U46617 (N_46617,N_42481,N_41894);
or U46618 (N_46618,N_42236,N_44584);
or U46619 (N_46619,N_43601,N_42400);
nor U46620 (N_46620,N_41925,N_42812);
xnor U46621 (N_46621,N_42323,N_43556);
xor U46622 (N_46622,N_40199,N_42998);
and U46623 (N_46623,N_40508,N_41897);
or U46624 (N_46624,N_44467,N_42698);
nor U46625 (N_46625,N_43895,N_42406);
and U46626 (N_46626,N_40032,N_41998);
and U46627 (N_46627,N_43179,N_42832);
and U46628 (N_46628,N_40798,N_40915);
nand U46629 (N_46629,N_42647,N_41586);
or U46630 (N_46630,N_40639,N_41601);
or U46631 (N_46631,N_44044,N_44739);
xor U46632 (N_46632,N_41973,N_44210);
xor U46633 (N_46633,N_43800,N_40975);
nand U46634 (N_46634,N_41584,N_44709);
nor U46635 (N_46635,N_41989,N_43779);
or U46636 (N_46636,N_41877,N_40830);
and U46637 (N_46637,N_44200,N_43725);
or U46638 (N_46638,N_42245,N_43870);
nand U46639 (N_46639,N_41517,N_43938);
xnor U46640 (N_46640,N_44167,N_40701);
nor U46641 (N_46641,N_40043,N_40474);
and U46642 (N_46642,N_42505,N_42565);
and U46643 (N_46643,N_41710,N_43974);
nand U46644 (N_46644,N_41847,N_41439);
and U46645 (N_46645,N_43808,N_42327);
nand U46646 (N_46646,N_42024,N_42488);
xor U46647 (N_46647,N_40050,N_42096);
and U46648 (N_46648,N_42549,N_40799);
and U46649 (N_46649,N_40626,N_43146);
xor U46650 (N_46650,N_44100,N_41403);
and U46651 (N_46651,N_43489,N_44681);
nor U46652 (N_46652,N_44912,N_40948);
nand U46653 (N_46653,N_42857,N_42997);
xnor U46654 (N_46654,N_40505,N_44277);
nor U46655 (N_46655,N_41325,N_43014);
xor U46656 (N_46656,N_42246,N_41095);
nor U46657 (N_46657,N_44041,N_40897);
nor U46658 (N_46658,N_44804,N_40893);
and U46659 (N_46659,N_43205,N_41049);
or U46660 (N_46660,N_43373,N_40069);
xor U46661 (N_46661,N_43664,N_41338);
xor U46662 (N_46662,N_41808,N_42293);
nand U46663 (N_46663,N_40193,N_43532);
or U46664 (N_46664,N_43659,N_43968);
nand U46665 (N_46665,N_43719,N_40313);
and U46666 (N_46666,N_44173,N_42843);
and U46667 (N_46667,N_43437,N_44223);
or U46668 (N_46668,N_40769,N_42140);
and U46669 (N_46669,N_43392,N_43363);
xor U46670 (N_46670,N_41324,N_44480);
nand U46671 (N_46671,N_41462,N_41738);
xor U46672 (N_46672,N_42799,N_44982);
nor U46673 (N_46673,N_43160,N_41253);
nor U46674 (N_46674,N_44539,N_44748);
and U46675 (N_46675,N_41128,N_44563);
nand U46676 (N_46676,N_41321,N_44863);
and U46677 (N_46677,N_41064,N_44209);
and U46678 (N_46678,N_40593,N_40787);
and U46679 (N_46679,N_40103,N_44424);
xor U46680 (N_46680,N_40793,N_44664);
nand U46681 (N_46681,N_43351,N_42922);
nand U46682 (N_46682,N_43220,N_41007);
nor U46683 (N_46683,N_41719,N_44906);
or U46684 (N_46684,N_42871,N_41614);
nor U46685 (N_46685,N_44745,N_43448);
or U46686 (N_46686,N_44695,N_42896);
or U46687 (N_46687,N_43005,N_44381);
and U46688 (N_46688,N_42431,N_44843);
and U46689 (N_46689,N_42563,N_41845);
and U46690 (N_46690,N_43832,N_41621);
xnor U46691 (N_46691,N_41420,N_41306);
or U46692 (N_46692,N_44198,N_40279);
nand U46693 (N_46693,N_40687,N_40813);
or U46694 (N_46694,N_41924,N_40762);
nor U46695 (N_46695,N_41316,N_41004);
xor U46696 (N_46696,N_40528,N_44349);
nor U46697 (N_46697,N_40560,N_41186);
nand U46698 (N_46698,N_41749,N_41863);
nand U46699 (N_46699,N_40641,N_44954);
nand U46700 (N_46700,N_40702,N_40903);
nand U46701 (N_46701,N_43152,N_41155);
xnor U46702 (N_46702,N_40911,N_40838);
and U46703 (N_46703,N_44676,N_40685);
and U46704 (N_46704,N_43242,N_42459);
nor U46705 (N_46705,N_43287,N_42061);
xnor U46706 (N_46706,N_41029,N_43530);
or U46707 (N_46707,N_42146,N_44595);
or U46708 (N_46708,N_44453,N_44226);
nand U46709 (N_46709,N_42528,N_43382);
xnor U46710 (N_46710,N_42757,N_43791);
xnor U46711 (N_46711,N_43402,N_42662);
and U46712 (N_46712,N_44542,N_42530);
and U46713 (N_46713,N_40883,N_41285);
nor U46714 (N_46714,N_42743,N_40921);
or U46715 (N_46715,N_42872,N_42112);
or U46716 (N_46716,N_40713,N_40249);
xnor U46717 (N_46717,N_44945,N_41765);
xor U46718 (N_46718,N_41568,N_44135);
and U46719 (N_46719,N_44633,N_41072);
and U46720 (N_46720,N_40668,N_43991);
xnor U46721 (N_46721,N_44760,N_40774);
nand U46722 (N_46722,N_41322,N_40460);
nand U46723 (N_46723,N_44015,N_44023);
xor U46724 (N_46724,N_43735,N_40861);
nor U46725 (N_46725,N_42547,N_43570);
and U46726 (N_46726,N_44286,N_40120);
or U46727 (N_46727,N_44789,N_40272);
nand U46728 (N_46728,N_40000,N_44495);
or U46729 (N_46729,N_40473,N_43752);
nand U46730 (N_46730,N_44473,N_41443);
nor U46731 (N_46731,N_42274,N_43549);
nand U46732 (N_46732,N_41582,N_42514);
and U46733 (N_46733,N_44234,N_43980);
nor U46734 (N_46734,N_44858,N_40405);
nand U46735 (N_46735,N_40214,N_42849);
xnor U46736 (N_46736,N_41881,N_44358);
xnor U46737 (N_46737,N_42882,N_44765);
xor U46738 (N_46738,N_44428,N_40744);
xor U46739 (N_46739,N_41844,N_40330);
and U46740 (N_46740,N_43506,N_43804);
or U46741 (N_46741,N_44718,N_44692);
or U46742 (N_46742,N_40852,N_40803);
and U46743 (N_46743,N_40912,N_44700);
or U46744 (N_46744,N_41670,N_41468);
and U46745 (N_46745,N_40592,N_42568);
and U46746 (N_46746,N_41979,N_41509);
xor U46747 (N_46747,N_41227,N_40376);
or U46748 (N_46748,N_40747,N_40806);
nand U46749 (N_46749,N_43523,N_42030);
or U46750 (N_46750,N_42976,N_42605);
nor U46751 (N_46751,N_43273,N_43944);
or U46752 (N_46752,N_40139,N_44523);
nand U46753 (N_46753,N_44899,N_40614);
nor U46754 (N_46754,N_41803,N_44359);
nand U46755 (N_46755,N_40825,N_42028);
xor U46756 (N_46756,N_41281,N_41570);
nor U46757 (N_46757,N_40845,N_44599);
and U46758 (N_46758,N_40708,N_43215);
or U46759 (N_46759,N_42143,N_40365);
nor U46760 (N_46760,N_41153,N_41864);
nand U46761 (N_46761,N_40633,N_42945);
or U46762 (N_46762,N_42347,N_44985);
nand U46763 (N_46763,N_43461,N_41762);
or U46764 (N_46764,N_42737,N_44812);
or U46765 (N_46765,N_40800,N_42574);
xnor U46766 (N_46766,N_41313,N_44725);
nor U46767 (N_46767,N_43191,N_41753);
nand U46768 (N_46768,N_43390,N_41745);
nand U46769 (N_46769,N_43972,N_44669);
and U46770 (N_46770,N_42394,N_42238);
nand U46771 (N_46771,N_43626,N_44610);
nor U46772 (N_46772,N_42863,N_43859);
and U46773 (N_46773,N_42623,N_40832);
and U46774 (N_46774,N_43140,N_42749);
or U46775 (N_46775,N_44348,N_41653);
nor U46776 (N_46776,N_42810,N_41033);
nor U46777 (N_46777,N_41858,N_44487);
nor U46778 (N_46778,N_41545,N_42924);
and U46779 (N_46779,N_40233,N_44136);
or U46780 (N_46780,N_44701,N_42234);
nor U46781 (N_46781,N_40077,N_43953);
nor U46782 (N_46782,N_44465,N_41199);
or U46783 (N_46783,N_40007,N_44636);
nor U46784 (N_46784,N_41484,N_43292);
nand U46785 (N_46785,N_40751,N_43063);
or U46786 (N_46786,N_40084,N_40242);
nor U46787 (N_46787,N_44969,N_44433);
and U46788 (N_46788,N_40097,N_42787);
and U46789 (N_46789,N_43711,N_42594);
xor U46790 (N_46790,N_40642,N_41909);
nor U46791 (N_46791,N_43187,N_41856);
xnor U46792 (N_46792,N_41573,N_43102);
xnor U46793 (N_46793,N_40106,N_42192);
or U46794 (N_46794,N_40757,N_44261);
xor U46795 (N_46795,N_43239,N_44637);
and U46796 (N_46796,N_41815,N_41819);
nand U46797 (N_46797,N_41171,N_43775);
nand U46798 (N_46798,N_43716,N_40908);
or U46799 (N_46799,N_40393,N_43558);
and U46800 (N_46800,N_40546,N_40556);
and U46801 (N_46801,N_41934,N_41122);
nand U46802 (N_46802,N_43795,N_42537);
or U46803 (N_46803,N_44494,N_42349);
nor U46804 (N_46804,N_43249,N_43361);
nand U46805 (N_46805,N_42768,N_43380);
or U46806 (N_46806,N_44250,N_42524);
nand U46807 (N_46807,N_40085,N_44170);
nor U46808 (N_46808,N_40971,N_43229);
xnor U46809 (N_46809,N_41638,N_44335);
and U46810 (N_46810,N_40209,N_44322);
and U46811 (N_46811,N_43542,N_43785);
xor U46812 (N_46812,N_44479,N_40860);
nand U46813 (N_46813,N_41996,N_43039);
nor U46814 (N_46814,N_44263,N_43113);
and U46815 (N_46815,N_40431,N_44706);
nor U46816 (N_46816,N_44443,N_44047);
or U46817 (N_46817,N_42845,N_44144);
nand U46818 (N_46818,N_41486,N_40048);
nor U46819 (N_46819,N_40607,N_42038);
nor U46820 (N_46820,N_43008,N_44337);
or U46821 (N_46821,N_43801,N_42260);
and U46822 (N_46822,N_41426,N_44122);
nand U46823 (N_46823,N_44401,N_43515);
and U46824 (N_46824,N_42289,N_42443);
or U46825 (N_46825,N_42117,N_43829);
and U46826 (N_46826,N_43709,N_40064);
xor U46827 (N_46827,N_44518,N_41981);
xnor U46828 (N_46828,N_43150,N_42548);
xnor U46829 (N_46829,N_40346,N_41606);
nand U46830 (N_46830,N_40736,N_44619);
nor U46831 (N_46831,N_40866,N_44410);
nor U46832 (N_46832,N_43891,N_40686);
and U46833 (N_46833,N_44704,N_40715);
xor U46834 (N_46834,N_42047,N_40956);
nand U46835 (N_46835,N_44541,N_42121);
nor U46836 (N_46836,N_41157,N_40251);
and U46837 (N_46837,N_41217,N_41265);
nand U46838 (N_46838,N_41011,N_41512);
nand U46839 (N_46839,N_40425,N_42282);
or U46840 (N_46840,N_44232,N_42240);
and U46841 (N_46841,N_41149,N_42071);
xnor U46842 (N_46842,N_41984,N_41705);
nand U46843 (N_46843,N_41304,N_44951);
and U46844 (N_46844,N_42569,N_44254);
nand U46845 (N_46845,N_40441,N_41503);
or U46846 (N_46846,N_44590,N_43212);
and U46847 (N_46847,N_41945,N_42823);
nand U46848 (N_46848,N_43480,N_40298);
nand U46849 (N_46849,N_44944,N_43952);
and U46850 (N_46850,N_43874,N_42315);
and U46851 (N_46851,N_40208,N_42880);
nand U46852 (N_46852,N_41563,N_43388);
nor U46853 (N_46853,N_40842,N_42955);
nor U46854 (N_46854,N_44246,N_43275);
xnor U46855 (N_46855,N_42848,N_41931);
nor U46856 (N_46856,N_43943,N_40504);
nor U46857 (N_46857,N_42324,N_44503);
nor U46858 (N_46858,N_41236,N_44757);
xor U46859 (N_46859,N_42673,N_40400);
or U46860 (N_46860,N_44463,N_40520);
xor U46861 (N_46861,N_44184,N_42629);
nand U46862 (N_46862,N_42129,N_41340);
nand U46863 (N_46863,N_40003,N_42085);
nand U46864 (N_46864,N_44291,N_41215);
or U46865 (N_46865,N_44565,N_44752);
nand U46866 (N_46866,N_43303,N_42093);
nor U46867 (N_46867,N_43876,N_41246);
or U46868 (N_46868,N_42753,N_40811);
nor U46869 (N_46869,N_41197,N_42649);
and U46870 (N_46870,N_42498,N_44603);
or U46871 (N_46871,N_44145,N_44111);
or U46872 (N_46872,N_43917,N_43838);
xnor U46873 (N_46873,N_43427,N_43283);
xnor U46874 (N_46874,N_43612,N_43218);
nor U46875 (N_46875,N_41769,N_42321);
xor U46876 (N_46876,N_40662,N_41348);
xnor U46877 (N_46877,N_44233,N_42056);
nand U46878 (N_46878,N_42744,N_40777);
and U46879 (N_46879,N_40291,N_44820);
nand U46880 (N_46880,N_41646,N_40102);
and U46881 (N_46881,N_44836,N_43093);
nor U46882 (N_46882,N_41387,N_44222);
xnor U46883 (N_46883,N_41031,N_40235);
nor U46884 (N_46884,N_40959,N_43940);
nor U46885 (N_46885,N_40478,N_43294);
nand U46886 (N_46886,N_43947,N_40211);
and U46887 (N_46887,N_40597,N_40217);
nor U46888 (N_46888,N_40154,N_44783);
or U46889 (N_46889,N_41196,N_40174);
or U46890 (N_46890,N_42920,N_42426);
and U46891 (N_46891,N_42738,N_44205);
or U46892 (N_46892,N_43258,N_44326);
or U46893 (N_46893,N_40558,N_43732);
nor U46894 (N_46894,N_44469,N_40099);
nand U46895 (N_46895,N_42127,N_40732);
nor U46896 (N_46896,N_44530,N_43248);
or U46897 (N_46897,N_41107,N_40746);
or U46898 (N_46898,N_43074,N_40501);
xnor U46899 (N_46899,N_44522,N_40663);
or U46900 (N_46900,N_44488,N_41326);
and U46901 (N_46901,N_40171,N_41701);
nor U46902 (N_46902,N_44151,N_41613);
nand U46903 (N_46903,N_44058,N_42355);
or U46904 (N_46904,N_44238,N_41498);
nor U46905 (N_46905,N_42190,N_43942);
nor U46906 (N_46906,N_42460,N_40495);
or U46907 (N_46907,N_43918,N_41271);
xor U46908 (N_46908,N_41040,N_41330);
nand U46909 (N_46909,N_44215,N_43848);
nand U46910 (N_46910,N_40336,N_43379);
nand U46911 (N_46911,N_44866,N_43988);
nor U46912 (N_46912,N_44353,N_40284);
nand U46913 (N_46913,N_40297,N_42248);
nand U46914 (N_46914,N_43613,N_40987);
nand U46915 (N_46915,N_44178,N_41542);
or U46916 (N_46916,N_44694,N_43977);
xnor U46917 (N_46917,N_43507,N_43521);
or U46918 (N_46918,N_41492,N_43646);
xnor U46919 (N_46919,N_44770,N_42244);
or U46920 (N_46920,N_42635,N_41990);
nand U46921 (N_46921,N_42879,N_41666);
nor U46922 (N_46922,N_42831,N_44882);
nor U46923 (N_46923,N_41161,N_44192);
nand U46924 (N_46924,N_41926,N_42790);
and U46925 (N_46925,N_41737,N_41722);
nand U46926 (N_46926,N_40594,N_42853);
or U46927 (N_46927,N_43155,N_43509);
nand U46928 (N_46928,N_43466,N_42865);
nor U46929 (N_46929,N_40350,N_40920);
nor U46930 (N_46930,N_43906,N_40859);
nor U46931 (N_46931,N_41736,N_40669);
or U46932 (N_46932,N_40196,N_44108);
xor U46933 (N_46933,N_42373,N_43470);
nor U46934 (N_46934,N_40629,N_41247);
nand U46935 (N_46935,N_42273,N_44420);
nor U46936 (N_46936,N_43460,N_43119);
and U46937 (N_46937,N_40863,N_40395);
or U46938 (N_46938,N_40962,N_43129);
nor U46939 (N_46939,N_44693,N_42025);
nand U46940 (N_46940,N_43308,N_43031);
or U46941 (N_46941,N_41623,N_42671);
or U46942 (N_46942,N_44873,N_41885);
nor U46943 (N_46943,N_42185,N_41156);
or U46944 (N_46944,N_43908,N_42847);
nor U46945 (N_46945,N_43951,N_44013);
nor U46946 (N_46946,N_42742,N_40172);
nor U46947 (N_46947,N_42781,N_40157);
nor U46948 (N_46948,N_42821,N_41198);
and U46949 (N_46949,N_43723,N_40561);
nor U46950 (N_46950,N_44127,N_42854);
or U46951 (N_46951,N_42198,N_44753);
or U46952 (N_46952,N_41277,N_42467);
xor U46953 (N_46953,N_43527,N_41698);
or U46954 (N_46954,N_40525,N_41202);
and U46955 (N_46955,N_42835,N_43551);
or U46956 (N_46956,N_41807,N_42365);
nand U46957 (N_46957,N_44663,N_42362);
or U46958 (N_46958,N_44067,N_43375);
xor U46959 (N_46959,N_43439,N_42852);
nand U46960 (N_46960,N_43061,N_40720);
nor U46961 (N_46961,N_43016,N_41785);
xor U46962 (N_46962,N_44698,N_42057);
and U46963 (N_46963,N_40914,N_40052);
nand U46964 (N_46964,N_43253,N_43787);
nand U46965 (N_46965,N_44006,N_43057);
or U46966 (N_46966,N_42211,N_43699);
nor U46967 (N_46967,N_44464,N_44803);
and U46968 (N_46968,N_44788,N_42546);
nand U46969 (N_46969,N_43173,N_41562);
xor U46970 (N_46970,N_43635,N_44627);
xor U46971 (N_46971,N_41997,N_43167);
and U46972 (N_46972,N_42932,N_44538);
xor U46973 (N_46973,N_44114,N_42695);
xor U46974 (N_46974,N_44889,N_41756);
xor U46975 (N_46975,N_40294,N_44869);
xnor U46976 (N_46976,N_44502,N_44573);
xnor U46977 (N_46977,N_44363,N_42007);
xnor U46978 (N_46978,N_43224,N_44703);
or U46979 (N_46979,N_44217,N_42792);
nor U46980 (N_46980,N_44435,N_41895);
or U46981 (N_46981,N_41001,N_43109);
or U46982 (N_46982,N_43897,N_40356);
or U46983 (N_46983,N_40540,N_40697);
xnor U46984 (N_46984,N_42862,N_44278);
nand U46985 (N_46985,N_40226,N_42177);
or U46986 (N_46986,N_43025,N_44588);
nor U46987 (N_46987,N_44751,N_42489);
nand U46988 (N_46988,N_42573,N_40681);
nor U46989 (N_46989,N_44955,N_42949);
and U46990 (N_46990,N_44119,N_41235);
nand U46991 (N_46991,N_43511,N_41566);
nor U46992 (N_46992,N_40728,N_40878);
nand U46993 (N_46993,N_42583,N_40204);
nand U46994 (N_46994,N_40335,N_41352);
or U46995 (N_46995,N_41466,N_40036);
nor U46996 (N_46996,N_42674,N_42466);
xor U46997 (N_46997,N_43516,N_44965);
nor U46998 (N_46998,N_44878,N_40324);
nor U46999 (N_46999,N_44149,N_43324);
nor U47000 (N_47000,N_42366,N_44772);
xnor U47001 (N_47001,N_41222,N_41427);
xor U47002 (N_47002,N_43706,N_44953);
nor U47003 (N_47003,N_42212,N_44742);
xnor U47004 (N_47004,N_41966,N_44672);
nor U47005 (N_47005,N_40699,N_43143);
nor U47006 (N_47006,N_44833,N_40933);
nand U47007 (N_47007,N_40595,N_43633);
or U47008 (N_47008,N_43856,N_41126);
nand U47009 (N_47009,N_42080,N_42503);
xnor U47010 (N_47010,N_40726,N_40683);
or U47011 (N_47011,N_44755,N_42710);
xnor U47012 (N_47012,N_43560,N_42614);
nor U47013 (N_47013,N_42221,N_41411);
nand U47014 (N_47014,N_41649,N_41008);
or U47015 (N_47015,N_41696,N_43528);
or U47016 (N_47016,N_42063,N_40189);
or U47017 (N_47017,N_41415,N_44033);
or U47018 (N_47018,N_44689,N_43903);
and U47019 (N_47019,N_42338,N_43927);
or U47020 (N_47020,N_44086,N_40130);
nor U47021 (N_47021,N_40256,N_42457);
nand U47022 (N_47022,N_42204,N_44395);
nand U47023 (N_47023,N_44877,N_40277);
nor U47024 (N_47024,N_41988,N_44855);
or U47025 (N_47025,N_43928,N_41497);
xor U47026 (N_47026,N_41091,N_43899);
or U47027 (N_47027,N_40873,N_41051);
nand U47028 (N_47028,N_41334,N_41759);
and U47029 (N_47029,N_43565,N_42250);
nor U47030 (N_47030,N_44646,N_43259);
and U47031 (N_47031,N_42669,N_41980);
nand U47032 (N_47032,N_44941,N_43124);
and U47033 (N_47033,N_44157,N_40698);
or U47034 (N_47034,N_40739,N_43861);
and U47035 (N_47035,N_40200,N_44849);
or U47036 (N_47036,N_43065,N_44970);
and U47037 (N_47037,N_42634,N_42150);
xor U47038 (N_47038,N_41232,N_41795);
and U47039 (N_47039,N_41936,N_44219);
or U47040 (N_47040,N_44647,N_44255);
xor U47041 (N_47041,N_42277,N_41546);
or U47042 (N_47042,N_41189,N_41951);
xor U47043 (N_47043,N_40940,N_41114);
and U47044 (N_47044,N_43737,N_42711);
nand U47045 (N_47045,N_43228,N_43631);
nor U47046 (N_47046,N_42062,N_42114);
and U47047 (N_47047,N_41971,N_43584);
or U47048 (N_47048,N_40587,N_43689);
xnor U47049 (N_47049,N_43442,N_41371);
xor U47050 (N_47050,N_41595,N_43070);
nor U47051 (N_47051,N_44072,N_44016);
and U47052 (N_47052,N_43069,N_40580);
or U47053 (N_47053,N_43623,N_40444);
nor U47054 (N_47054,N_41835,N_42290);
nand U47055 (N_47055,N_44871,N_44388);
nor U47056 (N_47056,N_44334,N_44470);
and U47057 (N_47057,N_44771,N_42956);
or U47058 (N_47058,N_44214,N_42510);
xor U47059 (N_47059,N_43587,N_41080);
and U47060 (N_47060,N_41527,N_41086);
nor U47061 (N_47061,N_41506,N_44148);
xor U47062 (N_47062,N_40926,N_42019);
xnor U47063 (N_47063,N_42009,N_40804);
nor U47064 (N_47064,N_40693,N_44116);
nor U47065 (N_47065,N_40665,N_43142);
xor U47066 (N_47066,N_40563,N_41880);
xor U47067 (N_47067,N_41337,N_40370);
xor U47068 (N_47068,N_42483,N_42005);
xnor U47069 (N_47069,N_40575,N_42276);
and U47070 (N_47070,N_42125,N_42173);
nor U47071 (N_47071,N_40347,N_44280);
nor U47072 (N_47072,N_41797,N_40725);
and U47073 (N_47073,N_41714,N_41746);
xor U47074 (N_47074,N_40420,N_41964);
and U47075 (N_47075,N_42693,N_43449);
or U47076 (N_47076,N_44840,N_44366);
and U47077 (N_47077,N_43456,N_41976);
nand U47078 (N_47078,N_41279,N_40755);
nand U47079 (N_47079,N_42227,N_44607);
and U47080 (N_47080,N_40536,N_44911);
or U47081 (N_47081,N_41206,N_40670);
nand U47082 (N_47082,N_40807,N_43126);
and U47083 (N_47083,N_42567,N_44247);
nand U47084 (N_47084,N_44498,N_42581);
xnor U47085 (N_47085,N_40213,N_42477);
nand U47086 (N_47086,N_41741,N_40511);
or U47087 (N_47087,N_42752,N_40624);
and U47088 (N_47088,N_44936,N_43651);
nor U47089 (N_47089,N_40406,N_41446);
nand U47090 (N_47090,N_43462,N_42219);
nor U47091 (N_47091,N_42756,N_43147);
nand U47092 (N_47092,N_40044,N_43423);
nor U47093 (N_47093,N_40338,N_44091);
and U47094 (N_47094,N_40030,N_44981);
or U47095 (N_47095,N_42126,N_43836);
nand U47096 (N_47096,N_44354,N_41300);
nor U47097 (N_47097,N_41651,N_43688);
nand U47098 (N_47098,N_41120,N_40410);
nand U47099 (N_47099,N_42318,N_40299);
nand U47100 (N_47100,N_40753,N_41906);
nand U47101 (N_47101,N_42722,N_44800);
xor U47102 (N_47102,N_43833,N_42541);
or U47103 (N_47103,N_42153,N_44290);
nor U47104 (N_47104,N_42345,N_43066);
xor U47105 (N_47105,N_44035,N_41140);
or U47106 (N_47106,N_43482,N_41943);
and U47107 (N_47107,N_44411,N_42430);
or U47108 (N_47108,N_43202,N_43376);
xor U47109 (N_47109,N_41543,N_41489);
nor U47110 (N_47110,N_42490,N_40274);
xor U47111 (N_47111,N_43346,N_40659);
nor U47112 (N_47112,N_41174,N_42416);
and U47113 (N_47113,N_43572,N_41690);
and U47114 (N_47114,N_42820,N_43964);
xnor U47115 (N_47115,N_40026,N_41388);
or U47116 (N_47116,N_43704,N_43997);
nor U47117 (N_47117,N_41825,N_43819);
xor U47118 (N_47118,N_44163,N_42137);
nor U47119 (N_47119,N_42272,N_41419);
nor U47120 (N_47120,N_43144,N_40716);
nor U47121 (N_47121,N_43640,N_41905);
nor U47122 (N_47122,N_43538,N_44641);
nor U47123 (N_47123,N_42717,N_41699);
xnor U47124 (N_47124,N_44377,N_44601);
xor U47125 (N_47125,N_40296,N_44512);
nor U47126 (N_47126,N_44750,N_44011);
or U47127 (N_47127,N_43096,N_44743);
and U47128 (N_47128,N_40259,N_43433);
and U47129 (N_47129,N_40913,N_42786);
xnor U47130 (N_47130,N_44837,N_42925);
and U47131 (N_47131,N_40136,N_44448);
nor U47132 (N_47132,N_44141,N_41233);
or U47133 (N_47133,N_40638,N_40688);
or U47134 (N_47134,N_40833,N_44583);
nor U47135 (N_47135,N_40567,N_44716);
nand U47136 (N_47136,N_44898,N_40191);
nor U47137 (N_47137,N_43842,N_41139);
nor U47138 (N_47138,N_43550,N_44040);
and U47139 (N_47139,N_42816,N_40020);
and U47140 (N_47140,N_44008,N_44946);
xor U47141 (N_47141,N_42357,N_40837);
or U47142 (N_47142,N_42341,N_43309);
nor U47143 (N_47143,N_41392,N_42859);
or U47144 (N_47144,N_42336,N_40375);
xnor U47145 (N_47145,N_43310,N_43855);
or U47146 (N_47146,N_43890,N_44846);
nor U47147 (N_47147,N_40275,N_41946);
nor U47148 (N_47148,N_43869,N_43839);
or U47149 (N_47149,N_42328,N_43326);
xnor U47150 (N_47150,N_41241,N_43471);
nand U47151 (N_47151,N_42225,N_42806);
or U47152 (N_47152,N_44028,N_40037);
or U47153 (N_47153,N_44199,N_41444);
nor U47154 (N_47154,N_41464,N_42658);
nand U47155 (N_47155,N_42991,N_44368);
nor U47156 (N_47156,N_42076,N_44434);
and U47157 (N_47157,N_43077,N_41867);
xnor U47158 (N_47158,N_42287,N_40541);
or U47159 (N_47159,N_43446,N_41618);
and U47160 (N_47160,N_43983,N_40302);
or U47161 (N_47161,N_41262,N_42544);
xnor U47162 (N_47162,N_44712,N_44396);
nor U47163 (N_47163,N_44394,N_40134);
xnor U47164 (N_47164,N_41036,N_41744);
nand U47165 (N_47165,N_44876,N_44298);
or U47166 (N_47166,N_43816,N_40773);
nor U47167 (N_47167,N_44972,N_44161);
or U47168 (N_47168,N_42309,N_41657);
and U47169 (N_47169,N_44083,N_40797);
xor U47170 (N_47170,N_40770,N_41537);
or U47171 (N_47171,N_43333,N_44012);
or U47172 (N_47172,N_42003,N_42232);
and U47173 (N_47173,N_41634,N_42385);
xnor U47174 (N_47174,N_43360,N_40632);
nand U47175 (N_47175,N_43788,N_43293);
and U47176 (N_47176,N_44867,N_40184);
or U47177 (N_47177,N_40805,N_43197);
and U47178 (N_47178,N_41947,N_43531);
nand U47179 (N_47179,N_42052,N_43814);
nand U47180 (N_47180,N_42881,N_40364);
xnor U47181 (N_47181,N_44132,N_44207);
nand U47182 (N_47182,N_44728,N_42566);
and U47183 (N_47183,N_42255,N_41335);
or U47184 (N_47184,N_41832,N_43101);
xor U47185 (N_47185,N_43052,N_42480);
and U47186 (N_47186,N_42762,N_41893);
xnor U47187 (N_47187,N_41784,N_41454);
or U47188 (N_47188,N_44537,N_44061);
nor U47189 (N_47189,N_43429,N_44875);
and U47190 (N_47190,N_42555,N_40559);
or U47191 (N_47191,N_42520,N_43914);
xnor U47192 (N_47192,N_44097,N_42691);
and U47193 (N_47193,N_41502,N_41950);
and U47194 (N_47194,N_42829,N_44943);
and U47195 (N_47195,N_43271,N_42758);
xor U47196 (N_47196,N_41405,N_44897);
or U47197 (N_47197,N_40168,N_40326);
and U47198 (N_47198,N_43050,N_41903);
and U47199 (N_47199,N_41414,N_40783);
nand U47200 (N_47200,N_41421,N_41915);
nand U47201 (N_47201,N_44007,N_42600);
and U47202 (N_47202,N_41117,N_41108);
and U47203 (N_47203,N_42653,N_40475);
nor U47204 (N_47204,N_42979,N_41045);
or U47205 (N_47205,N_44758,N_40394);
xnor U47206 (N_47206,N_40795,N_43369);
or U47207 (N_47207,N_41282,N_41780);
xor U47208 (N_47208,N_43301,N_44799);
nand U47209 (N_47209,N_41628,N_41799);
nor U47210 (N_47210,N_41465,N_41914);
and U47211 (N_47211,N_42060,N_41868);
nand U47212 (N_47212,N_43746,N_41299);
xor U47213 (N_47213,N_42941,N_41172);
nor U47214 (N_47214,N_42432,N_42580);
nor U47215 (N_47215,N_43850,N_40786);
and U47216 (N_47216,N_40552,N_40127);
nand U47217 (N_47217,N_41578,N_42626);
or U47218 (N_47218,N_41572,N_44872);
nor U47219 (N_47219,N_43592,N_44102);
xnor U47220 (N_47220,N_40534,N_41093);
xor U47221 (N_47221,N_41245,N_41507);
xnor U47222 (N_47222,N_43159,N_44120);
or U47223 (N_47223,N_41062,N_40255);
and U47224 (N_47224,N_40745,N_41846);
nand U47225 (N_47225,N_44237,N_42887);
nand U47226 (N_47226,N_41083,N_43614);
nand U47227 (N_47227,N_42058,N_41034);
nand U47228 (N_47228,N_41263,N_40374);
and U47229 (N_47229,N_43418,N_43821);
xor U47230 (N_47230,N_43792,N_40281);
nor U47231 (N_47231,N_41691,N_43686);
nor U47232 (N_47232,N_40794,N_40498);
xor U47233 (N_47233,N_42731,N_44362);
or U47234 (N_47234,N_40677,N_40351);
xnor U47235 (N_47235,N_42377,N_43835);
nor U47236 (N_47236,N_44281,N_40389);
xnor U47237 (N_47237,N_44125,N_41167);
xnor U47238 (N_47238,N_41385,N_41659);
nor U47239 (N_47239,N_41668,N_44493);
or U47240 (N_47240,N_43111,N_43976);
or U47241 (N_47241,N_41410,N_43559);
or U47242 (N_47242,N_40808,N_43186);
nor U47243 (N_47243,N_40584,N_40265);
or U47244 (N_47244,N_40427,N_40390);
nor U47245 (N_47245,N_43330,N_41141);
or U47246 (N_47246,N_41296,N_43280);
xor U47247 (N_47247,N_40283,N_41560);
or U47248 (N_47248,N_42391,N_40472);
xor U47249 (N_47249,N_44835,N_43815);
xnor U47250 (N_47250,N_43010,N_41314);
and U47251 (N_47251,N_44249,N_41244);
nor U47252 (N_47252,N_41602,N_42587);
nand U47253 (N_47253,N_44533,N_40682);
or U47254 (N_47254,N_42179,N_42266);
and U47255 (N_47255,N_44462,N_41717);
xnor U47256 (N_47256,N_40545,N_43673);
and U47257 (N_47257,N_42306,N_44797);
and U47258 (N_47258,N_42870,N_42633);
and U47259 (N_47259,N_41207,N_40054);
or U47260 (N_47260,N_43085,N_44513);
nor U47261 (N_47261,N_44761,N_43882);
or U47262 (N_47262,N_41088,N_42116);
xnor U47263 (N_47263,N_41660,N_43472);
or U47264 (N_47264,N_40380,N_40899);
nand U47265 (N_47265,N_44296,N_43067);
xor U47266 (N_47266,N_42108,N_40442);
xor U47267 (N_47267,N_40423,N_40937);
xnor U47268 (N_47268,N_44052,N_40309);
xor U47269 (N_47269,N_43337,N_40721);
xor U47270 (N_47270,N_41667,N_43416);
and U47271 (N_47271,N_41955,N_44859);
or U47272 (N_47272,N_43414,N_41076);
nand U47273 (N_47273,N_41381,N_44766);
nand U47274 (N_47274,N_40854,N_41195);
xnor U47275 (N_47275,N_44311,N_43761);
xor U47276 (N_47276,N_42571,N_41800);
and U47277 (N_47277,N_42607,N_41919);
xor U47278 (N_47278,N_41689,N_40672);
or U47279 (N_47279,N_43465,N_44299);
xnor U47280 (N_47280,N_41519,N_42588);
xnor U47281 (N_47281,N_42209,N_40954);
nand U47282 (N_47282,N_40352,N_40361);
nor U47283 (N_47283,N_41163,N_42410);
nor U47284 (N_47284,N_43825,N_44682);
nor U47285 (N_47285,N_44351,N_40818);
nand U47286 (N_47286,N_42224,N_44369);
nor U47287 (N_47287,N_42858,N_42934);
nor U47288 (N_47288,N_40014,N_43596);
nor U47289 (N_47289,N_40839,N_44629);
or U47290 (N_47290,N_41791,N_42511);
nand U47291 (N_47291,N_42380,N_42895);
or U47292 (N_47292,N_42423,N_42523);
or U47293 (N_47293,N_44661,N_42450);
and U47294 (N_47294,N_44318,N_44101);
or U47295 (N_47295,N_42590,N_40206);
nor U47296 (N_47296,N_41942,N_43896);
nor U47297 (N_47297,N_42771,N_43569);
and U47298 (N_47298,N_41026,N_43406);
nand U47299 (N_47299,N_40634,N_44074);
or U47300 (N_47300,N_42665,N_44815);
xnor U47301 (N_47301,N_40855,N_40618);
or U47302 (N_47302,N_43362,N_43438);
xnor U47303 (N_47303,N_42545,N_42554);
and U47304 (N_47304,N_42343,N_44598);
xnor U47305 (N_47305,N_42268,N_43169);
nand U47306 (N_47306,N_40530,N_41622);
nand U47307 (N_47307,N_42228,N_40707);
and U47308 (N_47308,N_43299,N_44162);
or U47309 (N_47309,N_44297,N_40648);
and U47310 (N_47310,N_43295,N_41533);
and U47311 (N_47311,N_41056,N_41680);
and U47312 (N_47312,N_44021,N_44596);
or U47313 (N_47313,N_44631,N_44346);
xnor U47314 (N_47314,N_42553,N_40107);
xor U47315 (N_47315,N_40079,N_40557);
nor U47316 (N_47316,N_41332,N_42601);
nor U47317 (N_47317,N_43589,N_44292);
and U47318 (N_47318,N_42989,N_42973);
xor U47319 (N_47319,N_42346,N_42608);
xnor U47320 (N_47320,N_44655,N_40381);
nand U47321 (N_47321,N_42935,N_41178);
and U47322 (N_47322,N_40045,N_41920);
nor U47323 (N_47323,N_40396,N_44183);
or U47324 (N_47324,N_42181,N_42360);
and U47325 (N_47325,N_44702,N_40826);
nor U47326 (N_47326,N_42668,N_42499);
nand U47327 (N_47327,N_41775,N_40714);
nor U47328 (N_47328,N_43924,N_42202);
xnor U47329 (N_47329,N_44482,N_42730);
and U47330 (N_47330,N_44861,N_44438);
and U47331 (N_47331,N_42284,N_42586);
nand U47332 (N_47332,N_41992,N_43045);
nor U47333 (N_47333,N_41871,N_40223);
xor U47334 (N_47334,N_41295,N_43827);
or U47335 (N_47335,N_44544,N_41302);
nand U47336 (N_47336,N_40467,N_42479);
or U47337 (N_47337,N_42721,N_44206);
and U47338 (N_47338,N_44527,N_41312);
xor U47339 (N_47339,N_42335,N_44105);
xor U47340 (N_47340,N_43419,N_44133);
nor U47341 (N_47341,N_42724,N_41496);
nand U47342 (N_47342,N_41982,N_44517);
xor U47343 (N_47343,N_44287,N_43501);
nand U47344 (N_47344,N_40445,N_44560);
xnor U47345 (N_47345,N_41396,N_40170);
xnor U47346 (N_47346,N_40218,N_42578);
and U47347 (N_47347,N_40150,N_41605);
nand U47348 (N_47348,N_43420,N_41985);
xnor U47349 (N_47349,N_41530,N_40814);
or U47350 (N_47350,N_40303,N_40700);
nand U47351 (N_47351,N_43702,N_44440);
nor U47352 (N_47352,N_44444,N_43860);
nand U47353 (N_47353,N_44400,N_43504);
or U47354 (N_47354,N_42029,N_44976);
nand U47355 (N_47355,N_43034,N_42267);
nand U47356 (N_47356,N_43265,N_42154);
nand U47357 (N_47357,N_43669,N_42216);
nor U47358 (N_47358,N_43141,N_40729);
xor U47359 (N_47359,N_41522,N_40062);
nand U47360 (N_47360,N_40286,N_42667);
xnor U47361 (N_47361,N_43717,N_42735);
or U47362 (N_47362,N_41416,N_44481);
nand U47363 (N_47363,N_40796,N_43852);
nand U47364 (N_47364,N_43608,N_44968);
xor U47365 (N_47365,N_43266,N_42977);
and U47366 (N_47366,N_44614,N_42447);
and U47367 (N_47367,N_42217,N_40574);
nand U47368 (N_47368,N_43021,N_44914);
and U47369 (N_47369,N_42890,N_41814);
nand U47370 (N_47370,N_41840,N_43639);
nand U47371 (N_47371,N_41096,N_41999);
and U47372 (N_47372,N_40320,N_44042);
nor U47373 (N_47373,N_43740,N_43641);
nand U47374 (N_47374,N_42094,N_40105);
or U47375 (N_47375,N_41581,N_43629);
or U47376 (N_47376,N_41702,N_41482);
or U47377 (N_47377,N_41303,N_43579);
nand U47378 (N_47378,N_42073,N_43949);
or U47379 (N_47379,N_40578,N_41449);
xnor U47380 (N_47380,N_41002,N_41286);
xor U47381 (N_47381,N_41490,N_42901);
and U47382 (N_47382,N_42543,N_40752);
and U47383 (N_47383,N_44456,N_44370);
nand U47384 (N_47384,N_41594,N_41393);
and U47385 (N_47385,N_41913,N_41993);
nand U47386 (N_47386,N_42943,N_40115);
nor U47387 (N_47387,N_40874,N_41787);
or U47388 (N_47388,N_43279,N_41000);
or U47389 (N_47389,N_41291,N_41694);
and U47390 (N_47390,N_41270,N_44404);
or U47391 (N_47391,N_41341,N_40113);
xor U47392 (N_47392,N_42152,N_44991);
nand U47393 (N_47393,N_43395,N_44547);
or U47394 (N_47394,N_44130,N_40573);
nand U47395 (N_47395,N_40673,N_43227);
xnor U47396 (N_47396,N_40004,N_40328);
nand U47397 (N_47397,N_40041,N_44853);
xnor U47398 (N_47398,N_42604,N_42651);
xnor U47399 (N_47399,N_44328,N_43778);
xnor U47400 (N_47400,N_41839,N_42818);
or U47401 (N_47401,N_41866,N_44471);
nand U47402 (N_47402,N_44313,N_41132);
nand U47403 (N_47403,N_41345,N_44901);
nor U47404 (N_47404,N_43391,N_40488);
nor U47405 (N_47405,N_41305,N_40538);
nand U47406 (N_47406,N_42953,N_44062);
nand U47407 (N_47407,N_42734,N_43172);
nor U47408 (N_47408,N_43100,N_41151);
xnor U47409 (N_47409,N_44066,N_42319);
xnor U47410 (N_47410,N_44391,N_40589);
xnor U47411 (N_47411,N_44511,N_43981);
xor U47412 (N_47412,N_40268,N_40132);
and U47413 (N_47413,N_40008,N_42135);
and U47414 (N_47414,N_41445,N_44176);
and U47415 (N_47415,N_42474,N_41821);
and U47416 (N_47416,N_41510,N_44243);
nand U47417 (N_47417,N_42873,N_44240);
nand U47418 (N_47418,N_44727,N_44948);
nand U47419 (N_47419,N_44644,N_41842);
or U47420 (N_47420,N_41963,N_40995);
or U47421 (N_47421,N_41014,N_43950);
nor U47422 (N_47422,N_42597,N_43332);
and U47423 (N_47423,N_43307,N_40544);
xnor U47424 (N_47424,N_44782,N_44741);
or U47425 (N_47425,N_41952,N_42160);
nand U47426 (N_47426,N_43724,N_41467);
and U47427 (N_47427,N_41339,N_44140);
nand U47428 (N_47428,N_40974,N_41400);
and U47429 (N_47429,N_40359,N_44345);
or U47430 (N_47430,N_43417,N_42755);
xor U47431 (N_47431,N_40667,N_44387);
xnor U47432 (N_47432,N_41250,N_40091);
and U47433 (N_47433,N_44080,N_43219);
and U47434 (N_47434,N_40865,N_43104);
nor U47435 (N_47435,N_44860,N_40943);
nor U47436 (N_47436,N_42612,N_44550);
nor U47437 (N_47437,N_44715,N_44504);
nand U47438 (N_47438,N_41574,N_40492);
and U47439 (N_47439,N_42011,N_40446);
nor U47440 (N_47440,N_44615,N_40983);
xor U47441 (N_47441,N_42957,N_41978);
and U47442 (N_47442,N_44374,N_42506);
nor U47443 (N_47443,N_40058,N_40145);
nor U47444 (N_47444,N_43671,N_40316);
and U47445 (N_47445,N_44412,N_44131);
nor U47446 (N_47446,N_42839,N_44551);
xnor U47447 (N_47447,N_43494,N_42754);
xnor U47448 (N_47448,N_41458,N_42878);
and U47449 (N_47449,N_42516,N_42993);
xor U47450 (N_47450,N_44604,N_41678);
or U47451 (N_47451,N_42877,N_40979);
nor U47452 (N_47452,N_41211,N_43682);
nand U47453 (N_47453,N_40051,N_42868);
nand U47454 (N_47454,N_40650,N_41615);
nor U47455 (N_47455,N_42559,N_41921);
or U47456 (N_47456,N_44308,N_42636);
and U47457 (N_47457,N_44687,N_44862);
nand U47458 (N_47458,N_40636,N_40121);
or U47459 (N_47459,N_43364,N_42800);
nand U47460 (N_47460,N_41703,N_42892);
nor U47461 (N_47461,N_43849,N_43182);
and U47462 (N_47462,N_44271,N_43637);
nand U47463 (N_47463,N_43797,N_43958);
and U47464 (N_47464,N_41734,N_40169);
nor U47465 (N_47465,N_41501,N_40458);
nand U47466 (N_47466,N_42785,N_43032);
xnor U47467 (N_47467,N_43561,N_44306);
and U47468 (N_47468,N_42652,N_44895);
xor U47469 (N_47469,N_42299,N_44917);
nand U47470 (N_47470,N_42023,N_42254);
nor U47471 (N_47471,N_43744,N_41290);
xor U47472 (N_47472,N_44327,N_41938);
nor U47473 (N_47473,N_40332,N_43854);
and U47474 (N_47474,N_42408,N_42694);
nor U47475 (N_47475,N_42281,N_40129);
nor U47476 (N_47476,N_43158,N_41589);
nor U47477 (N_47477,N_44069,N_41518);
or U47478 (N_47478,N_43496,N_40761);
xor U47479 (N_47479,N_40454,N_43582);
xnor U47480 (N_47480,N_41255,N_41802);
and U47481 (N_47481,N_40906,N_43653);
and U47482 (N_47482,N_42363,N_40022);
and U47483 (N_47483,N_41826,N_42314);
or U47484 (N_47484,N_41213,N_43278);
and U47485 (N_47485,N_41042,N_41764);
xnor U47486 (N_47486,N_43459,N_41767);
or U47487 (N_47487,N_40600,N_43796);
nor U47488 (N_47488,N_40212,N_43883);
and U47489 (N_47489,N_44030,N_41350);
nor U47490 (N_47490,N_41773,N_42840);
and U47491 (N_47491,N_44380,N_41857);
nor U47492 (N_47492,N_43881,N_42401);
and U47493 (N_47493,N_41899,N_40308);
xnor U47494 (N_47494,N_40219,N_42700);
and U47495 (N_47495,N_41548,N_44001);
or U47496 (N_47496,N_40925,N_42418);
or U47497 (N_47497,N_41418,N_44154);
and U47498 (N_47498,N_43692,N_44927);
nand U47499 (N_47499,N_41370,N_43226);
nand U47500 (N_47500,N_43087,N_42640);
nor U47501 (N_47501,N_41747,N_44706);
nand U47502 (N_47502,N_40122,N_44324);
xor U47503 (N_47503,N_44555,N_42057);
nor U47504 (N_47504,N_44209,N_42840);
or U47505 (N_47505,N_43574,N_42200);
or U47506 (N_47506,N_42242,N_44745);
or U47507 (N_47507,N_41489,N_41930);
nor U47508 (N_47508,N_41943,N_43242);
and U47509 (N_47509,N_40199,N_42518);
xnor U47510 (N_47510,N_41374,N_43419);
nand U47511 (N_47511,N_40309,N_44447);
or U47512 (N_47512,N_40893,N_42205);
nor U47513 (N_47513,N_41173,N_43052);
nor U47514 (N_47514,N_42269,N_43530);
nor U47515 (N_47515,N_43367,N_42703);
and U47516 (N_47516,N_40359,N_40440);
nor U47517 (N_47517,N_41034,N_41860);
xnor U47518 (N_47518,N_44215,N_40420);
nor U47519 (N_47519,N_42242,N_42018);
and U47520 (N_47520,N_43165,N_41554);
nor U47521 (N_47521,N_43723,N_42137);
nand U47522 (N_47522,N_44673,N_43433);
nand U47523 (N_47523,N_41341,N_44552);
nor U47524 (N_47524,N_40043,N_41939);
or U47525 (N_47525,N_44473,N_44782);
nor U47526 (N_47526,N_44385,N_41289);
and U47527 (N_47527,N_41083,N_40331);
nand U47528 (N_47528,N_44231,N_44971);
nand U47529 (N_47529,N_43177,N_42470);
and U47530 (N_47530,N_44480,N_40674);
or U47531 (N_47531,N_44304,N_43851);
nor U47532 (N_47532,N_40004,N_42530);
nand U47533 (N_47533,N_41096,N_44246);
and U47534 (N_47534,N_43171,N_41949);
nor U47535 (N_47535,N_44884,N_43679);
xnor U47536 (N_47536,N_41580,N_40751);
or U47537 (N_47537,N_40581,N_42921);
nor U47538 (N_47538,N_41909,N_40271);
xnor U47539 (N_47539,N_43490,N_42910);
or U47540 (N_47540,N_44785,N_43851);
xor U47541 (N_47541,N_40705,N_40604);
or U47542 (N_47542,N_40634,N_41305);
or U47543 (N_47543,N_43273,N_43517);
nor U47544 (N_47544,N_43515,N_44510);
nor U47545 (N_47545,N_42226,N_40070);
nor U47546 (N_47546,N_40980,N_43420);
or U47547 (N_47547,N_40633,N_40047);
and U47548 (N_47548,N_42839,N_44753);
nor U47549 (N_47549,N_40982,N_44190);
nand U47550 (N_47550,N_44638,N_40454);
nor U47551 (N_47551,N_42740,N_40166);
and U47552 (N_47552,N_42251,N_42794);
xnor U47553 (N_47553,N_41201,N_44867);
and U47554 (N_47554,N_42739,N_42537);
nor U47555 (N_47555,N_44894,N_41081);
and U47556 (N_47556,N_42462,N_41671);
and U47557 (N_47557,N_42202,N_44727);
and U47558 (N_47558,N_41559,N_41245);
or U47559 (N_47559,N_41267,N_40892);
or U47560 (N_47560,N_43646,N_41266);
nand U47561 (N_47561,N_42063,N_40536);
or U47562 (N_47562,N_44243,N_40387);
or U47563 (N_47563,N_40838,N_44523);
nand U47564 (N_47564,N_44072,N_42006);
xor U47565 (N_47565,N_44758,N_41902);
xor U47566 (N_47566,N_42688,N_40243);
or U47567 (N_47567,N_41026,N_42249);
and U47568 (N_47568,N_40469,N_44036);
nor U47569 (N_47569,N_40726,N_44272);
or U47570 (N_47570,N_43789,N_44469);
nor U47571 (N_47571,N_43069,N_41557);
or U47572 (N_47572,N_40032,N_41854);
or U47573 (N_47573,N_40999,N_42358);
nand U47574 (N_47574,N_44788,N_42718);
nor U47575 (N_47575,N_43889,N_44970);
and U47576 (N_47576,N_44493,N_41367);
nor U47577 (N_47577,N_40319,N_41829);
nand U47578 (N_47578,N_40225,N_40233);
or U47579 (N_47579,N_41809,N_42071);
or U47580 (N_47580,N_40595,N_44848);
xnor U47581 (N_47581,N_41856,N_44092);
xor U47582 (N_47582,N_43028,N_42849);
and U47583 (N_47583,N_44820,N_40060);
and U47584 (N_47584,N_40461,N_40656);
xor U47585 (N_47585,N_41275,N_44795);
or U47586 (N_47586,N_40772,N_41523);
and U47587 (N_47587,N_41721,N_42990);
and U47588 (N_47588,N_41896,N_40079);
nand U47589 (N_47589,N_42792,N_44918);
and U47590 (N_47590,N_44638,N_44344);
or U47591 (N_47591,N_43962,N_41834);
nor U47592 (N_47592,N_42957,N_44220);
nor U47593 (N_47593,N_44138,N_42579);
nand U47594 (N_47594,N_41721,N_42348);
xnor U47595 (N_47595,N_43879,N_44648);
nand U47596 (N_47596,N_40604,N_40492);
nand U47597 (N_47597,N_42387,N_41675);
or U47598 (N_47598,N_43258,N_42324);
nor U47599 (N_47599,N_42488,N_42019);
nor U47600 (N_47600,N_43017,N_44588);
nand U47601 (N_47601,N_42489,N_42662);
and U47602 (N_47602,N_41210,N_40737);
xnor U47603 (N_47603,N_44378,N_41608);
nor U47604 (N_47604,N_42180,N_40164);
nor U47605 (N_47605,N_44064,N_41135);
or U47606 (N_47606,N_42860,N_42524);
nor U47607 (N_47607,N_40522,N_43153);
nor U47608 (N_47608,N_42283,N_43994);
xnor U47609 (N_47609,N_41246,N_43559);
nor U47610 (N_47610,N_42043,N_43415);
and U47611 (N_47611,N_43405,N_41915);
nor U47612 (N_47612,N_43481,N_43790);
and U47613 (N_47613,N_41189,N_43506);
nor U47614 (N_47614,N_41559,N_40639);
or U47615 (N_47615,N_44577,N_41806);
and U47616 (N_47616,N_41816,N_44739);
nor U47617 (N_47617,N_40775,N_40164);
and U47618 (N_47618,N_43704,N_44074);
xor U47619 (N_47619,N_40738,N_43003);
nand U47620 (N_47620,N_40147,N_41883);
nor U47621 (N_47621,N_44165,N_43440);
nand U47622 (N_47622,N_41956,N_41766);
nand U47623 (N_47623,N_42399,N_40582);
nand U47624 (N_47624,N_42533,N_44425);
and U47625 (N_47625,N_41782,N_40996);
nor U47626 (N_47626,N_43164,N_44442);
nand U47627 (N_47627,N_44166,N_42193);
or U47628 (N_47628,N_42253,N_41332);
nor U47629 (N_47629,N_44280,N_40837);
nand U47630 (N_47630,N_44108,N_41405);
xnor U47631 (N_47631,N_43949,N_40457);
and U47632 (N_47632,N_44709,N_40038);
nand U47633 (N_47633,N_44451,N_41979);
and U47634 (N_47634,N_42749,N_40292);
nor U47635 (N_47635,N_44427,N_40176);
or U47636 (N_47636,N_42678,N_42955);
or U47637 (N_47637,N_40619,N_43791);
and U47638 (N_47638,N_42712,N_43736);
xor U47639 (N_47639,N_40484,N_40876);
nor U47640 (N_47640,N_41893,N_40696);
and U47641 (N_47641,N_43664,N_40923);
and U47642 (N_47642,N_41275,N_40052);
nor U47643 (N_47643,N_41608,N_42307);
nand U47644 (N_47644,N_44358,N_41189);
nor U47645 (N_47645,N_40424,N_43471);
nor U47646 (N_47646,N_44162,N_41275);
or U47647 (N_47647,N_42153,N_41090);
nor U47648 (N_47648,N_40917,N_43765);
nor U47649 (N_47649,N_42990,N_43131);
xnor U47650 (N_47650,N_42801,N_43788);
xor U47651 (N_47651,N_43474,N_42003);
xor U47652 (N_47652,N_44106,N_40989);
or U47653 (N_47653,N_43886,N_40072);
nand U47654 (N_47654,N_44111,N_44809);
nor U47655 (N_47655,N_41548,N_44498);
xor U47656 (N_47656,N_40021,N_43447);
or U47657 (N_47657,N_41370,N_41319);
nor U47658 (N_47658,N_42790,N_44519);
nand U47659 (N_47659,N_41022,N_41820);
nand U47660 (N_47660,N_40499,N_43211);
and U47661 (N_47661,N_44111,N_40130);
nor U47662 (N_47662,N_44466,N_41395);
nor U47663 (N_47663,N_43093,N_42533);
nor U47664 (N_47664,N_44301,N_41703);
nand U47665 (N_47665,N_42360,N_44723);
and U47666 (N_47666,N_43773,N_43309);
nand U47667 (N_47667,N_40549,N_41655);
or U47668 (N_47668,N_44744,N_41991);
nor U47669 (N_47669,N_40193,N_41090);
or U47670 (N_47670,N_42368,N_42098);
nand U47671 (N_47671,N_42003,N_43676);
or U47672 (N_47672,N_42014,N_40227);
or U47673 (N_47673,N_44792,N_42641);
nand U47674 (N_47674,N_40848,N_41704);
or U47675 (N_47675,N_41821,N_44390);
and U47676 (N_47676,N_40444,N_42387);
nand U47677 (N_47677,N_44904,N_40544);
or U47678 (N_47678,N_42105,N_40245);
nor U47679 (N_47679,N_42070,N_43607);
or U47680 (N_47680,N_42901,N_44097);
and U47681 (N_47681,N_41247,N_44770);
and U47682 (N_47682,N_42657,N_41795);
nand U47683 (N_47683,N_43820,N_44167);
xor U47684 (N_47684,N_44117,N_42012);
nor U47685 (N_47685,N_41063,N_41826);
or U47686 (N_47686,N_43431,N_43598);
and U47687 (N_47687,N_42875,N_43889);
or U47688 (N_47688,N_40972,N_42461);
nand U47689 (N_47689,N_42337,N_43784);
or U47690 (N_47690,N_44915,N_40094);
nand U47691 (N_47691,N_44940,N_44058);
and U47692 (N_47692,N_43507,N_41363);
or U47693 (N_47693,N_40497,N_43194);
xnor U47694 (N_47694,N_42685,N_43342);
and U47695 (N_47695,N_44416,N_41873);
and U47696 (N_47696,N_44305,N_41076);
or U47697 (N_47697,N_40853,N_44637);
nand U47698 (N_47698,N_41069,N_41996);
nand U47699 (N_47699,N_43338,N_41027);
nand U47700 (N_47700,N_42767,N_44965);
nor U47701 (N_47701,N_44556,N_43450);
or U47702 (N_47702,N_42965,N_43599);
or U47703 (N_47703,N_44535,N_43390);
nor U47704 (N_47704,N_43374,N_40553);
and U47705 (N_47705,N_40188,N_44937);
or U47706 (N_47706,N_43796,N_44133);
xnor U47707 (N_47707,N_40849,N_40208);
and U47708 (N_47708,N_44513,N_42475);
nand U47709 (N_47709,N_41879,N_41903);
or U47710 (N_47710,N_43311,N_41515);
nand U47711 (N_47711,N_43221,N_43991);
or U47712 (N_47712,N_41724,N_44495);
xnor U47713 (N_47713,N_43084,N_44064);
nor U47714 (N_47714,N_43585,N_43285);
nor U47715 (N_47715,N_42688,N_41287);
nand U47716 (N_47716,N_42934,N_41787);
nand U47717 (N_47717,N_43226,N_44798);
nor U47718 (N_47718,N_43379,N_40908);
nor U47719 (N_47719,N_42636,N_40944);
nand U47720 (N_47720,N_40103,N_44842);
nor U47721 (N_47721,N_41133,N_43199);
or U47722 (N_47722,N_41295,N_40309);
xor U47723 (N_47723,N_40097,N_40518);
and U47724 (N_47724,N_43368,N_43556);
nand U47725 (N_47725,N_43074,N_41384);
nand U47726 (N_47726,N_44686,N_43414);
nor U47727 (N_47727,N_41669,N_40338);
nand U47728 (N_47728,N_40305,N_44300);
xnor U47729 (N_47729,N_44308,N_41828);
nor U47730 (N_47730,N_42833,N_44478);
xor U47731 (N_47731,N_43731,N_43981);
and U47732 (N_47732,N_43291,N_40379);
and U47733 (N_47733,N_43316,N_44174);
xor U47734 (N_47734,N_42411,N_41360);
nor U47735 (N_47735,N_43646,N_42637);
nand U47736 (N_47736,N_44396,N_44836);
and U47737 (N_47737,N_44631,N_44344);
and U47738 (N_47738,N_44097,N_42308);
xor U47739 (N_47739,N_44631,N_44544);
or U47740 (N_47740,N_40166,N_42635);
or U47741 (N_47741,N_42254,N_40480);
nor U47742 (N_47742,N_40455,N_41790);
and U47743 (N_47743,N_42799,N_41751);
nand U47744 (N_47744,N_41630,N_41926);
xnor U47745 (N_47745,N_41072,N_41486);
nand U47746 (N_47746,N_40849,N_44188);
nor U47747 (N_47747,N_42765,N_40897);
and U47748 (N_47748,N_42137,N_44760);
xnor U47749 (N_47749,N_41300,N_44785);
nor U47750 (N_47750,N_44283,N_43291);
and U47751 (N_47751,N_40444,N_42072);
and U47752 (N_47752,N_42796,N_40933);
and U47753 (N_47753,N_44410,N_40021);
xnor U47754 (N_47754,N_41744,N_43979);
nor U47755 (N_47755,N_44375,N_42427);
and U47756 (N_47756,N_44122,N_42206);
and U47757 (N_47757,N_41155,N_40694);
nor U47758 (N_47758,N_40209,N_41970);
or U47759 (N_47759,N_40160,N_43284);
nand U47760 (N_47760,N_43763,N_44811);
xor U47761 (N_47761,N_44674,N_44044);
nor U47762 (N_47762,N_40664,N_41852);
nor U47763 (N_47763,N_44386,N_40213);
xor U47764 (N_47764,N_40335,N_40956);
and U47765 (N_47765,N_43846,N_42452);
nor U47766 (N_47766,N_42642,N_41024);
xnor U47767 (N_47767,N_43670,N_40224);
nor U47768 (N_47768,N_41444,N_41880);
nand U47769 (N_47769,N_43148,N_44837);
and U47770 (N_47770,N_40067,N_44837);
nor U47771 (N_47771,N_42514,N_44089);
nor U47772 (N_47772,N_41889,N_40342);
nand U47773 (N_47773,N_40581,N_44497);
nor U47774 (N_47774,N_41659,N_43159);
or U47775 (N_47775,N_40233,N_40530);
xor U47776 (N_47776,N_41575,N_41879);
or U47777 (N_47777,N_44466,N_41362);
or U47778 (N_47778,N_44933,N_42399);
nor U47779 (N_47779,N_44755,N_41255);
nand U47780 (N_47780,N_43061,N_43294);
nand U47781 (N_47781,N_42053,N_41009);
or U47782 (N_47782,N_43246,N_43761);
xor U47783 (N_47783,N_44344,N_40775);
or U47784 (N_47784,N_42205,N_40080);
or U47785 (N_47785,N_43657,N_40356);
and U47786 (N_47786,N_43120,N_43632);
or U47787 (N_47787,N_42181,N_41065);
or U47788 (N_47788,N_43433,N_43159);
xor U47789 (N_47789,N_40585,N_44381);
and U47790 (N_47790,N_43390,N_42482);
nand U47791 (N_47791,N_42086,N_43669);
nand U47792 (N_47792,N_44347,N_40443);
nand U47793 (N_47793,N_44961,N_41383);
or U47794 (N_47794,N_43295,N_44141);
xnor U47795 (N_47795,N_40253,N_41034);
nand U47796 (N_47796,N_40586,N_44509);
xor U47797 (N_47797,N_43979,N_41225);
nor U47798 (N_47798,N_44568,N_41823);
xor U47799 (N_47799,N_43212,N_43192);
nor U47800 (N_47800,N_43340,N_43931);
nand U47801 (N_47801,N_41432,N_44557);
xor U47802 (N_47802,N_40308,N_41905);
nor U47803 (N_47803,N_41163,N_40755);
nand U47804 (N_47804,N_44196,N_41065);
nor U47805 (N_47805,N_44011,N_42401);
or U47806 (N_47806,N_41952,N_40352);
xnor U47807 (N_47807,N_41499,N_41937);
and U47808 (N_47808,N_41397,N_44704);
xnor U47809 (N_47809,N_40660,N_43407);
xor U47810 (N_47810,N_43478,N_44931);
nor U47811 (N_47811,N_42462,N_44688);
xnor U47812 (N_47812,N_41301,N_43412);
and U47813 (N_47813,N_43861,N_44979);
and U47814 (N_47814,N_42512,N_41083);
nand U47815 (N_47815,N_43479,N_42231);
nor U47816 (N_47816,N_44620,N_42247);
or U47817 (N_47817,N_44546,N_43751);
nor U47818 (N_47818,N_44134,N_44216);
nand U47819 (N_47819,N_41215,N_43432);
and U47820 (N_47820,N_44790,N_40472);
xor U47821 (N_47821,N_41198,N_41775);
nor U47822 (N_47822,N_43898,N_40824);
or U47823 (N_47823,N_42777,N_42921);
nor U47824 (N_47824,N_41033,N_40954);
nand U47825 (N_47825,N_41807,N_40040);
nor U47826 (N_47826,N_43303,N_43551);
nand U47827 (N_47827,N_43077,N_43260);
nor U47828 (N_47828,N_42463,N_43633);
and U47829 (N_47829,N_41440,N_40262);
xor U47830 (N_47830,N_42039,N_41498);
xor U47831 (N_47831,N_41646,N_40590);
nand U47832 (N_47832,N_42425,N_41639);
and U47833 (N_47833,N_40080,N_42695);
nor U47834 (N_47834,N_43774,N_44681);
or U47835 (N_47835,N_44366,N_44850);
nand U47836 (N_47836,N_40826,N_40529);
and U47837 (N_47837,N_43689,N_41469);
or U47838 (N_47838,N_42004,N_40702);
nand U47839 (N_47839,N_43551,N_41218);
and U47840 (N_47840,N_42430,N_42476);
nor U47841 (N_47841,N_41260,N_40776);
and U47842 (N_47842,N_44682,N_44870);
nor U47843 (N_47843,N_43872,N_43383);
or U47844 (N_47844,N_41919,N_42482);
or U47845 (N_47845,N_41676,N_43407);
nand U47846 (N_47846,N_42936,N_44802);
and U47847 (N_47847,N_41667,N_44615);
and U47848 (N_47848,N_42575,N_43199);
xnor U47849 (N_47849,N_41620,N_40738);
nor U47850 (N_47850,N_42903,N_43644);
or U47851 (N_47851,N_44858,N_43357);
nor U47852 (N_47852,N_44384,N_41988);
or U47853 (N_47853,N_44322,N_41008);
or U47854 (N_47854,N_43781,N_40362);
and U47855 (N_47855,N_41352,N_42812);
or U47856 (N_47856,N_40989,N_40178);
or U47857 (N_47857,N_44516,N_42835);
nor U47858 (N_47858,N_40275,N_43725);
nor U47859 (N_47859,N_41396,N_41057);
nor U47860 (N_47860,N_41828,N_43207);
and U47861 (N_47861,N_44256,N_41003);
nor U47862 (N_47862,N_44420,N_40890);
nor U47863 (N_47863,N_41963,N_43755);
and U47864 (N_47864,N_43335,N_43884);
nand U47865 (N_47865,N_42665,N_43509);
xnor U47866 (N_47866,N_40864,N_43847);
nor U47867 (N_47867,N_44213,N_44233);
or U47868 (N_47868,N_40898,N_41601);
and U47869 (N_47869,N_40252,N_43864);
nand U47870 (N_47870,N_41306,N_43092);
and U47871 (N_47871,N_40833,N_43576);
and U47872 (N_47872,N_41428,N_41944);
xor U47873 (N_47873,N_43331,N_40544);
and U47874 (N_47874,N_44325,N_40672);
nor U47875 (N_47875,N_44410,N_40593);
nand U47876 (N_47876,N_43531,N_44165);
and U47877 (N_47877,N_44528,N_43481);
and U47878 (N_47878,N_43155,N_42402);
nor U47879 (N_47879,N_43196,N_43216);
or U47880 (N_47880,N_40946,N_41148);
nand U47881 (N_47881,N_43920,N_42276);
xnor U47882 (N_47882,N_44014,N_40975);
nand U47883 (N_47883,N_44540,N_40568);
or U47884 (N_47884,N_43263,N_41510);
nor U47885 (N_47885,N_41668,N_44137);
nor U47886 (N_47886,N_44447,N_41727);
or U47887 (N_47887,N_42685,N_44804);
nand U47888 (N_47888,N_41324,N_43156);
xnor U47889 (N_47889,N_43352,N_43949);
nor U47890 (N_47890,N_41249,N_41150);
or U47891 (N_47891,N_42981,N_43450);
nand U47892 (N_47892,N_44812,N_41310);
and U47893 (N_47893,N_41071,N_42475);
or U47894 (N_47894,N_43431,N_44408);
nand U47895 (N_47895,N_42013,N_43900);
xnor U47896 (N_47896,N_42352,N_44160);
nand U47897 (N_47897,N_41130,N_41439);
nand U47898 (N_47898,N_40783,N_43574);
xnor U47899 (N_47899,N_42429,N_44064);
nor U47900 (N_47900,N_40791,N_40905);
xor U47901 (N_47901,N_40123,N_44644);
nor U47902 (N_47902,N_41621,N_43039);
nand U47903 (N_47903,N_40507,N_43104);
nand U47904 (N_47904,N_44877,N_42517);
or U47905 (N_47905,N_44979,N_43204);
or U47906 (N_47906,N_43663,N_41413);
xnor U47907 (N_47907,N_43454,N_40550);
nand U47908 (N_47908,N_40994,N_40447);
xor U47909 (N_47909,N_43515,N_44703);
nand U47910 (N_47910,N_44699,N_43126);
or U47911 (N_47911,N_42788,N_42066);
and U47912 (N_47912,N_44601,N_44027);
nand U47913 (N_47913,N_44049,N_41683);
nand U47914 (N_47914,N_41194,N_44026);
or U47915 (N_47915,N_44148,N_43120);
nor U47916 (N_47916,N_44753,N_41712);
nor U47917 (N_47917,N_40459,N_41935);
and U47918 (N_47918,N_44968,N_42777);
nand U47919 (N_47919,N_43053,N_43932);
nand U47920 (N_47920,N_40430,N_40684);
or U47921 (N_47921,N_44070,N_42264);
or U47922 (N_47922,N_42958,N_41316);
xnor U47923 (N_47923,N_41732,N_41011);
and U47924 (N_47924,N_41438,N_44923);
nand U47925 (N_47925,N_43106,N_44821);
xnor U47926 (N_47926,N_44041,N_41157);
xnor U47927 (N_47927,N_42513,N_43472);
nand U47928 (N_47928,N_43069,N_41128);
and U47929 (N_47929,N_43745,N_44292);
xnor U47930 (N_47930,N_42938,N_41575);
or U47931 (N_47931,N_42399,N_41176);
nor U47932 (N_47932,N_42727,N_41372);
nand U47933 (N_47933,N_40213,N_41957);
xor U47934 (N_47934,N_40296,N_42980);
nor U47935 (N_47935,N_43166,N_40720);
nor U47936 (N_47936,N_42648,N_41113);
nor U47937 (N_47937,N_43610,N_42815);
nand U47938 (N_47938,N_43389,N_41181);
xnor U47939 (N_47939,N_41009,N_44120);
or U47940 (N_47940,N_43299,N_40434);
nand U47941 (N_47941,N_41402,N_40019);
xnor U47942 (N_47942,N_44121,N_43774);
or U47943 (N_47943,N_43237,N_42907);
or U47944 (N_47944,N_41192,N_40560);
nand U47945 (N_47945,N_41849,N_40796);
nor U47946 (N_47946,N_41903,N_41230);
nor U47947 (N_47947,N_42695,N_40669);
and U47948 (N_47948,N_42750,N_42310);
xor U47949 (N_47949,N_40219,N_42846);
nor U47950 (N_47950,N_40559,N_44012);
and U47951 (N_47951,N_41795,N_43422);
or U47952 (N_47952,N_42052,N_43331);
xnor U47953 (N_47953,N_44053,N_41496);
nor U47954 (N_47954,N_41139,N_41894);
nand U47955 (N_47955,N_42287,N_43637);
xnor U47956 (N_47956,N_40959,N_44084);
and U47957 (N_47957,N_41492,N_44412);
nor U47958 (N_47958,N_41415,N_40088);
and U47959 (N_47959,N_40237,N_41088);
or U47960 (N_47960,N_40151,N_40351);
xor U47961 (N_47961,N_44708,N_44904);
or U47962 (N_47962,N_43447,N_44480);
nand U47963 (N_47963,N_42599,N_43407);
and U47964 (N_47964,N_44738,N_44673);
xor U47965 (N_47965,N_42478,N_41824);
nand U47966 (N_47966,N_41828,N_43518);
or U47967 (N_47967,N_43333,N_41934);
xor U47968 (N_47968,N_41634,N_43549);
nand U47969 (N_47969,N_44520,N_41198);
or U47970 (N_47970,N_44414,N_42582);
or U47971 (N_47971,N_44216,N_43364);
nor U47972 (N_47972,N_43477,N_44499);
nor U47973 (N_47973,N_44619,N_42295);
xnor U47974 (N_47974,N_42841,N_44523);
nor U47975 (N_47975,N_41598,N_42185);
nand U47976 (N_47976,N_42212,N_44389);
or U47977 (N_47977,N_44193,N_42643);
or U47978 (N_47978,N_43651,N_44295);
nor U47979 (N_47979,N_41376,N_43590);
nor U47980 (N_47980,N_40103,N_43524);
or U47981 (N_47981,N_42304,N_41781);
or U47982 (N_47982,N_40276,N_44417);
nand U47983 (N_47983,N_41103,N_40826);
nand U47984 (N_47984,N_40769,N_44726);
xor U47985 (N_47985,N_43268,N_41935);
xor U47986 (N_47986,N_41907,N_44683);
nor U47987 (N_47987,N_40993,N_40754);
nor U47988 (N_47988,N_43778,N_43434);
or U47989 (N_47989,N_43798,N_43768);
and U47990 (N_47990,N_42894,N_43767);
or U47991 (N_47991,N_41644,N_44077);
xor U47992 (N_47992,N_40085,N_44270);
nand U47993 (N_47993,N_43981,N_41668);
or U47994 (N_47994,N_43856,N_42433);
nor U47995 (N_47995,N_40243,N_42997);
xor U47996 (N_47996,N_41242,N_43965);
xor U47997 (N_47997,N_41319,N_42682);
and U47998 (N_47998,N_42516,N_42379);
nor U47999 (N_47999,N_43752,N_42108);
and U48000 (N_48000,N_41945,N_41802);
and U48001 (N_48001,N_41167,N_42653);
or U48002 (N_48002,N_40619,N_44623);
nor U48003 (N_48003,N_43668,N_41111);
or U48004 (N_48004,N_41960,N_40621);
nor U48005 (N_48005,N_42085,N_43425);
or U48006 (N_48006,N_40154,N_44366);
or U48007 (N_48007,N_40164,N_44123);
or U48008 (N_48008,N_43570,N_43755);
nor U48009 (N_48009,N_41151,N_42941);
nand U48010 (N_48010,N_44474,N_43100);
nand U48011 (N_48011,N_41706,N_42443);
xnor U48012 (N_48012,N_42456,N_43789);
nor U48013 (N_48013,N_43184,N_41342);
nor U48014 (N_48014,N_44525,N_43821);
nor U48015 (N_48015,N_40902,N_43446);
nand U48016 (N_48016,N_43850,N_41681);
nand U48017 (N_48017,N_44515,N_43961);
or U48018 (N_48018,N_41239,N_42171);
nand U48019 (N_48019,N_40924,N_43709);
and U48020 (N_48020,N_41818,N_40610);
nor U48021 (N_48021,N_42081,N_42166);
and U48022 (N_48022,N_43912,N_43318);
and U48023 (N_48023,N_43189,N_41926);
nor U48024 (N_48024,N_43826,N_40857);
or U48025 (N_48025,N_43429,N_43783);
xnor U48026 (N_48026,N_40551,N_44690);
and U48027 (N_48027,N_43440,N_41386);
xor U48028 (N_48028,N_42803,N_44093);
xnor U48029 (N_48029,N_41484,N_41012);
and U48030 (N_48030,N_40171,N_44409);
or U48031 (N_48031,N_44349,N_44807);
xnor U48032 (N_48032,N_40645,N_42974);
xor U48033 (N_48033,N_41076,N_40881);
and U48034 (N_48034,N_40952,N_41157);
xor U48035 (N_48035,N_42327,N_41059);
xor U48036 (N_48036,N_42351,N_43453);
or U48037 (N_48037,N_40056,N_40667);
and U48038 (N_48038,N_44430,N_40508);
or U48039 (N_48039,N_41263,N_40782);
nand U48040 (N_48040,N_44050,N_40097);
and U48041 (N_48041,N_42942,N_41860);
xor U48042 (N_48042,N_43525,N_41783);
or U48043 (N_48043,N_44830,N_40236);
nor U48044 (N_48044,N_42014,N_42267);
or U48045 (N_48045,N_40081,N_42832);
and U48046 (N_48046,N_40860,N_44118);
nand U48047 (N_48047,N_44046,N_40763);
xnor U48048 (N_48048,N_40845,N_44074);
and U48049 (N_48049,N_43805,N_42321);
and U48050 (N_48050,N_41513,N_44300);
and U48051 (N_48051,N_43299,N_40488);
nand U48052 (N_48052,N_43225,N_40586);
nor U48053 (N_48053,N_42703,N_41040);
nand U48054 (N_48054,N_44351,N_40309);
and U48055 (N_48055,N_43353,N_40479);
nand U48056 (N_48056,N_44635,N_41834);
nor U48057 (N_48057,N_42656,N_42357);
nor U48058 (N_48058,N_40342,N_43333);
and U48059 (N_48059,N_40790,N_43537);
and U48060 (N_48060,N_41073,N_42022);
and U48061 (N_48061,N_41388,N_41696);
nand U48062 (N_48062,N_42010,N_40036);
nor U48063 (N_48063,N_40248,N_42783);
xnor U48064 (N_48064,N_44373,N_41373);
or U48065 (N_48065,N_44879,N_40657);
or U48066 (N_48066,N_44938,N_41827);
or U48067 (N_48067,N_43058,N_44293);
and U48068 (N_48068,N_42783,N_43681);
or U48069 (N_48069,N_41508,N_44076);
nand U48070 (N_48070,N_43936,N_42746);
and U48071 (N_48071,N_43926,N_43057);
xor U48072 (N_48072,N_44258,N_42518);
nor U48073 (N_48073,N_42854,N_40931);
and U48074 (N_48074,N_40606,N_41689);
nand U48075 (N_48075,N_44490,N_40078);
and U48076 (N_48076,N_43619,N_43758);
and U48077 (N_48077,N_43758,N_41231);
or U48078 (N_48078,N_44288,N_40621);
nor U48079 (N_48079,N_41446,N_44848);
nor U48080 (N_48080,N_41989,N_40846);
nand U48081 (N_48081,N_42436,N_44395);
or U48082 (N_48082,N_40351,N_40529);
nand U48083 (N_48083,N_42942,N_43955);
or U48084 (N_48084,N_42291,N_42003);
nor U48085 (N_48085,N_41728,N_44358);
or U48086 (N_48086,N_42337,N_41722);
or U48087 (N_48087,N_43292,N_41118);
nor U48088 (N_48088,N_41425,N_41796);
nand U48089 (N_48089,N_44501,N_43217);
or U48090 (N_48090,N_44424,N_42593);
xor U48091 (N_48091,N_41048,N_42734);
nand U48092 (N_48092,N_41391,N_43080);
and U48093 (N_48093,N_43797,N_41957);
xor U48094 (N_48094,N_43439,N_44087);
and U48095 (N_48095,N_41032,N_40708);
nand U48096 (N_48096,N_42363,N_40850);
nand U48097 (N_48097,N_42422,N_40792);
xnor U48098 (N_48098,N_44861,N_40934);
or U48099 (N_48099,N_42799,N_44130);
or U48100 (N_48100,N_41668,N_43270);
nor U48101 (N_48101,N_43972,N_41609);
nor U48102 (N_48102,N_43578,N_42890);
nand U48103 (N_48103,N_43352,N_43691);
nand U48104 (N_48104,N_40950,N_41562);
or U48105 (N_48105,N_41864,N_41509);
nand U48106 (N_48106,N_40053,N_41112);
nor U48107 (N_48107,N_43506,N_41797);
or U48108 (N_48108,N_44331,N_40157);
xnor U48109 (N_48109,N_42840,N_43183);
or U48110 (N_48110,N_40815,N_44116);
and U48111 (N_48111,N_44282,N_40280);
xor U48112 (N_48112,N_42767,N_42272);
or U48113 (N_48113,N_42727,N_44900);
or U48114 (N_48114,N_42222,N_41250);
nor U48115 (N_48115,N_43680,N_41058);
xor U48116 (N_48116,N_41005,N_40454);
and U48117 (N_48117,N_40071,N_43164);
and U48118 (N_48118,N_42603,N_44453);
xnor U48119 (N_48119,N_43796,N_42849);
xor U48120 (N_48120,N_40157,N_44596);
or U48121 (N_48121,N_42922,N_43316);
and U48122 (N_48122,N_44179,N_41061);
xnor U48123 (N_48123,N_43437,N_43430);
nor U48124 (N_48124,N_40788,N_44694);
and U48125 (N_48125,N_44700,N_42643);
and U48126 (N_48126,N_42403,N_40739);
nor U48127 (N_48127,N_41889,N_40301);
or U48128 (N_48128,N_44776,N_41713);
nor U48129 (N_48129,N_43241,N_44003);
and U48130 (N_48130,N_42429,N_44210);
nand U48131 (N_48131,N_44491,N_43692);
nor U48132 (N_48132,N_42574,N_40566);
nor U48133 (N_48133,N_44671,N_41063);
and U48134 (N_48134,N_42717,N_40470);
nand U48135 (N_48135,N_40108,N_44268);
nor U48136 (N_48136,N_43749,N_43707);
nand U48137 (N_48137,N_41676,N_40832);
and U48138 (N_48138,N_43397,N_44570);
nor U48139 (N_48139,N_41639,N_43720);
and U48140 (N_48140,N_40643,N_42074);
and U48141 (N_48141,N_43278,N_44247);
or U48142 (N_48142,N_41247,N_44872);
nand U48143 (N_48143,N_40641,N_43347);
nand U48144 (N_48144,N_40558,N_40744);
nor U48145 (N_48145,N_42802,N_40870);
nor U48146 (N_48146,N_42799,N_40103);
nor U48147 (N_48147,N_44698,N_42439);
nor U48148 (N_48148,N_42297,N_40689);
xnor U48149 (N_48149,N_41587,N_44087);
or U48150 (N_48150,N_44328,N_42986);
and U48151 (N_48151,N_41214,N_44972);
nand U48152 (N_48152,N_41165,N_44878);
nor U48153 (N_48153,N_40392,N_40703);
or U48154 (N_48154,N_40683,N_42263);
xnor U48155 (N_48155,N_41200,N_43554);
nor U48156 (N_48156,N_42007,N_41219);
xnor U48157 (N_48157,N_40634,N_43296);
xor U48158 (N_48158,N_43892,N_43108);
nor U48159 (N_48159,N_42808,N_42292);
nand U48160 (N_48160,N_40354,N_40448);
nand U48161 (N_48161,N_43407,N_42798);
and U48162 (N_48162,N_43140,N_40423);
xnor U48163 (N_48163,N_43927,N_42150);
xor U48164 (N_48164,N_43818,N_42026);
nor U48165 (N_48165,N_44119,N_44392);
xnor U48166 (N_48166,N_44147,N_44895);
or U48167 (N_48167,N_42863,N_42915);
or U48168 (N_48168,N_40338,N_43065);
nand U48169 (N_48169,N_41695,N_41197);
nand U48170 (N_48170,N_41891,N_44510);
xor U48171 (N_48171,N_41378,N_44860);
xor U48172 (N_48172,N_44941,N_43026);
nand U48173 (N_48173,N_42778,N_40160);
or U48174 (N_48174,N_44041,N_44104);
and U48175 (N_48175,N_43977,N_41233);
and U48176 (N_48176,N_40663,N_41933);
and U48177 (N_48177,N_40703,N_44058);
nand U48178 (N_48178,N_41300,N_42910);
xor U48179 (N_48179,N_43894,N_43343);
and U48180 (N_48180,N_43055,N_42774);
xnor U48181 (N_48181,N_43017,N_44639);
xnor U48182 (N_48182,N_41741,N_43463);
nor U48183 (N_48183,N_41043,N_43336);
xor U48184 (N_48184,N_44817,N_44950);
nor U48185 (N_48185,N_42309,N_43566);
and U48186 (N_48186,N_43173,N_41775);
nor U48187 (N_48187,N_43270,N_42039);
nor U48188 (N_48188,N_42714,N_41492);
and U48189 (N_48189,N_41556,N_41321);
nor U48190 (N_48190,N_41203,N_43657);
nand U48191 (N_48191,N_41486,N_44233);
and U48192 (N_48192,N_42201,N_44752);
xor U48193 (N_48193,N_42314,N_41223);
nor U48194 (N_48194,N_42598,N_40353);
and U48195 (N_48195,N_44065,N_41443);
nor U48196 (N_48196,N_40885,N_43487);
nand U48197 (N_48197,N_41431,N_40588);
xnor U48198 (N_48198,N_44566,N_40995);
or U48199 (N_48199,N_41882,N_44498);
xor U48200 (N_48200,N_42596,N_43764);
and U48201 (N_48201,N_44770,N_43517);
or U48202 (N_48202,N_41561,N_42260);
and U48203 (N_48203,N_41825,N_40651);
nand U48204 (N_48204,N_44584,N_44808);
nand U48205 (N_48205,N_44854,N_42930);
or U48206 (N_48206,N_42093,N_44455);
nor U48207 (N_48207,N_44207,N_41754);
and U48208 (N_48208,N_41350,N_40865);
and U48209 (N_48209,N_40312,N_42709);
nor U48210 (N_48210,N_40740,N_44196);
xor U48211 (N_48211,N_41869,N_44238);
and U48212 (N_48212,N_42211,N_42911);
and U48213 (N_48213,N_44131,N_44547);
xnor U48214 (N_48214,N_43544,N_40550);
and U48215 (N_48215,N_43154,N_40204);
xnor U48216 (N_48216,N_42224,N_43442);
nand U48217 (N_48217,N_41899,N_42833);
xor U48218 (N_48218,N_42295,N_40360);
nand U48219 (N_48219,N_43328,N_40976);
xor U48220 (N_48220,N_41563,N_40314);
xnor U48221 (N_48221,N_43947,N_41907);
or U48222 (N_48222,N_42801,N_43003);
nand U48223 (N_48223,N_40937,N_44362);
nand U48224 (N_48224,N_43684,N_40789);
and U48225 (N_48225,N_43562,N_42892);
and U48226 (N_48226,N_43017,N_43723);
and U48227 (N_48227,N_42323,N_41443);
nand U48228 (N_48228,N_42271,N_41673);
and U48229 (N_48229,N_44488,N_40168);
and U48230 (N_48230,N_44756,N_42922);
nand U48231 (N_48231,N_44264,N_42516);
and U48232 (N_48232,N_40413,N_40375);
nand U48233 (N_48233,N_40710,N_44364);
and U48234 (N_48234,N_40720,N_42734);
nor U48235 (N_48235,N_43226,N_44086);
xnor U48236 (N_48236,N_41985,N_40427);
nand U48237 (N_48237,N_41439,N_41536);
and U48238 (N_48238,N_41316,N_43612);
nand U48239 (N_48239,N_42600,N_44740);
nor U48240 (N_48240,N_44613,N_40862);
nor U48241 (N_48241,N_40322,N_41627);
nand U48242 (N_48242,N_41031,N_40883);
nand U48243 (N_48243,N_40222,N_44776);
nor U48244 (N_48244,N_41572,N_40086);
and U48245 (N_48245,N_44126,N_40768);
xnor U48246 (N_48246,N_43960,N_43795);
or U48247 (N_48247,N_42530,N_40741);
nor U48248 (N_48248,N_40876,N_43614);
xor U48249 (N_48249,N_40699,N_40303);
and U48250 (N_48250,N_41223,N_40605);
or U48251 (N_48251,N_44028,N_43510);
nor U48252 (N_48252,N_42423,N_43837);
or U48253 (N_48253,N_40137,N_42269);
or U48254 (N_48254,N_43729,N_41951);
xor U48255 (N_48255,N_44070,N_40945);
or U48256 (N_48256,N_43009,N_42359);
nor U48257 (N_48257,N_40476,N_41325);
xor U48258 (N_48258,N_42936,N_42009);
or U48259 (N_48259,N_40415,N_41569);
nand U48260 (N_48260,N_41010,N_40765);
nor U48261 (N_48261,N_42419,N_44475);
and U48262 (N_48262,N_44509,N_43887);
or U48263 (N_48263,N_40673,N_42409);
nor U48264 (N_48264,N_44522,N_42712);
and U48265 (N_48265,N_40559,N_44038);
nand U48266 (N_48266,N_41665,N_40696);
xnor U48267 (N_48267,N_40618,N_41414);
or U48268 (N_48268,N_43717,N_43966);
nor U48269 (N_48269,N_41527,N_42226);
or U48270 (N_48270,N_42986,N_43745);
and U48271 (N_48271,N_44793,N_44308);
and U48272 (N_48272,N_41986,N_44820);
nand U48273 (N_48273,N_40855,N_44553);
and U48274 (N_48274,N_42845,N_44247);
nand U48275 (N_48275,N_44969,N_40643);
xor U48276 (N_48276,N_42013,N_43493);
and U48277 (N_48277,N_40084,N_40649);
and U48278 (N_48278,N_43772,N_42793);
nor U48279 (N_48279,N_43165,N_44866);
nor U48280 (N_48280,N_41417,N_42121);
nand U48281 (N_48281,N_40651,N_41632);
or U48282 (N_48282,N_41576,N_42107);
and U48283 (N_48283,N_43141,N_44977);
xor U48284 (N_48284,N_43100,N_41142);
and U48285 (N_48285,N_44309,N_40702);
xor U48286 (N_48286,N_43531,N_40184);
or U48287 (N_48287,N_42778,N_41535);
and U48288 (N_48288,N_42121,N_44597);
and U48289 (N_48289,N_40446,N_42009);
nor U48290 (N_48290,N_40779,N_42741);
nand U48291 (N_48291,N_43746,N_42862);
xnor U48292 (N_48292,N_41746,N_41259);
or U48293 (N_48293,N_44646,N_43737);
or U48294 (N_48294,N_42220,N_43818);
nor U48295 (N_48295,N_41747,N_43424);
or U48296 (N_48296,N_42709,N_42752);
xnor U48297 (N_48297,N_44273,N_43320);
or U48298 (N_48298,N_44355,N_43040);
xnor U48299 (N_48299,N_41442,N_41325);
xnor U48300 (N_48300,N_43572,N_42897);
or U48301 (N_48301,N_40237,N_43154);
nand U48302 (N_48302,N_40964,N_41834);
xnor U48303 (N_48303,N_43427,N_41139);
nor U48304 (N_48304,N_43196,N_41038);
xor U48305 (N_48305,N_43291,N_43819);
xor U48306 (N_48306,N_40536,N_40018);
nand U48307 (N_48307,N_41734,N_41122);
or U48308 (N_48308,N_40279,N_40855);
and U48309 (N_48309,N_40557,N_40144);
or U48310 (N_48310,N_40305,N_43616);
xnor U48311 (N_48311,N_42909,N_42303);
nor U48312 (N_48312,N_40072,N_43965);
and U48313 (N_48313,N_44744,N_43595);
or U48314 (N_48314,N_44693,N_42728);
or U48315 (N_48315,N_41649,N_41212);
nand U48316 (N_48316,N_43232,N_42910);
or U48317 (N_48317,N_41687,N_44000);
nand U48318 (N_48318,N_40984,N_44065);
nand U48319 (N_48319,N_43413,N_44080);
nor U48320 (N_48320,N_43456,N_42603);
nand U48321 (N_48321,N_41237,N_42751);
nor U48322 (N_48322,N_40396,N_42339);
xor U48323 (N_48323,N_44767,N_42976);
nor U48324 (N_48324,N_42082,N_40675);
nor U48325 (N_48325,N_43442,N_44619);
xor U48326 (N_48326,N_44711,N_42343);
xnor U48327 (N_48327,N_43754,N_44420);
nand U48328 (N_48328,N_41882,N_42326);
nor U48329 (N_48329,N_42541,N_43943);
nor U48330 (N_48330,N_41807,N_40088);
nand U48331 (N_48331,N_41078,N_44466);
or U48332 (N_48332,N_43924,N_40666);
nor U48333 (N_48333,N_41706,N_41795);
nor U48334 (N_48334,N_41948,N_42663);
or U48335 (N_48335,N_40142,N_41213);
xor U48336 (N_48336,N_44227,N_42882);
and U48337 (N_48337,N_40005,N_42528);
nand U48338 (N_48338,N_40687,N_41911);
xnor U48339 (N_48339,N_42168,N_40709);
and U48340 (N_48340,N_42448,N_40810);
nand U48341 (N_48341,N_44621,N_41843);
nand U48342 (N_48342,N_41352,N_44544);
and U48343 (N_48343,N_40672,N_40717);
or U48344 (N_48344,N_40091,N_40264);
nor U48345 (N_48345,N_41742,N_43065);
or U48346 (N_48346,N_43227,N_44353);
nand U48347 (N_48347,N_40433,N_40159);
and U48348 (N_48348,N_42809,N_40476);
or U48349 (N_48349,N_41156,N_41574);
xor U48350 (N_48350,N_40330,N_42282);
nand U48351 (N_48351,N_44959,N_43532);
nor U48352 (N_48352,N_40889,N_40032);
and U48353 (N_48353,N_41877,N_41755);
and U48354 (N_48354,N_43531,N_40568);
nand U48355 (N_48355,N_40305,N_40756);
or U48356 (N_48356,N_43953,N_42655);
and U48357 (N_48357,N_40921,N_42832);
nor U48358 (N_48358,N_44533,N_43622);
or U48359 (N_48359,N_44950,N_42323);
and U48360 (N_48360,N_41037,N_43187);
and U48361 (N_48361,N_43045,N_40624);
nor U48362 (N_48362,N_41351,N_44320);
or U48363 (N_48363,N_40895,N_41695);
nand U48364 (N_48364,N_41121,N_44892);
nor U48365 (N_48365,N_44170,N_40145);
or U48366 (N_48366,N_44918,N_43527);
nor U48367 (N_48367,N_42264,N_42258);
nor U48368 (N_48368,N_40055,N_41006);
or U48369 (N_48369,N_41941,N_44001);
and U48370 (N_48370,N_42596,N_43497);
and U48371 (N_48371,N_42599,N_43028);
nand U48372 (N_48372,N_44729,N_44607);
or U48373 (N_48373,N_41079,N_42658);
nand U48374 (N_48374,N_40049,N_43116);
and U48375 (N_48375,N_42153,N_44824);
or U48376 (N_48376,N_44490,N_44753);
and U48377 (N_48377,N_42868,N_41810);
nand U48378 (N_48378,N_41169,N_41904);
nor U48379 (N_48379,N_42810,N_41320);
or U48380 (N_48380,N_43561,N_44547);
nand U48381 (N_48381,N_41463,N_44325);
nand U48382 (N_48382,N_42804,N_44084);
nor U48383 (N_48383,N_41085,N_41852);
and U48384 (N_48384,N_41625,N_44583);
xor U48385 (N_48385,N_44621,N_40859);
xor U48386 (N_48386,N_42244,N_40778);
nor U48387 (N_48387,N_42832,N_40309);
nor U48388 (N_48388,N_43683,N_41014);
xor U48389 (N_48389,N_40787,N_41308);
xnor U48390 (N_48390,N_41143,N_43011);
and U48391 (N_48391,N_44062,N_44107);
or U48392 (N_48392,N_42590,N_43397);
nand U48393 (N_48393,N_43244,N_44993);
nand U48394 (N_48394,N_42589,N_41604);
and U48395 (N_48395,N_41279,N_43497);
xor U48396 (N_48396,N_42923,N_44149);
and U48397 (N_48397,N_44230,N_43875);
and U48398 (N_48398,N_41129,N_42798);
nand U48399 (N_48399,N_42436,N_40258);
nand U48400 (N_48400,N_40113,N_42561);
and U48401 (N_48401,N_40478,N_44746);
nand U48402 (N_48402,N_43475,N_40720);
xnor U48403 (N_48403,N_43243,N_44340);
nor U48404 (N_48404,N_41315,N_44497);
xor U48405 (N_48405,N_42945,N_43264);
or U48406 (N_48406,N_42301,N_43787);
nand U48407 (N_48407,N_44387,N_42488);
nor U48408 (N_48408,N_43522,N_43716);
nor U48409 (N_48409,N_42229,N_42601);
or U48410 (N_48410,N_40574,N_43072);
or U48411 (N_48411,N_42588,N_42649);
nor U48412 (N_48412,N_42257,N_44469);
and U48413 (N_48413,N_43680,N_41031);
nand U48414 (N_48414,N_42895,N_42101);
and U48415 (N_48415,N_41269,N_43688);
and U48416 (N_48416,N_40722,N_41874);
nor U48417 (N_48417,N_40065,N_43513);
or U48418 (N_48418,N_44669,N_41181);
nand U48419 (N_48419,N_41685,N_41319);
and U48420 (N_48420,N_44655,N_42084);
and U48421 (N_48421,N_43811,N_42124);
and U48422 (N_48422,N_42404,N_42272);
nor U48423 (N_48423,N_40398,N_42982);
xor U48424 (N_48424,N_42021,N_44206);
and U48425 (N_48425,N_41855,N_43837);
xor U48426 (N_48426,N_40146,N_43229);
and U48427 (N_48427,N_41255,N_42258);
xnor U48428 (N_48428,N_41099,N_42175);
xnor U48429 (N_48429,N_40831,N_44848);
xnor U48430 (N_48430,N_44559,N_42547);
or U48431 (N_48431,N_41209,N_41924);
xor U48432 (N_48432,N_44973,N_41812);
and U48433 (N_48433,N_43524,N_40077);
and U48434 (N_48434,N_41284,N_44530);
nand U48435 (N_48435,N_43955,N_44739);
or U48436 (N_48436,N_41348,N_44968);
xnor U48437 (N_48437,N_43665,N_41295);
nor U48438 (N_48438,N_42825,N_40006);
xnor U48439 (N_48439,N_40712,N_41890);
or U48440 (N_48440,N_42918,N_43373);
xor U48441 (N_48441,N_41300,N_42798);
or U48442 (N_48442,N_41864,N_40038);
nand U48443 (N_48443,N_43679,N_41634);
or U48444 (N_48444,N_44239,N_44931);
and U48445 (N_48445,N_42813,N_42112);
and U48446 (N_48446,N_44274,N_44261);
or U48447 (N_48447,N_42796,N_43941);
and U48448 (N_48448,N_43358,N_43086);
and U48449 (N_48449,N_43828,N_44594);
or U48450 (N_48450,N_41179,N_41043);
and U48451 (N_48451,N_40977,N_41728);
nor U48452 (N_48452,N_42383,N_41752);
and U48453 (N_48453,N_40982,N_44279);
nor U48454 (N_48454,N_41482,N_44983);
nand U48455 (N_48455,N_41299,N_40084);
nand U48456 (N_48456,N_40969,N_43140);
nor U48457 (N_48457,N_40623,N_41836);
nand U48458 (N_48458,N_42246,N_43531);
xor U48459 (N_48459,N_43596,N_41393);
nand U48460 (N_48460,N_44344,N_43028);
nand U48461 (N_48461,N_44719,N_42004);
xor U48462 (N_48462,N_42411,N_40552);
and U48463 (N_48463,N_42292,N_44550);
nor U48464 (N_48464,N_43764,N_44629);
xor U48465 (N_48465,N_41246,N_42087);
nand U48466 (N_48466,N_41999,N_44185);
nand U48467 (N_48467,N_41052,N_42251);
nor U48468 (N_48468,N_44709,N_42371);
or U48469 (N_48469,N_44762,N_41350);
or U48470 (N_48470,N_42975,N_41312);
nand U48471 (N_48471,N_40545,N_40848);
nor U48472 (N_48472,N_43591,N_42640);
nand U48473 (N_48473,N_40112,N_43061);
or U48474 (N_48474,N_44153,N_42475);
or U48475 (N_48475,N_40613,N_43747);
or U48476 (N_48476,N_43672,N_44839);
xor U48477 (N_48477,N_43307,N_42937);
xor U48478 (N_48478,N_41451,N_41030);
nand U48479 (N_48479,N_43411,N_42356);
xor U48480 (N_48480,N_40772,N_43684);
and U48481 (N_48481,N_42708,N_44014);
xnor U48482 (N_48482,N_44895,N_40935);
nand U48483 (N_48483,N_44013,N_41968);
xnor U48484 (N_48484,N_40061,N_44297);
or U48485 (N_48485,N_41185,N_41796);
or U48486 (N_48486,N_44652,N_42279);
xor U48487 (N_48487,N_43034,N_44260);
and U48488 (N_48488,N_42947,N_44163);
nand U48489 (N_48489,N_41980,N_41887);
and U48490 (N_48490,N_42915,N_40995);
nand U48491 (N_48491,N_40538,N_41644);
xor U48492 (N_48492,N_41547,N_43635);
nor U48493 (N_48493,N_43714,N_42728);
or U48494 (N_48494,N_42718,N_44096);
xor U48495 (N_48495,N_42710,N_41406);
or U48496 (N_48496,N_44808,N_41479);
or U48497 (N_48497,N_43272,N_40970);
nand U48498 (N_48498,N_44604,N_44146);
nor U48499 (N_48499,N_41760,N_41474);
nor U48500 (N_48500,N_41376,N_40273);
or U48501 (N_48501,N_41148,N_42231);
xor U48502 (N_48502,N_40360,N_43547);
and U48503 (N_48503,N_42232,N_42106);
and U48504 (N_48504,N_43676,N_44819);
nand U48505 (N_48505,N_40095,N_44908);
or U48506 (N_48506,N_41375,N_42752);
and U48507 (N_48507,N_40315,N_40059);
xnor U48508 (N_48508,N_43708,N_40400);
and U48509 (N_48509,N_44461,N_43000);
nor U48510 (N_48510,N_44641,N_43932);
nand U48511 (N_48511,N_40454,N_44218);
xor U48512 (N_48512,N_44918,N_43255);
nand U48513 (N_48513,N_44113,N_44475);
nand U48514 (N_48514,N_42819,N_42234);
xor U48515 (N_48515,N_41950,N_40099);
nor U48516 (N_48516,N_43843,N_41401);
or U48517 (N_48517,N_40474,N_44402);
or U48518 (N_48518,N_42930,N_41810);
or U48519 (N_48519,N_40213,N_41753);
and U48520 (N_48520,N_43326,N_41300);
nand U48521 (N_48521,N_41297,N_41180);
or U48522 (N_48522,N_40126,N_40590);
nor U48523 (N_48523,N_44275,N_40193);
nor U48524 (N_48524,N_44298,N_40584);
xor U48525 (N_48525,N_43902,N_41253);
and U48526 (N_48526,N_40990,N_43579);
and U48527 (N_48527,N_44565,N_44857);
nand U48528 (N_48528,N_43608,N_40093);
or U48529 (N_48529,N_43929,N_43953);
nor U48530 (N_48530,N_44193,N_41312);
or U48531 (N_48531,N_42222,N_40128);
nor U48532 (N_48532,N_43091,N_40426);
xor U48533 (N_48533,N_42318,N_42507);
and U48534 (N_48534,N_44714,N_44052);
or U48535 (N_48535,N_42273,N_40483);
or U48536 (N_48536,N_41420,N_42702);
or U48537 (N_48537,N_40907,N_40152);
nor U48538 (N_48538,N_42546,N_42588);
or U48539 (N_48539,N_43604,N_41755);
and U48540 (N_48540,N_40471,N_44079);
or U48541 (N_48541,N_41306,N_40018);
or U48542 (N_48542,N_42720,N_43363);
and U48543 (N_48543,N_41660,N_42958);
xor U48544 (N_48544,N_41810,N_40137);
and U48545 (N_48545,N_43356,N_43612);
and U48546 (N_48546,N_44026,N_44719);
nand U48547 (N_48547,N_44776,N_42396);
nor U48548 (N_48548,N_44803,N_40247);
nand U48549 (N_48549,N_41845,N_42153);
nand U48550 (N_48550,N_41391,N_42504);
or U48551 (N_48551,N_42760,N_44841);
nand U48552 (N_48552,N_44487,N_40609);
xor U48553 (N_48553,N_41398,N_42948);
or U48554 (N_48554,N_43423,N_42025);
nand U48555 (N_48555,N_43668,N_41023);
and U48556 (N_48556,N_44244,N_44307);
nor U48557 (N_48557,N_43301,N_43076);
xnor U48558 (N_48558,N_43932,N_41258);
or U48559 (N_48559,N_43412,N_44565);
xnor U48560 (N_48560,N_40889,N_42235);
nand U48561 (N_48561,N_40509,N_40640);
and U48562 (N_48562,N_40444,N_43406);
nor U48563 (N_48563,N_43225,N_42799);
or U48564 (N_48564,N_40506,N_40781);
and U48565 (N_48565,N_42648,N_42658);
or U48566 (N_48566,N_43638,N_43135);
and U48567 (N_48567,N_41988,N_40515);
or U48568 (N_48568,N_40414,N_43609);
nor U48569 (N_48569,N_42911,N_41280);
xor U48570 (N_48570,N_41875,N_40972);
nor U48571 (N_48571,N_42670,N_43819);
or U48572 (N_48572,N_44254,N_41574);
and U48573 (N_48573,N_44641,N_43910);
and U48574 (N_48574,N_42947,N_41375);
nor U48575 (N_48575,N_40784,N_44759);
or U48576 (N_48576,N_42971,N_43072);
or U48577 (N_48577,N_44218,N_43096);
and U48578 (N_48578,N_40124,N_43295);
nand U48579 (N_48579,N_44119,N_44259);
and U48580 (N_48580,N_42848,N_41044);
nor U48581 (N_48581,N_43912,N_44416);
or U48582 (N_48582,N_40065,N_44877);
or U48583 (N_48583,N_43443,N_43726);
xor U48584 (N_48584,N_42421,N_41639);
nor U48585 (N_48585,N_41020,N_40801);
nor U48586 (N_48586,N_41520,N_43799);
or U48587 (N_48587,N_42725,N_40206);
nand U48588 (N_48588,N_43818,N_42795);
nor U48589 (N_48589,N_43015,N_42202);
or U48590 (N_48590,N_43837,N_42951);
or U48591 (N_48591,N_42156,N_42235);
nor U48592 (N_48592,N_44601,N_42173);
or U48593 (N_48593,N_44359,N_44066);
and U48594 (N_48594,N_41340,N_43684);
and U48595 (N_48595,N_42110,N_42058);
nand U48596 (N_48596,N_41163,N_42626);
nor U48597 (N_48597,N_40755,N_44891);
or U48598 (N_48598,N_43342,N_43983);
and U48599 (N_48599,N_43067,N_40459);
nor U48600 (N_48600,N_40378,N_40598);
nor U48601 (N_48601,N_40244,N_42551);
nor U48602 (N_48602,N_43668,N_40187);
nand U48603 (N_48603,N_41014,N_41996);
xor U48604 (N_48604,N_44242,N_40869);
and U48605 (N_48605,N_40670,N_44457);
and U48606 (N_48606,N_43627,N_41408);
xor U48607 (N_48607,N_44662,N_44064);
and U48608 (N_48608,N_40184,N_41238);
xnor U48609 (N_48609,N_43984,N_41679);
nor U48610 (N_48610,N_43659,N_40564);
xor U48611 (N_48611,N_41067,N_44077);
nor U48612 (N_48612,N_44907,N_43480);
nor U48613 (N_48613,N_40308,N_43397);
or U48614 (N_48614,N_41817,N_44725);
xor U48615 (N_48615,N_44046,N_40364);
nor U48616 (N_48616,N_44780,N_42992);
nor U48617 (N_48617,N_43828,N_40290);
or U48618 (N_48618,N_44600,N_43988);
or U48619 (N_48619,N_44958,N_43621);
nor U48620 (N_48620,N_42479,N_44000);
nor U48621 (N_48621,N_40790,N_40275);
or U48622 (N_48622,N_44807,N_41818);
nand U48623 (N_48623,N_44843,N_41848);
nor U48624 (N_48624,N_41555,N_42194);
nor U48625 (N_48625,N_44481,N_43073);
xnor U48626 (N_48626,N_42851,N_40949);
xor U48627 (N_48627,N_41923,N_40210);
xor U48628 (N_48628,N_42576,N_44439);
or U48629 (N_48629,N_41481,N_42398);
and U48630 (N_48630,N_43532,N_40735);
nor U48631 (N_48631,N_43566,N_40964);
or U48632 (N_48632,N_42638,N_43193);
nand U48633 (N_48633,N_44456,N_40727);
or U48634 (N_48634,N_40750,N_40373);
nor U48635 (N_48635,N_44645,N_40454);
xor U48636 (N_48636,N_42595,N_42817);
and U48637 (N_48637,N_43840,N_41141);
nand U48638 (N_48638,N_41687,N_42685);
and U48639 (N_48639,N_42272,N_40856);
and U48640 (N_48640,N_44222,N_42171);
nor U48641 (N_48641,N_40500,N_42645);
and U48642 (N_48642,N_44857,N_40564);
nor U48643 (N_48643,N_44266,N_41921);
or U48644 (N_48644,N_43897,N_43159);
nand U48645 (N_48645,N_42023,N_44522);
nand U48646 (N_48646,N_43192,N_41228);
nor U48647 (N_48647,N_44479,N_43155);
nor U48648 (N_48648,N_42354,N_41212);
and U48649 (N_48649,N_42070,N_44017);
nor U48650 (N_48650,N_44019,N_41322);
nand U48651 (N_48651,N_44781,N_42451);
xnor U48652 (N_48652,N_42161,N_42939);
and U48653 (N_48653,N_44232,N_42026);
and U48654 (N_48654,N_44572,N_42444);
nor U48655 (N_48655,N_43242,N_42136);
xor U48656 (N_48656,N_40039,N_40890);
and U48657 (N_48657,N_44285,N_40138);
or U48658 (N_48658,N_40023,N_44204);
nor U48659 (N_48659,N_40472,N_41114);
nor U48660 (N_48660,N_41290,N_44595);
or U48661 (N_48661,N_41612,N_41223);
or U48662 (N_48662,N_44681,N_40066);
nand U48663 (N_48663,N_44294,N_41083);
and U48664 (N_48664,N_41286,N_42398);
nand U48665 (N_48665,N_42334,N_41597);
and U48666 (N_48666,N_40660,N_43480);
or U48667 (N_48667,N_41257,N_43463);
nor U48668 (N_48668,N_40167,N_40260);
and U48669 (N_48669,N_43582,N_43110);
or U48670 (N_48670,N_42393,N_44062);
xor U48671 (N_48671,N_41055,N_41953);
nor U48672 (N_48672,N_42089,N_41569);
nor U48673 (N_48673,N_43353,N_43731);
xnor U48674 (N_48674,N_41571,N_42322);
and U48675 (N_48675,N_40313,N_41773);
xnor U48676 (N_48676,N_41185,N_44216);
and U48677 (N_48677,N_42033,N_40697);
nand U48678 (N_48678,N_42377,N_40214);
nand U48679 (N_48679,N_44225,N_42577);
nor U48680 (N_48680,N_44164,N_44866);
nand U48681 (N_48681,N_40576,N_44759);
nand U48682 (N_48682,N_43866,N_41296);
and U48683 (N_48683,N_44569,N_42553);
and U48684 (N_48684,N_44358,N_43347);
nor U48685 (N_48685,N_40225,N_43429);
and U48686 (N_48686,N_42217,N_42467);
and U48687 (N_48687,N_42100,N_41373);
nand U48688 (N_48688,N_41340,N_43721);
nor U48689 (N_48689,N_40880,N_43739);
and U48690 (N_48690,N_41804,N_40916);
and U48691 (N_48691,N_43900,N_41289);
and U48692 (N_48692,N_42614,N_41350);
xnor U48693 (N_48693,N_43786,N_43677);
and U48694 (N_48694,N_44006,N_42307);
nand U48695 (N_48695,N_42350,N_40197);
nor U48696 (N_48696,N_44808,N_42068);
or U48697 (N_48697,N_40512,N_42139);
xor U48698 (N_48698,N_44816,N_41858);
or U48699 (N_48699,N_44001,N_43236);
xnor U48700 (N_48700,N_42028,N_42921);
nand U48701 (N_48701,N_41360,N_44235);
xnor U48702 (N_48702,N_41126,N_42306);
xor U48703 (N_48703,N_40070,N_41189);
or U48704 (N_48704,N_41566,N_41055);
nor U48705 (N_48705,N_43339,N_43666);
and U48706 (N_48706,N_40517,N_42973);
nand U48707 (N_48707,N_42738,N_42327);
and U48708 (N_48708,N_41989,N_41353);
nand U48709 (N_48709,N_44852,N_43960);
and U48710 (N_48710,N_42153,N_41254);
nand U48711 (N_48711,N_44662,N_43371);
or U48712 (N_48712,N_44319,N_44858);
xor U48713 (N_48713,N_40598,N_41423);
nand U48714 (N_48714,N_41055,N_44734);
xnor U48715 (N_48715,N_41996,N_44751);
xnor U48716 (N_48716,N_42839,N_40469);
nor U48717 (N_48717,N_44933,N_42511);
or U48718 (N_48718,N_42771,N_40475);
nand U48719 (N_48719,N_43144,N_41039);
nor U48720 (N_48720,N_40460,N_41221);
and U48721 (N_48721,N_41910,N_40703);
nor U48722 (N_48722,N_44484,N_41421);
xor U48723 (N_48723,N_40536,N_43587);
xnor U48724 (N_48724,N_43290,N_41207);
xor U48725 (N_48725,N_40257,N_42678);
or U48726 (N_48726,N_42191,N_44617);
nand U48727 (N_48727,N_41282,N_40537);
nor U48728 (N_48728,N_41241,N_44561);
xor U48729 (N_48729,N_40722,N_41615);
and U48730 (N_48730,N_43268,N_42486);
nand U48731 (N_48731,N_44729,N_43610);
nand U48732 (N_48732,N_41579,N_41374);
or U48733 (N_48733,N_42483,N_40375);
nand U48734 (N_48734,N_44639,N_42324);
xnor U48735 (N_48735,N_40766,N_42434);
and U48736 (N_48736,N_40904,N_41657);
nand U48737 (N_48737,N_43839,N_41344);
nand U48738 (N_48738,N_42499,N_42245);
nor U48739 (N_48739,N_41088,N_43435);
nor U48740 (N_48740,N_42279,N_41400);
or U48741 (N_48741,N_44630,N_41010);
and U48742 (N_48742,N_43792,N_44382);
nand U48743 (N_48743,N_44675,N_43060);
or U48744 (N_48744,N_43007,N_42936);
or U48745 (N_48745,N_44093,N_43795);
nand U48746 (N_48746,N_40776,N_40073);
nand U48747 (N_48747,N_44470,N_42752);
and U48748 (N_48748,N_41111,N_40577);
nor U48749 (N_48749,N_42726,N_40691);
xnor U48750 (N_48750,N_40572,N_42689);
nor U48751 (N_48751,N_40219,N_41512);
nand U48752 (N_48752,N_43443,N_43260);
nand U48753 (N_48753,N_43535,N_41143);
and U48754 (N_48754,N_41191,N_41029);
and U48755 (N_48755,N_40933,N_42188);
or U48756 (N_48756,N_44601,N_44874);
nor U48757 (N_48757,N_41776,N_44360);
nor U48758 (N_48758,N_43289,N_41305);
and U48759 (N_48759,N_42317,N_44480);
or U48760 (N_48760,N_41284,N_40685);
nor U48761 (N_48761,N_41145,N_40817);
or U48762 (N_48762,N_42555,N_42778);
nand U48763 (N_48763,N_40742,N_41105);
and U48764 (N_48764,N_41226,N_44609);
and U48765 (N_48765,N_41413,N_44816);
nor U48766 (N_48766,N_43974,N_43082);
nand U48767 (N_48767,N_43232,N_41246);
nand U48768 (N_48768,N_44015,N_44268);
nand U48769 (N_48769,N_40864,N_41910);
or U48770 (N_48770,N_40119,N_40327);
or U48771 (N_48771,N_41143,N_41582);
nand U48772 (N_48772,N_41478,N_44028);
xor U48773 (N_48773,N_40078,N_40257);
nor U48774 (N_48774,N_43469,N_44464);
nor U48775 (N_48775,N_41418,N_43057);
nor U48776 (N_48776,N_40726,N_43508);
nand U48777 (N_48777,N_42084,N_42787);
or U48778 (N_48778,N_44835,N_43438);
nand U48779 (N_48779,N_41430,N_40087);
or U48780 (N_48780,N_40152,N_43724);
nor U48781 (N_48781,N_44697,N_43791);
xor U48782 (N_48782,N_41938,N_43671);
xnor U48783 (N_48783,N_42617,N_41406);
or U48784 (N_48784,N_40395,N_40553);
nor U48785 (N_48785,N_44568,N_43194);
nand U48786 (N_48786,N_40338,N_41071);
nor U48787 (N_48787,N_41250,N_42314);
xnor U48788 (N_48788,N_40589,N_44226);
nor U48789 (N_48789,N_43018,N_44335);
nand U48790 (N_48790,N_40744,N_40869);
or U48791 (N_48791,N_42130,N_42720);
or U48792 (N_48792,N_40050,N_43407);
nand U48793 (N_48793,N_40184,N_43974);
or U48794 (N_48794,N_43577,N_43866);
nand U48795 (N_48795,N_41141,N_40916);
and U48796 (N_48796,N_40289,N_43997);
or U48797 (N_48797,N_42541,N_42949);
and U48798 (N_48798,N_44312,N_40038);
nand U48799 (N_48799,N_44952,N_44707);
xor U48800 (N_48800,N_41532,N_44648);
xor U48801 (N_48801,N_43922,N_41544);
xnor U48802 (N_48802,N_40487,N_41265);
and U48803 (N_48803,N_43043,N_42057);
nand U48804 (N_48804,N_44913,N_41987);
xor U48805 (N_48805,N_42207,N_40901);
nand U48806 (N_48806,N_43950,N_43378);
xnor U48807 (N_48807,N_41514,N_42451);
nor U48808 (N_48808,N_41227,N_44504);
nor U48809 (N_48809,N_43890,N_42549);
xnor U48810 (N_48810,N_42771,N_41132);
or U48811 (N_48811,N_43768,N_42065);
and U48812 (N_48812,N_42155,N_40309);
nand U48813 (N_48813,N_41883,N_43583);
and U48814 (N_48814,N_43010,N_43507);
xor U48815 (N_48815,N_42368,N_42539);
nor U48816 (N_48816,N_41074,N_44392);
nand U48817 (N_48817,N_43920,N_42333);
nor U48818 (N_48818,N_42637,N_43830);
nor U48819 (N_48819,N_42244,N_42302);
nand U48820 (N_48820,N_41161,N_42653);
or U48821 (N_48821,N_40492,N_41316);
nor U48822 (N_48822,N_41945,N_42614);
xnor U48823 (N_48823,N_40591,N_44423);
nand U48824 (N_48824,N_44105,N_43274);
nand U48825 (N_48825,N_42480,N_43423);
or U48826 (N_48826,N_40236,N_44591);
nand U48827 (N_48827,N_40237,N_42791);
nor U48828 (N_48828,N_40039,N_42211);
and U48829 (N_48829,N_43520,N_43138);
or U48830 (N_48830,N_40643,N_42310);
nor U48831 (N_48831,N_43982,N_40504);
nor U48832 (N_48832,N_40279,N_42472);
and U48833 (N_48833,N_42627,N_40458);
or U48834 (N_48834,N_40969,N_44851);
nand U48835 (N_48835,N_42197,N_41221);
nor U48836 (N_48836,N_43309,N_43814);
nand U48837 (N_48837,N_41245,N_40840);
nand U48838 (N_48838,N_44323,N_42347);
or U48839 (N_48839,N_40655,N_44189);
xnor U48840 (N_48840,N_43382,N_40006);
xnor U48841 (N_48841,N_44992,N_40625);
nand U48842 (N_48842,N_41099,N_44027);
or U48843 (N_48843,N_44913,N_41059);
nor U48844 (N_48844,N_43269,N_43272);
or U48845 (N_48845,N_42937,N_40950);
or U48846 (N_48846,N_43694,N_41240);
and U48847 (N_48847,N_42974,N_44565);
nand U48848 (N_48848,N_43230,N_40959);
nand U48849 (N_48849,N_41231,N_42505);
and U48850 (N_48850,N_43637,N_44399);
nand U48851 (N_48851,N_42835,N_41011);
nor U48852 (N_48852,N_40453,N_42993);
nand U48853 (N_48853,N_42572,N_44566);
nor U48854 (N_48854,N_41171,N_43850);
and U48855 (N_48855,N_43578,N_44012);
xor U48856 (N_48856,N_42300,N_41878);
nand U48857 (N_48857,N_41406,N_43078);
or U48858 (N_48858,N_44126,N_44082);
xor U48859 (N_48859,N_41505,N_44863);
nand U48860 (N_48860,N_43785,N_42920);
nand U48861 (N_48861,N_42731,N_44797);
or U48862 (N_48862,N_43315,N_42782);
and U48863 (N_48863,N_42018,N_42345);
or U48864 (N_48864,N_40747,N_42702);
nor U48865 (N_48865,N_44647,N_41685);
and U48866 (N_48866,N_43307,N_41209);
nand U48867 (N_48867,N_44013,N_40968);
or U48868 (N_48868,N_43101,N_41086);
and U48869 (N_48869,N_42997,N_44990);
nand U48870 (N_48870,N_44763,N_41369);
nand U48871 (N_48871,N_44959,N_43805);
or U48872 (N_48872,N_44712,N_44577);
xor U48873 (N_48873,N_42585,N_40766);
nand U48874 (N_48874,N_44104,N_40236);
xnor U48875 (N_48875,N_42104,N_41395);
nor U48876 (N_48876,N_44995,N_40440);
nor U48877 (N_48877,N_40151,N_41821);
xnor U48878 (N_48878,N_43226,N_43858);
nor U48879 (N_48879,N_42912,N_42232);
and U48880 (N_48880,N_41516,N_43136);
xnor U48881 (N_48881,N_41927,N_42788);
xor U48882 (N_48882,N_41718,N_44518);
and U48883 (N_48883,N_42728,N_41603);
nor U48884 (N_48884,N_42377,N_42612);
xor U48885 (N_48885,N_40098,N_40241);
nand U48886 (N_48886,N_44071,N_42609);
xor U48887 (N_48887,N_40615,N_40020);
nor U48888 (N_48888,N_42948,N_40526);
or U48889 (N_48889,N_40464,N_40217);
nor U48890 (N_48890,N_42539,N_41611);
xnor U48891 (N_48891,N_42276,N_41622);
nor U48892 (N_48892,N_40925,N_41323);
xor U48893 (N_48893,N_41193,N_40110);
nand U48894 (N_48894,N_42716,N_41328);
xor U48895 (N_48895,N_41001,N_44863);
xnor U48896 (N_48896,N_40950,N_41158);
or U48897 (N_48897,N_40192,N_40965);
nand U48898 (N_48898,N_44945,N_43788);
nand U48899 (N_48899,N_44949,N_44505);
xor U48900 (N_48900,N_40698,N_43474);
nor U48901 (N_48901,N_43822,N_43079);
nand U48902 (N_48902,N_40596,N_40777);
xnor U48903 (N_48903,N_42839,N_42561);
or U48904 (N_48904,N_41830,N_44138);
nand U48905 (N_48905,N_44120,N_40656);
nor U48906 (N_48906,N_43391,N_41791);
xor U48907 (N_48907,N_44205,N_40722);
nor U48908 (N_48908,N_41007,N_42550);
nor U48909 (N_48909,N_42321,N_40857);
and U48910 (N_48910,N_44430,N_40739);
or U48911 (N_48911,N_44007,N_42130);
xor U48912 (N_48912,N_40305,N_42339);
xnor U48913 (N_48913,N_41855,N_43733);
nor U48914 (N_48914,N_44466,N_41224);
nor U48915 (N_48915,N_43120,N_44717);
and U48916 (N_48916,N_41686,N_40080);
xnor U48917 (N_48917,N_42349,N_42119);
and U48918 (N_48918,N_40800,N_43867);
and U48919 (N_48919,N_41269,N_44638);
or U48920 (N_48920,N_43172,N_43291);
nand U48921 (N_48921,N_41152,N_40298);
xor U48922 (N_48922,N_42016,N_40278);
or U48923 (N_48923,N_44278,N_42763);
xor U48924 (N_48924,N_40988,N_44314);
nor U48925 (N_48925,N_43801,N_44118);
or U48926 (N_48926,N_41521,N_41250);
and U48927 (N_48927,N_42655,N_43511);
nor U48928 (N_48928,N_42550,N_43178);
xnor U48929 (N_48929,N_42190,N_44142);
or U48930 (N_48930,N_42172,N_43835);
xor U48931 (N_48931,N_42963,N_43103);
nand U48932 (N_48932,N_41636,N_40693);
or U48933 (N_48933,N_40594,N_43631);
xnor U48934 (N_48934,N_40659,N_42512);
nand U48935 (N_48935,N_43647,N_43618);
xor U48936 (N_48936,N_44264,N_44832);
nor U48937 (N_48937,N_43014,N_43882);
nor U48938 (N_48938,N_40339,N_42910);
or U48939 (N_48939,N_40827,N_41510);
or U48940 (N_48940,N_40264,N_44292);
nand U48941 (N_48941,N_41669,N_44450);
nand U48942 (N_48942,N_41387,N_42949);
xor U48943 (N_48943,N_42348,N_44708);
xor U48944 (N_48944,N_42027,N_42450);
nor U48945 (N_48945,N_43704,N_43028);
nor U48946 (N_48946,N_44395,N_44718);
xor U48947 (N_48947,N_41022,N_43773);
nand U48948 (N_48948,N_41760,N_43666);
or U48949 (N_48949,N_43607,N_41472);
or U48950 (N_48950,N_41820,N_40881);
nand U48951 (N_48951,N_44829,N_42190);
nand U48952 (N_48952,N_43321,N_40926);
xnor U48953 (N_48953,N_43872,N_43581);
and U48954 (N_48954,N_41349,N_40926);
nor U48955 (N_48955,N_43082,N_41345);
and U48956 (N_48956,N_42458,N_41789);
and U48957 (N_48957,N_41333,N_44169);
or U48958 (N_48958,N_44471,N_42228);
and U48959 (N_48959,N_40874,N_43519);
and U48960 (N_48960,N_41359,N_43515);
and U48961 (N_48961,N_40845,N_43109);
and U48962 (N_48962,N_42291,N_42685);
and U48963 (N_48963,N_41593,N_44097);
nor U48964 (N_48964,N_44267,N_42542);
xnor U48965 (N_48965,N_41756,N_43721);
nor U48966 (N_48966,N_43130,N_44345);
or U48967 (N_48967,N_41562,N_44143);
nand U48968 (N_48968,N_40163,N_44196);
xor U48969 (N_48969,N_43649,N_40565);
and U48970 (N_48970,N_40609,N_41090);
nor U48971 (N_48971,N_40106,N_41941);
or U48972 (N_48972,N_40481,N_43266);
xor U48973 (N_48973,N_43250,N_42628);
nand U48974 (N_48974,N_43636,N_43264);
nand U48975 (N_48975,N_41842,N_40611);
or U48976 (N_48976,N_43192,N_42945);
nand U48977 (N_48977,N_43247,N_43194);
and U48978 (N_48978,N_42163,N_40856);
nor U48979 (N_48979,N_40418,N_42103);
nor U48980 (N_48980,N_43578,N_44638);
nor U48981 (N_48981,N_43583,N_44099);
and U48982 (N_48982,N_41237,N_43621);
nor U48983 (N_48983,N_40491,N_42189);
and U48984 (N_48984,N_44477,N_44786);
nand U48985 (N_48985,N_42593,N_43870);
nand U48986 (N_48986,N_44144,N_44459);
nand U48987 (N_48987,N_42701,N_40988);
or U48988 (N_48988,N_43712,N_41479);
or U48989 (N_48989,N_42620,N_42876);
nor U48990 (N_48990,N_40885,N_42937);
and U48991 (N_48991,N_43429,N_43125);
nand U48992 (N_48992,N_42247,N_42298);
xnor U48993 (N_48993,N_42276,N_41930);
nor U48994 (N_48994,N_41245,N_41493);
nor U48995 (N_48995,N_43042,N_42664);
or U48996 (N_48996,N_41141,N_40699);
nand U48997 (N_48997,N_44424,N_41509);
nor U48998 (N_48998,N_42801,N_44971);
xor U48999 (N_48999,N_42660,N_40334);
and U49000 (N_49000,N_40970,N_40532);
nand U49001 (N_49001,N_43158,N_43534);
xnor U49002 (N_49002,N_41435,N_40080);
nand U49003 (N_49003,N_41303,N_44626);
and U49004 (N_49004,N_40725,N_40708);
nor U49005 (N_49005,N_40386,N_44655);
nand U49006 (N_49006,N_40713,N_42462);
nor U49007 (N_49007,N_40875,N_44326);
xor U49008 (N_49008,N_42803,N_43364);
and U49009 (N_49009,N_40376,N_40123);
or U49010 (N_49010,N_41405,N_42433);
nor U49011 (N_49011,N_43675,N_41099);
or U49012 (N_49012,N_44058,N_41823);
nor U49013 (N_49013,N_42684,N_43080);
nand U49014 (N_49014,N_44743,N_41463);
or U49015 (N_49015,N_44968,N_42643);
xnor U49016 (N_49016,N_41462,N_44526);
or U49017 (N_49017,N_43512,N_43147);
or U49018 (N_49018,N_44559,N_40810);
or U49019 (N_49019,N_42531,N_42608);
xor U49020 (N_49020,N_40767,N_42237);
and U49021 (N_49021,N_41245,N_43787);
xnor U49022 (N_49022,N_44167,N_44723);
xnor U49023 (N_49023,N_43642,N_41967);
nand U49024 (N_49024,N_42748,N_40108);
or U49025 (N_49025,N_41183,N_44550);
and U49026 (N_49026,N_42528,N_44675);
nor U49027 (N_49027,N_40590,N_44698);
and U49028 (N_49028,N_40975,N_40776);
and U49029 (N_49029,N_41772,N_42969);
and U49030 (N_49030,N_40741,N_42787);
nor U49031 (N_49031,N_43189,N_43525);
and U49032 (N_49032,N_42500,N_42418);
or U49033 (N_49033,N_43924,N_43525);
and U49034 (N_49034,N_43609,N_41992);
and U49035 (N_49035,N_42433,N_43332);
xor U49036 (N_49036,N_42047,N_44493);
nor U49037 (N_49037,N_40996,N_41791);
and U49038 (N_49038,N_41512,N_41277);
and U49039 (N_49039,N_42509,N_41342);
xor U49040 (N_49040,N_44565,N_44387);
or U49041 (N_49041,N_42520,N_43511);
and U49042 (N_49042,N_40482,N_43520);
and U49043 (N_49043,N_42866,N_41021);
or U49044 (N_49044,N_43677,N_42191);
xor U49045 (N_49045,N_42175,N_44704);
or U49046 (N_49046,N_42161,N_44966);
xnor U49047 (N_49047,N_43390,N_44885);
and U49048 (N_49048,N_42373,N_40430);
and U49049 (N_49049,N_40078,N_40207);
xor U49050 (N_49050,N_42090,N_43987);
xor U49051 (N_49051,N_43563,N_42563);
and U49052 (N_49052,N_44849,N_43830);
and U49053 (N_49053,N_44797,N_41950);
nor U49054 (N_49054,N_43757,N_42760);
and U49055 (N_49055,N_43642,N_40069);
nor U49056 (N_49056,N_43142,N_43469);
nor U49057 (N_49057,N_40837,N_40107);
nand U49058 (N_49058,N_44775,N_41299);
nor U49059 (N_49059,N_44920,N_44205);
and U49060 (N_49060,N_42351,N_40917);
nor U49061 (N_49061,N_43559,N_41271);
nor U49062 (N_49062,N_40722,N_41799);
and U49063 (N_49063,N_43265,N_42410);
xnor U49064 (N_49064,N_43662,N_40125);
nor U49065 (N_49065,N_44723,N_41987);
nand U49066 (N_49066,N_41340,N_40702);
nor U49067 (N_49067,N_43585,N_44052);
or U49068 (N_49068,N_43851,N_43635);
nand U49069 (N_49069,N_44826,N_41384);
nand U49070 (N_49070,N_40097,N_44130);
and U49071 (N_49071,N_42777,N_41260);
nand U49072 (N_49072,N_42933,N_44359);
nor U49073 (N_49073,N_40423,N_40133);
nor U49074 (N_49074,N_43993,N_43048);
and U49075 (N_49075,N_41099,N_44149);
nor U49076 (N_49076,N_44947,N_44893);
and U49077 (N_49077,N_44185,N_43181);
xnor U49078 (N_49078,N_40638,N_44163);
nand U49079 (N_49079,N_40627,N_40323);
or U49080 (N_49080,N_42097,N_40899);
xnor U49081 (N_49081,N_41920,N_44978);
xor U49082 (N_49082,N_42153,N_41882);
xnor U49083 (N_49083,N_42573,N_42257);
nor U49084 (N_49084,N_44973,N_43413);
xor U49085 (N_49085,N_40594,N_43195);
and U49086 (N_49086,N_44016,N_42182);
nor U49087 (N_49087,N_42277,N_42570);
nor U49088 (N_49088,N_44162,N_43435);
and U49089 (N_49089,N_41094,N_42667);
or U49090 (N_49090,N_44127,N_44552);
xor U49091 (N_49091,N_40018,N_42102);
nor U49092 (N_49092,N_43839,N_43777);
and U49093 (N_49093,N_43176,N_44948);
or U49094 (N_49094,N_44790,N_44258);
xnor U49095 (N_49095,N_41198,N_42199);
or U49096 (N_49096,N_40357,N_40120);
and U49097 (N_49097,N_40442,N_44777);
xnor U49098 (N_49098,N_40714,N_44608);
nand U49099 (N_49099,N_43859,N_41591);
nand U49100 (N_49100,N_40598,N_40316);
nand U49101 (N_49101,N_41061,N_42456);
xor U49102 (N_49102,N_44519,N_41428);
and U49103 (N_49103,N_44524,N_42106);
xor U49104 (N_49104,N_41613,N_43804);
nand U49105 (N_49105,N_43257,N_41432);
or U49106 (N_49106,N_43042,N_42415);
nand U49107 (N_49107,N_40130,N_43690);
nor U49108 (N_49108,N_42169,N_42276);
nand U49109 (N_49109,N_42141,N_42646);
and U49110 (N_49110,N_44934,N_44792);
nor U49111 (N_49111,N_43585,N_40387);
or U49112 (N_49112,N_43147,N_41360);
and U49113 (N_49113,N_44528,N_40860);
xor U49114 (N_49114,N_41489,N_42582);
xnor U49115 (N_49115,N_42283,N_44065);
or U49116 (N_49116,N_42122,N_42789);
nand U49117 (N_49117,N_40118,N_42111);
nand U49118 (N_49118,N_44284,N_44650);
and U49119 (N_49119,N_43163,N_44338);
xor U49120 (N_49120,N_43068,N_41228);
nor U49121 (N_49121,N_44452,N_44900);
or U49122 (N_49122,N_44309,N_42598);
nor U49123 (N_49123,N_42406,N_40539);
or U49124 (N_49124,N_40349,N_44959);
nor U49125 (N_49125,N_43266,N_43337);
or U49126 (N_49126,N_42623,N_42807);
xnor U49127 (N_49127,N_41528,N_40484);
xor U49128 (N_49128,N_43220,N_41751);
or U49129 (N_49129,N_41982,N_40500);
xnor U49130 (N_49130,N_44802,N_42890);
nand U49131 (N_49131,N_44887,N_42938);
and U49132 (N_49132,N_40072,N_41889);
and U49133 (N_49133,N_41803,N_40627);
and U49134 (N_49134,N_41565,N_44161);
and U49135 (N_49135,N_41480,N_40673);
xor U49136 (N_49136,N_43860,N_41807);
xnor U49137 (N_49137,N_43342,N_42054);
nor U49138 (N_49138,N_41368,N_40632);
nand U49139 (N_49139,N_43875,N_40271);
nand U49140 (N_49140,N_42050,N_41182);
or U49141 (N_49141,N_42867,N_42174);
and U49142 (N_49142,N_41865,N_43826);
xnor U49143 (N_49143,N_41453,N_41484);
nand U49144 (N_49144,N_44861,N_44791);
nand U49145 (N_49145,N_44855,N_43964);
xnor U49146 (N_49146,N_44432,N_42804);
nand U49147 (N_49147,N_40298,N_42665);
nand U49148 (N_49148,N_40413,N_41506);
or U49149 (N_49149,N_40145,N_44676);
nand U49150 (N_49150,N_40119,N_44365);
nor U49151 (N_49151,N_41212,N_44095);
xnor U49152 (N_49152,N_41461,N_40692);
nor U49153 (N_49153,N_44058,N_43055);
or U49154 (N_49154,N_40052,N_41681);
nand U49155 (N_49155,N_42910,N_40375);
nor U49156 (N_49156,N_41917,N_44684);
xor U49157 (N_49157,N_42769,N_40881);
nand U49158 (N_49158,N_44654,N_40136);
nor U49159 (N_49159,N_43417,N_40843);
nor U49160 (N_49160,N_40919,N_43911);
nand U49161 (N_49161,N_44885,N_40120);
nor U49162 (N_49162,N_41741,N_40824);
and U49163 (N_49163,N_43424,N_44211);
or U49164 (N_49164,N_41545,N_44181);
and U49165 (N_49165,N_44455,N_41119);
and U49166 (N_49166,N_41702,N_42794);
or U49167 (N_49167,N_44459,N_43185);
and U49168 (N_49168,N_42614,N_41910);
xor U49169 (N_49169,N_41258,N_42221);
xnor U49170 (N_49170,N_41287,N_44117);
nand U49171 (N_49171,N_44622,N_44025);
nand U49172 (N_49172,N_42215,N_42168);
nand U49173 (N_49173,N_42282,N_44708);
xnor U49174 (N_49174,N_40744,N_42570);
xnor U49175 (N_49175,N_41309,N_43556);
nor U49176 (N_49176,N_40452,N_42765);
and U49177 (N_49177,N_42412,N_42912);
or U49178 (N_49178,N_43799,N_42626);
nor U49179 (N_49179,N_40293,N_44905);
xnor U49180 (N_49180,N_42133,N_43357);
xor U49181 (N_49181,N_43293,N_42385);
nand U49182 (N_49182,N_43110,N_41577);
and U49183 (N_49183,N_40437,N_40719);
and U49184 (N_49184,N_44930,N_43882);
nand U49185 (N_49185,N_43149,N_42964);
and U49186 (N_49186,N_40151,N_42922);
nand U49187 (N_49187,N_43740,N_41826);
nor U49188 (N_49188,N_40972,N_44376);
or U49189 (N_49189,N_43612,N_40037);
nor U49190 (N_49190,N_44115,N_40257);
or U49191 (N_49191,N_42206,N_43408);
and U49192 (N_49192,N_41418,N_41696);
nand U49193 (N_49193,N_43622,N_44657);
nand U49194 (N_49194,N_43589,N_40988);
and U49195 (N_49195,N_43558,N_43966);
or U49196 (N_49196,N_43586,N_40202);
nand U49197 (N_49197,N_44231,N_42989);
nor U49198 (N_49198,N_44755,N_42145);
and U49199 (N_49199,N_40807,N_41613);
or U49200 (N_49200,N_43410,N_41564);
nor U49201 (N_49201,N_42669,N_44880);
or U49202 (N_49202,N_44582,N_41031);
xnor U49203 (N_49203,N_43584,N_44660);
nor U49204 (N_49204,N_44560,N_43209);
or U49205 (N_49205,N_44777,N_42664);
xnor U49206 (N_49206,N_41127,N_42151);
nand U49207 (N_49207,N_42419,N_43868);
and U49208 (N_49208,N_43031,N_42204);
xnor U49209 (N_49209,N_42212,N_44082);
and U49210 (N_49210,N_42973,N_43851);
nor U49211 (N_49211,N_42188,N_40270);
xnor U49212 (N_49212,N_42306,N_44639);
and U49213 (N_49213,N_43596,N_42972);
nand U49214 (N_49214,N_42820,N_42398);
xor U49215 (N_49215,N_41901,N_43974);
nand U49216 (N_49216,N_42294,N_44134);
xor U49217 (N_49217,N_44525,N_42937);
or U49218 (N_49218,N_43211,N_44652);
or U49219 (N_49219,N_44693,N_41737);
and U49220 (N_49220,N_42509,N_41253);
or U49221 (N_49221,N_41100,N_41236);
or U49222 (N_49222,N_40958,N_41569);
and U49223 (N_49223,N_40928,N_40776);
xor U49224 (N_49224,N_40546,N_43157);
or U49225 (N_49225,N_41791,N_43992);
nor U49226 (N_49226,N_42597,N_42664);
and U49227 (N_49227,N_42676,N_43946);
nand U49228 (N_49228,N_40067,N_42791);
nor U49229 (N_49229,N_44228,N_41038);
nor U49230 (N_49230,N_41806,N_44198);
and U49231 (N_49231,N_41996,N_41864);
and U49232 (N_49232,N_44702,N_40418);
and U49233 (N_49233,N_41337,N_42171);
nor U49234 (N_49234,N_44158,N_42194);
xor U49235 (N_49235,N_42412,N_42677);
xor U49236 (N_49236,N_40957,N_41187);
nand U49237 (N_49237,N_42852,N_40073);
and U49238 (N_49238,N_43228,N_40994);
nor U49239 (N_49239,N_43116,N_42361);
nor U49240 (N_49240,N_40948,N_42526);
nor U49241 (N_49241,N_44161,N_43958);
and U49242 (N_49242,N_42484,N_44451);
nor U49243 (N_49243,N_40620,N_42750);
or U49244 (N_49244,N_40744,N_44646);
and U49245 (N_49245,N_43632,N_40282);
and U49246 (N_49246,N_41544,N_43469);
nand U49247 (N_49247,N_41190,N_40720);
xor U49248 (N_49248,N_42105,N_41923);
xor U49249 (N_49249,N_42685,N_44173);
xor U49250 (N_49250,N_43430,N_40329);
nand U49251 (N_49251,N_40565,N_44580);
xor U49252 (N_49252,N_43543,N_43128);
and U49253 (N_49253,N_41807,N_40619);
nand U49254 (N_49254,N_43386,N_43572);
and U49255 (N_49255,N_44868,N_40000);
xor U49256 (N_49256,N_41608,N_41262);
xnor U49257 (N_49257,N_43459,N_41227);
xnor U49258 (N_49258,N_41717,N_44266);
nor U49259 (N_49259,N_42124,N_44611);
nor U49260 (N_49260,N_40089,N_43368);
nand U49261 (N_49261,N_40842,N_42223);
xor U49262 (N_49262,N_44635,N_42082);
or U49263 (N_49263,N_40429,N_44235);
and U49264 (N_49264,N_42789,N_43956);
nor U49265 (N_49265,N_41662,N_41137);
and U49266 (N_49266,N_41499,N_43752);
xnor U49267 (N_49267,N_43829,N_41007);
or U49268 (N_49268,N_40313,N_42166);
and U49269 (N_49269,N_40206,N_44120);
or U49270 (N_49270,N_42183,N_40312);
or U49271 (N_49271,N_43655,N_42154);
nor U49272 (N_49272,N_42945,N_44813);
nor U49273 (N_49273,N_40343,N_43029);
or U49274 (N_49274,N_40225,N_42009);
xor U49275 (N_49275,N_43100,N_43256);
or U49276 (N_49276,N_43819,N_44719);
xnor U49277 (N_49277,N_41719,N_43833);
xor U49278 (N_49278,N_40491,N_41863);
and U49279 (N_49279,N_43954,N_40234);
xnor U49280 (N_49280,N_44593,N_44473);
or U49281 (N_49281,N_41243,N_43023);
nor U49282 (N_49282,N_42822,N_43307);
or U49283 (N_49283,N_42142,N_42544);
or U49284 (N_49284,N_43503,N_40599);
nor U49285 (N_49285,N_42479,N_42284);
or U49286 (N_49286,N_40642,N_44022);
nand U49287 (N_49287,N_42313,N_42139);
or U49288 (N_49288,N_40353,N_42784);
and U49289 (N_49289,N_42578,N_41034);
nand U49290 (N_49290,N_44670,N_44818);
and U49291 (N_49291,N_42685,N_42230);
and U49292 (N_49292,N_40652,N_44480);
xor U49293 (N_49293,N_41837,N_43785);
and U49294 (N_49294,N_41469,N_40668);
nand U49295 (N_49295,N_42611,N_42190);
nor U49296 (N_49296,N_41627,N_43181);
nand U49297 (N_49297,N_41913,N_44695);
xnor U49298 (N_49298,N_44555,N_42907);
and U49299 (N_49299,N_40675,N_41182);
and U49300 (N_49300,N_42587,N_43076);
nand U49301 (N_49301,N_42496,N_44306);
or U49302 (N_49302,N_40525,N_43940);
nand U49303 (N_49303,N_41248,N_42682);
nand U49304 (N_49304,N_41759,N_42522);
xor U49305 (N_49305,N_44136,N_41995);
nand U49306 (N_49306,N_41983,N_41610);
or U49307 (N_49307,N_41906,N_44381);
or U49308 (N_49308,N_42248,N_44072);
xor U49309 (N_49309,N_44560,N_44236);
xnor U49310 (N_49310,N_41167,N_44836);
or U49311 (N_49311,N_41772,N_41380);
and U49312 (N_49312,N_43587,N_44587);
nor U49313 (N_49313,N_41510,N_44379);
xor U49314 (N_49314,N_42795,N_41194);
or U49315 (N_49315,N_40696,N_43033);
xnor U49316 (N_49316,N_44267,N_41302);
nand U49317 (N_49317,N_44757,N_44807);
or U49318 (N_49318,N_40195,N_40664);
nand U49319 (N_49319,N_41870,N_41435);
xnor U49320 (N_49320,N_40047,N_40070);
and U49321 (N_49321,N_42417,N_42261);
xnor U49322 (N_49322,N_42194,N_42148);
or U49323 (N_49323,N_41339,N_42075);
nand U49324 (N_49324,N_41059,N_40683);
or U49325 (N_49325,N_43395,N_40226);
xnor U49326 (N_49326,N_42363,N_42307);
and U49327 (N_49327,N_40813,N_44829);
xnor U49328 (N_49328,N_43006,N_44063);
nor U49329 (N_49329,N_42574,N_44417);
or U49330 (N_49330,N_42077,N_44554);
nor U49331 (N_49331,N_43572,N_43349);
or U49332 (N_49332,N_42058,N_41468);
nand U49333 (N_49333,N_43966,N_41615);
nor U49334 (N_49334,N_43646,N_44193);
xor U49335 (N_49335,N_41962,N_42460);
nand U49336 (N_49336,N_43684,N_43862);
or U49337 (N_49337,N_41646,N_43746);
nor U49338 (N_49338,N_41336,N_43063);
xor U49339 (N_49339,N_40354,N_41301);
and U49340 (N_49340,N_42790,N_44321);
nor U49341 (N_49341,N_44212,N_40335);
or U49342 (N_49342,N_41451,N_42055);
nand U49343 (N_49343,N_43716,N_40628);
or U49344 (N_49344,N_42667,N_43972);
and U49345 (N_49345,N_42216,N_44771);
and U49346 (N_49346,N_44386,N_40287);
and U49347 (N_49347,N_43636,N_42272);
nor U49348 (N_49348,N_42784,N_40447);
xor U49349 (N_49349,N_44746,N_42588);
and U49350 (N_49350,N_40927,N_44351);
nand U49351 (N_49351,N_40844,N_40925);
or U49352 (N_49352,N_40919,N_44477);
xnor U49353 (N_49353,N_43865,N_42761);
xnor U49354 (N_49354,N_40730,N_44677);
or U49355 (N_49355,N_40754,N_41719);
and U49356 (N_49356,N_43970,N_40470);
or U49357 (N_49357,N_40726,N_44734);
xnor U49358 (N_49358,N_42842,N_42401);
nand U49359 (N_49359,N_42366,N_41635);
or U49360 (N_49360,N_43146,N_43715);
or U49361 (N_49361,N_42825,N_44698);
nand U49362 (N_49362,N_42954,N_43506);
xnor U49363 (N_49363,N_41207,N_42335);
xnor U49364 (N_49364,N_41736,N_42885);
nor U49365 (N_49365,N_42384,N_40632);
xor U49366 (N_49366,N_42409,N_43136);
or U49367 (N_49367,N_44874,N_44388);
nand U49368 (N_49368,N_41230,N_43608);
nand U49369 (N_49369,N_43063,N_44107);
or U49370 (N_49370,N_40250,N_43445);
and U49371 (N_49371,N_41541,N_42883);
and U49372 (N_49372,N_44645,N_42945);
and U49373 (N_49373,N_40155,N_41478);
or U49374 (N_49374,N_44299,N_43893);
nand U49375 (N_49375,N_43642,N_42621);
nand U49376 (N_49376,N_42992,N_43410);
nor U49377 (N_49377,N_43100,N_40540);
nand U49378 (N_49378,N_44425,N_42208);
nand U49379 (N_49379,N_44485,N_44111);
xor U49380 (N_49380,N_41173,N_41877);
nand U49381 (N_49381,N_42501,N_40858);
nand U49382 (N_49382,N_40305,N_41812);
and U49383 (N_49383,N_44753,N_42661);
xnor U49384 (N_49384,N_40597,N_40990);
or U49385 (N_49385,N_42409,N_42808);
nor U49386 (N_49386,N_43563,N_40415);
xor U49387 (N_49387,N_43096,N_43114);
nor U49388 (N_49388,N_42589,N_40909);
and U49389 (N_49389,N_44284,N_40545);
and U49390 (N_49390,N_43728,N_44393);
and U49391 (N_49391,N_40575,N_41882);
and U49392 (N_49392,N_40676,N_42242);
xor U49393 (N_49393,N_42931,N_40249);
and U49394 (N_49394,N_44174,N_43537);
and U49395 (N_49395,N_44955,N_41423);
xor U49396 (N_49396,N_40884,N_41317);
and U49397 (N_49397,N_41843,N_42806);
nor U49398 (N_49398,N_43396,N_41322);
and U49399 (N_49399,N_43379,N_44094);
nand U49400 (N_49400,N_40930,N_40456);
nor U49401 (N_49401,N_43683,N_42383);
and U49402 (N_49402,N_43887,N_41449);
and U49403 (N_49403,N_40359,N_41635);
nor U49404 (N_49404,N_44462,N_40191);
and U49405 (N_49405,N_44065,N_43456);
or U49406 (N_49406,N_43811,N_44402);
nor U49407 (N_49407,N_43668,N_41236);
nand U49408 (N_49408,N_40104,N_40272);
and U49409 (N_49409,N_41974,N_42922);
nor U49410 (N_49410,N_41671,N_41649);
or U49411 (N_49411,N_40619,N_40246);
nand U49412 (N_49412,N_44078,N_40553);
xor U49413 (N_49413,N_41338,N_42968);
nor U49414 (N_49414,N_42715,N_40042);
or U49415 (N_49415,N_42023,N_44354);
and U49416 (N_49416,N_41492,N_40280);
or U49417 (N_49417,N_40000,N_41173);
nor U49418 (N_49418,N_43216,N_40032);
nand U49419 (N_49419,N_41344,N_41492);
xor U49420 (N_49420,N_40089,N_42117);
and U49421 (N_49421,N_41077,N_41278);
nor U49422 (N_49422,N_42206,N_41308);
xor U49423 (N_49423,N_43918,N_40299);
and U49424 (N_49424,N_43648,N_44743);
nand U49425 (N_49425,N_43583,N_42792);
xnor U49426 (N_49426,N_44353,N_43888);
and U49427 (N_49427,N_41894,N_41963);
and U49428 (N_49428,N_44575,N_40177);
and U49429 (N_49429,N_42897,N_43288);
nor U49430 (N_49430,N_42686,N_43472);
xnor U49431 (N_49431,N_44772,N_44963);
xnor U49432 (N_49432,N_42245,N_44819);
nor U49433 (N_49433,N_43935,N_42691);
nor U49434 (N_49434,N_40855,N_43027);
nor U49435 (N_49435,N_42746,N_42516);
and U49436 (N_49436,N_42741,N_43054);
nand U49437 (N_49437,N_40956,N_41118);
nor U49438 (N_49438,N_44354,N_41244);
xnor U49439 (N_49439,N_40798,N_43850);
xor U49440 (N_49440,N_41147,N_40073);
xor U49441 (N_49441,N_41373,N_40247);
xor U49442 (N_49442,N_41559,N_44670);
nor U49443 (N_49443,N_40231,N_44929);
nand U49444 (N_49444,N_40462,N_40088);
and U49445 (N_49445,N_41318,N_41295);
or U49446 (N_49446,N_44113,N_41301);
nor U49447 (N_49447,N_43262,N_41252);
or U49448 (N_49448,N_40215,N_42955);
xnor U49449 (N_49449,N_42075,N_41424);
xor U49450 (N_49450,N_44701,N_41358);
or U49451 (N_49451,N_40538,N_42756);
and U49452 (N_49452,N_41090,N_41907);
xnor U49453 (N_49453,N_42070,N_44371);
nand U49454 (N_49454,N_40067,N_43309);
nand U49455 (N_49455,N_41963,N_44545);
and U49456 (N_49456,N_43475,N_40470);
nor U49457 (N_49457,N_41823,N_41409);
nor U49458 (N_49458,N_41726,N_42902);
xor U49459 (N_49459,N_43531,N_41191);
or U49460 (N_49460,N_40893,N_42241);
and U49461 (N_49461,N_43931,N_43744);
and U49462 (N_49462,N_44577,N_42265);
nor U49463 (N_49463,N_42569,N_42961);
nand U49464 (N_49464,N_40518,N_44483);
and U49465 (N_49465,N_43990,N_44668);
nand U49466 (N_49466,N_44446,N_40021);
nor U49467 (N_49467,N_44730,N_43823);
or U49468 (N_49468,N_42861,N_44329);
xor U49469 (N_49469,N_41824,N_40497);
xor U49470 (N_49470,N_44705,N_42530);
and U49471 (N_49471,N_43461,N_43316);
or U49472 (N_49472,N_41920,N_42382);
xor U49473 (N_49473,N_40668,N_42856);
xor U49474 (N_49474,N_42887,N_40915);
xnor U49475 (N_49475,N_41354,N_42506);
nand U49476 (N_49476,N_40730,N_44084);
nor U49477 (N_49477,N_42032,N_41976);
xor U49478 (N_49478,N_43286,N_44398);
or U49479 (N_49479,N_42874,N_44717);
or U49480 (N_49480,N_42114,N_44771);
xor U49481 (N_49481,N_41121,N_41436);
nor U49482 (N_49482,N_41746,N_43955);
xor U49483 (N_49483,N_40967,N_44115);
and U49484 (N_49484,N_44767,N_43691);
nor U49485 (N_49485,N_40417,N_43520);
or U49486 (N_49486,N_41971,N_40322);
or U49487 (N_49487,N_40633,N_40776);
nor U49488 (N_49488,N_41751,N_40443);
and U49489 (N_49489,N_42863,N_41890);
or U49490 (N_49490,N_41604,N_40006);
nor U49491 (N_49491,N_40610,N_41888);
xor U49492 (N_49492,N_40645,N_41566);
and U49493 (N_49493,N_44148,N_44321);
nor U49494 (N_49494,N_40508,N_40840);
or U49495 (N_49495,N_40285,N_43045);
xor U49496 (N_49496,N_40163,N_40632);
xnor U49497 (N_49497,N_41475,N_41117);
or U49498 (N_49498,N_42238,N_42955);
and U49499 (N_49499,N_43225,N_43817);
and U49500 (N_49500,N_43989,N_44263);
or U49501 (N_49501,N_41178,N_43468);
nor U49502 (N_49502,N_42679,N_42538);
xor U49503 (N_49503,N_41195,N_44361);
xnor U49504 (N_49504,N_43069,N_40394);
and U49505 (N_49505,N_40579,N_42591);
and U49506 (N_49506,N_41658,N_42790);
and U49507 (N_49507,N_41012,N_42668);
or U49508 (N_49508,N_44057,N_42205);
and U49509 (N_49509,N_40280,N_44896);
nor U49510 (N_49510,N_44220,N_44073);
or U49511 (N_49511,N_40866,N_41766);
nand U49512 (N_49512,N_40904,N_42429);
xnor U49513 (N_49513,N_41363,N_40398);
and U49514 (N_49514,N_43450,N_43601);
nand U49515 (N_49515,N_41440,N_41176);
xor U49516 (N_49516,N_42519,N_44205);
nor U49517 (N_49517,N_42006,N_42665);
and U49518 (N_49518,N_43143,N_44963);
nor U49519 (N_49519,N_43313,N_40412);
nor U49520 (N_49520,N_44012,N_44440);
or U49521 (N_49521,N_44781,N_41366);
nor U49522 (N_49522,N_43867,N_41404);
or U49523 (N_49523,N_44377,N_43417);
nor U49524 (N_49524,N_41786,N_43101);
or U49525 (N_49525,N_40821,N_44363);
nor U49526 (N_49526,N_41558,N_42097);
nand U49527 (N_49527,N_41712,N_43443);
and U49528 (N_49528,N_44643,N_43129);
xnor U49529 (N_49529,N_44754,N_44148);
xor U49530 (N_49530,N_42230,N_44513);
and U49531 (N_49531,N_41159,N_40074);
and U49532 (N_49532,N_43442,N_42377);
xnor U49533 (N_49533,N_44512,N_44881);
and U49534 (N_49534,N_41772,N_44847);
nand U49535 (N_49535,N_43663,N_40882);
nor U49536 (N_49536,N_41496,N_44041);
and U49537 (N_49537,N_41559,N_44569);
or U49538 (N_49538,N_41827,N_42506);
xor U49539 (N_49539,N_40093,N_42557);
or U49540 (N_49540,N_40884,N_43729);
and U49541 (N_49541,N_44861,N_43514);
and U49542 (N_49542,N_42096,N_43353);
and U49543 (N_49543,N_43906,N_42925);
nor U49544 (N_49544,N_43639,N_44944);
and U49545 (N_49545,N_43976,N_42316);
and U49546 (N_49546,N_44433,N_40196);
xor U49547 (N_49547,N_40015,N_43262);
xor U49548 (N_49548,N_43326,N_43617);
nor U49549 (N_49549,N_42031,N_40462);
and U49550 (N_49550,N_41540,N_42420);
xnor U49551 (N_49551,N_44028,N_42452);
xnor U49552 (N_49552,N_40238,N_41036);
nor U49553 (N_49553,N_40836,N_41276);
nand U49554 (N_49554,N_43470,N_41516);
or U49555 (N_49555,N_42933,N_42244);
nand U49556 (N_49556,N_42810,N_42258);
nor U49557 (N_49557,N_41663,N_42762);
nand U49558 (N_49558,N_42705,N_43051);
or U49559 (N_49559,N_43181,N_43670);
or U49560 (N_49560,N_44844,N_43513);
nand U49561 (N_49561,N_40115,N_41808);
nor U49562 (N_49562,N_41470,N_40849);
and U49563 (N_49563,N_40844,N_43737);
and U49564 (N_49564,N_43480,N_43109);
nor U49565 (N_49565,N_44896,N_40647);
nand U49566 (N_49566,N_40188,N_44887);
and U49567 (N_49567,N_41439,N_40220);
xnor U49568 (N_49568,N_44621,N_44348);
xnor U49569 (N_49569,N_40852,N_43175);
or U49570 (N_49570,N_40175,N_40375);
or U49571 (N_49571,N_41335,N_41219);
xnor U49572 (N_49572,N_41842,N_44106);
nor U49573 (N_49573,N_44524,N_42048);
or U49574 (N_49574,N_40326,N_40190);
nor U49575 (N_49575,N_40999,N_43369);
nand U49576 (N_49576,N_42547,N_41776);
nor U49577 (N_49577,N_44511,N_43953);
or U49578 (N_49578,N_40974,N_41558);
xnor U49579 (N_49579,N_43741,N_42330);
xor U49580 (N_49580,N_40308,N_42755);
nor U49581 (N_49581,N_41972,N_42239);
xnor U49582 (N_49582,N_41240,N_42245);
nand U49583 (N_49583,N_43321,N_42172);
xnor U49584 (N_49584,N_44846,N_44915);
and U49585 (N_49585,N_43426,N_41468);
or U49586 (N_49586,N_43056,N_41923);
nand U49587 (N_49587,N_40189,N_40951);
nand U49588 (N_49588,N_40488,N_40136);
xnor U49589 (N_49589,N_44440,N_41050);
xnor U49590 (N_49590,N_41254,N_44563);
nor U49591 (N_49591,N_44504,N_43051);
or U49592 (N_49592,N_40492,N_43647);
or U49593 (N_49593,N_40074,N_44456);
xnor U49594 (N_49594,N_42378,N_41778);
nor U49595 (N_49595,N_42766,N_44142);
or U49596 (N_49596,N_40448,N_44386);
and U49597 (N_49597,N_40609,N_40182);
and U49598 (N_49598,N_41854,N_42842);
nor U49599 (N_49599,N_41730,N_43930);
and U49600 (N_49600,N_41677,N_41421);
or U49601 (N_49601,N_40726,N_44572);
nand U49602 (N_49602,N_40030,N_44696);
and U49603 (N_49603,N_44842,N_44833);
or U49604 (N_49604,N_43515,N_43376);
nand U49605 (N_49605,N_41173,N_44778);
nor U49606 (N_49606,N_40383,N_44126);
nor U49607 (N_49607,N_43160,N_40678);
nand U49608 (N_49608,N_41110,N_44600);
nor U49609 (N_49609,N_42286,N_43642);
or U49610 (N_49610,N_43829,N_41880);
nand U49611 (N_49611,N_43890,N_43330);
xor U49612 (N_49612,N_43168,N_44815);
nand U49613 (N_49613,N_44065,N_44854);
or U49614 (N_49614,N_42503,N_41307);
nand U49615 (N_49615,N_43975,N_40940);
nor U49616 (N_49616,N_42621,N_40984);
or U49617 (N_49617,N_40913,N_43974);
nor U49618 (N_49618,N_42260,N_44681);
nor U49619 (N_49619,N_44143,N_43735);
xor U49620 (N_49620,N_42920,N_42115);
nand U49621 (N_49621,N_43942,N_40974);
nand U49622 (N_49622,N_42940,N_40693);
xnor U49623 (N_49623,N_40819,N_42892);
xor U49624 (N_49624,N_43411,N_41529);
xor U49625 (N_49625,N_42690,N_41123);
nor U49626 (N_49626,N_41793,N_40049);
nor U49627 (N_49627,N_42043,N_40037);
xnor U49628 (N_49628,N_44486,N_42555);
xor U49629 (N_49629,N_40814,N_40166);
or U49630 (N_49630,N_42505,N_41128);
or U49631 (N_49631,N_43099,N_44961);
xor U49632 (N_49632,N_43428,N_44426);
and U49633 (N_49633,N_43635,N_40454);
xnor U49634 (N_49634,N_42768,N_42660);
nand U49635 (N_49635,N_41668,N_42504);
nor U49636 (N_49636,N_43573,N_43665);
nor U49637 (N_49637,N_43390,N_41461);
nor U49638 (N_49638,N_43639,N_42239);
or U49639 (N_49639,N_43879,N_43731);
nor U49640 (N_49640,N_43415,N_42855);
xnor U49641 (N_49641,N_41828,N_40803);
or U49642 (N_49642,N_42045,N_43838);
or U49643 (N_49643,N_44076,N_44589);
or U49644 (N_49644,N_41290,N_40810);
and U49645 (N_49645,N_42046,N_43372);
or U49646 (N_49646,N_41781,N_43941);
or U49647 (N_49647,N_44900,N_44216);
or U49648 (N_49648,N_42207,N_40108);
and U49649 (N_49649,N_43392,N_44220);
or U49650 (N_49650,N_40594,N_43021);
nor U49651 (N_49651,N_40411,N_44507);
xor U49652 (N_49652,N_43803,N_44030);
xnor U49653 (N_49653,N_44738,N_43965);
nor U49654 (N_49654,N_41363,N_40053);
nor U49655 (N_49655,N_40206,N_43843);
and U49656 (N_49656,N_40585,N_43648);
xnor U49657 (N_49657,N_43311,N_43163);
and U49658 (N_49658,N_43551,N_40958);
and U49659 (N_49659,N_42859,N_42303);
and U49660 (N_49660,N_40080,N_43630);
and U49661 (N_49661,N_44901,N_41252);
or U49662 (N_49662,N_44481,N_42541);
nor U49663 (N_49663,N_41365,N_41537);
and U49664 (N_49664,N_42854,N_42086);
xnor U49665 (N_49665,N_44482,N_44625);
xor U49666 (N_49666,N_43396,N_44617);
xnor U49667 (N_49667,N_44292,N_43721);
xnor U49668 (N_49668,N_42320,N_44221);
xnor U49669 (N_49669,N_44924,N_43682);
nor U49670 (N_49670,N_41493,N_41430);
and U49671 (N_49671,N_42487,N_41072);
nor U49672 (N_49672,N_42758,N_40236);
xor U49673 (N_49673,N_43457,N_41332);
or U49674 (N_49674,N_44740,N_42998);
or U49675 (N_49675,N_40460,N_43648);
or U49676 (N_49676,N_43204,N_42616);
nand U49677 (N_49677,N_41647,N_43765);
nor U49678 (N_49678,N_41790,N_43534);
xnor U49679 (N_49679,N_40719,N_40030);
and U49680 (N_49680,N_42919,N_41628);
and U49681 (N_49681,N_44426,N_43301);
xnor U49682 (N_49682,N_43390,N_41761);
nor U49683 (N_49683,N_44491,N_43839);
xnor U49684 (N_49684,N_44648,N_41953);
or U49685 (N_49685,N_43221,N_40689);
or U49686 (N_49686,N_43057,N_42481);
xnor U49687 (N_49687,N_42889,N_42823);
nand U49688 (N_49688,N_44184,N_42188);
xnor U49689 (N_49689,N_44677,N_44025);
xnor U49690 (N_49690,N_41826,N_40795);
nand U49691 (N_49691,N_42978,N_42506);
nor U49692 (N_49692,N_44318,N_44674);
nand U49693 (N_49693,N_41130,N_44091);
xnor U49694 (N_49694,N_41359,N_43492);
nor U49695 (N_49695,N_40000,N_44350);
nor U49696 (N_49696,N_44574,N_41217);
and U49697 (N_49697,N_44349,N_42339);
xor U49698 (N_49698,N_44253,N_43613);
or U49699 (N_49699,N_44496,N_43134);
or U49700 (N_49700,N_44259,N_42871);
nor U49701 (N_49701,N_44920,N_43239);
and U49702 (N_49702,N_40246,N_43740);
or U49703 (N_49703,N_42681,N_43924);
nor U49704 (N_49704,N_43744,N_44823);
nor U49705 (N_49705,N_44012,N_41820);
and U49706 (N_49706,N_43842,N_40242);
nor U49707 (N_49707,N_40504,N_43758);
and U49708 (N_49708,N_40865,N_42802);
xor U49709 (N_49709,N_40992,N_40401);
nand U49710 (N_49710,N_42189,N_42465);
nor U49711 (N_49711,N_42005,N_41997);
and U49712 (N_49712,N_42658,N_41123);
and U49713 (N_49713,N_41438,N_42289);
and U49714 (N_49714,N_44091,N_41469);
or U49715 (N_49715,N_42628,N_41175);
xor U49716 (N_49716,N_41705,N_41234);
xor U49717 (N_49717,N_41432,N_40388);
or U49718 (N_49718,N_40590,N_40491);
nand U49719 (N_49719,N_42332,N_40533);
or U49720 (N_49720,N_42208,N_41250);
nor U49721 (N_49721,N_41426,N_42962);
and U49722 (N_49722,N_42363,N_44314);
or U49723 (N_49723,N_41580,N_40529);
xnor U49724 (N_49724,N_43622,N_41718);
xor U49725 (N_49725,N_42129,N_42702);
xor U49726 (N_49726,N_41724,N_44548);
and U49727 (N_49727,N_42916,N_40881);
or U49728 (N_49728,N_44816,N_43829);
or U49729 (N_49729,N_43977,N_43029);
nand U49730 (N_49730,N_44329,N_42004);
nor U49731 (N_49731,N_44959,N_43631);
and U49732 (N_49732,N_44058,N_41597);
xnor U49733 (N_49733,N_44520,N_42000);
nand U49734 (N_49734,N_42276,N_44293);
and U49735 (N_49735,N_43841,N_42055);
xnor U49736 (N_49736,N_41260,N_42584);
nor U49737 (N_49737,N_42584,N_43350);
and U49738 (N_49738,N_40517,N_40475);
or U49739 (N_49739,N_44185,N_43758);
xor U49740 (N_49740,N_44160,N_42176);
nor U49741 (N_49741,N_42163,N_40279);
xor U49742 (N_49742,N_40262,N_42602);
or U49743 (N_49743,N_41161,N_40918);
nand U49744 (N_49744,N_41769,N_41311);
and U49745 (N_49745,N_41986,N_42162);
nor U49746 (N_49746,N_44785,N_42834);
or U49747 (N_49747,N_40012,N_42581);
xnor U49748 (N_49748,N_44940,N_42671);
and U49749 (N_49749,N_43260,N_40641);
or U49750 (N_49750,N_43459,N_41507);
xnor U49751 (N_49751,N_41545,N_40697);
nand U49752 (N_49752,N_43922,N_40485);
nor U49753 (N_49753,N_41472,N_42779);
and U49754 (N_49754,N_43846,N_43563);
or U49755 (N_49755,N_41725,N_43230);
xnor U49756 (N_49756,N_44276,N_42376);
nand U49757 (N_49757,N_40434,N_44953);
nand U49758 (N_49758,N_41171,N_41360);
xnor U49759 (N_49759,N_42791,N_42819);
nand U49760 (N_49760,N_42419,N_40682);
xnor U49761 (N_49761,N_41685,N_40644);
or U49762 (N_49762,N_40967,N_42812);
nor U49763 (N_49763,N_40114,N_42925);
xnor U49764 (N_49764,N_41686,N_42863);
or U49765 (N_49765,N_40684,N_40973);
or U49766 (N_49766,N_40542,N_41404);
xor U49767 (N_49767,N_42673,N_40351);
or U49768 (N_49768,N_41899,N_40772);
or U49769 (N_49769,N_44415,N_44535);
xnor U49770 (N_49770,N_43006,N_41040);
or U49771 (N_49771,N_43744,N_41847);
nor U49772 (N_49772,N_41486,N_40632);
xnor U49773 (N_49773,N_40328,N_44813);
and U49774 (N_49774,N_42014,N_44642);
nand U49775 (N_49775,N_43124,N_43422);
xor U49776 (N_49776,N_44289,N_40135);
nor U49777 (N_49777,N_44859,N_44066);
nor U49778 (N_49778,N_44303,N_42530);
and U49779 (N_49779,N_41145,N_42880);
and U49780 (N_49780,N_41441,N_44076);
nor U49781 (N_49781,N_42626,N_44381);
and U49782 (N_49782,N_42796,N_44971);
nand U49783 (N_49783,N_42813,N_40023);
nor U49784 (N_49784,N_40867,N_41448);
or U49785 (N_49785,N_43678,N_42099);
or U49786 (N_49786,N_44356,N_41115);
and U49787 (N_49787,N_42528,N_41860);
nor U49788 (N_49788,N_41632,N_44052);
and U49789 (N_49789,N_41611,N_40568);
and U49790 (N_49790,N_40081,N_44517);
nor U49791 (N_49791,N_44685,N_44734);
and U49792 (N_49792,N_42651,N_41670);
nand U49793 (N_49793,N_43364,N_43131);
xnor U49794 (N_49794,N_41880,N_44911);
or U49795 (N_49795,N_42041,N_44430);
xor U49796 (N_49796,N_44360,N_42509);
or U49797 (N_49797,N_44783,N_44295);
nand U49798 (N_49798,N_41776,N_41720);
or U49799 (N_49799,N_41019,N_43967);
or U49800 (N_49800,N_42861,N_43480);
nand U49801 (N_49801,N_40548,N_40504);
and U49802 (N_49802,N_41263,N_43045);
and U49803 (N_49803,N_41731,N_44591);
and U49804 (N_49804,N_40945,N_42010);
or U49805 (N_49805,N_41966,N_41250);
xor U49806 (N_49806,N_43120,N_43426);
or U49807 (N_49807,N_40068,N_43983);
and U49808 (N_49808,N_41123,N_40922);
xnor U49809 (N_49809,N_43221,N_42213);
xnor U49810 (N_49810,N_40638,N_42344);
and U49811 (N_49811,N_42499,N_44985);
and U49812 (N_49812,N_40210,N_40039);
xnor U49813 (N_49813,N_40211,N_41907);
nand U49814 (N_49814,N_41815,N_40700);
xor U49815 (N_49815,N_42657,N_40499);
nand U49816 (N_49816,N_40089,N_44531);
or U49817 (N_49817,N_42497,N_44931);
and U49818 (N_49818,N_41237,N_41578);
xor U49819 (N_49819,N_42489,N_44767);
or U49820 (N_49820,N_44395,N_40522);
xor U49821 (N_49821,N_44592,N_42728);
and U49822 (N_49822,N_40908,N_40349);
nor U49823 (N_49823,N_40747,N_41827);
nand U49824 (N_49824,N_42769,N_43169);
nor U49825 (N_49825,N_41580,N_43492);
nor U49826 (N_49826,N_43610,N_44791);
nor U49827 (N_49827,N_40158,N_44495);
nand U49828 (N_49828,N_43633,N_43878);
nand U49829 (N_49829,N_42158,N_42665);
xor U49830 (N_49830,N_43780,N_41236);
nor U49831 (N_49831,N_43063,N_44630);
and U49832 (N_49832,N_40915,N_41702);
or U49833 (N_49833,N_40783,N_43100);
nand U49834 (N_49834,N_44572,N_40779);
nor U49835 (N_49835,N_43679,N_41865);
and U49836 (N_49836,N_40303,N_43903);
xnor U49837 (N_49837,N_42707,N_43966);
or U49838 (N_49838,N_43995,N_40166);
or U49839 (N_49839,N_40529,N_40391);
or U49840 (N_49840,N_41272,N_42809);
nand U49841 (N_49841,N_42246,N_42716);
nor U49842 (N_49842,N_42426,N_44709);
and U49843 (N_49843,N_43264,N_42014);
or U49844 (N_49844,N_42665,N_43583);
xor U49845 (N_49845,N_44902,N_43114);
xor U49846 (N_49846,N_42377,N_40930);
or U49847 (N_49847,N_40398,N_43121);
nand U49848 (N_49848,N_40834,N_42728);
nand U49849 (N_49849,N_44372,N_41747);
and U49850 (N_49850,N_44637,N_43854);
or U49851 (N_49851,N_40763,N_42444);
nor U49852 (N_49852,N_42232,N_43086);
nand U49853 (N_49853,N_41255,N_43444);
nand U49854 (N_49854,N_44728,N_41773);
and U49855 (N_49855,N_40256,N_42495);
or U49856 (N_49856,N_42369,N_41973);
and U49857 (N_49857,N_44834,N_42502);
nor U49858 (N_49858,N_43095,N_43177);
or U49859 (N_49859,N_43686,N_42021);
nand U49860 (N_49860,N_42234,N_42734);
nand U49861 (N_49861,N_44318,N_40757);
xor U49862 (N_49862,N_40682,N_41123);
and U49863 (N_49863,N_41291,N_44982);
or U49864 (N_49864,N_41230,N_40688);
xnor U49865 (N_49865,N_41596,N_41138);
and U49866 (N_49866,N_41096,N_40518);
nor U49867 (N_49867,N_40459,N_43194);
nand U49868 (N_49868,N_41811,N_44373);
xor U49869 (N_49869,N_40905,N_44596);
nor U49870 (N_49870,N_44883,N_43263);
nor U49871 (N_49871,N_41132,N_44589);
and U49872 (N_49872,N_44272,N_41524);
nand U49873 (N_49873,N_44344,N_40961);
xor U49874 (N_49874,N_44224,N_43461);
nand U49875 (N_49875,N_41505,N_40331);
xnor U49876 (N_49876,N_44526,N_41079);
or U49877 (N_49877,N_40035,N_40877);
xnor U49878 (N_49878,N_41646,N_42997);
nand U49879 (N_49879,N_44784,N_43221);
nor U49880 (N_49880,N_41489,N_40450);
nand U49881 (N_49881,N_41521,N_44519);
or U49882 (N_49882,N_41032,N_40984);
nand U49883 (N_49883,N_41853,N_41503);
nand U49884 (N_49884,N_43295,N_41083);
or U49885 (N_49885,N_42168,N_41355);
xor U49886 (N_49886,N_42846,N_41646);
nand U49887 (N_49887,N_40496,N_44126);
nand U49888 (N_49888,N_43620,N_43912);
nor U49889 (N_49889,N_42392,N_43363);
and U49890 (N_49890,N_41507,N_40811);
nand U49891 (N_49891,N_42549,N_41415);
and U49892 (N_49892,N_43554,N_42465);
xnor U49893 (N_49893,N_40017,N_40521);
nand U49894 (N_49894,N_40824,N_42015);
and U49895 (N_49895,N_43349,N_44270);
and U49896 (N_49896,N_41853,N_40988);
xnor U49897 (N_49897,N_41695,N_40983);
or U49898 (N_49898,N_44637,N_44636);
xnor U49899 (N_49899,N_43313,N_44827);
xnor U49900 (N_49900,N_41478,N_41717);
or U49901 (N_49901,N_41659,N_43522);
xor U49902 (N_49902,N_40667,N_40404);
or U49903 (N_49903,N_41481,N_42101);
nor U49904 (N_49904,N_43329,N_44491);
nand U49905 (N_49905,N_42506,N_43357);
nand U49906 (N_49906,N_43582,N_44318);
or U49907 (N_49907,N_43154,N_44679);
nand U49908 (N_49908,N_42373,N_43902);
xnor U49909 (N_49909,N_40021,N_43592);
nand U49910 (N_49910,N_43614,N_43929);
xnor U49911 (N_49911,N_40466,N_43285);
or U49912 (N_49912,N_44500,N_42834);
nand U49913 (N_49913,N_44926,N_43485);
and U49914 (N_49914,N_44084,N_43916);
nand U49915 (N_49915,N_42947,N_40981);
nand U49916 (N_49916,N_41489,N_43019);
and U49917 (N_49917,N_44389,N_42809);
nor U49918 (N_49918,N_43633,N_41682);
and U49919 (N_49919,N_42715,N_41715);
nand U49920 (N_49920,N_41425,N_43557);
and U49921 (N_49921,N_41112,N_42705);
and U49922 (N_49922,N_40970,N_40261);
nor U49923 (N_49923,N_42660,N_41778);
and U49924 (N_49924,N_41323,N_40214);
nor U49925 (N_49925,N_40981,N_44551);
xnor U49926 (N_49926,N_43857,N_40177);
nor U49927 (N_49927,N_42233,N_42421);
and U49928 (N_49928,N_40146,N_44868);
xnor U49929 (N_49929,N_40144,N_40459);
nand U49930 (N_49930,N_42717,N_43137);
xnor U49931 (N_49931,N_41703,N_40112);
nand U49932 (N_49932,N_42369,N_43765);
nor U49933 (N_49933,N_41594,N_43615);
xnor U49934 (N_49934,N_44537,N_41384);
nor U49935 (N_49935,N_43902,N_42748);
and U49936 (N_49936,N_44879,N_41674);
xor U49937 (N_49937,N_44210,N_43998);
xor U49938 (N_49938,N_41442,N_41979);
nor U49939 (N_49939,N_42277,N_42887);
xor U49940 (N_49940,N_41000,N_41650);
or U49941 (N_49941,N_42485,N_40121);
xor U49942 (N_49942,N_44101,N_44592);
nor U49943 (N_49943,N_41889,N_40341);
or U49944 (N_49944,N_40472,N_43512);
or U49945 (N_49945,N_40196,N_42009);
xnor U49946 (N_49946,N_41869,N_44572);
nor U49947 (N_49947,N_42942,N_42279);
nor U49948 (N_49948,N_44236,N_41331);
and U49949 (N_49949,N_40518,N_43221);
or U49950 (N_49950,N_41215,N_42319);
xnor U49951 (N_49951,N_43781,N_44403);
nand U49952 (N_49952,N_43278,N_40452);
xnor U49953 (N_49953,N_41036,N_43559);
nand U49954 (N_49954,N_40733,N_42192);
xnor U49955 (N_49955,N_44767,N_40230);
nand U49956 (N_49956,N_43493,N_43531);
nand U49957 (N_49957,N_44232,N_41958);
xor U49958 (N_49958,N_41926,N_40465);
nand U49959 (N_49959,N_40453,N_40773);
and U49960 (N_49960,N_42742,N_42708);
nor U49961 (N_49961,N_44645,N_42674);
or U49962 (N_49962,N_40163,N_42613);
nand U49963 (N_49963,N_43463,N_43428);
or U49964 (N_49964,N_43864,N_42244);
or U49965 (N_49965,N_44339,N_40745);
nand U49966 (N_49966,N_41187,N_42768);
and U49967 (N_49967,N_42133,N_41504);
or U49968 (N_49968,N_43498,N_42091);
nor U49969 (N_49969,N_41774,N_43541);
nand U49970 (N_49970,N_41285,N_42315);
or U49971 (N_49971,N_44913,N_41665);
nand U49972 (N_49972,N_40460,N_42111);
nor U49973 (N_49973,N_40525,N_40753);
and U49974 (N_49974,N_43269,N_40904);
nand U49975 (N_49975,N_44249,N_43125);
and U49976 (N_49976,N_42287,N_41175);
and U49977 (N_49977,N_42819,N_41061);
and U49978 (N_49978,N_41662,N_43672);
and U49979 (N_49979,N_44867,N_41526);
and U49980 (N_49980,N_44484,N_40324);
nor U49981 (N_49981,N_42848,N_43034);
and U49982 (N_49982,N_40054,N_44913);
nand U49983 (N_49983,N_43926,N_44270);
nor U49984 (N_49984,N_43398,N_41502);
nor U49985 (N_49985,N_44759,N_44465);
and U49986 (N_49986,N_43453,N_40559);
or U49987 (N_49987,N_40304,N_40860);
nor U49988 (N_49988,N_40423,N_43720);
and U49989 (N_49989,N_42978,N_41175);
xor U49990 (N_49990,N_41137,N_41954);
xor U49991 (N_49991,N_43379,N_44964);
nand U49992 (N_49992,N_44704,N_43112);
xor U49993 (N_49993,N_44461,N_41104);
nor U49994 (N_49994,N_43311,N_43513);
nand U49995 (N_49995,N_41023,N_43997);
nand U49996 (N_49996,N_41873,N_44707);
xnor U49997 (N_49997,N_41197,N_43140);
or U49998 (N_49998,N_40619,N_40965);
or U49999 (N_49999,N_42084,N_40861);
xor UO_0 (O_0,N_48327,N_47720);
or UO_1 (O_1,N_48521,N_47691);
nand UO_2 (O_2,N_45374,N_47578);
nor UO_3 (O_3,N_46768,N_46374);
xnor UO_4 (O_4,N_47853,N_45958);
xor UO_5 (O_5,N_48466,N_48787);
and UO_6 (O_6,N_47625,N_46359);
nand UO_7 (O_7,N_49239,N_46088);
or UO_8 (O_8,N_46093,N_45188);
or UO_9 (O_9,N_46746,N_45388);
nand UO_10 (O_10,N_45887,N_46355);
and UO_11 (O_11,N_45215,N_49347);
or UO_12 (O_12,N_45957,N_45244);
nor UO_13 (O_13,N_49204,N_45598);
xnor UO_14 (O_14,N_46849,N_49783);
xnor UO_15 (O_15,N_49839,N_46685);
xor UO_16 (O_16,N_46323,N_45753);
and UO_17 (O_17,N_46999,N_45892);
or UO_18 (O_18,N_48049,N_46959);
nor UO_19 (O_19,N_49006,N_45610);
or UO_20 (O_20,N_48695,N_47709);
nand UO_21 (O_21,N_45804,N_49688);
nor UO_22 (O_22,N_48829,N_48050);
nor UO_23 (O_23,N_45168,N_45255);
nor UO_24 (O_24,N_47995,N_48441);
nand UO_25 (O_25,N_46402,N_48813);
xor UO_26 (O_26,N_46405,N_47759);
xor UO_27 (O_27,N_48150,N_46448);
nor UO_28 (O_28,N_48863,N_46618);
xnor UO_29 (O_29,N_48627,N_48825);
and UO_30 (O_30,N_48751,N_47550);
xor UO_31 (O_31,N_49231,N_49293);
and UO_32 (O_32,N_49853,N_47809);
and UO_33 (O_33,N_48922,N_48262);
or UO_34 (O_34,N_47114,N_49241);
and UO_35 (O_35,N_48473,N_46884);
nor UO_36 (O_36,N_47538,N_46026);
or UO_37 (O_37,N_47074,N_49663);
nor UO_38 (O_38,N_48181,N_46115);
nand UO_39 (O_39,N_46923,N_49801);
nand UO_40 (O_40,N_46868,N_48556);
or UO_41 (O_41,N_49185,N_47327);
xnor UO_42 (O_42,N_49812,N_46726);
nand UO_43 (O_43,N_47476,N_49966);
nor UO_44 (O_44,N_46032,N_48896);
or UO_45 (O_45,N_49072,N_46737);
nand UO_46 (O_46,N_45888,N_49898);
or UO_47 (O_47,N_48294,N_46406);
or UO_48 (O_48,N_49904,N_49828);
nand UO_49 (O_49,N_45127,N_47480);
or UO_50 (O_50,N_49809,N_45770);
xor UO_51 (O_51,N_48229,N_46392);
or UO_52 (O_52,N_46921,N_48638);
or UO_53 (O_53,N_45429,N_49226);
nand UO_54 (O_54,N_46476,N_49404);
nor UO_55 (O_55,N_45692,N_46681);
nor UO_56 (O_56,N_48918,N_47879);
nand UO_57 (O_57,N_46461,N_48725);
and UO_58 (O_58,N_48457,N_47167);
or UO_59 (O_59,N_47004,N_45291);
nor UO_60 (O_60,N_47278,N_45984);
and UO_61 (O_61,N_46502,N_46544);
or UO_62 (O_62,N_49880,N_45752);
nor UO_63 (O_63,N_46975,N_46471);
or UO_64 (O_64,N_45740,N_46964);
nor UO_65 (O_65,N_49830,N_48368);
nand UO_66 (O_66,N_48405,N_48789);
nor UO_67 (O_67,N_48092,N_49013);
nor UO_68 (O_68,N_46809,N_46022);
and UO_69 (O_69,N_46435,N_46409);
and UO_70 (O_70,N_45851,N_49427);
nor UO_71 (O_71,N_47151,N_48268);
and UO_72 (O_72,N_45746,N_46066);
nor UO_73 (O_73,N_48464,N_45696);
xor UO_74 (O_74,N_48595,N_48481);
xnor UO_75 (O_75,N_48082,N_47650);
nor UO_76 (O_76,N_45924,N_46839);
and UO_77 (O_77,N_48037,N_45226);
xor UO_78 (O_78,N_49494,N_48867);
nor UO_79 (O_79,N_47745,N_45102);
nand UO_80 (O_80,N_45698,N_49713);
xor UO_81 (O_81,N_49129,N_48520);
or UO_82 (O_82,N_46492,N_45400);
xnor UO_83 (O_83,N_47039,N_46134);
xor UO_84 (O_84,N_47147,N_48646);
and UO_85 (O_85,N_48242,N_46948);
or UO_86 (O_86,N_46527,N_49173);
nor UO_87 (O_87,N_49701,N_47865);
nand UO_88 (O_88,N_49351,N_47703);
or UO_89 (O_89,N_48865,N_45837);
nand UO_90 (O_90,N_46697,N_49510);
nand UO_91 (O_91,N_49018,N_46947);
or UO_92 (O_92,N_48802,N_45196);
and UO_93 (O_93,N_47839,N_46447);
xnor UO_94 (O_94,N_49782,N_45259);
xor UO_95 (O_95,N_47467,N_49138);
and UO_96 (O_96,N_49375,N_49338);
nor UO_97 (O_97,N_46802,N_49779);
and UO_98 (O_98,N_48586,N_46113);
or UO_99 (O_99,N_45749,N_48764);
and UO_100 (O_100,N_49998,N_48271);
xor UO_101 (O_101,N_45541,N_47051);
nor UO_102 (O_102,N_47938,N_47402);
nand UO_103 (O_103,N_46514,N_47153);
nand UO_104 (O_104,N_46387,N_45809);
or UO_105 (O_105,N_47831,N_45287);
nor UO_106 (O_106,N_46680,N_47693);
nor UO_107 (O_107,N_48056,N_47719);
nand UO_108 (O_108,N_49551,N_45985);
and UO_109 (O_109,N_45395,N_46765);
and UO_110 (O_110,N_49340,N_47682);
nand UO_111 (O_111,N_46031,N_49916);
xnor UO_112 (O_112,N_49408,N_45830);
and UO_113 (O_113,N_46158,N_47785);
nor UO_114 (O_114,N_47953,N_49610);
nand UO_115 (O_115,N_46004,N_45921);
nor UO_116 (O_116,N_45640,N_47350);
nor UO_117 (O_117,N_46587,N_46952);
and UO_118 (O_118,N_45626,N_46080);
and UO_119 (O_119,N_48533,N_49482);
xnor UO_120 (O_120,N_46375,N_45040);
or UO_121 (O_121,N_46485,N_45021);
or UO_122 (O_122,N_49110,N_46979);
nand UO_123 (O_123,N_48276,N_45849);
xor UO_124 (O_124,N_47450,N_49332);
or UO_125 (O_125,N_49977,N_48618);
nand UO_126 (O_126,N_48354,N_48172);
xnor UO_127 (O_127,N_46752,N_49012);
nor UO_128 (O_128,N_46208,N_49039);
or UO_129 (O_129,N_48084,N_48514);
and UO_130 (O_130,N_47374,N_49542);
or UO_131 (O_131,N_49745,N_46102);
and UO_132 (O_132,N_47069,N_49169);
or UO_133 (O_133,N_45633,N_49228);
nand UO_134 (O_134,N_49974,N_49209);
xor UO_135 (O_135,N_46459,N_45185);
nand UO_136 (O_136,N_47415,N_47394);
and UO_137 (O_137,N_45258,N_47800);
xor UO_138 (O_138,N_45150,N_49448);
xnor UO_139 (O_139,N_47133,N_46248);
nor UO_140 (O_140,N_45909,N_45221);
or UO_141 (O_141,N_47332,N_46638);
nor UO_142 (O_142,N_46062,N_46785);
xnor UO_143 (O_143,N_46846,N_45109);
or UO_144 (O_144,N_46559,N_46541);
xor UO_145 (O_145,N_48509,N_48781);
and UO_146 (O_146,N_47873,N_46749);
nor UO_147 (O_147,N_48486,N_48662);
xnor UO_148 (O_148,N_49456,N_47922);
and UO_149 (O_149,N_46524,N_45392);
nor UO_150 (O_150,N_48002,N_48409);
nor UO_151 (O_151,N_48253,N_45889);
or UO_152 (O_152,N_49207,N_46076);
nor UO_153 (O_153,N_48961,N_47209);
nand UO_154 (O_154,N_47200,N_48610);
and UO_155 (O_155,N_49492,N_45521);
nand UO_156 (O_156,N_47213,N_46327);
and UO_157 (O_157,N_47508,N_47985);
and UO_158 (O_158,N_46647,N_46424);
xor UO_159 (O_159,N_45882,N_48573);
or UO_160 (O_160,N_49704,N_49754);
nand UO_161 (O_161,N_46596,N_48012);
and UO_162 (O_162,N_45209,N_47105);
nand UO_163 (O_163,N_48142,N_49158);
xor UO_164 (O_164,N_48542,N_46482);
nor UO_165 (O_165,N_46187,N_49706);
nor UO_166 (O_166,N_46859,N_45016);
or UO_167 (O_167,N_45760,N_48946);
nand UO_168 (O_168,N_47637,N_48782);
nand UO_169 (O_169,N_47596,N_45603);
nand UO_170 (O_170,N_45950,N_46018);
or UO_171 (O_171,N_47523,N_46404);
nand UO_172 (O_172,N_45754,N_46938);
xor UO_173 (O_173,N_45588,N_49046);
nor UO_174 (O_174,N_47323,N_49439);
or UO_175 (O_175,N_49937,N_49826);
nand UO_176 (O_176,N_47351,N_46108);
or UO_177 (O_177,N_45213,N_47822);
nor UO_178 (O_178,N_48231,N_45801);
nor UO_179 (O_179,N_46816,N_45101);
nor UO_180 (O_180,N_46757,N_49210);
nor UO_181 (O_181,N_45234,N_46799);
and UO_182 (O_182,N_48733,N_48664);
nand UO_183 (O_183,N_46645,N_49134);
nand UO_184 (O_184,N_49443,N_46515);
or UO_185 (O_185,N_46168,N_47748);
nand UO_186 (O_186,N_45207,N_45995);
xor UO_187 (O_187,N_48888,N_47806);
or UO_188 (O_188,N_47068,N_49617);
nor UO_189 (O_189,N_47072,N_45657);
nor UO_190 (O_190,N_49846,N_48046);
or UO_191 (O_191,N_48184,N_45805);
and UO_192 (O_192,N_48830,N_49768);
and UO_193 (O_193,N_46038,N_48552);
nand UO_194 (O_194,N_48298,N_47718);
nor UO_195 (O_195,N_49983,N_49730);
nand UO_196 (O_196,N_48728,N_46727);
and UO_197 (O_197,N_48854,N_45852);
or UO_198 (O_198,N_45261,N_46972);
nor UO_199 (O_199,N_47867,N_45061);
and UO_200 (O_200,N_49376,N_46543);
and UO_201 (O_201,N_47882,N_47575);
nand UO_202 (O_202,N_49690,N_46622);
and UO_203 (O_203,N_45821,N_45468);
nand UO_204 (O_204,N_45687,N_45780);
and UO_205 (O_205,N_48660,N_48244);
and UO_206 (O_206,N_47872,N_45620);
nor UO_207 (O_207,N_46565,N_47102);
nor UO_208 (O_208,N_49562,N_45378);
nand UO_209 (O_209,N_45664,N_47696);
or UO_210 (O_210,N_46794,N_48051);
nor UO_211 (O_211,N_49403,N_47216);
and UO_212 (O_212,N_45808,N_49067);
or UO_213 (O_213,N_48990,N_47076);
xor UO_214 (O_214,N_48176,N_45175);
xor UO_215 (O_215,N_45509,N_45491);
xor UO_216 (O_216,N_48350,N_49780);
nor UO_217 (O_217,N_47647,N_49246);
and UO_218 (O_218,N_46511,N_47285);
xor UO_219 (O_219,N_49003,N_47573);
nor UO_220 (O_220,N_47928,N_45294);
nand UO_221 (O_221,N_49008,N_47895);
and UO_222 (O_222,N_48379,N_49678);
or UO_223 (O_223,N_45057,N_46346);
or UO_224 (O_224,N_48450,N_47432);
nor UO_225 (O_225,N_49181,N_45013);
nand UO_226 (O_226,N_45033,N_46294);
and UO_227 (O_227,N_46210,N_49238);
xor UO_228 (O_228,N_49698,N_46370);
nor UO_229 (O_229,N_48841,N_47933);
xor UO_230 (O_230,N_47221,N_46739);
nand UO_231 (O_231,N_47203,N_48209);
xor UO_232 (O_232,N_45954,N_49788);
nand UO_233 (O_233,N_48394,N_48225);
or UO_234 (O_234,N_47701,N_46753);
and UO_235 (O_235,N_45671,N_48659);
nor UO_236 (O_236,N_47580,N_48330);
xnor UO_237 (O_237,N_47547,N_46103);
nor UO_238 (O_238,N_46955,N_45715);
or UO_239 (O_239,N_48054,N_48237);
and UO_240 (O_240,N_48147,N_49325);
nor UO_241 (O_241,N_49647,N_45273);
or UO_242 (O_242,N_47073,N_48622);
nand UO_243 (O_243,N_47871,N_47711);
xor UO_244 (O_244,N_45756,N_45326);
xnor UO_245 (O_245,N_47440,N_48360);
and UO_246 (O_246,N_46626,N_46637);
nand UO_247 (O_247,N_45638,N_49264);
nand UO_248 (O_248,N_49301,N_47658);
or UO_249 (O_249,N_46941,N_45063);
nor UO_250 (O_250,N_49422,N_46957);
nor UO_251 (O_251,N_48378,N_45815);
and UO_252 (O_252,N_49041,N_49545);
and UO_253 (O_253,N_49649,N_45078);
xor UO_254 (O_254,N_49381,N_48969);
nor UO_255 (O_255,N_48482,N_45048);
and UO_256 (O_256,N_46580,N_48236);
xnor UO_257 (O_257,N_48043,N_45001);
or UO_258 (O_258,N_49362,N_45110);
or UO_259 (O_259,N_45095,N_49417);
xnor UO_260 (O_260,N_48965,N_48203);
nand UO_261 (O_261,N_47568,N_48073);
nand UO_262 (O_262,N_48329,N_49787);
and UO_263 (O_263,N_49119,N_49412);
nor UO_264 (O_264,N_49064,N_46821);
and UO_265 (O_265,N_49807,N_46977);
nand UO_266 (O_266,N_45427,N_45365);
nor UO_267 (O_267,N_48310,N_48876);
and UO_268 (O_268,N_46017,N_48910);
and UO_269 (O_269,N_46176,N_47600);
or UO_270 (O_270,N_49988,N_48429);
and UO_271 (O_271,N_48083,N_45891);
or UO_272 (O_272,N_49589,N_45324);
nand UO_273 (O_273,N_49561,N_45141);
xnor UO_274 (O_274,N_45597,N_46316);
xor UO_275 (O_275,N_46853,N_47418);
or UO_276 (O_276,N_49789,N_49378);
nor UO_277 (O_277,N_47081,N_49515);
nand UO_278 (O_278,N_48469,N_48402);
nand UO_279 (O_279,N_47996,N_48044);
nand UO_280 (O_280,N_48315,N_45884);
nand UO_281 (O_281,N_48884,N_49434);
nor UO_282 (O_282,N_45777,N_47307);
and UO_283 (O_283,N_49445,N_47238);
xnor UO_284 (O_284,N_47875,N_45187);
nand UO_285 (O_285,N_47227,N_45785);
and UO_286 (O_286,N_45918,N_45907);
or UO_287 (O_287,N_45905,N_46260);
or UO_288 (O_288,N_47000,N_49976);
or UO_289 (O_289,N_45088,N_48065);
xnor UO_290 (O_290,N_48671,N_46564);
nor UO_291 (O_291,N_49089,N_45641);
xnor UO_292 (O_292,N_48059,N_47298);
nor UO_293 (O_293,N_49909,N_49478);
and UO_294 (O_294,N_45327,N_46686);
and UO_295 (O_295,N_48642,N_47405);
nor UO_296 (O_296,N_46312,N_45003);
xnor UO_297 (O_297,N_48691,N_49653);
or UO_298 (O_298,N_46886,N_47602);
and UO_299 (O_299,N_48839,N_46360);
or UO_300 (O_300,N_49092,N_49893);
or UO_301 (O_301,N_46220,N_47762);
or UO_302 (O_302,N_45113,N_48534);
and UO_303 (O_303,N_47470,N_48780);
nor UO_304 (O_304,N_47534,N_49393);
xnor UO_305 (O_305,N_46273,N_49184);
nand UO_306 (O_306,N_48614,N_49711);
and UO_307 (O_307,N_48631,N_45161);
nor UO_308 (O_308,N_47844,N_49842);
xor UO_309 (O_309,N_47964,N_49673);
and UO_310 (O_310,N_49843,N_45507);
or UO_311 (O_311,N_45178,N_46961);
and UO_312 (O_312,N_49600,N_47553);
or UO_313 (O_313,N_46116,N_48909);
nor UO_314 (O_314,N_48958,N_46568);
or UO_315 (O_315,N_45634,N_49464);
xnor UO_316 (O_316,N_47161,N_47764);
nand UO_317 (O_317,N_48899,N_45275);
and UO_318 (O_318,N_46071,N_46805);
and UO_319 (O_319,N_48222,N_48456);
xnor UO_320 (O_320,N_46378,N_45737);
and UO_321 (O_321,N_45650,N_48420);
and UO_322 (O_322,N_46046,N_49522);
or UO_323 (O_323,N_48738,N_48145);
nor UO_324 (O_324,N_49850,N_47737);
xnor UO_325 (O_325,N_49808,N_45282);
xor UO_326 (O_326,N_49763,N_49002);
xor UO_327 (O_327,N_47100,N_49044);
and UO_328 (O_328,N_47586,N_48777);
nand UO_329 (O_329,N_48160,N_49266);
and UO_330 (O_330,N_46480,N_47422);
or UO_331 (O_331,N_48701,N_47057);
and UO_332 (O_332,N_47788,N_49078);
nor UO_333 (O_333,N_47166,N_45596);
nand UO_334 (O_334,N_46945,N_46583);
xnor UO_335 (O_335,N_49004,N_45822);
xor UO_336 (O_336,N_45591,N_46048);
xor UO_337 (O_337,N_48407,N_47605);
nor UO_338 (O_338,N_47088,N_47025);
xor UO_339 (O_339,N_49071,N_48663);
nand UO_340 (O_340,N_45190,N_48301);
nor UO_341 (O_341,N_49987,N_46693);
xnor UO_342 (O_342,N_48364,N_48034);
or UO_343 (O_343,N_45159,N_47142);
nor UO_344 (O_344,N_46207,N_49700);
or UO_345 (O_345,N_45223,N_47368);
xnor UO_346 (O_346,N_49049,N_46875);
or UO_347 (O_347,N_46226,N_47828);
xor UO_348 (O_348,N_48216,N_48735);
xor UO_349 (O_349,N_46129,N_46254);
nor UO_350 (O_350,N_49658,N_49469);
nand UO_351 (O_351,N_46925,N_48166);
xnor UO_352 (O_352,N_49869,N_48131);
or UO_353 (O_353,N_48498,N_46439);
xor UO_354 (O_354,N_45879,N_49585);
xor UO_355 (O_355,N_47273,N_49720);
nor UO_356 (O_356,N_45967,N_48458);
nor UO_357 (O_357,N_45853,N_48041);
nand UO_358 (O_358,N_49888,N_48666);
or UO_359 (O_359,N_45212,N_46451);
nor UO_360 (O_360,N_48960,N_48328);
and UO_361 (O_361,N_49968,N_48974);
nand UO_362 (O_362,N_45842,N_45899);
or UO_363 (O_363,N_47846,N_48348);
nand UO_364 (O_364,N_47847,N_45557);
nand UO_365 (O_365,N_49892,N_47437);
and UO_366 (O_366,N_47798,N_46247);
xnor UO_367 (O_367,N_45080,N_48292);
xor UO_368 (O_368,N_48645,N_48722);
or UO_369 (O_369,N_45469,N_45656);
and UO_370 (O_370,N_45220,N_49513);
nand UO_371 (O_371,N_48565,N_46001);
xor UO_372 (O_372,N_48204,N_46237);
nand UO_373 (O_373,N_46735,N_47723);
nor UO_374 (O_374,N_47443,N_49689);
nor UO_375 (O_375,N_48655,N_47189);
and UO_376 (O_376,N_48568,N_45173);
nand UO_377 (O_377,N_49985,N_45039);
nand UO_378 (O_378,N_48243,N_45713);
nor UO_379 (O_379,N_49980,N_45116);
or UO_380 (O_380,N_48574,N_48729);
xnor UO_381 (O_381,N_46348,N_46969);
and UO_382 (O_382,N_48070,N_45124);
nor UO_383 (O_383,N_48791,N_46760);
xnor UO_384 (O_384,N_47681,N_49672);
nor UO_385 (O_385,N_48133,N_45508);
xor UO_386 (O_386,N_48956,N_48532);
or UO_387 (O_387,N_49452,N_46643);
xor UO_388 (O_388,N_45006,N_47661);
xor UO_389 (O_389,N_49066,N_48010);
and UO_390 (O_390,N_49302,N_46742);
nand UO_391 (O_391,N_48200,N_49642);
nor UO_392 (O_392,N_47548,N_48792);
xor UO_393 (O_393,N_48020,N_45075);
xnor UO_394 (O_394,N_46566,N_45736);
or UO_395 (O_395,N_47684,N_48470);
xnor UO_396 (O_396,N_47226,N_46530);
xnor UO_397 (O_397,N_47778,N_49159);
xor UO_398 (O_398,N_48019,N_49534);
or UO_399 (O_399,N_45914,N_46023);
nor UO_400 (O_400,N_49918,N_47266);
xnor UO_401 (O_401,N_48079,N_45913);
and UO_402 (O_402,N_45955,N_47358);
nor UO_403 (O_403,N_46282,N_47456);
and UO_404 (O_404,N_47910,N_45200);
xnor UO_405 (O_405,N_48366,N_45606);
nand UO_406 (O_406,N_47452,N_46156);
nand UO_407 (O_407,N_48355,N_46396);
xnor UO_408 (O_408,N_47997,N_47667);
nor UO_409 (O_409,N_46364,N_46648);
and UO_410 (O_410,N_48421,N_45272);
and UO_411 (O_411,N_47730,N_48986);
xnor UO_412 (O_412,N_48557,N_45701);
xnor UO_413 (O_413,N_45387,N_46438);
nor UO_414 (O_414,N_49391,N_49394);
xor UO_415 (O_415,N_46400,N_46732);
xnor UO_416 (O_416,N_49090,N_45845);
or UO_417 (O_417,N_45579,N_49122);
nor UO_418 (O_418,N_46692,N_45721);
or UO_419 (O_419,N_49731,N_47503);
and UO_420 (O_420,N_47228,N_47823);
xnor UO_421 (O_421,N_48577,N_49497);
and UO_422 (O_422,N_48847,N_49915);
nand UO_423 (O_423,N_46833,N_48260);
nor UO_424 (O_424,N_46497,N_46561);
or UO_425 (O_425,N_48480,N_46382);
nand UO_426 (O_426,N_47941,N_47724);
xor UO_427 (O_427,N_46716,N_49740);
xor UO_428 (O_428,N_48881,N_48518);
nand UO_429 (O_429,N_48649,N_45543);
or UO_430 (O_430,N_45465,N_45680);
nand UO_431 (O_431,N_48503,N_48592);
xor UO_432 (O_432,N_48424,N_45347);
and UO_433 (O_433,N_48793,N_45517);
and UO_434 (O_434,N_45270,N_45297);
or UO_435 (O_435,N_48241,N_46717);
and UO_436 (O_436,N_46545,N_49962);
nand UO_437 (O_437,N_48674,N_45236);
nand UO_438 (O_438,N_46971,N_46965);
nor UO_439 (O_439,N_47416,N_45566);
nor UO_440 (O_440,N_48687,N_49244);
xor UO_441 (O_441,N_48252,N_48119);
xnor UO_442 (O_442,N_49155,N_47117);
and UO_443 (O_443,N_47049,N_49162);
or UO_444 (O_444,N_48281,N_48988);
and UO_445 (O_445,N_49819,N_49724);
and UO_446 (O_446,N_48465,N_46173);
or UO_447 (O_447,N_49275,N_46223);
xnor UO_448 (O_448,N_49457,N_49527);
nor UO_449 (O_449,N_45489,N_48374);
and UO_450 (O_450,N_48270,N_48959);
xnor UO_451 (O_451,N_48304,N_49772);
nor UO_452 (O_452,N_45863,N_49292);
and UO_453 (O_453,N_48685,N_46363);
and UO_454 (O_454,N_49755,N_47631);
or UO_455 (O_455,N_45672,N_47319);
xnor UO_456 (O_456,N_46767,N_45038);
and UO_457 (O_457,N_47537,N_49854);
nor UO_458 (O_458,N_48652,N_49738);
or UO_459 (O_459,N_48640,N_47623);
nor UO_460 (O_460,N_48285,N_47763);
and UO_461 (O_461,N_45864,N_47482);
xnor UO_462 (O_462,N_46306,N_46719);
and UO_463 (O_463,N_49193,N_49733);
nand UO_464 (O_464,N_45162,N_45943);
nand UO_465 (O_465,N_47150,N_49967);
xor UO_466 (O_466,N_46027,N_48370);
xnor UO_467 (O_467,N_49009,N_46234);
nand UO_468 (O_468,N_47173,N_45703);
or UO_469 (O_469,N_47079,N_45371);
or UO_470 (O_470,N_47425,N_47207);
or UO_471 (O_471,N_46274,N_45055);
or UO_472 (O_472,N_46314,N_48197);
xor UO_473 (O_473,N_46611,N_48163);
or UO_474 (O_474,N_46161,N_47561);
and UO_475 (O_475,N_45874,N_49488);
or UO_476 (O_476,N_47324,N_48766);
or UO_477 (O_477,N_47218,N_49645);
nand UO_478 (O_478,N_47002,N_47583);
nand UO_479 (O_479,N_48399,N_45682);
and UO_480 (O_480,N_46495,N_48822);
and UO_481 (O_481,N_49657,N_47380);
xor UO_482 (O_482,N_47306,N_49214);
nand UO_483 (O_483,N_47981,N_48999);
and UO_484 (O_484,N_49715,N_46790);
nand UO_485 (O_485,N_49101,N_47199);
xnor UO_486 (O_486,N_46376,N_48836);
nand UO_487 (O_487,N_48962,N_45067);
and UO_488 (O_488,N_48408,N_48306);
nand UO_489 (O_489,N_48906,N_45046);
xor UO_490 (O_490,N_48263,N_45661);
and UO_491 (O_491,N_47957,N_49385);
nand UO_492 (O_492,N_47993,N_48156);
nor UO_493 (O_493,N_47126,N_49520);
and UO_494 (O_494,N_46718,N_49804);
xnor UO_495 (O_495,N_47121,N_48494);
nor UO_496 (O_496,N_46084,N_47733);
xor UO_497 (O_497,N_46204,N_46804);
xnor UO_498 (O_498,N_48063,N_48452);
and UO_499 (O_499,N_48319,N_47654);
and UO_500 (O_500,N_48601,N_47313);
or UO_501 (O_501,N_45164,N_46058);
xnor UO_502 (O_502,N_46005,N_46230);
xor UO_503 (O_503,N_47125,N_49868);
nand UO_504 (O_504,N_46198,N_46228);
nand UO_505 (O_505,N_46100,N_46155);
xnor UO_506 (O_506,N_46861,N_48290);
nor UO_507 (O_507,N_49666,N_47990);
xor UO_508 (O_508,N_46019,N_48217);
or UO_509 (O_509,N_45425,N_46548);
xor UO_510 (O_510,N_47094,N_46981);
or UO_511 (O_511,N_46410,N_48891);
xnor UO_512 (O_512,N_49272,N_46307);
nand UO_513 (O_513,N_47325,N_49276);
or UO_514 (O_514,N_45405,N_48015);
xnor UO_515 (O_515,N_49637,N_47888);
xor UO_516 (O_516,N_45382,N_45819);
and UO_517 (O_517,N_46578,N_46747);
and UO_518 (O_518,N_48396,N_46873);
or UO_519 (O_519,N_47356,N_46892);
xnor UO_520 (O_520,N_45857,N_46588);
and UO_521 (O_521,N_46595,N_47398);
nand UO_522 (O_522,N_46847,N_47795);
xor UO_523 (O_523,N_47275,N_47119);
and UO_524 (O_524,N_46987,N_46776);
nor UO_525 (O_525,N_46609,N_45422);
nor UO_526 (O_526,N_45086,N_46414);
nand UO_527 (O_527,N_46278,N_49632);
and UO_528 (O_528,N_47233,N_49692);
or UO_529 (O_529,N_46264,N_49618);
nor UO_530 (O_530,N_49567,N_48322);
nor UO_531 (O_531,N_48630,N_45343);
nor UO_532 (O_532,N_49170,N_48529);
xnor UO_533 (O_533,N_49794,N_49440);
nor UO_534 (O_534,N_49687,N_46653);
nand UO_535 (O_535,N_49015,N_47262);
and UO_536 (O_536,N_47477,N_47475);
xor UO_537 (O_537,N_49615,N_48393);
nor UO_538 (O_538,N_48702,N_49290);
xor UO_539 (O_539,N_45553,N_49486);
nor UO_540 (O_540,N_47768,N_45000);
or UO_541 (O_541,N_45781,N_48859);
nor UO_542 (O_542,N_48993,N_49269);
and UO_543 (O_543,N_49153,N_48517);
nor UO_544 (O_544,N_49373,N_47391);
nor UO_545 (O_545,N_45330,N_47695);
or UO_546 (O_546,N_45902,N_47390);
and UO_547 (O_547,N_45290,N_46296);
and UO_548 (O_548,N_46536,N_45961);
nand UO_549 (O_549,N_47489,N_48933);
nand UO_550 (O_550,N_46029,N_47773);
nor UO_551 (O_551,N_46593,N_48815);
nor UO_552 (O_552,N_47897,N_47987);
xnor UO_553 (O_553,N_46703,N_49307);
nand UO_554 (O_554,N_48584,N_46138);
nand UO_555 (O_555,N_48124,N_49017);
nor UO_556 (O_556,N_45045,N_48418);
nand UO_557 (O_557,N_49820,N_45938);
and UO_558 (O_558,N_45595,N_49416);
or UO_559 (O_559,N_48426,N_45306);
or UO_560 (O_560,N_47774,N_47946);
or UO_561 (O_561,N_46644,N_47817);
nand UO_562 (O_562,N_48324,N_48202);
nor UO_563 (O_563,N_45612,N_49308);
xnor UO_564 (O_564,N_49601,N_48192);
xor UO_565 (O_565,N_47739,N_49216);
nand UO_566 (O_566,N_47188,N_47407);
nand UO_567 (O_567,N_45227,N_46599);
xnor UO_568 (O_568,N_46834,N_45418);
or UO_569 (O_569,N_45019,N_48255);
or UO_570 (O_570,N_47729,N_45232);
xnor UO_571 (O_571,N_47137,N_48067);
nand UO_572 (O_572,N_46671,N_46783);
nor UO_573 (O_573,N_49526,N_47775);
nor UO_574 (O_574,N_47629,N_45604);
and UO_575 (O_575,N_45937,N_45983);
or UO_576 (O_576,N_45625,N_46368);
nand UO_577 (O_577,N_48914,N_49501);
nor UO_578 (O_578,N_49612,N_46956);
or UO_579 (O_579,N_46369,N_48114);
or UO_580 (O_580,N_45315,N_49144);
and UO_581 (O_581,N_46107,N_49126);
or UO_582 (O_582,N_49555,N_49735);
or UO_583 (O_583,N_48403,N_46429);
or UO_584 (O_584,N_49910,N_47533);
or UO_585 (O_585,N_46701,N_49659);
nor UO_586 (O_586,N_45247,N_45253);
nand UO_587 (O_587,N_49242,N_48570);
xor UO_588 (O_588,N_46256,N_49097);
nor UO_589 (O_589,N_46056,N_47454);
nor UO_590 (O_590,N_49674,N_47584);
or UO_591 (O_591,N_49750,N_46347);
nand UO_592 (O_592,N_47107,N_49198);
xnor UO_593 (O_593,N_47669,N_46788);
and UO_594 (O_594,N_46489,N_48018);
nand UO_595 (O_595,N_48179,N_46238);
nor UO_596 (O_596,N_48994,N_46063);
nor UO_597 (O_597,N_46146,N_48926);
nand UO_598 (O_598,N_49845,N_47138);
and UO_599 (O_599,N_45036,N_48763);
and UO_600 (O_600,N_46183,N_48719);
or UO_601 (O_601,N_47769,N_47793);
and UO_602 (O_602,N_47923,N_46232);
xor UO_603 (O_603,N_49278,N_46784);
and UO_604 (O_604,N_47825,N_48289);
nor UO_605 (O_605,N_45336,N_47083);
and UO_606 (O_606,N_49056,N_45470);
and UO_607 (O_607,N_47849,N_46993);
nor UO_608 (O_608,N_46771,N_47488);
xor UO_609 (O_609,N_45903,N_46197);
or UO_610 (O_610,N_47566,N_47265);
nand UO_611 (O_611,N_48036,N_46554);
or UO_612 (O_612,N_48925,N_47397);
nand UO_613 (O_613,N_48269,N_49083);
and UO_614 (O_614,N_47264,N_47960);
xor UO_615 (O_615,N_48849,N_45589);
nor UO_616 (O_616,N_47136,N_47291);
nand UO_617 (O_617,N_47522,N_48784);
nand UO_618 (O_618,N_45724,N_49778);
nor UO_619 (O_619,N_46055,N_49028);
nor UO_620 (O_620,N_45439,N_46724);
nand UO_621 (O_621,N_46678,N_49800);
and UO_622 (O_622,N_47024,N_46627);
or UO_623 (O_623,N_49407,N_47301);
xnor UO_624 (O_624,N_47009,N_48868);
xor UO_625 (O_625,N_46807,N_49584);
nand UO_626 (O_626,N_49007,N_47592);
or UO_627 (O_627,N_45042,N_49368);
or UO_628 (O_628,N_46562,N_47702);
xnor UO_629 (O_629,N_47512,N_49805);
nand UO_630 (O_630,N_46759,N_48492);
xor UO_631 (O_631,N_48654,N_47697);
or UO_632 (O_632,N_49529,N_49651);
xnor UO_633 (O_633,N_49221,N_45676);
nor UO_634 (O_634,N_48838,N_48483);
nor UO_635 (O_635,N_45839,N_46413);
xnor UO_636 (O_636,N_48776,N_48129);
or UO_637 (O_637,N_48647,N_48916);
xnor UO_638 (O_638,N_45939,N_48698);
nor UO_639 (O_639,N_46498,N_48616);
xnor UO_640 (O_640,N_47208,N_46332);
and UO_641 (O_641,N_46190,N_47980);
xnor UO_642 (O_642,N_49255,N_46280);
xnor UO_643 (O_643,N_49496,N_46258);
nor UO_644 (O_644,N_48146,N_48547);
or UO_645 (O_645,N_48300,N_45073);
and UO_646 (O_646,N_47215,N_48384);
nand UO_647 (O_647,N_47303,N_45923);
or UO_648 (O_648,N_48978,N_45428);
and UO_649 (O_649,N_49996,N_46054);
or UO_650 (O_650,N_46449,N_46640);
nor UO_651 (O_651,N_46009,N_48821);
xnor UO_652 (O_652,N_47782,N_47492);
xor UO_653 (O_653,N_47961,N_47500);
nor UO_654 (O_654,N_49172,N_47797);
nor UO_655 (O_655,N_46756,N_46000);
nand UO_656 (O_656,N_49965,N_48139);
or UO_657 (O_657,N_45283,N_46538);
nor UO_658 (O_658,N_47680,N_49157);
or UO_659 (O_659,N_47555,N_47031);
or UO_660 (O_660,N_45744,N_48487);
xnor UO_661 (O_661,N_48025,N_48955);
nand UO_662 (O_662,N_47506,N_48074);
xor UO_663 (O_663,N_46350,N_47026);
nor UO_664 (O_664,N_48524,N_48130);
xor UO_665 (O_665,N_45688,N_48710);
xor UO_666 (O_666,N_49886,N_48637);
xor UO_667 (O_667,N_49256,N_46344);
nand UO_668 (O_668,N_46911,N_49229);
xor UO_669 (O_669,N_46856,N_47544);
xnor UO_670 (O_670,N_47860,N_49729);
nor UO_671 (O_671,N_47261,N_45257);
nand UO_672 (O_672,N_47059,N_46750);
or UO_673 (O_673,N_47736,N_47281);
xnor UO_674 (O_674,N_49377,N_45202);
nor UO_675 (O_675,N_47921,N_47722);
nand UO_676 (O_676,N_47620,N_49984);
nand UO_677 (O_677,N_49346,N_45117);
nand UO_678 (O_678,N_47651,N_45573);
and UO_679 (O_679,N_49722,N_45645);
or UO_680 (O_680,N_45776,N_49354);
and UO_681 (O_681,N_48164,N_48943);
xnor UO_682 (O_682,N_46086,N_46391);
nand UO_683 (O_683,N_49840,N_47413);
xor UO_684 (O_684,N_48283,N_47182);
nand UO_685 (O_685,N_48811,N_49835);
xor UO_686 (O_686,N_49707,N_49953);
nand UO_687 (O_687,N_49662,N_45865);
or UO_688 (O_688,N_49359,N_45455);
and UO_689 (O_689,N_49115,N_46075);
xnor UO_690 (O_690,N_48461,N_45242);
nand UO_691 (O_691,N_48400,N_48325);
or UO_692 (O_692,N_48153,N_47758);
and UO_693 (O_693,N_45298,N_49776);
and UO_694 (O_694,N_48295,N_49837);
nand UO_695 (O_695,N_46650,N_45922);
and UO_696 (O_696,N_48076,N_45167);
nand UO_697 (O_697,N_47355,N_48143);
and UO_698 (O_698,N_47665,N_45079);
or UO_699 (O_699,N_47294,N_49533);
nand UO_700 (O_700,N_45940,N_47677);
or UO_701 (O_701,N_47591,N_46013);
nand UO_702 (O_702,N_46513,N_49043);
xor UO_703 (O_703,N_45007,N_49327);
or UO_704 (O_704,N_49922,N_46995);
xnor UO_705 (O_705,N_47880,N_47243);
xor UO_706 (O_706,N_45677,N_47246);
and UO_707 (O_707,N_48980,N_49311);
and UO_708 (O_708,N_45755,N_48757);
nand UO_709 (O_709,N_47824,N_45951);
nor UO_710 (O_710,N_46196,N_48109);
xor UO_711 (O_711,N_45476,N_49345);
and UO_712 (O_712,N_46477,N_47429);
or UO_713 (O_713,N_47363,N_48538);
and UO_714 (O_714,N_45997,N_47881);
or UO_715 (O_715,N_47463,N_48029);
xnor UO_716 (O_716,N_46488,N_46523);
nand UO_717 (O_717,N_49160,N_48797);
nand UO_718 (O_718,N_45126,N_49574);
nand UO_719 (O_719,N_48291,N_47241);
and UO_720 (O_720,N_48371,N_48998);
nor UO_721 (O_721,N_46723,N_48650);
nand UO_722 (O_722,N_47942,N_48670);
nand UO_723 (O_723,N_45910,N_49926);
nor UO_724 (O_724,N_48816,N_46366);
nand UO_725 (O_725,N_46077,N_47003);
nor UO_726 (O_726,N_45011,N_46629);
nand UO_727 (O_727,N_48436,N_49027);
nand UO_728 (O_728,N_48030,N_49315);
and UO_729 (O_729,N_47217,N_48369);
xor UO_730 (O_730,N_45363,N_47493);
and UO_731 (O_731,N_45734,N_45165);
or UO_732 (O_732,N_46339,N_45718);
nand UO_733 (O_733,N_46715,N_45312);
xor UO_734 (O_734,N_45195,N_45953);
nor UO_735 (O_735,N_49171,N_49285);
nand UO_736 (O_736,N_46194,N_48923);
nand UO_737 (O_737,N_46646,N_45145);
nand UO_738 (O_738,N_46143,N_48525);
nor UO_739 (O_739,N_47761,N_49247);
or UO_740 (O_740,N_46152,N_48161);
and UO_741 (O_741,N_46793,N_47999);
nor UO_742 (O_742,N_46135,N_49493);
xor UO_743 (O_743,N_45929,N_47685);
nand UO_744 (O_744,N_46577,N_46011);
or UO_745 (O_745,N_46002,N_49990);
and UO_746 (O_746,N_48651,N_45745);
or UO_747 (O_747,N_48915,N_45959);
and UO_748 (O_748,N_47149,N_48240);
nand UO_749 (O_749,N_48112,N_45099);
nor UO_750 (O_750,N_49186,N_47893);
xor UO_751 (O_751,N_47851,N_48001);
xnor UO_752 (O_752,N_46864,N_49459);
nor UO_753 (O_753,N_47939,N_47175);
nor UO_754 (O_754,N_47683,N_48341);
and UO_755 (O_755,N_49928,N_49829);
nand UO_756 (O_756,N_45570,N_48734);
xnor UO_757 (O_757,N_47572,N_46702);
xnor UO_758 (O_758,N_47108,N_49696);
nor UO_759 (O_759,N_46978,N_49449);
nand UO_760 (O_760,N_49194,N_46380);
xor UO_761 (O_761,N_48406,N_48795);
xnor UO_762 (O_762,N_45456,N_45156);
or UO_763 (O_763,N_48772,N_47460);
xnor UO_764 (O_764,N_47706,N_49372);
xnor UO_765 (O_765,N_46460,N_46537);
xnor UO_766 (O_766,N_45152,N_45933);
nand UO_767 (O_767,N_47916,N_49945);
xnor UO_768 (O_768,N_46335,N_49409);
nor UO_769 (O_769,N_45608,N_47237);
or UO_770 (O_770,N_46325,N_47799);
and UO_771 (O_771,N_46673,N_46153);
nor UO_772 (O_772,N_46758,N_46779);
nand UO_773 (O_773,N_45534,N_49259);
or UO_774 (O_774,N_46061,N_47389);
xnor UO_775 (O_775,N_46195,N_45383);
nor UO_776 (O_776,N_49477,N_48765);
nand UO_777 (O_777,N_46634,N_46552);
nand UO_778 (O_778,N_45397,N_47511);
or UO_779 (O_779,N_48796,N_46381);
or UO_780 (O_780,N_49832,N_45501);
or UO_781 (O_781,N_48254,N_48668);
xor UO_782 (O_782,N_48711,N_46652);
and UO_783 (O_783,N_47446,N_49728);
nor UO_784 (O_784,N_46555,N_45322);
xnor UO_785 (O_785,N_47392,N_45191);
xor UO_786 (O_786,N_47036,N_45344);
nor UO_787 (O_787,N_47412,N_46826);
or UO_788 (O_788,N_49337,N_47284);
and UO_789 (O_789,N_48446,N_46125);
nand UO_790 (O_790,N_49430,N_47504);
or UO_791 (O_791,N_45529,N_48113);
xnor UO_792 (O_792,N_47770,N_45120);
nor UO_793 (O_793,N_45966,N_48144);
or UO_794 (O_794,N_46601,N_45380);
nor UO_795 (O_795,N_45069,N_47449);
nor UO_796 (O_796,N_45349,N_49596);
and UO_797 (O_797,N_45148,N_45904);
or UO_798 (O_798,N_47314,N_49458);
or UO_799 (O_799,N_45411,N_45015);
or UO_800 (O_800,N_46430,N_45340);
nand UO_801 (O_801,N_48779,N_48042);
nand UO_802 (O_802,N_45833,N_48810);
nor UO_803 (O_803,N_49636,N_45497);
xor UO_804 (O_804,N_46929,N_45062);
or UO_805 (O_805,N_45044,N_46067);
nand UO_806 (O_806,N_48005,N_45471);
or UO_807 (O_807,N_45252,N_47565);
xnor UO_808 (O_808,N_47712,N_47131);
or UO_809 (O_809,N_45719,N_45345);
nand UO_810 (O_810,N_48072,N_45952);
nand UO_811 (O_811,N_45877,N_48539);
nor UO_812 (O_812,N_49305,N_47757);
nor UO_813 (O_813,N_48188,N_48963);
xnor UO_814 (O_814,N_45854,N_45473);
or UO_815 (O_815,N_49164,N_48338);
or UO_816 (O_816,N_48827,N_48756);
or UO_817 (O_817,N_46014,N_47988);
xnor UO_818 (O_818,N_49352,N_46843);
nor UO_819 (O_819,N_49023,N_47163);
or UO_820 (O_820,N_48992,N_46458);
nor UO_821 (O_821,N_46872,N_47856);
xor UO_822 (O_822,N_48693,N_46585);
nand UO_823 (O_823,N_47842,N_46808);
and UO_824 (O_824,N_47603,N_47760);
nor UO_825 (O_825,N_49312,N_48856);
or UO_826 (O_826,N_45653,N_47643);
and UO_827 (O_827,N_45683,N_46124);
nor UO_828 (O_828,N_49793,N_49491);
or UO_829 (O_829,N_47191,N_45129);
and UO_830 (O_830,N_49330,N_47160);
and UO_831 (O_831,N_45817,N_45115);
xor UO_832 (O_832,N_48238,N_46288);
nand UO_833 (O_833,N_46612,N_49969);
xnor UO_834 (O_834,N_47630,N_46474);
or UO_835 (O_835,N_49350,N_48506);
nand UO_836 (O_836,N_49761,N_48721);
or UO_837 (O_837,N_48860,N_46824);
and UO_838 (O_838,N_46479,N_48716);
nand UO_839 (O_839,N_47562,N_49894);
nand UO_840 (O_840,N_47195,N_48682);
nor UO_841 (O_841,N_46231,N_48412);
nor UO_842 (O_842,N_49355,N_46191);
xor UO_843 (O_843,N_45460,N_45971);
and UO_844 (O_844,N_45847,N_48249);
and UO_845 (O_845,N_49603,N_49625);
xor UO_846 (O_846,N_49060,N_47917);
nor UO_847 (O_847,N_45201,N_49798);
nor UO_848 (O_848,N_46281,N_48609);
xor UO_849 (O_849,N_49553,N_48226);
nor UO_850 (O_850,N_48902,N_47316);
xor UO_851 (O_851,N_49135,N_47787);
and UO_852 (O_852,N_49531,N_45091);
and UO_853 (O_853,N_48932,N_47184);
nor UO_854 (O_854,N_47103,N_47353);
xor UO_855 (O_855,N_49147,N_47717);
nor UO_856 (O_856,N_49865,N_45944);
and UO_857 (O_857,N_47514,N_46751);
nor UO_858 (O_858,N_45419,N_45875);
nor UO_859 (O_859,N_46177,N_46175);
nor UO_860 (O_860,N_48945,N_47614);
xor UO_861 (O_861,N_46827,N_45858);
nand UO_862 (O_862,N_48367,N_47892);
and UO_863 (O_863,N_48345,N_46434);
or UO_864 (O_864,N_46455,N_48442);
nor UO_865 (O_865,N_46371,N_46496);
nand UO_866 (O_866,N_45783,N_48024);
nor UO_867 (O_867,N_48286,N_49877);
or UO_868 (O_868,N_49415,N_46229);
or UO_869 (O_869,N_45458,N_47965);
nand UO_870 (O_870,N_48233,N_46462);
xnor UO_871 (O_871,N_45401,N_49621);
and UO_872 (O_872,N_47975,N_45293);
and UO_873 (O_873,N_48607,N_49085);
xor UO_874 (O_874,N_49287,N_45368);
and UO_875 (O_875,N_46922,N_49528);
xor UO_876 (O_876,N_45614,N_49435);
xnor UO_877 (O_877,N_45390,N_49823);
nor UO_878 (O_878,N_45441,N_45510);
or UO_879 (O_879,N_45034,N_48490);
nand UO_880 (O_880,N_46814,N_49298);
xnor UO_881 (O_881,N_46579,N_48275);
xnor UO_882 (O_882,N_48433,N_45803);
or UO_883 (O_883,N_49903,N_46879);
or UO_884 (O_884,N_45020,N_49363);
or UO_885 (O_885,N_49190,N_45757);
nand UO_886 (O_886,N_46006,N_46491);
or UO_887 (O_887,N_47850,N_47900);
nand UO_888 (O_888,N_47571,N_47976);
and UO_889 (O_889,N_49187,N_49441);
or UO_890 (O_890,N_48997,N_47364);
xor UO_891 (O_891,N_45818,N_49114);
or UO_892 (O_892,N_46699,N_47043);
nor UO_893 (O_893,N_48011,N_49758);
and UO_894 (O_894,N_48386,N_46535);
nand UO_895 (O_895,N_46951,N_47633);
and UO_896 (O_896,N_46044,N_47542);
or UO_897 (O_897,N_48519,N_45748);
xor UO_898 (O_898,N_48463,N_45176);
xnor UO_899 (O_899,N_47903,N_48069);
nand UO_900 (O_900,N_46698,N_49716);
nor UO_901 (O_901,N_45978,N_45233);
xor UO_902 (O_902,N_48760,N_49146);
nor UO_903 (O_903,N_48390,N_46035);
nor UO_904 (O_904,N_47344,N_47524);
nor UO_905 (O_905,N_49383,N_46934);
xor UO_906 (O_906,N_48930,N_48852);
or UO_907 (O_907,N_49577,N_49125);
and UO_908 (O_908,N_45963,N_45160);
and UO_909 (O_909,N_45739,N_47197);
xor UO_910 (O_910,N_46736,N_46233);
nor UO_911 (O_911,N_49576,N_45706);
and UO_912 (O_912,N_45663,N_48207);
or UO_913 (O_913,N_48459,N_47185);
and UO_914 (O_914,N_45488,N_47139);
nand UO_915 (O_915,N_48605,N_46915);
or UO_916 (O_916,N_49471,N_46299);
nand UO_917 (O_917,N_47519,N_46694);
nor UO_918 (O_918,N_47257,N_47343);
nand UO_919 (O_919,N_46976,N_48410);
xor UO_920 (O_920,N_49997,N_49024);
or UO_921 (O_921,N_47192,N_47190);
xnor UO_922 (O_922,N_45799,N_46763);
xnor UO_923 (O_923,N_45163,N_48851);
or UO_924 (O_924,N_48388,N_46057);
and UO_925 (O_925,N_45546,N_49708);
nand UO_926 (O_926,N_46908,N_49180);
or UO_927 (O_927,N_48871,N_47334);
xor UO_928 (O_928,N_47061,N_49547);
and UO_929 (O_929,N_46453,N_49014);
or UO_930 (O_930,N_47288,N_48343);
nor UO_931 (O_931,N_48351,N_46213);
or UO_932 (O_932,N_48747,N_49906);
and UO_933 (O_933,N_49336,N_47455);
nand UO_934 (O_934,N_47436,N_47019);
xnor UO_935 (O_935,N_46292,N_49237);
nand UO_936 (O_936,N_48086,N_46898);
nand UO_937 (O_937,N_48718,N_49150);
nand UO_938 (O_938,N_45729,N_45975);
nor UO_939 (O_939,N_46432,N_46040);
nor UO_940 (O_940,N_48175,N_45452);
nor UO_941 (O_941,N_48387,N_47668);
nor UO_942 (O_942,N_49905,N_48023);
nand UO_943 (O_943,N_46666,N_48976);
xor UO_944 (O_944,N_46249,N_49638);
xor UO_945 (O_945,N_45498,N_47699);
or UO_946 (O_946,N_46245,N_48855);
xor UO_947 (O_947,N_46745,N_47231);
or UO_948 (O_948,N_45065,N_47649);
xor UO_949 (O_949,N_48221,N_46505);
or UO_950 (O_950,N_47859,N_48773);
xor UO_951 (O_951,N_48578,N_47168);
nand UO_952 (O_952,N_49851,N_47030);
and UO_953 (O_953,N_46221,N_45094);
or UO_954 (O_954,N_47206,N_48448);
nand UO_955 (O_955,N_45081,N_45886);
or UO_956 (O_956,N_47767,N_46526);
nor UO_957 (O_957,N_46709,N_45563);
nand UO_958 (O_958,N_47790,N_49370);
nand UO_959 (O_959,N_49016,N_45530);
and UO_960 (O_960,N_49117,N_46028);
and UO_961 (O_961,N_46345,N_48526);
xnor UO_962 (O_962,N_46743,N_47116);
or UO_963 (O_963,N_49631,N_49310);
xor UO_964 (O_964,N_48581,N_48786);
nand UO_965 (O_965,N_47372,N_46822);
or UO_966 (O_966,N_48879,N_45292);
nor UO_967 (O_967,N_49294,N_49862);
xor UO_968 (O_968,N_48353,N_48045);
or UO_969 (O_969,N_48515,N_46620);
nor UO_970 (O_970,N_47590,N_46734);
or UO_971 (O_971,N_47230,N_49946);
or UO_972 (O_972,N_47354,N_49670);
nand UO_973 (O_973,N_49300,N_48383);
nand UO_974 (O_974,N_47918,N_46365);
or UO_975 (O_975,N_49810,N_47595);
xnor UO_976 (O_976,N_49989,N_48755);
xor UO_977 (O_977,N_47687,N_48091);
nor UO_978 (O_978,N_48727,N_49899);
nand UO_979 (O_979,N_49767,N_45690);
and UO_980 (O_980,N_45339,N_45685);
or UO_981 (O_981,N_47827,N_46517);
xor UO_982 (O_982,N_46604,N_49644);
and UO_983 (O_983,N_46433,N_47223);
or UO_984 (O_984,N_46603,N_45026);
xnor UO_985 (O_985,N_45704,N_49834);
or UO_986 (O_986,N_46270,N_49156);
and UO_987 (O_987,N_46506,N_45364);
xnor UO_988 (O_988,N_45577,N_49699);
nand UO_989 (O_989,N_45582,N_45569);
nor UO_990 (O_990,N_49005,N_46101);
xnor UO_991 (O_991,N_48404,N_47090);
nand UO_992 (O_992,N_48451,N_48303);
and UO_993 (O_993,N_45871,N_47037);
nand UO_994 (O_994,N_49695,N_47920);
nand UO_995 (O_995,N_46172,N_47092);
and UO_996 (O_996,N_48274,N_46803);
nor UO_997 (O_997,N_45505,N_49944);
or UO_998 (O_998,N_46748,N_45464);
xnor UO_999 (O_999,N_47224,N_47001);
xnor UO_1000 (O_1000,N_47210,N_48297);
nand UO_1001 (O_1001,N_48554,N_47145);
and UO_1002 (O_1002,N_47251,N_49624);
xnor UO_1003 (O_1003,N_46286,N_45433);
and UO_1004 (O_1004,N_45481,N_47202);
or UO_1005 (O_1005,N_47008,N_45357);
or UO_1006 (O_1006,N_46683,N_47010);
and UO_1007 (O_1007,N_46837,N_48000);
or UO_1008 (O_1008,N_46927,N_48522);
and UO_1009 (O_1009,N_47815,N_47468);
xor UO_1010 (O_1010,N_49149,N_45908);
or UO_1011 (O_1011,N_45192,N_46882);
nor UO_1012 (O_1012,N_45313,N_49251);
nand UO_1013 (O_1013,N_48089,N_46354);
or UO_1014 (O_1014,N_48929,N_45155);
nand UO_1015 (O_1015,N_47588,N_48726);
nand UO_1016 (O_1016,N_47984,N_49034);
or UO_1017 (O_1017,N_49329,N_48478);
nand UO_1018 (O_1018,N_49366,N_47383);
nand UO_1019 (O_1019,N_46854,N_46891);
nand UO_1020 (O_1020,N_45962,N_45490);
nor UO_1021 (O_1021,N_47732,N_47531);
and UO_1022 (O_1022,N_48280,N_45056);
xnor UO_1023 (O_1023,N_46494,N_46171);
xor UO_1024 (O_1024,N_49942,N_48340);
nand UO_1025 (O_1025,N_48759,N_47540);
or UO_1026 (O_1026,N_48804,N_47027);
nand UO_1027 (O_1027,N_46722,N_45615);
nor UO_1028 (O_1028,N_45691,N_47513);
and UO_1029 (O_1029,N_46073,N_47930);
or UO_1030 (O_1030,N_46398,N_46182);
and UO_1031 (O_1031,N_46870,N_45267);
or UO_1032 (O_1032,N_47528,N_48528);
nor UO_1033 (O_1033,N_47924,N_45172);
or UO_1034 (O_1034,N_49054,N_49855);
nand UO_1035 (O_1035,N_45670,N_47433);
nand UO_1036 (O_1036,N_48356,N_47021);
or UO_1037 (O_1037,N_46880,N_45068);
nand UO_1038 (O_1038,N_47559,N_47086);
nand UO_1039 (O_1039,N_47338,N_48560);
and UO_1040 (O_1040,N_49920,N_48127);
nor UO_1041 (O_1041,N_48700,N_48703);
xnor UO_1042 (O_1042,N_46942,N_47746);
and UO_1043 (O_1043,N_49917,N_49744);
xor UO_1044 (O_1044,N_46900,N_48061);
or UO_1045 (O_1045,N_49467,N_46200);
nor UO_1046 (O_1046,N_45514,N_45502);
xor UO_1047 (O_1047,N_49331,N_45710);
nor UO_1048 (O_1048,N_49871,N_48081);
or UO_1049 (O_1049,N_48583,N_47624);
and UO_1050 (O_1050,N_47835,N_45702);
xor UO_1051 (O_1051,N_45868,N_48264);
or UO_1052 (O_1052,N_47992,N_46313);
or UO_1053 (O_1053,N_49367,N_46126);
or UO_1054 (O_1054,N_47577,N_45965);
and UO_1055 (O_1055,N_46361,N_48165);
xor UO_1056 (O_1056,N_49199,N_48125);
and UO_1057 (O_1057,N_47300,N_46770);
xor UO_1058 (O_1058,N_47606,N_45587);
and UO_1059 (O_1059,N_48947,N_46324);
nor UO_1060 (O_1060,N_48633,N_48500);
nand UO_1061 (O_1061,N_49650,N_49232);
nand UO_1062 (O_1062,N_49519,N_45179);
or UO_1063 (O_1063,N_46192,N_48247);
nand UO_1064 (O_1064,N_46285,N_46656);
and UO_1065 (O_1065,N_47317,N_49723);
nor UO_1066 (O_1066,N_45666,N_48033);
nor UO_1067 (O_1067,N_49200,N_46792);
or UO_1068 (O_1068,N_46051,N_47517);
xor UO_1069 (O_1069,N_48256,N_49136);
xnor UO_1070 (O_1070,N_47385,N_48883);
nor UO_1071 (O_1071,N_46250,N_48309);
or UO_1072 (O_1072,N_46528,N_45264);
or UO_1073 (O_1073,N_47686,N_46099);
nor UO_1074 (O_1074,N_45600,N_47063);
or UO_1075 (O_1075,N_45434,N_49038);
nor UO_1076 (O_1076,N_49314,N_46276);
or UO_1077 (O_1077,N_46320,N_45208);
xor UO_1078 (O_1078,N_48055,N_47937);
nand UO_1079 (O_1079,N_46343,N_45873);
xnor UO_1080 (O_1080,N_48382,N_46636);
nor UO_1081 (O_1081,N_47130,N_46820);
nand UO_1082 (O_1082,N_49088,N_47913);
xnor UO_1083 (O_1083,N_48035,N_47752);
nor UO_1084 (O_1084,N_48928,N_46211);
or UO_1085 (O_1085,N_46336,N_46287);
nor UO_1086 (O_1086,N_49552,N_47347);
and UO_1087 (O_1087,N_45585,N_45426);
or UO_1088 (O_1088,N_48939,N_47956);
nor UO_1089 (O_1089,N_48422,N_47023);
xnor UO_1090 (O_1090,N_49774,N_46812);
or UO_1091 (O_1091,N_45399,N_49986);
nor UO_1092 (O_1092,N_49098,N_48215);
nor UO_1093 (O_1093,N_45482,N_45635);
nand UO_1094 (O_1094,N_49222,N_48060);
nor UO_1095 (O_1095,N_46654,N_47989);
and UO_1096 (O_1096,N_49379,N_47628);
xnor UO_1097 (O_1097,N_45435,N_45028);
xnor UO_1098 (O_1098,N_48116,N_47322);
nor UO_1099 (O_1099,N_47099,N_46881);
or UO_1100 (O_1100,N_47194,N_49390);
and UO_1101 (O_1101,N_45424,N_47359);
xor UO_1102 (O_1102,N_45972,N_46147);
xnor UO_1103 (O_1103,N_46300,N_47157);
nand UO_1104 (O_1104,N_46920,N_47952);
and UO_1105 (O_1105,N_45747,N_47541);
and UO_1106 (O_1106,N_45052,N_46050);
or UO_1107 (O_1107,N_49921,N_45342);
xor UO_1108 (O_1108,N_48477,N_45520);
nand UO_1109 (O_1109,N_45605,N_46714);
nand UO_1110 (O_1110,N_46082,N_49675);
and UO_1111 (O_1111,N_48549,N_46970);
nand UO_1112 (O_1112,N_45732,N_47931);
or UO_1113 (O_1113,N_48894,N_48331);
or UO_1114 (O_1114,N_45695,N_46179);
xnor UO_1115 (O_1115,N_48569,N_46775);
and UO_1116 (O_1116,N_46131,N_47959);
nand UO_1117 (O_1117,N_47340,N_49406);
and UO_1118 (O_1118,N_47458,N_49213);
xnor UO_1119 (O_1119,N_49523,N_47062);
xor UO_1120 (O_1120,N_47180,N_45012);
or UO_1121 (O_1121,N_49769,N_47979);
or UO_1122 (O_1122,N_45072,N_49825);
xor UO_1123 (O_1123,N_47304,N_49112);
nand UO_1124 (O_1124,N_46731,N_46120);
or UO_1125 (O_1125,N_48541,N_46144);
and UO_1126 (O_1126,N_49263,N_46142);
and UO_1127 (O_1127,N_48191,N_49323);
nor UO_1128 (O_1128,N_47474,N_47756);
xnor UO_1129 (O_1129,N_45956,N_45437);
nand UO_1130 (O_1130,N_47330,N_47841);
nor UO_1131 (O_1131,N_45066,N_49912);
and UO_1132 (O_1132,N_47902,N_48571);
or UO_1133 (O_1133,N_46935,N_48423);
nand UO_1134 (O_1134,N_45725,N_45412);
xor UO_1135 (O_1135,N_47060,N_47678);
or UO_1136 (O_1136,N_45931,N_47970);
and UO_1137 (O_1137,N_47616,N_45193);
nand UO_1138 (O_1138,N_47201,N_48527);
xor UO_1139 (O_1139,N_48613,N_49914);
nand UO_1140 (O_1140,N_46574,N_46532);
or UO_1141 (O_1141,N_49872,N_45386);
nand UO_1142 (O_1142,N_49291,N_49499);
nor UO_1143 (O_1143,N_47070,N_46167);
or UO_1144 (O_1144,N_45583,N_45385);
xnor UO_1145 (O_1145,N_49489,N_47594);
nand UO_1146 (O_1146,N_49925,N_48110);
nand UO_1147 (O_1147,N_46904,N_48606);
nor UO_1148 (O_1148,N_46777,N_45070);
nand UO_1149 (O_1149,N_49654,N_49011);
nor UO_1150 (O_1150,N_49504,N_48278);
xor UO_1151 (O_1151,N_47626,N_48880);
and UO_1152 (O_1152,N_48924,N_49289);
nor UO_1153 (O_1153,N_49993,N_47012);
nor UO_1154 (O_1154,N_49437,N_45051);
or UO_1155 (O_1155,N_46889,N_47387);
or UO_1156 (O_1156,N_45493,N_47601);
or UO_1157 (O_1157,N_47447,N_45667);
and UO_1158 (O_1158,N_49261,N_45218);
xnor UO_1159 (O_1159,N_49208,N_49560);
nor UO_1160 (O_1160,N_45370,N_45607);
nor UO_1161 (O_1161,N_45658,N_46043);
and UO_1162 (O_1162,N_48604,N_47708);
nand UO_1163 (O_1163,N_48497,N_49901);
xor UO_1164 (O_1164,N_45133,N_49382);
and UO_1165 (O_1165,N_46277,N_47113);
xor UO_1166 (O_1166,N_47636,N_49411);
nand UO_1167 (O_1167,N_49818,N_46261);
or UO_1168 (O_1168,N_45981,N_48907);
nor UO_1169 (O_1169,N_48775,N_46876);
xor UO_1170 (O_1170,N_48159,N_49324);
nand UO_1171 (O_1171,N_49433,N_47444);
and UO_1172 (O_1172,N_45613,N_46259);
and UO_1173 (O_1173,N_49815,N_45136);
nor UO_1174 (O_1174,N_47170,N_46586);
xnor UO_1175 (O_1175,N_45611,N_49070);
or UO_1176 (O_1176,N_48212,N_49705);
or UO_1177 (O_1177,N_46862,N_46857);
or UO_1178 (O_1178,N_47527,N_49475);
and UO_1179 (O_1179,N_48675,N_49484);
nand UO_1180 (O_1180,N_46109,N_46575);
nand UO_1181 (O_1181,N_49371,N_48293);
or UO_1182 (O_1182,N_46189,N_49949);
nand UO_1183 (O_1183,N_49958,N_46386);
xor UO_1184 (O_1184,N_46907,N_47406);
and UO_1185 (O_1185,N_49543,N_46980);
nand UO_1186 (O_1186,N_45561,N_48720);
nand UO_1187 (O_1187,N_46800,N_45277);
and UO_1188 (O_1188,N_49514,N_45675);
or UO_1189 (O_1189,N_48694,N_48177);
or UO_1190 (O_1190,N_49575,N_45554);
and UO_1191 (O_1191,N_48320,N_48661);
xor UO_1192 (O_1192,N_47803,N_48449);
or UO_1193 (O_1193,N_48801,N_45532);
nand UO_1194 (O_1194,N_47423,N_46209);
xor UO_1195 (O_1195,N_45897,N_49356);
nor UO_1196 (O_1196,N_49341,N_48732);
nand UO_1197 (O_1197,N_49535,N_45361);
and UO_1198 (O_1198,N_47484,N_49762);
xor UO_1199 (O_1199,N_46590,N_45632);
nor UO_1200 (O_1200,N_45697,N_45767);
nand UO_1201 (O_1201,N_47248,N_46740);
or UO_1202 (O_1202,N_49630,N_49030);
nand UO_1203 (O_1203,N_47925,N_46606);
nand UO_1204 (O_1204,N_48047,N_46105);
nand UO_1205 (O_1205,N_48111,N_46141);
nor UO_1206 (O_1206,N_45533,N_49900);
or UO_1207 (O_1207,N_47948,N_49402);
nor UO_1208 (O_1208,N_47857,N_46738);
xnor UO_1209 (O_1209,N_46484,N_46937);
or UO_1210 (O_1210,N_47829,N_45030);
or UO_1211 (O_1211,N_47260,N_48803);
xor UO_1212 (O_1212,N_49580,N_47075);
or UO_1213 (O_1213,N_47378,N_47465);
xnor UO_1214 (O_1214,N_49725,N_47496);
nor UO_1215 (O_1215,N_45430,N_46996);
or UO_1216 (O_1216,N_49262,N_49252);
xnor UO_1217 (O_1217,N_47315,N_45800);
nand UO_1218 (O_1218,N_47843,N_49844);
and UO_1219 (O_1219,N_49579,N_47710);
nor UO_1220 (O_1220,N_46607,N_45643);
or UO_1221 (O_1221,N_47362,N_47557);
or UO_1222 (O_1222,N_46500,N_47894);
xor UO_1223 (O_1223,N_46720,N_47840);
nand UO_1224 (O_1224,N_46483,N_49450);
xnor UO_1225 (O_1225,N_48603,N_48158);
nand UO_1226 (O_1226,N_48180,N_45211);
or UO_1227 (O_1227,N_48673,N_46215);
nand UO_1228 (O_1228,N_46944,N_48862);
nand UO_1229 (O_1229,N_47478,N_48809);
xnor UO_1230 (O_1230,N_48745,N_46591);
nand UO_1231 (O_1231,N_45572,N_48866);
or UO_1232 (O_1232,N_48696,N_45602);
and UO_1233 (O_1233,N_46639,N_46110);
or UO_1234 (O_1234,N_46655,N_46407);
nor UO_1235 (O_1235,N_49726,N_46016);
nor UO_1236 (O_1236,N_48495,N_48206);
and UO_1237 (O_1237,N_49245,N_47891);
or UO_1238 (O_1238,N_46542,N_47109);
and UO_1239 (O_1239,N_47838,N_45154);
nand UO_1240 (O_1240,N_45479,N_45182);
and UO_1241 (O_1241,N_45883,N_49864);
or UO_1242 (O_1242,N_46540,N_46428);
nand UO_1243 (O_1243,N_47878,N_47154);
and UO_1244 (O_1244,N_46225,N_45125);
nor UO_1245 (O_1245,N_47639,N_46351);
nand UO_1246 (O_1246,N_46367,N_48155);
nand UO_1247 (O_1247,N_47564,N_46810);
nand UO_1248 (O_1248,N_49059,N_45423);
and UO_1249 (O_1249,N_46539,N_45278);
nor UO_1250 (O_1250,N_45093,N_45317);
and UO_1251 (O_1251,N_48704,N_47219);
xnor UO_1252 (O_1252,N_46974,N_49792);
nand UO_1253 (O_1253,N_45140,N_47525);
xor UO_1254 (O_1254,N_47804,N_45731);
xor UO_1255 (O_1255,N_49077,N_45137);
nand UO_1256 (O_1256,N_48987,N_49145);
xnor UO_1257 (O_1257,N_45031,N_47420);
and UO_1258 (O_1258,N_49813,N_47906);
xnor UO_1259 (O_1259,N_46151,N_48690);
xor UO_1260 (O_1260,N_49248,N_48643);
or UO_1261 (O_1261,N_48794,N_46918);
nand UO_1262 (O_1262,N_49712,N_48126);
nand UO_1263 (O_1263,N_47742,N_48752);
nand UO_1264 (O_1264,N_46512,N_45025);
nand UO_1265 (O_1265,N_47384,N_47236);
xnor UO_1266 (O_1266,N_48966,N_48430);
nor UO_1267 (O_1267,N_47973,N_49544);
and UO_1268 (O_1268,N_47805,N_49559);
or UO_1269 (O_1269,N_45448,N_47751);
nand UO_1270 (O_1270,N_46140,N_49451);
nor UO_1271 (O_1271,N_47134,N_46321);
nor UO_1272 (O_1272,N_49438,N_45813);
nand UO_1273 (O_1273,N_47295,N_45478);
or UO_1274 (O_1274,N_47032,N_45796);
or UO_1275 (O_1275,N_49749,N_49640);
and UO_1276 (O_1276,N_45122,N_48590);
nor UO_1277 (O_1277,N_48826,N_48983);
nand UO_1278 (O_1278,N_48951,N_48850);
or UO_1279 (O_1279,N_47832,N_45406);
nand UO_1280 (O_1280,N_45228,N_46265);
nor UO_1281 (O_1281,N_45369,N_47510);
nor UO_1282 (O_1282,N_47267,N_47735);
nand UO_1283 (O_1283,N_45229,N_49281);
nand UO_1284 (O_1284,N_47848,N_49322);
nor UO_1285 (O_1285,N_48199,N_45064);
nand UO_1286 (O_1286,N_47491,N_48105);
and UO_1287 (O_1287,N_47863,N_46478);
or UO_1288 (O_1288,N_46533,N_47604);
nand UO_1289 (O_1289,N_48877,N_46613);
or UO_1290 (O_1290,N_46761,N_49058);
nor UO_1291 (O_1291,N_49413,N_45335);
xnor UO_1292 (O_1292,N_45977,N_45758);
nand UO_1293 (O_1293,N_47644,N_45665);
nand UO_1294 (O_1294,N_48644,N_49790);
nand UO_1295 (O_1295,N_47945,N_47321);
or UO_1296 (O_1296,N_47587,N_49206);
or UO_1297 (O_1297,N_47448,N_49667);
xor UO_1298 (O_1298,N_45834,N_47054);
or UO_1299 (O_1299,N_45249,N_46136);
xnor UO_1300 (O_1300,N_45023,N_47963);
and UO_1301 (O_1301,N_45555,N_46416);
or UO_1302 (O_1302,N_48031,N_46796);
and UO_1303 (O_1303,N_46660,N_48624);
xor UO_1304 (O_1304,N_45262,N_48996);
nand UO_1305 (O_1305,N_45708,N_46330);
nor UO_1306 (O_1306,N_48540,N_47582);
and UO_1307 (O_1307,N_49414,N_45869);
and UO_1308 (O_1308,N_46353,N_46989);
nor UO_1309 (O_1309,N_47084,N_49747);
nor UO_1310 (O_1310,N_47904,N_45810);
xnor UO_1311 (O_1311,N_46623,N_45005);
nor UO_1312 (O_1312,N_48381,N_46906);
and UO_1313 (O_1313,N_48641,N_48743);
or UO_1314 (O_1314,N_48798,N_48302);
xnor UO_1315 (O_1315,N_47439,N_46871);
or UO_1316 (O_1316,N_47310,N_49686);
and UO_1317 (O_1317,N_46630,N_45318);
nand UO_1318 (O_1318,N_45254,N_47727);
xnor UO_1319 (O_1319,N_48754,N_49087);
and UO_1320 (O_1320,N_47884,N_48977);
xor UO_1321 (O_1321,N_48676,N_45827);
and UO_1322 (O_1322,N_49943,N_45022);
nand UO_1323 (O_1323,N_49453,N_48228);
nor UO_1324 (O_1324,N_48505,N_48626);
nand UO_1325 (O_1325,N_45089,N_45686);
and UO_1326 (O_1326,N_48401,N_48502);
and UO_1327 (O_1327,N_47494,N_45571);
or UO_1328 (O_1328,N_46089,N_47485);
or UO_1329 (O_1329,N_48968,N_46493);
xnor UO_1330 (O_1330,N_47045,N_45027);
xor UO_1331 (O_1331,N_49432,N_48979);
xor UO_1332 (O_1332,N_48699,N_47662);
xnor UO_1333 (O_1333,N_49094,N_48117);
xor UO_1334 (O_1334,N_46085,N_45299);
or UO_1335 (O_1335,N_49271,N_46372);
nand UO_1336 (O_1336,N_46773,N_46520);
xnor UO_1337 (O_1337,N_49466,N_49604);
nand UO_1338 (O_1338,N_48799,N_48817);
or UO_1339 (O_1339,N_45205,N_48075);
xnor UO_1340 (O_1340,N_47411,N_46902);
nor UO_1341 (O_1341,N_49568,N_48501);
or UO_1342 (O_1342,N_49052,N_49032);
nor UO_1343 (O_1343,N_49999,N_49188);
nand UO_1344 (O_1344,N_48919,N_48488);
xnor UO_1345 (O_1345,N_45074,N_45673);
and UO_1346 (O_1346,N_45147,N_46267);
xnor UO_1347 (O_1347,N_46600,N_49019);
or UO_1348 (O_1348,N_48874,N_48741);
and UO_1349 (O_1349,N_47165,N_47609);
nor UO_1350 (O_1350,N_46170,N_47994);
nand UO_1351 (O_1351,N_49831,N_46079);
xnor UO_1352 (O_1352,N_45353,N_45894);
and UO_1353 (O_1353,N_48689,N_49029);
or UO_1354 (O_1354,N_45824,N_46518);
or UO_1355 (O_1355,N_49911,N_47250);
xnor UO_1356 (O_1356,N_48313,N_49399);
nor UO_1357 (O_1357,N_47403,N_47983);
nor UO_1358 (O_1358,N_46465,N_45949);
or UO_1359 (O_1359,N_48995,N_49973);
and UO_1360 (O_1360,N_47158,N_45018);
nor UO_1361 (O_1361,N_45723,N_46930);
or UO_1362 (O_1362,N_47927,N_49791);
or UO_1363 (O_1363,N_45241,N_46178);
or UO_1364 (O_1364,N_49127,N_49339);
and UO_1365 (O_1365,N_47789,N_48235);
or UO_1366 (O_1366,N_49652,N_45782);
or UO_1367 (O_1367,N_46729,N_48858);
nand UO_1368 (O_1368,N_45712,N_49971);
nor UO_1369 (O_1369,N_45684,N_46469);
nand UO_1370 (O_1370,N_47652,N_47714);
nand UO_1371 (O_1371,N_47483,N_47435);
and UO_1372 (O_1372,N_48981,N_46150);
nand UO_1373 (O_1373,N_49856,N_48597);
nand UO_1374 (O_1374,N_46373,N_45565);
and UO_1375 (O_1375,N_46319,N_46417);
or UO_1376 (O_1376,N_47292,N_45054);
nand UO_1377 (O_1377,N_46305,N_45485);
and UO_1378 (O_1378,N_49786,N_49759);
or UO_1379 (O_1379,N_47016,N_46065);
nor UO_1380 (O_1380,N_45784,N_49785);
xor UO_1381 (O_1381,N_45631,N_49254);
nor UO_1382 (O_1382,N_48705,N_49606);
and UO_1383 (O_1383,N_45214,N_48665);
nor UO_1384 (O_1384,N_45870,N_45444);
nand UO_1385 (O_1385,N_47256,N_46581);
xnor UO_1386 (O_1386,N_49128,N_47178);
xor UO_1387 (O_1387,N_46874,N_45945);
and UO_1388 (O_1388,N_45654,N_48190);
nand UO_1389 (O_1389,N_45942,N_47038);
nor UO_1390 (O_1390,N_46635,N_49929);
xnor UO_1391 (O_1391,N_46060,N_45999);
or UO_1392 (O_1392,N_48428,N_49288);
nand UO_1393 (O_1393,N_48068,N_49454);
xor UO_1394 (O_1394,N_49130,N_49349);
and UO_1395 (O_1395,N_45925,N_48395);
or UO_1396 (O_1396,N_49418,N_46700);
nor UO_1397 (O_1397,N_45766,N_49884);
and UO_1398 (O_1398,N_46384,N_45123);
or UO_1399 (O_1399,N_46616,N_47277);
and UO_1400 (O_1400,N_47883,N_46037);
xnor UO_1401 (O_1401,N_48612,N_47242);
xor UO_1402 (O_1402,N_45403,N_46910);
nor UO_1403 (O_1403,N_49212,N_46214);
or UO_1404 (O_1404,N_49936,N_47091);
xor UO_1405 (O_1405,N_48152,N_45238);
nor UO_1406 (O_1406,N_45941,N_45798);
nand UO_1407 (O_1407,N_46615,N_48416);
and UO_1408 (O_1408,N_49267,N_45235);
and UO_1409 (O_1409,N_48800,N_46890);
nor UO_1410 (O_1410,N_48750,N_48952);
nor UO_1411 (O_1411,N_49195,N_47308);
xor UO_1412 (O_1412,N_45791,N_47690);
xnor UO_1413 (O_1413,N_49010,N_48989);
nor UO_1414 (O_1414,N_46467,N_46677);
or UO_1415 (O_1415,N_46825,N_49863);
xnor UO_1416 (O_1416,N_45276,N_48251);
xnor UO_1417 (O_1417,N_45463,N_47014);
and UO_1418 (O_1418,N_47653,N_45351);
nand UO_1419 (O_1419,N_48912,N_45526);
nand UO_1420 (O_1420,N_47743,N_49799);
or UO_1421 (O_1421,N_49891,N_49660);
nor UO_1422 (O_1422,N_45743,N_46721);
xnor UO_1423 (O_1423,N_48284,N_46844);
and UO_1424 (O_1424,N_49702,N_47744);
nand UO_1425 (O_1425,N_45281,N_48103);
xor UO_1426 (O_1426,N_45302,N_48903);
and UO_1427 (O_1427,N_48101,N_45860);
xnor UO_1428 (O_1428,N_48021,N_46007);
xor UO_1429 (O_1429,N_45584,N_47141);
and UO_1430 (O_1430,N_48843,N_49727);
nand UO_1431 (O_1431,N_47543,N_45443);
nor UO_1432 (O_1432,N_48934,N_49616);
xor UO_1433 (O_1433,N_48085,N_48953);
xor UO_1434 (O_1434,N_48678,N_47048);
or UO_1435 (O_1435,N_45183,N_49137);
or UO_1436 (O_1436,N_48123,N_45210);
nand UO_1437 (O_1437,N_49057,N_46389);
nand UO_1438 (O_1438,N_49474,N_46968);
nand UO_1439 (O_1439,N_49876,N_46012);
and UO_1440 (O_1440,N_47118,N_48844);
nand UO_1441 (O_1441,N_47047,N_46393);
nor UO_1442 (O_1442,N_47560,N_45286);
xor UO_1443 (O_1443,N_49599,N_48239);
nand UO_1444 (O_1444,N_46470,N_46531);
xor UO_1445 (O_1445,N_47672,N_49108);
nor UO_1446 (O_1446,N_49483,N_47471);
nand UO_1447 (O_1447,N_46909,N_49105);
xnor UO_1448 (O_1448,N_45898,N_46010);
xnor UO_1449 (O_1449,N_47290,N_46117);
or UO_1450 (O_1450,N_49620,N_45700);
nand UO_1451 (O_1451,N_47707,N_45296);
xor UO_1452 (O_1452,N_49392,N_45170);
nor UO_1453 (O_1453,N_48559,N_49656);
xnor UO_1454 (O_1454,N_47935,N_49694);
and UO_1455 (O_1455,N_46074,N_45415);
nor UO_1456 (O_1456,N_45901,N_48471);
nand UO_1457 (O_1457,N_45576,N_46631);
and UO_1458 (O_1458,N_47451,N_46235);
or UO_1459 (O_1459,N_46984,N_49682);
nor UO_1460 (O_1460,N_45358,N_48296);
or UO_1461 (O_1461,N_49557,N_47255);
nor UO_1462 (O_1462,N_49177,N_49895);
nor UO_1463 (O_1463,N_45623,N_48555);
or UO_1464 (O_1464,N_49369,N_49283);
nand UO_1465 (O_1465,N_49069,N_48749);
xor UO_1466 (O_1466,N_47589,N_49963);
and UO_1467 (O_1467,N_47052,N_48413);
xnor UO_1468 (O_1468,N_49586,N_46592);
xnor UO_1469 (O_1469,N_45500,N_49274);
nor UO_1470 (O_1470,N_49353,N_46795);
or UO_1471 (O_1471,N_46845,N_48608);
or UO_1472 (O_1472,N_45820,N_46725);
xnor UO_1473 (O_1473,N_48887,N_48135);
and UO_1474 (O_1474,N_46547,N_45319);
nor UO_1475 (O_1475,N_47634,N_49468);
and UO_1476 (O_1476,N_48066,N_45096);
or UO_1477 (O_1477,N_48746,N_48543);
nand UO_1478 (O_1478,N_46337,N_48344);
nand UO_1479 (O_1479,N_46394,N_48258);
or UO_1480 (O_1480,N_49952,N_48173);
nor UO_1481 (O_1481,N_46308,N_45537);
xor UO_1482 (O_1482,N_49260,N_47794);
xor UO_1483 (O_1483,N_46769,N_45516);
nand UO_1484 (O_1484,N_47112,N_45639);
or UO_1485 (O_1485,N_46436,N_46570);
and UO_1486 (O_1486,N_45032,N_48246);
xnor UO_1487 (O_1487,N_46632,N_47734);
or UO_1488 (O_1488,N_46481,N_46521);
nand UO_1489 (O_1489,N_45310,N_47053);
or UO_1490 (O_1490,N_45769,N_45104);
xnor UO_1491 (O_1491,N_49410,N_48326);
nand UO_1492 (O_1492,N_49470,N_49498);
or UO_1493 (O_1493,N_48600,N_48198);
nand UO_1494 (O_1494,N_45778,N_47870);
nor UO_1495 (O_1495,N_47320,N_45300);
or UO_1496 (O_1496,N_47754,N_46858);
nand UO_1497 (O_1497,N_46422,N_49521);
or UO_1498 (O_1498,N_49026,N_48944);
nand UO_1499 (O_1499,N_46401,N_49578);
nor UO_1500 (O_1500,N_49431,N_46954);
xnor UO_1501 (O_1501,N_49766,N_49476);
and UO_1502 (O_1502,N_45900,N_48769);
nor UO_1503 (O_1503,N_48349,N_47361);
xnor UO_1504 (O_1504,N_48920,N_47908);
and UO_1505 (O_1505,N_45084,N_47283);
or UO_1506 (O_1506,N_47497,N_48257);
and UO_1507 (O_1507,N_45308,N_47546);
nor UO_1508 (O_1508,N_47357,N_46688);
nand UO_1509 (O_1509,N_46098,N_48299);
xor UO_1510 (O_1510,N_49176,N_46781);
xnor UO_1511 (O_1511,N_49594,N_49118);
or UO_1512 (O_1512,N_49102,N_49361);
or UO_1513 (O_1513,N_45527,N_48567);
xor UO_1514 (O_1514,N_49163,N_46356);
or UO_1515 (O_1515,N_45627,N_47186);
nor UO_1516 (O_1516,N_47986,N_47962);
nor UO_1517 (O_1517,N_47339,N_48724);
or UO_1518 (O_1518,N_45564,N_47287);
nand UO_1519 (O_1519,N_49316,N_49677);
nor UO_1520 (O_1520,N_47058,N_49270);
xor UO_1521 (O_1521,N_47698,N_47885);
nor UO_1522 (O_1522,N_49852,N_46782);
or UO_1523 (O_1523,N_49512,N_46272);
nand UO_1524 (O_1524,N_49485,N_49773);
or UO_1525 (O_1525,N_49111,N_46917);
xnor UO_1526 (O_1526,N_49627,N_48771);
or UO_1527 (O_1527,N_49068,N_49096);
nand UO_1528 (O_1528,N_49191,N_49037);
nor UO_1529 (O_1529,N_45197,N_45377);
xor UO_1530 (O_1530,N_45367,N_46464);
nor UO_1531 (O_1531,N_47198,N_49802);
and UO_1532 (O_1532,N_48389,N_48183);
and UO_1533 (O_1533,N_48208,N_45539);
and UO_1534 (O_1534,N_46670,N_45506);
and UO_1535 (O_1535,N_48564,N_45928);
xnor UO_1536 (O_1536,N_45738,N_46529);
nor UO_1537 (O_1537,N_45764,N_47272);
nand UO_1538 (O_1538,N_49629,N_46468);
nand UO_1539 (O_1539,N_46504,N_45268);
and UO_1540 (O_1540,N_47671,N_47078);
nand UO_1541 (O_1541,N_48840,N_48087);
xnor UO_1542 (O_1542,N_46442,N_45856);
nand UO_1543 (O_1543,N_49444,N_46507);
nand UO_1544 (O_1544,N_49896,N_49770);
nand UO_1545 (O_1545,N_47140,N_45848);
nor UO_1546 (O_1546,N_45642,N_47635);
nor UO_1547 (O_1547,N_49875,N_45993);
nand UO_1548 (O_1548,N_47716,N_49303);
nand UO_1549 (O_1549,N_46509,N_46352);
xor UO_1550 (O_1550,N_45303,N_45217);
nand UO_1551 (O_1551,N_48272,N_48485);
nor UO_1552 (O_1552,N_48385,N_46663);
nand UO_1553 (O_1553,N_48013,N_48714);
and UO_1554 (O_1554,N_48377,N_46092);
or UO_1555 (O_1555,N_49387,N_48038);
xor UO_1556 (O_1556,N_49421,N_47245);
nand UO_1557 (O_1557,N_46621,N_46149);
nor UO_1558 (O_1558,N_47670,N_46817);
nor UO_1559 (O_1559,N_45043,N_45143);
nor UO_1560 (O_1560,N_46665,N_47518);
xnor UO_1561 (O_1561,N_46457,N_47978);
and UO_1562 (O_1562,N_47144,N_45332);
or UO_1563 (O_1563,N_47179,N_48683);
and UO_1564 (O_1564,N_47969,N_48375);
xor UO_1565 (O_1565,N_45513,N_45968);
xnor UO_1566 (O_1566,N_45669,N_46145);
or UO_1567 (O_1567,N_45649,N_49948);
and UO_1568 (O_1568,N_46992,N_45355);
xor UO_1569 (O_1569,N_48937,N_47254);
nand UO_1570 (O_1570,N_47648,N_46275);
nor UO_1571 (O_1571,N_46895,N_49537);
nand UO_1572 (O_1572,N_49703,N_46836);
nor UO_1573 (O_1573,N_49655,N_45862);
or UO_1574 (O_1574,N_46605,N_47821);
nand UO_1575 (O_1575,N_49249,N_48053);
nor UO_1576 (O_1576,N_48731,N_49420);
and UO_1577 (O_1577,N_45121,N_48886);
xor UO_1578 (O_1578,N_45890,N_49348);
nand UO_1579 (O_1579,N_48398,N_49635);
nor UO_1580 (O_1580,N_47526,N_46928);
nor UO_1581 (O_1581,N_47212,N_49091);
xor UO_1582 (O_1582,N_45727,N_45599);
nand UO_1583 (O_1583,N_47784,N_49540);
nand UO_1584 (O_1584,N_45551,N_46174);
and UO_1585 (O_1585,N_47501,N_45288);
xnor UO_1586 (O_1586,N_49756,N_46130);
or UO_1587 (O_1587,N_46551,N_46069);
nor UO_1588 (O_1588,N_48017,N_49595);
nand UO_1589 (O_1589,N_48380,N_45574);
and UO_1590 (O_1590,N_49633,N_48984);
or UO_1591 (O_1591,N_45590,N_47115);
xor UO_1592 (O_1592,N_48648,N_49907);
nor UO_1593 (O_1593,N_47466,N_45790);
and UO_1594 (O_1594,N_47046,N_47020);
xnor UO_1595 (O_1595,N_47106,N_47396);
nand UO_1596 (O_1596,N_47373,N_49022);
nand UO_1597 (O_1597,N_49236,N_46242);
and UO_1598 (O_1598,N_46094,N_46311);
xnor UO_1599 (O_1599,N_45829,N_49495);
or UO_1600 (O_1600,N_45730,N_48432);
nand UO_1601 (O_1601,N_45307,N_45646);
or UO_1602 (O_1602,N_49243,N_48006);
and UO_1603 (O_1603,N_45445,N_48440);
and UO_1604 (O_1604,N_47619,N_48546);
or UO_1605 (O_1605,N_45562,N_47034);
xor UO_1606 (O_1606,N_49268,N_47235);
and UO_1607 (O_1607,N_45836,N_49174);
nor UO_1608 (O_1608,N_45935,N_45994);
xor UO_1609 (O_1609,N_48213,N_48016);
nor UO_1610 (O_1610,N_49220,N_46798);
nor UO_1611 (O_1611,N_47164,N_49964);
or UO_1612 (O_1612,N_47017,N_49857);
nand UO_1613 (O_1613,N_49428,N_48679);
and UO_1614 (O_1614,N_49426,N_47638);
and UO_1615 (O_1615,N_46791,N_49882);
xnor UO_1616 (O_1616,N_49093,N_48715);
nand UO_1617 (O_1617,N_46295,N_45171);
nor UO_1618 (O_1618,N_46188,N_47104);
xor UO_1619 (O_1619,N_45372,N_46780);
xnor UO_1620 (O_1620,N_48305,N_45189);
xor UO_1621 (O_1621,N_47312,N_45996);
xnor UO_1622 (O_1622,N_48052,N_47951);
nor UO_1623 (O_1623,N_48157,N_49573);
nand UO_1624 (O_1624,N_48599,N_45720);
xnor UO_1625 (O_1625,N_46628,N_45647);
or UO_1626 (O_1626,N_49824,N_47005);
and UO_1627 (O_1627,N_45134,N_47689);
nand UO_1628 (O_1628,N_46625,N_47615);
nor UO_1629 (O_1629,N_45314,N_47434);
xor UO_1630 (O_1630,N_46081,N_48973);
or UO_1631 (O_1631,N_45681,N_47258);
or UO_1632 (O_1632,N_46255,N_47419);
or UO_1633 (O_1633,N_46203,N_49167);
nor UO_1634 (O_1634,N_47947,N_45593);
nand UO_1635 (O_1635,N_48635,N_47280);
or UO_1636 (O_1636,N_47472,N_49563);
nor UO_1637 (O_1637,N_49203,N_47065);
xor UO_1638 (O_1638,N_45896,N_46446);
nand UO_1639 (O_1639,N_49530,N_49342);
nor UO_1640 (O_1640,N_45475,N_45859);
nor UO_1641 (O_1641,N_47028,N_49442);
nand UO_1642 (O_1642,N_47400,N_45131);
nor UO_1643 (O_1643,N_45936,N_49760);
nand UO_1644 (O_1644,N_45002,N_49223);
xor UO_1645 (O_1645,N_49192,N_46602);
nor UO_1646 (O_1646,N_48039,N_48415);
nand UO_1647 (O_1647,N_46383,N_49151);
xnor UO_1648 (O_1648,N_48102,N_46340);
and UO_1649 (O_1649,N_47386,N_47229);
nor UO_1650 (O_1650,N_48445,N_47222);
and UO_1651 (O_1651,N_49979,N_48508);
xnor UO_1652 (O_1652,N_45325,N_46239);
and UO_1653 (O_1653,N_47613,N_49668);
and UO_1654 (O_1654,N_48493,N_47551);
nand UO_1655 (O_1655,N_46241,N_46708);
or UO_1656 (O_1656,N_48819,N_49104);
nand UO_1657 (O_1657,N_45466,N_49317);
xor UO_1658 (O_1658,N_47441,N_49240);
nand UO_1659 (O_1659,N_47731,N_49334);
or UO_1660 (O_1660,N_49396,N_49423);
or UO_1661 (O_1661,N_46133,N_49035);
and UO_1662 (O_1662,N_47169,N_46163);
and UO_1663 (O_1663,N_48141,N_45432);
or UO_1664 (O_1664,N_46008,N_46301);
xnor UO_1665 (O_1665,N_47529,N_49277);
nor UO_1666 (O_1666,N_48582,N_48187);
and UO_1667 (O_1667,N_49250,N_49033);
xnor UO_1668 (O_1668,N_48572,N_47490);
and UO_1669 (O_1669,N_47302,N_46997);
nor UO_1670 (O_1670,N_48230,N_45630);
nor UO_1671 (O_1671,N_45826,N_46914);
or UO_1672 (O_1672,N_49388,N_46420);
nor UO_1673 (O_1673,N_48361,N_49784);
nor UO_1674 (O_1674,N_45487,N_46675);
nand UO_1675 (O_1675,N_48708,N_48214);
or UO_1676 (O_1676,N_45373,N_48149);
nand UO_1677 (O_1677,N_47936,N_46166);
nand UO_1678 (O_1678,N_47858,N_47056);
nand UO_1679 (O_1679,N_47854,N_48824);
xnor UO_1680 (O_1680,N_48594,N_48365);
nor UO_1681 (O_1681,N_47187,N_47966);
and UO_1682 (O_1682,N_49509,N_49109);
xnor UO_1683 (O_1683,N_45480,N_45964);
nor UO_1684 (O_1684,N_45524,N_45449);
xor UO_1685 (O_1685,N_48831,N_48837);
or UO_1686 (O_1686,N_46395,N_46905);
and UO_1687 (O_1687,N_45153,N_49036);
and UO_1688 (O_1688,N_49436,N_47193);
nand UO_1689 (O_1689,N_48096,N_45948);
nand UO_1690 (O_1690,N_49939,N_45166);
and UO_1691 (O_1691,N_45828,N_47876);
and UO_1692 (O_1692,N_49508,N_48975);
nor UO_1693 (O_1693,N_46982,N_49950);
and UO_1694 (O_1694,N_45774,N_47410);
or UO_1695 (O_1695,N_45309,N_47367);
xor UO_1696 (O_1696,N_47820,N_45041);
or UO_1697 (O_1697,N_47607,N_47085);
nor UO_1698 (O_1698,N_49849,N_48629);
nor UO_1699 (O_1699,N_49161,N_45451);
nor UO_1700 (O_1700,N_47715,N_49230);
nor UO_1701 (O_1701,N_49507,N_48132);
or UO_1702 (O_1702,N_46931,N_46899);
or UO_1703 (O_1703,N_48182,N_45169);
nand UO_1704 (O_1704,N_47905,N_45245);
or UO_1705 (O_1705,N_46224,N_48397);
nor UO_1706 (O_1706,N_45601,N_49429);
and UO_1707 (O_1707,N_46949,N_45402);
nor UO_1708 (O_1708,N_48205,N_46111);
nand UO_1709 (O_1709,N_49541,N_45880);
xnor UO_1710 (O_1710,N_45881,N_47365);
xnor UO_1711 (O_1711,N_47940,N_46894);
nand UO_1712 (O_1712,N_47915,N_45409);
xnor UO_1713 (O_1713,N_46916,N_47700);
or UO_1714 (O_1714,N_45135,N_45492);
nor UO_1715 (O_1715,N_47404,N_45835);
nor UO_1716 (O_1716,N_49582,N_46205);
or UO_1717 (O_1717,N_48587,N_49506);
and UO_1718 (O_1718,N_47155,N_48004);
nor UO_1719 (O_1719,N_47796,N_48093);
nand UO_1720 (O_1720,N_48878,N_49103);
or UO_1721 (O_1721,N_46310,N_47830);
nand UO_1722 (O_1722,N_49395,N_45472);
and UO_1723 (O_1723,N_47934,N_46823);
xor UO_1724 (O_1724,N_46811,N_45916);
nor UO_1725 (O_1725,N_49908,N_49360);
and UO_1726 (O_1726,N_48333,N_46083);
and UO_1727 (O_1727,N_49503,N_49741);
nor UO_1728 (O_1728,N_48686,N_48857);
nand UO_1729 (O_1729,N_45076,N_49479);
nand UO_1730 (O_1730,N_48443,N_48591);
and UO_1731 (O_1731,N_46679,N_49867);
xnor UO_1732 (O_1732,N_46651,N_46983);
or UO_1733 (O_1733,N_45519,N_49123);
or UO_1734 (O_1734,N_48137,N_46710);
xnor UO_1735 (O_1735,N_48468,N_49765);
or UO_1736 (O_1736,N_47196,N_48790);
or UO_1737 (O_1737,N_46806,N_48484);
and UO_1738 (O_1738,N_45050,N_48935);
and UO_1739 (O_1739,N_49717,N_49816);
xnor UO_1740 (O_1740,N_47329,N_45436);
xor UO_1741 (O_1741,N_49736,N_48971);
or UO_1742 (O_1742,N_45323,N_45394);
nand UO_1743 (O_1743,N_46641,N_49107);
and UO_1744 (O_1744,N_45416,N_46689);
nand UO_1745 (O_1745,N_45866,N_45413);
nand UO_1746 (O_1746,N_46379,N_45410);
and UO_1747 (O_1747,N_47066,N_48118);
nor UO_1748 (O_1748,N_46556,N_47377);
nor UO_1749 (O_1749,N_48174,N_46114);
or UO_1750 (O_1750,N_45008,N_46097);
nor UO_1751 (O_1751,N_47515,N_45969);
and UO_1752 (O_1752,N_49048,N_49951);
xor UO_1753 (O_1753,N_45149,N_45103);
nand UO_1754 (O_1754,N_48890,N_45991);
nor UO_1755 (O_1755,N_47852,N_45047);
nor UO_1756 (O_1756,N_46597,N_48625);
nor UO_1757 (O_1757,N_47855,N_47297);
nor UO_1758 (O_1758,N_49490,N_45927);
nor UO_1759 (O_1759,N_46851,N_48474);
nand UO_1760 (O_1760,N_48991,N_46357);
xnor UO_1761 (O_1761,N_47833,N_47826);
and UO_1762 (O_1762,N_46594,N_48940);
or UO_1763 (O_1763,N_45825,N_46118);
xnor UO_1764 (O_1764,N_48580,N_45118);
xnor UO_1765 (O_1765,N_47426,N_49581);
or UO_1766 (O_1766,N_49465,N_48210);
xor UO_1767 (O_1767,N_45280,N_47499);
xor UO_1768 (O_1768,N_46869,N_47296);
or UO_1769 (O_1769,N_48954,N_45823);
nor UO_1770 (O_1770,N_47096,N_48510);
xor UO_1771 (O_1771,N_46546,N_47220);
nor UO_1772 (O_1772,N_49664,N_46091);
nor UO_1773 (O_1773,N_45376,N_47814);
nand UO_1774 (O_1774,N_45662,N_48467);
nand UO_1775 (O_1775,N_47556,N_49679);
or UO_1776 (O_1776,N_46563,N_48417);
nand UO_1777 (O_1777,N_48288,N_47205);
nor UO_1778 (O_1778,N_47877,N_46893);
nand UO_1779 (O_1779,N_49714,N_49991);
and UO_1780 (O_1780,N_48593,N_49955);
xnor UO_1781 (O_1781,N_48936,N_47545);
nand UO_1782 (O_1782,N_45811,N_46403);
and UO_1783 (O_1783,N_47366,N_45876);
nand UO_1784 (O_1784,N_45773,N_48088);
nand UO_1785 (O_1785,N_45787,N_45219);
or UO_1786 (O_1786,N_45284,N_45260);
xor UO_1787 (O_1787,N_49462,N_47311);
or UO_1788 (O_1788,N_48168,N_45248);
or UO_1789 (O_1789,N_47998,N_46883);
or UO_1790 (O_1790,N_47143,N_49205);
nor UO_1791 (O_1791,N_45105,N_45911);
nor UO_1792 (O_1792,N_47753,N_45789);
xnor UO_1793 (O_1793,N_47417,N_48523);
and UO_1794 (O_1794,N_47172,N_47679);
nor UO_1795 (O_1795,N_47694,N_46201);
nor UO_1796 (O_1796,N_46649,N_45814);
nor UO_1797 (O_1797,N_48544,N_47371);
nand UO_1798 (O_1798,N_48372,N_49811);
and UO_1799 (O_1799,N_48680,N_48964);
nand UO_1800 (O_1800,N_45982,N_49697);
xnor UO_1801 (O_1801,N_47123,N_49927);
xnor UO_1802 (O_1802,N_48489,N_46284);
and UO_1803 (O_1803,N_47949,N_46463);
and UO_1804 (O_1804,N_49803,N_46499);
and UO_1805 (O_1805,N_49935,N_48122);
xnor UO_1806 (O_1806,N_48563,N_48970);
or UO_1807 (O_1807,N_47808,N_45816);
nand UO_1808 (O_1808,N_45157,N_47674);
nand UO_1809 (O_1809,N_49152,N_49225);
nor UO_1810 (O_1810,N_48736,N_49040);
nand UO_1811 (O_1811,N_45628,N_48108);
xnor UO_1812 (O_1812,N_46598,N_45980);
or UO_1813 (O_1813,N_46619,N_47813);
nand UO_1814 (O_1814,N_48219,N_46185);
and UO_1815 (O_1815,N_45622,N_49866);
xor UO_1816 (O_1816,N_48335,N_45379);
xnor UO_1817 (O_1817,N_48454,N_46733);
nand UO_1818 (O_1818,N_49591,N_47862);
or UO_1819 (O_1819,N_47688,N_48332);
or UO_1820 (O_1820,N_48120,N_49795);
xnor UO_1821 (O_1821,N_46349,N_47552);
and UO_1822 (O_1822,N_47558,N_45100);
xnor UO_1823 (O_1823,N_47481,N_49710);
xor UO_1824 (O_1824,N_45243,N_46452);
nand UO_1825 (O_1825,N_47269,N_48562);
xor UO_1826 (O_1826,N_47127,N_47299);
xnor UO_1827 (O_1827,N_46263,N_48195);
nand UO_1828 (O_1828,N_48882,N_48740);
or UO_1829 (O_1829,N_48312,N_49219);
and UO_1830 (O_1830,N_49947,N_49084);
nand UO_1831 (O_1831,N_46450,N_46755);
nand UO_1832 (O_1832,N_47776,N_45831);
and UO_1833 (O_1833,N_49669,N_49847);
nand UO_1834 (O_1834,N_47783,N_48677);
nand UO_1835 (O_1835,N_49841,N_47617);
xnor UO_1836 (O_1836,N_48917,N_45930);
nand UO_1837 (O_1837,N_49693,N_47253);
and UO_1838 (O_1838,N_46473,N_46385);
and UO_1839 (O_1839,N_46388,N_46164);
nor UO_1840 (O_1840,N_46059,N_48022);
nor UO_1841 (O_1841,N_46041,N_49796);
and UO_1842 (O_1842,N_45979,N_49887);
nor UO_1843 (O_1843,N_49665,N_47326);
nor UO_1844 (O_1844,N_47345,N_48507);
and UO_1845 (O_1845,N_46444,N_46045);
and UO_1846 (O_1846,N_48762,N_48684);
nand UO_1847 (O_1847,N_49743,N_48927);
nand UO_1848 (O_1848,N_47234,N_49079);
xor UO_1849 (O_1849,N_45846,N_48895);
xnor UO_1850 (O_1850,N_48062,N_49565);
nor UO_1851 (O_1851,N_46377,N_46487);
xnor UO_1852 (O_1852,N_45059,N_46291);
nor UO_1853 (O_1853,N_45269,N_46684);
nand UO_1854 (O_1854,N_48658,N_47530);
nand UO_1855 (O_1855,N_46139,N_47766);
and UO_1856 (O_1856,N_49848,N_45083);
nand UO_1857 (O_1857,N_46696,N_48712);
and UO_1858 (O_1858,N_45538,N_49051);
nor UO_1859 (O_1859,N_47869,N_47692);
xor UO_1860 (O_1860,N_47509,N_48639);
nor UO_1861 (O_1861,N_46047,N_47457);
nor UO_1862 (O_1862,N_46608,N_45567);
and UO_1863 (O_1863,N_47811,N_49556);
nor UO_1864 (O_1864,N_46516,N_49333);
nand UO_1865 (O_1865,N_49897,N_46024);
nor UO_1866 (O_1866,N_45843,N_48479);
nand UO_1867 (O_1867,N_46033,N_47780);
or UO_1868 (O_1868,N_49588,N_47660);
nor UO_1869 (O_1869,N_47982,N_49472);
and UO_1870 (O_1870,N_45926,N_48106);
xor UO_1871 (O_1871,N_46199,N_47110);
or UO_1872 (O_1872,N_46852,N_48818);
nor UO_1873 (O_1873,N_46289,N_47156);
nor UO_1874 (O_1874,N_46217,N_48064);
and UO_1875 (O_1875,N_47459,N_46411);
nand UO_1876 (O_1876,N_49684,N_49063);
nor UO_1877 (O_1877,N_45239,N_45558);
nand UO_1878 (O_1878,N_46052,N_45090);
or UO_1879 (O_1879,N_46633,N_47887);
and UO_1880 (O_1880,N_49611,N_47249);
nor UO_1881 (O_1881,N_47268,N_49746);
nor UO_1882 (O_1882,N_46865,N_49505);
nor UO_1883 (O_1883,N_49536,N_48931);
xnor UO_1884 (O_1884,N_47943,N_45806);
nor UO_1885 (O_1885,N_45138,N_47890);
xor UO_1886 (O_1886,N_46202,N_46658);
nand UO_1887 (O_1887,N_46020,N_45644);
and UO_1888 (O_1888,N_45771,N_47159);
nor UO_1889 (O_1889,N_47738,N_45225);
nor UO_1890 (O_1890,N_48201,N_46271);
nand UO_1891 (O_1891,N_49047,N_47244);
nand UO_1892 (O_1892,N_48713,N_49001);
or UO_1893 (O_1893,N_46317,N_45651);
and UO_1894 (O_1894,N_46127,N_46986);
nor UO_1895 (O_1895,N_49978,N_46087);
or UO_1896 (O_1896,N_48516,N_46456);
and UO_1897 (O_1897,N_49959,N_46181);
and UO_1898 (O_1898,N_49932,N_48589);
nor UO_1899 (O_1899,N_49461,N_46885);
xor UO_1900 (O_1900,N_45442,N_45279);
nand UO_1901 (O_1901,N_45861,N_48905);
and UO_1902 (O_1902,N_46070,N_48897);
xnor UO_1903 (O_1903,N_48189,N_49870);
nand UO_1904 (O_1904,N_49737,N_45119);
nand UO_1905 (O_1905,N_47771,N_49546);
nor UO_1906 (O_1906,N_47807,N_46584);
xor UO_1907 (O_1907,N_47211,N_48669);
nor UO_1908 (O_1908,N_45142,N_46860);
and UO_1909 (O_1909,N_49757,N_48232);
or UO_1910 (O_1910,N_47040,N_49132);
nor UO_1911 (O_1911,N_47950,N_45174);
xnor UO_1912 (O_1912,N_47399,N_47507);
nand UO_1913 (O_1913,N_49764,N_48077);
or UO_1914 (O_1914,N_46342,N_48814);
nor UO_1915 (O_1915,N_49739,N_49050);
and UO_1916 (O_1916,N_49148,N_47621);
and UO_1917 (O_1917,N_46318,N_46472);
xnor UO_1918 (O_1918,N_45024,N_48261);
xor UO_1919 (O_1919,N_49956,N_48475);
xor UO_1920 (O_1920,N_47834,N_49284);
or UO_1921 (O_1921,N_49550,N_45917);
nand UO_1922 (O_1922,N_45181,N_49685);
xnor UO_1923 (O_1923,N_47089,N_46888);
xnor UO_1924 (O_1924,N_45594,N_45832);
nor UO_1925 (O_1925,N_47346,N_49320);
and UO_1926 (O_1926,N_49075,N_49280);
and UO_1927 (O_1927,N_48438,N_45934);
and UO_1928 (O_1928,N_48823,N_49335);
nor UO_1929 (O_1929,N_49817,N_47128);
nand UO_1930 (O_1930,N_49622,N_48460);
nor UO_1931 (O_1931,N_46162,N_45071);
and UO_1932 (O_1932,N_46712,N_47214);
nand UO_1933 (O_1933,N_47424,N_49885);
nor UO_1934 (O_1934,N_45932,N_47728);
and UO_1935 (O_1935,N_46475,N_47035);
and UO_1936 (O_1936,N_46657,N_49814);
xor UO_1937 (O_1937,N_45499,N_45536);
xor UO_1938 (O_1938,N_48623,N_49397);
xnor UO_1939 (O_1939,N_46830,N_49931);
and UO_1940 (O_1940,N_45973,N_45354);
nand UO_1941 (O_1941,N_46988,N_45586);
or UO_1942 (O_1942,N_47369,N_45049);
xor UO_1943 (O_1943,N_47676,N_48250);
nand UO_1944 (O_1944,N_46309,N_46674);
or UO_1945 (O_1945,N_46106,N_48788);
xnor UO_1946 (O_1946,N_48785,N_48435);
or UO_1947 (O_1947,N_48007,N_47135);
and UO_1948 (O_1948,N_46572,N_47837);
and UO_1949 (O_1949,N_49883,N_49566);
nand UO_1950 (O_1950,N_48551,N_45431);
or UO_1951 (O_1951,N_49748,N_45111);
nand UO_1952 (O_1952,N_46490,N_46582);
or UO_1953 (O_1953,N_47567,N_49328);
xor UO_1954 (O_1954,N_47077,N_47570);
and UO_1955 (O_1955,N_48707,N_46706);
xnor UO_1956 (O_1956,N_49082,N_47270);
nand UO_1957 (O_1957,N_48373,N_45477);
nand UO_1958 (O_1958,N_46148,N_48833);
nor UO_1959 (O_1959,N_49296,N_49623);
and UO_1960 (O_1960,N_45295,N_49319);
nor UO_1961 (O_1961,N_46664,N_48576);
nor UO_1962 (O_1962,N_49211,N_46549);
nand UO_1963 (O_1963,N_47263,N_47641);
or UO_1964 (O_1964,N_47129,N_45709);
xor UO_1965 (O_1965,N_46815,N_48748);
or UO_1966 (O_1966,N_45733,N_46789);
or UO_1967 (O_1967,N_49182,N_45575);
or UO_1968 (O_1968,N_47802,N_48845);
nor UO_1969 (O_1969,N_45467,N_48512);
nor UO_1970 (O_1970,N_47328,N_48362);
xnor UO_1971 (O_1971,N_47725,N_45550);
and UO_1972 (O_1972,N_47713,N_47498);
or UO_1973 (O_1973,N_46946,N_48846);
or UO_1974 (O_1974,N_49139,N_48848);
nand UO_1975 (O_1975,N_49781,N_49175);
nand UO_1976 (O_1976,N_46466,N_45092);
nor UO_1977 (O_1977,N_45618,N_47977);
nor UO_1978 (O_1978,N_45341,N_45414);
or UO_1979 (O_1979,N_48842,N_47579);
nor UO_1980 (O_1980,N_49357,N_47462);
xor UO_1981 (O_1981,N_47836,N_49538);
xnor UO_1982 (O_1982,N_45237,N_46128);
nor UO_1983 (O_1983,N_48472,N_46326);
xnor UO_1984 (O_1984,N_48148,N_49941);
xor UO_1985 (O_1985,N_47642,N_46068);
xnor UO_1986 (O_1986,N_47554,N_46766);
or UO_1987 (O_1987,N_45384,N_49608);
nand UO_1988 (O_1988,N_47177,N_47535);
nand UO_1989 (O_1989,N_49215,N_48447);
xnor UO_1990 (O_1990,N_45728,N_45285);
and UO_1991 (O_1991,N_46334,N_48170);
nor UO_1992 (O_1992,N_49295,N_45841);
nor UO_1993 (O_1993,N_45990,N_46427);
nor UO_1994 (O_1994,N_47176,N_49055);
xnor UO_1995 (O_1995,N_47896,N_47183);
or UO_1996 (O_1996,N_47608,N_49861);
or UO_1997 (O_1997,N_46119,N_48550);
nand UO_1998 (O_1998,N_48080,N_47502);
nand UO_1999 (O_1999,N_45578,N_49628);
or UO_2000 (O_2000,N_45391,N_47453);
and UO_2001 (O_2001,N_46764,N_48496);
nor UO_2002 (O_2002,N_47655,N_47395);
nand UO_2003 (O_2003,N_47610,N_49873);
or UO_2004 (O_2004,N_47932,N_48553);
and UO_2005 (O_2005,N_48504,N_45263);
and UO_2006 (O_2006,N_49106,N_46508);
and UO_2007 (O_2007,N_49020,N_49930);
nor UO_2008 (O_2008,N_47479,N_45592);
nand UO_2009 (O_2009,N_46426,N_46896);
or UO_2010 (O_2010,N_47657,N_49511);
xor UO_2011 (O_2011,N_49646,N_45231);
nor UO_2012 (O_2012,N_46901,N_48621);
or UO_2013 (O_2013,N_49141,N_46445);
nor UO_2014 (O_2014,N_46774,N_47749);
nand UO_2015 (O_2015,N_49165,N_45112);
nor UO_2016 (O_2016,N_48681,N_49923);
and UO_2017 (O_2017,N_46903,N_46939);
nor UO_2018 (O_2018,N_48889,N_45844);
or UO_2019 (O_2019,N_48347,N_46443);
xnor UO_2020 (O_2020,N_45333,N_49970);
nand UO_2021 (O_2021,N_45992,N_45348);
and UO_2022 (O_2022,N_48314,N_46236);
and UO_2023 (O_2023,N_46887,N_48154);
and UO_2024 (O_2024,N_49227,N_45779);
or UO_2025 (O_2025,N_48094,N_47376);
xor UO_2026 (O_2026,N_47282,N_45362);
and UO_2027 (O_2027,N_47563,N_47042);
and UO_2028 (O_2028,N_49643,N_45525);
nand UO_2029 (O_2029,N_48334,N_46206);
nand UO_2030 (O_2030,N_45146,N_47810);
or UO_2031 (O_2031,N_47914,N_46842);
nor UO_2032 (O_2032,N_45077,N_47955);
or UO_2033 (O_2033,N_45407,N_48511);
nor UO_2034 (O_2034,N_47919,N_48028);
nand UO_2035 (O_2035,N_49380,N_45029);
or UO_2036 (O_2036,N_46829,N_45797);
or UO_2037 (O_2037,N_48391,N_47473);
or UO_2038 (O_2038,N_48352,N_46571);
or UO_2039 (O_2039,N_46711,N_47382);
nand UO_2040 (O_2040,N_46990,N_49045);
nand UO_2041 (O_2041,N_47393,N_45230);
xnor UO_2042 (O_2042,N_45974,N_49775);
or UO_2043 (O_2043,N_46362,N_49463);
nand UO_2044 (O_2044,N_48040,N_46617);
nor UO_2045 (O_2045,N_47252,N_46036);
and UO_2046 (O_2046,N_49518,N_49374);
nor UO_2047 (O_2047,N_48967,N_45408);
nor UO_2048 (O_2048,N_49306,N_47532);
nor UO_2049 (O_2049,N_46662,N_48444);
and UO_2050 (O_2050,N_45396,N_46304);
nand UO_2051 (O_2051,N_48267,N_47505);
nor UO_2052 (O_2052,N_47388,N_46240);
and UO_2053 (O_2053,N_49751,N_46877);
xor UO_2054 (O_2054,N_47861,N_46160);
nor UO_2055 (O_2055,N_48611,N_49607);
and UO_2056 (O_2056,N_48861,N_45768);
xor UO_2057 (O_2057,N_47868,N_48363);
or UO_2058 (O_2058,N_46257,N_46064);
and UO_2059 (O_2059,N_45389,N_46078);
or UO_2060 (O_2060,N_48431,N_47663);
nand UO_2061 (O_2061,N_48265,N_46953);
or UO_2062 (O_2062,N_49838,N_48835);
nand UO_2063 (O_2063,N_47029,N_45203);
xor UO_2064 (O_2064,N_45765,N_48317);
nand UO_2065 (O_2065,N_49938,N_45206);
xnor UO_2066 (O_2066,N_45106,N_48834);
nor UO_2067 (O_2067,N_48337,N_49133);
and UO_2068 (O_2068,N_47352,N_46819);
xor UO_2069 (O_2069,N_49065,N_49641);
or UO_2070 (O_2070,N_49074,N_48100);
nand UO_2071 (O_2071,N_49168,N_46973);
nand UO_2072 (O_2072,N_45462,N_46534);
or UO_2073 (O_2073,N_48535,N_45523);
or UO_2074 (O_2074,N_47469,N_49042);
or UO_2075 (O_2075,N_47569,N_45763);
xor UO_2076 (O_2076,N_46614,N_45674);
xnor UO_2077 (O_2077,N_48941,N_48566);
nor UO_2078 (O_2078,N_48737,N_45694);
nor UO_2079 (O_2079,N_48194,N_46744);
and UO_2080 (O_2080,N_47659,N_47747);
nor UO_2081 (O_2081,N_48870,N_47348);
xor UO_2082 (O_2082,N_49619,N_49235);
and UO_2083 (O_2083,N_46159,N_45311);
nor UO_2084 (O_2084,N_46960,N_46216);
and UO_2085 (O_2085,N_47971,N_47461);
or UO_2086 (O_2086,N_47071,N_49062);
nand UO_2087 (O_2087,N_48908,N_47991);
xnor UO_2088 (O_2088,N_46154,N_49233);
and UO_2089 (O_2089,N_48911,N_45878);
or UO_2090 (O_2090,N_46832,N_47612);
and UO_2091 (O_2091,N_46963,N_47593);
nand UO_2092 (O_2092,N_49994,N_48248);
nor UO_2093 (O_2093,N_48615,N_45775);
nor UO_2094 (O_2094,N_46418,N_49502);
nor UO_2095 (O_2095,N_49099,N_47335);
or UO_2096 (O_2096,N_49836,N_45316);
xor UO_2097 (O_2097,N_48342,N_47464);
or UO_2098 (O_2098,N_45807,N_46550);
nand UO_2099 (O_2099,N_48071,N_46358);
nand UO_2100 (O_2100,N_45180,N_46243);
or UO_2101 (O_2101,N_45915,N_49179);
xnor UO_2102 (O_2102,N_45256,N_45556);
and UO_2103 (O_2103,N_48245,N_45678);
nor UO_2104 (O_2104,N_45454,N_49178);
nand UO_2105 (O_2105,N_48938,N_48864);
nand UO_2106 (O_2106,N_46415,N_46251);
or UO_2107 (O_2107,N_47666,N_48057);
nor UO_2108 (O_2108,N_46912,N_48672);
or UO_2109 (O_2109,N_48758,N_49253);
xor UO_2110 (O_2110,N_48282,N_48602);
nor UO_2111 (O_2111,N_49593,N_45919);
nor UO_2112 (O_2112,N_47122,N_48536);
or UO_2113 (O_2113,N_45717,N_48950);
nor UO_2114 (O_2114,N_45659,N_46786);
or UO_2115 (O_2115,N_46298,N_49597);
nor UO_2116 (O_2116,N_49516,N_46840);
or UO_2117 (O_2117,N_45855,N_46039);
nand UO_2118 (O_2118,N_48266,N_47279);
and UO_2119 (O_2119,N_49299,N_49583);
xor UO_2120 (O_2120,N_49860,N_47018);
xor UO_2121 (O_2121,N_48009,N_47597);
nor UO_2122 (O_2122,N_49218,N_48730);
or UO_2123 (O_2123,N_49053,N_45417);
nand UO_2124 (O_2124,N_48739,N_45895);
and UO_2125 (O_2125,N_45450,N_46691);
nand UO_2126 (O_2126,N_49881,N_45271);
nand UO_2127 (O_2127,N_45398,N_46157);
nor UO_2128 (O_2128,N_45329,N_47013);
or UO_2129 (O_2129,N_45251,N_49121);
or UO_2130 (O_2130,N_49752,N_48499);
nor UO_2131 (O_2131,N_45568,N_45511);
or UO_2132 (O_2132,N_46933,N_47818);
or UO_2133 (O_2133,N_45872,N_45289);
and UO_2134 (O_2134,N_49570,N_45741);
xor UO_2135 (O_2135,N_46419,N_47225);
and UO_2136 (O_2136,N_48359,N_45250);
or UO_2137 (O_2137,N_45240,N_45420);
or UO_2138 (O_2138,N_45486,N_47656);
nor UO_2139 (O_2139,N_46624,N_45989);
xnor UO_2140 (O_2140,N_46642,N_49455);
nor UO_2141 (O_2141,N_47640,N_47442);
nor UO_2142 (O_2142,N_45946,N_49282);
and UO_2143 (O_2143,N_47146,N_47664);
xnor UO_2144 (O_2144,N_46193,N_46682);
nor UO_2145 (O_2145,N_47082,N_47011);
xor UO_2146 (O_2146,N_45544,N_48619);
nor UO_2147 (O_2147,N_45474,N_49154);
xnor UO_2148 (O_2148,N_49124,N_47271);
nor UO_2149 (O_2149,N_45216,N_46184);
nor UO_2150 (O_2150,N_48346,N_48008);
and UO_2151 (O_2151,N_49992,N_48948);
and UO_2152 (O_2152,N_46707,N_45772);
nand UO_2153 (O_2153,N_49525,N_48316);
nand UO_2154 (O_2154,N_46503,N_49981);
nor UO_2155 (O_2155,N_45535,N_49602);
or UO_2156 (O_2156,N_46180,N_48744);
nand UO_2157 (O_2157,N_48434,N_49189);
and UO_2158 (O_2158,N_46279,N_47750);
nor UO_2159 (O_2159,N_48090,N_49197);
or UO_2160 (O_2160,N_46950,N_48875);
xor UO_2161 (O_2161,N_45504,N_49234);
and UO_2162 (O_2162,N_47741,N_48709);
and UO_2163 (O_2163,N_47675,N_47929);
and UO_2164 (O_2164,N_46741,N_49609);
nor UO_2165 (O_2165,N_48425,N_46049);
xnor UO_2166 (O_2166,N_48136,N_47007);
xor UO_2167 (O_2167,N_48537,N_49031);
or UO_2168 (O_2168,N_46269,N_46072);
and UO_2169 (O_2169,N_45139,N_49961);
nor UO_2170 (O_2170,N_47576,N_45265);
and UO_2171 (O_2171,N_48167,N_45906);
nand UO_2172 (O_2172,N_45158,N_46962);
nand UO_2173 (O_2173,N_45515,N_46669);
nand UO_2174 (O_2174,N_47899,N_45186);
or UO_2175 (O_2175,N_49183,N_46754);
and UO_2176 (O_2176,N_46095,N_47958);
and UO_2177 (O_2177,N_49683,N_48323);
xnor UO_2178 (O_2178,N_47431,N_49389);
xor UO_2179 (O_2179,N_49806,N_49571);
and UO_2180 (O_2180,N_47430,N_46253);
and UO_2181 (O_2181,N_45496,N_47705);
nand UO_2182 (O_2182,N_47148,N_48921);
xnor UO_2183 (O_2183,N_45693,N_46053);
or UO_2184 (O_2184,N_47792,N_46818);
nor UO_2185 (O_2185,N_48058,N_46940);
and UO_2186 (O_2186,N_49401,N_47801);
or UO_2187 (O_2187,N_48853,N_46713);
nand UO_2188 (O_2188,N_45440,N_48196);
nand UO_2189 (O_2189,N_47445,N_48427);
and UO_2190 (O_2190,N_46440,N_49614);
and UO_2191 (O_2191,N_45381,N_45483);
and UO_2192 (O_2192,N_45014,N_47521);
or UO_2193 (O_2193,N_48872,N_47098);
or UO_2194 (O_2194,N_48913,N_49718);
nand UO_2195 (O_2195,N_46122,N_46408);
or UO_2196 (O_2196,N_45446,N_45893);
nand UO_2197 (O_2197,N_49120,N_46897);
or UO_2198 (O_2198,N_45132,N_46132);
xnor UO_2199 (O_2199,N_48376,N_46519);
nor UO_2200 (O_2200,N_45560,N_46728);
xnor UO_2201 (O_2201,N_49734,N_49569);
or UO_2202 (O_2202,N_47064,N_45531);
nor UO_2203 (O_2203,N_46222,N_46283);
or UO_2204 (O_2204,N_46268,N_49721);
or UO_2205 (O_2205,N_49095,N_47414);
nor UO_2206 (O_2206,N_48171,N_46828);
nand UO_2207 (O_2207,N_45750,N_49100);
xor UO_2208 (O_2208,N_48476,N_48098);
xnor UO_2209 (O_2209,N_46557,N_47886);
or UO_2210 (O_2210,N_48985,N_45559);
nor UO_2211 (O_2211,N_47276,N_49258);
nor UO_2212 (O_2212,N_45484,N_49532);
or UO_2213 (O_2213,N_46672,N_48636);
xor UO_2214 (O_2214,N_48869,N_46338);
and UO_2215 (O_2215,N_48437,N_49587);
xor UO_2216 (O_2216,N_47427,N_45707);
or UO_2217 (O_2217,N_46331,N_47632);
nand UO_2218 (O_2218,N_48218,N_46831);
or UO_2219 (O_2219,N_48321,N_49081);
xnor UO_2220 (O_2220,N_45998,N_49753);
xnor UO_2221 (O_2221,N_48667,N_49957);
nor UO_2222 (O_2222,N_45986,N_47740);
and UO_2223 (O_2223,N_47240,N_45338);
and UO_2224 (O_2224,N_48048,N_46926);
xor UO_2225 (O_2225,N_49613,N_49661);
or UO_2226 (O_2226,N_45624,N_47428);
nor UO_2227 (O_2227,N_48585,N_45010);
nand UO_2228 (O_2228,N_47645,N_47259);
xor UO_2229 (O_2229,N_47781,N_45375);
nor UO_2230 (O_2230,N_46695,N_46123);
nand UO_2231 (O_2231,N_47549,N_45058);
nand UO_2232 (O_2232,N_46866,N_49858);
xor UO_2233 (O_2233,N_45960,N_47111);
nand UO_2234 (O_2234,N_47866,N_45494);
xnor UO_2235 (O_2235,N_45547,N_48439);
nor UO_2236 (O_2236,N_49590,N_46924);
nor UO_2237 (O_2237,N_46659,N_48783);
nand UO_2238 (O_2238,N_48545,N_47611);
and UO_2239 (O_2239,N_47174,N_49365);
nor UO_2240 (O_2240,N_46772,N_48634);
and UO_2241 (O_2241,N_48900,N_49797);
xnor UO_2242 (O_2242,N_47486,N_48227);
nor UO_2243 (O_2243,N_45699,N_47646);
xnor UO_2244 (O_2244,N_48598,N_49265);
nor UO_2245 (O_2245,N_45679,N_46762);
nor UO_2246 (O_2246,N_48308,N_47786);
and UO_2247 (O_2247,N_46985,N_48530);
nor UO_2248 (O_2248,N_46855,N_46668);
nand UO_2249 (O_2249,N_47379,N_45461);
or UO_2250 (O_2250,N_46262,N_45920);
nor UO_2251 (O_2251,N_46867,N_47232);
or UO_2252 (O_2252,N_45528,N_47673);
and UO_2253 (O_2253,N_47779,N_49318);
and UO_2254 (O_2254,N_46687,N_49954);
nand UO_2255 (O_2255,N_47755,N_45144);
and UO_2256 (O_2256,N_45360,N_47912);
nand UO_2257 (O_2257,N_46302,N_47954);
xnor UO_2258 (O_2258,N_45337,N_49384);
or UO_2259 (O_2259,N_48806,N_48901);
or UO_2260 (O_2260,N_49598,N_45004);
nand UO_2261 (O_2261,N_49321,N_46423);
xor UO_2262 (O_2262,N_47336,N_47409);
xnor UO_2263 (O_2263,N_47015,N_48805);
nand UO_2264 (O_2264,N_45495,N_48491);
and UO_2265 (O_2265,N_49995,N_45788);
and UO_2266 (O_2266,N_46878,N_45648);
nor UO_2267 (O_2267,N_46015,N_46025);
nor UO_2268 (O_2268,N_49073,N_49480);
nor UO_2269 (O_2269,N_45867,N_45542);
and UO_2270 (O_2270,N_48561,N_45840);
nor UO_2271 (O_2271,N_49626,N_46137);
and UO_2272 (O_2272,N_48575,N_47926);
nand UO_2273 (O_2273,N_48558,N_46397);
nor UO_2274 (O_2274,N_45518,N_49140);
nor UO_2275 (O_2275,N_45617,N_49076);
xnor UO_2276 (O_2276,N_47095,N_46042);
and UO_2277 (O_2277,N_45838,N_46850);
nor UO_2278 (O_2278,N_49681,N_49061);
and UO_2279 (O_2279,N_45130,N_49473);
and UO_2280 (O_2280,N_47816,N_45786);
xor UO_2281 (O_2281,N_48942,N_45549);
nor UO_2282 (O_2282,N_45987,N_46186);
nand UO_2283 (O_2283,N_49446,N_49691);
nor UO_2284 (O_2284,N_46034,N_49940);
and UO_2285 (O_2285,N_45705,N_48820);
xnor UO_2286 (O_2286,N_45988,N_48832);
xnor UO_2287 (O_2287,N_48358,N_48455);
nor UO_2288 (O_2288,N_46218,N_48692);
nand UO_2289 (O_2289,N_46676,N_49481);
or UO_2290 (O_2290,N_45107,N_46412);
xnor UO_2291 (O_2291,N_45621,N_49257);
nand UO_2292 (O_2292,N_47909,N_47360);
nor UO_2293 (O_2293,N_49676,N_47845);
nor UO_2294 (O_2294,N_49279,N_46112);
nor UO_2295 (O_2295,N_49386,N_46522);
or UO_2296 (O_2296,N_48193,N_46322);
or UO_2297 (O_2297,N_49343,N_47247);
or UO_2298 (O_2298,N_48656,N_45616);
or UO_2299 (O_2299,N_49572,N_46390);
nor UO_2300 (O_2300,N_48706,N_46787);
or UO_2301 (O_2301,N_49166,N_47819);
and UO_2302 (O_2302,N_45204,N_45085);
and UO_2303 (O_2303,N_47438,N_46841);
or UO_2304 (O_2304,N_46021,N_45301);
or UO_2305 (O_2305,N_49400,N_46437);
xnor UO_2306 (O_2306,N_47171,N_45177);
xor UO_2307 (O_2307,N_48311,N_49500);
xnor UO_2308 (O_2308,N_49405,N_46303);
nor UO_2309 (O_2309,N_47726,N_45199);
xor UO_2310 (O_2310,N_48097,N_49732);
or UO_2311 (O_2311,N_48287,N_45947);
nor UO_2312 (O_2312,N_47370,N_47050);
nand UO_2313 (O_2313,N_48211,N_45359);
and UO_2314 (O_2314,N_45716,N_46998);
and UO_2315 (O_2315,N_48357,N_47309);
nand UO_2316 (O_2316,N_48178,N_48121);
nor UO_2317 (O_2317,N_48753,N_47516);
nand UO_2318 (O_2318,N_46003,N_48162);
or UO_2319 (O_2319,N_46801,N_48411);
nor UO_2320 (O_2320,N_48972,N_47772);
xnor UO_2321 (O_2321,N_45438,N_47401);
nor UO_2322 (O_2322,N_47599,N_47033);
or UO_2323 (O_2323,N_46558,N_48770);
xor UO_2324 (O_2324,N_49539,N_47487);
or UO_2325 (O_2325,N_45246,N_46341);
nor UO_2326 (O_2326,N_48234,N_47618);
xnor UO_2327 (O_2327,N_48873,N_45404);
nand UO_2328 (O_2328,N_47093,N_47331);
and UO_2329 (O_2329,N_48778,N_45503);
and UO_2330 (O_2330,N_48099,N_48807);
or UO_2331 (O_2331,N_46943,N_47874);
xnor UO_2332 (O_2332,N_45459,N_46244);
nand UO_2333 (O_2333,N_46165,N_45795);
or UO_2334 (O_2334,N_49960,N_45689);
xor UO_2335 (O_2335,N_49202,N_48003);
or UO_2336 (O_2336,N_46553,N_47911);
xnor UO_2337 (O_2337,N_49919,N_45751);
nand UO_2338 (O_2338,N_45636,N_48628);
nor UO_2339 (O_2339,N_49304,N_46705);
nor UO_2340 (O_2340,N_48898,N_46252);
xnor UO_2341 (O_2341,N_48904,N_47721);
or UO_2342 (O_2342,N_47907,N_46913);
nand UO_2343 (O_2343,N_48336,N_47381);
nand UO_2344 (O_2344,N_45761,N_45722);
and UO_2345 (O_2345,N_49131,N_48742);
xor UO_2346 (O_2346,N_45421,N_45305);
nand UO_2347 (O_2347,N_48026,N_48893);
or UO_2348 (O_2348,N_48462,N_48761);
xor UO_2349 (O_2349,N_46576,N_46525);
nand UO_2350 (O_2350,N_47239,N_46569);
or UO_2351 (O_2351,N_48027,N_46293);
nor UO_2352 (O_2352,N_46246,N_45304);
xnor UO_2353 (O_2353,N_47162,N_47120);
nand UO_2354 (O_2354,N_48134,N_46030);
xnor UO_2355 (O_2355,N_46290,N_45060);
xor UO_2356 (O_2356,N_47152,N_47375);
nand UO_2357 (O_2357,N_47704,N_46667);
and UO_2358 (O_2358,N_45320,N_47622);
xnor UO_2359 (O_2359,N_47581,N_47087);
or UO_2360 (O_2360,N_45812,N_48259);
nand UO_2361 (O_2361,N_46813,N_45331);
or UO_2362 (O_2362,N_48717,N_48169);
nor UO_2363 (O_2363,N_46333,N_46328);
and UO_2364 (O_2364,N_47132,N_49424);
and UO_2365 (O_2365,N_49874,N_48220);
nor UO_2366 (O_2366,N_46560,N_46966);
nand UO_2367 (O_2367,N_46690,N_46589);
xor UO_2368 (O_2368,N_47536,N_48419);
nor UO_2369 (O_2369,N_46399,N_49142);
nand UO_2370 (O_2370,N_48620,N_47889);
and UO_2371 (O_2371,N_47274,N_45224);
xor UO_2372 (O_2372,N_45082,N_46227);
nand UO_2373 (O_2373,N_49358,N_49447);
and UO_2374 (O_2374,N_45912,N_49592);
xor UO_2375 (O_2375,N_47585,N_48812);
nor UO_2376 (O_2376,N_47898,N_49398);
nand UO_2377 (O_2377,N_48513,N_48032);
or UO_2378 (O_2378,N_48885,N_48078);
or UO_2379 (O_2379,N_46315,N_47333);
nand UO_2380 (O_2380,N_49605,N_49297);
or UO_2381 (O_2381,N_45009,N_48223);
xnor UO_2382 (O_2382,N_45637,N_46212);
or UO_2383 (O_2383,N_47765,N_48579);
or UO_2384 (O_2384,N_46266,N_49827);
xor UO_2385 (O_2385,N_49924,N_47305);
or UO_2386 (O_2386,N_48531,N_49554);
and UO_2387 (O_2387,N_45609,N_48768);
nor UO_2388 (O_2388,N_47097,N_45512);
and UO_2389 (O_2389,N_47055,N_49821);
xnor UO_2390 (O_2390,N_45266,N_45457);
or UO_2391 (O_2391,N_45198,N_48273);
or UO_2392 (O_2392,N_45334,N_47864);
nor UO_2393 (O_2393,N_48632,N_45802);
xnor UO_2394 (O_2394,N_49364,N_45581);
nand UO_2395 (O_2395,N_45087,N_46932);
nor UO_2396 (O_2396,N_49080,N_49113);
and UO_2397 (O_2397,N_49889,N_45453);
and UO_2398 (O_2398,N_49648,N_45194);
and UO_2399 (O_2399,N_49549,N_49822);
and UO_2400 (O_2400,N_47598,N_45035);
xnor UO_2401 (O_2401,N_48414,N_45742);
nand UO_2402 (O_2402,N_49671,N_48697);
nor UO_2403 (O_2403,N_45184,N_47022);
or UO_2404 (O_2404,N_49273,N_47124);
and UO_2405 (O_2405,N_47574,N_45053);
nor UO_2406 (O_2406,N_48808,N_49639);
or UO_2407 (O_2407,N_46936,N_45652);
xor UO_2408 (O_2408,N_46090,N_45762);
or UO_2409 (O_2409,N_49224,N_48307);
and UO_2410 (O_2410,N_46991,N_45711);
or UO_2411 (O_2411,N_46567,N_49879);
or UO_2412 (O_2412,N_49021,N_48548);
or UO_2413 (O_2413,N_45540,N_46219);
xnor UO_2414 (O_2414,N_48949,N_46848);
or UO_2415 (O_2415,N_49833,N_47101);
and UO_2416 (O_2416,N_48588,N_46486);
or UO_2417 (O_2417,N_49982,N_49286);
or UO_2418 (O_2418,N_46425,N_49313);
nor UO_2419 (O_2419,N_48185,N_49913);
nor UO_2420 (O_2420,N_49217,N_46778);
or UO_2421 (O_2421,N_48279,N_49517);
and UO_2422 (O_2422,N_45017,N_45668);
and UO_2423 (O_2423,N_47318,N_45970);
nand UO_2424 (O_2424,N_47293,N_45793);
or UO_2425 (O_2425,N_47341,N_48095);
or UO_2426 (O_2426,N_47974,N_45548);
xnor UO_2427 (O_2427,N_45759,N_46730);
nor UO_2428 (O_2428,N_47286,N_47421);
nor UO_2429 (O_2429,N_49344,N_47791);
and UO_2430 (O_2430,N_49890,N_47337);
nand UO_2431 (O_2431,N_46919,N_46994);
and UO_2432 (O_2432,N_46121,N_49902);
nor UO_2433 (O_2433,N_48957,N_46863);
or UO_2434 (O_2434,N_48115,N_47006);
nor UO_2435 (O_2435,N_47067,N_48277);
xnor UO_2436 (O_2436,N_46454,N_49196);
and UO_2437 (O_2437,N_47539,N_46610);
xnor UO_2438 (O_2438,N_45850,N_46838);
xnor UO_2439 (O_2439,N_48892,N_46835);
nor UO_2440 (O_2440,N_48688,N_48657);
and UO_2441 (O_2441,N_49878,N_46704);
or UO_2442 (O_2442,N_47968,N_49558);
and UO_2443 (O_2443,N_45545,N_47901);
nand UO_2444 (O_2444,N_49000,N_45726);
nand UO_2445 (O_2445,N_45108,N_48186);
xnor UO_2446 (O_2446,N_49564,N_46573);
nor UO_2447 (O_2447,N_47408,N_48617);
xnor UO_2448 (O_2448,N_46421,N_46958);
nand UO_2449 (O_2449,N_45356,N_49309);
nand UO_2450 (O_2450,N_49487,N_48392);
nor UO_2451 (O_2451,N_49086,N_47044);
xor UO_2452 (O_2452,N_45714,N_45735);
xor UO_2453 (O_2453,N_49143,N_46104);
nand UO_2454 (O_2454,N_49975,N_48318);
and UO_2455 (O_2455,N_49771,N_45393);
xnor UO_2456 (O_2456,N_48596,N_45328);
or UO_2457 (O_2457,N_49025,N_45794);
xor UO_2458 (O_2458,N_45097,N_46501);
and UO_2459 (O_2459,N_45660,N_45350);
nor UO_2460 (O_2460,N_46441,N_45098);
nor UO_2461 (O_2461,N_45580,N_49680);
and UO_2462 (O_2462,N_49524,N_45366);
xor UO_2463 (O_2463,N_47967,N_45447);
and UO_2464 (O_2464,N_47944,N_49548);
nor UO_2465 (O_2465,N_46510,N_49972);
nor UO_2466 (O_2466,N_45976,N_46797);
nand UO_2467 (O_2467,N_45321,N_47080);
nor UO_2468 (O_2468,N_49419,N_49709);
nand UO_2469 (O_2469,N_48138,N_47627);
nand UO_2470 (O_2470,N_47181,N_48104);
nand UO_2471 (O_2471,N_48723,N_45885);
or UO_2472 (O_2472,N_48453,N_45037);
nor UO_2473 (O_2473,N_46169,N_47520);
or UO_2474 (O_2474,N_49719,N_45274);
nor UO_2475 (O_2475,N_48828,N_45552);
or UO_2476 (O_2476,N_49742,N_48107);
nor UO_2477 (O_2477,N_45522,N_48774);
and UO_2478 (O_2478,N_47342,N_46096);
xnor UO_2479 (O_2479,N_49326,N_45128);
nand UO_2480 (O_2480,N_47812,N_46661);
and UO_2481 (O_2481,N_49460,N_49201);
nand UO_2482 (O_2482,N_45346,N_45619);
or UO_2483 (O_2483,N_47289,N_49933);
xnor UO_2484 (O_2484,N_45792,N_48151);
or UO_2485 (O_2485,N_48140,N_48653);
or UO_2486 (O_2486,N_45629,N_46431);
xnor UO_2487 (O_2487,N_45655,N_48224);
nand UO_2488 (O_2488,N_47777,N_47041);
nand UO_2489 (O_2489,N_49777,N_47972);
and UO_2490 (O_2490,N_49116,N_49425);
nand UO_2491 (O_2491,N_48128,N_48982);
nand UO_2492 (O_2492,N_48767,N_47204);
and UO_2493 (O_2493,N_49859,N_45151);
and UO_2494 (O_2494,N_47349,N_46967);
or UO_2495 (O_2495,N_47495,N_49634);
nor UO_2496 (O_2496,N_45352,N_48339);
and UO_2497 (O_2497,N_46297,N_48014);
or UO_2498 (O_2498,N_49934,N_46329);
xnor UO_2499 (O_2499,N_45222,N_45114);
nor UO_2500 (O_2500,N_48741,N_46190);
nand UO_2501 (O_2501,N_48716,N_47456);
or UO_2502 (O_2502,N_45772,N_46083);
or UO_2503 (O_2503,N_48900,N_45694);
and UO_2504 (O_2504,N_45297,N_46511);
xor UO_2505 (O_2505,N_46525,N_48772);
and UO_2506 (O_2506,N_47967,N_48709);
xnor UO_2507 (O_2507,N_49273,N_45342);
nor UO_2508 (O_2508,N_49649,N_47777);
or UO_2509 (O_2509,N_45356,N_45451);
or UO_2510 (O_2510,N_47918,N_46114);
and UO_2511 (O_2511,N_46254,N_48356);
nor UO_2512 (O_2512,N_46446,N_47974);
nor UO_2513 (O_2513,N_47271,N_46897);
or UO_2514 (O_2514,N_48591,N_47216);
nand UO_2515 (O_2515,N_46775,N_46312);
or UO_2516 (O_2516,N_46868,N_47661);
or UO_2517 (O_2517,N_47177,N_48434);
or UO_2518 (O_2518,N_46243,N_47659);
nand UO_2519 (O_2519,N_45398,N_46821);
nand UO_2520 (O_2520,N_49187,N_48928);
nand UO_2521 (O_2521,N_45261,N_45328);
nand UO_2522 (O_2522,N_47830,N_49308);
nor UO_2523 (O_2523,N_49097,N_46134);
nand UO_2524 (O_2524,N_45199,N_47564);
or UO_2525 (O_2525,N_46477,N_46734);
nor UO_2526 (O_2526,N_47030,N_47148);
or UO_2527 (O_2527,N_46751,N_45830);
xnor UO_2528 (O_2528,N_47361,N_45434);
nor UO_2529 (O_2529,N_48378,N_46956);
xnor UO_2530 (O_2530,N_48002,N_48888);
xor UO_2531 (O_2531,N_46860,N_48090);
xor UO_2532 (O_2532,N_45081,N_46965);
xor UO_2533 (O_2533,N_45423,N_46503);
xnor UO_2534 (O_2534,N_47360,N_46247);
nand UO_2535 (O_2535,N_47642,N_45238);
and UO_2536 (O_2536,N_45628,N_49552);
xnor UO_2537 (O_2537,N_46894,N_46507);
xnor UO_2538 (O_2538,N_48632,N_45151);
xor UO_2539 (O_2539,N_45877,N_45672);
and UO_2540 (O_2540,N_45363,N_46376);
and UO_2541 (O_2541,N_46629,N_47456);
nor UO_2542 (O_2542,N_49388,N_49758);
or UO_2543 (O_2543,N_49732,N_47825);
and UO_2544 (O_2544,N_46232,N_46602);
nor UO_2545 (O_2545,N_46000,N_46853);
nand UO_2546 (O_2546,N_48270,N_48271);
nor UO_2547 (O_2547,N_45167,N_49438);
xor UO_2548 (O_2548,N_48403,N_49746);
or UO_2549 (O_2549,N_48096,N_45185);
or UO_2550 (O_2550,N_49369,N_46816);
and UO_2551 (O_2551,N_48057,N_45457);
or UO_2552 (O_2552,N_49903,N_48624);
nor UO_2553 (O_2553,N_45969,N_48882);
nand UO_2554 (O_2554,N_45799,N_49728);
xnor UO_2555 (O_2555,N_48434,N_47300);
or UO_2556 (O_2556,N_49005,N_46981);
nand UO_2557 (O_2557,N_48512,N_47657);
nor UO_2558 (O_2558,N_45997,N_49656);
and UO_2559 (O_2559,N_47842,N_46766);
or UO_2560 (O_2560,N_49639,N_49761);
nand UO_2561 (O_2561,N_45211,N_48405);
nor UO_2562 (O_2562,N_46706,N_49581);
xnor UO_2563 (O_2563,N_49703,N_46833);
xor UO_2564 (O_2564,N_47550,N_49874);
nor UO_2565 (O_2565,N_48563,N_45952);
xnor UO_2566 (O_2566,N_48198,N_47221);
xnor UO_2567 (O_2567,N_48389,N_49941);
nand UO_2568 (O_2568,N_46394,N_49097);
xnor UO_2569 (O_2569,N_47994,N_46754);
or UO_2570 (O_2570,N_49887,N_49192);
or UO_2571 (O_2571,N_46491,N_45215);
and UO_2572 (O_2572,N_49398,N_46430);
nor UO_2573 (O_2573,N_48464,N_49121);
and UO_2574 (O_2574,N_48322,N_45542);
nand UO_2575 (O_2575,N_45883,N_48665);
xor UO_2576 (O_2576,N_47887,N_46925);
xnor UO_2577 (O_2577,N_48982,N_47676);
or UO_2578 (O_2578,N_45336,N_45172);
or UO_2579 (O_2579,N_46010,N_48004);
nand UO_2580 (O_2580,N_47003,N_47418);
nor UO_2581 (O_2581,N_49964,N_48296);
xor UO_2582 (O_2582,N_46626,N_47786);
nand UO_2583 (O_2583,N_46874,N_48353);
nor UO_2584 (O_2584,N_45454,N_46328);
and UO_2585 (O_2585,N_49486,N_45816);
and UO_2586 (O_2586,N_45013,N_46341);
and UO_2587 (O_2587,N_46093,N_47152);
nand UO_2588 (O_2588,N_49418,N_45824);
xor UO_2589 (O_2589,N_46734,N_46452);
xor UO_2590 (O_2590,N_45123,N_45014);
nor UO_2591 (O_2591,N_46948,N_46530);
or UO_2592 (O_2592,N_45404,N_46503);
nand UO_2593 (O_2593,N_47878,N_48428);
nand UO_2594 (O_2594,N_47513,N_48828);
xnor UO_2595 (O_2595,N_49625,N_47927);
nor UO_2596 (O_2596,N_46126,N_48407);
and UO_2597 (O_2597,N_47053,N_45222);
nand UO_2598 (O_2598,N_49248,N_47477);
xor UO_2599 (O_2599,N_49337,N_47408);
nand UO_2600 (O_2600,N_45676,N_46406);
xor UO_2601 (O_2601,N_45789,N_46105);
or UO_2602 (O_2602,N_48312,N_48934);
or UO_2603 (O_2603,N_49161,N_45673);
nand UO_2604 (O_2604,N_48108,N_45514);
nor UO_2605 (O_2605,N_48157,N_48879);
nand UO_2606 (O_2606,N_47933,N_46797);
xor UO_2607 (O_2607,N_45092,N_49492);
or UO_2608 (O_2608,N_48700,N_49184);
nor UO_2609 (O_2609,N_45744,N_45612);
xnor UO_2610 (O_2610,N_49705,N_47533);
or UO_2611 (O_2611,N_47984,N_47744);
nor UO_2612 (O_2612,N_46159,N_46841);
nor UO_2613 (O_2613,N_45738,N_49898);
nand UO_2614 (O_2614,N_49077,N_49042);
nor UO_2615 (O_2615,N_45135,N_46787);
nand UO_2616 (O_2616,N_47802,N_46041);
or UO_2617 (O_2617,N_46516,N_48801);
nor UO_2618 (O_2618,N_49453,N_48410);
or UO_2619 (O_2619,N_47121,N_45348);
nand UO_2620 (O_2620,N_48299,N_46404);
nor UO_2621 (O_2621,N_49736,N_45488);
and UO_2622 (O_2622,N_48273,N_46520);
xnor UO_2623 (O_2623,N_49821,N_46601);
and UO_2624 (O_2624,N_47242,N_46007);
xnor UO_2625 (O_2625,N_48488,N_45765);
xnor UO_2626 (O_2626,N_47491,N_45108);
and UO_2627 (O_2627,N_49886,N_45301);
nor UO_2628 (O_2628,N_45518,N_48644);
nor UO_2629 (O_2629,N_49473,N_48445);
nor UO_2630 (O_2630,N_46619,N_46464);
xor UO_2631 (O_2631,N_46198,N_46019);
nor UO_2632 (O_2632,N_48376,N_45937);
nor UO_2633 (O_2633,N_46840,N_45313);
nor UO_2634 (O_2634,N_48995,N_46232);
or UO_2635 (O_2635,N_46275,N_49284);
nand UO_2636 (O_2636,N_48510,N_47767);
nor UO_2637 (O_2637,N_46259,N_49731);
nor UO_2638 (O_2638,N_48775,N_45877);
xor UO_2639 (O_2639,N_49759,N_46303);
and UO_2640 (O_2640,N_48512,N_48381);
nor UO_2641 (O_2641,N_45522,N_47346);
or UO_2642 (O_2642,N_48863,N_48400);
and UO_2643 (O_2643,N_48309,N_46716);
nor UO_2644 (O_2644,N_48423,N_48025);
nand UO_2645 (O_2645,N_45465,N_45213);
xor UO_2646 (O_2646,N_49138,N_45893);
or UO_2647 (O_2647,N_47679,N_46286);
or UO_2648 (O_2648,N_47674,N_45895);
and UO_2649 (O_2649,N_47316,N_46937);
or UO_2650 (O_2650,N_45244,N_46649);
nor UO_2651 (O_2651,N_47468,N_46653);
or UO_2652 (O_2652,N_45229,N_49077);
nand UO_2653 (O_2653,N_45170,N_47727);
xor UO_2654 (O_2654,N_49641,N_47152);
and UO_2655 (O_2655,N_49832,N_48404);
xor UO_2656 (O_2656,N_47167,N_46770);
nand UO_2657 (O_2657,N_47488,N_46466);
xnor UO_2658 (O_2658,N_46551,N_47683);
nor UO_2659 (O_2659,N_47143,N_49164);
or UO_2660 (O_2660,N_45702,N_47516);
and UO_2661 (O_2661,N_49212,N_45774);
nor UO_2662 (O_2662,N_47145,N_49510);
or UO_2663 (O_2663,N_47230,N_47682);
and UO_2664 (O_2664,N_49222,N_48413);
nand UO_2665 (O_2665,N_49546,N_47787);
or UO_2666 (O_2666,N_47223,N_46764);
nand UO_2667 (O_2667,N_46768,N_45312);
or UO_2668 (O_2668,N_46738,N_45005);
and UO_2669 (O_2669,N_48338,N_49015);
or UO_2670 (O_2670,N_48804,N_47764);
and UO_2671 (O_2671,N_48404,N_46607);
xnor UO_2672 (O_2672,N_48282,N_49622);
nor UO_2673 (O_2673,N_46908,N_49658);
nand UO_2674 (O_2674,N_48397,N_47175);
xnor UO_2675 (O_2675,N_49554,N_48794);
or UO_2676 (O_2676,N_48129,N_49521);
nor UO_2677 (O_2677,N_46164,N_49782);
xnor UO_2678 (O_2678,N_47687,N_48965);
xnor UO_2679 (O_2679,N_45904,N_46346);
or UO_2680 (O_2680,N_45984,N_45385);
xnor UO_2681 (O_2681,N_48672,N_49801);
or UO_2682 (O_2682,N_48687,N_46052);
xnor UO_2683 (O_2683,N_45507,N_47684);
xor UO_2684 (O_2684,N_47680,N_46401);
and UO_2685 (O_2685,N_45806,N_47472);
and UO_2686 (O_2686,N_49630,N_47219);
or UO_2687 (O_2687,N_47300,N_48859);
nor UO_2688 (O_2688,N_49072,N_45607);
xor UO_2689 (O_2689,N_48959,N_47382);
or UO_2690 (O_2690,N_48157,N_49125);
xnor UO_2691 (O_2691,N_49222,N_48245);
nand UO_2692 (O_2692,N_45917,N_48586);
and UO_2693 (O_2693,N_48170,N_49858);
nor UO_2694 (O_2694,N_48488,N_46213);
and UO_2695 (O_2695,N_48405,N_45638);
and UO_2696 (O_2696,N_47914,N_49388);
or UO_2697 (O_2697,N_47074,N_45626);
and UO_2698 (O_2698,N_49332,N_47291);
or UO_2699 (O_2699,N_48731,N_45651);
or UO_2700 (O_2700,N_46251,N_45964);
xnor UO_2701 (O_2701,N_49099,N_47790);
and UO_2702 (O_2702,N_46359,N_48683);
and UO_2703 (O_2703,N_47184,N_45344);
xor UO_2704 (O_2704,N_46802,N_45226);
nor UO_2705 (O_2705,N_48168,N_48890);
xor UO_2706 (O_2706,N_49359,N_48138);
nor UO_2707 (O_2707,N_46224,N_49766);
or UO_2708 (O_2708,N_46005,N_47536);
nor UO_2709 (O_2709,N_45046,N_46456);
nand UO_2710 (O_2710,N_46768,N_49076);
nor UO_2711 (O_2711,N_47686,N_49235);
nor UO_2712 (O_2712,N_47733,N_48046);
or UO_2713 (O_2713,N_48757,N_46248);
nor UO_2714 (O_2714,N_49849,N_49864);
nor UO_2715 (O_2715,N_46890,N_46328);
or UO_2716 (O_2716,N_49401,N_49746);
and UO_2717 (O_2717,N_48146,N_47641);
nand UO_2718 (O_2718,N_46157,N_48218);
xnor UO_2719 (O_2719,N_45681,N_49568);
nand UO_2720 (O_2720,N_49937,N_46464);
nor UO_2721 (O_2721,N_49044,N_49507);
or UO_2722 (O_2722,N_47318,N_49248);
and UO_2723 (O_2723,N_47042,N_45135);
nor UO_2724 (O_2724,N_46377,N_45752);
or UO_2725 (O_2725,N_48555,N_45435);
nor UO_2726 (O_2726,N_48487,N_45254);
and UO_2727 (O_2727,N_47541,N_46964);
nand UO_2728 (O_2728,N_45392,N_46830);
xnor UO_2729 (O_2729,N_45092,N_49273);
xor UO_2730 (O_2730,N_48899,N_49209);
nand UO_2731 (O_2731,N_46324,N_47719);
nor UO_2732 (O_2732,N_48759,N_49118);
xor UO_2733 (O_2733,N_45718,N_47184);
or UO_2734 (O_2734,N_46128,N_46865);
xnor UO_2735 (O_2735,N_49471,N_49525);
nand UO_2736 (O_2736,N_45818,N_46895);
or UO_2737 (O_2737,N_47756,N_47454);
and UO_2738 (O_2738,N_45943,N_49480);
or UO_2739 (O_2739,N_48575,N_49412);
nor UO_2740 (O_2740,N_46674,N_48118);
xnor UO_2741 (O_2741,N_47371,N_46642);
nand UO_2742 (O_2742,N_47982,N_48641);
and UO_2743 (O_2743,N_49142,N_49648);
nand UO_2744 (O_2744,N_49713,N_45299);
xnor UO_2745 (O_2745,N_49305,N_48855);
xor UO_2746 (O_2746,N_45722,N_45743);
and UO_2747 (O_2747,N_49276,N_45452);
nor UO_2748 (O_2748,N_45114,N_47558);
and UO_2749 (O_2749,N_47664,N_49859);
and UO_2750 (O_2750,N_45652,N_47992);
and UO_2751 (O_2751,N_47331,N_47257);
nor UO_2752 (O_2752,N_46576,N_46740);
or UO_2753 (O_2753,N_48163,N_45347);
or UO_2754 (O_2754,N_45055,N_46282);
xor UO_2755 (O_2755,N_49745,N_47391);
xnor UO_2756 (O_2756,N_47206,N_48319);
and UO_2757 (O_2757,N_45211,N_45328);
xnor UO_2758 (O_2758,N_45409,N_47251);
xnor UO_2759 (O_2759,N_48597,N_47013);
or UO_2760 (O_2760,N_45742,N_46998);
nand UO_2761 (O_2761,N_49974,N_45276);
and UO_2762 (O_2762,N_46028,N_46890);
or UO_2763 (O_2763,N_46573,N_46213);
and UO_2764 (O_2764,N_45494,N_45516);
or UO_2765 (O_2765,N_46691,N_48368);
or UO_2766 (O_2766,N_47543,N_46221);
xnor UO_2767 (O_2767,N_45910,N_47729);
nor UO_2768 (O_2768,N_49433,N_46003);
or UO_2769 (O_2769,N_45023,N_48339);
xnor UO_2770 (O_2770,N_47747,N_47300);
or UO_2771 (O_2771,N_49577,N_46177);
and UO_2772 (O_2772,N_48056,N_49756);
xor UO_2773 (O_2773,N_49605,N_48703);
and UO_2774 (O_2774,N_46977,N_45536);
xor UO_2775 (O_2775,N_46923,N_47375);
nor UO_2776 (O_2776,N_46158,N_48195);
nor UO_2777 (O_2777,N_46656,N_49901);
nor UO_2778 (O_2778,N_48208,N_45490);
or UO_2779 (O_2779,N_47935,N_47232);
nor UO_2780 (O_2780,N_45956,N_46882);
and UO_2781 (O_2781,N_48387,N_47652);
nor UO_2782 (O_2782,N_46899,N_46396);
or UO_2783 (O_2783,N_45622,N_46630);
xnor UO_2784 (O_2784,N_46573,N_47348);
nand UO_2785 (O_2785,N_48329,N_45637);
nand UO_2786 (O_2786,N_47712,N_47860);
nor UO_2787 (O_2787,N_49389,N_47198);
and UO_2788 (O_2788,N_45966,N_49883);
or UO_2789 (O_2789,N_48471,N_45573);
or UO_2790 (O_2790,N_47789,N_48980);
xnor UO_2791 (O_2791,N_45699,N_49022);
nand UO_2792 (O_2792,N_48208,N_48909);
or UO_2793 (O_2793,N_46313,N_46375);
nor UO_2794 (O_2794,N_48825,N_49377);
nor UO_2795 (O_2795,N_47946,N_46839);
xor UO_2796 (O_2796,N_46547,N_48340);
xor UO_2797 (O_2797,N_46234,N_48214);
or UO_2798 (O_2798,N_45096,N_47687);
or UO_2799 (O_2799,N_47716,N_46697);
nor UO_2800 (O_2800,N_48898,N_49260);
nand UO_2801 (O_2801,N_49080,N_45844);
and UO_2802 (O_2802,N_45632,N_47359);
nand UO_2803 (O_2803,N_48310,N_48161);
and UO_2804 (O_2804,N_48330,N_46218);
nand UO_2805 (O_2805,N_49377,N_45141);
or UO_2806 (O_2806,N_46044,N_49935);
or UO_2807 (O_2807,N_48298,N_45185);
and UO_2808 (O_2808,N_48356,N_47097);
or UO_2809 (O_2809,N_46789,N_45701);
and UO_2810 (O_2810,N_46680,N_48836);
nor UO_2811 (O_2811,N_45741,N_46169);
and UO_2812 (O_2812,N_47492,N_49828);
and UO_2813 (O_2813,N_48077,N_45495);
or UO_2814 (O_2814,N_45421,N_46791);
and UO_2815 (O_2815,N_45776,N_49889);
nor UO_2816 (O_2816,N_48292,N_46318);
and UO_2817 (O_2817,N_49587,N_45142);
or UO_2818 (O_2818,N_48921,N_47353);
or UO_2819 (O_2819,N_46472,N_49213);
nand UO_2820 (O_2820,N_45993,N_49949);
or UO_2821 (O_2821,N_47653,N_45050);
nor UO_2822 (O_2822,N_49269,N_47830);
or UO_2823 (O_2823,N_45070,N_46639);
nor UO_2824 (O_2824,N_47247,N_47706);
nor UO_2825 (O_2825,N_46846,N_47289);
or UO_2826 (O_2826,N_48810,N_48504);
xor UO_2827 (O_2827,N_49413,N_47511);
xor UO_2828 (O_2828,N_49173,N_45811);
nor UO_2829 (O_2829,N_48559,N_48388);
nand UO_2830 (O_2830,N_46670,N_47759);
nand UO_2831 (O_2831,N_48985,N_47282);
nand UO_2832 (O_2832,N_45106,N_48816);
nand UO_2833 (O_2833,N_45146,N_48908);
nor UO_2834 (O_2834,N_46345,N_49692);
nor UO_2835 (O_2835,N_49718,N_47972);
and UO_2836 (O_2836,N_48977,N_46875);
nand UO_2837 (O_2837,N_45560,N_49444);
or UO_2838 (O_2838,N_49387,N_48014);
or UO_2839 (O_2839,N_48949,N_45894);
nor UO_2840 (O_2840,N_46909,N_49153);
nand UO_2841 (O_2841,N_45743,N_46814);
nor UO_2842 (O_2842,N_48614,N_49868);
xnor UO_2843 (O_2843,N_48079,N_49492);
and UO_2844 (O_2844,N_47516,N_48875);
or UO_2845 (O_2845,N_47741,N_48608);
or UO_2846 (O_2846,N_47662,N_49906);
xnor UO_2847 (O_2847,N_47571,N_46336);
nand UO_2848 (O_2848,N_47005,N_48635);
nor UO_2849 (O_2849,N_47939,N_45543);
nor UO_2850 (O_2850,N_45108,N_47719);
xnor UO_2851 (O_2851,N_46782,N_49176);
and UO_2852 (O_2852,N_45800,N_47243);
nand UO_2853 (O_2853,N_48749,N_48557);
and UO_2854 (O_2854,N_48125,N_49724);
xor UO_2855 (O_2855,N_45880,N_48549);
and UO_2856 (O_2856,N_45341,N_47913);
or UO_2857 (O_2857,N_49330,N_47987);
nor UO_2858 (O_2858,N_45491,N_49920);
nand UO_2859 (O_2859,N_49861,N_49335);
or UO_2860 (O_2860,N_46872,N_48794);
nor UO_2861 (O_2861,N_45083,N_48096);
and UO_2862 (O_2862,N_46795,N_49081);
xnor UO_2863 (O_2863,N_45623,N_45636);
xor UO_2864 (O_2864,N_46591,N_48493);
or UO_2865 (O_2865,N_49856,N_48710);
nor UO_2866 (O_2866,N_48673,N_47682);
or UO_2867 (O_2867,N_47178,N_47068);
and UO_2868 (O_2868,N_47979,N_47358);
nand UO_2869 (O_2869,N_49533,N_49753);
and UO_2870 (O_2870,N_47896,N_49324);
or UO_2871 (O_2871,N_47268,N_46665);
and UO_2872 (O_2872,N_45586,N_45850);
or UO_2873 (O_2873,N_45253,N_47792);
nand UO_2874 (O_2874,N_47334,N_46281);
and UO_2875 (O_2875,N_46898,N_46641);
nor UO_2876 (O_2876,N_49404,N_45957);
nand UO_2877 (O_2877,N_47096,N_45435);
xor UO_2878 (O_2878,N_49382,N_48698);
and UO_2879 (O_2879,N_49927,N_48752);
nor UO_2880 (O_2880,N_48118,N_49822);
nand UO_2881 (O_2881,N_48132,N_45689);
or UO_2882 (O_2882,N_48969,N_48951);
xor UO_2883 (O_2883,N_45893,N_46862);
and UO_2884 (O_2884,N_48157,N_46656);
nor UO_2885 (O_2885,N_48425,N_49344);
nand UO_2886 (O_2886,N_45018,N_45242);
or UO_2887 (O_2887,N_49629,N_49471);
nand UO_2888 (O_2888,N_46935,N_47004);
nand UO_2889 (O_2889,N_48635,N_49427);
nand UO_2890 (O_2890,N_45198,N_49831);
or UO_2891 (O_2891,N_46973,N_46482);
xor UO_2892 (O_2892,N_47015,N_45579);
nor UO_2893 (O_2893,N_48473,N_45100);
and UO_2894 (O_2894,N_49622,N_47894);
and UO_2895 (O_2895,N_46900,N_45237);
xnor UO_2896 (O_2896,N_49218,N_45521);
nor UO_2897 (O_2897,N_45050,N_45403);
xnor UO_2898 (O_2898,N_49200,N_46378);
or UO_2899 (O_2899,N_48140,N_46852);
nor UO_2900 (O_2900,N_49190,N_45102);
nor UO_2901 (O_2901,N_48171,N_45018);
and UO_2902 (O_2902,N_46063,N_46396);
and UO_2903 (O_2903,N_46778,N_49839);
nor UO_2904 (O_2904,N_48509,N_49340);
xor UO_2905 (O_2905,N_45058,N_45362);
xnor UO_2906 (O_2906,N_45157,N_45329);
nor UO_2907 (O_2907,N_46195,N_46296);
nand UO_2908 (O_2908,N_48545,N_46478);
xor UO_2909 (O_2909,N_46079,N_47496);
xor UO_2910 (O_2910,N_45376,N_48603);
or UO_2911 (O_2911,N_46216,N_45889);
and UO_2912 (O_2912,N_48295,N_47546);
xnor UO_2913 (O_2913,N_45930,N_48807);
xor UO_2914 (O_2914,N_47371,N_45454);
xor UO_2915 (O_2915,N_48101,N_47319);
xor UO_2916 (O_2916,N_46515,N_49470);
xnor UO_2917 (O_2917,N_45147,N_48942);
xnor UO_2918 (O_2918,N_45963,N_48665);
and UO_2919 (O_2919,N_49391,N_45485);
nand UO_2920 (O_2920,N_45032,N_45053);
nor UO_2921 (O_2921,N_48707,N_48623);
or UO_2922 (O_2922,N_45678,N_49656);
nand UO_2923 (O_2923,N_46269,N_46298);
nand UO_2924 (O_2924,N_48366,N_47385);
xnor UO_2925 (O_2925,N_46372,N_48775);
and UO_2926 (O_2926,N_45862,N_45013);
and UO_2927 (O_2927,N_45183,N_49196);
nand UO_2928 (O_2928,N_48643,N_49504);
nor UO_2929 (O_2929,N_48988,N_49250);
or UO_2930 (O_2930,N_45618,N_49455);
and UO_2931 (O_2931,N_47688,N_45836);
xnor UO_2932 (O_2932,N_46185,N_48422);
or UO_2933 (O_2933,N_49532,N_48821);
and UO_2934 (O_2934,N_48184,N_45956);
nor UO_2935 (O_2935,N_48884,N_46935);
and UO_2936 (O_2936,N_49145,N_46811);
and UO_2937 (O_2937,N_47268,N_48099);
nor UO_2938 (O_2938,N_47711,N_47603);
or UO_2939 (O_2939,N_45557,N_46236);
nand UO_2940 (O_2940,N_49396,N_47721);
nor UO_2941 (O_2941,N_46125,N_47675);
nand UO_2942 (O_2942,N_49341,N_48765);
or UO_2943 (O_2943,N_48155,N_46347);
nor UO_2944 (O_2944,N_45374,N_45685);
nor UO_2945 (O_2945,N_49474,N_47799);
xnor UO_2946 (O_2946,N_49184,N_47025);
nand UO_2947 (O_2947,N_45190,N_46947);
xnor UO_2948 (O_2948,N_46471,N_46886);
nand UO_2949 (O_2949,N_49490,N_45433);
xor UO_2950 (O_2950,N_47798,N_45371);
nor UO_2951 (O_2951,N_48785,N_47573);
nand UO_2952 (O_2952,N_48936,N_46055);
nand UO_2953 (O_2953,N_49308,N_45491);
xor UO_2954 (O_2954,N_48162,N_45838);
nor UO_2955 (O_2955,N_46839,N_47536);
nand UO_2956 (O_2956,N_48736,N_45239);
and UO_2957 (O_2957,N_48548,N_47370);
or UO_2958 (O_2958,N_45423,N_48070);
or UO_2959 (O_2959,N_49354,N_47624);
or UO_2960 (O_2960,N_47523,N_47023);
xor UO_2961 (O_2961,N_45067,N_48083);
or UO_2962 (O_2962,N_47983,N_48595);
nand UO_2963 (O_2963,N_47231,N_49078);
or UO_2964 (O_2964,N_46563,N_49473);
nor UO_2965 (O_2965,N_45782,N_49583);
xor UO_2966 (O_2966,N_49104,N_48773);
nor UO_2967 (O_2967,N_48999,N_46768);
and UO_2968 (O_2968,N_48604,N_48432);
nand UO_2969 (O_2969,N_49912,N_47299);
nor UO_2970 (O_2970,N_49303,N_46452);
nand UO_2971 (O_2971,N_45931,N_47753);
xor UO_2972 (O_2972,N_48851,N_48330);
and UO_2973 (O_2973,N_49930,N_49050);
or UO_2974 (O_2974,N_47764,N_48936);
or UO_2975 (O_2975,N_48924,N_49770);
xnor UO_2976 (O_2976,N_49902,N_46398);
and UO_2977 (O_2977,N_46583,N_48230);
xor UO_2978 (O_2978,N_45870,N_47028);
nand UO_2979 (O_2979,N_46919,N_49259);
or UO_2980 (O_2980,N_45720,N_49712);
or UO_2981 (O_2981,N_47131,N_49221);
nand UO_2982 (O_2982,N_45984,N_47266);
nand UO_2983 (O_2983,N_45209,N_49411);
nor UO_2984 (O_2984,N_46095,N_49393);
nand UO_2985 (O_2985,N_47962,N_45844);
nor UO_2986 (O_2986,N_45301,N_48822);
xor UO_2987 (O_2987,N_46938,N_46669);
xor UO_2988 (O_2988,N_45851,N_47975);
or UO_2989 (O_2989,N_48640,N_45592);
or UO_2990 (O_2990,N_47929,N_47763);
xnor UO_2991 (O_2991,N_46830,N_49754);
xnor UO_2992 (O_2992,N_48643,N_45932);
or UO_2993 (O_2993,N_46575,N_49524);
xnor UO_2994 (O_2994,N_45707,N_46554);
and UO_2995 (O_2995,N_47169,N_47526);
xor UO_2996 (O_2996,N_47194,N_48127);
or UO_2997 (O_2997,N_45941,N_49958);
xnor UO_2998 (O_2998,N_49127,N_47469);
nor UO_2999 (O_2999,N_45423,N_45221);
or UO_3000 (O_3000,N_45131,N_47669);
nand UO_3001 (O_3001,N_47716,N_45642);
nand UO_3002 (O_3002,N_46776,N_47307);
nand UO_3003 (O_3003,N_45907,N_48720);
nand UO_3004 (O_3004,N_46654,N_45540);
and UO_3005 (O_3005,N_47402,N_46817);
nor UO_3006 (O_3006,N_45982,N_48644);
or UO_3007 (O_3007,N_47506,N_48342);
and UO_3008 (O_3008,N_47273,N_45621);
nand UO_3009 (O_3009,N_46275,N_49440);
nand UO_3010 (O_3010,N_45751,N_47251);
and UO_3011 (O_3011,N_49275,N_49415);
xnor UO_3012 (O_3012,N_48934,N_48860);
nand UO_3013 (O_3013,N_47764,N_49116);
nand UO_3014 (O_3014,N_46766,N_48970);
and UO_3015 (O_3015,N_47995,N_46068);
xnor UO_3016 (O_3016,N_45871,N_45272);
nor UO_3017 (O_3017,N_49097,N_46668);
or UO_3018 (O_3018,N_47808,N_48591);
nand UO_3019 (O_3019,N_46933,N_49721);
nand UO_3020 (O_3020,N_45250,N_49143);
and UO_3021 (O_3021,N_49153,N_47735);
nor UO_3022 (O_3022,N_48652,N_48758);
or UO_3023 (O_3023,N_48412,N_47557);
or UO_3024 (O_3024,N_49507,N_46003);
xnor UO_3025 (O_3025,N_47630,N_48205);
or UO_3026 (O_3026,N_47379,N_48130);
xnor UO_3027 (O_3027,N_48187,N_48683);
xnor UO_3028 (O_3028,N_48136,N_49090);
and UO_3029 (O_3029,N_48665,N_45290);
xor UO_3030 (O_3030,N_47897,N_46395);
nor UO_3031 (O_3031,N_48811,N_48117);
nor UO_3032 (O_3032,N_47900,N_45763);
xor UO_3033 (O_3033,N_47874,N_48149);
nand UO_3034 (O_3034,N_46624,N_47801);
and UO_3035 (O_3035,N_49138,N_46887);
nor UO_3036 (O_3036,N_47822,N_48505);
nand UO_3037 (O_3037,N_46172,N_48762);
xnor UO_3038 (O_3038,N_46488,N_49128);
nand UO_3039 (O_3039,N_45326,N_47211);
or UO_3040 (O_3040,N_45807,N_49694);
and UO_3041 (O_3041,N_46076,N_48091);
nand UO_3042 (O_3042,N_46773,N_48706);
nand UO_3043 (O_3043,N_45472,N_49311);
or UO_3044 (O_3044,N_45552,N_46778);
nand UO_3045 (O_3045,N_49093,N_48189);
xor UO_3046 (O_3046,N_49967,N_47883);
nand UO_3047 (O_3047,N_45363,N_48178);
xnor UO_3048 (O_3048,N_47069,N_47828);
nor UO_3049 (O_3049,N_48668,N_49630);
and UO_3050 (O_3050,N_46713,N_48527);
or UO_3051 (O_3051,N_45522,N_47827);
or UO_3052 (O_3052,N_49693,N_46367);
xnor UO_3053 (O_3053,N_48396,N_48263);
nand UO_3054 (O_3054,N_46221,N_47787);
or UO_3055 (O_3055,N_46413,N_47392);
xor UO_3056 (O_3056,N_46653,N_47371);
nor UO_3057 (O_3057,N_48239,N_48735);
or UO_3058 (O_3058,N_46375,N_47567);
xnor UO_3059 (O_3059,N_47108,N_49489);
nor UO_3060 (O_3060,N_48958,N_47835);
nor UO_3061 (O_3061,N_47891,N_45019);
nor UO_3062 (O_3062,N_49725,N_45608);
xor UO_3063 (O_3063,N_47800,N_49898);
or UO_3064 (O_3064,N_49933,N_47425);
xnor UO_3065 (O_3065,N_46471,N_46211);
nand UO_3066 (O_3066,N_49601,N_47038);
xor UO_3067 (O_3067,N_49190,N_49743);
and UO_3068 (O_3068,N_49542,N_46618);
nor UO_3069 (O_3069,N_48028,N_48376);
nor UO_3070 (O_3070,N_46038,N_49120);
nor UO_3071 (O_3071,N_49441,N_47640);
or UO_3072 (O_3072,N_49273,N_45992);
xnor UO_3073 (O_3073,N_47140,N_49480);
xnor UO_3074 (O_3074,N_45730,N_48679);
nand UO_3075 (O_3075,N_45867,N_47242);
and UO_3076 (O_3076,N_49593,N_46489);
nor UO_3077 (O_3077,N_45436,N_47641);
or UO_3078 (O_3078,N_46135,N_48920);
or UO_3079 (O_3079,N_46534,N_49241);
or UO_3080 (O_3080,N_46072,N_46713);
and UO_3081 (O_3081,N_45963,N_49790);
nor UO_3082 (O_3082,N_46228,N_46316);
nand UO_3083 (O_3083,N_46171,N_45846);
or UO_3084 (O_3084,N_49284,N_45990);
or UO_3085 (O_3085,N_46849,N_47248);
xnor UO_3086 (O_3086,N_49408,N_48923);
nor UO_3087 (O_3087,N_47964,N_46067);
and UO_3088 (O_3088,N_48191,N_45603);
and UO_3089 (O_3089,N_46849,N_45355);
nand UO_3090 (O_3090,N_45498,N_46475);
nor UO_3091 (O_3091,N_46330,N_49467);
and UO_3092 (O_3092,N_48223,N_47122);
nand UO_3093 (O_3093,N_48858,N_45252);
nand UO_3094 (O_3094,N_45417,N_46145);
nand UO_3095 (O_3095,N_46426,N_47436);
xor UO_3096 (O_3096,N_45890,N_48930);
nor UO_3097 (O_3097,N_47785,N_47014);
or UO_3098 (O_3098,N_49140,N_49680);
nand UO_3099 (O_3099,N_49617,N_45067);
nand UO_3100 (O_3100,N_46382,N_48172);
xor UO_3101 (O_3101,N_49007,N_49124);
nor UO_3102 (O_3102,N_45913,N_48259);
nor UO_3103 (O_3103,N_48855,N_48105);
nand UO_3104 (O_3104,N_45658,N_46237);
xnor UO_3105 (O_3105,N_48917,N_46255);
xor UO_3106 (O_3106,N_47272,N_46869);
and UO_3107 (O_3107,N_48375,N_46837);
nor UO_3108 (O_3108,N_49275,N_46268);
nand UO_3109 (O_3109,N_49798,N_46741);
or UO_3110 (O_3110,N_47378,N_46694);
or UO_3111 (O_3111,N_49762,N_49441);
nand UO_3112 (O_3112,N_49300,N_46450);
or UO_3113 (O_3113,N_48699,N_45821);
xnor UO_3114 (O_3114,N_47949,N_46076);
nand UO_3115 (O_3115,N_49863,N_47564);
nor UO_3116 (O_3116,N_47876,N_48697);
nor UO_3117 (O_3117,N_48875,N_46977);
and UO_3118 (O_3118,N_49664,N_46854);
nand UO_3119 (O_3119,N_49730,N_48210);
xnor UO_3120 (O_3120,N_46996,N_49283);
nor UO_3121 (O_3121,N_45404,N_46067);
and UO_3122 (O_3122,N_47379,N_49709);
nor UO_3123 (O_3123,N_45759,N_48022);
and UO_3124 (O_3124,N_47781,N_48890);
or UO_3125 (O_3125,N_45304,N_45267);
and UO_3126 (O_3126,N_45443,N_49426);
xnor UO_3127 (O_3127,N_47020,N_49750);
or UO_3128 (O_3128,N_49413,N_45000);
nor UO_3129 (O_3129,N_47348,N_45233);
nor UO_3130 (O_3130,N_46507,N_45732);
nor UO_3131 (O_3131,N_48471,N_46786);
nor UO_3132 (O_3132,N_45413,N_46507);
nor UO_3133 (O_3133,N_45632,N_46488);
and UO_3134 (O_3134,N_48070,N_47784);
or UO_3135 (O_3135,N_46311,N_48602);
xor UO_3136 (O_3136,N_47256,N_47797);
nor UO_3137 (O_3137,N_49849,N_49950);
and UO_3138 (O_3138,N_45241,N_45060);
nand UO_3139 (O_3139,N_46848,N_45412);
nand UO_3140 (O_3140,N_49349,N_49060);
and UO_3141 (O_3141,N_47080,N_49597);
xnor UO_3142 (O_3142,N_48853,N_45453);
and UO_3143 (O_3143,N_47410,N_48512);
nand UO_3144 (O_3144,N_46286,N_48966);
nand UO_3145 (O_3145,N_49468,N_47873);
nand UO_3146 (O_3146,N_46277,N_47984);
xnor UO_3147 (O_3147,N_47584,N_46399);
xor UO_3148 (O_3148,N_49087,N_48621);
nor UO_3149 (O_3149,N_49349,N_46123);
xor UO_3150 (O_3150,N_47018,N_45610);
or UO_3151 (O_3151,N_49043,N_45702);
nand UO_3152 (O_3152,N_45297,N_48777);
or UO_3153 (O_3153,N_48239,N_45865);
nor UO_3154 (O_3154,N_47163,N_49280);
or UO_3155 (O_3155,N_45750,N_45028);
and UO_3156 (O_3156,N_49466,N_49150);
or UO_3157 (O_3157,N_48346,N_48204);
or UO_3158 (O_3158,N_47843,N_46044);
nor UO_3159 (O_3159,N_48043,N_47456);
and UO_3160 (O_3160,N_46307,N_45620);
nor UO_3161 (O_3161,N_46626,N_47154);
nand UO_3162 (O_3162,N_47104,N_45578);
nor UO_3163 (O_3163,N_49948,N_49527);
nor UO_3164 (O_3164,N_45351,N_47749);
nand UO_3165 (O_3165,N_47597,N_45053);
nand UO_3166 (O_3166,N_46183,N_48543);
nand UO_3167 (O_3167,N_48685,N_48631);
or UO_3168 (O_3168,N_46178,N_47635);
and UO_3169 (O_3169,N_46609,N_45723);
xnor UO_3170 (O_3170,N_49576,N_49899);
nand UO_3171 (O_3171,N_47950,N_45630);
nand UO_3172 (O_3172,N_47607,N_47115);
or UO_3173 (O_3173,N_46467,N_46253);
or UO_3174 (O_3174,N_49672,N_48578);
and UO_3175 (O_3175,N_48944,N_47053);
nor UO_3176 (O_3176,N_48537,N_45181);
or UO_3177 (O_3177,N_47371,N_46007);
or UO_3178 (O_3178,N_49281,N_45742);
nor UO_3179 (O_3179,N_49010,N_48778);
xnor UO_3180 (O_3180,N_46259,N_47157);
nor UO_3181 (O_3181,N_49706,N_48619);
xor UO_3182 (O_3182,N_48134,N_47472);
or UO_3183 (O_3183,N_46842,N_46801);
nand UO_3184 (O_3184,N_47040,N_47278);
xor UO_3185 (O_3185,N_45148,N_46756);
or UO_3186 (O_3186,N_47514,N_48950);
nor UO_3187 (O_3187,N_47067,N_45682);
nor UO_3188 (O_3188,N_46031,N_49575);
and UO_3189 (O_3189,N_45072,N_46997);
and UO_3190 (O_3190,N_45386,N_48613);
or UO_3191 (O_3191,N_47793,N_48147);
or UO_3192 (O_3192,N_46936,N_46975);
and UO_3193 (O_3193,N_45208,N_48266);
nor UO_3194 (O_3194,N_46457,N_48592);
and UO_3195 (O_3195,N_47287,N_47681);
or UO_3196 (O_3196,N_48257,N_45228);
nand UO_3197 (O_3197,N_49132,N_45883);
or UO_3198 (O_3198,N_48859,N_48408);
xor UO_3199 (O_3199,N_48267,N_49598);
or UO_3200 (O_3200,N_46269,N_47642);
or UO_3201 (O_3201,N_49869,N_48368);
or UO_3202 (O_3202,N_45195,N_49051);
and UO_3203 (O_3203,N_47917,N_46100);
xor UO_3204 (O_3204,N_46501,N_46844);
nor UO_3205 (O_3205,N_45109,N_48706);
nor UO_3206 (O_3206,N_47870,N_47595);
nand UO_3207 (O_3207,N_46211,N_47621);
and UO_3208 (O_3208,N_49212,N_48179);
or UO_3209 (O_3209,N_47976,N_49777);
and UO_3210 (O_3210,N_45516,N_46264);
or UO_3211 (O_3211,N_48932,N_48097);
nor UO_3212 (O_3212,N_47741,N_46611);
and UO_3213 (O_3213,N_47397,N_46642);
or UO_3214 (O_3214,N_47243,N_46460);
nand UO_3215 (O_3215,N_49072,N_47700);
nand UO_3216 (O_3216,N_46148,N_45862);
or UO_3217 (O_3217,N_49374,N_47890);
and UO_3218 (O_3218,N_46552,N_49637);
and UO_3219 (O_3219,N_49559,N_48150);
nand UO_3220 (O_3220,N_46689,N_48819);
nor UO_3221 (O_3221,N_45538,N_47830);
or UO_3222 (O_3222,N_49913,N_49313);
and UO_3223 (O_3223,N_47376,N_49155);
and UO_3224 (O_3224,N_48857,N_46526);
nand UO_3225 (O_3225,N_48909,N_48064);
nor UO_3226 (O_3226,N_47983,N_46137);
and UO_3227 (O_3227,N_49323,N_48248);
and UO_3228 (O_3228,N_46609,N_45941);
nand UO_3229 (O_3229,N_46352,N_49319);
and UO_3230 (O_3230,N_47719,N_45912);
nor UO_3231 (O_3231,N_46330,N_47611);
nand UO_3232 (O_3232,N_45772,N_45571);
nand UO_3233 (O_3233,N_46555,N_48655);
nand UO_3234 (O_3234,N_49725,N_47138);
nand UO_3235 (O_3235,N_45820,N_45221);
xnor UO_3236 (O_3236,N_45490,N_47197);
or UO_3237 (O_3237,N_46694,N_45051);
xnor UO_3238 (O_3238,N_46871,N_47302);
nand UO_3239 (O_3239,N_46596,N_49925);
nand UO_3240 (O_3240,N_46464,N_47976);
nor UO_3241 (O_3241,N_49503,N_48926);
nor UO_3242 (O_3242,N_48072,N_47735);
and UO_3243 (O_3243,N_46804,N_48296);
nand UO_3244 (O_3244,N_49982,N_49113);
xnor UO_3245 (O_3245,N_47336,N_47827);
xor UO_3246 (O_3246,N_46553,N_46875);
nand UO_3247 (O_3247,N_46190,N_47293);
nand UO_3248 (O_3248,N_49040,N_48959);
and UO_3249 (O_3249,N_46525,N_49551);
nand UO_3250 (O_3250,N_48364,N_45157);
xor UO_3251 (O_3251,N_47693,N_48452);
or UO_3252 (O_3252,N_45017,N_46363);
and UO_3253 (O_3253,N_47648,N_46510);
nand UO_3254 (O_3254,N_45636,N_49306);
xnor UO_3255 (O_3255,N_46149,N_46039);
and UO_3256 (O_3256,N_48306,N_45289);
nor UO_3257 (O_3257,N_45163,N_48444);
nand UO_3258 (O_3258,N_46896,N_48968);
xnor UO_3259 (O_3259,N_49944,N_45037);
and UO_3260 (O_3260,N_48269,N_45306);
or UO_3261 (O_3261,N_45456,N_45219);
xor UO_3262 (O_3262,N_49949,N_46465);
and UO_3263 (O_3263,N_47455,N_48692);
nand UO_3264 (O_3264,N_45683,N_46502);
and UO_3265 (O_3265,N_45675,N_47659);
or UO_3266 (O_3266,N_46271,N_49422);
nand UO_3267 (O_3267,N_46496,N_48406);
nand UO_3268 (O_3268,N_45531,N_45199);
nand UO_3269 (O_3269,N_46286,N_47576);
or UO_3270 (O_3270,N_47030,N_45545);
and UO_3271 (O_3271,N_46857,N_45071);
or UO_3272 (O_3272,N_47689,N_48917);
or UO_3273 (O_3273,N_45163,N_47371);
and UO_3274 (O_3274,N_46621,N_49365);
nor UO_3275 (O_3275,N_46509,N_47771);
nand UO_3276 (O_3276,N_48340,N_49497);
nor UO_3277 (O_3277,N_46353,N_45864);
nand UO_3278 (O_3278,N_48985,N_46671);
or UO_3279 (O_3279,N_48214,N_47371);
nor UO_3280 (O_3280,N_48004,N_47815);
nor UO_3281 (O_3281,N_45166,N_45426);
or UO_3282 (O_3282,N_47430,N_45425);
nor UO_3283 (O_3283,N_47374,N_48749);
xnor UO_3284 (O_3284,N_48775,N_49006);
nand UO_3285 (O_3285,N_47480,N_46659);
nor UO_3286 (O_3286,N_45380,N_47277);
or UO_3287 (O_3287,N_47413,N_46559);
nand UO_3288 (O_3288,N_47251,N_45487);
or UO_3289 (O_3289,N_47664,N_47331);
xnor UO_3290 (O_3290,N_46945,N_49215);
and UO_3291 (O_3291,N_49621,N_46168);
xor UO_3292 (O_3292,N_45878,N_45246);
and UO_3293 (O_3293,N_47293,N_45610);
xnor UO_3294 (O_3294,N_47746,N_48472);
xnor UO_3295 (O_3295,N_49110,N_45058);
xor UO_3296 (O_3296,N_46331,N_46360);
nand UO_3297 (O_3297,N_45807,N_45742);
nor UO_3298 (O_3298,N_46626,N_45864);
xor UO_3299 (O_3299,N_47805,N_49671);
or UO_3300 (O_3300,N_46081,N_47634);
nand UO_3301 (O_3301,N_49935,N_45815);
xor UO_3302 (O_3302,N_48904,N_47724);
or UO_3303 (O_3303,N_45586,N_49355);
nor UO_3304 (O_3304,N_46986,N_49979);
nor UO_3305 (O_3305,N_47654,N_48452);
nand UO_3306 (O_3306,N_47120,N_45809);
and UO_3307 (O_3307,N_49282,N_46746);
nor UO_3308 (O_3308,N_47710,N_47919);
and UO_3309 (O_3309,N_45689,N_46208);
or UO_3310 (O_3310,N_48266,N_47764);
xor UO_3311 (O_3311,N_46336,N_47313);
nor UO_3312 (O_3312,N_47990,N_45859);
and UO_3313 (O_3313,N_47738,N_48302);
and UO_3314 (O_3314,N_49675,N_45926);
or UO_3315 (O_3315,N_48494,N_47342);
or UO_3316 (O_3316,N_49453,N_45216);
nor UO_3317 (O_3317,N_45908,N_47686);
nand UO_3318 (O_3318,N_48334,N_48931);
nor UO_3319 (O_3319,N_49946,N_47346);
nand UO_3320 (O_3320,N_45925,N_48494);
or UO_3321 (O_3321,N_46515,N_47952);
nand UO_3322 (O_3322,N_46295,N_48151);
and UO_3323 (O_3323,N_46654,N_46588);
nor UO_3324 (O_3324,N_49539,N_48652);
nor UO_3325 (O_3325,N_47618,N_46723);
nor UO_3326 (O_3326,N_47020,N_46176);
nand UO_3327 (O_3327,N_46165,N_49909);
xor UO_3328 (O_3328,N_46042,N_49815);
or UO_3329 (O_3329,N_48896,N_48957);
xnor UO_3330 (O_3330,N_46018,N_46929);
xnor UO_3331 (O_3331,N_48525,N_49795);
nand UO_3332 (O_3332,N_49906,N_48448);
or UO_3333 (O_3333,N_45284,N_46206);
nand UO_3334 (O_3334,N_46713,N_49883);
xor UO_3335 (O_3335,N_47102,N_45706);
and UO_3336 (O_3336,N_46674,N_47670);
nand UO_3337 (O_3337,N_46812,N_47427);
and UO_3338 (O_3338,N_49342,N_49100);
and UO_3339 (O_3339,N_47008,N_46437);
xor UO_3340 (O_3340,N_49687,N_49328);
or UO_3341 (O_3341,N_49543,N_47244);
or UO_3342 (O_3342,N_46356,N_46705);
and UO_3343 (O_3343,N_48390,N_47637);
xnor UO_3344 (O_3344,N_48025,N_48593);
and UO_3345 (O_3345,N_48160,N_45088);
or UO_3346 (O_3346,N_45521,N_48587);
or UO_3347 (O_3347,N_45621,N_47331);
or UO_3348 (O_3348,N_45589,N_46180);
and UO_3349 (O_3349,N_49906,N_47467);
nor UO_3350 (O_3350,N_49893,N_45078);
xor UO_3351 (O_3351,N_47294,N_46441);
and UO_3352 (O_3352,N_45009,N_45386);
xnor UO_3353 (O_3353,N_46067,N_47267);
and UO_3354 (O_3354,N_46666,N_46073);
nand UO_3355 (O_3355,N_49705,N_48299);
nand UO_3356 (O_3356,N_46082,N_46215);
nand UO_3357 (O_3357,N_45874,N_46580);
and UO_3358 (O_3358,N_47350,N_45227);
xnor UO_3359 (O_3359,N_49394,N_48607);
or UO_3360 (O_3360,N_47475,N_45812);
and UO_3361 (O_3361,N_47054,N_48523);
and UO_3362 (O_3362,N_46520,N_47550);
and UO_3363 (O_3363,N_45784,N_47728);
xor UO_3364 (O_3364,N_46900,N_45290);
nor UO_3365 (O_3365,N_48154,N_46660);
xor UO_3366 (O_3366,N_47835,N_49735);
or UO_3367 (O_3367,N_48233,N_45149);
nor UO_3368 (O_3368,N_46405,N_45062);
xor UO_3369 (O_3369,N_46961,N_45058);
xnor UO_3370 (O_3370,N_48027,N_45080);
nor UO_3371 (O_3371,N_49825,N_47683);
nand UO_3372 (O_3372,N_48211,N_49260);
xnor UO_3373 (O_3373,N_47522,N_47669);
xor UO_3374 (O_3374,N_48938,N_46682);
xnor UO_3375 (O_3375,N_49604,N_45768);
or UO_3376 (O_3376,N_48632,N_48473);
or UO_3377 (O_3377,N_49369,N_49641);
nand UO_3378 (O_3378,N_49243,N_45949);
nand UO_3379 (O_3379,N_48475,N_47744);
or UO_3380 (O_3380,N_49975,N_46030);
nand UO_3381 (O_3381,N_45305,N_48536);
nand UO_3382 (O_3382,N_45639,N_47553);
xnor UO_3383 (O_3383,N_49919,N_48053);
and UO_3384 (O_3384,N_45494,N_47976);
xor UO_3385 (O_3385,N_46236,N_47987);
and UO_3386 (O_3386,N_48096,N_46029);
nand UO_3387 (O_3387,N_46162,N_45054);
nor UO_3388 (O_3388,N_47470,N_45905);
xnor UO_3389 (O_3389,N_49098,N_49929);
nand UO_3390 (O_3390,N_45662,N_49267);
nor UO_3391 (O_3391,N_48470,N_49361);
nor UO_3392 (O_3392,N_45387,N_49024);
and UO_3393 (O_3393,N_47848,N_46011);
nand UO_3394 (O_3394,N_45482,N_49144);
and UO_3395 (O_3395,N_49210,N_46821);
or UO_3396 (O_3396,N_45256,N_49412);
xnor UO_3397 (O_3397,N_45061,N_49247);
and UO_3398 (O_3398,N_47720,N_45131);
nor UO_3399 (O_3399,N_46855,N_45126);
or UO_3400 (O_3400,N_47860,N_45318);
and UO_3401 (O_3401,N_48538,N_48169);
nand UO_3402 (O_3402,N_49790,N_49105);
and UO_3403 (O_3403,N_47972,N_48033);
and UO_3404 (O_3404,N_45062,N_48245);
nor UO_3405 (O_3405,N_48235,N_49967);
nor UO_3406 (O_3406,N_45371,N_45818);
and UO_3407 (O_3407,N_46194,N_49058);
xnor UO_3408 (O_3408,N_47924,N_46218);
nor UO_3409 (O_3409,N_45128,N_49955);
or UO_3410 (O_3410,N_45457,N_47818);
and UO_3411 (O_3411,N_48285,N_46144);
xnor UO_3412 (O_3412,N_47297,N_47537);
nor UO_3413 (O_3413,N_47797,N_47810);
nor UO_3414 (O_3414,N_45678,N_48049);
or UO_3415 (O_3415,N_48475,N_45942);
xnor UO_3416 (O_3416,N_46410,N_46239);
and UO_3417 (O_3417,N_48175,N_48299);
nor UO_3418 (O_3418,N_45139,N_48830);
and UO_3419 (O_3419,N_46736,N_49668);
xor UO_3420 (O_3420,N_48276,N_46313);
nor UO_3421 (O_3421,N_47102,N_47930);
xor UO_3422 (O_3422,N_45732,N_48429);
or UO_3423 (O_3423,N_48779,N_48928);
or UO_3424 (O_3424,N_45442,N_48602);
or UO_3425 (O_3425,N_49554,N_49959);
xor UO_3426 (O_3426,N_46053,N_45757);
nor UO_3427 (O_3427,N_49472,N_45472);
and UO_3428 (O_3428,N_47926,N_45588);
and UO_3429 (O_3429,N_47187,N_49442);
nor UO_3430 (O_3430,N_48131,N_49407);
xnor UO_3431 (O_3431,N_46536,N_48523);
nor UO_3432 (O_3432,N_46278,N_49451);
nor UO_3433 (O_3433,N_45139,N_46321);
or UO_3434 (O_3434,N_49377,N_46803);
or UO_3435 (O_3435,N_49569,N_47333);
nand UO_3436 (O_3436,N_47368,N_46794);
and UO_3437 (O_3437,N_49515,N_45934);
nand UO_3438 (O_3438,N_48790,N_47508);
nor UO_3439 (O_3439,N_46330,N_46307);
or UO_3440 (O_3440,N_45737,N_46017);
and UO_3441 (O_3441,N_47677,N_47482);
and UO_3442 (O_3442,N_47325,N_49915);
xnor UO_3443 (O_3443,N_45634,N_47060);
xnor UO_3444 (O_3444,N_49955,N_46330);
or UO_3445 (O_3445,N_48230,N_47844);
xor UO_3446 (O_3446,N_47811,N_46704);
or UO_3447 (O_3447,N_45823,N_46215);
and UO_3448 (O_3448,N_46513,N_45331);
nand UO_3449 (O_3449,N_49863,N_49302);
nor UO_3450 (O_3450,N_46043,N_49336);
or UO_3451 (O_3451,N_47742,N_48143);
or UO_3452 (O_3452,N_45903,N_46514);
nand UO_3453 (O_3453,N_49936,N_46478);
nand UO_3454 (O_3454,N_45401,N_49587);
and UO_3455 (O_3455,N_48575,N_47448);
and UO_3456 (O_3456,N_49815,N_49481);
and UO_3457 (O_3457,N_48662,N_49966);
and UO_3458 (O_3458,N_48079,N_46409);
or UO_3459 (O_3459,N_47074,N_45823);
and UO_3460 (O_3460,N_45463,N_49583);
or UO_3461 (O_3461,N_47201,N_45062);
xor UO_3462 (O_3462,N_45282,N_45147);
xnor UO_3463 (O_3463,N_47848,N_49653);
or UO_3464 (O_3464,N_46428,N_49741);
nand UO_3465 (O_3465,N_47811,N_45598);
and UO_3466 (O_3466,N_47456,N_45170);
and UO_3467 (O_3467,N_49802,N_46224);
and UO_3468 (O_3468,N_48271,N_49134);
nand UO_3469 (O_3469,N_49570,N_46649);
nor UO_3470 (O_3470,N_47809,N_47396);
or UO_3471 (O_3471,N_49984,N_48534);
nor UO_3472 (O_3472,N_49718,N_49222);
or UO_3473 (O_3473,N_48639,N_47458);
or UO_3474 (O_3474,N_47154,N_49087);
nor UO_3475 (O_3475,N_49236,N_48527);
nand UO_3476 (O_3476,N_45809,N_47713);
nand UO_3477 (O_3477,N_46637,N_46479);
nand UO_3478 (O_3478,N_46278,N_47633);
or UO_3479 (O_3479,N_48916,N_45953);
and UO_3480 (O_3480,N_46431,N_48626);
nor UO_3481 (O_3481,N_45491,N_49837);
nor UO_3482 (O_3482,N_47006,N_45374);
or UO_3483 (O_3483,N_46345,N_48481);
and UO_3484 (O_3484,N_46204,N_48248);
and UO_3485 (O_3485,N_49513,N_49599);
nand UO_3486 (O_3486,N_48783,N_49566);
and UO_3487 (O_3487,N_47404,N_48496);
nor UO_3488 (O_3488,N_45692,N_45000);
and UO_3489 (O_3489,N_47660,N_48975);
or UO_3490 (O_3490,N_49501,N_48117);
and UO_3491 (O_3491,N_49728,N_49168);
and UO_3492 (O_3492,N_47278,N_45227);
or UO_3493 (O_3493,N_47569,N_46049);
xor UO_3494 (O_3494,N_46679,N_46218);
or UO_3495 (O_3495,N_45752,N_47449);
nand UO_3496 (O_3496,N_49943,N_48460);
and UO_3497 (O_3497,N_49828,N_49429);
nor UO_3498 (O_3498,N_45651,N_45225);
or UO_3499 (O_3499,N_47532,N_46074);
or UO_3500 (O_3500,N_49767,N_48253);
nor UO_3501 (O_3501,N_46750,N_49629);
xnor UO_3502 (O_3502,N_46629,N_49312);
xnor UO_3503 (O_3503,N_48111,N_46447);
xnor UO_3504 (O_3504,N_45586,N_45396);
nand UO_3505 (O_3505,N_45421,N_45742);
xnor UO_3506 (O_3506,N_49553,N_49847);
nor UO_3507 (O_3507,N_48291,N_47154);
or UO_3508 (O_3508,N_49024,N_47368);
xnor UO_3509 (O_3509,N_46838,N_48347);
and UO_3510 (O_3510,N_45775,N_49116);
nor UO_3511 (O_3511,N_45683,N_48933);
nand UO_3512 (O_3512,N_48745,N_45930);
or UO_3513 (O_3513,N_45376,N_46331);
nand UO_3514 (O_3514,N_49319,N_48736);
nand UO_3515 (O_3515,N_45827,N_46924);
xnor UO_3516 (O_3516,N_49342,N_49379);
or UO_3517 (O_3517,N_47091,N_46126);
nand UO_3518 (O_3518,N_47297,N_49916);
nor UO_3519 (O_3519,N_49769,N_48886);
and UO_3520 (O_3520,N_49180,N_49541);
and UO_3521 (O_3521,N_47790,N_48564);
and UO_3522 (O_3522,N_49608,N_47738);
and UO_3523 (O_3523,N_45226,N_46075);
xnor UO_3524 (O_3524,N_48920,N_49021);
or UO_3525 (O_3525,N_49985,N_45324);
and UO_3526 (O_3526,N_45019,N_47185);
xnor UO_3527 (O_3527,N_47775,N_47011);
nor UO_3528 (O_3528,N_47165,N_47086);
nand UO_3529 (O_3529,N_49246,N_47526);
nand UO_3530 (O_3530,N_45177,N_48957);
nor UO_3531 (O_3531,N_46493,N_48808);
and UO_3532 (O_3532,N_47340,N_49875);
nand UO_3533 (O_3533,N_47304,N_49987);
nand UO_3534 (O_3534,N_49274,N_46164);
and UO_3535 (O_3535,N_49601,N_47625);
nand UO_3536 (O_3536,N_45892,N_48417);
xnor UO_3537 (O_3537,N_45267,N_47339);
nand UO_3538 (O_3538,N_45245,N_49709);
nor UO_3539 (O_3539,N_49544,N_49868);
nand UO_3540 (O_3540,N_46767,N_45080);
or UO_3541 (O_3541,N_48804,N_46038);
nor UO_3542 (O_3542,N_49511,N_48201);
xnor UO_3543 (O_3543,N_45882,N_47766);
nand UO_3544 (O_3544,N_49302,N_48671);
xnor UO_3545 (O_3545,N_48141,N_48348);
and UO_3546 (O_3546,N_47850,N_46219);
nand UO_3547 (O_3547,N_48985,N_49145);
nand UO_3548 (O_3548,N_49816,N_49518);
nor UO_3549 (O_3549,N_45691,N_45203);
nand UO_3550 (O_3550,N_49422,N_49493);
and UO_3551 (O_3551,N_46698,N_46549);
and UO_3552 (O_3552,N_45340,N_46449);
and UO_3553 (O_3553,N_45579,N_46355);
xor UO_3554 (O_3554,N_48948,N_49506);
nor UO_3555 (O_3555,N_45867,N_45159);
nand UO_3556 (O_3556,N_45173,N_45432);
nor UO_3557 (O_3557,N_49345,N_48936);
nor UO_3558 (O_3558,N_46625,N_49572);
xor UO_3559 (O_3559,N_48443,N_46516);
xnor UO_3560 (O_3560,N_47025,N_45198);
or UO_3561 (O_3561,N_48568,N_47888);
and UO_3562 (O_3562,N_45044,N_46035);
and UO_3563 (O_3563,N_47517,N_45143);
nor UO_3564 (O_3564,N_49223,N_47482);
or UO_3565 (O_3565,N_49117,N_48483);
or UO_3566 (O_3566,N_45369,N_46282);
nor UO_3567 (O_3567,N_49206,N_49613);
or UO_3568 (O_3568,N_49479,N_45128);
nand UO_3569 (O_3569,N_49055,N_47587);
nand UO_3570 (O_3570,N_45135,N_45669);
xnor UO_3571 (O_3571,N_49226,N_46392);
nor UO_3572 (O_3572,N_48604,N_45212);
or UO_3573 (O_3573,N_48328,N_48915);
and UO_3574 (O_3574,N_48634,N_45913);
nand UO_3575 (O_3575,N_45723,N_47996);
and UO_3576 (O_3576,N_49729,N_49492);
nand UO_3577 (O_3577,N_45428,N_48834);
and UO_3578 (O_3578,N_45384,N_48432);
or UO_3579 (O_3579,N_48222,N_49904);
nor UO_3580 (O_3580,N_49227,N_49607);
xnor UO_3581 (O_3581,N_49983,N_45570);
nand UO_3582 (O_3582,N_46716,N_48851);
nand UO_3583 (O_3583,N_49350,N_45425);
nand UO_3584 (O_3584,N_47521,N_48901);
nand UO_3585 (O_3585,N_47025,N_48170);
and UO_3586 (O_3586,N_45226,N_48861);
and UO_3587 (O_3587,N_46946,N_46450);
nor UO_3588 (O_3588,N_48091,N_48367);
xor UO_3589 (O_3589,N_48887,N_47621);
nand UO_3590 (O_3590,N_47559,N_48238);
and UO_3591 (O_3591,N_45474,N_48610);
xor UO_3592 (O_3592,N_48064,N_47674);
nand UO_3593 (O_3593,N_47873,N_46895);
xor UO_3594 (O_3594,N_47931,N_47373);
or UO_3595 (O_3595,N_46034,N_49498);
nor UO_3596 (O_3596,N_45354,N_48174);
xor UO_3597 (O_3597,N_47650,N_48228);
nor UO_3598 (O_3598,N_46307,N_46224);
xor UO_3599 (O_3599,N_48644,N_47609);
nor UO_3600 (O_3600,N_47786,N_48451);
nor UO_3601 (O_3601,N_45809,N_47742);
or UO_3602 (O_3602,N_47458,N_45383);
nor UO_3603 (O_3603,N_47741,N_49121);
and UO_3604 (O_3604,N_47226,N_45814);
nor UO_3605 (O_3605,N_49229,N_48540);
nand UO_3606 (O_3606,N_47618,N_45977);
nand UO_3607 (O_3607,N_45183,N_48344);
nor UO_3608 (O_3608,N_48642,N_47339);
nand UO_3609 (O_3609,N_46232,N_46749);
xnor UO_3610 (O_3610,N_47793,N_47135);
xor UO_3611 (O_3611,N_49870,N_46425);
nor UO_3612 (O_3612,N_49599,N_49085);
or UO_3613 (O_3613,N_49479,N_48296);
and UO_3614 (O_3614,N_49856,N_48669);
and UO_3615 (O_3615,N_48620,N_49930);
and UO_3616 (O_3616,N_48811,N_48992);
or UO_3617 (O_3617,N_49717,N_46278);
or UO_3618 (O_3618,N_47031,N_45422);
nand UO_3619 (O_3619,N_47004,N_49774);
and UO_3620 (O_3620,N_48258,N_45895);
or UO_3621 (O_3621,N_48038,N_48931);
nand UO_3622 (O_3622,N_47355,N_47060);
nor UO_3623 (O_3623,N_46042,N_46361);
or UO_3624 (O_3624,N_45126,N_45895);
nor UO_3625 (O_3625,N_46324,N_45268);
nand UO_3626 (O_3626,N_48646,N_48792);
and UO_3627 (O_3627,N_47455,N_48649);
or UO_3628 (O_3628,N_45721,N_45955);
and UO_3629 (O_3629,N_46702,N_47393);
xor UO_3630 (O_3630,N_46554,N_48219);
nor UO_3631 (O_3631,N_49564,N_47220);
and UO_3632 (O_3632,N_46346,N_48078);
nand UO_3633 (O_3633,N_45863,N_48034);
nand UO_3634 (O_3634,N_49523,N_47542);
or UO_3635 (O_3635,N_47099,N_45320);
xor UO_3636 (O_3636,N_45068,N_46863);
or UO_3637 (O_3637,N_48459,N_48975);
xnor UO_3638 (O_3638,N_45890,N_48771);
xor UO_3639 (O_3639,N_49401,N_49489);
and UO_3640 (O_3640,N_49268,N_46003);
nand UO_3641 (O_3641,N_45011,N_48535);
xor UO_3642 (O_3642,N_46611,N_45422);
or UO_3643 (O_3643,N_47142,N_49472);
nand UO_3644 (O_3644,N_47912,N_47647);
xnor UO_3645 (O_3645,N_46937,N_46115);
or UO_3646 (O_3646,N_45233,N_49486);
nand UO_3647 (O_3647,N_49781,N_48400);
nor UO_3648 (O_3648,N_49514,N_45263);
nor UO_3649 (O_3649,N_47542,N_45403);
or UO_3650 (O_3650,N_47527,N_45519);
xor UO_3651 (O_3651,N_49839,N_48714);
xnor UO_3652 (O_3652,N_46471,N_46851);
or UO_3653 (O_3653,N_45365,N_47287);
and UO_3654 (O_3654,N_45131,N_46798);
or UO_3655 (O_3655,N_46231,N_49099);
nand UO_3656 (O_3656,N_48453,N_45590);
xor UO_3657 (O_3657,N_46173,N_46736);
nor UO_3658 (O_3658,N_45727,N_48563);
and UO_3659 (O_3659,N_49223,N_46172);
xor UO_3660 (O_3660,N_46266,N_48172);
nor UO_3661 (O_3661,N_45410,N_46834);
xnor UO_3662 (O_3662,N_48490,N_47152);
and UO_3663 (O_3663,N_49624,N_49848);
nand UO_3664 (O_3664,N_48550,N_48956);
xor UO_3665 (O_3665,N_47836,N_46139);
nand UO_3666 (O_3666,N_46441,N_48409);
nand UO_3667 (O_3667,N_49604,N_46422);
xor UO_3668 (O_3668,N_45963,N_47825);
or UO_3669 (O_3669,N_48914,N_49736);
nor UO_3670 (O_3670,N_48161,N_48163);
xnor UO_3671 (O_3671,N_46040,N_48961);
and UO_3672 (O_3672,N_47587,N_49509);
and UO_3673 (O_3673,N_49956,N_46168);
nand UO_3674 (O_3674,N_47032,N_47128);
or UO_3675 (O_3675,N_46510,N_48594);
nand UO_3676 (O_3676,N_46807,N_49617);
nor UO_3677 (O_3677,N_49637,N_45245);
and UO_3678 (O_3678,N_46877,N_49289);
xor UO_3679 (O_3679,N_45571,N_46327);
nand UO_3680 (O_3680,N_45729,N_48723);
or UO_3681 (O_3681,N_45994,N_47930);
xor UO_3682 (O_3682,N_45111,N_46603);
and UO_3683 (O_3683,N_49469,N_48411);
nand UO_3684 (O_3684,N_47662,N_48394);
and UO_3685 (O_3685,N_48116,N_45473);
and UO_3686 (O_3686,N_48338,N_45199);
and UO_3687 (O_3687,N_46157,N_45900);
xor UO_3688 (O_3688,N_46945,N_49303);
nand UO_3689 (O_3689,N_47060,N_46104);
and UO_3690 (O_3690,N_45544,N_48426);
nor UO_3691 (O_3691,N_47447,N_46851);
and UO_3692 (O_3692,N_49763,N_49291);
or UO_3693 (O_3693,N_45748,N_49827);
nand UO_3694 (O_3694,N_47001,N_49336);
nor UO_3695 (O_3695,N_49591,N_45011);
xnor UO_3696 (O_3696,N_46472,N_46031);
and UO_3697 (O_3697,N_48052,N_49984);
xnor UO_3698 (O_3698,N_47108,N_47811);
nor UO_3699 (O_3699,N_49094,N_47081);
and UO_3700 (O_3700,N_46345,N_45823);
nor UO_3701 (O_3701,N_49777,N_48835);
or UO_3702 (O_3702,N_45698,N_47061);
nor UO_3703 (O_3703,N_47788,N_46936);
or UO_3704 (O_3704,N_47684,N_46179);
nand UO_3705 (O_3705,N_46605,N_46008);
or UO_3706 (O_3706,N_46871,N_47323);
or UO_3707 (O_3707,N_48413,N_46433);
nor UO_3708 (O_3708,N_45133,N_47963);
and UO_3709 (O_3709,N_49545,N_47494);
or UO_3710 (O_3710,N_48237,N_46843);
or UO_3711 (O_3711,N_47459,N_45042);
nor UO_3712 (O_3712,N_46945,N_47407);
nor UO_3713 (O_3713,N_47015,N_45631);
and UO_3714 (O_3714,N_47695,N_47832);
nor UO_3715 (O_3715,N_47903,N_45228);
nand UO_3716 (O_3716,N_49635,N_49640);
and UO_3717 (O_3717,N_48175,N_48657);
xnor UO_3718 (O_3718,N_45640,N_47695);
nand UO_3719 (O_3719,N_49137,N_45217);
nor UO_3720 (O_3720,N_46149,N_49130);
nor UO_3721 (O_3721,N_48092,N_48498);
nor UO_3722 (O_3722,N_49421,N_46612);
nor UO_3723 (O_3723,N_49986,N_47614);
xnor UO_3724 (O_3724,N_49190,N_47776);
and UO_3725 (O_3725,N_46680,N_47666);
nor UO_3726 (O_3726,N_47508,N_49155);
xnor UO_3727 (O_3727,N_48959,N_45800);
nand UO_3728 (O_3728,N_48950,N_47747);
or UO_3729 (O_3729,N_48887,N_45157);
nor UO_3730 (O_3730,N_45912,N_46443);
and UO_3731 (O_3731,N_45261,N_48574);
xor UO_3732 (O_3732,N_46637,N_48658);
and UO_3733 (O_3733,N_47798,N_47279);
or UO_3734 (O_3734,N_45470,N_45175);
and UO_3735 (O_3735,N_46573,N_45471);
xnor UO_3736 (O_3736,N_49931,N_48611);
nor UO_3737 (O_3737,N_46800,N_47623);
or UO_3738 (O_3738,N_47630,N_45586);
or UO_3739 (O_3739,N_45582,N_49423);
nand UO_3740 (O_3740,N_49552,N_46771);
and UO_3741 (O_3741,N_45886,N_46985);
or UO_3742 (O_3742,N_48611,N_48782);
nor UO_3743 (O_3743,N_47780,N_46294);
or UO_3744 (O_3744,N_48254,N_45724);
nand UO_3745 (O_3745,N_49635,N_49915);
nor UO_3746 (O_3746,N_48239,N_46548);
and UO_3747 (O_3747,N_47396,N_46510);
and UO_3748 (O_3748,N_46676,N_45762);
nor UO_3749 (O_3749,N_49853,N_47392);
or UO_3750 (O_3750,N_45444,N_47296);
and UO_3751 (O_3751,N_48056,N_49770);
and UO_3752 (O_3752,N_45676,N_45632);
xor UO_3753 (O_3753,N_47252,N_49897);
or UO_3754 (O_3754,N_45054,N_49211);
nor UO_3755 (O_3755,N_46327,N_48831);
xnor UO_3756 (O_3756,N_48801,N_45487);
nand UO_3757 (O_3757,N_45966,N_47923);
xor UO_3758 (O_3758,N_48928,N_46212);
or UO_3759 (O_3759,N_49313,N_48273);
or UO_3760 (O_3760,N_46135,N_45535);
nand UO_3761 (O_3761,N_48942,N_49877);
nand UO_3762 (O_3762,N_48468,N_48842);
or UO_3763 (O_3763,N_49177,N_48812);
nor UO_3764 (O_3764,N_47465,N_45688);
nand UO_3765 (O_3765,N_46257,N_48750);
xor UO_3766 (O_3766,N_48201,N_47721);
nand UO_3767 (O_3767,N_48989,N_49869);
nor UO_3768 (O_3768,N_46208,N_49875);
and UO_3769 (O_3769,N_49043,N_45950);
and UO_3770 (O_3770,N_48211,N_48849);
nand UO_3771 (O_3771,N_48546,N_46755);
xor UO_3772 (O_3772,N_48205,N_45644);
and UO_3773 (O_3773,N_47725,N_46746);
or UO_3774 (O_3774,N_46849,N_48167);
nor UO_3775 (O_3775,N_49346,N_47417);
nor UO_3776 (O_3776,N_49294,N_47519);
xnor UO_3777 (O_3777,N_47663,N_49634);
or UO_3778 (O_3778,N_46971,N_46547);
or UO_3779 (O_3779,N_48986,N_48424);
and UO_3780 (O_3780,N_46142,N_46141);
or UO_3781 (O_3781,N_45531,N_45366);
nor UO_3782 (O_3782,N_47957,N_48644);
or UO_3783 (O_3783,N_45414,N_48440);
nor UO_3784 (O_3784,N_46523,N_46093);
xor UO_3785 (O_3785,N_49199,N_49963);
and UO_3786 (O_3786,N_46132,N_47560);
nand UO_3787 (O_3787,N_45318,N_49943);
nor UO_3788 (O_3788,N_49909,N_45713);
and UO_3789 (O_3789,N_47872,N_46466);
nor UO_3790 (O_3790,N_46361,N_46545);
or UO_3791 (O_3791,N_47638,N_49787);
xnor UO_3792 (O_3792,N_48117,N_45887);
nor UO_3793 (O_3793,N_48489,N_45530);
or UO_3794 (O_3794,N_46369,N_45265);
or UO_3795 (O_3795,N_45935,N_46253);
and UO_3796 (O_3796,N_45170,N_47324);
or UO_3797 (O_3797,N_45694,N_45952);
and UO_3798 (O_3798,N_49643,N_48765);
or UO_3799 (O_3799,N_48625,N_49058);
or UO_3800 (O_3800,N_49006,N_46337);
and UO_3801 (O_3801,N_45764,N_48937);
nor UO_3802 (O_3802,N_47583,N_45326);
or UO_3803 (O_3803,N_48587,N_45056);
nor UO_3804 (O_3804,N_45170,N_45151);
xor UO_3805 (O_3805,N_47042,N_48781);
xnor UO_3806 (O_3806,N_48965,N_47140);
or UO_3807 (O_3807,N_48437,N_47825);
and UO_3808 (O_3808,N_47856,N_48892);
or UO_3809 (O_3809,N_48038,N_47457);
nand UO_3810 (O_3810,N_46503,N_46344);
or UO_3811 (O_3811,N_49503,N_45229);
xnor UO_3812 (O_3812,N_49985,N_46815);
xor UO_3813 (O_3813,N_46576,N_46284);
xnor UO_3814 (O_3814,N_49288,N_48578);
nand UO_3815 (O_3815,N_49311,N_47584);
nand UO_3816 (O_3816,N_47242,N_46167);
xor UO_3817 (O_3817,N_47576,N_47987);
or UO_3818 (O_3818,N_48813,N_48274);
xnor UO_3819 (O_3819,N_45304,N_45025);
or UO_3820 (O_3820,N_45655,N_48396);
and UO_3821 (O_3821,N_46545,N_45071);
xor UO_3822 (O_3822,N_47543,N_49622);
or UO_3823 (O_3823,N_48230,N_47464);
nor UO_3824 (O_3824,N_48380,N_46795);
xnor UO_3825 (O_3825,N_45005,N_47712);
or UO_3826 (O_3826,N_46922,N_49721);
and UO_3827 (O_3827,N_49427,N_47624);
nand UO_3828 (O_3828,N_45651,N_49853);
nor UO_3829 (O_3829,N_45283,N_47082);
xor UO_3830 (O_3830,N_45552,N_45747);
xor UO_3831 (O_3831,N_49566,N_49141);
nand UO_3832 (O_3832,N_49019,N_45608);
nand UO_3833 (O_3833,N_48700,N_46179);
and UO_3834 (O_3834,N_48640,N_45622);
nand UO_3835 (O_3835,N_48004,N_48466);
or UO_3836 (O_3836,N_49638,N_47241);
xor UO_3837 (O_3837,N_48935,N_48826);
or UO_3838 (O_3838,N_48675,N_46139);
nor UO_3839 (O_3839,N_48137,N_49911);
nor UO_3840 (O_3840,N_47888,N_47474);
and UO_3841 (O_3841,N_46887,N_48273);
nor UO_3842 (O_3842,N_46059,N_47205);
xor UO_3843 (O_3843,N_46291,N_49858);
or UO_3844 (O_3844,N_46314,N_48213);
nor UO_3845 (O_3845,N_48725,N_46469);
or UO_3846 (O_3846,N_47024,N_45306);
xor UO_3847 (O_3847,N_49808,N_47209);
and UO_3848 (O_3848,N_46051,N_46934);
and UO_3849 (O_3849,N_49672,N_49647);
xnor UO_3850 (O_3850,N_48135,N_45235);
nand UO_3851 (O_3851,N_47779,N_47768);
or UO_3852 (O_3852,N_47633,N_46838);
or UO_3853 (O_3853,N_49499,N_47745);
nand UO_3854 (O_3854,N_49085,N_48572);
and UO_3855 (O_3855,N_46328,N_48987);
nor UO_3856 (O_3856,N_48510,N_45783);
and UO_3857 (O_3857,N_46536,N_48246);
nor UO_3858 (O_3858,N_48608,N_47918);
and UO_3859 (O_3859,N_46651,N_48237);
xor UO_3860 (O_3860,N_47726,N_47221);
and UO_3861 (O_3861,N_48179,N_49802);
xor UO_3862 (O_3862,N_46516,N_47425);
nor UO_3863 (O_3863,N_46565,N_46288);
nor UO_3864 (O_3864,N_46346,N_48445);
and UO_3865 (O_3865,N_47982,N_46975);
and UO_3866 (O_3866,N_45832,N_46199);
nor UO_3867 (O_3867,N_45587,N_49929);
nand UO_3868 (O_3868,N_46680,N_46620);
nand UO_3869 (O_3869,N_48133,N_45408);
nand UO_3870 (O_3870,N_45317,N_45293);
xor UO_3871 (O_3871,N_48290,N_49163);
and UO_3872 (O_3872,N_46562,N_45954);
and UO_3873 (O_3873,N_47761,N_48449);
xor UO_3874 (O_3874,N_48405,N_47174);
or UO_3875 (O_3875,N_45435,N_45918);
or UO_3876 (O_3876,N_48169,N_48567);
nor UO_3877 (O_3877,N_46365,N_46011);
nor UO_3878 (O_3878,N_48254,N_49254);
nor UO_3879 (O_3879,N_47574,N_49224);
xor UO_3880 (O_3880,N_49679,N_46182);
nand UO_3881 (O_3881,N_48328,N_45988);
and UO_3882 (O_3882,N_48154,N_47745);
and UO_3883 (O_3883,N_47984,N_45094);
and UO_3884 (O_3884,N_46061,N_47080);
or UO_3885 (O_3885,N_47112,N_47641);
nand UO_3886 (O_3886,N_48285,N_46852);
and UO_3887 (O_3887,N_46008,N_48876);
nor UO_3888 (O_3888,N_45896,N_46965);
nand UO_3889 (O_3889,N_46703,N_48270);
nor UO_3890 (O_3890,N_46351,N_49309);
nand UO_3891 (O_3891,N_46539,N_45987);
xor UO_3892 (O_3892,N_49198,N_45350);
and UO_3893 (O_3893,N_47745,N_47482);
nor UO_3894 (O_3894,N_45757,N_48603);
or UO_3895 (O_3895,N_45285,N_48628);
or UO_3896 (O_3896,N_45098,N_45095);
or UO_3897 (O_3897,N_48410,N_46540);
xnor UO_3898 (O_3898,N_46465,N_47188);
or UO_3899 (O_3899,N_47367,N_49952);
and UO_3900 (O_3900,N_47830,N_49726);
and UO_3901 (O_3901,N_45903,N_46343);
nand UO_3902 (O_3902,N_49265,N_48118);
xor UO_3903 (O_3903,N_45367,N_45665);
or UO_3904 (O_3904,N_46075,N_47874);
nand UO_3905 (O_3905,N_49100,N_49822);
nand UO_3906 (O_3906,N_46440,N_48042);
and UO_3907 (O_3907,N_45014,N_46780);
and UO_3908 (O_3908,N_47531,N_46816);
nor UO_3909 (O_3909,N_48706,N_49608);
nand UO_3910 (O_3910,N_49002,N_48418);
xor UO_3911 (O_3911,N_47027,N_48026);
nand UO_3912 (O_3912,N_46932,N_49063);
nor UO_3913 (O_3913,N_48385,N_47068);
nor UO_3914 (O_3914,N_47030,N_46968);
nor UO_3915 (O_3915,N_46862,N_46443);
or UO_3916 (O_3916,N_47694,N_47102);
nand UO_3917 (O_3917,N_47274,N_48083);
nor UO_3918 (O_3918,N_47336,N_46428);
nor UO_3919 (O_3919,N_47024,N_45683);
or UO_3920 (O_3920,N_48255,N_46836);
xor UO_3921 (O_3921,N_48072,N_46614);
xnor UO_3922 (O_3922,N_46013,N_46162);
or UO_3923 (O_3923,N_45833,N_46606);
and UO_3924 (O_3924,N_49784,N_47214);
nor UO_3925 (O_3925,N_48470,N_48836);
and UO_3926 (O_3926,N_48891,N_48922);
and UO_3927 (O_3927,N_48194,N_48113);
nor UO_3928 (O_3928,N_49405,N_49144);
xnor UO_3929 (O_3929,N_48040,N_47415);
nand UO_3930 (O_3930,N_49309,N_48452);
or UO_3931 (O_3931,N_45737,N_49333);
and UO_3932 (O_3932,N_47198,N_47731);
nand UO_3933 (O_3933,N_49614,N_49394);
nor UO_3934 (O_3934,N_46132,N_49066);
nor UO_3935 (O_3935,N_47994,N_48180);
and UO_3936 (O_3936,N_49303,N_45847);
or UO_3937 (O_3937,N_45382,N_49026);
nand UO_3938 (O_3938,N_45893,N_48308);
and UO_3939 (O_3939,N_49827,N_49957);
and UO_3940 (O_3940,N_46531,N_46742);
xnor UO_3941 (O_3941,N_46219,N_48355);
and UO_3942 (O_3942,N_49372,N_48758);
nand UO_3943 (O_3943,N_46771,N_45956);
and UO_3944 (O_3944,N_48615,N_45090);
nand UO_3945 (O_3945,N_48701,N_45776);
xor UO_3946 (O_3946,N_48134,N_46017);
or UO_3947 (O_3947,N_49253,N_49801);
xnor UO_3948 (O_3948,N_48457,N_45813);
nand UO_3949 (O_3949,N_47456,N_48114);
nor UO_3950 (O_3950,N_47173,N_49354);
or UO_3951 (O_3951,N_49243,N_47545);
nand UO_3952 (O_3952,N_47701,N_48092);
xor UO_3953 (O_3953,N_49843,N_47190);
and UO_3954 (O_3954,N_49096,N_47272);
and UO_3955 (O_3955,N_49979,N_46522);
xor UO_3956 (O_3956,N_47709,N_45961);
nand UO_3957 (O_3957,N_47293,N_48174);
or UO_3958 (O_3958,N_47260,N_45577);
and UO_3959 (O_3959,N_45435,N_46586);
or UO_3960 (O_3960,N_47901,N_47163);
and UO_3961 (O_3961,N_46253,N_48197);
nor UO_3962 (O_3962,N_47494,N_48687);
nand UO_3963 (O_3963,N_46942,N_47239);
xor UO_3964 (O_3964,N_49648,N_49514);
xnor UO_3965 (O_3965,N_49324,N_47960);
or UO_3966 (O_3966,N_46268,N_49583);
xnor UO_3967 (O_3967,N_48108,N_46691);
nor UO_3968 (O_3968,N_49012,N_45077);
nor UO_3969 (O_3969,N_46455,N_45233);
and UO_3970 (O_3970,N_48332,N_45157);
and UO_3971 (O_3971,N_48279,N_46173);
nor UO_3972 (O_3972,N_46773,N_47526);
and UO_3973 (O_3973,N_45986,N_49007);
nand UO_3974 (O_3974,N_47825,N_47648);
or UO_3975 (O_3975,N_49715,N_46401);
nand UO_3976 (O_3976,N_47972,N_48160);
or UO_3977 (O_3977,N_48836,N_47545);
nor UO_3978 (O_3978,N_49706,N_49273);
xor UO_3979 (O_3979,N_47372,N_49421);
xnor UO_3980 (O_3980,N_48020,N_49107);
and UO_3981 (O_3981,N_47599,N_46768);
nor UO_3982 (O_3982,N_49973,N_48713);
nor UO_3983 (O_3983,N_48138,N_47131);
nand UO_3984 (O_3984,N_47338,N_46760);
xnor UO_3985 (O_3985,N_47508,N_48525);
nand UO_3986 (O_3986,N_49320,N_48367);
nand UO_3987 (O_3987,N_47280,N_47175);
nor UO_3988 (O_3988,N_47422,N_45016);
and UO_3989 (O_3989,N_48471,N_48563);
and UO_3990 (O_3990,N_49720,N_48006);
xnor UO_3991 (O_3991,N_48966,N_49195);
nor UO_3992 (O_3992,N_45651,N_48496);
xnor UO_3993 (O_3993,N_47296,N_47300);
and UO_3994 (O_3994,N_47086,N_49203);
nand UO_3995 (O_3995,N_45592,N_48146);
nand UO_3996 (O_3996,N_48978,N_45514);
and UO_3997 (O_3997,N_46101,N_45231);
xnor UO_3998 (O_3998,N_49689,N_47103);
or UO_3999 (O_3999,N_47653,N_48652);
and UO_4000 (O_4000,N_48652,N_45325);
nor UO_4001 (O_4001,N_48681,N_46477);
and UO_4002 (O_4002,N_46210,N_47034);
nor UO_4003 (O_4003,N_48510,N_48691);
or UO_4004 (O_4004,N_45676,N_49644);
xor UO_4005 (O_4005,N_45577,N_46311);
or UO_4006 (O_4006,N_48749,N_48689);
xor UO_4007 (O_4007,N_48841,N_45334);
nand UO_4008 (O_4008,N_45985,N_46683);
or UO_4009 (O_4009,N_46663,N_48745);
nor UO_4010 (O_4010,N_49676,N_46104);
nor UO_4011 (O_4011,N_47477,N_45075);
or UO_4012 (O_4012,N_47028,N_45613);
xor UO_4013 (O_4013,N_46057,N_48207);
nand UO_4014 (O_4014,N_47869,N_47249);
nand UO_4015 (O_4015,N_49451,N_48536);
and UO_4016 (O_4016,N_49027,N_45092);
xor UO_4017 (O_4017,N_49493,N_46328);
or UO_4018 (O_4018,N_48709,N_47042);
nor UO_4019 (O_4019,N_46244,N_47048);
nor UO_4020 (O_4020,N_46548,N_47545);
or UO_4021 (O_4021,N_45149,N_49623);
xor UO_4022 (O_4022,N_49611,N_46265);
nor UO_4023 (O_4023,N_45485,N_49686);
xor UO_4024 (O_4024,N_48477,N_49161);
and UO_4025 (O_4025,N_49312,N_48047);
nand UO_4026 (O_4026,N_49222,N_45501);
nand UO_4027 (O_4027,N_47106,N_48382);
nor UO_4028 (O_4028,N_47513,N_47715);
nand UO_4029 (O_4029,N_45369,N_49735);
xnor UO_4030 (O_4030,N_45372,N_46618);
xnor UO_4031 (O_4031,N_48469,N_49212);
and UO_4032 (O_4032,N_48116,N_45793);
and UO_4033 (O_4033,N_45484,N_45728);
xnor UO_4034 (O_4034,N_49139,N_48781);
nor UO_4035 (O_4035,N_47457,N_46989);
xnor UO_4036 (O_4036,N_49677,N_49269);
nand UO_4037 (O_4037,N_45144,N_47926);
nand UO_4038 (O_4038,N_49077,N_49320);
nand UO_4039 (O_4039,N_46578,N_47629);
and UO_4040 (O_4040,N_49395,N_45506);
or UO_4041 (O_4041,N_49868,N_47118);
nor UO_4042 (O_4042,N_46959,N_46524);
nand UO_4043 (O_4043,N_46379,N_47318);
xnor UO_4044 (O_4044,N_47323,N_49051);
and UO_4045 (O_4045,N_46611,N_45471);
xor UO_4046 (O_4046,N_49800,N_46534);
nand UO_4047 (O_4047,N_49733,N_47107);
xor UO_4048 (O_4048,N_47674,N_46166);
or UO_4049 (O_4049,N_49963,N_45657);
and UO_4050 (O_4050,N_47590,N_48299);
xnor UO_4051 (O_4051,N_46773,N_49801);
and UO_4052 (O_4052,N_46743,N_49050);
xor UO_4053 (O_4053,N_46495,N_46129);
nand UO_4054 (O_4054,N_49183,N_48339);
nor UO_4055 (O_4055,N_49772,N_46738);
xnor UO_4056 (O_4056,N_47245,N_45143);
xnor UO_4057 (O_4057,N_48442,N_45670);
and UO_4058 (O_4058,N_47021,N_48590);
nand UO_4059 (O_4059,N_49861,N_48402);
and UO_4060 (O_4060,N_47561,N_45672);
nor UO_4061 (O_4061,N_45112,N_49205);
xor UO_4062 (O_4062,N_47035,N_47456);
and UO_4063 (O_4063,N_49033,N_47014);
xor UO_4064 (O_4064,N_46620,N_45866);
xor UO_4065 (O_4065,N_48849,N_45324);
nand UO_4066 (O_4066,N_45488,N_49323);
nor UO_4067 (O_4067,N_45929,N_47775);
nor UO_4068 (O_4068,N_45705,N_49592);
and UO_4069 (O_4069,N_49687,N_47314);
nand UO_4070 (O_4070,N_48630,N_48538);
nor UO_4071 (O_4071,N_47445,N_46835);
xor UO_4072 (O_4072,N_49047,N_48892);
nand UO_4073 (O_4073,N_49476,N_47115);
nor UO_4074 (O_4074,N_48278,N_47490);
and UO_4075 (O_4075,N_45331,N_45298);
nor UO_4076 (O_4076,N_48312,N_46529);
or UO_4077 (O_4077,N_45902,N_45775);
nor UO_4078 (O_4078,N_48464,N_47696);
nand UO_4079 (O_4079,N_48295,N_48898);
xor UO_4080 (O_4080,N_49630,N_46061);
or UO_4081 (O_4081,N_47864,N_48555);
xnor UO_4082 (O_4082,N_47208,N_45885);
nand UO_4083 (O_4083,N_47721,N_48776);
and UO_4084 (O_4084,N_49824,N_48986);
nand UO_4085 (O_4085,N_49670,N_48001);
xnor UO_4086 (O_4086,N_47072,N_48506);
nand UO_4087 (O_4087,N_46168,N_47106);
and UO_4088 (O_4088,N_45118,N_47856);
and UO_4089 (O_4089,N_46423,N_48254);
nand UO_4090 (O_4090,N_47462,N_45425);
or UO_4091 (O_4091,N_49030,N_49577);
nor UO_4092 (O_4092,N_46171,N_49291);
nand UO_4093 (O_4093,N_46582,N_47073);
nor UO_4094 (O_4094,N_45285,N_49164);
xnor UO_4095 (O_4095,N_45583,N_49127);
or UO_4096 (O_4096,N_45492,N_49778);
and UO_4097 (O_4097,N_46554,N_45443);
or UO_4098 (O_4098,N_45612,N_49570);
or UO_4099 (O_4099,N_48055,N_46411);
or UO_4100 (O_4100,N_48862,N_47430);
or UO_4101 (O_4101,N_48983,N_48561);
nor UO_4102 (O_4102,N_45195,N_48624);
xnor UO_4103 (O_4103,N_47214,N_48419);
or UO_4104 (O_4104,N_46443,N_48778);
or UO_4105 (O_4105,N_47364,N_46994);
and UO_4106 (O_4106,N_45088,N_45340);
nand UO_4107 (O_4107,N_48005,N_49167);
xnor UO_4108 (O_4108,N_47406,N_46671);
or UO_4109 (O_4109,N_48918,N_47679);
or UO_4110 (O_4110,N_47581,N_49825);
nand UO_4111 (O_4111,N_48925,N_47390);
nand UO_4112 (O_4112,N_49421,N_46336);
or UO_4113 (O_4113,N_47715,N_45589);
and UO_4114 (O_4114,N_47992,N_46233);
nand UO_4115 (O_4115,N_48288,N_45514);
xnor UO_4116 (O_4116,N_48073,N_48511);
nand UO_4117 (O_4117,N_45276,N_46409);
or UO_4118 (O_4118,N_45332,N_49624);
xnor UO_4119 (O_4119,N_49803,N_46450);
nand UO_4120 (O_4120,N_49378,N_46955);
xnor UO_4121 (O_4121,N_48187,N_45835);
and UO_4122 (O_4122,N_47572,N_48515);
or UO_4123 (O_4123,N_46376,N_46462);
nor UO_4124 (O_4124,N_45564,N_49471);
nor UO_4125 (O_4125,N_47759,N_45247);
or UO_4126 (O_4126,N_47386,N_48598);
nor UO_4127 (O_4127,N_46915,N_48764);
or UO_4128 (O_4128,N_45675,N_47781);
or UO_4129 (O_4129,N_47938,N_47888);
and UO_4130 (O_4130,N_46820,N_48297);
or UO_4131 (O_4131,N_49659,N_48647);
xnor UO_4132 (O_4132,N_46036,N_48625);
or UO_4133 (O_4133,N_47539,N_45939);
xor UO_4134 (O_4134,N_49456,N_48044);
xnor UO_4135 (O_4135,N_48246,N_45934);
nor UO_4136 (O_4136,N_46316,N_46583);
and UO_4137 (O_4137,N_48631,N_47657);
nor UO_4138 (O_4138,N_49271,N_47273);
or UO_4139 (O_4139,N_49859,N_47004);
or UO_4140 (O_4140,N_45684,N_46821);
or UO_4141 (O_4141,N_49539,N_49004);
xor UO_4142 (O_4142,N_48853,N_46746);
or UO_4143 (O_4143,N_48246,N_48330);
nand UO_4144 (O_4144,N_49956,N_48790);
and UO_4145 (O_4145,N_47077,N_46654);
or UO_4146 (O_4146,N_49867,N_45871);
nor UO_4147 (O_4147,N_49040,N_49707);
nor UO_4148 (O_4148,N_46633,N_46626);
nor UO_4149 (O_4149,N_45665,N_47881);
nand UO_4150 (O_4150,N_48566,N_49089);
nand UO_4151 (O_4151,N_48409,N_45022);
xnor UO_4152 (O_4152,N_47865,N_49327);
or UO_4153 (O_4153,N_47522,N_49541);
or UO_4154 (O_4154,N_47231,N_45800);
xor UO_4155 (O_4155,N_46550,N_48108);
and UO_4156 (O_4156,N_45618,N_48879);
and UO_4157 (O_4157,N_49031,N_48445);
xnor UO_4158 (O_4158,N_49519,N_48258);
nor UO_4159 (O_4159,N_47871,N_48066);
xnor UO_4160 (O_4160,N_46398,N_48034);
xor UO_4161 (O_4161,N_45117,N_46718);
and UO_4162 (O_4162,N_46279,N_46388);
or UO_4163 (O_4163,N_45313,N_46333);
and UO_4164 (O_4164,N_49282,N_46925);
nand UO_4165 (O_4165,N_45697,N_47036);
nand UO_4166 (O_4166,N_49520,N_48922);
nand UO_4167 (O_4167,N_47450,N_45777);
nor UO_4168 (O_4168,N_46708,N_46351);
or UO_4169 (O_4169,N_48697,N_49402);
xnor UO_4170 (O_4170,N_45460,N_45694);
or UO_4171 (O_4171,N_45120,N_47024);
nor UO_4172 (O_4172,N_47529,N_49252);
and UO_4173 (O_4173,N_46023,N_47167);
nand UO_4174 (O_4174,N_47581,N_45754);
and UO_4175 (O_4175,N_45429,N_48626);
nor UO_4176 (O_4176,N_47287,N_47286);
xnor UO_4177 (O_4177,N_46988,N_46673);
and UO_4178 (O_4178,N_46391,N_48182);
xnor UO_4179 (O_4179,N_46498,N_46788);
nor UO_4180 (O_4180,N_46733,N_47786);
xor UO_4181 (O_4181,N_46990,N_48231);
xnor UO_4182 (O_4182,N_45031,N_47313);
and UO_4183 (O_4183,N_45088,N_45245);
xor UO_4184 (O_4184,N_46726,N_49166);
nor UO_4185 (O_4185,N_45628,N_46814);
or UO_4186 (O_4186,N_48807,N_46901);
xnor UO_4187 (O_4187,N_45407,N_45421);
and UO_4188 (O_4188,N_45851,N_48248);
or UO_4189 (O_4189,N_47923,N_47114);
or UO_4190 (O_4190,N_46560,N_46459);
xnor UO_4191 (O_4191,N_46914,N_47247);
nor UO_4192 (O_4192,N_45841,N_49168);
and UO_4193 (O_4193,N_46955,N_46790);
xor UO_4194 (O_4194,N_46645,N_49687);
nor UO_4195 (O_4195,N_49055,N_47283);
nor UO_4196 (O_4196,N_45016,N_47945);
nand UO_4197 (O_4197,N_45813,N_46511);
nand UO_4198 (O_4198,N_46259,N_48118);
nand UO_4199 (O_4199,N_45028,N_49444);
xnor UO_4200 (O_4200,N_49748,N_45531);
nor UO_4201 (O_4201,N_45731,N_46145);
nand UO_4202 (O_4202,N_49251,N_49257);
nand UO_4203 (O_4203,N_49753,N_46653);
or UO_4204 (O_4204,N_45480,N_49863);
or UO_4205 (O_4205,N_47931,N_47228);
xnor UO_4206 (O_4206,N_46051,N_46268);
nor UO_4207 (O_4207,N_48232,N_46016);
nor UO_4208 (O_4208,N_45276,N_46627);
nand UO_4209 (O_4209,N_45967,N_48845);
xnor UO_4210 (O_4210,N_45211,N_46878);
xor UO_4211 (O_4211,N_48668,N_46691);
or UO_4212 (O_4212,N_49660,N_46964);
nand UO_4213 (O_4213,N_47148,N_46720);
or UO_4214 (O_4214,N_47652,N_47632);
xor UO_4215 (O_4215,N_47360,N_47663);
nand UO_4216 (O_4216,N_48330,N_46209);
and UO_4217 (O_4217,N_47705,N_49098);
or UO_4218 (O_4218,N_45293,N_48051);
xnor UO_4219 (O_4219,N_45773,N_48902);
nor UO_4220 (O_4220,N_45521,N_49122);
or UO_4221 (O_4221,N_46624,N_48744);
and UO_4222 (O_4222,N_45659,N_48641);
nor UO_4223 (O_4223,N_46903,N_46782);
and UO_4224 (O_4224,N_46732,N_45680);
or UO_4225 (O_4225,N_46127,N_49791);
and UO_4226 (O_4226,N_47115,N_47877);
or UO_4227 (O_4227,N_45890,N_48984);
and UO_4228 (O_4228,N_46089,N_47186);
and UO_4229 (O_4229,N_47413,N_49465);
and UO_4230 (O_4230,N_46658,N_48634);
or UO_4231 (O_4231,N_48397,N_49816);
nand UO_4232 (O_4232,N_49821,N_46933);
and UO_4233 (O_4233,N_48392,N_49490);
nand UO_4234 (O_4234,N_47996,N_45543);
or UO_4235 (O_4235,N_46976,N_45541);
or UO_4236 (O_4236,N_48678,N_46771);
or UO_4237 (O_4237,N_49926,N_47302);
and UO_4238 (O_4238,N_48417,N_48265);
nand UO_4239 (O_4239,N_48433,N_48609);
nor UO_4240 (O_4240,N_49400,N_48227);
and UO_4241 (O_4241,N_46341,N_45215);
nor UO_4242 (O_4242,N_49298,N_47758);
nand UO_4243 (O_4243,N_47192,N_45884);
nand UO_4244 (O_4244,N_46299,N_48800);
nand UO_4245 (O_4245,N_46255,N_46655);
nand UO_4246 (O_4246,N_49920,N_49849);
or UO_4247 (O_4247,N_47721,N_47779);
xor UO_4248 (O_4248,N_48749,N_48365);
nor UO_4249 (O_4249,N_45969,N_47676);
or UO_4250 (O_4250,N_48165,N_47155);
and UO_4251 (O_4251,N_46413,N_45499);
nor UO_4252 (O_4252,N_46399,N_49145);
nand UO_4253 (O_4253,N_46677,N_47166);
nor UO_4254 (O_4254,N_49336,N_49682);
xor UO_4255 (O_4255,N_48765,N_45549);
nor UO_4256 (O_4256,N_49314,N_49045);
nand UO_4257 (O_4257,N_49538,N_47260);
nor UO_4258 (O_4258,N_47960,N_47490);
nand UO_4259 (O_4259,N_49579,N_46269);
nand UO_4260 (O_4260,N_49695,N_45449);
nand UO_4261 (O_4261,N_47283,N_45867);
and UO_4262 (O_4262,N_47229,N_46282);
nand UO_4263 (O_4263,N_48836,N_48425);
nor UO_4264 (O_4264,N_49203,N_47764);
xnor UO_4265 (O_4265,N_48042,N_45603);
and UO_4266 (O_4266,N_45584,N_47001);
nor UO_4267 (O_4267,N_45758,N_49778);
xor UO_4268 (O_4268,N_45302,N_49377);
nand UO_4269 (O_4269,N_45202,N_48344);
nand UO_4270 (O_4270,N_48935,N_49639);
nand UO_4271 (O_4271,N_45769,N_45158);
nand UO_4272 (O_4272,N_47920,N_46592);
or UO_4273 (O_4273,N_47132,N_46594);
xnor UO_4274 (O_4274,N_45833,N_45225);
xnor UO_4275 (O_4275,N_49635,N_48502);
nor UO_4276 (O_4276,N_49867,N_45349);
and UO_4277 (O_4277,N_45518,N_47006);
nand UO_4278 (O_4278,N_45052,N_45842);
and UO_4279 (O_4279,N_46132,N_46062);
and UO_4280 (O_4280,N_47175,N_49436);
nand UO_4281 (O_4281,N_47547,N_46709);
nand UO_4282 (O_4282,N_45107,N_47272);
nor UO_4283 (O_4283,N_48391,N_49219);
or UO_4284 (O_4284,N_49116,N_45498);
and UO_4285 (O_4285,N_47143,N_46923);
xnor UO_4286 (O_4286,N_48828,N_48291);
or UO_4287 (O_4287,N_46924,N_48108);
nand UO_4288 (O_4288,N_46632,N_45035);
nand UO_4289 (O_4289,N_46287,N_47441);
or UO_4290 (O_4290,N_48989,N_45945);
and UO_4291 (O_4291,N_48495,N_45143);
or UO_4292 (O_4292,N_48948,N_47929);
or UO_4293 (O_4293,N_49168,N_46489);
or UO_4294 (O_4294,N_47743,N_47958);
and UO_4295 (O_4295,N_47881,N_47070);
or UO_4296 (O_4296,N_45271,N_46386);
and UO_4297 (O_4297,N_45801,N_47338);
nor UO_4298 (O_4298,N_47385,N_48725);
nor UO_4299 (O_4299,N_47689,N_48283);
xor UO_4300 (O_4300,N_45642,N_45559);
nor UO_4301 (O_4301,N_49073,N_46598);
and UO_4302 (O_4302,N_48300,N_48746);
and UO_4303 (O_4303,N_45121,N_47418);
or UO_4304 (O_4304,N_47676,N_49607);
or UO_4305 (O_4305,N_49565,N_45736);
or UO_4306 (O_4306,N_46952,N_49831);
nand UO_4307 (O_4307,N_45958,N_49844);
nand UO_4308 (O_4308,N_49744,N_48198);
or UO_4309 (O_4309,N_47007,N_48947);
and UO_4310 (O_4310,N_46727,N_46216);
nor UO_4311 (O_4311,N_49574,N_48464);
or UO_4312 (O_4312,N_49844,N_46849);
or UO_4313 (O_4313,N_48756,N_48393);
and UO_4314 (O_4314,N_47786,N_46845);
nor UO_4315 (O_4315,N_45430,N_46707);
nand UO_4316 (O_4316,N_46693,N_47000);
or UO_4317 (O_4317,N_48745,N_45893);
nor UO_4318 (O_4318,N_47714,N_49568);
nor UO_4319 (O_4319,N_47592,N_47101);
xor UO_4320 (O_4320,N_47433,N_45163);
nor UO_4321 (O_4321,N_46192,N_48564);
and UO_4322 (O_4322,N_49864,N_46002);
nand UO_4323 (O_4323,N_46047,N_46538);
and UO_4324 (O_4324,N_45377,N_49811);
nand UO_4325 (O_4325,N_45681,N_48818);
and UO_4326 (O_4326,N_46752,N_45330);
xor UO_4327 (O_4327,N_49423,N_46176);
xor UO_4328 (O_4328,N_49075,N_48219);
xnor UO_4329 (O_4329,N_48107,N_45032);
xor UO_4330 (O_4330,N_47468,N_45993);
xor UO_4331 (O_4331,N_47566,N_49803);
xnor UO_4332 (O_4332,N_48351,N_48752);
nor UO_4333 (O_4333,N_46802,N_49745);
or UO_4334 (O_4334,N_48299,N_48087);
or UO_4335 (O_4335,N_46729,N_45045);
nand UO_4336 (O_4336,N_48702,N_45065);
and UO_4337 (O_4337,N_46497,N_48092);
or UO_4338 (O_4338,N_45981,N_46636);
nand UO_4339 (O_4339,N_45194,N_49010);
or UO_4340 (O_4340,N_49491,N_48330);
nor UO_4341 (O_4341,N_49260,N_49751);
and UO_4342 (O_4342,N_48797,N_47645);
and UO_4343 (O_4343,N_46571,N_46432);
xor UO_4344 (O_4344,N_45300,N_48666);
or UO_4345 (O_4345,N_46697,N_47526);
and UO_4346 (O_4346,N_47057,N_48221);
nand UO_4347 (O_4347,N_49934,N_47825);
nor UO_4348 (O_4348,N_49913,N_49060);
nor UO_4349 (O_4349,N_49470,N_47637);
and UO_4350 (O_4350,N_46399,N_47419);
xnor UO_4351 (O_4351,N_49833,N_46571);
nand UO_4352 (O_4352,N_49989,N_45490);
nand UO_4353 (O_4353,N_45708,N_47110);
xor UO_4354 (O_4354,N_49986,N_45555);
nand UO_4355 (O_4355,N_48828,N_47116);
nor UO_4356 (O_4356,N_47612,N_45573);
or UO_4357 (O_4357,N_45778,N_47191);
xor UO_4358 (O_4358,N_48200,N_47129);
nor UO_4359 (O_4359,N_47730,N_46399);
nand UO_4360 (O_4360,N_46999,N_49703);
nor UO_4361 (O_4361,N_47756,N_48249);
xnor UO_4362 (O_4362,N_46725,N_45177);
nand UO_4363 (O_4363,N_47489,N_47419);
xnor UO_4364 (O_4364,N_48441,N_48488);
xnor UO_4365 (O_4365,N_46108,N_46570);
and UO_4366 (O_4366,N_47999,N_47105);
nor UO_4367 (O_4367,N_48412,N_46735);
nand UO_4368 (O_4368,N_48962,N_45815);
or UO_4369 (O_4369,N_45691,N_48365);
nand UO_4370 (O_4370,N_48381,N_45094);
nor UO_4371 (O_4371,N_45227,N_49139);
nor UO_4372 (O_4372,N_47202,N_46446);
and UO_4373 (O_4373,N_48089,N_46085);
nand UO_4374 (O_4374,N_45503,N_48432);
nand UO_4375 (O_4375,N_49299,N_48762);
or UO_4376 (O_4376,N_49496,N_47184);
nor UO_4377 (O_4377,N_48241,N_47164);
and UO_4378 (O_4378,N_46736,N_45233);
or UO_4379 (O_4379,N_49361,N_48840);
nand UO_4380 (O_4380,N_49987,N_48565);
xor UO_4381 (O_4381,N_49233,N_45237);
nand UO_4382 (O_4382,N_48596,N_47324);
or UO_4383 (O_4383,N_47969,N_48331);
nor UO_4384 (O_4384,N_45169,N_45448);
xor UO_4385 (O_4385,N_49189,N_49983);
xor UO_4386 (O_4386,N_48795,N_48997);
or UO_4387 (O_4387,N_45551,N_45377);
nand UO_4388 (O_4388,N_47814,N_45370);
and UO_4389 (O_4389,N_46045,N_47528);
xnor UO_4390 (O_4390,N_49871,N_46073);
nor UO_4391 (O_4391,N_46858,N_46030);
and UO_4392 (O_4392,N_47702,N_45894);
nor UO_4393 (O_4393,N_47546,N_45451);
xor UO_4394 (O_4394,N_49568,N_46770);
and UO_4395 (O_4395,N_46737,N_45391);
nor UO_4396 (O_4396,N_47843,N_45642);
xor UO_4397 (O_4397,N_48487,N_47601);
xnor UO_4398 (O_4398,N_47237,N_45384);
nor UO_4399 (O_4399,N_45945,N_47453);
nand UO_4400 (O_4400,N_49265,N_47116);
or UO_4401 (O_4401,N_47719,N_45251);
nand UO_4402 (O_4402,N_46732,N_49582);
or UO_4403 (O_4403,N_45417,N_45920);
nand UO_4404 (O_4404,N_47925,N_48281);
nor UO_4405 (O_4405,N_48777,N_49799);
nand UO_4406 (O_4406,N_49382,N_47403);
and UO_4407 (O_4407,N_45342,N_49657);
nand UO_4408 (O_4408,N_46692,N_47503);
xor UO_4409 (O_4409,N_47164,N_47589);
and UO_4410 (O_4410,N_47757,N_45818);
nand UO_4411 (O_4411,N_46162,N_45350);
xor UO_4412 (O_4412,N_45147,N_45965);
nand UO_4413 (O_4413,N_47127,N_49259);
or UO_4414 (O_4414,N_47868,N_49100);
nand UO_4415 (O_4415,N_46816,N_49905);
nor UO_4416 (O_4416,N_48629,N_49654);
and UO_4417 (O_4417,N_45119,N_46918);
nand UO_4418 (O_4418,N_47502,N_46926);
or UO_4419 (O_4419,N_46092,N_47394);
and UO_4420 (O_4420,N_48671,N_47668);
or UO_4421 (O_4421,N_49861,N_45484);
and UO_4422 (O_4422,N_48143,N_48842);
or UO_4423 (O_4423,N_48623,N_45552);
nor UO_4424 (O_4424,N_45656,N_48326);
xnor UO_4425 (O_4425,N_46758,N_48090);
nand UO_4426 (O_4426,N_47757,N_47664);
xnor UO_4427 (O_4427,N_46675,N_45140);
nand UO_4428 (O_4428,N_47424,N_49249);
xor UO_4429 (O_4429,N_48806,N_46848);
nand UO_4430 (O_4430,N_48861,N_47456);
xor UO_4431 (O_4431,N_45271,N_45693);
nor UO_4432 (O_4432,N_49891,N_45073);
xnor UO_4433 (O_4433,N_49825,N_45285);
xnor UO_4434 (O_4434,N_45314,N_45450);
nand UO_4435 (O_4435,N_49424,N_47975);
nand UO_4436 (O_4436,N_45989,N_47745);
nor UO_4437 (O_4437,N_49049,N_46272);
or UO_4438 (O_4438,N_46071,N_45503);
and UO_4439 (O_4439,N_49111,N_47912);
and UO_4440 (O_4440,N_45457,N_47742);
nor UO_4441 (O_4441,N_49378,N_47703);
and UO_4442 (O_4442,N_47532,N_45574);
nor UO_4443 (O_4443,N_49500,N_49676);
and UO_4444 (O_4444,N_47228,N_49133);
xor UO_4445 (O_4445,N_47601,N_49258);
and UO_4446 (O_4446,N_47010,N_48540);
xor UO_4447 (O_4447,N_49514,N_45760);
xor UO_4448 (O_4448,N_47719,N_46567);
nor UO_4449 (O_4449,N_48979,N_45781);
nor UO_4450 (O_4450,N_46301,N_45304);
or UO_4451 (O_4451,N_45971,N_49670);
nor UO_4452 (O_4452,N_49915,N_47068);
nor UO_4453 (O_4453,N_46124,N_48756);
or UO_4454 (O_4454,N_47392,N_47377);
xor UO_4455 (O_4455,N_46876,N_45569);
and UO_4456 (O_4456,N_47409,N_49722);
nand UO_4457 (O_4457,N_49787,N_46805);
and UO_4458 (O_4458,N_45518,N_48653);
nand UO_4459 (O_4459,N_47617,N_45177);
or UO_4460 (O_4460,N_47015,N_49359);
xnor UO_4461 (O_4461,N_49432,N_47049);
xor UO_4462 (O_4462,N_49056,N_49873);
nand UO_4463 (O_4463,N_45701,N_48400);
nand UO_4464 (O_4464,N_45198,N_49770);
xnor UO_4465 (O_4465,N_46592,N_49513);
nor UO_4466 (O_4466,N_45469,N_49785);
and UO_4467 (O_4467,N_48461,N_45072);
nor UO_4468 (O_4468,N_46862,N_45239);
or UO_4469 (O_4469,N_47420,N_48202);
nor UO_4470 (O_4470,N_46339,N_46739);
and UO_4471 (O_4471,N_47068,N_47262);
or UO_4472 (O_4472,N_47819,N_46914);
or UO_4473 (O_4473,N_46959,N_47840);
xor UO_4474 (O_4474,N_48000,N_48359);
xnor UO_4475 (O_4475,N_45980,N_47101);
nand UO_4476 (O_4476,N_49772,N_45125);
xnor UO_4477 (O_4477,N_47261,N_48565);
and UO_4478 (O_4478,N_45270,N_49918);
xor UO_4479 (O_4479,N_45259,N_47070);
or UO_4480 (O_4480,N_48219,N_46853);
nor UO_4481 (O_4481,N_49725,N_48751);
nand UO_4482 (O_4482,N_48541,N_45273);
or UO_4483 (O_4483,N_47080,N_46157);
and UO_4484 (O_4484,N_47302,N_46122);
and UO_4485 (O_4485,N_46458,N_48971);
nor UO_4486 (O_4486,N_48767,N_46076);
and UO_4487 (O_4487,N_45553,N_46594);
xnor UO_4488 (O_4488,N_47001,N_48428);
or UO_4489 (O_4489,N_45209,N_49587);
nand UO_4490 (O_4490,N_47403,N_49376);
nor UO_4491 (O_4491,N_46743,N_46420);
or UO_4492 (O_4492,N_45802,N_46682);
nor UO_4493 (O_4493,N_47429,N_46852);
or UO_4494 (O_4494,N_47694,N_46431);
nor UO_4495 (O_4495,N_46622,N_45113);
and UO_4496 (O_4496,N_45060,N_45462);
nor UO_4497 (O_4497,N_46616,N_47326);
and UO_4498 (O_4498,N_45728,N_47368);
nand UO_4499 (O_4499,N_48973,N_45233);
nand UO_4500 (O_4500,N_49988,N_46048);
xnor UO_4501 (O_4501,N_48178,N_45138);
and UO_4502 (O_4502,N_46910,N_48101);
xor UO_4503 (O_4503,N_47795,N_45520);
or UO_4504 (O_4504,N_49653,N_48545);
and UO_4505 (O_4505,N_45716,N_49682);
or UO_4506 (O_4506,N_47787,N_48371);
xor UO_4507 (O_4507,N_49845,N_46986);
and UO_4508 (O_4508,N_47943,N_47828);
nor UO_4509 (O_4509,N_48975,N_47286);
nor UO_4510 (O_4510,N_49052,N_46732);
or UO_4511 (O_4511,N_48152,N_48461);
nor UO_4512 (O_4512,N_49685,N_46073);
xor UO_4513 (O_4513,N_47257,N_49140);
xor UO_4514 (O_4514,N_47239,N_48743);
and UO_4515 (O_4515,N_47184,N_48790);
nand UO_4516 (O_4516,N_45544,N_46154);
or UO_4517 (O_4517,N_45849,N_47070);
nand UO_4518 (O_4518,N_46637,N_45431);
nor UO_4519 (O_4519,N_47541,N_45975);
xnor UO_4520 (O_4520,N_48739,N_49654);
or UO_4521 (O_4521,N_47297,N_49901);
nand UO_4522 (O_4522,N_47403,N_45692);
xnor UO_4523 (O_4523,N_46814,N_49985);
or UO_4524 (O_4524,N_46750,N_49764);
nand UO_4525 (O_4525,N_46577,N_48056);
or UO_4526 (O_4526,N_48380,N_47387);
nand UO_4527 (O_4527,N_46105,N_48851);
nor UO_4528 (O_4528,N_46606,N_47210);
nor UO_4529 (O_4529,N_46379,N_49623);
nor UO_4530 (O_4530,N_45064,N_49254);
and UO_4531 (O_4531,N_48234,N_46743);
xnor UO_4532 (O_4532,N_48386,N_47233);
xnor UO_4533 (O_4533,N_46278,N_45041);
xor UO_4534 (O_4534,N_46041,N_45824);
or UO_4535 (O_4535,N_46363,N_48526);
xnor UO_4536 (O_4536,N_49836,N_49557);
nand UO_4537 (O_4537,N_45383,N_45514);
xor UO_4538 (O_4538,N_46767,N_46418);
nor UO_4539 (O_4539,N_45918,N_49382);
and UO_4540 (O_4540,N_49432,N_46632);
xor UO_4541 (O_4541,N_45844,N_46608);
xor UO_4542 (O_4542,N_47671,N_47034);
nand UO_4543 (O_4543,N_48542,N_47352);
nand UO_4544 (O_4544,N_48549,N_49301);
or UO_4545 (O_4545,N_46512,N_45253);
or UO_4546 (O_4546,N_46959,N_47898);
nand UO_4547 (O_4547,N_49664,N_49938);
nand UO_4548 (O_4548,N_49397,N_46005);
xnor UO_4549 (O_4549,N_47417,N_47938);
or UO_4550 (O_4550,N_47996,N_49069);
nor UO_4551 (O_4551,N_46766,N_49132);
nand UO_4552 (O_4552,N_47819,N_47539);
and UO_4553 (O_4553,N_48243,N_47548);
and UO_4554 (O_4554,N_46063,N_46567);
nor UO_4555 (O_4555,N_47228,N_48437);
nor UO_4556 (O_4556,N_45879,N_49668);
nand UO_4557 (O_4557,N_47094,N_47634);
or UO_4558 (O_4558,N_49051,N_46270);
or UO_4559 (O_4559,N_49706,N_47564);
nand UO_4560 (O_4560,N_47154,N_48503);
and UO_4561 (O_4561,N_45528,N_46114);
and UO_4562 (O_4562,N_48267,N_45169);
and UO_4563 (O_4563,N_47495,N_45876);
nand UO_4564 (O_4564,N_46422,N_49316);
xor UO_4565 (O_4565,N_45313,N_47178);
xnor UO_4566 (O_4566,N_46946,N_49761);
nand UO_4567 (O_4567,N_46088,N_48835);
nand UO_4568 (O_4568,N_49819,N_45703);
or UO_4569 (O_4569,N_49325,N_45062);
nor UO_4570 (O_4570,N_48166,N_48514);
nand UO_4571 (O_4571,N_49252,N_47815);
xor UO_4572 (O_4572,N_49224,N_47951);
nor UO_4573 (O_4573,N_47301,N_48434);
xor UO_4574 (O_4574,N_47605,N_49132);
xnor UO_4575 (O_4575,N_46091,N_45453);
nand UO_4576 (O_4576,N_49991,N_45553);
and UO_4577 (O_4577,N_48767,N_46257);
and UO_4578 (O_4578,N_49649,N_48967);
nor UO_4579 (O_4579,N_46294,N_49794);
and UO_4580 (O_4580,N_48817,N_49539);
xnor UO_4581 (O_4581,N_45299,N_46737);
xnor UO_4582 (O_4582,N_48446,N_47858);
xnor UO_4583 (O_4583,N_45140,N_46545);
xor UO_4584 (O_4584,N_46349,N_49892);
or UO_4585 (O_4585,N_46189,N_47758);
nand UO_4586 (O_4586,N_47383,N_45574);
nor UO_4587 (O_4587,N_45371,N_47925);
and UO_4588 (O_4588,N_45256,N_45965);
nand UO_4589 (O_4589,N_46586,N_47192);
or UO_4590 (O_4590,N_46306,N_45033);
nand UO_4591 (O_4591,N_48575,N_48938);
nand UO_4592 (O_4592,N_46421,N_46398);
nand UO_4593 (O_4593,N_47562,N_49639);
and UO_4594 (O_4594,N_45541,N_45671);
or UO_4595 (O_4595,N_47018,N_49374);
nor UO_4596 (O_4596,N_47733,N_45941);
and UO_4597 (O_4597,N_47005,N_47676);
nand UO_4598 (O_4598,N_46015,N_47009);
nor UO_4599 (O_4599,N_46772,N_49832);
xor UO_4600 (O_4600,N_46945,N_48875);
xnor UO_4601 (O_4601,N_49205,N_48256);
nand UO_4602 (O_4602,N_45948,N_47030);
and UO_4603 (O_4603,N_45268,N_48261);
nor UO_4604 (O_4604,N_47597,N_48017);
or UO_4605 (O_4605,N_49486,N_48031);
nand UO_4606 (O_4606,N_49670,N_49117);
and UO_4607 (O_4607,N_49088,N_48040);
and UO_4608 (O_4608,N_47846,N_48528);
or UO_4609 (O_4609,N_45227,N_49577);
nor UO_4610 (O_4610,N_46705,N_49276);
nor UO_4611 (O_4611,N_46370,N_45067);
nor UO_4612 (O_4612,N_47173,N_47248);
and UO_4613 (O_4613,N_46263,N_45523);
nand UO_4614 (O_4614,N_47516,N_46115);
and UO_4615 (O_4615,N_48961,N_47885);
nand UO_4616 (O_4616,N_49948,N_48270);
nand UO_4617 (O_4617,N_46565,N_46890);
nor UO_4618 (O_4618,N_47203,N_48082);
xnor UO_4619 (O_4619,N_46766,N_46579);
xor UO_4620 (O_4620,N_45868,N_46962);
nor UO_4621 (O_4621,N_49730,N_48320);
nand UO_4622 (O_4622,N_47852,N_47198);
nor UO_4623 (O_4623,N_46346,N_46805);
and UO_4624 (O_4624,N_45707,N_45115);
nand UO_4625 (O_4625,N_46690,N_48308);
nor UO_4626 (O_4626,N_45460,N_47470);
or UO_4627 (O_4627,N_47803,N_49598);
nor UO_4628 (O_4628,N_48089,N_46916);
nor UO_4629 (O_4629,N_45291,N_49001);
or UO_4630 (O_4630,N_46375,N_47254);
xnor UO_4631 (O_4631,N_48894,N_47879);
nand UO_4632 (O_4632,N_49856,N_46763);
nor UO_4633 (O_4633,N_45274,N_46061);
and UO_4634 (O_4634,N_47355,N_47725);
or UO_4635 (O_4635,N_48698,N_45026);
or UO_4636 (O_4636,N_49177,N_45836);
nor UO_4637 (O_4637,N_46714,N_46267);
or UO_4638 (O_4638,N_49313,N_46228);
xnor UO_4639 (O_4639,N_45812,N_45357);
xor UO_4640 (O_4640,N_49784,N_47549);
or UO_4641 (O_4641,N_49265,N_45117);
nor UO_4642 (O_4642,N_49875,N_45237);
nor UO_4643 (O_4643,N_46664,N_45402);
or UO_4644 (O_4644,N_46700,N_47315);
or UO_4645 (O_4645,N_48521,N_47802);
and UO_4646 (O_4646,N_49701,N_49077);
or UO_4647 (O_4647,N_48616,N_45585);
and UO_4648 (O_4648,N_47890,N_48004);
nor UO_4649 (O_4649,N_49408,N_46294);
and UO_4650 (O_4650,N_47551,N_47822);
nor UO_4651 (O_4651,N_46820,N_46238);
nand UO_4652 (O_4652,N_45128,N_45254);
nor UO_4653 (O_4653,N_49191,N_49193);
nor UO_4654 (O_4654,N_45134,N_47184);
or UO_4655 (O_4655,N_47208,N_45556);
nand UO_4656 (O_4656,N_48350,N_46265);
or UO_4657 (O_4657,N_49911,N_48144);
nand UO_4658 (O_4658,N_45465,N_49829);
nand UO_4659 (O_4659,N_47895,N_49815);
or UO_4660 (O_4660,N_46263,N_49578);
and UO_4661 (O_4661,N_47179,N_47442);
nor UO_4662 (O_4662,N_48969,N_45604);
or UO_4663 (O_4663,N_48421,N_46924);
and UO_4664 (O_4664,N_48239,N_47832);
nor UO_4665 (O_4665,N_49211,N_48190);
or UO_4666 (O_4666,N_45694,N_48972);
xor UO_4667 (O_4667,N_46206,N_45264);
and UO_4668 (O_4668,N_49649,N_48523);
xnor UO_4669 (O_4669,N_47474,N_48387);
nor UO_4670 (O_4670,N_46658,N_48714);
xnor UO_4671 (O_4671,N_46384,N_46706);
nor UO_4672 (O_4672,N_45758,N_47579);
nor UO_4673 (O_4673,N_48416,N_46533);
or UO_4674 (O_4674,N_47732,N_47491);
xor UO_4675 (O_4675,N_49721,N_49315);
nand UO_4676 (O_4676,N_45711,N_48720);
or UO_4677 (O_4677,N_46247,N_49170);
and UO_4678 (O_4678,N_46640,N_46082);
nor UO_4679 (O_4679,N_47536,N_45885);
and UO_4680 (O_4680,N_47611,N_48869);
nand UO_4681 (O_4681,N_48783,N_45980);
xor UO_4682 (O_4682,N_45056,N_49519);
nand UO_4683 (O_4683,N_46824,N_47169);
nor UO_4684 (O_4684,N_46000,N_46663);
xor UO_4685 (O_4685,N_48129,N_45743);
nand UO_4686 (O_4686,N_47055,N_49021);
xor UO_4687 (O_4687,N_48543,N_49009);
nor UO_4688 (O_4688,N_47523,N_49842);
nor UO_4689 (O_4689,N_49495,N_48074);
nor UO_4690 (O_4690,N_45461,N_47947);
and UO_4691 (O_4691,N_45377,N_49641);
xnor UO_4692 (O_4692,N_49894,N_45233);
xor UO_4693 (O_4693,N_48079,N_48262);
and UO_4694 (O_4694,N_49888,N_47486);
and UO_4695 (O_4695,N_46090,N_46945);
and UO_4696 (O_4696,N_49019,N_49324);
and UO_4697 (O_4697,N_49114,N_48784);
and UO_4698 (O_4698,N_45184,N_45013);
nand UO_4699 (O_4699,N_46924,N_49811);
or UO_4700 (O_4700,N_46686,N_46398);
and UO_4701 (O_4701,N_48119,N_47553);
xnor UO_4702 (O_4702,N_46487,N_45811);
xnor UO_4703 (O_4703,N_49839,N_49897);
nand UO_4704 (O_4704,N_49185,N_47691);
nand UO_4705 (O_4705,N_49021,N_49564);
nand UO_4706 (O_4706,N_49723,N_48500);
and UO_4707 (O_4707,N_49777,N_46062);
or UO_4708 (O_4708,N_47201,N_45691);
nor UO_4709 (O_4709,N_49880,N_47981);
or UO_4710 (O_4710,N_49623,N_48396);
and UO_4711 (O_4711,N_45977,N_47817);
nand UO_4712 (O_4712,N_45923,N_48707);
or UO_4713 (O_4713,N_47683,N_49493);
nor UO_4714 (O_4714,N_45151,N_48982);
xnor UO_4715 (O_4715,N_45888,N_48402);
xnor UO_4716 (O_4716,N_49197,N_45874);
nor UO_4717 (O_4717,N_47535,N_45184);
xnor UO_4718 (O_4718,N_46575,N_48256);
or UO_4719 (O_4719,N_46440,N_47399);
and UO_4720 (O_4720,N_49188,N_46685);
xor UO_4721 (O_4721,N_46485,N_48852);
nor UO_4722 (O_4722,N_48667,N_45806);
or UO_4723 (O_4723,N_46695,N_48682);
or UO_4724 (O_4724,N_49641,N_45738);
nand UO_4725 (O_4725,N_47196,N_49142);
xor UO_4726 (O_4726,N_45806,N_46867);
nand UO_4727 (O_4727,N_47586,N_48329);
and UO_4728 (O_4728,N_48380,N_49388);
and UO_4729 (O_4729,N_46874,N_47775);
and UO_4730 (O_4730,N_49409,N_47081);
nor UO_4731 (O_4731,N_45202,N_48626);
xor UO_4732 (O_4732,N_45779,N_48574);
xor UO_4733 (O_4733,N_48193,N_49863);
or UO_4734 (O_4734,N_49966,N_47782);
nand UO_4735 (O_4735,N_45697,N_45009);
and UO_4736 (O_4736,N_46242,N_48370);
and UO_4737 (O_4737,N_49074,N_45813);
xnor UO_4738 (O_4738,N_48820,N_49476);
or UO_4739 (O_4739,N_48192,N_47145);
nor UO_4740 (O_4740,N_46635,N_45659);
nand UO_4741 (O_4741,N_49335,N_45929);
nor UO_4742 (O_4742,N_45284,N_49468);
nand UO_4743 (O_4743,N_48765,N_47392);
nor UO_4744 (O_4744,N_45210,N_48590);
nor UO_4745 (O_4745,N_47485,N_45080);
xnor UO_4746 (O_4746,N_49682,N_48063);
nor UO_4747 (O_4747,N_46937,N_49968);
or UO_4748 (O_4748,N_46738,N_45317);
or UO_4749 (O_4749,N_46942,N_45017);
xor UO_4750 (O_4750,N_45177,N_48334);
nand UO_4751 (O_4751,N_49018,N_47440);
or UO_4752 (O_4752,N_46076,N_45389);
xor UO_4753 (O_4753,N_47741,N_45333);
and UO_4754 (O_4754,N_47467,N_46789);
and UO_4755 (O_4755,N_47757,N_47276);
xor UO_4756 (O_4756,N_49095,N_47814);
nand UO_4757 (O_4757,N_47233,N_49631);
nand UO_4758 (O_4758,N_48929,N_48347);
and UO_4759 (O_4759,N_45201,N_46991);
and UO_4760 (O_4760,N_49843,N_46305);
nor UO_4761 (O_4761,N_46999,N_49429);
xnor UO_4762 (O_4762,N_47854,N_47746);
or UO_4763 (O_4763,N_45133,N_47956);
and UO_4764 (O_4764,N_45203,N_47055);
or UO_4765 (O_4765,N_48153,N_48691);
and UO_4766 (O_4766,N_46103,N_45115);
and UO_4767 (O_4767,N_47051,N_47381);
xnor UO_4768 (O_4768,N_47151,N_48498);
xor UO_4769 (O_4769,N_49726,N_49177);
xnor UO_4770 (O_4770,N_45804,N_48491);
and UO_4771 (O_4771,N_45958,N_46121);
xnor UO_4772 (O_4772,N_47570,N_47213);
or UO_4773 (O_4773,N_45311,N_45538);
or UO_4774 (O_4774,N_45194,N_46353);
and UO_4775 (O_4775,N_49631,N_47271);
or UO_4776 (O_4776,N_45329,N_47773);
or UO_4777 (O_4777,N_48707,N_47872);
or UO_4778 (O_4778,N_48829,N_48163);
nand UO_4779 (O_4779,N_48042,N_46367);
nand UO_4780 (O_4780,N_49326,N_45568);
nand UO_4781 (O_4781,N_47066,N_48044);
nor UO_4782 (O_4782,N_47014,N_46072);
nand UO_4783 (O_4783,N_46673,N_48053);
or UO_4784 (O_4784,N_46056,N_46428);
xor UO_4785 (O_4785,N_48092,N_49753);
xnor UO_4786 (O_4786,N_47101,N_49344);
xor UO_4787 (O_4787,N_46591,N_48321);
nand UO_4788 (O_4788,N_46351,N_45075);
and UO_4789 (O_4789,N_48293,N_46156);
nor UO_4790 (O_4790,N_46126,N_46972);
and UO_4791 (O_4791,N_46918,N_48498);
xnor UO_4792 (O_4792,N_49803,N_49642);
nand UO_4793 (O_4793,N_49751,N_49068);
and UO_4794 (O_4794,N_46990,N_48075);
nor UO_4795 (O_4795,N_47352,N_47473);
xor UO_4796 (O_4796,N_48156,N_47507);
xnor UO_4797 (O_4797,N_46622,N_49583);
nand UO_4798 (O_4798,N_49084,N_45431);
and UO_4799 (O_4799,N_48104,N_49553);
nor UO_4800 (O_4800,N_48497,N_46890);
and UO_4801 (O_4801,N_46890,N_46103);
nand UO_4802 (O_4802,N_45415,N_49259);
nand UO_4803 (O_4803,N_49958,N_49321);
nor UO_4804 (O_4804,N_45078,N_46505);
xnor UO_4805 (O_4805,N_49110,N_46207);
or UO_4806 (O_4806,N_46437,N_45472);
nor UO_4807 (O_4807,N_47690,N_49412);
nor UO_4808 (O_4808,N_47993,N_49841);
or UO_4809 (O_4809,N_48371,N_46790);
and UO_4810 (O_4810,N_45858,N_46929);
nand UO_4811 (O_4811,N_48047,N_48645);
or UO_4812 (O_4812,N_48203,N_49886);
xor UO_4813 (O_4813,N_49215,N_49557);
nand UO_4814 (O_4814,N_47821,N_45485);
and UO_4815 (O_4815,N_47198,N_46887);
nand UO_4816 (O_4816,N_49579,N_46054);
nand UO_4817 (O_4817,N_47659,N_45640);
nand UO_4818 (O_4818,N_47610,N_48656);
and UO_4819 (O_4819,N_45258,N_46772);
xnor UO_4820 (O_4820,N_48263,N_49139);
nand UO_4821 (O_4821,N_48662,N_45324);
or UO_4822 (O_4822,N_46491,N_49701);
or UO_4823 (O_4823,N_49586,N_48322);
xor UO_4824 (O_4824,N_46446,N_45316);
or UO_4825 (O_4825,N_45166,N_49271);
xnor UO_4826 (O_4826,N_46538,N_49104);
nand UO_4827 (O_4827,N_48444,N_46765);
and UO_4828 (O_4828,N_48607,N_45865);
nand UO_4829 (O_4829,N_45257,N_48525);
nor UO_4830 (O_4830,N_48381,N_47050);
and UO_4831 (O_4831,N_45489,N_49488);
xor UO_4832 (O_4832,N_49025,N_49104);
or UO_4833 (O_4833,N_47260,N_49192);
or UO_4834 (O_4834,N_47252,N_45958);
and UO_4835 (O_4835,N_46037,N_47693);
and UO_4836 (O_4836,N_45788,N_49770);
xnor UO_4837 (O_4837,N_47788,N_46694);
nor UO_4838 (O_4838,N_49520,N_47332);
nor UO_4839 (O_4839,N_49449,N_45362);
xnor UO_4840 (O_4840,N_47058,N_45300);
nor UO_4841 (O_4841,N_49351,N_49898);
nand UO_4842 (O_4842,N_49400,N_47458);
and UO_4843 (O_4843,N_49855,N_45131);
or UO_4844 (O_4844,N_46874,N_47690);
or UO_4845 (O_4845,N_45767,N_49919);
or UO_4846 (O_4846,N_46583,N_49415);
nand UO_4847 (O_4847,N_49032,N_47980);
xor UO_4848 (O_4848,N_48982,N_49616);
xor UO_4849 (O_4849,N_47078,N_45425);
and UO_4850 (O_4850,N_45671,N_48533);
nand UO_4851 (O_4851,N_45161,N_49213);
nand UO_4852 (O_4852,N_47207,N_46759);
and UO_4853 (O_4853,N_48351,N_46533);
xor UO_4854 (O_4854,N_46937,N_48517);
nor UO_4855 (O_4855,N_48507,N_45521);
nor UO_4856 (O_4856,N_49804,N_49046);
xnor UO_4857 (O_4857,N_47784,N_45697);
nor UO_4858 (O_4858,N_46423,N_46283);
nand UO_4859 (O_4859,N_45132,N_46268);
nor UO_4860 (O_4860,N_47171,N_46582);
nand UO_4861 (O_4861,N_45673,N_49541);
xor UO_4862 (O_4862,N_48325,N_46075);
and UO_4863 (O_4863,N_47371,N_48653);
or UO_4864 (O_4864,N_45912,N_46071);
nand UO_4865 (O_4865,N_46779,N_45137);
xor UO_4866 (O_4866,N_45203,N_47918);
nand UO_4867 (O_4867,N_47512,N_45465);
and UO_4868 (O_4868,N_46657,N_48696);
and UO_4869 (O_4869,N_49462,N_47237);
xnor UO_4870 (O_4870,N_48881,N_49859);
nand UO_4871 (O_4871,N_49586,N_46066);
and UO_4872 (O_4872,N_46057,N_45458);
or UO_4873 (O_4873,N_49153,N_48831);
and UO_4874 (O_4874,N_49501,N_45442);
xor UO_4875 (O_4875,N_47395,N_46589);
and UO_4876 (O_4876,N_49308,N_47502);
nor UO_4877 (O_4877,N_45752,N_49129);
and UO_4878 (O_4878,N_47770,N_45934);
and UO_4879 (O_4879,N_48988,N_47961);
xor UO_4880 (O_4880,N_47705,N_45348);
nor UO_4881 (O_4881,N_47212,N_47673);
or UO_4882 (O_4882,N_49442,N_45065);
xor UO_4883 (O_4883,N_48002,N_46824);
or UO_4884 (O_4884,N_49237,N_48240);
and UO_4885 (O_4885,N_45654,N_47949);
or UO_4886 (O_4886,N_47528,N_48527);
xnor UO_4887 (O_4887,N_46992,N_46581);
or UO_4888 (O_4888,N_48768,N_45429);
nand UO_4889 (O_4889,N_49536,N_48904);
nor UO_4890 (O_4890,N_47021,N_45676);
and UO_4891 (O_4891,N_48870,N_46655);
and UO_4892 (O_4892,N_47209,N_45707);
xnor UO_4893 (O_4893,N_45297,N_47399);
nand UO_4894 (O_4894,N_47431,N_47662);
xnor UO_4895 (O_4895,N_46763,N_49928);
or UO_4896 (O_4896,N_46206,N_49272);
xor UO_4897 (O_4897,N_45577,N_48307);
xor UO_4898 (O_4898,N_48374,N_47746);
or UO_4899 (O_4899,N_47124,N_48892);
or UO_4900 (O_4900,N_49549,N_47317);
nor UO_4901 (O_4901,N_49583,N_48434);
nor UO_4902 (O_4902,N_45077,N_46168);
or UO_4903 (O_4903,N_48763,N_47557);
xnor UO_4904 (O_4904,N_45079,N_45235);
nor UO_4905 (O_4905,N_47047,N_48002);
xor UO_4906 (O_4906,N_48309,N_46116);
nand UO_4907 (O_4907,N_47939,N_46585);
or UO_4908 (O_4908,N_48778,N_47767);
xor UO_4909 (O_4909,N_47247,N_47677);
nor UO_4910 (O_4910,N_45548,N_48228);
xnor UO_4911 (O_4911,N_48818,N_45556);
or UO_4912 (O_4912,N_45360,N_45039);
xor UO_4913 (O_4913,N_48952,N_45306);
nor UO_4914 (O_4914,N_49011,N_49797);
or UO_4915 (O_4915,N_47139,N_46815);
or UO_4916 (O_4916,N_49732,N_46497);
and UO_4917 (O_4917,N_45208,N_46363);
or UO_4918 (O_4918,N_49327,N_47326);
nand UO_4919 (O_4919,N_48152,N_48525);
nand UO_4920 (O_4920,N_47261,N_49744);
and UO_4921 (O_4921,N_46257,N_46262);
nand UO_4922 (O_4922,N_48081,N_46341);
nand UO_4923 (O_4923,N_45299,N_46034);
or UO_4924 (O_4924,N_49787,N_47680);
or UO_4925 (O_4925,N_47030,N_49552);
nand UO_4926 (O_4926,N_46402,N_45011);
nand UO_4927 (O_4927,N_47058,N_49170);
and UO_4928 (O_4928,N_49215,N_48961);
or UO_4929 (O_4929,N_49120,N_46034);
nor UO_4930 (O_4930,N_49366,N_45254);
xnor UO_4931 (O_4931,N_46660,N_46843);
nand UO_4932 (O_4932,N_46361,N_49150);
xnor UO_4933 (O_4933,N_48223,N_46746);
or UO_4934 (O_4934,N_45052,N_46605);
nor UO_4935 (O_4935,N_46208,N_48081);
and UO_4936 (O_4936,N_46226,N_46720);
nor UO_4937 (O_4937,N_45400,N_45430);
xor UO_4938 (O_4938,N_46549,N_47781);
nand UO_4939 (O_4939,N_48172,N_45525);
xnor UO_4940 (O_4940,N_46418,N_47996);
xor UO_4941 (O_4941,N_49324,N_47701);
nand UO_4942 (O_4942,N_47809,N_49401);
or UO_4943 (O_4943,N_48675,N_45774);
nor UO_4944 (O_4944,N_48877,N_48028);
xor UO_4945 (O_4945,N_46810,N_48879);
and UO_4946 (O_4946,N_46845,N_45255);
or UO_4947 (O_4947,N_47982,N_45525);
nand UO_4948 (O_4948,N_46711,N_45711);
xor UO_4949 (O_4949,N_45338,N_49461);
xnor UO_4950 (O_4950,N_47766,N_49047);
xor UO_4951 (O_4951,N_47767,N_46507);
xnor UO_4952 (O_4952,N_45972,N_48243);
or UO_4953 (O_4953,N_48530,N_48981);
and UO_4954 (O_4954,N_47807,N_46418);
nand UO_4955 (O_4955,N_45106,N_46926);
or UO_4956 (O_4956,N_46323,N_49870);
xor UO_4957 (O_4957,N_49870,N_45894);
xnor UO_4958 (O_4958,N_48766,N_48276);
xor UO_4959 (O_4959,N_45687,N_48745);
nor UO_4960 (O_4960,N_49358,N_47034);
or UO_4961 (O_4961,N_47564,N_48369);
xnor UO_4962 (O_4962,N_45991,N_46567);
nor UO_4963 (O_4963,N_48171,N_46993);
and UO_4964 (O_4964,N_48774,N_48300);
nand UO_4965 (O_4965,N_46214,N_49635);
and UO_4966 (O_4966,N_45295,N_49585);
or UO_4967 (O_4967,N_45331,N_45278);
or UO_4968 (O_4968,N_46303,N_45737);
nand UO_4969 (O_4969,N_47686,N_45046);
or UO_4970 (O_4970,N_47420,N_48464);
nand UO_4971 (O_4971,N_45990,N_46691);
or UO_4972 (O_4972,N_49778,N_49088);
nor UO_4973 (O_4973,N_46115,N_45771);
or UO_4974 (O_4974,N_48572,N_48068);
nand UO_4975 (O_4975,N_45597,N_47183);
nor UO_4976 (O_4976,N_49277,N_45421);
xnor UO_4977 (O_4977,N_46595,N_45711);
nand UO_4978 (O_4978,N_47166,N_49905);
xnor UO_4979 (O_4979,N_47672,N_45049);
xnor UO_4980 (O_4980,N_48407,N_46511);
nor UO_4981 (O_4981,N_49830,N_49479);
or UO_4982 (O_4982,N_47826,N_46687);
xor UO_4983 (O_4983,N_47849,N_49288);
nor UO_4984 (O_4984,N_47281,N_49399);
or UO_4985 (O_4985,N_49673,N_48636);
nor UO_4986 (O_4986,N_48558,N_47946);
or UO_4987 (O_4987,N_49923,N_46534);
or UO_4988 (O_4988,N_45193,N_49347);
nor UO_4989 (O_4989,N_46739,N_46064);
and UO_4990 (O_4990,N_47585,N_48991);
or UO_4991 (O_4991,N_47681,N_45485);
and UO_4992 (O_4992,N_48737,N_48829);
xor UO_4993 (O_4993,N_49456,N_48246);
xor UO_4994 (O_4994,N_45714,N_46756);
and UO_4995 (O_4995,N_46945,N_46206);
or UO_4996 (O_4996,N_49826,N_46431);
nand UO_4997 (O_4997,N_47174,N_49966);
nor UO_4998 (O_4998,N_47273,N_48629);
or UO_4999 (O_4999,N_47883,N_47211);
endmodule