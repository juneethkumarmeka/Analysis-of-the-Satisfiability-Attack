module basic_500_3000_500_4_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_26,In_128);
nand U1 (N_1,In_486,In_246);
and U2 (N_2,In_100,In_400);
or U3 (N_3,In_472,In_393);
or U4 (N_4,In_176,In_69);
nand U5 (N_5,In_76,In_271);
or U6 (N_6,In_249,In_291);
and U7 (N_7,In_195,In_52);
and U8 (N_8,In_413,In_315);
or U9 (N_9,In_442,In_468);
nor U10 (N_10,In_253,In_70);
or U11 (N_11,In_132,In_384);
or U12 (N_12,In_302,In_415);
nand U13 (N_13,In_106,In_337);
and U14 (N_14,In_117,In_165);
nand U15 (N_15,In_45,In_133);
and U16 (N_16,In_268,In_435);
nor U17 (N_17,In_462,In_159);
nor U18 (N_18,In_463,In_47);
nor U19 (N_19,In_467,In_104);
or U20 (N_20,In_43,In_200);
or U21 (N_21,In_428,In_382);
nor U22 (N_22,In_493,In_346);
or U23 (N_23,In_158,In_326);
and U24 (N_24,In_251,In_7);
or U25 (N_25,In_345,In_171);
or U26 (N_26,In_398,In_114);
or U27 (N_27,In_82,In_269);
and U28 (N_28,In_460,In_0);
nor U29 (N_29,In_180,In_239);
and U30 (N_30,In_138,In_207);
nor U31 (N_31,In_322,In_408);
nor U32 (N_32,In_116,In_371);
nand U33 (N_33,In_369,In_135);
nand U34 (N_34,In_381,In_110);
and U35 (N_35,In_277,In_81);
or U36 (N_36,In_388,In_163);
and U37 (N_37,In_262,In_314);
nand U38 (N_38,In_166,In_361);
nand U39 (N_39,In_57,In_49);
nor U40 (N_40,In_419,In_457);
and U41 (N_41,In_464,In_305);
and U42 (N_42,In_150,In_236);
or U43 (N_43,In_245,In_333);
or U44 (N_44,In_88,In_225);
nor U45 (N_45,In_340,In_375);
and U46 (N_46,In_372,In_102);
nor U47 (N_47,In_276,In_13);
or U48 (N_48,In_141,In_488);
or U49 (N_49,In_160,In_256);
and U50 (N_50,In_264,In_492);
and U51 (N_51,In_196,In_449);
nand U52 (N_52,In_29,In_53);
nor U53 (N_53,In_257,In_46);
or U54 (N_54,In_281,In_194);
and U55 (N_55,In_235,In_212);
xor U56 (N_56,In_365,In_349);
or U57 (N_57,In_494,In_332);
or U58 (N_58,In_1,In_229);
nand U59 (N_59,In_55,In_499);
nand U60 (N_60,In_204,In_108);
nor U61 (N_61,In_175,In_323);
nor U62 (N_62,In_164,In_273);
nand U63 (N_63,In_260,In_111);
or U64 (N_64,In_320,In_185);
or U65 (N_65,In_161,In_206);
and U66 (N_66,In_448,In_339);
or U67 (N_67,In_199,In_351);
nor U68 (N_68,In_367,In_137);
or U69 (N_69,In_490,In_99);
and U70 (N_70,In_437,In_401);
or U71 (N_71,In_122,In_342);
nor U72 (N_72,In_168,In_495);
nor U73 (N_73,In_385,In_412);
nor U74 (N_74,In_211,In_170);
or U75 (N_75,In_218,In_41);
and U76 (N_76,In_197,In_37);
nand U77 (N_77,In_485,In_379);
nor U78 (N_78,In_131,In_444);
or U79 (N_79,In_290,In_316);
xnor U80 (N_80,In_354,In_22);
and U81 (N_81,In_68,In_360);
or U82 (N_82,In_98,In_250);
or U83 (N_83,In_350,In_344);
or U84 (N_84,In_425,In_397);
nor U85 (N_85,In_429,In_42);
nor U86 (N_86,In_152,In_147);
or U87 (N_87,In_34,In_31);
nand U88 (N_88,In_16,In_282);
nand U89 (N_89,In_312,In_383);
and U90 (N_90,In_307,In_358);
or U91 (N_91,In_456,In_478);
nand U92 (N_92,In_258,In_112);
nor U93 (N_93,In_248,In_470);
nor U94 (N_94,In_423,In_453);
and U95 (N_95,In_411,In_418);
or U96 (N_96,In_134,In_420);
or U97 (N_97,In_479,In_489);
nand U98 (N_98,In_189,In_21);
and U99 (N_99,In_123,In_107);
nand U100 (N_100,In_178,In_473);
nor U101 (N_101,In_275,In_343);
nand U102 (N_102,In_461,In_85);
or U103 (N_103,In_145,In_390);
nand U104 (N_104,In_399,In_433);
and U105 (N_105,In_482,In_474);
nand U106 (N_106,In_172,In_455);
or U107 (N_107,In_94,In_301);
nand U108 (N_108,In_77,In_409);
or U109 (N_109,In_353,In_202);
or U110 (N_110,In_18,In_79);
nor U111 (N_111,In_402,In_267);
nor U112 (N_112,In_363,In_190);
xnor U113 (N_113,In_186,In_40);
nor U114 (N_114,In_115,In_450);
nor U115 (N_115,In_292,In_51);
or U116 (N_116,In_296,In_237);
nor U117 (N_117,In_24,In_265);
or U118 (N_118,In_173,In_498);
and U119 (N_119,In_432,In_373);
or U120 (N_120,In_311,In_148);
and U121 (N_121,In_255,In_87);
or U122 (N_122,In_272,In_174);
or U123 (N_123,In_215,In_93);
nand U124 (N_124,In_86,In_366);
nor U125 (N_125,In_146,In_233);
nand U126 (N_126,In_427,In_438);
nand U127 (N_127,In_223,In_56);
or U128 (N_128,In_244,In_459);
nor U129 (N_129,In_72,In_232);
nand U130 (N_130,In_434,In_193);
or U131 (N_131,In_188,In_226);
nand U132 (N_132,In_240,In_210);
nor U133 (N_133,In_405,In_20);
or U134 (N_134,In_64,In_286);
xor U135 (N_135,In_480,In_19);
or U136 (N_136,In_392,In_497);
nand U137 (N_137,In_395,In_252);
or U138 (N_138,In_295,In_4);
nand U139 (N_139,In_357,In_387);
and U140 (N_140,In_410,In_201);
and U141 (N_141,In_203,In_347);
and U142 (N_142,In_451,In_9);
nand U143 (N_143,In_3,In_317);
or U144 (N_144,In_118,In_130);
or U145 (N_145,In_139,In_91);
nor U146 (N_146,In_11,In_12);
nor U147 (N_147,In_297,In_289);
nand U148 (N_148,In_105,In_441);
nor U149 (N_149,In_270,In_169);
and U150 (N_150,In_280,In_213);
or U151 (N_151,In_220,In_153);
nor U152 (N_152,In_162,In_352);
nor U153 (N_153,In_319,In_140);
nand U154 (N_154,In_380,In_209);
and U155 (N_155,In_370,In_101);
nand U156 (N_156,In_294,In_143);
nor U157 (N_157,In_127,In_234);
nand U158 (N_158,In_238,In_376);
and U159 (N_159,In_65,In_466);
nand U160 (N_160,In_121,In_491);
and U161 (N_161,In_436,In_25);
xor U162 (N_162,In_288,In_334);
and U163 (N_163,In_414,In_216);
nor U164 (N_164,In_327,In_309);
nor U165 (N_165,In_192,In_299);
nor U166 (N_166,In_446,In_476);
nand U167 (N_167,In_440,In_62);
and U168 (N_168,In_109,In_330);
nand U169 (N_169,In_120,In_136);
nand U170 (N_170,In_404,In_391);
or U171 (N_171,In_119,In_205);
nor U172 (N_172,In_483,In_407);
nor U173 (N_173,In_228,In_27);
or U174 (N_174,In_80,In_247);
nor U175 (N_175,In_241,In_181);
and U176 (N_176,In_426,In_208);
or U177 (N_177,In_95,In_274);
nor U178 (N_178,In_30,In_191);
nor U179 (N_179,In_126,In_59);
nand U180 (N_180,In_298,In_33);
and U181 (N_181,In_443,In_187);
or U182 (N_182,In_156,In_39);
and U183 (N_183,In_454,In_61);
nand U184 (N_184,In_458,In_417);
or U185 (N_185,In_324,In_155);
nor U186 (N_186,In_355,In_32);
or U187 (N_187,In_430,In_48);
and U188 (N_188,In_475,In_89);
and U189 (N_189,In_230,In_28);
or U190 (N_190,In_304,In_278);
xnor U191 (N_191,In_154,In_124);
xor U192 (N_192,In_67,In_8);
or U193 (N_193,In_328,In_243);
nor U194 (N_194,In_129,In_359);
or U195 (N_195,In_329,In_125);
and U196 (N_196,In_151,In_184);
xnor U197 (N_197,In_58,In_331);
or U198 (N_198,In_263,In_284);
nand U199 (N_199,In_325,In_63);
and U200 (N_200,In_335,In_266);
and U201 (N_201,In_66,In_487);
or U202 (N_202,In_54,In_318);
and U203 (N_203,In_283,In_157);
nor U204 (N_204,In_313,In_224);
nand U205 (N_205,In_445,In_465);
or U206 (N_206,In_217,In_341);
and U207 (N_207,In_90,In_481);
nand U208 (N_208,In_424,In_219);
or U209 (N_209,In_396,In_50);
nand U210 (N_210,In_389,In_103);
nor U211 (N_211,In_73,In_259);
nor U212 (N_212,In_394,In_377);
and U213 (N_213,In_84,In_338);
and U214 (N_214,In_416,In_386);
and U215 (N_215,In_421,In_2);
and U216 (N_216,In_97,In_71);
and U217 (N_217,In_368,In_293);
or U218 (N_218,In_198,In_287);
or U219 (N_219,In_183,In_306);
nor U220 (N_220,In_78,In_452);
xnor U221 (N_221,In_231,In_348);
nor U222 (N_222,In_374,In_14);
or U223 (N_223,In_310,In_261);
or U224 (N_224,In_179,In_364);
or U225 (N_225,In_92,In_17);
or U226 (N_226,In_113,In_221);
nor U227 (N_227,In_321,In_144);
nand U228 (N_228,In_469,In_96);
nor U229 (N_229,In_177,In_285);
or U230 (N_230,In_142,In_378);
nor U231 (N_231,In_83,In_422);
nor U232 (N_232,In_471,In_403);
nand U233 (N_233,In_484,In_356);
nor U234 (N_234,In_477,In_15);
or U235 (N_235,In_496,In_439);
and U236 (N_236,In_44,In_38);
or U237 (N_237,In_222,In_447);
nor U238 (N_238,In_35,In_214);
and U239 (N_239,In_303,In_149);
or U240 (N_240,In_242,In_6);
or U241 (N_241,In_431,In_36);
nor U242 (N_242,In_60,In_5);
and U243 (N_243,In_182,In_362);
nand U244 (N_244,In_406,In_308);
nor U245 (N_245,In_300,In_74);
nand U246 (N_246,In_10,In_279);
nand U247 (N_247,In_336,In_75);
or U248 (N_248,In_167,In_254);
nor U249 (N_249,In_227,In_23);
or U250 (N_250,In_5,In_69);
nand U251 (N_251,In_300,In_350);
or U252 (N_252,In_197,In_496);
and U253 (N_253,In_317,In_28);
and U254 (N_254,In_139,In_93);
nor U255 (N_255,In_225,In_212);
nor U256 (N_256,In_144,In_360);
and U257 (N_257,In_443,In_254);
and U258 (N_258,In_301,In_127);
nand U259 (N_259,In_369,In_355);
nor U260 (N_260,In_247,In_338);
or U261 (N_261,In_272,In_177);
and U262 (N_262,In_320,In_98);
xnor U263 (N_263,In_220,In_147);
or U264 (N_264,In_323,In_84);
nand U265 (N_265,In_370,In_497);
and U266 (N_266,In_235,In_40);
and U267 (N_267,In_308,In_81);
nor U268 (N_268,In_30,In_430);
nor U269 (N_269,In_60,In_311);
or U270 (N_270,In_202,In_214);
and U271 (N_271,In_289,In_114);
nand U272 (N_272,In_465,In_30);
and U273 (N_273,In_70,In_161);
nand U274 (N_274,In_452,In_14);
nand U275 (N_275,In_214,In_87);
nand U276 (N_276,In_455,In_162);
nor U277 (N_277,In_163,In_44);
nand U278 (N_278,In_426,In_488);
or U279 (N_279,In_176,In_47);
nand U280 (N_280,In_498,In_340);
nand U281 (N_281,In_256,In_114);
or U282 (N_282,In_441,In_136);
nand U283 (N_283,In_17,In_472);
and U284 (N_284,In_384,In_406);
nand U285 (N_285,In_159,In_157);
nor U286 (N_286,In_433,In_8);
or U287 (N_287,In_176,In_487);
nand U288 (N_288,In_28,In_412);
or U289 (N_289,In_353,In_177);
or U290 (N_290,In_458,In_444);
nor U291 (N_291,In_153,In_213);
or U292 (N_292,In_178,In_161);
nand U293 (N_293,In_452,In_409);
or U294 (N_294,In_13,In_0);
and U295 (N_295,In_404,In_17);
or U296 (N_296,In_112,In_208);
or U297 (N_297,In_61,In_336);
and U298 (N_298,In_362,In_415);
xnor U299 (N_299,In_265,In_105);
nor U300 (N_300,In_218,In_376);
xor U301 (N_301,In_457,In_431);
or U302 (N_302,In_428,In_199);
or U303 (N_303,In_139,In_131);
nand U304 (N_304,In_187,In_57);
nor U305 (N_305,In_378,In_364);
and U306 (N_306,In_41,In_339);
nand U307 (N_307,In_366,In_5);
and U308 (N_308,In_10,In_271);
nor U309 (N_309,In_215,In_192);
and U310 (N_310,In_459,In_13);
nor U311 (N_311,In_64,In_223);
nand U312 (N_312,In_135,In_54);
nor U313 (N_313,In_9,In_7);
nor U314 (N_314,In_387,In_247);
or U315 (N_315,In_7,In_374);
or U316 (N_316,In_381,In_38);
nor U317 (N_317,In_163,In_401);
and U318 (N_318,In_280,In_332);
nor U319 (N_319,In_211,In_387);
and U320 (N_320,In_415,In_105);
and U321 (N_321,In_87,In_139);
nand U322 (N_322,In_80,In_446);
nand U323 (N_323,In_324,In_466);
nand U324 (N_324,In_349,In_447);
and U325 (N_325,In_291,In_355);
and U326 (N_326,In_98,In_357);
or U327 (N_327,In_391,In_442);
or U328 (N_328,In_419,In_472);
or U329 (N_329,In_45,In_389);
or U330 (N_330,In_77,In_119);
and U331 (N_331,In_385,In_168);
or U332 (N_332,In_80,In_418);
nand U333 (N_333,In_403,In_481);
nor U334 (N_334,In_470,In_379);
nand U335 (N_335,In_385,In_237);
or U336 (N_336,In_93,In_105);
or U337 (N_337,In_126,In_447);
and U338 (N_338,In_228,In_358);
nand U339 (N_339,In_225,In_49);
nor U340 (N_340,In_375,In_155);
nand U341 (N_341,In_414,In_20);
and U342 (N_342,In_399,In_264);
and U343 (N_343,In_143,In_124);
nand U344 (N_344,In_260,In_110);
and U345 (N_345,In_332,In_226);
and U346 (N_346,In_23,In_68);
nand U347 (N_347,In_420,In_313);
or U348 (N_348,In_210,In_469);
xnor U349 (N_349,In_485,In_250);
nor U350 (N_350,In_390,In_228);
nand U351 (N_351,In_427,In_49);
nor U352 (N_352,In_373,In_168);
or U353 (N_353,In_373,In_26);
or U354 (N_354,In_98,In_97);
nor U355 (N_355,In_291,In_486);
nand U356 (N_356,In_250,In_112);
and U357 (N_357,In_466,In_253);
and U358 (N_358,In_112,In_162);
or U359 (N_359,In_402,In_182);
and U360 (N_360,In_170,In_493);
and U361 (N_361,In_136,In_306);
or U362 (N_362,In_396,In_453);
or U363 (N_363,In_477,In_445);
nand U364 (N_364,In_481,In_247);
and U365 (N_365,In_498,In_57);
nor U366 (N_366,In_87,In_237);
nand U367 (N_367,In_76,In_400);
and U368 (N_368,In_432,In_153);
nor U369 (N_369,In_285,In_315);
nor U370 (N_370,In_83,In_382);
nor U371 (N_371,In_443,In_266);
nand U372 (N_372,In_173,In_151);
or U373 (N_373,In_27,In_324);
nor U374 (N_374,In_407,In_369);
and U375 (N_375,In_171,In_232);
and U376 (N_376,In_445,In_370);
or U377 (N_377,In_205,In_462);
and U378 (N_378,In_195,In_324);
nand U379 (N_379,In_105,In_257);
or U380 (N_380,In_45,In_172);
nor U381 (N_381,In_141,In_230);
nor U382 (N_382,In_220,In_339);
or U383 (N_383,In_465,In_154);
nand U384 (N_384,In_67,In_233);
nand U385 (N_385,In_32,In_257);
nor U386 (N_386,In_433,In_378);
or U387 (N_387,In_16,In_201);
or U388 (N_388,In_259,In_228);
nand U389 (N_389,In_437,In_433);
nand U390 (N_390,In_10,In_22);
and U391 (N_391,In_320,In_458);
nand U392 (N_392,In_166,In_135);
nor U393 (N_393,In_123,In_179);
and U394 (N_394,In_409,In_282);
nor U395 (N_395,In_150,In_100);
nor U396 (N_396,In_307,In_335);
and U397 (N_397,In_489,In_86);
nor U398 (N_398,In_410,In_144);
nand U399 (N_399,In_388,In_351);
nand U400 (N_400,In_284,In_48);
and U401 (N_401,In_271,In_471);
or U402 (N_402,In_425,In_108);
and U403 (N_403,In_456,In_286);
or U404 (N_404,In_55,In_211);
nor U405 (N_405,In_298,In_123);
xnor U406 (N_406,In_336,In_482);
nand U407 (N_407,In_112,In_384);
nor U408 (N_408,In_485,In_62);
or U409 (N_409,In_293,In_412);
or U410 (N_410,In_345,In_433);
nor U411 (N_411,In_18,In_108);
or U412 (N_412,In_80,In_399);
and U413 (N_413,In_441,In_356);
and U414 (N_414,In_375,In_73);
nand U415 (N_415,In_440,In_241);
and U416 (N_416,In_105,In_181);
nand U417 (N_417,In_149,In_338);
nand U418 (N_418,In_400,In_373);
or U419 (N_419,In_296,In_397);
nor U420 (N_420,In_456,In_2);
and U421 (N_421,In_25,In_397);
nand U422 (N_422,In_359,In_109);
and U423 (N_423,In_116,In_78);
or U424 (N_424,In_405,In_88);
nand U425 (N_425,In_463,In_369);
nor U426 (N_426,In_236,In_422);
or U427 (N_427,In_57,In_350);
and U428 (N_428,In_118,In_497);
nor U429 (N_429,In_8,In_198);
or U430 (N_430,In_477,In_211);
and U431 (N_431,In_261,In_115);
and U432 (N_432,In_456,In_487);
and U433 (N_433,In_396,In_455);
xnor U434 (N_434,In_220,In_461);
nand U435 (N_435,In_76,In_455);
nor U436 (N_436,In_300,In_21);
nor U437 (N_437,In_367,In_161);
and U438 (N_438,In_242,In_204);
nand U439 (N_439,In_350,In_391);
and U440 (N_440,In_470,In_407);
and U441 (N_441,In_56,In_485);
and U442 (N_442,In_429,In_441);
and U443 (N_443,In_396,In_351);
nor U444 (N_444,In_194,In_315);
and U445 (N_445,In_50,In_128);
nor U446 (N_446,In_461,In_198);
and U447 (N_447,In_401,In_435);
or U448 (N_448,In_1,In_7);
nand U449 (N_449,In_226,In_196);
or U450 (N_450,In_287,In_197);
nor U451 (N_451,In_28,In_443);
or U452 (N_452,In_449,In_331);
or U453 (N_453,In_16,In_85);
or U454 (N_454,In_312,In_456);
nand U455 (N_455,In_403,In_445);
and U456 (N_456,In_386,In_460);
and U457 (N_457,In_399,In_232);
nand U458 (N_458,In_236,In_356);
nor U459 (N_459,In_357,In_257);
and U460 (N_460,In_174,In_456);
and U461 (N_461,In_205,In_319);
and U462 (N_462,In_38,In_110);
and U463 (N_463,In_94,In_484);
xor U464 (N_464,In_177,In_189);
and U465 (N_465,In_247,In_5);
nor U466 (N_466,In_33,In_171);
nand U467 (N_467,In_277,In_98);
nor U468 (N_468,In_94,In_355);
nor U469 (N_469,In_28,In_205);
nand U470 (N_470,In_19,In_390);
nor U471 (N_471,In_230,In_279);
and U472 (N_472,In_140,In_6);
or U473 (N_473,In_343,In_397);
nor U474 (N_474,In_206,In_407);
nand U475 (N_475,In_250,In_52);
and U476 (N_476,In_444,In_320);
and U477 (N_477,In_223,In_5);
and U478 (N_478,In_82,In_6);
or U479 (N_479,In_493,In_366);
nor U480 (N_480,In_420,In_7);
nor U481 (N_481,In_406,In_282);
nand U482 (N_482,In_471,In_125);
nor U483 (N_483,In_201,In_235);
nor U484 (N_484,In_126,In_133);
nand U485 (N_485,In_352,In_217);
nor U486 (N_486,In_108,In_220);
and U487 (N_487,In_421,In_30);
xor U488 (N_488,In_39,In_15);
nor U489 (N_489,In_253,In_469);
and U490 (N_490,In_204,In_441);
or U491 (N_491,In_108,In_433);
or U492 (N_492,In_129,In_183);
and U493 (N_493,In_354,In_240);
or U494 (N_494,In_43,In_78);
nand U495 (N_495,In_424,In_26);
or U496 (N_496,In_122,In_327);
nor U497 (N_497,In_336,In_277);
and U498 (N_498,In_23,In_287);
or U499 (N_499,In_158,In_205);
nor U500 (N_500,In_370,In_211);
nor U501 (N_501,In_306,In_384);
and U502 (N_502,In_221,In_93);
nor U503 (N_503,In_139,In_219);
xor U504 (N_504,In_266,In_192);
nand U505 (N_505,In_70,In_18);
nand U506 (N_506,In_28,In_455);
and U507 (N_507,In_374,In_153);
nor U508 (N_508,In_284,In_16);
xor U509 (N_509,In_373,In_474);
nand U510 (N_510,In_37,In_373);
nand U511 (N_511,In_458,In_428);
nor U512 (N_512,In_134,In_136);
nor U513 (N_513,In_450,In_386);
nor U514 (N_514,In_387,In_106);
or U515 (N_515,In_35,In_8);
or U516 (N_516,In_497,In_246);
nand U517 (N_517,In_374,In_410);
or U518 (N_518,In_48,In_132);
and U519 (N_519,In_463,In_290);
nand U520 (N_520,In_213,In_86);
or U521 (N_521,In_367,In_153);
and U522 (N_522,In_402,In_463);
or U523 (N_523,In_487,In_39);
nor U524 (N_524,In_450,In_214);
and U525 (N_525,In_207,In_298);
or U526 (N_526,In_116,In_437);
nand U527 (N_527,In_171,In_354);
or U528 (N_528,In_439,In_363);
and U529 (N_529,In_364,In_293);
and U530 (N_530,In_320,In_291);
nand U531 (N_531,In_419,In_465);
nand U532 (N_532,In_69,In_170);
or U533 (N_533,In_160,In_288);
and U534 (N_534,In_491,In_387);
nor U535 (N_535,In_0,In_359);
and U536 (N_536,In_221,In_42);
nand U537 (N_537,In_109,In_231);
nor U538 (N_538,In_349,In_384);
and U539 (N_539,In_330,In_310);
nand U540 (N_540,In_148,In_422);
or U541 (N_541,In_15,In_158);
or U542 (N_542,In_20,In_380);
xnor U543 (N_543,In_487,In_404);
or U544 (N_544,In_122,In_315);
or U545 (N_545,In_403,In_385);
xnor U546 (N_546,In_198,In_188);
or U547 (N_547,In_417,In_188);
or U548 (N_548,In_490,In_383);
and U549 (N_549,In_117,In_293);
or U550 (N_550,In_122,In_271);
xor U551 (N_551,In_134,In_21);
nor U552 (N_552,In_311,In_90);
and U553 (N_553,In_46,In_58);
and U554 (N_554,In_162,In_315);
or U555 (N_555,In_401,In_324);
and U556 (N_556,In_377,In_309);
nor U557 (N_557,In_249,In_460);
nand U558 (N_558,In_286,In_429);
nor U559 (N_559,In_46,In_366);
nand U560 (N_560,In_413,In_57);
or U561 (N_561,In_287,In_279);
or U562 (N_562,In_423,In_439);
nor U563 (N_563,In_27,In_248);
and U564 (N_564,In_281,In_476);
nand U565 (N_565,In_73,In_195);
and U566 (N_566,In_359,In_162);
nor U567 (N_567,In_425,In_211);
nand U568 (N_568,In_145,In_39);
and U569 (N_569,In_229,In_384);
xor U570 (N_570,In_173,In_257);
xor U571 (N_571,In_278,In_84);
or U572 (N_572,In_111,In_238);
and U573 (N_573,In_38,In_496);
nor U574 (N_574,In_221,In_300);
and U575 (N_575,In_253,In_398);
nand U576 (N_576,In_357,In_297);
xor U577 (N_577,In_98,In_243);
nand U578 (N_578,In_445,In_213);
nor U579 (N_579,In_241,In_6);
or U580 (N_580,In_410,In_352);
and U581 (N_581,In_440,In_232);
or U582 (N_582,In_164,In_73);
nor U583 (N_583,In_165,In_68);
or U584 (N_584,In_5,In_139);
or U585 (N_585,In_378,In_108);
nand U586 (N_586,In_70,In_202);
and U587 (N_587,In_352,In_494);
and U588 (N_588,In_326,In_121);
or U589 (N_589,In_498,In_490);
and U590 (N_590,In_361,In_308);
nor U591 (N_591,In_302,In_203);
nor U592 (N_592,In_134,In_301);
nor U593 (N_593,In_446,In_390);
nand U594 (N_594,In_477,In_158);
nand U595 (N_595,In_481,In_18);
and U596 (N_596,In_30,In_416);
and U597 (N_597,In_410,In_427);
xnor U598 (N_598,In_366,In_89);
and U599 (N_599,In_467,In_69);
nand U600 (N_600,In_266,In_184);
nand U601 (N_601,In_180,In_38);
nor U602 (N_602,In_341,In_194);
nand U603 (N_603,In_205,In_325);
nor U604 (N_604,In_352,In_114);
nand U605 (N_605,In_487,In_305);
nor U606 (N_606,In_225,In_324);
nor U607 (N_607,In_492,In_250);
or U608 (N_608,In_77,In_182);
xor U609 (N_609,In_177,In_301);
nand U610 (N_610,In_137,In_65);
or U611 (N_611,In_297,In_183);
nand U612 (N_612,In_33,In_135);
xnor U613 (N_613,In_139,In_372);
nor U614 (N_614,In_465,In_460);
nor U615 (N_615,In_228,In_185);
or U616 (N_616,In_119,In_236);
or U617 (N_617,In_449,In_41);
or U618 (N_618,In_315,In_135);
and U619 (N_619,In_437,In_287);
or U620 (N_620,In_162,In_54);
nor U621 (N_621,In_471,In_79);
and U622 (N_622,In_328,In_487);
nand U623 (N_623,In_210,In_170);
and U624 (N_624,In_166,In_37);
nor U625 (N_625,In_315,In_252);
nand U626 (N_626,In_73,In_127);
and U627 (N_627,In_196,In_130);
nor U628 (N_628,In_453,In_429);
and U629 (N_629,In_373,In_140);
nand U630 (N_630,In_497,In_323);
and U631 (N_631,In_254,In_245);
and U632 (N_632,In_187,In_435);
or U633 (N_633,In_462,In_385);
nand U634 (N_634,In_116,In_420);
nand U635 (N_635,In_486,In_435);
nand U636 (N_636,In_485,In_156);
or U637 (N_637,In_487,In_293);
or U638 (N_638,In_207,In_36);
and U639 (N_639,In_39,In_251);
nor U640 (N_640,In_327,In_286);
and U641 (N_641,In_240,In_496);
nor U642 (N_642,In_250,In_51);
and U643 (N_643,In_393,In_0);
nor U644 (N_644,In_433,In_69);
or U645 (N_645,In_392,In_481);
and U646 (N_646,In_471,In_142);
or U647 (N_647,In_321,In_34);
or U648 (N_648,In_421,In_113);
nand U649 (N_649,In_56,In_345);
or U650 (N_650,In_56,In_33);
and U651 (N_651,In_202,In_147);
nor U652 (N_652,In_164,In_199);
nor U653 (N_653,In_387,In_225);
nor U654 (N_654,In_402,In_289);
nand U655 (N_655,In_350,In_162);
and U656 (N_656,In_15,In_79);
and U657 (N_657,In_424,In_218);
nor U658 (N_658,In_406,In_352);
or U659 (N_659,In_90,In_436);
xor U660 (N_660,In_198,In_104);
xnor U661 (N_661,In_464,In_466);
or U662 (N_662,In_192,In_496);
or U663 (N_663,In_488,In_245);
and U664 (N_664,In_73,In_386);
and U665 (N_665,In_101,In_214);
and U666 (N_666,In_162,In_300);
and U667 (N_667,In_383,In_127);
or U668 (N_668,In_95,In_373);
or U669 (N_669,In_456,In_139);
nor U670 (N_670,In_41,In_442);
nand U671 (N_671,In_85,In_233);
nand U672 (N_672,In_5,In_343);
nand U673 (N_673,In_313,In_492);
or U674 (N_674,In_394,In_383);
and U675 (N_675,In_143,In_449);
nand U676 (N_676,In_467,In_87);
nand U677 (N_677,In_192,In_135);
and U678 (N_678,In_105,In_399);
xnor U679 (N_679,In_453,In_32);
or U680 (N_680,In_476,In_200);
and U681 (N_681,In_172,In_176);
or U682 (N_682,In_22,In_159);
and U683 (N_683,In_17,In_115);
nand U684 (N_684,In_110,In_496);
or U685 (N_685,In_245,In_28);
nand U686 (N_686,In_271,In_111);
nor U687 (N_687,In_168,In_84);
nand U688 (N_688,In_194,In_492);
nand U689 (N_689,In_37,In_322);
and U690 (N_690,In_170,In_232);
nand U691 (N_691,In_255,In_468);
nor U692 (N_692,In_380,In_438);
nor U693 (N_693,In_435,In_17);
nand U694 (N_694,In_12,In_64);
nand U695 (N_695,In_246,In_263);
or U696 (N_696,In_22,In_168);
nand U697 (N_697,In_127,In_149);
nand U698 (N_698,In_263,In_391);
nor U699 (N_699,In_92,In_424);
or U700 (N_700,In_390,In_238);
and U701 (N_701,In_494,In_172);
nor U702 (N_702,In_478,In_127);
nor U703 (N_703,In_59,In_456);
nor U704 (N_704,In_168,In_395);
or U705 (N_705,In_75,In_188);
nor U706 (N_706,In_337,In_111);
and U707 (N_707,In_356,In_286);
nand U708 (N_708,In_398,In_347);
or U709 (N_709,In_190,In_380);
or U710 (N_710,In_180,In_101);
nor U711 (N_711,In_398,In_223);
nand U712 (N_712,In_445,In_216);
or U713 (N_713,In_455,In_266);
nand U714 (N_714,In_448,In_61);
nand U715 (N_715,In_237,In_193);
nor U716 (N_716,In_210,In_493);
xnor U717 (N_717,In_183,In_71);
nand U718 (N_718,In_97,In_375);
nor U719 (N_719,In_231,In_474);
nand U720 (N_720,In_29,In_16);
nor U721 (N_721,In_140,In_52);
or U722 (N_722,In_392,In_43);
nor U723 (N_723,In_108,In_217);
nor U724 (N_724,In_222,In_176);
or U725 (N_725,In_281,In_54);
or U726 (N_726,In_194,In_56);
nand U727 (N_727,In_422,In_204);
and U728 (N_728,In_128,In_80);
or U729 (N_729,In_406,In_225);
nor U730 (N_730,In_255,In_78);
nand U731 (N_731,In_14,In_370);
nor U732 (N_732,In_95,In_5);
nor U733 (N_733,In_458,In_84);
and U734 (N_734,In_341,In_57);
or U735 (N_735,In_26,In_200);
or U736 (N_736,In_355,In_401);
and U737 (N_737,In_134,In_0);
nand U738 (N_738,In_24,In_65);
or U739 (N_739,In_141,In_472);
nand U740 (N_740,In_198,In_433);
nand U741 (N_741,In_320,In_356);
or U742 (N_742,In_4,In_421);
nor U743 (N_743,In_20,In_116);
and U744 (N_744,In_449,In_491);
nor U745 (N_745,In_299,In_20);
or U746 (N_746,In_157,In_385);
xor U747 (N_747,In_65,In_258);
nand U748 (N_748,In_424,In_498);
nor U749 (N_749,In_481,In_265);
nand U750 (N_750,N_51,N_110);
nor U751 (N_751,N_44,N_282);
nand U752 (N_752,N_156,N_731);
nor U753 (N_753,N_718,N_422);
and U754 (N_754,N_648,N_467);
nand U755 (N_755,N_745,N_186);
nand U756 (N_756,N_142,N_414);
nor U757 (N_757,N_598,N_637);
and U758 (N_758,N_443,N_602);
and U759 (N_759,N_178,N_650);
or U760 (N_760,N_504,N_742);
or U761 (N_761,N_542,N_558);
and U762 (N_762,N_644,N_366);
nand U763 (N_763,N_684,N_502);
and U764 (N_764,N_495,N_344);
or U765 (N_765,N_340,N_324);
or U766 (N_766,N_357,N_212);
xnor U767 (N_767,N_410,N_534);
or U768 (N_768,N_310,N_74);
or U769 (N_769,N_375,N_354);
nor U770 (N_770,N_226,N_79);
nand U771 (N_771,N_84,N_45);
nor U772 (N_772,N_332,N_436);
nand U773 (N_773,N_729,N_677);
or U774 (N_774,N_307,N_128);
or U775 (N_775,N_148,N_672);
nor U776 (N_776,N_540,N_36);
nand U777 (N_777,N_639,N_293);
and U778 (N_778,N_615,N_479);
nand U779 (N_779,N_336,N_359);
and U780 (N_780,N_596,N_185);
or U781 (N_781,N_601,N_23);
nor U782 (N_782,N_719,N_68);
nor U783 (N_783,N_261,N_193);
nor U784 (N_784,N_576,N_712);
and U785 (N_785,N_232,N_485);
nor U786 (N_786,N_591,N_651);
xor U787 (N_787,N_123,N_720);
nand U788 (N_788,N_508,N_646);
and U789 (N_789,N_64,N_420);
and U790 (N_790,N_56,N_722);
or U791 (N_791,N_364,N_413);
nand U792 (N_792,N_384,N_380);
and U793 (N_793,N_63,N_303);
and U794 (N_794,N_312,N_175);
xnor U795 (N_795,N_716,N_647);
nand U796 (N_796,N_626,N_333);
nor U797 (N_797,N_693,N_360);
and U798 (N_798,N_533,N_2);
nor U799 (N_799,N_329,N_9);
nor U800 (N_800,N_468,N_610);
nand U801 (N_801,N_0,N_683);
and U802 (N_802,N_179,N_377);
or U803 (N_803,N_92,N_283);
or U804 (N_804,N_196,N_445);
and U805 (N_805,N_545,N_539);
and U806 (N_806,N_448,N_21);
nand U807 (N_807,N_476,N_277);
and U808 (N_808,N_341,N_29);
or U809 (N_809,N_163,N_486);
and U810 (N_810,N_73,N_229);
nand U811 (N_811,N_515,N_511);
nor U812 (N_812,N_484,N_151);
nor U813 (N_813,N_386,N_519);
nor U814 (N_814,N_348,N_734);
or U815 (N_815,N_580,N_560);
and U816 (N_816,N_138,N_117);
nor U817 (N_817,N_318,N_292);
nor U818 (N_818,N_126,N_274);
or U819 (N_819,N_496,N_201);
and U820 (N_820,N_260,N_331);
nand U821 (N_821,N_500,N_416);
nand U822 (N_822,N_154,N_525);
nand U823 (N_823,N_408,N_40);
or U824 (N_824,N_81,N_262);
nand U825 (N_825,N_369,N_258);
nor U826 (N_826,N_425,N_412);
or U827 (N_827,N_586,N_714);
nor U828 (N_828,N_55,N_240);
nand U829 (N_829,N_191,N_707);
or U830 (N_830,N_670,N_505);
nand U831 (N_831,N_509,N_234);
nand U832 (N_832,N_593,N_271);
nor U833 (N_833,N_299,N_306);
nor U834 (N_834,N_571,N_118);
nand U835 (N_835,N_256,N_204);
or U836 (N_836,N_272,N_326);
nand U837 (N_837,N_673,N_434);
nand U838 (N_838,N_103,N_302);
and U839 (N_839,N_723,N_286);
xor U840 (N_840,N_327,N_739);
and U841 (N_841,N_451,N_218);
or U842 (N_842,N_624,N_101);
nor U843 (N_843,N_389,N_49);
nor U844 (N_844,N_182,N_219);
nor U845 (N_845,N_184,N_708);
or U846 (N_846,N_465,N_634);
and U847 (N_847,N_95,N_675);
nor U848 (N_848,N_150,N_619);
or U849 (N_849,N_135,N_664);
or U850 (N_850,N_529,N_442);
nand U851 (N_851,N_305,N_62);
nor U852 (N_852,N_304,N_400);
and U853 (N_853,N_605,N_630);
and U854 (N_854,N_402,N_134);
or U855 (N_855,N_544,N_613);
nand U856 (N_856,N_12,N_665);
nand U857 (N_857,N_518,N_347);
and U858 (N_858,N_112,N_311);
nor U859 (N_859,N_704,N_177);
nor U860 (N_860,N_97,N_245);
and U861 (N_861,N_512,N_301);
nor U862 (N_862,N_162,N_695);
and U863 (N_863,N_243,N_116);
and U864 (N_864,N_674,N_238);
nor U865 (N_865,N_317,N_463);
or U866 (N_866,N_440,N_659);
nand U867 (N_867,N_435,N_546);
nor U868 (N_868,N_82,N_633);
nor U869 (N_869,N_568,N_456);
and U870 (N_870,N_666,N_600);
nand U871 (N_871,N_146,N_67);
nor U872 (N_872,N_33,N_202);
nor U873 (N_873,N_614,N_257);
nor U874 (N_874,N_109,N_749);
and U875 (N_875,N_503,N_685);
nand U876 (N_876,N_144,N_160);
nand U877 (N_877,N_165,N_290);
and U878 (N_878,N_661,N_481);
nor U879 (N_879,N_566,N_527);
or U880 (N_880,N_432,N_501);
and U881 (N_881,N_641,N_345);
and U882 (N_882,N_556,N_78);
and U883 (N_883,N_526,N_567);
and U884 (N_884,N_421,N_444);
nand U885 (N_885,N_631,N_114);
and U886 (N_886,N_635,N_132);
and U887 (N_887,N_570,N_423);
nor U888 (N_888,N_220,N_174);
or U889 (N_889,N_622,N_342);
or U890 (N_890,N_139,N_363);
nand U891 (N_891,N_237,N_246);
xnor U892 (N_892,N_645,N_592);
nor U893 (N_893,N_741,N_668);
and U894 (N_894,N_25,N_288);
or U895 (N_895,N_57,N_550);
nand U896 (N_896,N_190,N_93);
or U897 (N_897,N_352,N_211);
or U898 (N_898,N_457,N_100);
nand U899 (N_899,N_141,N_689);
and U900 (N_900,N_740,N_300);
and U901 (N_901,N_39,N_16);
nand U902 (N_902,N_690,N_99);
nor U903 (N_903,N_725,N_35);
and U904 (N_904,N_129,N_607);
or U905 (N_905,N_627,N_70);
or U906 (N_906,N_210,N_53);
nand U907 (N_907,N_582,N_379);
nor U908 (N_908,N_250,N_143);
or U909 (N_909,N_266,N_309);
or U910 (N_910,N_548,N_276);
and U911 (N_911,N_430,N_662);
and U912 (N_912,N_398,N_325);
nor U913 (N_913,N_553,N_280);
or U914 (N_914,N_699,N_543);
nor U915 (N_915,N_642,N_239);
nand U916 (N_916,N_603,N_427);
or U917 (N_917,N_72,N_166);
or U918 (N_918,N_285,N_131);
nor U919 (N_919,N_252,N_13);
or U920 (N_920,N_322,N_48);
nor U921 (N_921,N_573,N_287);
nand U922 (N_922,N_381,N_321);
and U923 (N_923,N_58,N_632);
nand U924 (N_924,N_506,N_473);
nor U925 (N_925,N_471,N_371);
nand U926 (N_926,N_730,N_102);
or U927 (N_927,N_50,N_426);
or U928 (N_928,N_89,N_295);
or U929 (N_929,N_200,N_676);
nand U930 (N_930,N_735,N_450);
xor U931 (N_931,N_270,N_554);
and U932 (N_932,N_696,N_279);
and U933 (N_933,N_28,N_517);
and U934 (N_934,N_71,N_667);
nand U935 (N_935,N_358,N_663);
nand U936 (N_936,N_681,N_459);
nor U937 (N_937,N_194,N_120);
or U938 (N_938,N_638,N_584);
and U939 (N_939,N_26,N_628);
nor U940 (N_940,N_597,N_581);
nor U941 (N_941,N_374,N_176);
or U942 (N_942,N_335,N_487);
nor U943 (N_943,N_715,N_281);
nand U944 (N_944,N_611,N_536);
or U945 (N_945,N_604,N_572);
or U946 (N_946,N_406,N_215);
nand U947 (N_947,N_528,N_216);
nand U948 (N_948,N_587,N_30);
and U949 (N_949,N_296,N_706);
or U950 (N_950,N_217,N_15);
nor U951 (N_951,N_319,N_390);
nor U952 (N_952,N_315,N_122);
and U953 (N_953,N_617,N_688);
or U954 (N_954,N_253,N_458);
and U955 (N_955,N_140,N_475);
nor U956 (N_956,N_606,N_431);
and U957 (N_957,N_222,N_578);
nand U958 (N_958,N_743,N_589);
and U959 (N_959,N_181,N_199);
and U960 (N_960,N_531,N_124);
nand U961 (N_961,N_441,N_727);
and U962 (N_962,N_612,N_3);
or U963 (N_963,N_577,N_658);
and U964 (N_964,N_76,N_499);
or U965 (N_965,N_460,N_694);
or U966 (N_966,N_61,N_490);
nor U967 (N_967,N_653,N_152);
or U968 (N_968,N_541,N_255);
and U969 (N_969,N_744,N_549);
nor U970 (N_970,N_244,N_655);
nor U971 (N_971,N_405,N_565);
nor U972 (N_972,N_187,N_362);
or U973 (N_973,N_24,N_313);
and U974 (N_974,N_314,N_136);
or U975 (N_975,N_407,N_705);
xnor U976 (N_976,N_86,N_214);
or U977 (N_977,N_251,N_284);
nor U978 (N_978,N_488,N_370);
nor U979 (N_979,N_449,N_429);
nand U980 (N_980,N_455,N_209);
xor U981 (N_981,N_569,N_17);
nand U982 (N_982,N_157,N_119);
or U983 (N_983,N_47,N_483);
or U984 (N_984,N_497,N_328);
nand U985 (N_985,N_579,N_98);
nor U986 (N_986,N_158,N_230);
and U987 (N_987,N_361,N_149);
nand U988 (N_988,N_514,N_404);
nor U989 (N_989,N_588,N_249);
nand U990 (N_990,N_267,N_575);
nor U991 (N_991,N_552,N_530);
nand U992 (N_992,N_520,N_713);
nor U993 (N_993,N_88,N_654);
nor U994 (N_994,N_547,N_248);
and U995 (N_995,N_583,N_590);
and U996 (N_996,N_339,N_298);
or U997 (N_997,N_669,N_428);
nor U998 (N_998,N_372,N_107);
or U999 (N_999,N_438,N_608);
nor U1000 (N_1000,N_738,N_656);
nor U1001 (N_1001,N_409,N_643);
and U1002 (N_1002,N_660,N_223);
nand U1003 (N_1003,N_137,N_297);
nor U1004 (N_1004,N_563,N_167);
or U1005 (N_1005,N_717,N_636);
nor U1006 (N_1006,N_424,N_640);
or U1007 (N_1007,N_382,N_197);
nor U1008 (N_1008,N_491,N_417);
or U1009 (N_1009,N_269,N_1);
and U1010 (N_1010,N_105,N_564);
or U1011 (N_1011,N_77,N_153);
or U1012 (N_1012,N_687,N_206);
nand U1013 (N_1013,N_41,N_649);
and U1014 (N_1014,N_701,N_351);
nand U1015 (N_1015,N_555,N_316);
nor U1016 (N_1016,N_106,N_145);
and U1017 (N_1017,N_671,N_164);
nand U1018 (N_1018,N_10,N_625);
nor U1019 (N_1019,N_353,N_87);
nor U1020 (N_1020,N_396,N_559);
nor U1021 (N_1021,N_337,N_170);
nand U1022 (N_1022,N_205,N_65);
xnor U1023 (N_1023,N_748,N_395);
nand U1024 (N_1024,N_397,N_213);
and U1025 (N_1025,N_383,N_171);
nor U1026 (N_1026,N_391,N_494);
or U1027 (N_1027,N_482,N_121);
and U1028 (N_1028,N_513,N_94);
and U1029 (N_1029,N_721,N_378);
or U1030 (N_1030,N_388,N_42);
nor U1031 (N_1031,N_59,N_724);
or U1032 (N_1032,N_228,N_493);
and U1033 (N_1033,N_532,N_259);
and U1034 (N_1034,N_192,N_510);
nor U1035 (N_1035,N_437,N_733);
nor U1036 (N_1036,N_155,N_236);
or U1037 (N_1037,N_657,N_399);
and U1038 (N_1038,N_629,N_368);
or U1039 (N_1039,N_189,N_320);
nand U1040 (N_1040,N_537,N_330);
nor U1041 (N_1041,N_574,N_221);
and U1042 (N_1042,N_195,N_20);
nor U1043 (N_1043,N_133,N_447);
nor U1044 (N_1044,N_14,N_710);
nand U1045 (N_1045,N_172,N_711);
or U1046 (N_1046,N_367,N_609);
nor U1047 (N_1047,N_401,N_235);
or U1048 (N_1048,N_478,N_679);
nor U1049 (N_1049,N_551,N_454);
nand U1050 (N_1050,N_180,N_680);
or U1051 (N_1051,N_538,N_470);
nand U1052 (N_1052,N_96,N_11);
nor U1053 (N_1053,N_60,N_4);
nor U1054 (N_1054,N_461,N_108);
nand U1055 (N_1055,N_241,N_376);
and U1056 (N_1056,N_746,N_585);
xnor U1057 (N_1057,N_173,N_231);
and U1058 (N_1058,N_535,N_480);
or U1059 (N_1059,N_32,N_85);
and U1060 (N_1060,N_356,N_621);
nand U1061 (N_1061,N_198,N_737);
or U1062 (N_1062,N_466,N_678);
and U1063 (N_1063,N_43,N_373);
nand U1064 (N_1064,N_161,N_524);
nor U1065 (N_1065,N_91,N_446);
nand U1066 (N_1066,N_323,N_385);
or U1067 (N_1067,N_66,N_709);
nand U1068 (N_1068,N_355,N_159);
and U1069 (N_1069,N_294,N_620);
or U1070 (N_1070,N_308,N_265);
nand U1071 (N_1071,N_523,N_130);
or U1072 (N_1072,N_365,N_268);
nand U1073 (N_1073,N_90,N_702);
nand U1074 (N_1074,N_522,N_599);
or U1075 (N_1075,N_289,N_732);
or U1076 (N_1076,N_27,N_264);
nor U1077 (N_1077,N_224,N_477);
or U1078 (N_1078,N_557,N_52);
nor U1079 (N_1079,N_462,N_747);
and U1080 (N_1080,N_225,N_127);
or U1081 (N_1081,N_169,N_698);
and U1082 (N_1082,N_18,N_334);
and U1083 (N_1083,N_692,N_394);
nor U1084 (N_1084,N_691,N_291);
nand U1085 (N_1085,N_623,N_54);
or U1086 (N_1086,N_498,N_492);
nand U1087 (N_1087,N_387,N_349);
and U1088 (N_1088,N_452,N_594);
nand U1089 (N_1089,N_273,N_38);
or U1090 (N_1090,N_111,N_343);
and U1091 (N_1091,N_227,N_168);
nand U1092 (N_1092,N_275,N_147);
and U1093 (N_1093,N_207,N_433);
nand U1094 (N_1094,N_697,N_415);
nand U1095 (N_1095,N_726,N_125);
nor U1096 (N_1096,N_8,N_7);
xor U1097 (N_1097,N_203,N_392);
nand U1098 (N_1098,N_46,N_188);
or U1099 (N_1099,N_682,N_507);
and U1100 (N_1100,N_263,N_472);
and U1101 (N_1101,N_115,N_19);
nand U1102 (N_1102,N_521,N_419);
or U1103 (N_1103,N_393,N_562);
or U1104 (N_1104,N_595,N_474);
nor U1105 (N_1105,N_104,N_22);
nand U1106 (N_1106,N_34,N_561);
nand U1107 (N_1107,N_703,N_686);
or U1108 (N_1108,N_464,N_736);
nor U1109 (N_1109,N_75,N_489);
and U1110 (N_1110,N_83,N_208);
or U1111 (N_1111,N_6,N_439);
nor U1112 (N_1112,N_652,N_411);
nor U1113 (N_1113,N_254,N_80);
nor U1114 (N_1114,N_338,N_37);
or U1115 (N_1115,N_618,N_346);
nor U1116 (N_1116,N_278,N_453);
nand U1117 (N_1117,N_728,N_616);
nor U1118 (N_1118,N_247,N_350);
nand U1119 (N_1119,N_5,N_469);
and U1120 (N_1120,N_418,N_69);
nor U1121 (N_1121,N_403,N_183);
and U1122 (N_1122,N_242,N_31);
and U1123 (N_1123,N_516,N_113);
and U1124 (N_1124,N_233,N_700);
or U1125 (N_1125,N_94,N_307);
xnor U1126 (N_1126,N_416,N_591);
nor U1127 (N_1127,N_354,N_314);
nor U1128 (N_1128,N_577,N_135);
and U1129 (N_1129,N_393,N_124);
nor U1130 (N_1130,N_703,N_70);
nand U1131 (N_1131,N_260,N_597);
nand U1132 (N_1132,N_388,N_744);
nor U1133 (N_1133,N_268,N_74);
or U1134 (N_1134,N_29,N_392);
or U1135 (N_1135,N_237,N_619);
nor U1136 (N_1136,N_382,N_81);
nand U1137 (N_1137,N_331,N_397);
and U1138 (N_1138,N_581,N_218);
or U1139 (N_1139,N_661,N_734);
and U1140 (N_1140,N_441,N_432);
or U1141 (N_1141,N_432,N_691);
or U1142 (N_1142,N_526,N_746);
nor U1143 (N_1143,N_507,N_625);
and U1144 (N_1144,N_365,N_332);
nor U1145 (N_1145,N_248,N_151);
nor U1146 (N_1146,N_730,N_362);
nand U1147 (N_1147,N_421,N_487);
nor U1148 (N_1148,N_474,N_463);
or U1149 (N_1149,N_717,N_504);
and U1150 (N_1150,N_174,N_0);
and U1151 (N_1151,N_126,N_406);
or U1152 (N_1152,N_178,N_161);
and U1153 (N_1153,N_129,N_216);
and U1154 (N_1154,N_416,N_142);
and U1155 (N_1155,N_354,N_149);
or U1156 (N_1156,N_600,N_607);
nand U1157 (N_1157,N_194,N_442);
or U1158 (N_1158,N_457,N_435);
nor U1159 (N_1159,N_211,N_35);
or U1160 (N_1160,N_224,N_168);
nor U1161 (N_1161,N_190,N_233);
nor U1162 (N_1162,N_296,N_574);
and U1163 (N_1163,N_572,N_83);
or U1164 (N_1164,N_516,N_302);
nor U1165 (N_1165,N_225,N_666);
nand U1166 (N_1166,N_192,N_462);
nand U1167 (N_1167,N_467,N_67);
and U1168 (N_1168,N_337,N_663);
nor U1169 (N_1169,N_462,N_396);
nand U1170 (N_1170,N_180,N_379);
nor U1171 (N_1171,N_500,N_234);
or U1172 (N_1172,N_506,N_574);
nor U1173 (N_1173,N_571,N_323);
and U1174 (N_1174,N_47,N_11);
nor U1175 (N_1175,N_459,N_325);
or U1176 (N_1176,N_527,N_451);
and U1177 (N_1177,N_513,N_666);
nand U1178 (N_1178,N_533,N_153);
nor U1179 (N_1179,N_502,N_399);
or U1180 (N_1180,N_529,N_480);
or U1181 (N_1181,N_268,N_515);
nand U1182 (N_1182,N_225,N_106);
nand U1183 (N_1183,N_28,N_584);
or U1184 (N_1184,N_476,N_669);
nand U1185 (N_1185,N_533,N_630);
xnor U1186 (N_1186,N_573,N_144);
nand U1187 (N_1187,N_373,N_78);
nor U1188 (N_1188,N_631,N_14);
nand U1189 (N_1189,N_266,N_108);
nor U1190 (N_1190,N_274,N_504);
nand U1191 (N_1191,N_224,N_27);
and U1192 (N_1192,N_600,N_689);
nor U1193 (N_1193,N_338,N_403);
or U1194 (N_1194,N_559,N_389);
nor U1195 (N_1195,N_249,N_742);
nor U1196 (N_1196,N_412,N_244);
nor U1197 (N_1197,N_621,N_359);
or U1198 (N_1198,N_116,N_654);
nand U1199 (N_1199,N_660,N_316);
and U1200 (N_1200,N_34,N_531);
or U1201 (N_1201,N_566,N_240);
or U1202 (N_1202,N_382,N_237);
nor U1203 (N_1203,N_485,N_42);
nand U1204 (N_1204,N_344,N_120);
and U1205 (N_1205,N_188,N_347);
nand U1206 (N_1206,N_687,N_489);
nor U1207 (N_1207,N_18,N_24);
nor U1208 (N_1208,N_375,N_48);
and U1209 (N_1209,N_3,N_282);
nand U1210 (N_1210,N_187,N_735);
or U1211 (N_1211,N_502,N_119);
nand U1212 (N_1212,N_206,N_741);
or U1213 (N_1213,N_148,N_430);
nand U1214 (N_1214,N_279,N_536);
and U1215 (N_1215,N_539,N_638);
and U1216 (N_1216,N_600,N_488);
or U1217 (N_1217,N_170,N_679);
or U1218 (N_1218,N_295,N_579);
and U1219 (N_1219,N_294,N_649);
and U1220 (N_1220,N_427,N_457);
and U1221 (N_1221,N_399,N_689);
nor U1222 (N_1222,N_345,N_529);
and U1223 (N_1223,N_593,N_517);
and U1224 (N_1224,N_78,N_522);
or U1225 (N_1225,N_622,N_715);
nand U1226 (N_1226,N_609,N_270);
nor U1227 (N_1227,N_168,N_610);
and U1228 (N_1228,N_79,N_668);
and U1229 (N_1229,N_73,N_381);
and U1230 (N_1230,N_430,N_77);
or U1231 (N_1231,N_476,N_282);
nor U1232 (N_1232,N_368,N_482);
nor U1233 (N_1233,N_92,N_561);
nor U1234 (N_1234,N_400,N_559);
nand U1235 (N_1235,N_749,N_10);
nor U1236 (N_1236,N_232,N_124);
or U1237 (N_1237,N_414,N_594);
nand U1238 (N_1238,N_113,N_419);
nor U1239 (N_1239,N_237,N_420);
nor U1240 (N_1240,N_244,N_261);
nand U1241 (N_1241,N_497,N_597);
or U1242 (N_1242,N_142,N_128);
and U1243 (N_1243,N_643,N_373);
nand U1244 (N_1244,N_35,N_668);
and U1245 (N_1245,N_225,N_24);
or U1246 (N_1246,N_667,N_459);
or U1247 (N_1247,N_464,N_149);
or U1248 (N_1248,N_549,N_706);
or U1249 (N_1249,N_688,N_33);
nand U1250 (N_1250,N_414,N_375);
and U1251 (N_1251,N_224,N_245);
and U1252 (N_1252,N_443,N_170);
or U1253 (N_1253,N_652,N_597);
nor U1254 (N_1254,N_163,N_323);
or U1255 (N_1255,N_743,N_308);
and U1256 (N_1256,N_258,N_598);
or U1257 (N_1257,N_503,N_321);
nand U1258 (N_1258,N_323,N_253);
nor U1259 (N_1259,N_45,N_324);
nor U1260 (N_1260,N_494,N_748);
nor U1261 (N_1261,N_409,N_730);
and U1262 (N_1262,N_572,N_694);
nand U1263 (N_1263,N_454,N_289);
and U1264 (N_1264,N_626,N_185);
nor U1265 (N_1265,N_319,N_1);
nand U1266 (N_1266,N_552,N_567);
nand U1267 (N_1267,N_388,N_566);
nor U1268 (N_1268,N_367,N_600);
nor U1269 (N_1269,N_732,N_158);
or U1270 (N_1270,N_210,N_545);
nand U1271 (N_1271,N_380,N_350);
or U1272 (N_1272,N_431,N_314);
nor U1273 (N_1273,N_330,N_572);
nor U1274 (N_1274,N_163,N_379);
nor U1275 (N_1275,N_420,N_623);
nor U1276 (N_1276,N_430,N_521);
xnor U1277 (N_1277,N_62,N_177);
or U1278 (N_1278,N_652,N_385);
and U1279 (N_1279,N_458,N_211);
and U1280 (N_1280,N_18,N_586);
xnor U1281 (N_1281,N_503,N_370);
nand U1282 (N_1282,N_700,N_27);
nor U1283 (N_1283,N_607,N_298);
or U1284 (N_1284,N_418,N_458);
nand U1285 (N_1285,N_31,N_16);
or U1286 (N_1286,N_492,N_529);
nand U1287 (N_1287,N_490,N_67);
nand U1288 (N_1288,N_657,N_105);
nor U1289 (N_1289,N_118,N_208);
or U1290 (N_1290,N_97,N_462);
nor U1291 (N_1291,N_208,N_613);
and U1292 (N_1292,N_483,N_508);
nor U1293 (N_1293,N_71,N_149);
nand U1294 (N_1294,N_497,N_219);
nand U1295 (N_1295,N_219,N_57);
nor U1296 (N_1296,N_333,N_631);
and U1297 (N_1297,N_547,N_486);
nand U1298 (N_1298,N_344,N_584);
and U1299 (N_1299,N_42,N_244);
xnor U1300 (N_1300,N_662,N_528);
nand U1301 (N_1301,N_183,N_575);
or U1302 (N_1302,N_116,N_80);
or U1303 (N_1303,N_497,N_691);
or U1304 (N_1304,N_474,N_710);
nand U1305 (N_1305,N_489,N_469);
and U1306 (N_1306,N_417,N_640);
or U1307 (N_1307,N_456,N_543);
nor U1308 (N_1308,N_660,N_635);
nor U1309 (N_1309,N_191,N_187);
nand U1310 (N_1310,N_589,N_407);
or U1311 (N_1311,N_365,N_677);
and U1312 (N_1312,N_282,N_562);
nor U1313 (N_1313,N_707,N_295);
and U1314 (N_1314,N_601,N_397);
and U1315 (N_1315,N_696,N_664);
nor U1316 (N_1316,N_699,N_315);
nor U1317 (N_1317,N_310,N_543);
or U1318 (N_1318,N_679,N_583);
or U1319 (N_1319,N_244,N_430);
nand U1320 (N_1320,N_222,N_64);
nand U1321 (N_1321,N_499,N_131);
and U1322 (N_1322,N_547,N_224);
xor U1323 (N_1323,N_737,N_189);
nor U1324 (N_1324,N_70,N_572);
nand U1325 (N_1325,N_631,N_369);
nand U1326 (N_1326,N_463,N_402);
or U1327 (N_1327,N_252,N_158);
and U1328 (N_1328,N_132,N_383);
and U1329 (N_1329,N_226,N_20);
nor U1330 (N_1330,N_221,N_638);
nand U1331 (N_1331,N_538,N_510);
nor U1332 (N_1332,N_192,N_274);
nand U1333 (N_1333,N_419,N_445);
nor U1334 (N_1334,N_354,N_388);
or U1335 (N_1335,N_356,N_724);
or U1336 (N_1336,N_227,N_86);
nand U1337 (N_1337,N_350,N_457);
nand U1338 (N_1338,N_126,N_78);
or U1339 (N_1339,N_229,N_176);
nor U1340 (N_1340,N_270,N_480);
nor U1341 (N_1341,N_301,N_42);
nand U1342 (N_1342,N_422,N_63);
xnor U1343 (N_1343,N_431,N_427);
and U1344 (N_1344,N_38,N_570);
nor U1345 (N_1345,N_441,N_123);
nand U1346 (N_1346,N_382,N_379);
and U1347 (N_1347,N_645,N_272);
nand U1348 (N_1348,N_565,N_415);
or U1349 (N_1349,N_598,N_38);
nor U1350 (N_1350,N_100,N_566);
nor U1351 (N_1351,N_496,N_477);
nor U1352 (N_1352,N_351,N_419);
xor U1353 (N_1353,N_89,N_32);
nor U1354 (N_1354,N_75,N_132);
nor U1355 (N_1355,N_436,N_378);
or U1356 (N_1356,N_696,N_156);
nor U1357 (N_1357,N_597,N_481);
or U1358 (N_1358,N_686,N_185);
and U1359 (N_1359,N_475,N_71);
or U1360 (N_1360,N_220,N_360);
or U1361 (N_1361,N_232,N_652);
and U1362 (N_1362,N_319,N_7);
nand U1363 (N_1363,N_23,N_494);
or U1364 (N_1364,N_369,N_189);
nor U1365 (N_1365,N_136,N_429);
nand U1366 (N_1366,N_60,N_344);
xor U1367 (N_1367,N_711,N_570);
nor U1368 (N_1368,N_83,N_213);
nor U1369 (N_1369,N_596,N_151);
or U1370 (N_1370,N_701,N_252);
or U1371 (N_1371,N_120,N_418);
nand U1372 (N_1372,N_107,N_393);
nand U1373 (N_1373,N_601,N_251);
nand U1374 (N_1374,N_694,N_714);
xnor U1375 (N_1375,N_4,N_63);
nand U1376 (N_1376,N_680,N_125);
and U1377 (N_1377,N_172,N_261);
nor U1378 (N_1378,N_372,N_447);
nor U1379 (N_1379,N_631,N_351);
and U1380 (N_1380,N_11,N_614);
and U1381 (N_1381,N_505,N_238);
or U1382 (N_1382,N_178,N_198);
and U1383 (N_1383,N_308,N_89);
and U1384 (N_1384,N_493,N_127);
nor U1385 (N_1385,N_630,N_731);
nand U1386 (N_1386,N_264,N_276);
nor U1387 (N_1387,N_675,N_641);
nor U1388 (N_1388,N_221,N_209);
or U1389 (N_1389,N_85,N_526);
nor U1390 (N_1390,N_234,N_3);
xnor U1391 (N_1391,N_261,N_680);
xor U1392 (N_1392,N_168,N_282);
and U1393 (N_1393,N_653,N_678);
and U1394 (N_1394,N_293,N_311);
or U1395 (N_1395,N_422,N_341);
nand U1396 (N_1396,N_623,N_126);
and U1397 (N_1397,N_729,N_70);
nand U1398 (N_1398,N_273,N_622);
or U1399 (N_1399,N_474,N_103);
nand U1400 (N_1400,N_671,N_577);
or U1401 (N_1401,N_359,N_571);
nor U1402 (N_1402,N_521,N_141);
nand U1403 (N_1403,N_214,N_588);
or U1404 (N_1404,N_674,N_213);
nor U1405 (N_1405,N_356,N_22);
nand U1406 (N_1406,N_708,N_644);
nor U1407 (N_1407,N_6,N_618);
nand U1408 (N_1408,N_3,N_360);
and U1409 (N_1409,N_452,N_98);
nand U1410 (N_1410,N_655,N_734);
and U1411 (N_1411,N_97,N_51);
or U1412 (N_1412,N_2,N_47);
and U1413 (N_1413,N_14,N_239);
nand U1414 (N_1414,N_257,N_599);
nand U1415 (N_1415,N_625,N_319);
or U1416 (N_1416,N_120,N_694);
or U1417 (N_1417,N_19,N_139);
nand U1418 (N_1418,N_285,N_609);
and U1419 (N_1419,N_226,N_132);
nor U1420 (N_1420,N_89,N_511);
or U1421 (N_1421,N_646,N_85);
nand U1422 (N_1422,N_679,N_97);
nand U1423 (N_1423,N_577,N_263);
xnor U1424 (N_1424,N_686,N_605);
and U1425 (N_1425,N_185,N_396);
and U1426 (N_1426,N_378,N_275);
and U1427 (N_1427,N_523,N_211);
nand U1428 (N_1428,N_39,N_749);
nor U1429 (N_1429,N_264,N_553);
nor U1430 (N_1430,N_372,N_99);
or U1431 (N_1431,N_694,N_61);
nand U1432 (N_1432,N_492,N_244);
nand U1433 (N_1433,N_572,N_613);
or U1434 (N_1434,N_350,N_647);
nor U1435 (N_1435,N_639,N_554);
nor U1436 (N_1436,N_731,N_705);
or U1437 (N_1437,N_54,N_605);
and U1438 (N_1438,N_458,N_563);
nand U1439 (N_1439,N_406,N_548);
and U1440 (N_1440,N_524,N_408);
nand U1441 (N_1441,N_242,N_234);
and U1442 (N_1442,N_715,N_212);
and U1443 (N_1443,N_37,N_716);
or U1444 (N_1444,N_343,N_664);
and U1445 (N_1445,N_132,N_46);
nor U1446 (N_1446,N_345,N_609);
nand U1447 (N_1447,N_159,N_24);
nor U1448 (N_1448,N_382,N_538);
nand U1449 (N_1449,N_318,N_200);
nand U1450 (N_1450,N_27,N_676);
and U1451 (N_1451,N_536,N_13);
nor U1452 (N_1452,N_265,N_242);
nand U1453 (N_1453,N_563,N_674);
nand U1454 (N_1454,N_479,N_387);
and U1455 (N_1455,N_459,N_394);
nand U1456 (N_1456,N_205,N_735);
nand U1457 (N_1457,N_671,N_677);
nand U1458 (N_1458,N_513,N_42);
nand U1459 (N_1459,N_533,N_228);
and U1460 (N_1460,N_9,N_476);
or U1461 (N_1461,N_154,N_666);
or U1462 (N_1462,N_388,N_77);
nor U1463 (N_1463,N_695,N_418);
nor U1464 (N_1464,N_319,N_592);
nand U1465 (N_1465,N_87,N_629);
nand U1466 (N_1466,N_90,N_18);
nor U1467 (N_1467,N_353,N_414);
nor U1468 (N_1468,N_374,N_517);
or U1469 (N_1469,N_449,N_347);
xnor U1470 (N_1470,N_702,N_511);
nor U1471 (N_1471,N_269,N_560);
nand U1472 (N_1472,N_19,N_355);
nor U1473 (N_1473,N_401,N_198);
and U1474 (N_1474,N_209,N_407);
and U1475 (N_1475,N_600,N_720);
and U1476 (N_1476,N_198,N_703);
nor U1477 (N_1477,N_172,N_741);
nor U1478 (N_1478,N_587,N_305);
or U1479 (N_1479,N_476,N_56);
and U1480 (N_1480,N_298,N_108);
and U1481 (N_1481,N_18,N_207);
or U1482 (N_1482,N_301,N_514);
or U1483 (N_1483,N_176,N_283);
and U1484 (N_1484,N_169,N_442);
xor U1485 (N_1485,N_429,N_418);
nor U1486 (N_1486,N_490,N_692);
nand U1487 (N_1487,N_30,N_507);
and U1488 (N_1488,N_641,N_627);
or U1489 (N_1489,N_282,N_555);
or U1490 (N_1490,N_46,N_747);
or U1491 (N_1491,N_511,N_245);
nand U1492 (N_1492,N_434,N_739);
nand U1493 (N_1493,N_184,N_325);
and U1494 (N_1494,N_464,N_671);
and U1495 (N_1495,N_575,N_635);
or U1496 (N_1496,N_448,N_125);
and U1497 (N_1497,N_363,N_724);
nor U1498 (N_1498,N_676,N_720);
nor U1499 (N_1499,N_221,N_544);
or U1500 (N_1500,N_853,N_1069);
nor U1501 (N_1501,N_1048,N_817);
or U1502 (N_1502,N_1274,N_1297);
xor U1503 (N_1503,N_949,N_1340);
xnor U1504 (N_1504,N_1271,N_866);
xnor U1505 (N_1505,N_854,N_1146);
nor U1506 (N_1506,N_861,N_1250);
and U1507 (N_1507,N_1483,N_1093);
nand U1508 (N_1508,N_1468,N_1411);
nor U1509 (N_1509,N_1195,N_1349);
or U1510 (N_1510,N_1212,N_1078);
and U1511 (N_1511,N_998,N_926);
or U1512 (N_1512,N_1403,N_1181);
nor U1513 (N_1513,N_1236,N_992);
and U1514 (N_1514,N_1438,N_818);
or U1515 (N_1515,N_1138,N_1272);
or U1516 (N_1516,N_1261,N_1049);
or U1517 (N_1517,N_1301,N_1154);
nand U1518 (N_1518,N_1270,N_1105);
and U1519 (N_1519,N_1159,N_1267);
xnor U1520 (N_1520,N_1035,N_1022);
nor U1521 (N_1521,N_1453,N_1056);
nand U1522 (N_1522,N_907,N_968);
nor U1523 (N_1523,N_1055,N_1444);
nor U1524 (N_1524,N_1322,N_922);
nor U1525 (N_1525,N_1439,N_1366);
nand U1526 (N_1526,N_1149,N_912);
nor U1527 (N_1527,N_1188,N_852);
nor U1528 (N_1528,N_1239,N_945);
or U1529 (N_1529,N_1133,N_890);
nor U1530 (N_1530,N_1217,N_782);
nor U1531 (N_1531,N_971,N_1039);
nor U1532 (N_1532,N_1449,N_1058);
nand U1533 (N_1533,N_906,N_751);
and U1534 (N_1534,N_878,N_1112);
nand U1535 (N_1535,N_1163,N_1458);
nor U1536 (N_1536,N_1382,N_1354);
nor U1537 (N_1537,N_1399,N_975);
and U1538 (N_1538,N_842,N_1356);
nor U1539 (N_1539,N_1156,N_1174);
or U1540 (N_1540,N_1185,N_1479);
nor U1541 (N_1541,N_1276,N_851);
nand U1542 (N_1542,N_1030,N_934);
nor U1543 (N_1543,N_1214,N_1355);
or U1544 (N_1544,N_924,N_1189);
or U1545 (N_1545,N_997,N_899);
or U1546 (N_1546,N_1073,N_1344);
nand U1547 (N_1547,N_1464,N_1235);
or U1548 (N_1548,N_1300,N_1173);
or U1549 (N_1549,N_859,N_1027);
nand U1550 (N_1550,N_919,N_913);
nand U1551 (N_1551,N_1298,N_1440);
nor U1552 (N_1552,N_895,N_909);
and U1553 (N_1553,N_1315,N_994);
nand U1554 (N_1554,N_1002,N_1160);
or U1555 (N_1555,N_1392,N_1342);
or U1556 (N_1556,N_1364,N_1243);
and U1557 (N_1557,N_1409,N_1213);
nand U1558 (N_1558,N_1478,N_1273);
or U1559 (N_1559,N_1321,N_921);
or U1560 (N_1560,N_1038,N_1068);
nor U1561 (N_1561,N_929,N_1117);
nor U1562 (N_1562,N_1254,N_1119);
nor U1563 (N_1563,N_1095,N_777);
and U1564 (N_1564,N_980,N_769);
and U1565 (N_1565,N_1305,N_1125);
or U1566 (N_1566,N_1000,N_1231);
and U1567 (N_1567,N_1140,N_1359);
nand U1568 (N_1568,N_858,N_939);
nor U1569 (N_1569,N_1345,N_1278);
or U1570 (N_1570,N_819,N_938);
and U1571 (N_1571,N_954,N_843);
nor U1572 (N_1572,N_1425,N_902);
nand U1573 (N_1573,N_1215,N_821);
nor U1574 (N_1574,N_1040,N_1318);
nand U1575 (N_1575,N_1207,N_1017);
nand U1576 (N_1576,N_1263,N_1186);
and U1577 (N_1577,N_1171,N_814);
and U1578 (N_1578,N_811,N_1020);
nor U1579 (N_1579,N_1323,N_1152);
nor U1580 (N_1580,N_1240,N_1131);
and U1581 (N_1581,N_776,N_809);
nor U1582 (N_1582,N_753,N_754);
nor U1583 (N_1583,N_1103,N_1208);
nor U1584 (N_1584,N_1075,N_1437);
xor U1585 (N_1585,N_1130,N_959);
and U1586 (N_1586,N_1484,N_1268);
nand U1587 (N_1587,N_1311,N_765);
nand U1588 (N_1588,N_1158,N_1187);
nand U1589 (N_1589,N_856,N_993);
or U1590 (N_1590,N_836,N_1225);
nand U1591 (N_1591,N_885,N_1378);
and U1592 (N_1592,N_1367,N_1481);
and U1593 (N_1593,N_1441,N_1150);
and U1594 (N_1594,N_1447,N_812);
nand U1595 (N_1595,N_847,N_1129);
nand U1596 (N_1596,N_1386,N_797);
nor U1597 (N_1597,N_1423,N_862);
xor U1598 (N_1598,N_974,N_824);
nor U1599 (N_1599,N_1398,N_1269);
nand U1600 (N_1600,N_958,N_1396);
nor U1601 (N_1601,N_1059,N_1353);
nor U1602 (N_1602,N_822,N_793);
xnor U1603 (N_1603,N_1196,N_867);
or U1604 (N_1604,N_850,N_1326);
nand U1605 (N_1605,N_1294,N_1029);
nand U1606 (N_1606,N_927,N_1127);
nor U1607 (N_1607,N_1142,N_1332);
nand U1608 (N_1608,N_1486,N_760);
or U1609 (N_1609,N_1256,N_877);
and U1610 (N_1610,N_1111,N_1167);
nor U1611 (N_1611,N_1408,N_1110);
nor U1612 (N_1612,N_1108,N_764);
or U1613 (N_1613,N_1106,N_807);
nor U1614 (N_1614,N_1116,N_1287);
or U1615 (N_1615,N_1026,N_957);
nand U1616 (N_1616,N_1216,N_1090);
nor U1617 (N_1617,N_961,N_1404);
nor U1618 (N_1618,N_991,N_1406);
xnor U1619 (N_1619,N_955,N_804);
nor U1620 (N_1620,N_1184,N_1044);
or U1621 (N_1621,N_1424,N_872);
nor U1622 (N_1622,N_1050,N_780);
nor U1623 (N_1623,N_984,N_1472);
nand U1624 (N_1624,N_1168,N_1065);
nor U1625 (N_1625,N_1005,N_799);
or U1626 (N_1626,N_1368,N_1452);
nand U1627 (N_1627,N_1202,N_1200);
or U1628 (N_1628,N_1348,N_1400);
or U1629 (N_1629,N_865,N_1247);
nor U1630 (N_1630,N_1289,N_838);
nor U1631 (N_1631,N_1052,N_1114);
or U1632 (N_1632,N_946,N_1204);
xnor U1633 (N_1633,N_1081,N_966);
and U1634 (N_1634,N_792,N_983);
nor U1635 (N_1635,N_1191,N_933);
nor U1636 (N_1636,N_800,N_1120);
or U1637 (N_1637,N_1221,N_857);
nand U1638 (N_1638,N_916,N_1285);
and U1639 (N_1639,N_805,N_1016);
or U1640 (N_1640,N_1141,N_1320);
nor U1641 (N_1641,N_1019,N_1024);
nand U1642 (N_1642,N_988,N_1015);
or U1643 (N_1643,N_1197,N_940);
or U1644 (N_1644,N_1061,N_1257);
nor U1645 (N_1645,N_1262,N_1288);
nand U1646 (N_1646,N_1265,N_1280);
nand U1647 (N_1647,N_1079,N_875);
nor U1648 (N_1648,N_1242,N_823);
nor U1649 (N_1649,N_1162,N_1165);
nor U1650 (N_1650,N_1302,N_953);
and U1651 (N_1651,N_1067,N_1362);
nor U1652 (N_1652,N_869,N_896);
nand U1653 (N_1653,N_1429,N_759);
nor U1654 (N_1654,N_1192,N_1246);
xor U1655 (N_1655,N_825,N_1018);
or U1656 (N_1656,N_1376,N_766);
nand U1657 (N_1657,N_1380,N_1226);
nand U1658 (N_1658,N_1476,N_1066);
nand U1659 (N_1659,N_967,N_1175);
nor U1660 (N_1660,N_794,N_1477);
nor U1661 (N_1661,N_999,N_964);
or U1662 (N_1662,N_1091,N_1033);
or U1663 (N_1663,N_1292,N_1474);
nor U1664 (N_1664,N_889,N_1222);
xnor U1665 (N_1665,N_1054,N_876);
nor U1666 (N_1666,N_950,N_1490);
or U1667 (N_1667,N_860,N_874);
nor U1668 (N_1668,N_1194,N_841);
and U1669 (N_1669,N_910,N_1172);
or U1670 (N_1670,N_786,N_802);
nand U1671 (N_1671,N_1405,N_844);
nor U1672 (N_1672,N_1281,N_918);
nor U1673 (N_1673,N_1233,N_1180);
nand U1674 (N_1674,N_960,N_773);
nand U1675 (N_1675,N_1433,N_1334);
nor U1676 (N_1676,N_1494,N_925);
nand U1677 (N_1677,N_1388,N_1104);
nand U1678 (N_1678,N_1137,N_1060);
nand U1679 (N_1679,N_1198,N_1369);
or U1680 (N_1680,N_880,N_1465);
nand U1681 (N_1681,N_1488,N_1014);
nand U1682 (N_1682,N_1331,N_1128);
or U1683 (N_1683,N_1459,N_1211);
nand U1684 (N_1684,N_774,N_1365);
nor U1685 (N_1685,N_1357,N_1309);
nor U1686 (N_1686,N_1275,N_1199);
nand U1687 (N_1687,N_813,N_790);
and U1688 (N_1688,N_1312,N_1493);
nor U1689 (N_1689,N_1361,N_1329);
nor U1690 (N_1690,N_952,N_1304);
nand U1691 (N_1691,N_1469,N_1012);
nor U1692 (N_1692,N_898,N_914);
or U1693 (N_1693,N_995,N_1371);
nor U1694 (N_1694,N_928,N_830);
nor U1695 (N_1695,N_1126,N_1134);
nor U1696 (N_1696,N_1201,N_936);
or U1697 (N_1697,N_1179,N_868);
and U1698 (N_1698,N_923,N_1397);
nand U1699 (N_1699,N_1383,N_848);
and U1700 (N_1700,N_1417,N_943);
and U1701 (N_1701,N_1025,N_1006);
nor U1702 (N_1702,N_970,N_1284);
or U1703 (N_1703,N_911,N_1489);
and U1704 (N_1704,N_944,N_1370);
or U1705 (N_1705,N_1454,N_1295);
nor U1706 (N_1706,N_1121,N_1031);
and U1707 (N_1707,N_1456,N_1251);
and U1708 (N_1708,N_973,N_1496);
or U1709 (N_1709,N_881,N_932);
and U1710 (N_1710,N_1495,N_837);
and U1711 (N_1711,N_1099,N_781);
or U1712 (N_1712,N_1237,N_1339);
and U1713 (N_1713,N_835,N_750);
or U1714 (N_1714,N_1123,N_976);
or U1715 (N_1715,N_1161,N_789);
nor U1716 (N_1716,N_1085,N_1100);
nand U1717 (N_1717,N_1087,N_1457);
nand U1718 (N_1718,N_829,N_761);
or U1719 (N_1719,N_1375,N_1310);
nand U1720 (N_1720,N_900,N_979);
nor U1721 (N_1721,N_864,N_1144);
and U1722 (N_1722,N_1410,N_1177);
nor U1723 (N_1723,N_904,N_1442);
nand U1724 (N_1724,N_1135,N_1455);
or U1725 (N_1725,N_1166,N_1157);
or U1726 (N_1726,N_963,N_1415);
and U1727 (N_1727,N_1307,N_886);
and U1728 (N_1728,N_1228,N_1450);
or U1729 (N_1729,N_1098,N_1283);
nor U1730 (N_1730,N_1374,N_1259);
and U1731 (N_1731,N_1363,N_1151);
nand U1732 (N_1732,N_1028,N_1462);
nor U1733 (N_1733,N_972,N_1080);
or U1734 (N_1734,N_1210,N_1487);
nor U1735 (N_1735,N_969,N_1064);
nand U1736 (N_1736,N_1043,N_1070);
xnor U1737 (N_1737,N_1384,N_1206);
or U1738 (N_1738,N_756,N_1325);
xor U1739 (N_1739,N_948,N_752);
and U1740 (N_1740,N_810,N_1482);
and U1741 (N_1741,N_834,N_808);
and U1742 (N_1742,N_803,N_771);
xor U1743 (N_1743,N_1096,N_1203);
and U1744 (N_1744,N_1248,N_1143);
and U1745 (N_1745,N_775,N_1467);
nand U1746 (N_1746,N_1277,N_1394);
or U1747 (N_1747,N_1351,N_1083);
and U1748 (N_1748,N_1491,N_1074);
or U1749 (N_1749,N_1021,N_1088);
nor U1750 (N_1750,N_1153,N_1385);
or U1751 (N_1751,N_1390,N_1232);
or U1752 (N_1752,N_871,N_1089);
nor U1753 (N_1753,N_883,N_870);
and U1754 (N_1754,N_798,N_1443);
or U1755 (N_1755,N_1042,N_1145);
nor U1756 (N_1756,N_1051,N_1109);
nor U1757 (N_1757,N_917,N_1244);
or U1758 (N_1758,N_796,N_863);
nand U1759 (N_1759,N_996,N_1499);
nor U1760 (N_1760,N_1234,N_1279);
xor U1761 (N_1761,N_941,N_981);
and U1762 (N_1762,N_1473,N_951);
nand U1763 (N_1763,N_956,N_828);
and U1764 (N_1764,N_1107,N_1422);
and U1765 (N_1765,N_840,N_772);
nand U1766 (N_1766,N_1148,N_1092);
or U1767 (N_1767,N_1498,N_1076);
and U1768 (N_1768,N_1434,N_1224);
xor U1769 (N_1769,N_1402,N_1346);
nand U1770 (N_1770,N_1497,N_755);
nand U1771 (N_1771,N_1072,N_1249);
xor U1772 (N_1772,N_891,N_1082);
nor U1773 (N_1773,N_1164,N_831);
nand U1774 (N_1774,N_901,N_1373);
and U1775 (N_1775,N_937,N_1293);
or U1776 (N_1776,N_1391,N_1102);
nand U1777 (N_1777,N_990,N_816);
or U1778 (N_1778,N_1466,N_985);
nor U1779 (N_1779,N_1001,N_1034);
nor U1780 (N_1780,N_845,N_833);
nand U1781 (N_1781,N_849,N_1436);
or U1782 (N_1782,N_1299,N_1448);
nor U1783 (N_1783,N_1182,N_1347);
nand U1784 (N_1784,N_1238,N_1337);
nor U1785 (N_1785,N_768,N_884);
nand U1786 (N_1786,N_1253,N_894);
nor U1787 (N_1787,N_762,N_1046);
or U1788 (N_1788,N_783,N_931);
or U1789 (N_1789,N_1336,N_1350);
or U1790 (N_1790,N_1183,N_1328);
and U1791 (N_1791,N_965,N_1147);
or U1792 (N_1792,N_1245,N_987);
nand U1793 (N_1793,N_1229,N_815);
xor U1794 (N_1794,N_1352,N_1430);
nor U1795 (N_1795,N_1389,N_1011);
and U1796 (N_1796,N_1319,N_826);
xnor U1797 (N_1797,N_935,N_1032);
and U1798 (N_1798,N_1264,N_1372);
nor U1799 (N_1799,N_767,N_1314);
or U1800 (N_1800,N_1115,N_893);
nor U1801 (N_1801,N_1062,N_1266);
and U1802 (N_1802,N_977,N_905);
nor U1803 (N_1803,N_1013,N_1252);
or U1804 (N_1804,N_1041,N_779);
nor U1805 (N_1805,N_806,N_788);
or U1806 (N_1806,N_1308,N_1053);
and U1807 (N_1807,N_1463,N_791);
nor U1808 (N_1808,N_763,N_920);
nand U1809 (N_1809,N_787,N_1341);
nand U1810 (N_1810,N_1071,N_1139);
nor U1811 (N_1811,N_1057,N_1136);
nor U1812 (N_1812,N_1471,N_1333);
or U1813 (N_1813,N_1255,N_989);
nand U1814 (N_1814,N_1037,N_1023);
or U1815 (N_1815,N_1327,N_1230);
nor U1816 (N_1816,N_1063,N_1227);
and U1817 (N_1817,N_1432,N_1418);
nor U1818 (N_1818,N_1475,N_942);
nand U1819 (N_1819,N_846,N_820);
nor U1820 (N_1820,N_1176,N_1492);
and U1821 (N_1821,N_1451,N_1086);
and U1822 (N_1822,N_1101,N_1335);
nor U1823 (N_1823,N_1324,N_1047);
or U1824 (N_1824,N_1155,N_1036);
nand U1825 (N_1825,N_1313,N_982);
or U1826 (N_1826,N_1045,N_1113);
nand U1827 (N_1827,N_770,N_1218);
nor U1828 (N_1828,N_801,N_757);
nand U1829 (N_1829,N_1132,N_1084);
nand U1830 (N_1830,N_1077,N_1220);
nor U1831 (N_1831,N_839,N_1330);
nand U1832 (N_1832,N_778,N_1395);
or U1833 (N_1833,N_882,N_1306);
nand U1834 (N_1834,N_1343,N_1407);
or U1835 (N_1835,N_1009,N_962);
and U1836 (N_1836,N_1461,N_1205);
nor U1837 (N_1837,N_1446,N_827);
or U1838 (N_1838,N_1427,N_1122);
nor U1839 (N_1839,N_1097,N_784);
nand U1840 (N_1840,N_873,N_1416);
and U1841 (N_1841,N_947,N_1169);
or U1842 (N_1842,N_1094,N_1170);
and U1843 (N_1843,N_1413,N_1421);
and U1844 (N_1844,N_1178,N_1010);
nor U1845 (N_1845,N_1435,N_879);
nand U1846 (N_1846,N_795,N_1379);
and U1847 (N_1847,N_1412,N_915);
and U1848 (N_1848,N_1485,N_978);
or U1849 (N_1849,N_758,N_930);
nor U1850 (N_1850,N_897,N_1286);
nand U1851 (N_1851,N_1316,N_1401);
nor U1852 (N_1852,N_1008,N_1260);
or U1853 (N_1853,N_1124,N_1282);
or U1854 (N_1854,N_1426,N_888);
nand U1855 (N_1855,N_1358,N_1381);
or U1856 (N_1856,N_1419,N_892);
or U1857 (N_1857,N_887,N_1007);
nor U1858 (N_1858,N_1190,N_1480);
nor U1859 (N_1859,N_1193,N_855);
nor U1860 (N_1860,N_785,N_1291);
nor U1861 (N_1861,N_1338,N_1303);
or U1862 (N_1862,N_1460,N_1360);
or U1863 (N_1863,N_1470,N_1420);
or U1864 (N_1864,N_1377,N_1223);
or U1865 (N_1865,N_1003,N_908);
and U1866 (N_1866,N_903,N_1118);
or U1867 (N_1867,N_1317,N_1296);
or U1868 (N_1868,N_1241,N_1393);
or U1869 (N_1869,N_832,N_1004);
nand U1870 (N_1870,N_1290,N_1445);
nor U1871 (N_1871,N_1431,N_1209);
nand U1872 (N_1872,N_1258,N_986);
and U1873 (N_1873,N_1219,N_1428);
or U1874 (N_1874,N_1387,N_1414);
nand U1875 (N_1875,N_1364,N_797);
nor U1876 (N_1876,N_751,N_1498);
or U1877 (N_1877,N_1037,N_1355);
and U1878 (N_1878,N_1147,N_1300);
or U1879 (N_1879,N_865,N_965);
or U1880 (N_1880,N_1085,N_1222);
nand U1881 (N_1881,N_1256,N_1429);
nand U1882 (N_1882,N_1070,N_1327);
and U1883 (N_1883,N_1335,N_1395);
or U1884 (N_1884,N_1477,N_956);
and U1885 (N_1885,N_1324,N_805);
nor U1886 (N_1886,N_1266,N_995);
and U1887 (N_1887,N_999,N_1092);
nand U1888 (N_1888,N_1312,N_1462);
nor U1889 (N_1889,N_1003,N_1012);
and U1890 (N_1890,N_846,N_1122);
or U1891 (N_1891,N_1386,N_864);
nor U1892 (N_1892,N_1301,N_1345);
and U1893 (N_1893,N_1343,N_948);
or U1894 (N_1894,N_916,N_982);
or U1895 (N_1895,N_1059,N_1026);
and U1896 (N_1896,N_1202,N_1381);
or U1897 (N_1897,N_801,N_1425);
xor U1898 (N_1898,N_1031,N_1373);
or U1899 (N_1899,N_1306,N_1275);
xor U1900 (N_1900,N_922,N_1309);
or U1901 (N_1901,N_1000,N_785);
or U1902 (N_1902,N_1438,N_977);
or U1903 (N_1903,N_876,N_1345);
or U1904 (N_1904,N_1397,N_878);
nand U1905 (N_1905,N_1385,N_1393);
xnor U1906 (N_1906,N_1384,N_1439);
nand U1907 (N_1907,N_1212,N_1182);
or U1908 (N_1908,N_959,N_1028);
nor U1909 (N_1909,N_1388,N_1010);
or U1910 (N_1910,N_1484,N_1458);
nand U1911 (N_1911,N_1034,N_970);
nand U1912 (N_1912,N_1215,N_1022);
or U1913 (N_1913,N_1351,N_776);
nor U1914 (N_1914,N_822,N_1426);
and U1915 (N_1915,N_1439,N_857);
nor U1916 (N_1916,N_843,N_1479);
nor U1917 (N_1917,N_861,N_939);
and U1918 (N_1918,N_998,N_891);
nand U1919 (N_1919,N_808,N_935);
and U1920 (N_1920,N_1133,N_780);
and U1921 (N_1921,N_1120,N_893);
nor U1922 (N_1922,N_1119,N_1395);
and U1923 (N_1923,N_1498,N_1353);
nor U1924 (N_1924,N_1191,N_1018);
or U1925 (N_1925,N_1394,N_1439);
nor U1926 (N_1926,N_843,N_1024);
or U1927 (N_1927,N_1066,N_1273);
and U1928 (N_1928,N_1184,N_1167);
nand U1929 (N_1929,N_879,N_1498);
nand U1930 (N_1930,N_1046,N_1389);
nand U1931 (N_1931,N_1031,N_997);
nand U1932 (N_1932,N_1319,N_1358);
nand U1933 (N_1933,N_1113,N_831);
and U1934 (N_1934,N_813,N_1113);
and U1935 (N_1935,N_1083,N_930);
nor U1936 (N_1936,N_829,N_1443);
nand U1937 (N_1937,N_1309,N_1092);
nor U1938 (N_1938,N_755,N_972);
or U1939 (N_1939,N_1301,N_1102);
and U1940 (N_1940,N_951,N_1320);
and U1941 (N_1941,N_785,N_1129);
nor U1942 (N_1942,N_1265,N_1491);
nand U1943 (N_1943,N_948,N_888);
and U1944 (N_1944,N_1042,N_1468);
nor U1945 (N_1945,N_825,N_1034);
and U1946 (N_1946,N_850,N_1156);
and U1947 (N_1947,N_1381,N_1257);
or U1948 (N_1948,N_1240,N_1394);
nor U1949 (N_1949,N_1214,N_1253);
nand U1950 (N_1950,N_1492,N_818);
and U1951 (N_1951,N_840,N_1366);
nor U1952 (N_1952,N_1131,N_806);
and U1953 (N_1953,N_1281,N_884);
nor U1954 (N_1954,N_1385,N_934);
and U1955 (N_1955,N_1299,N_1307);
nor U1956 (N_1956,N_1019,N_891);
nor U1957 (N_1957,N_1287,N_1262);
nand U1958 (N_1958,N_850,N_768);
and U1959 (N_1959,N_846,N_1126);
nand U1960 (N_1960,N_1064,N_1201);
or U1961 (N_1961,N_1158,N_898);
nor U1962 (N_1962,N_1319,N_814);
and U1963 (N_1963,N_1306,N_1337);
and U1964 (N_1964,N_785,N_1377);
and U1965 (N_1965,N_1217,N_1483);
nor U1966 (N_1966,N_1414,N_888);
nand U1967 (N_1967,N_1210,N_794);
xor U1968 (N_1968,N_1330,N_1244);
nand U1969 (N_1969,N_896,N_1081);
or U1970 (N_1970,N_1409,N_858);
and U1971 (N_1971,N_1111,N_1308);
and U1972 (N_1972,N_1365,N_1419);
nor U1973 (N_1973,N_1117,N_1232);
nand U1974 (N_1974,N_862,N_1201);
nand U1975 (N_1975,N_893,N_916);
and U1976 (N_1976,N_1043,N_1337);
nand U1977 (N_1977,N_1379,N_931);
nand U1978 (N_1978,N_1107,N_1068);
nor U1979 (N_1979,N_1419,N_1432);
or U1980 (N_1980,N_1007,N_823);
and U1981 (N_1981,N_1238,N_1381);
nand U1982 (N_1982,N_797,N_1435);
and U1983 (N_1983,N_1270,N_854);
or U1984 (N_1984,N_1427,N_1494);
or U1985 (N_1985,N_1006,N_1382);
and U1986 (N_1986,N_911,N_1268);
or U1987 (N_1987,N_1392,N_1352);
nor U1988 (N_1988,N_1191,N_825);
or U1989 (N_1989,N_967,N_769);
nand U1990 (N_1990,N_1076,N_1228);
nor U1991 (N_1991,N_773,N_1319);
or U1992 (N_1992,N_1191,N_1102);
nand U1993 (N_1993,N_1473,N_1324);
and U1994 (N_1994,N_1001,N_1057);
or U1995 (N_1995,N_1061,N_817);
nand U1996 (N_1996,N_785,N_1083);
and U1997 (N_1997,N_892,N_1310);
and U1998 (N_1998,N_1113,N_1275);
nor U1999 (N_1999,N_1104,N_1298);
nor U2000 (N_2000,N_762,N_964);
nor U2001 (N_2001,N_981,N_993);
or U2002 (N_2002,N_1238,N_1087);
or U2003 (N_2003,N_1483,N_1245);
nand U2004 (N_2004,N_1298,N_1452);
nor U2005 (N_2005,N_1074,N_1137);
nand U2006 (N_2006,N_894,N_1333);
and U2007 (N_2007,N_1331,N_915);
nand U2008 (N_2008,N_768,N_1292);
or U2009 (N_2009,N_817,N_961);
or U2010 (N_2010,N_1357,N_1381);
nor U2011 (N_2011,N_941,N_1072);
and U2012 (N_2012,N_853,N_1432);
nor U2013 (N_2013,N_823,N_1075);
nor U2014 (N_2014,N_1213,N_1076);
and U2015 (N_2015,N_767,N_1483);
nand U2016 (N_2016,N_997,N_1020);
xnor U2017 (N_2017,N_1304,N_1179);
nor U2018 (N_2018,N_1065,N_1095);
nand U2019 (N_2019,N_1367,N_1049);
and U2020 (N_2020,N_1346,N_1383);
or U2021 (N_2021,N_1097,N_1068);
or U2022 (N_2022,N_938,N_1002);
nand U2023 (N_2023,N_842,N_1343);
nand U2024 (N_2024,N_1105,N_1254);
or U2025 (N_2025,N_1347,N_1069);
and U2026 (N_2026,N_959,N_1356);
and U2027 (N_2027,N_1308,N_1043);
and U2028 (N_2028,N_1432,N_1460);
or U2029 (N_2029,N_1407,N_1242);
nor U2030 (N_2030,N_1398,N_890);
or U2031 (N_2031,N_777,N_751);
nor U2032 (N_2032,N_960,N_1022);
nand U2033 (N_2033,N_875,N_837);
nor U2034 (N_2034,N_1482,N_848);
and U2035 (N_2035,N_913,N_1127);
xnor U2036 (N_2036,N_1178,N_1264);
and U2037 (N_2037,N_836,N_1405);
or U2038 (N_2038,N_793,N_1321);
nor U2039 (N_2039,N_1437,N_1050);
or U2040 (N_2040,N_1402,N_1426);
nand U2041 (N_2041,N_1057,N_1394);
nor U2042 (N_2042,N_849,N_975);
nand U2043 (N_2043,N_1088,N_1228);
and U2044 (N_2044,N_1458,N_881);
nand U2045 (N_2045,N_964,N_876);
xor U2046 (N_2046,N_1047,N_1153);
nor U2047 (N_2047,N_1159,N_953);
or U2048 (N_2048,N_1367,N_988);
nand U2049 (N_2049,N_1403,N_1233);
nor U2050 (N_2050,N_1355,N_1193);
or U2051 (N_2051,N_1071,N_1395);
and U2052 (N_2052,N_1035,N_1442);
nand U2053 (N_2053,N_1240,N_1379);
nand U2054 (N_2054,N_1156,N_1420);
xor U2055 (N_2055,N_1000,N_930);
nand U2056 (N_2056,N_1341,N_1398);
and U2057 (N_2057,N_1346,N_1164);
and U2058 (N_2058,N_1443,N_1274);
nor U2059 (N_2059,N_1410,N_883);
or U2060 (N_2060,N_1254,N_1427);
nand U2061 (N_2061,N_978,N_1319);
or U2062 (N_2062,N_1153,N_819);
nor U2063 (N_2063,N_1002,N_784);
nand U2064 (N_2064,N_1298,N_905);
nor U2065 (N_2065,N_1030,N_1317);
or U2066 (N_2066,N_1491,N_818);
and U2067 (N_2067,N_1417,N_1110);
nor U2068 (N_2068,N_1095,N_1273);
nor U2069 (N_2069,N_770,N_1012);
nor U2070 (N_2070,N_1390,N_959);
or U2071 (N_2071,N_1373,N_840);
or U2072 (N_2072,N_1264,N_1022);
or U2073 (N_2073,N_1331,N_812);
or U2074 (N_2074,N_1105,N_890);
and U2075 (N_2075,N_799,N_797);
and U2076 (N_2076,N_1000,N_1295);
nand U2077 (N_2077,N_1272,N_1436);
and U2078 (N_2078,N_1395,N_1032);
nor U2079 (N_2079,N_990,N_1031);
nor U2080 (N_2080,N_1136,N_931);
or U2081 (N_2081,N_1468,N_997);
and U2082 (N_2082,N_1240,N_988);
nor U2083 (N_2083,N_1491,N_769);
and U2084 (N_2084,N_1193,N_773);
nor U2085 (N_2085,N_1462,N_1355);
or U2086 (N_2086,N_1118,N_1095);
nand U2087 (N_2087,N_1107,N_763);
or U2088 (N_2088,N_1098,N_755);
nor U2089 (N_2089,N_1256,N_1407);
nor U2090 (N_2090,N_1476,N_1076);
nand U2091 (N_2091,N_1029,N_876);
nor U2092 (N_2092,N_797,N_1246);
or U2093 (N_2093,N_1159,N_1107);
nand U2094 (N_2094,N_1348,N_1106);
and U2095 (N_2095,N_1005,N_1310);
or U2096 (N_2096,N_903,N_1025);
nand U2097 (N_2097,N_824,N_1085);
nand U2098 (N_2098,N_947,N_917);
nand U2099 (N_2099,N_1326,N_858);
xor U2100 (N_2100,N_1345,N_895);
and U2101 (N_2101,N_820,N_1446);
xnor U2102 (N_2102,N_1343,N_1078);
nor U2103 (N_2103,N_1128,N_1469);
or U2104 (N_2104,N_1195,N_946);
nand U2105 (N_2105,N_864,N_1327);
nand U2106 (N_2106,N_1105,N_879);
nand U2107 (N_2107,N_1046,N_1077);
nand U2108 (N_2108,N_866,N_1369);
nor U2109 (N_2109,N_897,N_954);
or U2110 (N_2110,N_1477,N_1249);
nand U2111 (N_2111,N_1459,N_1289);
nor U2112 (N_2112,N_999,N_1498);
and U2113 (N_2113,N_1406,N_1130);
nand U2114 (N_2114,N_816,N_1454);
nor U2115 (N_2115,N_1380,N_1078);
and U2116 (N_2116,N_931,N_1231);
or U2117 (N_2117,N_921,N_1483);
and U2118 (N_2118,N_1224,N_796);
nor U2119 (N_2119,N_1057,N_1023);
nand U2120 (N_2120,N_768,N_990);
or U2121 (N_2121,N_817,N_950);
and U2122 (N_2122,N_922,N_862);
nor U2123 (N_2123,N_1200,N_1001);
nand U2124 (N_2124,N_1073,N_1044);
or U2125 (N_2125,N_1085,N_1044);
or U2126 (N_2126,N_1288,N_867);
nand U2127 (N_2127,N_1112,N_1401);
and U2128 (N_2128,N_985,N_1071);
and U2129 (N_2129,N_868,N_1397);
nand U2130 (N_2130,N_1292,N_1014);
or U2131 (N_2131,N_1168,N_936);
nand U2132 (N_2132,N_888,N_930);
nand U2133 (N_2133,N_1374,N_1303);
nor U2134 (N_2134,N_1304,N_810);
or U2135 (N_2135,N_925,N_1485);
nor U2136 (N_2136,N_849,N_1245);
nand U2137 (N_2137,N_1104,N_801);
and U2138 (N_2138,N_898,N_1011);
or U2139 (N_2139,N_1154,N_1482);
and U2140 (N_2140,N_1316,N_1344);
xnor U2141 (N_2141,N_1232,N_825);
nor U2142 (N_2142,N_1102,N_1221);
nand U2143 (N_2143,N_841,N_1184);
and U2144 (N_2144,N_1421,N_950);
or U2145 (N_2145,N_1489,N_1472);
nor U2146 (N_2146,N_1008,N_1038);
nor U2147 (N_2147,N_1349,N_1194);
and U2148 (N_2148,N_1211,N_1143);
nor U2149 (N_2149,N_1022,N_884);
or U2150 (N_2150,N_1104,N_1336);
nor U2151 (N_2151,N_759,N_1192);
and U2152 (N_2152,N_1123,N_777);
nor U2153 (N_2153,N_1142,N_1274);
and U2154 (N_2154,N_849,N_1009);
or U2155 (N_2155,N_1152,N_1307);
nand U2156 (N_2156,N_1087,N_1167);
nand U2157 (N_2157,N_1456,N_968);
or U2158 (N_2158,N_1305,N_815);
and U2159 (N_2159,N_887,N_1233);
nand U2160 (N_2160,N_1204,N_1404);
and U2161 (N_2161,N_897,N_913);
nand U2162 (N_2162,N_1238,N_978);
or U2163 (N_2163,N_1012,N_1106);
or U2164 (N_2164,N_945,N_1191);
nor U2165 (N_2165,N_789,N_819);
nor U2166 (N_2166,N_1073,N_1256);
or U2167 (N_2167,N_1435,N_1453);
nand U2168 (N_2168,N_1448,N_906);
or U2169 (N_2169,N_1141,N_855);
nor U2170 (N_2170,N_1288,N_1263);
or U2171 (N_2171,N_922,N_1099);
or U2172 (N_2172,N_959,N_1113);
or U2173 (N_2173,N_905,N_1090);
and U2174 (N_2174,N_880,N_1485);
nor U2175 (N_2175,N_956,N_947);
nand U2176 (N_2176,N_1055,N_1253);
and U2177 (N_2177,N_1275,N_982);
nand U2178 (N_2178,N_1049,N_1395);
nand U2179 (N_2179,N_1490,N_1416);
or U2180 (N_2180,N_1342,N_943);
nor U2181 (N_2181,N_912,N_1194);
or U2182 (N_2182,N_928,N_934);
nor U2183 (N_2183,N_1056,N_1495);
nand U2184 (N_2184,N_1243,N_760);
or U2185 (N_2185,N_1349,N_1255);
or U2186 (N_2186,N_1426,N_1301);
nor U2187 (N_2187,N_937,N_780);
and U2188 (N_2188,N_1186,N_1200);
nand U2189 (N_2189,N_1328,N_910);
nand U2190 (N_2190,N_1253,N_854);
nand U2191 (N_2191,N_1058,N_1136);
and U2192 (N_2192,N_1451,N_1478);
nand U2193 (N_2193,N_1462,N_869);
or U2194 (N_2194,N_1373,N_956);
nand U2195 (N_2195,N_1254,N_999);
nor U2196 (N_2196,N_1278,N_1389);
nor U2197 (N_2197,N_816,N_796);
nand U2198 (N_2198,N_1190,N_1408);
and U2199 (N_2199,N_1346,N_1267);
nor U2200 (N_2200,N_1037,N_1416);
nor U2201 (N_2201,N_933,N_1392);
and U2202 (N_2202,N_1020,N_1354);
and U2203 (N_2203,N_1302,N_796);
or U2204 (N_2204,N_1395,N_1425);
or U2205 (N_2205,N_1197,N_1205);
and U2206 (N_2206,N_1210,N_1034);
nand U2207 (N_2207,N_1016,N_904);
and U2208 (N_2208,N_1402,N_1068);
or U2209 (N_2209,N_1086,N_1328);
and U2210 (N_2210,N_867,N_1176);
and U2211 (N_2211,N_772,N_937);
or U2212 (N_2212,N_1377,N_1099);
nor U2213 (N_2213,N_1423,N_1149);
or U2214 (N_2214,N_1472,N_852);
or U2215 (N_2215,N_812,N_1253);
nor U2216 (N_2216,N_845,N_1342);
nand U2217 (N_2217,N_1484,N_1013);
nor U2218 (N_2218,N_1286,N_931);
xor U2219 (N_2219,N_923,N_1027);
nand U2220 (N_2220,N_1187,N_805);
nand U2221 (N_2221,N_1121,N_1360);
nor U2222 (N_2222,N_1086,N_778);
nand U2223 (N_2223,N_1415,N_1485);
nand U2224 (N_2224,N_776,N_1256);
and U2225 (N_2225,N_1123,N_1195);
nand U2226 (N_2226,N_1391,N_1078);
or U2227 (N_2227,N_1022,N_1123);
and U2228 (N_2228,N_1129,N_1435);
and U2229 (N_2229,N_764,N_1062);
and U2230 (N_2230,N_1400,N_959);
nand U2231 (N_2231,N_799,N_1169);
or U2232 (N_2232,N_1153,N_1124);
nand U2233 (N_2233,N_1336,N_1270);
nand U2234 (N_2234,N_944,N_775);
nor U2235 (N_2235,N_1063,N_1283);
nand U2236 (N_2236,N_1113,N_1342);
nor U2237 (N_2237,N_777,N_899);
nand U2238 (N_2238,N_1006,N_1122);
nand U2239 (N_2239,N_1014,N_1313);
or U2240 (N_2240,N_1358,N_1457);
nand U2241 (N_2241,N_847,N_1107);
nand U2242 (N_2242,N_1497,N_1050);
xor U2243 (N_2243,N_1084,N_983);
nor U2244 (N_2244,N_1162,N_799);
and U2245 (N_2245,N_779,N_1410);
or U2246 (N_2246,N_840,N_789);
nor U2247 (N_2247,N_1292,N_1056);
and U2248 (N_2248,N_814,N_1191);
or U2249 (N_2249,N_1055,N_1100);
nor U2250 (N_2250,N_1521,N_1977);
or U2251 (N_2251,N_1864,N_2133);
or U2252 (N_2252,N_2076,N_2097);
nand U2253 (N_2253,N_1631,N_1790);
and U2254 (N_2254,N_2113,N_1553);
or U2255 (N_2255,N_2221,N_1670);
or U2256 (N_2256,N_1513,N_2209);
nand U2257 (N_2257,N_2173,N_1593);
nor U2258 (N_2258,N_2112,N_2036);
nand U2259 (N_2259,N_1587,N_2199);
and U2260 (N_2260,N_2163,N_1711);
nor U2261 (N_2261,N_2081,N_2176);
or U2262 (N_2262,N_1761,N_2156);
nor U2263 (N_2263,N_1556,N_1571);
nand U2264 (N_2264,N_1895,N_2120);
or U2265 (N_2265,N_2145,N_1552);
or U2266 (N_2266,N_2087,N_1902);
nor U2267 (N_2267,N_1502,N_1503);
and U2268 (N_2268,N_1615,N_1898);
and U2269 (N_2269,N_1850,N_1769);
nor U2270 (N_2270,N_2009,N_1836);
or U2271 (N_2271,N_1765,N_1572);
nor U2272 (N_2272,N_1921,N_1937);
and U2273 (N_2273,N_2110,N_2001);
xor U2274 (N_2274,N_1661,N_2062);
nand U2275 (N_2275,N_1669,N_2063);
and U2276 (N_2276,N_2045,N_1942);
nor U2277 (N_2277,N_1881,N_1815);
nand U2278 (N_2278,N_2083,N_2054);
xor U2279 (N_2279,N_2189,N_1771);
nand U2280 (N_2280,N_2164,N_2055);
xnor U2281 (N_2281,N_1967,N_2240);
or U2282 (N_2282,N_2118,N_1601);
nor U2283 (N_2283,N_1824,N_1905);
or U2284 (N_2284,N_1695,N_1520);
nand U2285 (N_2285,N_1996,N_1994);
or U2286 (N_2286,N_1692,N_1889);
nor U2287 (N_2287,N_2091,N_2033);
nand U2288 (N_2288,N_1971,N_2030);
nand U2289 (N_2289,N_1979,N_1775);
and U2290 (N_2290,N_2231,N_1506);
or U2291 (N_2291,N_1768,N_1893);
and U2292 (N_2292,N_1558,N_1726);
nor U2293 (N_2293,N_1704,N_1728);
nand U2294 (N_2294,N_1635,N_1651);
or U2295 (N_2295,N_2249,N_1604);
and U2296 (N_2296,N_2034,N_1746);
nand U2297 (N_2297,N_2024,N_1969);
and U2298 (N_2298,N_1973,N_2238);
or U2299 (N_2299,N_1993,N_2020);
and U2300 (N_2300,N_2123,N_1602);
nor U2301 (N_2301,N_1808,N_1701);
nand U2302 (N_2302,N_1913,N_2155);
nor U2303 (N_2303,N_1772,N_1823);
and U2304 (N_2304,N_1583,N_1774);
or U2305 (N_2305,N_1694,N_1674);
nor U2306 (N_2306,N_2053,N_1813);
nand U2307 (N_2307,N_1678,N_2038);
nor U2308 (N_2308,N_1589,N_1640);
or U2309 (N_2309,N_1968,N_2138);
nor U2310 (N_2310,N_1840,N_2211);
and U2311 (N_2311,N_2010,N_1956);
nand U2312 (N_2312,N_1609,N_2213);
nor U2313 (N_2313,N_1624,N_1700);
and U2314 (N_2314,N_1725,N_2170);
nor U2315 (N_2315,N_1684,N_1858);
or U2316 (N_2316,N_2245,N_2180);
or U2317 (N_2317,N_1707,N_1755);
nor U2318 (N_2318,N_1871,N_2247);
and U2319 (N_2319,N_1702,N_1687);
or U2320 (N_2320,N_1783,N_2071);
xnor U2321 (N_2321,N_2139,N_1561);
nand U2322 (N_2322,N_1779,N_1839);
and U2323 (N_2323,N_1547,N_1734);
nand U2324 (N_2324,N_1612,N_1985);
nor U2325 (N_2325,N_1543,N_2184);
or U2326 (N_2326,N_2108,N_1546);
or U2327 (N_2327,N_2142,N_1952);
nor U2328 (N_2328,N_1983,N_1744);
and U2329 (N_2329,N_2102,N_1809);
nand U2330 (N_2330,N_1667,N_2227);
nor U2331 (N_2331,N_1512,N_1819);
or U2332 (N_2332,N_2204,N_1965);
nand U2333 (N_2333,N_1685,N_1782);
or U2334 (N_2334,N_1507,N_2089);
nand U2335 (N_2335,N_1794,N_1557);
and U2336 (N_2336,N_2094,N_2151);
nand U2337 (N_2337,N_1584,N_1720);
nor U2338 (N_2338,N_1933,N_1890);
and U2339 (N_2339,N_2007,N_2185);
and U2340 (N_2340,N_2143,N_1785);
or U2341 (N_2341,N_1595,N_2157);
nand U2342 (N_2342,N_2186,N_1811);
and U2343 (N_2343,N_1975,N_2165);
and U2344 (N_2344,N_1796,N_2125);
and U2345 (N_2345,N_1800,N_2106);
and U2346 (N_2346,N_2017,N_1865);
nor U2347 (N_2347,N_1619,N_2146);
and U2348 (N_2348,N_2066,N_1888);
or U2349 (N_2349,N_1565,N_2127);
nand U2350 (N_2350,N_1723,N_2057);
nand U2351 (N_2351,N_2047,N_2107);
or U2352 (N_2352,N_1645,N_1843);
nor U2353 (N_2353,N_1943,N_1988);
and U2354 (N_2354,N_1647,N_2093);
nand U2355 (N_2355,N_1931,N_1622);
and U2356 (N_2356,N_1570,N_1999);
nand U2357 (N_2357,N_1784,N_1856);
or U2358 (N_2358,N_1925,N_2079);
or U2359 (N_2359,N_2198,N_1860);
or U2360 (N_2360,N_1880,N_2169);
or U2361 (N_2361,N_1737,N_1603);
or U2362 (N_2362,N_1665,N_1699);
and U2363 (N_2363,N_1945,N_1625);
nand U2364 (N_2364,N_1821,N_1501);
nand U2365 (N_2365,N_1677,N_2195);
or U2366 (N_2366,N_1526,N_1534);
nor U2367 (N_2367,N_1671,N_1524);
and U2368 (N_2368,N_1891,N_1878);
nand U2369 (N_2369,N_2080,N_1934);
nand U2370 (N_2370,N_2014,N_1829);
nor U2371 (N_2371,N_1909,N_1541);
nand U2372 (N_2372,N_1632,N_2100);
nand U2373 (N_2373,N_2052,N_2043);
and U2374 (N_2374,N_1830,N_1846);
or U2375 (N_2375,N_1868,N_2210);
and U2376 (N_2376,N_2166,N_1847);
and U2377 (N_2377,N_1500,N_1545);
and U2378 (N_2378,N_1703,N_1867);
nor U2379 (N_2379,N_1953,N_1714);
and U2380 (N_2380,N_2004,N_1751);
and U2381 (N_2381,N_1706,N_2104);
and U2382 (N_2382,N_1528,N_1733);
nor U2383 (N_2383,N_1582,N_1532);
or U2384 (N_2384,N_1927,N_1801);
or U2385 (N_2385,N_2220,N_1740);
nand U2386 (N_2386,N_1533,N_1688);
nor U2387 (N_2387,N_1987,N_2148);
nor U2388 (N_2388,N_2131,N_2167);
nand U2389 (N_2389,N_1636,N_2069);
or U2390 (N_2390,N_1992,N_2074);
and U2391 (N_2391,N_1818,N_1932);
or U2392 (N_2392,N_2194,N_1915);
or U2393 (N_2393,N_1510,N_2075);
and U2394 (N_2394,N_1986,N_1656);
nor U2395 (N_2395,N_2214,N_1862);
or U2396 (N_2396,N_1752,N_1568);
or U2397 (N_2397,N_1777,N_2042);
and U2398 (N_2398,N_1696,N_2215);
nor U2399 (N_2399,N_2206,N_1638);
nand U2400 (N_2400,N_2022,N_1873);
nand U2401 (N_2401,N_1792,N_2061);
nand U2402 (N_2402,N_1797,N_1957);
nand U2403 (N_2403,N_2121,N_2224);
nor U2404 (N_2404,N_1892,N_1525);
nand U2405 (N_2405,N_2239,N_1509);
and U2406 (N_2406,N_1854,N_1569);
and U2407 (N_2407,N_1770,N_2056);
nand U2408 (N_2408,N_1575,N_2019);
and U2409 (N_2409,N_2078,N_1901);
nand U2410 (N_2410,N_2124,N_1691);
nor U2411 (N_2411,N_2129,N_1807);
nand U2412 (N_2412,N_1566,N_1946);
and U2413 (N_2413,N_1982,N_1802);
nand U2414 (N_2414,N_2144,N_1544);
or U2415 (N_2415,N_2196,N_2064);
nor U2416 (N_2416,N_2025,N_2023);
nand U2417 (N_2417,N_1722,N_1920);
nand U2418 (N_2418,N_2188,N_2202);
nor U2419 (N_2419,N_2200,N_2119);
or U2420 (N_2420,N_1941,N_1837);
and U2421 (N_2421,N_1581,N_1884);
or U2422 (N_2422,N_1853,N_1991);
or U2423 (N_2423,N_1745,N_1786);
nor U2424 (N_2424,N_1773,N_1812);
nand U2425 (N_2425,N_1623,N_1519);
or U2426 (N_2426,N_2132,N_1935);
and U2427 (N_2427,N_1610,N_1579);
nand U2428 (N_2428,N_1820,N_1923);
or U2429 (N_2429,N_1650,N_1580);
nand U2430 (N_2430,N_1872,N_1620);
or U2431 (N_2431,N_1567,N_1793);
or U2432 (N_2432,N_1764,N_2225);
or U2433 (N_2433,N_2044,N_1530);
nor U2434 (N_2434,N_1531,N_1781);
or U2435 (N_2435,N_1885,N_1958);
and U2436 (N_2436,N_1637,N_1551);
xor U2437 (N_2437,N_1577,N_2149);
nand U2438 (N_2438,N_1538,N_2135);
nand U2439 (N_2439,N_1922,N_1539);
nor U2440 (N_2440,N_1592,N_2177);
nand U2441 (N_2441,N_1715,N_1762);
nor U2442 (N_2442,N_1944,N_1634);
and U2443 (N_2443,N_2218,N_1759);
nor U2444 (N_2444,N_1563,N_2222);
nand U2445 (N_2445,N_2050,N_2219);
nand U2446 (N_2446,N_1693,N_1748);
or U2447 (N_2447,N_2232,N_1559);
and U2448 (N_2448,N_1698,N_2128);
nor U2449 (N_2449,N_1641,N_1652);
nand U2450 (N_2450,N_1896,N_2242);
or U2451 (N_2451,N_1828,N_1976);
or U2452 (N_2452,N_1834,N_2116);
nand U2453 (N_2453,N_2117,N_1536);
nand U2454 (N_2454,N_1527,N_1505);
nand U2455 (N_2455,N_2197,N_2217);
or U2456 (N_2456,N_1866,N_1574);
or U2457 (N_2457,N_1766,N_1928);
nor U2458 (N_2458,N_1708,N_2048);
or U2459 (N_2459,N_1747,N_1529);
and U2460 (N_2460,N_1845,N_1537);
or U2461 (N_2461,N_1787,N_1731);
nand U2462 (N_2462,N_1826,N_1876);
nor U2463 (N_2463,N_1668,N_1599);
nor U2464 (N_2464,N_1936,N_1917);
and U2465 (N_2465,N_2178,N_1817);
nand U2466 (N_2466,N_1899,N_1960);
nand U2467 (N_2467,N_2006,N_1621);
nand U2468 (N_2468,N_2183,N_1562);
nand U2469 (N_2469,N_1814,N_1657);
and U2470 (N_2470,N_1626,N_1600);
or U2471 (N_2471,N_1964,N_1805);
xor U2472 (N_2472,N_2150,N_1646);
nor U2473 (N_2473,N_1831,N_2029);
or U2474 (N_2474,N_1676,N_1910);
or U2475 (N_2475,N_1679,N_2028);
and U2476 (N_2476,N_1738,N_1887);
nand U2477 (N_2477,N_2060,N_2193);
nor U2478 (N_2478,N_1628,N_1825);
or U2479 (N_2479,N_2190,N_1719);
and U2480 (N_2480,N_1978,N_1954);
or U2481 (N_2481,N_2012,N_2008);
and U2482 (N_2482,N_1754,N_1649);
and U2483 (N_2483,N_1857,N_1950);
nor U2484 (N_2484,N_2248,N_2162);
nor U2485 (N_2485,N_1763,N_1816);
nand U2486 (N_2486,N_2021,N_1972);
and U2487 (N_2487,N_2152,N_1717);
xor U2488 (N_2488,N_1804,N_1757);
or U2489 (N_2489,N_1861,N_2159);
nor U2490 (N_2490,N_1948,N_2115);
nand U2491 (N_2491,N_1886,N_1970);
xor U2492 (N_2492,N_1672,N_1682);
nand U2493 (N_2493,N_1535,N_1966);
nor U2494 (N_2494,N_1799,N_2137);
nor U2495 (N_2495,N_2174,N_2141);
nand U2496 (N_2496,N_1903,N_1833);
and U2497 (N_2497,N_2015,N_1877);
nand U2498 (N_2498,N_2084,N_2158);
or U2499 (N_2499,N_2243,N_2111);
and U2500 (N_2500,N_1875,N_1511);
nand U2501 (N_2501,N_1633,N_1844);
nor U2502 (N_2502,N_1659,N_2032);
or U2503 (N_2503,N_2096,N_1712);
nor U2504 (N_2504,N_1838,N_2099);
nand U2505 (N_2505,N_1930,N_1990);
nand U2506 (N_2506,N_1729,N_1666);
nor U2507 (N_2507,N_2072,N_1963);
or U2508 (N_2508,N_1705,N_2136);
xnor U2509 (N_2509,N_1642,N_1739);
nand U2510 (N_2510,N_1907,N_1736);
nor U2511 (N_2511,N_2105,N_2122);
nand U2512 (N_2512,N_2236,N_1591);
or U2513 (N_2513,N_1605,N_2126);
and U2514 (N_2514,N_1560,N_1586);
or U2515 (N_2515,N_1697,N_2179);
nand U2516 (N_2516,N_2230,N_1980);
or U2517 (N_2517,N_2086,N_1630);
nand U2518 (N_2518,N_1753,N_1806);
or U2519 (N_2519,N_1616,N_1835);
or U2520 (N_2520,N_2095,N_1997);
nand U2521 (N_2521,N_2208,N_2046);
nor U2522 (N_2522,N_2077,N_1908);
nor U2523 (N_2523,N_2191,N_1750);
nand U2524 (N_2524,N_2201,N_1949);
or U2525 (N_2525,N_1981,N_2026);
or U2526 (N_2526,N_2246,N_1710);
nand U2527 (N_2527,N_1690,N_1962);
or U2528 (N_2528,N_1658,N_1655);
and U2529 (N_2529,N_1554,N_1732);
or U2530 (N_2530,N_1906,N_1741);
nor U2531 (N_2531,N_1718,N_2098);
nand U2532 (N_2532,N_1742,N_2154);
or U2533 (N_2533,N_1550,N_1743);
nand U2534 (N_2534,N_1673,N_1596);
nand U2535 (N_2535,N_1897,N_1578);
or U2536 (N_2536,N_1852,N_2241);
nand U2537 (N_2537,N_1675,N_2229);
nor U2538 (N_2538,N_1919,N_2182);
nand U2539 (N_2539,N_1776,N_1998);
nor U2540 (N_2540,N_2041,N_1959);
nor U2541 (N_2541,N_2160,N_1851);
and U2542 (N_2542,N_1618,N_1863);
nand U2543 (N_2543,N_1724,N_1680);
or U2544 (N_2544,N_1548,N_1951);
and U2545 (N_2545,N_1540,N_2109);
nor U2546 (N_2546,N_2031,N_2171);
nor U2547 (N_2547,N_1924,N_2039);
and U2548 (N_2548,N_2073,N_2027);
nor U2549 (N_2549,N_2082,N_2058);
or U2550 (N_2550,N_1542,N_2226);
nor U2551 (N_2551,N_1789,N_1882);
nand U2552 (N_2552,N_2134,N_1611);
or U2553 (N_2553,N_1778,N_1974);
and U2554 (N_2554,N_2233,N_1918);
and U2555 (N_2555,N_1516,N_1938);
or U2556 (N_2556,N_1607,N_2140);
and U2557 (N_2557,N_2090,N_1549);
nor U2558 (N_2558,N_1795,N_2085);
nor U2559 (N_2559,N_1827,N_2114);
xnor U2560 (N_2560,N_1841,N_1514);
nor U2561 (N_2561,N_2147,N_1629);
or U2562 (N_2562,N_2002,N_1939);
nand U2563 (N_2563,N_2103,N_2051);
and U2564 (N_2564,N_1947,N_1758);
and U2565 (N_2565,N_1522,N_1660);
nor U2566 (N_2566,N_1916,N_1749);
nand U2567 (N_2567,N_1689,N_1713);
nand U2568 (N_2568,N_1798,N_1686);
nor U2569 (N_2569,N_1585,N_2228);
and U2570 (N_2570,N_1874,N_2013);
or U2571 (N_2571,N_2187,N_2175);
xnor U2572 (N_2572,N_1955,N_1859);
nor U2573 (N_2573,N_1555,N_1894);
nor U2574 (N_2574,N_2207,N_1788);
nor U2575 (N_2575,N_1756,N_1995);
nand U2576 (N_2576,N_2018,N_1617);
and U2577 (N_2577,N_2216,N_1627);
nand U2578 (N_2578,N_2092,N_1576);
nor U2579 (N_2579,N_2003,N_1573);
nand U2580 (N_2580,N_2203,N_1590);
or U2581 (N_2581,N_1517,N_1912);
nand U2582 (N_2582,N_1848,N_2205);
nand U2583 (N_2583,N_1832,N_1883);
and U2584 (N_2584,N_1681,N_1849);
nand U2585 (N_2585,N_1515,N_2237);
nand U2586 (N_2586,N_1606,N_2130);
nand U2587 (N_2587,N_2234,N_1594);
or U2588 (N_2588,N_1523,N_2040);
or U2589 (N_2589,N_2212,N_1879);
nand U2590 (N_2590,N_1810,N_1653);
nor U2591 (N_2591,N_1822,N_1760);
nand U2592 (N_2592,N_1654,N_1613);
nand U2593 (N_2593,N_2065,N_1961);
nor U2594 (N_2594,N_1643,N_1648);
and U2595 (N_2595,N_1730,N_1926);
nand U2596 (N_2596,N_2101,N_2223);
nor U2597 (N_2597,N_2067,N_2192);
xnor U2598 (N_2598,N_1735,N_1940);
nor U2599 (N_2599,N_2181,N_1639);
nor U2600 (N_2600,N_1984,N_2161);
or U2601 (N_2601,N_1683,N_1504);
and U2602 (N_2602,N_2168,N_1929);
and U2603 (N_2603,N_1989,N_1644);
or U2604 (N_2604,N_2059,N_1664);
and U2605 (N_2605,N_2011,N_2070);
nand U2606 (N_2606,N_1709,N_2068);
and U2607 (N_2607,N_1780,N_1803);
and U2608 (N_2608,N_1508,N_1791);
nand U2609 (N_2609,N_1614,N_1855);
or U2610 (N_2610,N_2035,N_1914);
nor U2611 (N_2611,N_2016,N_2037);
nand U2612 (N_2612,N_1588,N_1911);
nand U2613 (N_2613,N_1767,N_1564);
and U2614 (N_2614,N_1904,N_2000);
or U2615 (N_2615,N_1869,N_2244);
xnor U2616 (N_2616,N_2088,N_1716);
nor U2617 (N_2617,N_1870,N_1608);
and U2618 (N_2618,N_2172,N_1900);
xor U2619 (N_2619,N_1842,N_2005);
or U2620 (N_2620,N_1662,N_1727);
nand U2621 (N_2621,N_2049,N_1663);
and U2622 (N_2622,N_1597,N_1518);
and U2623 (N_2623,N_2235,N_2153);
nor U2624 (N_2624,N_1721,N_1598);
nand U2625 (N_2625,N_1991,N_1868);
or U2626 (N_2626,N_1798,N_2037);
nand U2627 (N_2627,N_1568,N_1647);
nand U2628 (N_2628,N_1911,N_1528);
nand U2629 (N_2629,N_1561,N_2003);
and U2630 (N_2630,N_2025,N_2223);
or U2631 (N_2631,N_2112,N_1564);
nor U2632 (N_2632,N_1919,N_1577);
nor U2633 (N_2633,N_1863,N_2063);
nor U2634 (N_2634,N_1746,N_1825);
or U2635 (N_2635,N_1785,N_1524);
and U2636 (N_2636,N_1753,N_1741);
nor U2637 (N_2637,N_1582,N_1681);
nand U2638 (N_2638,N_1684,N_2071);
nand U2639 (N_2639,N_1848,N_1928);
xor U2640 (N_2640,N_2191,N_1993);
nand U2641 (N_2641,N_2119,N_1523);
nand U2642 (N_2642,N_2046,N_1979);
or U2643 (N_2643,N_1572,N_1559);
nand U2644 (N_2644,N_1905,N_1810);
and U2645 (N_2645,N_2060,N_1727);
nor U2646 (N_2646,N_1637,N_2071);
and U2647 (N_2647,N_2143,N_1851);
and U2648 (N_2648,N_1846,N_1609);
and U2649 (N_2649,N_1621,N_2114);
or U2650 (N_2650,N_1923,N_1667);
nor U2651 (N_2651,N_1626,N_1595);
and U2652 (N_2652,N_1525,N_1569);
or U2653 (N_2653,N_1772,N_1809);
or U2654 (N_2654,N_2027,N_2144);
nor U2655 (N_2655,N_2050,N_2108);
and U2656 (N_2656,N_1515,N_1897);
nand U2657 (N_2657,N_1650,N_1573);
nand U2658 (N_2658,N_1647,N_1585);
nor U2659 (N_2659,N_1820,N_1990);
and U2660 (N_2660,N_1564,N_1899);
nor U2661 (N_2661,N_1895,N_2050);
nand U2662 (N_2662,N_1597,N_1715);
nor U2663 (N_2663,N_2131,N_1600);
nor U2664 (N_2664,N_1952,N_1616);
xnor U2665 (N_2665,N_1761,N_1776);
and U2666 (N_2666,N_1924,N_2112);
or U2667 (N_2667,N_2077,N_1872);
nor U2668 (N_2668,N_1536,N_1767);
and U2669 (N_2669,N_1997,N_1643);
or U2670 (N_2670,N_1946,N_1510);
or U2671 (N_2671,N_1593,N_1928);
and U2672 (N_2672,N_1814,N_1860);
and U2673 (N_2673,N_1625,N_1842);
and U2674 (N_2674,N_1569,N_1561);
nand U2675 (N_2675,N_1936,N_2234);
nor U2676 (N_2676,N_1997,N_2156);
or U2677 (N_2677,N_2185,N_1828);
and U2678 (N_2678,N_2081,N_1997);
nor U2679 (N_2679,N_1526,N_1775);
and U2680 (N_2680,N_1822,N_2156);
and U2681 (N_2681,N_2189,N_2159);
nand U2682 (N_2682,N_2034,N_1942);
nand U2683 (N_2683,N_1913,N_1535);
nor U2684 (N_2684,N_1634,N_1670);
nand U2685 (N_2685,N_2239,N_1661);
nand U2686 (N_2686,N_2045,N_1616);
nand U2687 (N_2687,N_2161,N_1805);
nor U2688 (N_2688,N_1870,N_2012);
or U2689 (N_2689,N_2131,N_1942);
or U2690 (N_2690,N_1709,N_2226);
nor U2691 (N_2691,N_1927,N_1869);
nor U2692 (N_2692,N_2221,N_1883);
nand U2693 (N_2693,N_1690,N_1697);
and U2694 (N_2694,N_2200,N_1884);
nand U2695 (N_2695,N_1699,N_1598);
nor U2696 (N_2696,N_1754,N_2144);
and U2697 (N_2697,N_2112,N_2123);
and U2698 (N_2698,N_2216,N_1653);
or U2699 (N_2699,N_2189,N_1676);
nor U2700 (N_2700,N_2038,N_2124);
nand U2701 (N_2701,N_1732,N_2243);
or U2702 (N_2702,N_1641,N_2105);
and U2703 (N_2703,N_1878,N_1698);
nand U2704 (N_2704,N_1888,N_1706);
nor U2705 (N_2705,N_2156,N_2111);
or U2706 (N_2706,N_2224,N_2036);
nor U2707 (N_2707,N_1915,N_1914);
and U2708 (N_2708,N_2183,N_1863);
and U2709 (N_2709,N_2012,N_2102);
and U2710 (N_2710,N_1597,N_1737);
nand U2711 (N_2711,N_2024,N_2087);
or U2712 (N_2712,N_1540,N_2008);
nor U2713 (N_2713,N_1802,N_1952);
and U2714 (N_2714,N_1549,N_1917);
nor U2715 (N_2715,N_1701,N_2156);
nand U2716 (N_2716,N_1601,N_1710);
nand U2717 (N_2717,N_1512,N_1693);
nand U2718 (N_2718,N_2069,N_2037);
or U2719 (N_2719,N_1973,N_1590);
nor U2720 (N_2720,N_1918,N_1832);
nor U2721 (N_2721,N_2048,N_1573);
and U2722 (N_2722,N_1952,N_1956);
nand U2723 (N_2723,N_1587,N_1545);
or U2724 (N_2724,N_2150,N_1603);
or U2725 (N_2725,N_2201,N_1767);
nor U2726 (N_2726,N_2032,N_1603);
nor U2727 (N_2727,N_2244,N_2127);
nor U2728 (N_2728,N_1587,N_1525);
nand U2729 (N_2729,N_1703,N_1543);
and U2730 (N_2730,N_1909,N_2226);
nor U2731 (N_2731,N_1768,N_1733);
and U2732 (N_2732,N_1601,N_1645);
nor U2733 (N_2733,N_1561,N_2133);
nor U2734 (N_2734,N_2241,N_1616);
nor U2735 (N_2735,N_1501,N_1928);
nand U2736 (N_2736,N_1675,N_1721);
and U2737 (N_2737,N_1858,N_1905);
and U2738 (N_2738,N_2015,N_1828);
and U2739 (N_2739,N_1516,N_2241);
nand U2740 (N_2740,N_2086,N_1747);
nor U2741 (N_2741,N_1655,N_1735);
nand U2742 (N_2742,N_1607,N_1670);
or U2743 (N_2743,N_2046,N_1597);
xor U2744 (N_2744,N_2127,N_1880);
and U2745 (N_2745,N_1898,N_1978);
xnor U2746 (N_2746,N_1792,N_2241);
and U2747 (N_2747,N_2149,N_2157);
and U2748 (N_2748,N_1536,N_1772);
and U2749 (N_2749,N_2189,N_2109);
nand U2750 (N_2750,N_2181,N_1706);
nor U2751 (N_2751,N_1615,N_1668);
nand U2752 (N_2752,N_1687,N_1910);
xnor U2753 (N_2753,N_1856,N_2248);
and U2754 (N_2754,N_1601,N_1594);
and U2755 (N_2755,N_1841,N_2233);
nand U2756 (N_2756,N_1737,N_2013);
nand U2757 (N_2757,N_1624,N_2036);
or U2758 (N_2758,N_1592,N_2090);
or U2759 (N_2759,N_2239,N_1534);
nand U2760 (N_2760,N_1996,N_2229);
or U2761 (N_2761,N_1933,N_1600);
nand U2762 (N_2762,N_1915,N_2053);
nand U2763 (N_2763,N_1515,N_2204);
nand U2764 (N_2764,N_1611,N_2204);
xor U2765 (N_2765,N_1819,N_2112);
or U2766 (N_2766,N_1886,N_2062);
or U2767 (N_2767,N_1836,N_2107);
and U2768 (N_2768,N_1797,N_2106);
or U2769 (N_2769,N_2109,N_1575);
nor U2770 (N_2770,N_2206,N_1617);
nand U2771 (N_2771,N_1627,N_1652);
and U2772 (N_2772,N_1556,N_1975);
or U2773 (N_2773,N_1733,N_2168);
nor U2774 (N_2774,N_2108,N_1609);
nor U2775 (N_2775,N_2009,N_1627);
or U2776 (N_2776,N_1808,N_1510);
and U2777 (N_2777,N_1875,N_2143);
nand U2778 (N_2778,N_2009,N_2190);
or U2779 (N_2779,N_1599,N_1979);
nand U2780 (N_2780,N_2220,N_1862);
and U2781 (N_2781,N_1932,N_1769);
and U2782 (N_2782,N_1634,N_1814);
nor U2783 (N_2783,N_1669,N_1757);
and U2784 (N_2784,N_1790,N_1930);
nand U2785 (N_2785,N_1596,N_1740);
and U2786 (N_2786,N_1895,N_1622);
or U2787 (N_2787,N_1550,N_1707);
nand U2788 (N_2788,N_2119,N_2189);
nor U2789 (N_2789,N_2077,N_1612);
and U2790 (N_2790,N_1809,N_1603);
and U2791 (N_2791,N_2059,N_1660);
or U2792 (N_2792,N_1544,N_1547);
nand U2793 (N_2793,N_2232,N_2111);
nor U2794 (N_2794,N_2164,N_2020);
nor U2795 (N_2795,N_1623,N_1715);
nor U2796 (N_2796,N_1926,N_1991);
and U2797 (N_2797,N_1894,N_1576);
and U2798 (N_2798,N_1511,N_2146);
or U2799 (N_2799,N_1700,N_1587);
nand U2800 (N_2800,N_1529,N_1722);
or U2801 (N_2801,N_1756,N_1626);
and U2802 (N_2802,N_1568,N_1807);
nand U2803 (N_2803,N_1581,N_1599);
and U2804 (N_2804,N_2091,N_1513);
nor U2805 (N_2805,N_2063,N_1759);
nor U2806 (N_2806,N_2107,N_2090);
nand U2807 (N_2807,N_2069,N_2096);
nand U2808 (N_2808,N_1574,N_2226);
or U2809 (N_2809,N_1994,N_1747);
nor U2810 (N_2810,N_1861,N_2203);
nand U2811 (N_2811,N_2011,N_2205);
nor U2812 (N_2812,N_1869,N_1696);
and U2813 (N_2813,N_2088,N_1987);
nor U2814 (N_2814,N_1528,N_2133);
nor U2815 (N_2815,N_2080,N_2099);
and U2816 (N_2816,N_2162,N_2059);
nand U2817 (N_2817,N_1969,N_1922);
or U2818 (N_2818,N_2249,N_2102);
or U2819 (N_2819,N_1719,N_2131);
or U2820 (N_2820,N_2124,N_1656);
nand U2821 (N_2821,N_1945,N_2152);
or U2822 (N_2822,N_1551,N_1857);
or U2823 (N_2823,N_1785,N_1841);
or U2824 (N_2824,N_1519,N_1773);
nor U2825 (N_2825,N_1661,N_1691);
nor U2826 (N_2826,N_1895,N_1621);
nor U2827 (N_2827,N_1622,N_1604);
nand U2828 (N_2828,N_1691,N_1837);
nand U2829 (N_2829,N_2078,N_1828);
or U2830 (N_2830,N_1533,N_2096);
and U2831 (N_2831,N_1694,N_1991);
or U2832 (N_2832,N_1800,N_2157);
nand U2833 (N_2833,N_1778,N_1927);
or U2834 (N_2834,N_1799,N_1939);
or U2835 (N_2835,N_2188,N_1658);
nor U2836 (N_2836,N_1571,N_1579);
nor U2837 (N_2837,N_1898,N_1581);
and U2838 (N_2838,N_1868,N_1766);
nor U2839 (N_2839,N_1714,N_1534);
nor U2840 (N_2840,N_2032,N_1538);
nand U2841 (N_2841,N_1640,N_2060);
nor U2842 (N_2842,N_1504,N_1509);
nor U2843 (N_2843,N_2077,N_1632);
nor U2844 (N_2844,N_1794,N_2231);
and U2845 (N_2845,N_1842,N_1948);
or U2846 (N_2846,N_2081,N_1781);
and U2847 (N_2847,N_1729,N_1935);
nand U2848 (N_2848,N_1815,N_1893);
and U2849 (N_2849,N_1687,N_2049);
nor U2850 (N_2850,N_1665,N_1870);
nand U2851 (N_2851,N_1702,N_2225);
nand U2852 (N_2852,N_1643,N_2033);
nand U2853 (N_2853,N_2109,N_2183);
nand U2854 (N_2854,N_1948,N_1631);
xnor U2855 (N_2855,N_1702,N_1603);
or U2856 (N_2856,N_1935,N_1809);
nand U2857 (N_2857,N_1832,N_1624);
nor U2858 (N_2858,N_1978,N_2073);
nor U2859 (N_2859,N_1647,N_1622);
nand U2860 (N_2860,N_1564,N_1974);
and U2861 (N_2861,N_1732,N_2207);
and U2862 (N_2862,N_2175,N_1667);
nor U2863 (N_2863,N_2155,N_1547);
nand U2864 (N_2864,N_1876,N_2027);
nand U2865 (N_2865,N_1845,N_1957);
or U2866 (N_2866,N_1637,N_1902);
or U2867 (N_2867,N_2108,N_2179);
nand U2868 (N_2868,N_1825,N_1791);
nor U2869 (N_2869,N_1569,N_1709);
and U2870 (N_2870,N_2081,N_1802);
and U2871 (N_2871,N_2235,N_2168);
and U2872 (N_2872,N_2132,N_2026);
and U2873 (N_2873,N_1843,N_1916);
and U2874 (N_2874,N_1608,N_1702);
and U2875 (N_2875,N_1691,N_1922);
and U2876 (N_2876,N_2212,N_1986);
nor U2877 (N_2877,N_2176,N_1523);
nor U2878 (N_2878,N_1517,N_1855);
or U2879 (N_2879,N_2161,N_2135);
nor U2880 (N_2880,N_1783,N_1631);
nor U2881 (N_2881,N_1898,N_1539);
nor U2882 (N_2882,N_1577,N_1722);
nor U2883 (N_2883,N_1691,N_2103);
or U2884 (N_2884,N_1662,N_2058);
nand U2885 (N_2885,N_2080,N_2150);
nor U2886 (N_2886,N_1606,N_1648);
and U2887 (N_2887,N_1985,N_1664);
nor U2888 (N_2888,N_1757,N_2202);
or U2889 (N_2889,N_1815,N_1611);
nand U2890 (N_2890,N_1623,N_1910);
nand U2891 (N_2891,N_2042,N_1558);
nor U2892 (N_2892,N_2081,N_1731);
or U2893 (N_2893,N_1634,N_1898);
nor U2894 (N_2894,N_1942,N_1517);
nor U2895 (N_2895,N_1986,N_1525);
nand U2896 (N_2896,N_2063,N_1944);
nand U2897 (N_2897,N_1939,N_1789);
and U2898 (N_2898,N_1942,N_1725);
or U2899 (N_2899,N_1619,N_1868);
and U2900 (N_2900,N_1936,N_2123);
nor U2901 (N_2901,N_1827,N_2022);
nor U2902 (N_2902,N_1867,N_2152);
and U2903 (N_2903,N_2086,N_2117);
and U2904 (N_2904,N_2131,N_1604);
and U2905 (N_2905,N_1805,N_1817);
nor U2906 (N_2906,N_1922,N_1835);
or U2907 (N_2907,N_1524,N_1819);
or U2908 (N_2908,N_1769,N_1856);
nor U2909 (N_2909,N_1630,N_1520);
nand U2910 (N_2910,N_2038,N_2081);
or U2911 (N_2911,N_1908,N_2035);
nor U2912 (N_2912,N_2166,N_1838);
or U2913 (N_2913,N_2066,N_1737);
nand U2914 (N_2914,N_1644,N_2151);
nand U2915 (N_2915,N_2163,N_1708);
or U2916 (N_2916,N_2016,N_1912);
or U2917 (N_2917,N_1511,N_1765);
and U2918 (N_2918,N_2142,N_1970);
nand U2919 (N_2919,N_1984,N_2035);
and U2920 (N_2920,N_1710,N_1629);
and U2921 (N_2921,N_1884,N_1640);
or U2922 (N_2922,N_2042,N_2142);
nor U2923 (N_2923,N_1757,N_1520);
nand U2924 (N_2924,N_1585,N_1809);
nor U2925 (N_2925,N_2155,N_1791);
xor U2926 (N_2926,N_1923,N_1798);
or U2927 (N_2927,N_2139,N_2091);
nor U2928 (N_2928,N_2231,N_1634);
nand U2929 (N_2929,N_2089,N_1852);
and U2930 (N_2930,N_1975,N_2018);
nand U2931 (N_2931,N_1716,N_1893);
xnor U2932 (N_2932,N_1786,N_1931);
and U2933 (N_2933,N_1606,N_1549);
nand U2934 (N_2934,N_2123,N_1501);
or U2935 (N_2935,N_1590,N_1697);
nand U2936 (N_2936,N_2165,N_2098);
nand U2937 (N_2937,N_2074,N_1740);
nand U2938 (N_2938,N_1951,N_1786);
or U2939 (N_2939,N_1702,N_1971);
and U2940 (N_2940,N_1544,N_2151);
and U2941 (N_2941,N_1617,N_1916);
or U2942 (N_2942,N_2111,N_2102);
and U2943 (N_2943,N_2115,N_2060);
or U2944 (N_2944,N_1563,N_1554);
nor U2945 (N_2945,N_1695,N_1789);
or U2946 (N_2946,N_1536,N_1944);
nor U2947 (N_2947,N_2054,N_1677);
nand U2948 (N_2948,N_2218,N_2191);
nor U2949 (N_2949,N_1983,N_1756);
nand U2950 (N_2950,N_1594,N_1745);
nor U2951 (N_2951,N_1852,N_1645);
or U2952 (N_2952,N_2071,N_2203);
or U2953 (N_2953,N_2139,N_1589);
and U2954 (N_2954,N_1659,N_1839);
or U2955 (N_2955,N_2081,N_1563);
nand U2956 (N_2956,N_2193,N_1815);
nand U2957 (N_2957,N_1785,N_1727);
or U2958 (N_2958,N_2198,N_1747);
or U2959 (N_2959,N_1663,N_1775);
nor U2960 (N_2960,N_1778,N_1918);
and U2961 (N_2961,N_2042,N_2202);
nor U2962 (N_2962,N_2076,N_1810);
or U2963 (N_2963,N_1564,N_1814);
and U2964 (N_2964,N_1796,N_1726);
xor U2965 (N_2965,N_2107,N_2144);
nand U2966 (N_2966,N_1529,N_1543);
or U2967 (N_2967,N_1594,N_1951);
or U2968 (N_2968,N_2244,N_1737);
nand U2969 (N_2969,N_2025,N_2019);
nand U2970 (N_2970,N_2159,N_1504);
nand U2971 (N_2971,N_1508,N_1855);
nand U2972 (N_2972,N_2001,N_1946);
or U2973 (N_2973,N_1777,N_1686);
nor U2974 (N_2974,N_2160,N_1636);
nand U2975 (N_2975,N_2238,N_1929);
xnor U2976 (N_2976,N_1929,N_1896);
nand U2977 (N_2977,N_2196,N_2155);
nand U2978 (N_2978,N_2161,N_1853);
or U2979 (N_2979,N_1664,N_1876);
nor U2980 (N_2980,N_1526,N_1906);
and U2981 (N_2981,N_1674,N_2132);
nor U2982 (N_2982,N_1854,N_1509);
or U2983 (N_2983,N_1837,N_2000);
or U2984 (N_2984,N_1631,N_1630);
or U2985 (N_2985,N_2145,N_1660);
nand U2986 (N_2986,N_1601,N_1637);
or U2987 (N_2987,N_1835,N_1955);
nor U2988 (N_2988,N_1671,N_2085);
or U2989 (N_2989,N_1783,N_1829);
nand U2990 (N_2990,N_2240,N_1877);
nand U2991 (N_2991,N_1892,N_1702);
nor U2992 (N_2992,N_2038,N_1734);
nand U2993 (N_2993,N_1920,N_2070);
nand U2994 (N_2994,N_1794,N_2014);
nand U2995 (N_2995,N_1522,N_2084);
nand U2996 (N_2996,N_1729,N_2029);
nand U2997 (N_2997,N_1653,N_1999);
and U2998 (N_2998,N_1797,N_1544);
and U2999 (N_2999,N_1903,N_2204);
and UO_0 (O_0,N_2839,N_2554);
or UO_1 (O_1,N_2685,N_2584);
nor UO_2 (O_2,N_2760,N_2336);
nor UO_3 (O_3,N_2774,N_2759);
nor UO_4 (O_4,N_2934,N_2904);
nand UO_5 (O_5,N_2855,N_2930);
xor UO_6 (O_6,N_2828,N_2507);
and UO_7 (O_7,N_2258,N_2427);
nand UO_8 (O_8,N_2426,N_2923);
or UO_9 (O_9,N_2947,N_2681);
nor UO_10 (O_10,N_2732,N_2827);
and UO_11 (O_11,N_2561,N_2946);
nand UO_12 (O_12,N_2562,N_2739);
and UO_13 (O_13,N_2656,N_2603);
and UO_14 (O_14,N_2495,N_2919);
nor UO_15 (O_15,N_2910,N_2675);
or UO_16 (O_16,N_2830,N_2566);
and UO_17 (O_17,N_2880,N_2349);
nor UO_18 (O_18,N_2465,N_2509);
nand UO_19 (O_19,N_2678,N_2911);
and UO_20 (O_20,N_2390,N_2639);
and UO_21 (O_21,N_2963,N_2458);
and UO_22 (O_22,N_2474,N_2416);
and UO_23 (O_23,N_2557,N_2850);
nor UO_24 (O_24,N_2403,N_2446);
and UO_25 (O_25,N_2411,N_2410);
or UO_26 (O_26,N_2303,N_2327);
and UO_27 (O_27,N_2516,N_2255);
xnor UO_28 (O_28,N_2280,N_2356);
and UO_29 (O_29,N_2782,N_2973);
nor UO_30 (O_30,N_2553,N_2482);
or UO_31 (O_31,N_2877,N_2582);
and UO_32 (O_32,N_2740,N_2938);
and UO_33 (O_33,N_2615,N_2799);
nand UO_34 (O_34,N_2648,N_2695);
or UO_35 (O_35,N_2837,N_2472);
nand UO_36 (O_36,N_2369,N_2770);
nand UO_37 (O_37,N_2409,N_2951);
or UO_38 (O_38,N_2699,N_2662);
or UO_39 (O_39,N_2252,N_2490);
nand UO_40 (O_40,N_2568,N_2835);
nor UO_41 (O_41,N_2622,N_2560);
nand UO_42 (O_42,N_2676,N_2667);
nor UO_43 (O_43,N_2275,N_2831);
and UO_44 (O_44,N_2351,N_2338);
or UO_45 (O_45,N_2840,N_2539);
xor UO_46 (O_46,N_2371,N_2790);
or UO_47 (O_47,N_2886,N_2479);
nand UO_48 (O_48,N_2316,N_2592);
nand UO_49 (O_49,N_2632,N_2926);
and UO_50 (O_50,N_2550,N_2786);
or UO_51 (O_51,N_2612,N_2892);
or UO_52 (O_52,N_2305,N_2956);
or UO_53 (O_53,N_2538,N_2521);
and UO_54 (O_54,N_2888,N_2979);
nor UO_55 (O_55,N_2254,N_2259);
or UO_56 (O_56,N_2391,N_2668);
or UO_57 (O_57,N_2251,N_2396);
nor UO_58 (O_58,N_2948,N_2337);
xnor UO_59 (O_59,N_2765,N_2727);
nor UO_60 (O_60,N_2298,N_2986);
nor UO_61 (O_61,N_2464,N_2436);
nand UO_62 (O_62,N_2621,N_2975);
nor UO_63 (O_63,N_2704,N_2581);
nand UO_64 (O_64,N_2440,N_2586);
nor UO_65 (O_65,N_2310,N_2463);
nand UO_66 (O_66,N_2354,N_2763);
or UO_67 (O_67,N_2385,N_2984);
nor UO_68 (O_68,N_2449,N_2265);
nor UO_69 (O_69,N_2494,N_2319);
or UO_70 (O_70,N_2949,N_2715);
and UO_71 (O_71,N_2833,N_2994);
xor UO_72 (O_72,N_2536,N_2412);
and UO_73 (O_73,N_2646,N_2891);
and UO_74 (O_74,N_2279,N_2829);
or UO_75 (O_75,N_2483,N_2708);
nand UO_76 (O_76,N_2944,N_2964);
and UO_77 (O_77,N_2459,N_2764);
nor UO_78 (O_78,N_2524,N_2519);
nor UO_79 (O_79,N_2296,N_2787);
and UO_80 (O_80,N_2709,N_2659);
and UO_81 (O_81,N_2991,N_2533);
nand UO_82 (O_82,N_2617,N_2600);
nand UO_83 (O_83,N_2731,N_2977);
or UO_84 (O_84,N_2375,N_2299);
and UO_85 (O_85,N_2711,N_2522);
and UO_86 (O_86,N_2278,N_2544);
nand UO_87 (O_87,N_2578,N_2547);
or UO_88 (O_88,N_2325,N_2362);
nand UO_89 (O_89,N_2384,N_2901);
and UO_90 (O_90,N_2377,N_2443);
nor UO_91 (O_91,N_2328,N_2771);
and UO_92 (O_92,N_2344,N_2959);
nor UO_93 (O_93,N_2329,N_2801);
and UO_94 (O_94,N_2331,N_2957);
nand UO_95 (O_95,N_2271,N_2781);
nand UO_96 (O_96,N_2323,N_2549);
or UO_97 (O_97,N_2373,N_2276);
or UO_98 (O_98,N_2398,N_2756);
and UO_99 (O_99,N_2969,N_2990);
and UO_100 (O_100,N_2431,N_2253);
and UO_101 (O_101,N_2473,N_2574);
nand UO_102 (O_102,N_2264,N_2625);
nand UO_103 (O_103,N_2419,N_2348);
nand UO_104 (O_104,N_2691,N_2650);
nand UO_105 (O_105,N_2793,N_2707);
nor UO_106 (O_106,N_2909,N_2618);
or UO_107 (O_107,N_2942,N_2623);
and UO_108 (O_108,N_2908,N_2274);
nand UO_109 (O_109,N_2841,N_2383);
and UO_110 (O_110,N_2388,N_2597);
and UO_111 (O_111,N_2652,N_2526);
nand UO_112 (O_112,N_2752,N_2713);
nor UO_113 (O_113,N_2614,N_2960);
or UO_114 (O_114,N_2847,N_2610);
or UO_115 (O_115,N_2882,N_2601);
nor UO_116 (O_116,N_2360,N_2821);
nor UO_117 (O_117,N_2370,N_2480);
or UO_118 (O_118,N_2637,N_2414);
and UO_119 (O_119,N_2397,N_2726);
nand UO_120 (O_120,N_2696,N_2497);
nand UO_121 (O_121,N_2394,N_2689);
or UO_122 (O_122,N_2380,N_2750);
and UO_123 (O_123,N_2687,N_2269);
nand UO_124 (O_124,N_2697,N_2309);
nor UO_125 (O_125,N_2736,N_2452);
nand UO_126 (O_126,N_2506,N_2293);
nor UO_127 (O_127,N_2813,N_2435);
or UO_128 (O_128,N_2364,N_2492);
and UO_129 (O_129,N_2834,N_2466);
nor UO_130 (O_130,N_2643,N_2366);
nor UO_131 (O_131,N_2609,N_2447);
nand UO_132 (O_132,N_2552,N_2635);
nand UO_133 (O_133,N_2422,N_2745);
nor UO_134 (O_134,N_2250,N_2467);
nand UO_135 (O_135,N_2588,N_2896);
or UO_136 (O_136,N_2415,N_2683);
nor UO_137 (O_137,N_2933,N_2393);
nand UO_138 (O_138,N_2499,N_2401);
nor UO_139 (O_139,N_2496,N_2718);
or UO_140 (O_140,N_2912,N_2461);
or UO_141 (O_141,N_2503,N_2429);
or UO_142 (O_142,N_2334,N_2619);
nor UO_143 (O_143,N_2758,N_2874);
nand UO_144 (O_144,N_2903,N_2789);
or UO_145 (O_145,N_2970,N_2669);
or UO_146 (O_146,N_2961,N_2796);
nand UO_147 (O_147,N_2502,N_2742);
nand UO_148 (O_148,N_2780,N_2545);
nor UO_149 (O_149,N_2379,N_2674);
or UO_150 (O_150,N_2939,N_2535);
and UO_151 (O_151,N_2686,N_2700);
nor UO_152 (O_152,N_2872,N_2641);
or UO_153 (O_153,N_2341,N_2701);
or UO_154 (O_154,N_2857,N_2551);
or UO_155 (O_155,N_2894,N_2433);
nand UO_156 (O_156,N_2866,N_2854);
and UO_157 (O_157,N_2491,N_2462);
nand UO_158 (O_158,N_2734,N_2856);
or UO_159 (O_159,N_2649,N_2315);
and UO_160 (O_160,N_2442,N_2844);
or UO_161 (O_161,N_2907,N_2300);
nor UO_162 (O_162,N_2607,N_2591);
nor UO_163 (O_163,N_2605,N_2543);
nor UO_164 (O_164,N_2693,N_2540);
and UO_165 (O_165,N_2382,N_2753);
nor UO_166 (O_166,N_2558,N_2378);
nor UO_167 (O_167,N_2457,N_2852);
or UO_168 (O_168,N_2940,N_2478);
nand UO_169 (O_169,N_2846,N_2826);
or UO_170 (O_170,N_2735,N_2883);
nand UO_171 (O_171,N_2339,N_2313);
nor UO_172 (O_172,N_2448,N_2914);
or UO_173 (O_173,N_2613,N_2717);
nor UO_174 (O_174,N_2372,N_2776);
nor UO_175 (O_175,N_2363,N_2399);
nor UO_176 (O_176,N_2738,N_2406);
and UO_177 (O_177,N_2998,N_2895);
and UO_178 (O_178,N_2809,N_2873);
nor UO_179 (O_179,N_2598,N_2918);
nand UO_180 (O_180,N_2794,N_2484);
or UO_181 (O_181,N_2863,N_2505);
nand UO_182 (O_182,N_2631,N_2783);
and UO_183 (O_183,N_2875,N_2858);
nor UO_184 (O_184,N_2749,N_2455);
nor UO_185 (O_185,N_2468,N_2630);
or UO_186 (O_186,N_2870,N_2283);
or UO_187 (O_187,N_2860,N_2477);
or UO_188 (O_188,N_2267,N_2945);
nor UO_189 (O_189,N_2817,N_2470);
nand UO_190 (O_190,N_2306,N_2571);
nor UO_191 (O_191,N_2282,N_2802);
or UO_192 (O_192,N_2332,N_2376);
nor UO_193 (O_193,N_2546,N_2666);
nand UO_194 (O_194,N_2583,N_2260);
and UO_195 (O_195,N_2869,N_2511);
xnor UO_196 (O_196,N_2359,N_2292);
and UO_197 (O_197,N_2564,N_2823);
nor UO_198 (O_198,N_2723,N_2672);
and UO_199 (O_199,N_2653,N_2485);
or UO_200 (O_200,N_2798,N_2616);
and UO_201 (O_201,N_2285,N_2811);
nor UO_202 (O_202,N_2537,N_2413);
and UO_203 (O_203,N_2922,N_2510);
and UO_204 (O_204,N_2476,N_2532);
nor UO_205 (O_205,N_2889,N_2899);
nor UO_206 (O_206,N_2848,N_2647);
or UO_207 (O_207,N_2952,N_2885);
or UO_208 (O_208,N_2772,N_2761);
nor UO_209 (O_209,N_2287,N_2663);
nor UO_210 (O_210,N_2716,N_2743);
or UO_211 (O_211,N_2580,N_2441);
and UO_212 (O_212,N_2575,N_2859);
and UO_213 (O_213,N_2714,N_2682);
nor UO_214 (O_214,N_2651,N_2270);
nor UO_215 (O_215,N_2967,N_2958);
or UO_216 (O_216,N_2974,N_2818);
or UO_217 (O_217,N_2881,N_2679);
or UO_218 (O_218,N_2773,N_2816);
or UO_219 (O_219,N_2488,N_2905);
and UO_220 (O_220,N_2788,N_2897);
and UO_221 (O_221,N_2996,N_2262);
nand UO_222 (O_222,N_2450,N_2744);
nor UO_223 (O_223,N_2527,N_2481);
or UO_224 (O_224,N_2321,N_2767);
nand UO_225 (O_225,N_2966,N_2797);
nand UO_226 (O_226,N_2965,N_2565);
or UO_227 (O_227,N_2531,N_2792);
nand UO_228 (O_228,N_2754,N_2902);
nor UO_229 (O_229,N_2981,N_2320);
and UO_230 (O_230,N_2627,N_2638);
xnor UO_231 (O_231,N_2314,N_2824);
nand UO_232 (O_232,N_2365,N_2710);
nand UO_233 (O_233,N_2748,N_2555);
nand UO_234 (O_234,N_2322,N_2324);
nand UO_235 (O_235,N_2290,N_2460);
xor UO_236 (O_236,N_2628,N_2421);
nand UO_237 (O_237,N_2864,N_2405);
nand UO_238 (O_238,N_2921,N_2453);
or UO_239 (O_239,N_2528,N_2281);
nand UO_240 (O_240,N_2418,N_2862);
or UO_241 (O_241,N_2924,N_2836);
nor UO_242 (O_242,N_2705,N_2311);
nand UO_243 (O_243,N_2645,N_2268);
nand UO_244 (O_244,N_2815,N_2346);
nor UO_245 (O_245,N_2876,N_2728);
nand UO_246 (O_246,N_2721,N_2680);
nand UO_247 (O_247,N_2301,N_2374);
xor UO_248 (O_248,N_2755,N_2719);
nor UO_249 (O_249,N_2400,N_2832);
nor UO_250 (O_250,N_2318,N_2444);
nor UO_251 (O_251,N_2791,N_2567);
and UO_252 (O_252,N_2640,N_2887);
nand UO_253 (O_253,N_2636,N_2517);
nor UO_254 (O_254,N_2992,N_2983);
nor UO_255 (O_255,N_2579,N_2347);
nor UO_256 (O_256,N_2746,N_2404);
nand UO_257 (O_257,N_2670,N_2518);
nor UO_258 (O_258,N_2694,N_2294);
or UO_259 (O_259,N_2692,N_2751);
and UO_260 (O_260,N_2703,N_2784);
nand UO_261 (O_261,N_2730,N_2954);
nor UO_262 (O_262,N_2928,N_2775);
and UO_263 (O_263,N_2658,N_2589);
nand UO_264 (O_264,N_2424,N_2330);
or UO_265 (O_265,N_2548,N_2995);
and UO_266 (O_266,N_2387,N_2563);
and UO_267 (O_267,N_2778,N_2962);
or UO_268 (O_268,N_2993,N_2684);
and UO_269 (O_269,N_2420,N_2810);
or UO_270 (O_270,N_2438,N_2489);
nor UO_271 (O_271,N_2512,N_2395);
or UO_272 (O_272,N_2849,N_2900);
or UO_273 (O_273,N_2808,N_2871);
xor UO_274 (O_274,N_2498,N_2985);
or UO_275 (O_275,N_2368,N_2820);
nor UO_276 (O_276,N_2381,N_2915);
and UO_277 (O_277,N_2596,N_2757);
nand UO_278 (O_278,N_2814,N_2988);
and UO_279 (O_279,N_2302,N_2392);
or UO_280 (O_280,N_2577,N_2762);
nand UO_281 (O_281,N_2277,N_2724);
nor UO_282 (O_282,N_2657,N_2291);
nor UO_283 (O_283,N_2978,N_2980);
nor UO_284 (O_284,N_2295,N_2769);
nor UO_285 (O_285,N_2853,N_2602);
nor UO_286 (O_286,N_2432,N_2916);
and UO_287 (O_287,N_2576,N_2456);
or UO_288 (O_288,N_2599,N_2932);
nand UO_289 (O_289,N_2943,N_2297);
nand UO_290 (O_290,N_2508,N_2825);
nand UO_291 (O_291,N_2879,N_2304);
nand UO_292 (O_292,N_2971,N_2671);
and UO_293 (O_293,N_2272,N_2702);
or UO_294 (O_294,N_2935,N_2342);
or UO_295 (O_295,N_2690,N_2335);
and UO_296 (O_296,N_2941,N_2729);
or UO_297 (O_297,N_2286,N_2556);
and UO_298 (O_298,N_2804,N_2805);
nand UO_299 (O_299,N_2430,N_2608);
nand UO_300 (O_300,N_2661,N_2529);
and UO_301 (O_301,N_2785,N_2343);
and UO_302 (O_302,N_2606,N_2861);
and UO_303 (O_303,N_2737,N_2677);
nor UO_304 (O_304,N_2803,N_2634);
nor UO_305 (O_305,N_2806,N_2288);
and UO_306 (O_306,N_2523,N_2633);
or UO_307 (O_307,N_2722,N_2644);
nand UO_308 (O_308,N_2843,N_2439);
nand UO_309 (O_309,N_2624,N_2307);
nor UO_310 (O_310,N_2819,N_2428);
nand UO_311 (O_311,N_2865,N_2587);
nor UO_312 (O_312,N_2720,N_2664);
nor UO_313 (O_313,N_2504,N_2987);
nor UO_314 (O_314,N_2357,N_2997);
nor UO_315 (O_315,N_2851,N_2263);
nor UO_316 (O_316,N_2929,N_2273);
nand UO_317 (O_317,N_2367,N_2515);
nand UO_318 (O_318,N_2266,N_2913);
nor UO_319 (O_319,N_2779,N_2595);
or UO_320 (O_320,N_2386,N_2358);
nand UO_321 (O_321,N_2890,N_2570);
nand UO_322 (O_322,N_2712,N_2402);
or UO_323 (O_323,N_2673,N_2345);
nand UO_324 (O_324,N_2698,N_2408);
xnor UO_325 (O_325,N_2868,N_2807);
or UO_326 (O_326,N_2256,N_2594);
and UO_327 (O_327,N_2471,N_2423);
or UO_328 (O_328,N_2654,N_2514);
nor UO_329 (O_329,N_2917,N_2741);
and UO_330 (O_330,N_2884,N_2620);
or UO_331 (O_331,N_2626,N_2454);
and UO_332 (O_332,N_2437,N_2572);
and UO_333 (O_333,N_2766,N_2257);
xnor UO_334 (O_334,N_2660,N_2326);
nor UO_335 (O_335,N_2800,N_2655);
nor UO_336 (O_336,N_2333,N_2534);
nand UO_337 (O_337,N_2573,N_2733);
nor UO_338 (O_338,N_2434,N_2469);
and UO_339 (O_339,N_2989,N_2340);
xor UO_340 (O_340,N_2352,N_2525);
nand UO_341 (O_341,N_2317,N_2665);
nor UO_342 (O_342,N_2593,N_2867);
and UO_343 (O_343,N_2604,N_2590);
nand UO_344 (O_344,N_2289,N_2936);
nand UO_345 (O_345,N_2768,N_2747);
nor UO_346 (O_346,N_2389,N_2999);
or UO_347 (O_347,N_2925,N_2611);
nand UO_348 (O_348,N_2451,N_2937);
nand UO_349 (O_349,N_2706,N_2355);
nor UO_350 (O_350,N_2878,N_2898);
nand UO_351 (O_351,N_2353,N_2893);
or UO_352 (O_352,N_2972,N_2425);
and UO_353 (O_353,N_2445,N_2688);
or UO_354 (O_354,N_2284,N_2795);
and UO_355 (O_355,N_2493,N_2725);
or UO_356 (O_356,N_2920,N_2976);
or UO_357 (O_357,N_2541,N_2312);
nor UO_358 (O_358,N_2842,N_2822);
nand UO_359 (O_359,N_2812,N_2530);
and UO_360 (O_360,N_2845,N_2906);
nand UO_361 (O_361,N_2931,N_2261);
and UO_362 (O_362,N_2642,N_2953);
nand UO_363 (O_363,N_2777,N_2982);
nand UO_364 (O_364,N_2501,N_2968);
or UO_365 (O_365,N_2487,N_2950);
nand UO_366 (O_366,N_2361,N_2513);
and UO_367 (O_367,N_2475,N_2585);
nand UO_368 (O_368,N_2417,N_2838);
nand UO_369 (O_369,N_2520,N_2308);
nand UO_370 (O_370,N_2927,N_2407);
xor UO_371 (O_371,N_2542,N_2955);
nor UO_372 (O_372,N_2486,N_2500);
or UO_373 (O_373,N_2350,N_2559);
nand UO_374 (O_374,N_2569,N_2629);
xor UO_375 (O_375,N_2680,N_2554);
and UO_376 (O_376,N_2520,N_2433);
nand UO_377 (O_377,N_2466,N_2399);
nand UO_378 (O_378,N_2592,N_2751);
nand UO_379 (O_379,N_2282,N_2517);
and UO_380 (O_380,N_2488,N_2335);
nor UO_381 (O_381,N_2941,N_2758);
and UO_382 (O_382,N_2467,N_2970);
or UO_383 (O_383,N_2583,N_2325);
nor UO_384 (O_384,N_2411,N_2835);
nand UO_385 (O_385,N_2521,N_2834);
and UO_386 (O_386,N_2889,N_2770);
or UO_387 (O_387,N_2871,N_2250);
and UO_388 (O_388,N_2310,N_2299);
and UO_389 (O_389,N_2460,N_2326);
nor UO_390 (O_390,N_2456,N_2847);
and UO_391 (O_391,N_2839,N_2551);
or UO_392 (O_392,N_2630,N_2401);
or UO_393 (O_393,N_2370,N_2951);
nor UO_394 (O_394,N_2818,N_2514);
or UO_395 (O_395,N_2736,N_2408);
xor UO_396 (O_396,N_2749,N_2853);
nand UO_397 (O_397,N_2991,N_2905);
nor UO_398 (O_398,N_2840,N_2527);
or UO_399 (O_399,N_2345,N_2744);
and UO_400 (O_400,N_2669,N_2792);
nor UO_401 (O_401,N_2405,N_2308);
nor UO_402 (O_402,N_2499,N_2882);
nand UO_403 (O_403,N_2325,N_2954);
nand UO_404 (O_404,N_2662,N_2265);
nand UO_405 (O_405,N_2555,N_2526);
and UO_406 (O_406,N_2805,N_2283);
and UO_407 (O_407,N_2356,N_2418);
or UO_408 (O_408,N_2397,N_2681);
nand UO_409 (O_409,N_2847,N_2268);
nand UO_410 (O_410,N_2869,N_2761);
nor UO_411 (O_411,N_2328,N_2505);
nand UO_412 (O_412,N_2921,N_2995);
nor UO_413 (O_413,N_2529,N_2997);
or UO_414 (O_414,N_2435,N_2385);
and UO_415 (O_415,N_2361,N_2617);
or UO_416 (O_416,N_2435,N_2629);
or UO_417 (O_417,N_2270,N_2805);
nand UO_418 (O_418,N_2899,N_2483);
and UO_419 (O_419,N_2624,N_2346);
nand UO_420 (O_420,N_2851,N_2523);
xnor UO_421 (O_421,N_2746,N_2453);
and UO_422 (O_422,N_2259,N_2979);
or UO_423 (O_423,N_2423,N_2934);
and UO_424 (O_424,N_2275,N_2795);
nand UO_425 (O_425,N_2812,N_2672);
nor UO_426 (O_426,N_2753,N_2446);
nand UO_427 (O_427,N_2544,N_2778);
and UO_428 (O_428,N_2263,N_2620);
or UO_429 (O_429,N_2264,N_2704);
nand UO_430 (O_430,N_2906,N_2638);
nand UO_431 (O_431,N_2895,N_2721);
and UO_432 (O_432,N_2500,N_2875);
or UO_433 (O_433,N_2388,N_2289);
nor UO_434 (O_434,N_2383,N_2343);
xnor UO_435 (O_435,N_2857,N_2562);
nor UO_436 (O_436,N_2833,N_2523);
nor UO_437 (O_437,N_2548,N_2849);
or UO_438 (O_438,N_2647,N_2940);
xor UO_439 (O_439,N_2328,N_2801);
nand UO_440 (O_440,N_2739,N_2301);
or UO_441 (O_441,N_2964,N_2608);
nor UO_442 (O_442,N_2721,N_2553);
and UO_443 (O_443,N_2613,N_2503);
nand UO_444 (O_444,N_2667,N_2778);
or UO_445 (O_445,N_2756,N_2417);
nand UO_446 (O_446,N_2768,N_2324);
nor UO_447 (O_447,N_2743,N_2787);
nor UO_448 (O_448,N_2765,N_2826);
nand UO_449 (O_449,N_2726,N_2838);
nand UO_450 (O_450,N_2618,N_2636);
or UO_451 (O_451,N_2731,N_2413);
nand UO_452 (O_452,N_2412,N_2631);
or UO_453 (O_453,N_2511,N_2550);
nor UO_454 (O_454,N_2748,N_2731);
and UO_455 (O_455,N_2575,N_2423);
nand UO_456 (O_456,N_2375,N_2709);
and UO_457 (O_457,N_2609,N_2991);
nand UO_458 (O_458,N_2785,N_2718);
nor UO_459 (O_459,N_2583,N_2651);
nand UO_460 (O_460,N_2946,N_2283);
nand UO_461 (O_461,N_2285,N_2573);
nor UO_462 (O_462,N_2974,N_2826);
or UO_463 (O_463,N_2759,N_2630);
nand UO_464 (O_464,N_2584,N_2911);
nor UO_465 (O_465,N_2514,N_2756);
or UO_466 (O_466,N_2811,N_2764);
and UO_467 (O_467,N_2797,N_2748);
and UO_468 (O_468,N_2878,N_2948);
and UO_469 (O_469,N_2725,N_2805);
and UO_470 (O_470,N_2837,N_2342);
or UO_471 (O_471,N_2597,N_2250);
and UO_472 (O_472,N_2499,N_2269);
and UO_473 (O_473,N_2603,N_2320);
or UO_474 (O_474,N_2628,N_2987);
or UO_475 (O_475,N_2542,N_2882);
nor UO_476 (O_476,N_2512,N_2610);
and UO_477 (O_477,N_2878,N_2915);
or UO_478 (O_478,N_2542,N_2736);
and UO_479 (O_479,N_2264,N_2885);
or UO_480 (O_480,N_2497,N_2699);
or UO_481 (O_481,N_2732,N_2534);
nand UO_482 (O_482,N_2600,N_2286);
nand UO_483 (O_483,N_2953,N_2545);
nand UO_484 (O_484,N_2601,N_2833);
or UO_485 (O_485,N_2647,N_2335);
nor UO_486 (O_486,N_2615,N_2603);
xor UO_487 (O_487,N_2803,N_2425);
or UO_488 (O_488,N_2407,N_2514);
and UO_489 (O_489,N_2809,N_2573);
or UO_490 (O_490,N_2961,N_2782);
or UO_491 (O_491,N_2404,N_2327);
nor UO_492 (O_492,N_2323,N_2776);
or UO_493 (O_493,N_2991,N_2500);
nor UO_494 (O_494,N_2876,N_2837);
nand UO_495 (O_495,N_2956,N_2355);
and UO_496 (O_496,N_2588,N_2386);
or UO_497 (O_497,N_2889,N_2552);
and UO_498 (O_498,N_2621,N_2324);
or UO_499 (O_499,N_2323,N_2693);
endmodule