module basic_2500_25000_3000_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1459,In_608);
and U1 (N_1,In_1791,In_1476);
nor U2 (N_2,In_530,In_2103);
or U3 (N_3,In_1626,In_2138);
or U4 (N_4,In_221,In_489);
or U5 (N_5,In_1087,In_2302);
nand U6 (N_6,In_481,In_1207);
nor U7 (N_7,In_809,In_2193);
xor U8 (N_8,In_1224,In_1462);
xor U9 (N_9,In_1072,In_2203);
and U10 (N_10,In_1311,In_1983);
or U11 (N_11,In_1096,In_898);
or U12 (N_12,In_1604,In_2378);
xor U13 (N_13,In_1810,In_714);
or U14 (N_14,In_1873,In_1113);
nand U15 (N_15,In_86,In_230);
and U16 (N_16,In_239,In_2145);
nor U17 (N_17,In_1473,In_93);
or U18 (N_18,In_2278,In_1013);
nand U19 (N_19,In_829,In_296);
xor U20 (N_20,In_1858,In_1898);
and U21 (N_21,In_2197,In_2347);
xnor U22 (N_22,In_499,In_2326);
nor U23 (N_23,In_1758,In_1310);
or U24 (N_24,In_1723,In_1931);
and U25 (N_25,In_1914,In_633);
xnor U26 (N_26,In_219,In_2035);
and U27 (N_27,In_207,In_1895);
or U28 (N_28,In_1583,In_2421);
or U29 (N_29,In_2364,In_1512);
or U30 (N_30,In_1998,In_1492);
nor U31 (N_31,In_1920,In_1141);
and U32 (N_32,In_1707,In_312);
nor U33 (N_33,In_1692,In_779);
nor U34 (N_34,In_2221,In_1897);
and U35 (N_35,In_1672,In_1102);
xor U36 (N_36,In_2062,In_1718);
and U37 (N_37,In_1896,In_145);
nand U38 (N_38,In_233,In_399);
xor U39 (N_39,In_2122,In_1260);
nor U40 (N_40,In_1043,In_163);
xor U41 (N_41,In_1855,In_990);
or U42 (N_42,In_1901,In_1019);
nor U43 (N_43,In_242,In_1635);
or U44 (N_44,In_1467,In_492);
or U45 (N_45,In_1805,In_2011);
or U46 (N_46,In_1244,In_869);
nand U47 (N_47,In_1384,In_2482);
nor U48 (N_48,In_2371,In_862);
or U49 (N_49,In_18,In_453);
or U50 (N_50,In_2411,In_20);
or U51 (N_51,In_2432,In_1843);
nor U52 (N_52,In_1757,In_143);
or U53 (N_53,In_903,In_335);
nor U54 (N_54,In_1793,In_1768);
nand U55 (N_55,In_1077,In_1232);
xor U56 (N_56,In_1204,In_2446);
xnor U57 (N_57,In_1331,In_635);
nor U58 (N_58,In_1688,In_120);
nand U59 (N_59,In_2340,In_2318);
nand U60 (N_60,In_1504,In_2042);
or U61 (N_61,In_877,In_1383);
or U62 (N_62,In_403,In_2236);
and U63 (N_63,In_988,In_2419);
nor U64 (N_64,In_117,In_1676);
nand U65 (N_65,In_2324,In_951);
or U66 (N_66,In_1779,In_2405);
nand U67 (N_67,In_2451,In_1618);
nor U68 (N_68,In_1689,In_2273);
or U69 (N_69,In_309,In_1407);
nor U70 (N_70,In_1036,In_1411);
nand U71 (N_71,In_54,In_109);
and U72 (N_72,In_1554,In_1521);
nor U73 (N_73,In_2356,In_1927);
or U74 (N_74,In_2161,In_11);
nand U75 (N_75,In_1817,In_613);
nor U76 (N_76,In_1069,In_618);
or U77 (N_77,In_1208,In_2438);
nand U78 (N_78,In_2399,In_843);
nand U79 (N_79,In_1929,In_2168);
xor U80 (N_80,In_1155,In_2157);
and U81 (N_81,In_213,In_616);
and U82 (N_82,In_2296,In_1250);
nor U83 (N_83,In_1441,In_388);
nand U84 (N_84,In_730,In_1164);
and U85 (N_85,In_2165,In_1661);
nor U86 (N_86,In_1387,In_1888);
nand U87 (N_87,In_2447,In_470);
and U88 (N_88,In_577,In_1321);
and U89 (N_89,In_1477,In_900);
nand U90 (N_90,In_151,In_2458);
nand U91 (N_91,In_1559,In_421);
and U92 (N_92,In_115,In_1416);
and U93 (N_93,In_1478,In_544);
nand U94 (N_94,In_1022,In_505);
nand U95 (N_95,In_1788,In_1389);
nor U96 (N_96,In_1205,In_2316);
nand U97 (N_97,In_1760,In_643);
nand U98 (N_98,In_1668,In_2417);
and U99 (N_99,In_2362,In_136);
nor U100 (N_100,In_1913,In_2250);
and U101 (N_101,In_1842,In_1453);
or U102 (N_102,In_1307,In_1582);
and U103 (N_103,In_1191,In_264);
nor U104 (N_104,In_1484,In_169);
xnor U105 (N_105,In_302,In_2144);
or U106 (N_106,In_1755,In_756);
xnor U107 (N_107,In_992,In_1217);
or U108 (N_108,In_1014,In_1370);
xnor U109 (N_109,In_2409,In_45);
nor U110 (N_110,In_1654,In_1883);
xor U111 (N_111,In_1868,In_1497);
and U112 (N_112,In_2338,In_1825);
xnor U113 (N_113,In_275,In_2243);
or U114 (N_114,In_1976,In_1192);
nor U115 (N_115,In_2276,In_1295);
xnor U116 (N_116,In_611,In_217);
nand U117 (N_117,In_153,In_2357);
nor U118 (N_118,In_1093,In_92);
or U119 (N_119,In_974,In_197);
or U120 (N_120,In_95,In_2418);
xnor U121 (N_121,In_2480,In_1899);
xnor U122 (N_122,In_2190,In_251);
nand U123 (N_123,In_673,In_2379);
nor U124 (N_124,In_1270,In_2189);
nor U125 (N_125,In_979,In_1274);
xnor U126 (N_126,In_462,In_1405);
nand U127 (N_127,In_2292,In_171);
nor U128 (N_128,In_2381,In_376);
nand U129 (N_129,In_2436,In_989);
nand U130 (N_130,In_1592,In_268);
or U131 (N_131,In_812,In_2075);
or U132 (N_132,In_1452,In_939);
nor U133 (N_133,In_280,In_1126);
xor U134 (N_134,In_1774,In_1990);
nand U135 (N_135,In_1082,In_460);
xor U136 (N_136,In_2218,In_1738);
and U137 (N_137,In_849,In_389);
and U138 (N_138,In_1349,In_2228);
nor U139 (N_139,In_2283,In_1677);
and U140 (N_140,In_2044,In_2286);
or U141 (N_141,In_2487,In_2472);
and U142 (N_142,In_2014,In_634);
or U143 (N_143,In_728,In_435);
and U144 (N_144,In_114,In_1359);
and U145 (N_145,In_517,In_46);
xnor U146 (N_146,In_1992,In_579);
xnor U147 (N_147,In_1061,In_1534);
or U148 (N_148,In_667,In_290);
nand U149 (N_149,In_347,In_1719);
and U150 (N_150,In_814,In_2137);
nor U151 (N_151,In_407,In_484);
nor U152 (N_152,In_1801,In_285);
and U153 (N_153,In_1440,In_628);
and U154 (N_154,In_64,In_234);
nand U155 (N_155,In_953,In_1458);
nand U156 (N_156,In_1622,In_1764);
nand U157 (N_157,In_589,In_1769);
nor U158 (N_158,In_2212,In_455);
or U159 (N_159,In_2425,In_998);
or U160 (N_160,In_1797,In_610);
nor U161 (N_161,In_1656,In_2476);
or U162 (N_162,In_1045,In_412);
nor U163 (N_163,In_1814,In_2106);
nor U164 (N_164,In_1860,In_1978);
nand U165 (N_165,In_59,In_1246);
xor U166 (N_166,In_1300,In_68);
or U167 (N_167,In_2028,In_2146);
nor U168 (N_168,In_195,In_2252);
xor U169 (N_169,In_2444,In_886);
and U170 (N_170,In_2257,In_336);
and U171 (N_171,In_1881,In_63);
xor U172 (N_172,In_1848,In_612);
nor U173 (N_173,In_1366,In_2462);
nand U174 (N_174,In_1979,In_2009);
and U175 (N_175,In_1112,In_522);
and U176 (N_176,In_2491,In_1563);
and U177 (N_177,In_1678,In_2439);
nand U178 (N_178,In_2047,In_1051);
and U179 (N_179,In_334,In_2017);
xnor U180 (N_180,In_644,In_1123);
or U181 (N_181,In_539,In_1569);
nand U182 (N_182,In_969,In_1067);
nor U183 (N_183,In_1722,In_413);
and U184 (N_184,In_214,In_260);
and U185 (N_185,In_905,In_1221);
nand U186 (N_186,In_1047,In_983);
nor U187 (N_187,In_1390,In_734);
xnor U188 (N_188,In_1413,In_1294);
nand U189 (N_189,In_825,In_894);
nor U190 (N_190,In_270,In_1227);
nor U191 (N_191,In_493,In_2427);
nand U192 (N_192,In_1536,In_999);
nand U193 (N_193,In_382,In_946);
nand U194 (N_194,In_1892,In_231);
nor U195 (N_195,In_1524,In_2021);
nand U196 (N_196,In_1851,In_1510);
nor U197 (N_197,In_1776,In_1857);
nor U198 (N_198,In_1275,In_1790);
and U199 (N_199,In_1555,In_1258);
nor U200 (N_200,In_875,In_1601);
xor U201 (N_201,In_368,In_273);
and U202 (N_202,In_2064,In_1172);
or U203 (N_203,In_101,In_1968);
nand U204 (N_204,In_1507,In_556);
and U205 (N_205,In_2385,In_911);
nand U206 (N_206,In_344,In_71);
xnor U207 (N_207,In_1131,In_2130);
xnor U208 (N_208,In_586,In_626);
nor U209 (N_209,In_1392,In_1753);
nand U210 (N_210,In_427,In_181);
nor U211 (N_211,In_768,In_1616);
and U212 (N_212,In_1171,In_1924);
and U213 (N_213,In_2060,In_1345);
and U214 (N_214,In_430,In_198);
and U215 (N_215,In_524,In_1007);
and U216 (N_216,In_1229,In_787);
nor U217 (N_217,In_56,In_1731);
nor U218 (N_218,In_1354,In_594);
xor U219 (N_219,In_1403,In_2051);
xnor U220 (N_220,In_777,In_2262);
nor U221 (N_221,In_2019,In_947);
or U222 (N_222,In_1283,In_1659);
xor U223 (N_223,In_1828,In_1176);
nor U224 (N_224,In_1190,In_884);
nand U225 (N_225,In_1298,In_237);
xor U226 (N_226,In_1775,In_1461);
or U227 (N_227,In_1949,In_1648);
or U228 (N_228,In_2117,In_994);
or U229 (N_229,In_627,In_856);
xnor U230 (N_230,In_1284,In_2241);
nand U231 (N_231,In_917,In_2374);
nand U232 (N_232,In_326,In_861);
xor U233 (N_233,In_2498,In_23);
nor U234 (N_234,In_1612,In_1840);
or U235 (N_235,In_2333,In_915);
or U236 (N_236,In_362,In_2183);
nor U237 (N_237,In_1375,In_2158);
nor U238 (N_238,In_1887,In_1641);
and U239 (N_239,In_1362,In_1412);
nor U240 (N_240,In_1038,In_1450);
nand U241 (N_241,In_1026,In_1308);
xor U242 (N_242,In_374,In_919);
or U243 (N_243,In_1079,In_229);
and U244 (N_244,In_2054,In_2494);
nor U245 (N_245,In_1188,In_416);
nand U246 (N_246,In_2251,In_2429);
xnor U247 (N_247,In_2109,In_99);
or U248 (N_248,In_1186,In_395);
and U249 (N_249,In_672,In_2084);
xor U250 (N_250,In_822,In_75);
xor U251 (N_251,In_28,In_749);
nand U252 (N_252,In_1291,In_1097);
or U253 (N_253,In_941,In_803);
xor U254 (N_254,In_1647,In_2320);
and U255 (N_255,In_1379,In_107);
xor U256 (N_256,In_257,In_1008);
nand U257 (N_257,In_425,In_929);
or U258 (N_258,In_1076,In_1593);
nand U259 (N_259,In_699,In_1455);
or U260 (N_260,In_1735,In_1746);
nand U261 (N_261,In_646,In_811);
nor U262 (N_262,In_641,In_318);
nand U263 (N_263,In_355,In_933);
and U264 (N_264,In_906,In_1620);
and U265 (N_265,In_10,In_2369);
nand U266 (N_266,In_161,In_1212);
xor U267 (N_267,In_2431,In_1649);
xnor U268 (N_268,In_702,In_450);
nor U269 (N_269,In_1596,In_2152);
and U270 (N_270,In_1865,In_1074);
nor U271 (N_271,In_661,In_110);
or U272 (N_272,In_924,In_441);
or U273 (N_273,In_78,In_1815);
nand U274 (N_274,In_935,In_27);
nor U275 (N_275,In_1919,In_743);
and U276 (N_276,In_418,In_540);
and U277 (N_277,In_658,In_1962);
or U278 (N_278,In_736,In_49);
nand U279 (N_279,In_1875,In_1189);
nor U280 (N_280,In_357,In_420);
nor U281 (N_281,In_1617,In_1488);
xnor U282 (N_282,In_194,In_546);
nor U283 (N_283,In_1154,In_2070);
and U284 (N_284,In_1326,In_629);
and U285 (N_285,In_1419,In_2355);
or U286 (N_286,In_2155,In_1947);
xnor U287 (N_287,In_1558,In_1121);
nand U288 (N_288,In_1959,In_1471);
xnor U289 (N_289,In_2058,In_695);
or U290 (N_290,In_2287,In_2202);
nand U291 (N_291,In_2255,In_1342);
and U292 (N_292,In_1629,In_536);
xnor U293 (N_293,In_1553,In_2323);
xnor U294 (N_294,In_1704,In_483);
nor U295 (N_295,In_1290,In_1634);
nand U296 (N_296,In_1351,In_864);
or U297 (N_297,In_909,In_1705);
nand U298 (N_298,In_1631,In_2353);
or U299 (N_299,In_34,In_1786);
and U300 (N_300,In_896,In_1133);
nor U301 (N_301,In_750,In_445);
nand U302 (N_302,In_2050,In_2459);
and U303 (N_303,In_246,In_1950);
and U304 (N_304,In_837,In_866);
nand U305 (N_305,In_1422,In_914);
and U306 (N_306,In_1847,In_600);
and U307 (N_307,In_1348,In_1528);
nand U308 (N_308,In_188,In_904);
or U309 (N_309,In_428,In_1060);
nand U310 (N_310,In_391,In_1444);
nand U311 (N_311,In_254,In_2211);
nor U312 (N_312,In_1989,In_1970);
nor U313 (N_313,In_4,In_72);
nand U314 (N_314,In_851,In_839);
nand U315 (N_315,In_1385,In_1119);
and U316 (N_316,In_2141,In_2092);
and U317 (N_317,In_2235,In_2031);
xor U318 (N_318,In_859,In_2331);
and U319 (N_319,In_2184,In_1454);
nand U320 (N_320,In_2238,In_716);
xor U321 (N_321,In_76,In_1235);
or U322 (N_322,In_465,In_2032);
nor U323 (N_323,In_2408,In_2082);
or U324 (N_324,In_2121,In_1627);
xnor U325 (N_325,In_1261,In_575);
and U326 (N_326,In_183,In_352);
xnor U327 (N_327,In_1430,In_1834);
and U328 (N_328,In_620,In_1516);
or U329 (N_329,In_2359,In_1566);
and U330 (N_330,In_104,In_179);
or U331 (N_331,In_967,In_1339);
xor U332 (N_332,In_1703,In_984);
or U333 (N_333,In_1690,In_590);
xor U334 (N_334,In_1490,In_1174);
or U335 (N_335,In_343,In_1799);
and U336 (N_336,In_593,In_2346);
xnor U337 (N_337,In_43,In_2467);
and U338 (N_338,In_1509,In_2253);
and U339 (N_339,In_823,In_1195);
xor U340 (N_340,In_1715,In_799);
xor U341 (N_341,In_1772,In_396);
and U342 (N_342,In_2013,In_69);
xnor U343 (N_343,In_2052,In_2);
or U344 (N_344,In_645,In_199);
nor U345 (N_345,In_860,In_1431);
xor U346 (N_346,In_2401,In_731);
and U347 (N_347,In_791,In_449);
and U348 (N_348,In_571,In_1286);
or U349 (N_349,In_187,In_2167);
or U350 (N_350,In_1198,In_1474);
or U351 (N_351,In_2328,In_350);
or U352 (N_352,In_842,In_631);
or U353 (N_353,In_781,In_835);
or U354 (N_354,In_541,In_621);
nand U355 (N_355,In_1015,In_1139);
nand U356 (N_356,In_226,In_2475);
and U357 (N_357,In_1748,In_2100);
or U358 (N_358,In_558,In_1251);
xor U359 (N_359,In_1663,In_82);
and U360 (N_360,In_1729,In_278);
xnor U361 (N_361,In_1151,In_180);
xnor U362 (N_362,In_1505,In_2342);
or U363 (N_363,In_2478,In_1495);
xnor U364 (N_364,In_1382,In_1150);
xor U365 (N_365,In_139,In_261);
xnor U366 (N_366,In_2305,In_380);
nand U367 (N_367,In_1075,In_1900);
and U368 (N_368,In_2023,In_1680);
nand U369 (N_369,In_985,In_2209);
nor U370 (N_370,In_360,In_328);
and U371 (N_371,In_310,In_1143);
nand U372 (N_372,In_1269,In_2002);
xor U373 (N_373,In_1686,In_689);
or U374 (N_374,In_783,In_1942);
or U375 (N_375,In_2249,In_1822);
and U376 (N_376,In_675,In_2005);
nor U377 (N_377,In_2123,In_1049);
nor U378 (N_378,In_166,In_1885);
and U379 (N_379,In_542,In_1570);
or U380 (N_380,In_751,In_1357);
nor U381 (N_381,In_1967,In_1698);
xor U382 (N_382,In_390,In_1052);
and U383 (N_383,In_1262,In_1891);
or U384 (N_384,In_1009,In_314);
or U385 (N_385,In_1381,In_474);
or U386 (N_386,In_2410,In_668);
and U387 (N_387,In_912,In_307);
nand U388 (N_388,In_501,In_2341);
or U389 (N_389,In_1856,In_1089);
and U390 (N_390,In_2350,In_1000);
or U391 (N_391,In_1011,In_2481);
xnor U392 (N_392,In_323,In_1081);
xor U393 (N_393,In_1029,In_426);
xnor U394 (N_394,In_1564,In_1702);
or U395 (N_395,In_209,In_1048);
nor U396 (N_396,In_2149,In_2282);
xnor U397 (N_397,In_2456,In_480);
and U398 (N_398,In_458,In_1526);
or U399 (N_399,In_1464,In_252);
nor U400 (N_400,In_1273,In_1882);
or U401 (N_401,In_778,In_1845);
or U402 (N_402,In_175,In_1918);
and U403 (N_403,In_2003,In_434);
or U404 (N_404,In_1030,In_2453);
nand U405 (N_405,In_2396,In_792);
or U406 (N_406,In_372,In_2300);
and U407 (N_407,In_341,In_840);
xnor U408 (N_408,In_2339,In_555);
and U409 (N_409,In_1584,In_1378);
or U410 (N_410,In_1827,In_545);
and U411 (N_411,In_2440,In_981);
and U412 (N_412,In_141,In_255);
xnor U413 (N_413,In_2483,In_1182);
or U414 (N_414,In_1577,In_2389);
xnor U415 (N_415,In_732,In_519);
or U416 (N_416,In_476,In_1912);
or U417 (N_417,In_680,In_17);
xor U418 (N_418,In_1608,In_282);
xnor U419 (N_419,In_1499,In_1181);
nor U420 (N_420,In_882,In_1988);
xnor U421 (N_421,In_1289,In_1325);
nand U422 (N_422,In_1070,In_1073);
and U423 (N_423,In_411,In_306);
xor U424 (N_424,In_1439,In_332);
and U425 (N_425,In_960,In_1006);
and U426 (N_426,In_1522,In_2204);
xor U427 (N_427,In_885,In_1021);
and U428 (N_428,In_665,In_982);
and U429 (N_429,In_406,In_2315);
or U430 (N_430,In_1266,In_614);
or U431 (N_431,In_1624,In_1646);
or U432 (N_432,In_2071,In_692);
and U433 (N_433,In_1819,In_1614);
nand U434 (N_434,In_1402,In_29);
and U435 (N_435,In_574,In_1055);
and U436 (N_436,In_1434,In_683);
nand U437 (N_437,In_523,In_1278);
nand U438 (N_438,In_2312,In_2397);
and U439 (N_439,In_1201,In_2216);
xor U440 (N_440,In_1889,In_1813);
nor U441 (N_441,In_2336,In_97);
or U442 (N_442,In_440,In_433);
and U443 (N_443,In_482,In_720);
nor U444 (N_444,In_2102,In_1849);
and U445 (N_445,In_2056,In_1046);
nor U446 (N_446,In_681,In_124);
xor U447 (N_447,In_1682,In_1546);
xnor U448 (N_448,In_1020,In_955);
xor U449 (N_449,In_794,In_2244);
xor U450 (N_450,In_22,In_1724);
nand U451 (N_451,In_35,In_1018);
and U452 (N_452,In_375,In_1727);
nand U453 (N_453,In_1025,In_1866);
nand U454 (N_454,In_2053,In_70);
and U455 (N_455,In_1800,In_444);
nand U456 (N_456,In_1833,In_1784);
and U457 (N_457,In_1694,In_24);
nand U458 (N_458,In_804,In_503);
or U459 (N_459,In_707,In_2027);
and U460 (N_460,In_518,In_2465);
or U461 (N_461,In_438,In_2259);
nor U462 (N_462,In_2104,In_1309);
nor U463 (N_463,In_1406,In_284);
nor U464 (N_464,In_1196,In_2348);
nand U465 (N_465,In_1780,In_202);
xnor U466 (N_466,In_2010,In_2065);
nand U467 (N_467,In_2126,In_1508);
nor U468 (N_468,In_744,In_930);
nor U469 (N_469,In_494,In_2461);
nor U470 (N_470,In_1223,In_2437);
or U471 (N_471,In_1475,In_977);
nor U472 (N_472,In_201,In_1130);
xor U473 (N_473,In_1589,In_588);
nor U474 (N_474,In_1581,In_1306);
xor U475 (N_475,In_304,In_604);
or U476 (N_476,In_685,In_2469);
xor U477 (N_477,In_773,In_1216);
or U478 (N_478,In_1766,In_561);
and U479 (N_479,In_325,In_549);
and U480 (N_480,In_42,In_2435);
or U481 (N_481,In_1579,In_220);
or U482 (N_482,In_2140,In_1761);
and U483 (N_483,In_782,In_648);
xnor U484 (N_484,In_2069,In_1092);
or U485 (N_485,In_578,In_1368);
xnor U486 (N_486,In_2055,In_1798);
xor U487 (N_487,In_9,In_2365);
xor U488 (N_488,In_2358,In_508);
and U489 (N_489,In_826,In_1482);
xnor U490 (N_490,In_1533,In_329);
xnor U491 (N_491,In_666,In_77);
xnor U492 (N_492,In_2008,In_770);
and U493 (N_493,In_1436,In_2059);
or U494 (N_494,In_709,In_1973);
nand U495 (N_495,In_580,In_509);
nand U496 (N_496,In_2068,In_1869);
nor U497 (N_497,In_932,In_934);
nand U498 (N_498,In_31,In_1206);
or U499 (N_499,In_507,In_2386);
nand U500 (N_500,In_1759,In_487);
nand U501 (N_501,In_1573,In_85);
and U502 (N_502,In_448,In_1829);
or U503 (N_503,In_2463,In_700);
nor U504 (N_504,In_1446,In_287);
xnor U505 (N_505,In_562,In_2006);
or U506 (N_506,In_1256,In_1619);
and U507 (N_507,In_581,In_203);
xor U508 (N_508,In_1085,In_1183);
and U509 (N_509,In_870,In_2034);
or U510 (N_510,In_1108,In_155);
nand U511 (N_511,In_1997,In_1447);
or U512 (N_512,In_1481,In_2087);
nor U513 (N_513,In_1744,In_1320);
and U514 (N_514,In_2373,In_1347);
and U515 (N_515,In_1863,In_1921);
nor U516 (N_516,In_240,In_1315);
xnor U517 (N_517,In_2242,In_1605);
nor U518 (N_518,In_543,In_1388);
xnor U519 (N_519,In_13,In_592);
nand U520 (N_520,In_303,In_660);
and U521 (N_521,In_622,In_122);
nand U522 (N_522,In_937,In_2085);
or U523 (N_523,In_1170,In_60);
nor U524 (N_524,In_664,In_2232);
or U525 (N_525,In_2185,In_300);
and U526 (N_526,In_1145,In_841);
xnor U527 (N_527,In_1099,In_40);
nor U528 (N_528,In_1606,In_291);
xnor U529 (N_529,In_1001,In_2061);
or U530 (N_530,In_1638,In_1494);
nand U531 (N_531,In_1886,In_1936);
xor U532 (N_532,In_688,In_916);
nand U533 (N_533,In_1934,In_1485);
nand U534 (N_534,In_1303,In_824);
and U535 (N_535,In_936,In_81);
nor U536 (N_536,In_748,In_1541);
xor U537 (N_537,In_1428,In_649);
xnor U538 (N_538,In_1358,In_491);
xnor U539 (N_539,In_1118,In_1532);
and U540 (N_540,In_922,In_2131);
xor U541 (N_541,In_2317,In_1337);
nand U542 (N_542,In_65,In_975);
xnor U543 (N_543,In_830,In_553);
xor U544 (N_544,In_653,In_2490);
and U545 (N_545,In_1429,In_477);
xnor U546 (N_546,In_2119,In_2217);
xnor U547 (N_547,In_701,In_1807);
and U548 (N_548,In_185,In_2370);
nand U549 (N_549,In_1252,In_112);
nand U550 (N_550,In_1037,In_383);
and U551 (N_551,In_1518,In_316);
nor U552 (N_552,In_1129,In_962);
xnor U553 (N_553,In_2154,In_512);
and U554 (N_554,In_2135,In_1696);
nor U555 (N_555,In_1946,In_1408);
nand U556 (N_556,In_1529,In_1911);
nor U557 (N_557,In_2423,In_1041);
and U558 (N_558,In_2309,In_637);
and U559 (N_559,In_2147,In_1971);
and U560 (N_560,In_398,In_1418);
nor U561 (N_561,In_1163,In_2443);
and U562 (N_562,In_1115,In_1489);
nand U563 (N_563,In_2192,In_774);
and U564 (N_564,In_146,In_1410);
or U565 (N_565,In_1457,In_1820);
nor U566 (N_566,In_1271,In_1161);
nand U567 (N_567,In_892,In_2097);
or U568 (N_568,In_506,In_339);
nor U569 (N_569,In_520,In_2395);
xnor U570 (N_570,In_1935,In_2208);
or U571 (N_571,In_1916,In_2114);
or U572 (N_572,In_573,In_1657);
and U573 (N_573,In_2254,In_1249);
nor U574 (N_574,In_1053,In_1111);
or U575 (N_575,In_2016,In_1173);
nand U576 (N_576,In_2392,In_1169);
and U577 (N_577,In_1465,In_1233);
nand U578 (N_578,In_1838,In_971);
and U579 (N_579,In_105,In_2363);
nor U580 (N_580,In_1180,In_1336);
and U581 (N_581,In_1225,In_923);
and U582 (N_582,In_2188,In_1670);
nor U583 (N_583,In_2433,In_1024);
or U584 (N_584,In_1660,In_1501);
nor U585 (N_585,In_2288,In_2036);
nand U586 (N_586,In_1101,In_2383);
xor U587 (N_587,In_1480,In_696);
nand U588 (N_588,In_2388,In_315);
nand U589 (N_589,In_2311,In_415);
xnor U590 (N_590,In_1613,In_467);
and U591 (N_591,In_1005,In_1142);
xor U592 (N_592,In_55,In_2270);
xor U593 (N_593,In_910,In_36);
nor U594 (N_594,In_2403,In_342);
nand U595 (N_595,In_1871,In_281);
xor U596 (N_596,In_927,In_2175);
nor U597 (N_597,In_2230,In_1159);
nor U598 (N_598,In_1056,In_2025);
or U599 (N_599,In_1630,In_2073);
and U600 (N_600,In_1110,In_1137);
nand U601 (N_601,In_942,In_2215);
nor U602 (N_602,In_2310,In_1669);
or U603 (N_603,In_2337,In_2063);
xor U604 (N_604,In_345,In_2332);
and U605 (N_605,In_2182,In_2136);
xnor U606 (N_606,In_2489,In_1083);
nor U607 (N_607,In_1364,In_190);
or U608 (N_608,In_91,In_2004);
nor U609 (N_609,In_1928,In_2284);
nor U610 (N_610,In_832,In_414);
or U611 (N_611,In_1215,In_2390);
nor U612 (N_612,In_1932,In_1487);
or U613 (N_613,In_2285,In_807);
nand U614 (N_614,In_2248,In_2445);
nor U615 (N_615,In_1726,In_1796);
xor U616 (N_616,In_1127,In_2290);
or U617 (N_617,In_1222,In_1218);
or U618 (N_618,In_1373,In_2205);
xor U619 (N_619,In_557,In_2039);
nand U620 (N_620,In_2279,In_657);
nor U621 (N_621,In_1255,In_1837);
and U622 (N_622,In_1763,In_855);
nor U623 (N_623,In_1296,In_496);
and U624 (N_624,In_2261,In_378);
or U625 (N_625,In_2180,In_1531);
nor U626 (N_626,In_1878,In_486);
xnor U627 (N_627,In_2349,In_330);
nor U628 (N_628,In_2012,In_806);
and U629 (N_629,In_1503,In_116);
xor U630 (N_630,In_62,In_1071);
xor U631 (N_631,In_1078,In_2086);
nor U632 (N_632,In_1506,In_844);
and U633 (N_633,In_754,In_1693);
xnor U634 (N_634,In_853,In_1340);
or U635 (N_635,In_595,In_498);
and U636 (N_636,In_446,In_1313);
nand U637 (N_637,In_1114,In_289);
nor U638 (N_638,In_1655,In_568);
or U639 (N_639,In_215,In_1821);
or U640 (N_640,In_1639,In_454);
nor U641 (N_641,In_1185,In_1352);
xnor U642 (N_642,In_2468,In_691);
nor U643 (N_643,In_276,In_1542);
or U644 (N_644,In_1044,In_761);
nand U645 (N_645,In_1398,In_1832);
or U646 (N_646,In_1219,In_2046);
or U647 (N_647,In_1652,In_241);
xor U648 (N_648,In_1804,In_108);
and U649 (N_649,In_205,In_2402);
or U650 (N_650,In_2234,In_2413);
nand U651 (N_651,In_2162,In_1977);
xor U652 (N_652,In_2280,In_891);
xor U653 (N_653,In_684,In_513);
xor U654 (N_654,In_1653,In_996);
xor U655 (N_655,In_719,In_607);
or U656 (N_656,In_16,In_619);
nand U657 (N_657,In_2354,In_928);
nand U658 (N_658,In_959,In_2345);
and U659 (N_659,In_1124,In_443);
and U660 (N_660,In_758,In_2343);
xnor U661 (N_661,In_1502,In_2231);
nor U662 (N_662,In_599,In_2210);
and U663 (N_663,In_351,In_1369);
or U664 (N_664,In_1239,In_817);
or U665 (N_665,In_880,In_1586);
nand U666 (N_666,In_1771,In_1443);
xor U667 (N_667,In_674,In_1623);
nor U668 (N_668,In_126,In_1933);
nand U669 (N_669,In_652,In_401);
or U670 (N_670,In_51,In_1841);
xnor U671 (N_671,In_150,In_1720);
nand U672 (N_672,In_678,In_2398);
nor U673 (N_673,In_2414,In_495);
nand U674 (N_674,In_2266,In_80);
or U675 (N_675,In_1965,In_2030);
nor U676 (N_676,In_956,In_165);
nor U677 (N_677,In_478,In_582);
nor U678 (N_678,In_361,In_1116);
nor U679 (N_679,In_845,In_1697);
xnor U680 (N_680,In_887,In_693);
nand U681 (N_681,In_1765,In_379);
or U682 (N_682,In_1609,In_1469);
xnor U683 (N_683,In_147,In_2291);
nand U684 (N_684,In_48,In_2260);
or U685 (N_685,In_819,In_1292);
nand U686 (N_686,In_1567,In_127);
xor U687 (N_687,In_2173,In_1433);
nand U688 (N_688,In_847,In_61);
or U689 (N_689,In_2496,In_410);
and U690 (N_690,In_1211,In_1199);
or U691 (N_691,In_1751,In_1789);
nor U692 (N_692,In_1050,In_1602);
nor U693 (N_693,In_1809,In_1177);
and U694 (N_694,In_1844,In_196);
xor U695 (N_695,In_815,In_1);
nand U696 (N_696,In_663,In_584);
nand U697 (N_697,In_908,In_1874);
and U698 (N_698,In_526,In_1880);
or U699 (N_699,In_1109,In_572);
nor U700 (N_700,In_1297,In_2351);
nand U701 (N_701,In_1941,In_1802);
and U702 (N_702,In_1386,In_1166);
or U703 (N_703,In_1367,In_2313);
or U704 (N_704,In_1621,In_1394);
or U705 (N_705,In_497,In_895);
nor U706 (N_706,In_2029,In_2187);
nor U707 (N_707,In_1344,In_852);
xnor U708 (N_708,In_2464,In_1420);
or U709 (N_709,In_500,In_2297);
or U710 (N_710,In_767,In_2470);
xor U711 (N_711,In_1335,In_2471);
or U712 (N_712,In_152,In_1572);
nor U713 (N_713,In_1923,In_1535);
xnor U714 (N_714,In_827,In_2420);
nor U715 (N_715,In_2387,In_1107);
and U716 (N_716,In_2038,In_128);
xnor U717 (N_717,In_818,In_1323);
nand U718 (N_718,In_1513,In_980);
nand U719 (N_719,In_451,In_550);
and U720 (N_720,In_1777,In_140);
nand U721 (N_721,In_1565,In_686);
nand U722 (N_722,In_795,In_769);
nor U723 (N_723,In_1104,In_1371);
xor U724 (N_724,In_1835,In_1088);
nor U725 (N_725,In_1539,In_2477);
nor U726 (N_726,In_790,In_2382);
nor U727 (N_727,In_26,In_2037);
nor U728 (N_728,In_1794,In_760);
or U729 (N_729,In_247,In_135);
nand U730 (N_730,In_2223,In_1922);
and U731 (N_731,In_1228,In_2077);
or U732 (N_732,In_363,In_2493);
nor U733 (N_733,In_2299,In_1240);
nand U734 (N_734,In_1674,In_370);
and U735 (N_735,In_757,In_565);
xor U736 (N_736,In_1867,In_1035);
and U737 (N_737,In_156,In_2272);
or U738 (N_738,In_2449,In_331);
xor U739 (N_739,In_1175,In_1523);
nand U740 (N_740,In_1514,In_793);
nand U741 (N_741,In_1243,In_776);
xnor U742 (N_742,In_364,In_1580);
nor U743 (N_743,In_679,In_2160);
or U744 (N_744,In_1679,In_1318);
or U745 (N_745,In_1353,In_353);
xnor U746 (N_746,In_1762,In_1823);
nor U747 (N_747,In_1710,In_2171);
nor U748 (N_748,In_888,In_970);
or U749 (N_749,In_1836,In_1544);
or U750 (N_750,In_918,In_1153);
nor U751 (N_751,In_881,In_525);
nand U752 (N_752,In_1187,In_1066);
nor U753 (N_753,In_272,In_2394);
and U754 (N_754,In_1633,In_676);
nand U755 (N_755,In_1034,In_1343);
and U756 (N_756,In_1448,In_258);
nand U757 (N_757,In_1254,In_2268);
and U758 (N_758,In_1591,In_1437);
xor U759 (N_759,In_2099,In_1330);
and U760 (N_760,In_299,In_987);
xnor U761 (N_761,In_1515,In_718);
xnor U762 (N_762,In_763,In_2352);
xnor U763 (N_763,In_1953,In_2081);
nor U764 (N_764,In_2452,In_1346);
xor U765 (N_765,In_1363,In_1894);
or U766 (N_766,In_1377,In_514);
and U767 (N_767,In_528,In_961);
and U768 (N_768,In_447,In_1039);
xnor U769 (N_769,In_1545,In_236);
and U770 (N_770,In_392,In_1328);
xor U771 (N_771,In_642,In_468);
or U772 (N_772,In_397,In_436);
and U773 (N_773,In_560,In_1905);
nand U774 (N_774,In_327,In_473);
and U775 (N_775,In_1496,In_2450);
and U776 (N_776,In_2442,In_206);
nor U777 (N_777,In_338,In_1332);
nor U778 (N_778,In_1716,In_2415);
or U779 (N_779,In_1236,In_459);
nand U780 (N_780,In_1826,In_204);
or U781 (N_781,In_172,In_1562);
and U782 (N_782,In_245,In_1691);
and U783 (N_783,In_38,In_1095);
xnor U784 (N_784,In_2306,In_2486);
nor U785 (N_785,In_872,In_597);
or U786 (N_786,In_957,In_986);
and U787 (N_787,In_563,In_765);
or U788 (N_788,In_1695,In_2176);
xor U789 (N_789,In_948,In_2441);
and U790 (N_790,In_533,In_2281);
and U791 (N_791,In_1750,In_2169);
xnor U792 (N_792,In_88,In_243);
xor U793 (N_793,In_132,In_670);
nor U794 (N_794,In_1852,In_973);
nand U795 (N_795,In_1687,In_464);
or U796 (N_796,In_2422,In_2194);
or U797 (N_797,In_587,In_997);
and U798 (N_798,In_305,In_1662);
nor U799 (N_799,In_1355,In_591);
or U800 (N_800,In_2001,In_2247);
nor U801 (N_801,In_1194,In_2072);
nand U802 (N_802,In_944,In_271);
nand U803 (N_803,In_2199,In_369);
xor U804 (N_804,In_893,In_178);
nand U805 (N_805,In_2033,In_1728);
xnor U806 (N_806,In_698,In_250);
and U807 (N_807,In_266,In_784);
or U808 (N_808,In_2107,In_954);
nor U809 (N_809,In_377,In_2303);
xnor U810 (N_810,In_253,In_671);
and U811 (N_811,In_2024,In_1925);
nand U812 (N_812,In_2319,In_349);
nand U813 (N_813,In_697,In_2304);
nor U814 (N_814,In_53,In_2293);
or U815 (N_815,In_2164,In_2133);
and U816 (N_816,In_1879,In_2366);
and U817 (N_817,In_79,In_1981);
nand U818 (N_818,In_1908,In_943);
or U819 (N_819,In_1831,In_2116);
xor U820 (N_820,In_265,In_1948);
or U821 (N_821,In_1721,In_1966);
and U822 (N_822,In_724,In_2224);
nand U823 (N_823,In_2294,In_348);
xnor U824 (N_824,In_96,In_1811);
nand U825 (N_825,In_1016,In_2258);
or U826 (N_826,In_2049,In_1012);
nor U827 (N_827,In_1128,In_2226);
xor U828 (N_828,In_2473,In_1242);
and U829 (N_829,In_2020,In_2112);
nor U830 (N_830,In_262,In_1517);
nand U831 (N_831,In_192,In_1425);
xor U832 (N_832,In_1893,In_1237);
or U833 (N_833,In_387,In_836);
and U834 (N_834,In_1611,In_6);
or U835 (N_835,In_1057,In_1319);
nor U836 (N_836,In_1754,In_2094);
xor U837 (N_837,In_2295,In_712);
nand U838 (N_838,In_2150,In_423);
and U839 (N_839,In_1417,In_1210);
nand U840 (N_840,In_687,In_256);
nor U841 (N_841,In_479,In_958);
xnor U842 (N_842,In_1146,In_2091);
xnor U843 (N_843,In_1238,In_39);
or U844 (N_844,In_3,In_1954);
nor U845 (N_845,In_301,In_1598);
and U846 (N_846,In_1312,In_1850);
xnor U847 (N_847,In_940,In_1282);
or U848 (N_848,In_159,In_1603);
nor U849 (N_849,In_1449,In_1288);
and U850 (N_850,In_2045,In_708);
xnor U851 (N_851,In_1700,In_1717);
or U852 (N_852,In_529,In_424);
nand U853 (N_853,In_677,In_1664);
xor U854 (N_854,In_288,In_1125);
nand U855 (N_855,In_547,In_949);
nor U856 (N_856,In_212,In_1299);
nand U857 (N_857,In_1374,In_726);
nand U858 (N_858,In_755,In_129);
or U859 (N_859,In_2089,In_883);
or U860 (N_860,In_1147,In_1930);
nand U861 (N_861,In_871,In_402);
nor U862 (N_862,In_1595,In_715);
nand U863 (N_863,In_1264,In_2172);
or U864 (N_864,In_2108,In_419);
nand U865 (N_865,In_224,In_1745);
and U866 (N_866,In_1540,In_1165);
nor U867 (N_867,In_890,In_1160);
nor U868 (N_868,In_2080,In_1736);
nand U869 (N_869,In_12,In_1571);
or U870 (N_870,In_2074,In_2151);
nor U871 (N_871,In_2344,In_2163);
nand U872 (N_872,In_615,In_800);
nor U873 (N_873,In_1329,In_184);
xnor U874 (N_874,In_1122,In_1903);
nand U875 (N_875,In_1600,In_2191);
nor U876 (N_876,In_1767,In_1951);
xnor U877 (N_877,In_991,In_1643);
and U878 (N_878,In_472,In_125);
nand U879 (N_879,In_938,In_488);
or U880 (N_880,In_995,In_191);
xnor U881 (N_881,In_952,In_218);
or U882 (N_882,In_654,In_638);
and U883 (N_883,In_1132,In_1247);
nor U884 (N_884,In_1756,In_1773);
nand U885 (N_885,In_52,In_138);
and U886 (N_886,In_1675,In_1945);
and U887 (N_887,In_2040,In_405);
and U888 (N_888,In_532,In_2178);
xor U889 (N_889,In_789,In_925);
xnor U890 (N_890,In_422,In_1301);
or U891 (N_891,In_805,In_2098);
nor U892 (N_892,In_1451,In_810);
or U893 (N_893,In_311,In_1213);
and U894 (N_894,In_2129,In_1574);
nor U895 (N_895,In_1456,In_2043);
nor U896 (N_896,In_907,In_650);
nand U897 (N_897,In_798,In_2289);
nand U898 (N_898,In_1002,In_1556);
nand U899 (N_899,In_286,In_534);
xor U900 (N_900,In_429,In_1588);
nand U901 (N_901,In_2384,In_238);
nor U902 (N_902,In_1961,In_274);
and U903 (N_903,In_15,In_2067);
xor U904 (N_904,In_1839,In_137);
or U905 (N_905,In_704,In_1969);
or U906 (N_906,In_1642,In_682);
and U907 (N_907,In_865,In_879);
or U908 (N_908,In_764,In_1525);
or U909 (N_909,In_740,In_1902);
and U910 (N_910,In_1956,In_2412);
nor U911 (N_911,In_2301,In_1877);
nor U912 (N_912,In_964,In_1267);
and U913 (N_913,In_1876,In_1519);
and U914 (N_914,In_2095,In_1575);
nand U915 (N_915,In_1594,In_457);
nor U916 (N_916,In_1859,In_554);
nand U917 (N_917,In_130,In_1004);
and U918 (N_918,In_1714,In_738);
nand U919 (N_919,In_1483,In_431);
nor U920 (N_920,In_1547,In_102);
nor U921 (N_921,In_729,In_2174);
nor U922 (N_922,In_2220,In_2206);
xor U923 (N_923,In_1421,In_44);
or U924 (N_924,In_2156,In_2041);
or U925 (N_925,In_913,In_576);
nor U926 (N_926,In_1749,In_340);
nor U927 (N_927,In_385,In_2222);
or U928 (N_928,In_1200,In_1442);
or U929 (N_929,In_439,In_2391);
nor U930 (N_930,In_2404,In_537);
or U931 (N_931,In_2265,In_227);
nor U932 (N_932,In_2377,In_308);
nand U933 (N_933,In_47,In_2275);
or U934 (N_934,In_228,In_1438);
xnor U935 (N_935,In_2110,In_1156);
or U936 (N_936,In_2321,In_1220);
xnor U937 (N_937,In_490,In_1792);
and U938 (N_938,In_235,In_394);
or U939 (N_939,In_511,In_123);
xnor U940 (N_940,In_1561,In_1787);
nand U941 (N_941,In_2088,In_617);
or U942 (N_942,In_1610,In_950);
nand U943 (N_943,In_2132,In_1742);
nor U944 (N_944,In_244,In_1673);
nor U945 (N_945,In_1033,In_1202);
xor U946 (N_946,In_2368,In_1415);
or U947 (N_947,In_1987,In_1733);
or U948 (N_948,In_504,In_1560);
nand U949 (N_949,In_33,In_1952);
xor U950 (N_950,In_1996,In_2330);
xor U951 (N_951,In_1498,In_2213);
and U952 (N_952,In_149,In_838);
and U953 (N_953,In_1100,In_850);
and U954 (N_954,In_1599,In_1080);
nor U955 (N_955,In_2460,In_1285);
or U956 (N_956,In_725,In_746);
and U957 (N_957,In_775,In_1785);
or U958 (N_958,In_1027,In_267);
xnor U959 (N_959,In_747,In_632);
and U960 (N_960,In_1511,In_721);
nor U961 (N_961,In_1117,In_651);
nand U962 (N_962,In_828,In_2214);
xor U963 (N_963,In_874,In_131);
nor U964 (N_964,In_1491,In_1683);
nor U965 (N_965,In_222,In_8);
nor U966 (N_966,In_1460,In_1576);
xnor U967 (N_967,In_2327,In_762);
nor U968 (N_968,In_87,In_1197);
and U969 (N_969,In_1701,In_820);
nand U970 (N_970,In_32,In_98);
nor U971 (N_971,In_2159,In_2196);
nor U972 (N_972,In_596,In_1062);
or U973 (N_973,In_2153,In_2148);
or U974 (N_974,In_739,In_834);
or U975 (N_975,In_89,In_100);
and U976 (N_976,In_2329,In_1972);
or U977 (N_977,In_1910,In_2499);
xor U978 (N_978,In_1955,In_2066);
nand U979 (N_979,In_210,In_1615);
nand U980 (N_980,In_1327,In_2400);
or U981 (N_981,In_1904,In_564);
and U982 (N_982,In_2227,In_160);
xnor U983 (N_983,In_710,In_1665);
nor U984 (N_984,In_694,In_662);
nand U985 (N_985,In_1709,In_1527);
and U986 (N_986,In_1752,In_2376);
and U987 (N_987,In_1550,In_1032);
nor U988 (N_988,In_1994,In_1257);
or U989 (N_989,In_2120,In_103);
xor U990 (N_990,In_1372,In_945);
nand U991 (N_991,In_1708,In_1543);
and U992 (N_992,In_1268,In_384);
or U993 (N_993,In_1783,In_1557);
or U994 (N_994,In_796,In_346);
or U995 (N_995,In_1391,In_1090);
or U996 (N_996,In_2455,In_263);
nand U997 (N_997,In_1468,In_1058);
nor U998 (N_998,In_1023,In_647);
and U999 (N_999,In_1824,In_1003);
and U1000 (N_1000,In_322,In_356);
and U1001 (N_1001,In_797,In_1263);
nand U1002 (N_1002,In_320,In_1265);
or U1003 (N_1003,In_2479,In_786);
or U1004 (N_1004,In_208,In_527);
and U1005 (N_1005,In_292,In_1287);
nand U1006 (N_1006,In_1149,In_1140);
nand U1007 (N_1007,In_1915,In_1684);
and U1008 (N_1008,In_1091,In_2018);
and U1009 (N_1009,In_1741,In_1472);
and U1010 (N_1010,In_2113,In_854);
or U1011 (N_1011,In_1862,In_1548);
xor U1012 (N_1012,In_2125,In_2367);
nand U1013 (N_1013,In_2057,In_1304);
or U1014 (N_1014,In_232,In_1530);
xnor U1015 (N_1015,In_1334,In_659);
nand U1016 (N_1016,In_66,In_1414);
nand U1017 (N_1017,In_294,In_2142);
xnor U1018 (N_1018,In_976,In_1830);
or U1019 (N_1019,In_1549,In_83);
xor U1020 (N_1020,In_780,In_1350);
nand U1021 (N_1021,In_2000,In_1158);
nand U1022 (N_1022,In_189,In_639);
nand U1023 (N_1023,In_690,In_1552);
or U1024 (N_1024,In_1241,In_106);
and U1025 (N_1025,In_1193,In_1203);
or U1026 (N_1026,In_1861,In_25);
xor U1027 (N_1027,In_2118,In_656);
xnor U1028 (N_1028,In_5,In_259);
nor U1029 (N_1029,In_167,In_878);
or U1030 (N_1030,In_531,In_1734);
and U1031 (N_1031,In_2267,In_1178);
xnor U1032 (N_1032,In_873,In_1214);
nor U1033 (N_1033,In_1816,In_1985);
xnor U1034 (N_1034,In_1184,In_722);
or U1035 (N_1035,In_2239,In_902);
nor U1036 (N_1036,In_1393,In_978);
xor U1037 (N_1037,In_1168,In_669);
nand U1038 (N_1038,In_2079,In_7);
or U1039 (N_1039,In_2426,In_1272);
nor U1040 (N_1040,In_802,In_1376);
nand U1041 (N_1041,In_1725,In_1739);
nor U1042 (N_1042,In_623,In_133);
or U1043 (N_1043,In_2334,In_1975);
xor U1044 (N_1044,In_164,In_1361);
and U1045 (N_1045,In_1086,In_148);
xor U1046 (N_1046,In_1094,In_1500);
or U1047 (N_1047,In_1658,In_2406);
nor U1048 (N_1048,In_1435,In_2179);
and U1049 (N_1049,In_118,In_1148);
or U1050 (N_1050,In_386,In_605);
and U1051 (N_1051,In_1040,In_2207);
nor U1052 (N_1052,In_1671,In_1064);
xnor U1053 (N_1053,In_2115,In_1135);
nor U1054 (N_1054,In_1864,In_1426);
or U1055 (N_1055,In_1711,In_2263);
and U1056 (N_1056,In_437,In_373);
and U1057 (N_1057,In_548,In_515);
or U1058 (N_1058,In_566,In_119);
xnor U1059 (N_1059,In_144,In_279);
nand U1060 (N_1060,In_2322,In_463);
nor U1061 (N_1061,In_636,In_863);
and U1062 (N_1062,In_1105,In_73);
nand U1063 (N_1063,In_1063,In_1907);
and U1064 (N_1064,In_1578,In_703);
and U1065 (N_1065,In_1138,In_1854);
and U1066 (N_1066,In_404,In_2225);
xnor U1067 (N_1067,In_1537,In_1747);
xnor U1068 (N_1068,In_1607,In_1645);
nand U1069 (N_1069,In_442,In_2007);
and U1070 (N_1070,In_157,In_1423);
or U1071 (N_1071,In_1974,In_899);
nor U1072 (N_1072,In_1259,In_1280);
and U1073 (N_1073,In_1248,In_1054);
nand U1074 (N_1074,In_766,In_2229);
and U1075 (N_1075,In_1853,In_1713);
nand U1076 (N_1076,In_640,In_2200);
nor U1077 (N_1077,In_1681,In_2277);
nand U1078 (N_1078,In_1993,In_2240);
or U1079 (N_1079,In_1926,In_1597);
nand U1080 (N_1080,In_269,In_400);
or U1081 (N_1081,In_1466,In_771);
or U1082 (N_1082,In_585,In_624);
xor U1083 (N_1083,In_2201,In_1028);
nor U1084 (N_1084,In_0,In_466);
nor U1085 (N_1085,In_1010,In_1059);
and U1086 (N_1086,In_319,In_813);
nand U1087 (N_1087,In_1068,In_705);
and U1088 (N_1088,In_741,In_2393);
nand U1089 (N_1089,In_2090,In_186);
and U1090 (N_1090,In_170,In_625);
and U1091 (N_1091,In_510,In_2245);
and U1092 (N_1092,In_1396,In_1245);
nor U1093 (N_1093,In_2407,In_2308);
xor U1094 (N_1094,In_200,In_1917);
nor U1095 (N_1095,In_1980,In_867);
or U1096 (N_1096,In_1632,In_134);
or U1097 (N_1097,In_1231,In_2166);
nor U1098 (N_1098,In_655,In_1982);
nor U1099 (N_1099,In_2170,In_2361);
nand U1100 (N_1100,In_84,In_1640);
and U1101 (N_1101,In_772,In_1781);
and U1102 (N_1102,In_1316,In_921);
nor U1103 (N_1103,In_1806,In_1399);
and U1104 (N_1104,In_1890,In_1305);
nand U1105 (N_1105,In_966,In_211);
nor U1106 (N_1106,In_1134,In_745);
xnor U1107 (N_1107,In_723,In_1338);
nor U1108 (N_1108,In_931,In_317);
or U1109 (N_1109,In_1963,In_1958);
nand U1110 (N_1110,In_857,In_2195);
xnor U1111 (N_1111,In_182,In_1432);
or U1112 (N_1112,In_2497,In_1940);
or U1113 (N_1113,In_121,In_1818);
nor U1114 (N_1114,In_2093,In_926);
xnor U1115 (N_1115,In_1031,In_1984);
or U1116 (N_1116,In_816,In_801);
and U1117 (N_1117,In_706,In_2428);
nand U1118 (N_1118,In_1986,In_1380);
and U1119 (N_1119,In_759,In_248);
and U1120 (N_1120,In_1712,In_2495);
or U1121 (N_1121,In_41,In_2416);
or U1122 (N_1122,In_2457,In_808);
nor U1123 (N_1123,In_2026,In_2083);
or U1124 (N_1124,In_337,In_2274);
xor U1125 (N_1125,In_333,In_831);
nor U1126 (N_1126,In_1395,In_174);
and U1127 (N_1127,In_225,In_742);
xor U1128 (N_1128,In_1463,In_50);
or U1129 (N_1129,In_1400,In_1493);
nor U1130 (N_1130,In_2198,In_30);
xor U1131 (N_1131,In_432,In_452);
xnor U1132 (N_1132,In_1743,In_1341);
nor U1133 (N_1133,In_94,In_1324);
and U1134 (N_1134,In_846,In_1628);
xnor U1135 (N_1135,In_283,In_630);
or U1136 (N_1136,In_2485,In_1644);
or U1137 (N_1137,In_920,In_1106);
or U1138 (N_1138,In_570,In_359);
and U1139 (N_1139,In_277,In_1906);
or U1140 (N_1140,In_1293,In_1944);
and U1141 (N_1141,In_559,In_1957);
xor U1142 (N_1142,In_727,In_408);
or U1143 (N_1143,In_1084,In_90);
nand U1144 (N_1144,In_471,In_74);
xnor U1145 (N_1145,In_2492,In_1960);
and U1146 (N_1146,In_2015,In_1103);
nor U1147 (N_1147,In_1803,In_158);
xor U1148 (N_1148,In_393,In_2372);
nor U1149 (N_1149,In_2186,In_1120);
or U1150 (N_1150,In_1587,In_1042);
nor U1151 (N_1151,In_1520,In_193);
xnor U1152 (N_1152,In_968,In_417);
and U1153 (N_1153,In_293,In_1846);
and U1154 (N_1154,In_2466,In_737);
or U1155 (N_1155,In_1167,In_1884);
or U1156 (N_1156,In_2448,In_876);
nand U1157 (N_1157,In_2022,In_2454);
xor U1158 (N_1158,In_2314,In_2380);
nand U1159 (N_1159,In_785,In_298);
nor U1160 (N_1160,In_297,In_57);
nor U1161 (N_1161,In_2219,In_538);
and U1162 (N_1162,In_1333,In_1230);
nor U1163 (N_1163,In_1365,In_965);
xor U1164 (N_1164,In_475,In_1017);
nand U1165 (N_1165,In_569,In_1445);
nand U1166 (N_1166,In_2143,In_1666);
nor U1167 (N_1167,In_1999,In_2430);
xor U1168 (N_1168,In_713,In_1302);
nand U1169 (N_1169,In_516,In_313);
xnor U1170 (N_1170,In_1964,In_1538);
and U1171 (N_1171,In_1685,In_1226);
nand U1172 (N_1172,In_889,In_1778);
and U1173 (N_1173,In_1699,In_223);
nand U1174 (N_1174,In_2264,In_502);
and U1175 (N_1175,In_606,In_371);
or U1176 (N_1176,In_1568,In_2271);
xnor U1177 (N_1177,In_521,In_2298);
nand U1178 (N_1178,In_2237,In_14);
or U1179 (N_1179,In_1404,In_1360);
and U1180 (N_1180,In_897,In_381);
xnor U1181 (N_1181,In_2335,In_848);
xnor U1182 (N_1182,In_1732,In_1234);
nor U1183 (N_1183,In_2111,In_1281);
nor U1184 (N_1184,In_1939,In_142);
nand U1185 (N_1185,In_901,In_551);
nand U1186 (N_1186,In_19,In_21);
or U1187 (N_1187,In_1401,In_2375);
or U1188 (N_1188,In_1943,In_1253);
and U1189 (N_1189,In_603,In_295);
xor U1190 (N_1190,In_1812,In_2134);
nand U1191 (N_1191,In_37,In_113);
xor U1192 (N_1192,In_365,In_2488);
and U1193 (N_1193,In_1098,In_324);
and U1194 (N_1194,In_354,In_1424);
xor U1195 (N_1195,In_67,In_173);
and U1196 (N_1196,In_2360,In_1636);
nor U1197 (N_1197,In_1991,In_1909);
xnor U1198 (N_1198,In_1065,In_2139);
or U1199 (N_1199,In_154,In_58);
or U1200 (N_1200,In_1938,In_216);
nand U1201 (N_1201,In_469,In_1740);
or U1202 (N_1202,In_735,In_1356);
or U1203 (N_1203,In_1590,In_485);
nor U1204 (N_1204,In_358,In_717);
or U1205 (N_1205,In_2078,In_567);
nor U1206 (N_1206,In_1470,In_1157);
or U1207 (N_1207,In_602,In_2484);
nand U1208 (N_1208,In_249,In_1209);
or U1209 (N_1209,In_1179,In_711);
xnor U1210 (N_1210,In_1397,In_1585);
xnor U1211 (N_1211,In_409,In_2128);
or U1212 (N_1212,In_1551,In_972);
xor U1213 (N_1213,In_2076,In_366);
or U1214 (N_1214,In_552,In_2177);
xnor U1215 (N_1215,In_2096,In_1706);
or U1216 (N_1216,In_788,In_1795);
nor U1217 (N_1217,In_535,In_2127);
or U1218 (N_1218,In_1625,In_2256);
nand U1219 (N_1219,In_2474,In_598);
nor U1220 (N_1220,In_111,In_1782);
or U1221 (N_1221,In_1162,In_1937);
nor U1222 (N_1222,In_1322,In_456);
or U1223 (N_1223,In_2233,In_2307);
nand U1224 (N_1224,In_1870,In_1136);
or U1225 (N_1225,In_1409,In_367);
xnor U1226 (N_1226,In_2124,In_993);
xnor U1227 (N_1227,In_1279,In_1770);
or U1228 (N_1228,In_821,In_2424);
and U1229 (N_1229,In_1730,In_1651);
and U1230 (N_1230,In_1995,In_1650);
and U1231 (N_1231,In_2048,In_1872);
or U1232 (N_1232,In_162,In_583);
nor U1233 (N_1233,In_1314,In_1276);
nor U1234 (N_1234,In_176,In_1808);
and U1235 (N_1235,In_2181,In_168);
and U1236 (N_1236,In_733,In_1486);
xnor U1237 (N_1237,In_461,In_2434);
nand U1238 (N_1238,In_1277,In_1637);
and U1239 (N_1239,In_753,In_609);
xnor U1240 (N_1240,In_963,In_2269);
nand U1241 (N_1241,In_858,In_321);
nand U1242 (N_1242,In_752,In_2325);
xor U1243 (N_1243,In_177,In_601);
nor U1244 (N_1244,In_2101,In_1667);
xor U1245 (N_1245,In_1317,In_2105);
nand U1246 (N_1246,In_1737,In_1144);
nand U1247 (N_1247,In_1427,In_1479);
xnor U1248 (N_1248,In_1152,In_833);
or U1249 (N_1249,In_2246,In_868);
and U1250 (N_1250,In_1190,In_1518);
nand U1251 (N_1251,In_2373,In_1983);
or U1252 (N_1252,In_2021,In_2408);
nor U1253 (N_1253,In_1968,In_1211);
xnor U1254 (N_1254,In_560,In_1067);
nand U1255 (N_1255,In_310,In_2438);
nor U1256 (N_1256,In_351,In_1851);
and U1257 (N_1257,In_1211,In_2478);
and U1258 (N_1258,In_893,In_2076);
or U1259 (N_1259,In_1616,In_582);
or U1260 (N_1260,In_1096,In_1556);
nand U1261 (N_1261,In_1286,In_1549);
and U1262 (N_1262,In_1524,In_2058);
xor U1263 (N_1263,In_60,In_1899);
nand U1264 (N_1264,In_1183,In_1755);
nand U1265 (N_1265,In_1328,In_2319);
or U1266 (N_1266,In_1515,In_443);
xor U1267 (N_1267,In_1630,In_2270);
nor U1268 (N_1268,In_135,In_1429);
or U1269 (N_1269,In_378,In_2066);
nor U1270 (N_1270,In_1910,In_1592);
and U1271 (N_1271,In_2173,In_166);
nor U1272 (N_1272,In_1014,In_607);
nand U1273 (N_1273,In_530,In_1223);
xor U1274 (N_1274,In_567,In_326);
nand U1275 (N_1275,In_2298,In_1777);
nor U1276 (N_1276,In_766,In_843);
nand U1277 (N_1277,In_425,In_1989);
nor U1278 (N_1278,In_211,In_1351);
and U1279 (N_1279,In_1195,In_2156);
nor U1280 (N_1280,In_618,In_562);
and U1281 (N_1281,In_1086,In_277);
or U1282 (N_1282,In_1255,In_2406);
and U1283 (N_1283,In_384,In_2110);
or U1284 (N_1284,In_1230,In_68);
and U1285 (N_1285,In_169,In_793);
or U1286 (N_1286,In_246,In_703);
nor U1287 (N_1287,In_1126,In_356);
xor U1288 (N_1288,In_954,In_2313);
nand U1289 (N_1289,In_2313,In_2368);
xor U1290 (N_1290,In_1805,In_855);
and U1291 (N_1291,In_424,In_1504);
nor U1292 (N_1292,In_672,In_683);
and U1293 (N_1293,In_1744,In_167);
or U1294 (N_1294,In_256,In_2427);
and U1295 (N_1295,In_15,In_2480);
nor U1296 (N_1296,In_1508,In_2141);
and U1297 (N_1297,In_1837,In_1813);
and U1298 (N_1298,In_278,In_2173);
or U1299 (N_1299,In_1045,In_2211);
xor U1300 (N_1300,In_996,In_775);
nand U1301 (N_1301,In_1912,In_107);
or U1302 (N_1302,In_73,In_311);
and U1303 (N_1303,In_1913,In_464);
and U1304 (N_1304,In_1227,In_1459);
xnor U1305 (N_1305,In_1739,In_1358);
nor U1306 (N_1306,In_2080,In_1296);
xor U1307 (N_1307,In_1627,In_2083);
xnor U1308 (N_1308,In_1686,In_495);
xor U1309 (N_1309,In_528,In_959);
or U1310 (N_1310,In_2176,In_2000);
nand U1311 (N_1311,In_83,In_1112);
xnor U1312 (N_1312,In_559,In_1883);
or U1313 (N_1313,In_1478,In_508);
xnor U1314 (N_1314,In_2169,In_1480);
nand U1315 (N_1315,In_286,In_1551);
or U1316 (N_1316,In_2231,In_109);
or U1317 (N_1317,In_684,In_1163);
xnor U1318 (N_1318,In_2359,In_1330);
nand U1319 (N_1319,In_2117,In_1922);
nor U1320 (N_1320,In_1100,In_2108);
nand U1321 (N_1321,In_2466,In_91);
nand U1322 (N_1322,In_146,In_2170);
nor U1323 (N_1323,In_938,In_43);
nand U1324 (N_1324,In_2215,In_2262);
nor U1325 (N_1325,In_1202,In_2163);
and U1326 (N_1326,In_2028,In_2229);
and U1327 (N_1327,In_725,In_1100);
nor U1328 (N_1328,In_1779,In_387);
nand U1329 (N_1329,In_439,In_2070);
xnor U1330 (N_1330,In_768,In_120);
xnor U1331 (N_1331,In_2489,In_1268);
or U1332 (N_1332,In_1828,In_2202);
and U1333 (N_1333,In_296,In_392);
xor U1334 (N_1334,In_1076,In_2089);
nor U1335 (N_1335,In_2077,In_1009);
or U1336 (N_1336,In_278,In_1933);
or U1337 (N_1337,In_1807,In_1696);
nor U1338 (N_1338,In_1631,In_978);
xnor U1339 (N_1339,In_1332,In_2255);
or U1340 (N_1340,In_911,In_609);
nand U1341 (N_1341,In_1526,In_1509);
or U1342 (N_1342,In_901,In_416);
or U1343 (N_1343,In_229,In_693);
nand U1344 (N_1344,In_1137,In_161);
nand U1345 (N_1345,In_2485,In_915);
or U1346 (N_1346,In_640,In_2433);
nor U1347 (N_1347,In_301,In_1743);
xor U1348 (N_1348,In_1269,In_411);
and U1349 (N_1349,In_1473,In_1082);
and U1350 (N_1350,In_489,In_1300);
or U1351 (N_1351,In_988,In_748);
nor U1352 (N_1352,In_1070,In_231);
xor U1353 (N_1353,In_1962,In_2276);
nand U1354 (N_1354,In_211,In_1257);
xor U1355 (N_1355,In_484,In_1717);
or U1356 (N_1356,In_2295,In_114);
xnor U1357 (N_1357,In_739,In_1487);
xor U1358 (N_1358,In_524,In_1395);
and U1359 (N_1359,In_2327,In_469);
or U1360 (N_1360,In_2359,In_1909);
and U1361 (N_1361,In_2119,In_1231);
nor U1362 (N_1362,In_647,In_1216);
or U1363 (N_1363,In_602,In_1275);
and U1364 (N_1364,In_1705,In_1027);
or U1365 (N_1365,In_1567,In_647);
or U1366 (N_1366,In_2053,In_1641);
xnor U1367 (N_1367,In_676,In_1019);
and U1368 (N_1368,In_2496,In_434);
or U1369 (N_1369,In_2152,In_2261);
or U1370 (N_1370,In_675,In_409);
or U1371 (N_1371,In_768,In_389);
and U1372 (N_1372,In_828,In_2167);
nor U1373 (N_1373,In_919,In_1744);
nor U1374 (N_1374,In_375,In_159);
or U1375 (N_1375,In_102,In_1820);
xor U1376 (N_1376,In_1226,In_1155);
or U1377 (N_1377,In_1389,In_1367);
nand U1378 (N_1378,In_295,In_93);
xnor U1379 (N_1379,In_1557,In_1385);
nand U1380 (N_1380,In_438,In_329);
nand U1381 (N_1381,In_66,In_1266);
nor U1382 (N_1382,In_1715,In_1351);
and U1383 (N_1383,In_336,In_1846);
nor U1384 (N_1384,In_809,In_863);
xnor U1385 (N_1385,In_1993,In_120);
or U1386 (N_1386,In_1604,In_4);
nand U1387 (N_1387,In_1978,In_770);
or U1388 (N_1388,In_1002,In_1916);
nor U1389 (N_1389,In_2029,In_532);
and U1390 (N_1390,In_790,In_791);
or U1391 (N_1391,In_984,In_689);
nor U1392 (N_1392,In_105,In_601);
nand U1393 (N_1393,In_2452,In_2261);
and U1394 (N_1394,In_977,In_2447);
and U1395 (N_1395,In_2198,In_1687);
and U1396 (N_1396,In_1446,In_1805);
or U1397 (N_1397,In_1902,In_33);
or U1398 (N_1398,In_184,In_1080);
nand U1399 (N_1399,In_930,In_80);
or U1400 (N_1400,In_866,In_148);
and U1401 (N_1401,In_2289,In_480);
or U1402 (N_1402,In_2347,In_725);
nand U1403 (N_1403,In_2373,In_108);
nor U1404 (N_1404,In_1134,In_859);
nand U1405 (N_1405,In_408,In_2494);
or U1406 (N_1406,In_48,In_40);
nand U1407 (N_1407,In_2243,In_630);
nor U1408 (N_1408,In_2321,In_1437);
or U1409 (N_1409,In_1445,In_1690);
xnor U1410 (N_1410,In_1825,In_2261);
nand U1411 (N_1411,In_67,In_171);
nor U1412 (N_1412,In_1871,In_1207);
xor U1413 (N_1413,In_944,In_336);
nor U1414 (N_1414,In_2494,In_501);
nand U1415 (N_1415,In_301,In_199);
nand U1416 (N_1416,In_863,In_29);
xor U1417 (N_1417,In_269,In_1628);
nor U1418 (N_1418,In_900,In_2427);
and U1419 (N_1419,In_908,In_2056);
or U1420 (N_1420,In_881,In_378);
or U1421 (N_1421,In_1203,In_1055);
and U1422 (N_1422,In_36,In_528);
or U1423 (N_1423,In_2471,In_450);
or U1424 (N_1424,In_1395,In_1327);
nand U1425 (N_1425,In_1071,In_1021);
xnor U1426 (N_1426,In_495,In_1142);
nand U1427 (N_1427,In_376,In_2195);
xnor U1428 (N_1428,In_1582,In_1276);
nor U1429 (N_1429,In_1530,In_1845);
nand U1430 (N_1430,In_882,In_2370);
nor U1431 (N_1431,In_176,In_423);
or U1432 (N_1432,In_326,In_525);
nand U1433 (N_1433,In_2137,In_276);
nor U1434 (N_1434,In_89,In_573);
and U1435 (N_1435,In_412,In_512);
and U1436 (N_1436,In_652,In_2035);
xor U1437 (N_1437,In_1370,In_1220);
nor U1438 (N_1438,In_1616,In_1350);
nand U1439 (N_1439,In_2491,In_2022);
xnor U1440 (N_1440,In_2199,In_1010);
xnor U1441 (N_1441,In_1893,In_2056);
nand U1442 (N_1442,In_477,In_1935);
and U1443 (N_1443,In_2338,In_949);
and U1444 (N_1444,In_2441,In_1821);
nand U1445 (N_1445,In_799,In_1869);
nand U1446 (N_1446,In_1979,In_1394);
nand U1447 (N_1447,In_1494,In_2462);
and U1448 (N_1448,In_2105,In_619);
and U1449 (N_1449,In_1827,In_2134);
nand U1450 (N_1450,In_622,In_487);
xnor U1451 (N_1451,In_411,In_2493);
and U1452 (N_1452,In_2223,In_2033);
or U1453 (N_1453,In_467,In_2220);
or U1454 (N_1454,In_2417,In_1030);
and U1455 (N_1455,In_178,In_1509);
and U1456 (N_1456,In_2096,In_1546);
nor U1457 (N_1457,In_721,In_2390);
and U1458 (N_1458,In_2347,In_1198);
xor U1459 (N_1459,In_2158,In_2196);
or U1460 (N_1460,In_893,In_1816);
nand U1461 (N_1461,In_413,In_97);
nor U1462 (N_1462,In_933,In_1354);
or U1463 (N_1463,In_1970,In_1117);
or U1464 (N_1464,In_1664,In_2149);
nand U1465 (N_1465,In_772,In_1786);
or U1466 (N_1466,In_1227,In_1435);
xnor U1467 (N_1467,In_105,In_242);
and U1468 (N_1468,In_2175,In_369);
xnor U1469 (N_1469,In_1041,In_2205);
or U1470 (N_1470,In_1952,In_312);
and U1471 (N_1471,In_187,In_318);
nor U1472 (N_1472,In_128,In_537);
xnor U1473 (N_1473,In_1837,In_1386);
xor U1474 (N_1474,In_191,In_1308);
and U1475 (N_1475,In_2339,In_2005);
and U1476 (N_1476,In_790,In_2085);
and U1477 (N_1477,In_1205,In_2248);
nand U1478 (N_1478,In_1786,In_1281);
nand U1479 (N_1479,In_990,In_1572);
or U1480 (N_1480,In_2009,In_2121);
nand U1481 (N_1481,In_2083,In_856);
nand U1482 (N_1482,In_694,In_309);
or U1483 (N_1483,In_1188,In_240);
xor U1484 (N_1484,In_996,In_1476);
nand U1485 (N_1485,In_739,In_1253);
nand U1486 (N_1486,In_578,In_822);
and U1487 (N_1487,In_504,In_532);
and U1488 (N_1488,In_1222,In_2038);
nand U1489 (N_1489,In_476,In_1945);
nand U1490 (N_1490,In_92,In_2321);
xnor U1491 (N_1491,In_2005,In_397);
nand U1492 (N_1492,In_1064,In_611);
and U1493 (N_1493,In_2354,In_150);
or U1494 (N_1494,In_956,In_1062);
nand U1495 (N_1495,In_154,In_602);
or U1496 (N_1496,In_1721,In_815);
or U1497 (N_1497,In_848,In_1307);
or U1498 (N_1498,In_705,In_321);
xnor U1499 (N_1499,In_1714,In_553);
or U1500 (N_1500,In_2323,In_65);
or U1501 (N_1501,In_363,In_345);
nor U1502 (N_1502,In_1562,In_252);
or U1503 (N_1503,In_2200,In_1051);
or U1504 (N_1504,In_979,In_322);
or U1505 (N_1505,In_806,In_852);
nor U1506 (N_1506,In_610,In_2440);
nor U1507 (N_1507,In_1469,In_1610);
nor U1508 (N_1508,In_1435,In_1953);
nand U1509 (N_1509,In_2211,In_581);
nand U1510 (N_1510,In_1175,In_1314);
nand U1511 (N_1511,In_2129,In_1293);
nor U1512 (N_1512,In_2397,In_1421);
nand U1513 (N_1513,In_165,In_256);
xnor U1514 (N_1514,In_272,In_1909);
or U1515 (N_1515,In_1923,In_474);
nor U1516 (N_1516,In_843,In_1957);
xor U1517 (N_1517,In_104,In_2044);
xnor U1518 (N_1518,In_2243,In_1655);
nand U1519 (N_1519,In_994,In_920);
or U1520 (N_1520,In_938,In_1539);
nor U1521 (N_1521,In_1480,In_111);
and U1522 (N_1522,In_2086,In_444);
xnor U1523 (N_1523,In_443,In_129);
nand U1524 (N_1524,In_1696,In_779);
xnor U1525 (N_1525,In_55,In_2324);
xnor U1526 (N_1526,In_1258,In_94);
nand U1527 (N_1527,In_737,In_232);
nor U1528 (N_1528,In_538,In_1376);
or U1529 (N_1529,In_319,In_1462);
xnor U1530 (N_1530,In_939,In_1800);
xor U1531 (N_1531,In_344,In_565);
or U1532 (N_1532,In_657,In_1450);
xor U1533 (N_1533,In_1141,In_1164);
or U1534 (N_1534,In_91,In_1824);
or U1535 (N_1535,In_639,In_2394);
nor U1536 (N_1536,In_1363,In_613);
and U1537 (N_1537,In_843,In_2341);
and U1538 (N_1538,In_361,In_445);
nor U1539 (N_1539,In_1521,In_329);
and U1540 (N_1540,In_270,In_284);
xnor U1541 (N_1541,In_1385,In_910);
or U1542 (N_1542,In_1780,In_13);
xnor U1543 (N_1543,In_2000,In_1252);
and U1544 (N_1544,In_1431,In_1115);
nor U1545 (N_1545,In_2086,In_1256);
or U1546 (N_1546,In_1583,In_676);
nor U1547 (N_1547,In_564,In_1210);
and U1548 (N_1548,In_510,In_891);
xor U1549 (N_1549,In_2019,In_2187);
nand U1550 (N_1550,In_56,In_396);
nand U1551 (N_1551,In_625,In_2068);
and U1552 (N_1552,In_844,In_1125);
and U1553 (N_1553,In_1441,In_840);
and U1554 (N_1554,In_283,In_177);
or U1555 (N_1555,In_1536,In_13);
xnor U1556 (N_1556,In_2145,In_1437);
nor U1557 (N_1557,In_668,In_637);
or U1558 (N_1558,In_1870,In_1890);
nand U1559 (N_1559,In_2352,In_1856);
nor U1560 (N_1560,In_2478,In_1193);
nor U1561 (N_1561,In_1071,In_703);
nand U1562 (N_1562,In_1950,In_2022);
nor U1563 (N_1563,In_917,In_2200);
xor U1564 (N_1564,In_784,In_2098);
xor U1565 (N_1565,In_1484,In_1038);
nor U1566 (N_1566,In_1233,In_1522);
xnor U1567 (N_1567,In_1196,In_1657);
nand U1568 (N_1568,In_241,In_2279);
nor U1569 (N_1569,In_2109,In_2166);
nor U1570 (N_1570,In_1981,In_1562);
or U1571 (N_1571,In_654,In_1134);
and U1572 (N_1572,In_1087,In_1535);
nand U1573 (N_1573,In_1029,In_1477);
or U1574 (N_1574,In_1210,In_1043);
or U1575 (N_1575,In_1388,In_1166);
nand U1576 (N_1576,In_603,In_1997);
nor U1577 (N_1577,In_1793,In_510);
xor U1578 (N_1578,In_2277,In_1777);
nor U1579 (N_1579,In_1725,In_1298);
or U1580 (N_1580,In_253,In_307);
xor U1581 (N_1581,In_466,In_262);
or U1582 (N_1582,In_371,In_2173);
nor U1583 (N_1583,In_475,In_733);
and U1584 (N_1584,In_2195,In_820);
nor U1585 (N_1585,In_231,In_2032);
or U1586 (N_1586,In_2171,In_2106);
or U1587 (N_1587,In_451,In_2335);
nand U1588 (N_1588,In_1330,In_1312);
or U1589 (N_1589,In_434,In_2346);
xnor U1590 (N_1590,In_2270,In_1811);
or U1591 (N_1591,In_1049,In_2333);
nor U1592 (N_1592,In_1939,In_2360);
or U1593 (N_1593,In_311,In_394);
nor U1594 (N_1594,In_1384,In_355);
nor U1595 (N_1595,In_1182,In_121);
nor U1596 (N_1596,In_1029,In_2186);
or U1597 (N_1597,In_1021,In_1042);
nand U1598 (N_1598,In_2284,In_1706);
nand U1599 (N_1599,In_571,In_105);
nor U1600 (N_1600,In_2210,In_1310);
nor U1601 (N_1601,In_122,In_1936);
or U1602 (N_1602,In_1994,In_2314);
or U1603 (N_1603,In_1581,In_2402);
or U1604 (N_1604,In_1715,In_1067);
nor U1605 (N_1605,In_204,In_382);
xnor U1606 (N_1606,In_653,In_1588);
and U1607 (N_1607,In_587,In_2471);
and U1608 (N_1608,In_734,In_222);
and U1609 (N_1609,In_1086,In_12);
nand U1610 (N_1610,In_1093,In_1264);
or U1611 (N_1611,In_923,In_105);
or U1612 (N_1612,In_2483,In_2221);
nor U1613 (N_1613,In_1000,In_922);
and U1614 (N_1614,In_140,In_879);
or U1615 (N_1615,In_2480,In_1931);
nand U1616 (N_1616,In_1538,In_2045);
xnor U1617 (N_1617,In_1624,In_1104);
nand U1618 (N_1618,In_1248,In_541);
and U1619 (N_1619,In_1770,In_858);
or U1620 (N_1620,In_1017,In_2390);
or U1621 (N_1621,In_1215,In_1468);
and U1622 (N_1622,In_230,In_180);
nor U1623 (N_1623,In_2487,In_170);
or U1624 (N_1624,In_2148,In_2137);
and U1625 (N_1625,In_1321,In_1934);
or U1626 (N_1626,In_990,In_2099);
or U1627 (N_1627,In_117,In_1441);
nor U1628 (N_1628,In_2464,In_1710);
xnor U1629 (N_1629,In_1829,In_1164);
and U1630 (N_1630,In_1084,In_1970);
nor U1631 (N_1631,In_1264,In_1162);
or U1632 (N_1632,In_815,In_2441);
nand U1633 (N_1633,In_2323,In_359);
nand U1634 (N_1634,In_1701,In_1044);
or U1635 (N_1635,In_1194,In_1934);
xnor U1636 (N_1636,In_301,In_1075);
and U1637 (N_1637,In_1071,In_1262);
xor U1638 (N_1638,In_335,In_2159);
or U1639 (N_1639,In_1345,In_2401);
or U1640 (N_1640,In_1520,In_81);
nand U1641 (N_1641,In_1007,In_261);
or U1642 (N_1642,In_2485,In_699);
nor U1643 (N_1643,In_570,In_904);
or U1644 (N_1644,In_2071,In_1418);
and U1645 (N_1645,In_1387,In_2324);
xnor U1646 (N_1646,In_1202,In_783);
and U1647 (N_1647,In_2419,In_103);
nor U1648 (N_1648,In_2233,In_79);
or U1649 (N_1649,In_1894,In_1234);
or U1650 (N_1650,In_1253,In_394);
and U1651 (N_1651,In_1776,In_933);
or U1652 (N_1652,In_2393,In_2077);
nand U1653 (N_1653,In_2377,In_2474);
or U1654 (N_1654,In_861,In_1514);
xnor U1655 (N_1655,In_1603,In_1281);
and U1656 (N_1656,In_783,In_1234);
or U1657 (N_1657,In_1171,In_1754);
xnor U1658 (N_1658,In_773,In_1731);
or U1659 (N_1659,In_2155,In_1556);
and U1660 (N_1660,In_468,In_2395);
and U1661 (N_1661,In_352,In_2133);
or U1662 (N_1662,In_2039,In_1735);
nand U1663 (N_1663,In_1157,In_1666);
or U1664 (N_1664,In_1565,In_951);
nor U1665 (N_1665,In_45,In_741);
and U1666 (N_1666,In_101,In_1461);
nor U1667 (N_1667,In_1388,In_745);
and U1668 (N_1668,In_2109,In_1007);
xor U1669 (N_1669,In_2422,In_473);
or U1670 (N_1670,In_1653,In_1038);
nor U1671 (N_1671,In_1622,In_2321);
xnor U1672 (N_1672,In_1178,In_552);
xor U1673 (N_1673,In_797,In_403);
xor U1674 (N_1674,In_49,In_964);
nand U1675 (N_1675,In_1345,In_1321);
or U1676 (N_1676,In_2275,In_570);
nand U1677 (N_1677,In_1349,In_1695);
or U1678 (N_1678,In_2118,In_1789);
xor U1679 (N_1679,In_2118,In_1753);
and U1680 (N_1680,In_722,In_1730);
nand U1681 (N_1681,In_1957,In_2059);
xnor U1682 (N_1682,In_777,In_2296);
nor U1683 (N_1683,In_475,In_2065);
xor U1684 (N_1684,In_1284,In_1578);
nor U1685 (N_1685,In_920,In_2426);
nor U1686 (N_1686,In_1936,In_107);
nand U1687 (N_1687,In_2219,In_516);
xor U1688 (N_1688,In_944,In_20);
nor U1689 (N_1689,In_2179,In_657);
and U1690 (N_1690,In_667,In_676);
xor U1691 (N_1691,In_2464,In_1657);
xnor U1692 (N_1692,In_1858,In_1402);
and U1693 (N_1693,In_2220,In_2394);
nor U1694 (N_1694,In_1267,In_462);
or U1695 (N_1695,In_1542,In_1616);
xnor U1696 (N_1696,In_1504,In_1730);
nand U1697 (N_1697,In_622,In_1238);
and U1698 (N_1698,In_2108,In_1973);
xnor U1699 (N_1699,In_1975,In_664);
nor U1700 (N_1700,In_1886,In_1334);
xor U1701 (N_1701,In_1569,In_502);
nand U1702 (N_1702,In_791,In_1420);
xnor U1703 (N_1703,In_553,In_2187);
xnor U1704 (N_1704,In_1876,In_1068);
xor U1705 (N_1705,In_510,In_1034);
and U1706 (N_1706,In_573,In_802);
xor U1707 (N_1707,In_420,In_417);
nand U1708 (N_1708,In_1868,In_278);
xor U1709 (N_1709,In_1318,In_416);
nor U1710 (N_1710,In_1487,In_1242);
xnor U1711 (N_1711,In_622,In_1192);
and U1712 (N_1712,In_1901,In_1333);
or U1713 (N_1713,In_1660,In_528);
and U1714 (N_1714,In_1900,In_837);
and U1715 (N_1715,In_170,In_852);
nor U1716 (N_1716,In_50,In_1540);
and U1717 (N_1717,In_347,In_664);
or U1718 (N_1718,In_997,In_1565);
nand U1719 (N_1719,In_244,In_1937);
xor U1720 (N_1720,In_1934,In_1307);
nor U1721 (N_1721,In_1375,In_1420);
and U1722 (N_1722,In_2086,In_1945);
or U1723 (N_1723,In_2195,In_590);
nor U1724 (N_1724,In_1033,In_2406);
nor U1725 (N_1725,In_1521,In_402);
xnor U1726 (N_1726,In_2199,In_586);
or U1727 (N_1727,In_2188,In_976);
nand U1728 (N_1728,In_1325,In_196);
xnor U1729 (N_1729,In_1523,In_693);
xnor U1730 (N_1730,In_1886,In_1757);
or U1731 (N_1731,In_1216,In_1563);
nor U1732 (N_1732,In_1558,In_1868);
nand U1733 (N_1733,In_730,In_639);
or U1734 (N_1734,In_1378,In_875);
nand U1735 (N_1735,In_189,In_1754);
nor U1736 (N_1736,In_1331,In_1967);
or U1737 (N_1737,In_2085,In_2463);
nand U1738 (N_1738,In_2350,In_1685);
nor U1739 (N_1739,In_664,In_1641);
or U1740 (N_1740,In_193,In_427);
nor U1741 (N_1741,In_1831,In_235);
and U1742 (N_1742,In_2443,In_1012);
nand U1743 (N_1743,In_884,In_1216);
nor U1744 (N_1744,In_283,In_256);
xnor U1745 (N_1745,In_764,In_1150);
or U1746 (N_1746,In_1210,In_2047);
xor U1747 (N_1747,In_1472,In_587);
nor U1748 (N_1748,In_1856,In_23);
or U1749 (N_1749,In_2060,In_742);
nor U1750 (N_1750,In_260,In_81);
nand U1751 (N_1751,In_78,In_981);
and U1752 (N_1752,In_1482,In_1337);
nor U1753 (N_1753,In_1017,In_2160);
nand U1754 (N_1754,In_1586,In_375);
nor U1755 (N_1755,In_2036,In_2267);
or U1756 (N_1756,In_2108,In_1907);
nor U1757 (N_1757,In_159,In_1317);
and U1758 (N_1758,In_1119,In_910);
nand U1759 (N_1759,In_1866,In_1130);
nor U1760 (N_1760,In_1580,In_219);
nand U1761 (N_1761,In_311,In_2366);
nor U1762 (N_1762,In_0,In_2229);
nor U1763 (N_1763,In_2045,In_653);
or U1764 (N_1764,In_201,In_902);
nand U1765 (N_1765,In_2314,In_1995);
xnor U1766 (N_1766,In_2102,In_52);
nor U1767 (N_1767,In_848,In_1265);
and U1768 (N_1768,In_1698,In_520);
and U1769 (N_1769,In_1734,In_1725);
nor U1770 (N_1770,In_590,In_2266);
or U1771 (N_1771,In_1107,In_1945);
or U1772 (N_1772,In_1226,In_882);
nand U1773 (N_1773,In_1460,In_1404);
nor U1774 (N_1774,In_1923,In_2101);
nor U1775 (N_1775,In_420,In_1927);
and U1776 (N_1776,In_1576,In_1868);
nand U1777 (N_1777,In_92,In_390);
and U1778 (N_1778,In_1543,In_922);
nor U1779 (N_1779,In_1593,In_519);
and U1780 (N_1780,In_1458,In_812);
nand U1781 (N_1781,In_343,In_947);
nand U1782 (N_1782,In_1601,In_2266);
nor U1783 (N_1783,In_1849,In_482);
xor U1784 (N_1784,In_39,In_1579);
xnor U1785 (N_1785,In_2102,In_215);
and U1786 (N_1786,In_210,In_1614);
xnor U1787 (N_1787,In_1884,In_1219);
or U1788 (N_1788,In_105,In_1062);
nor U1789 (N_1789,In_930,In_675);
or U1790 (N_1790,In_2221,In_2329);
xnor U1791 (N_1791,In_2176,In_733);
nand U1792 (N_1792,In_409,In_221);
xor U1793 (N_1793,In_496,In_961);
xor U1794 (N_1794,In_1138,In_181);
xor U1795 (N_1795,In_278,In_783);
and U1796 (N_1796,In_213,In_716);
or U1797 (N_1797,In_1933,In_2183);
and U1798 (N_1798,In_2342,In_231);
nor U1799 (N_1799,In_2128,In_1426);
xor U1800 (N_1800,In_1489,In_579);
nand U1801 (N_1801,In_177,In_176);
or U1802 (N_1802,In_1415,In_865);
xor U1803 (N_1803,In_228,In_2126);
nor U1804 (N_1804,In_2383,In_213);
nand U1805 (N_1805,In_415,In_1565);
or U1806 (N_1806,In_1152,In_211);
nor U1807 (N_1807,In_1835,In_1078);
nor U1808 (N_1808,In_1249,In_76);
and U1809 (N_1809,In_2464,In_719);
nor U1810 (N_1810,In_1458,In_1477);
nand U1811 (N_1811,In_2475,In_2339);
nor U1812 (N_1812,In_1725,In_1604);
or U1813 (N_1813,In_2217,In_1876);
and U1814 (N_1814,In_2447,In_931);
nand U1815 (N_1815,In_332,In_1943);
or U1816 (N_1816,In_2061,In_1464);
xor U1817 (N_1817,In_524,In_1844);
xor U1818 (N_1818,In_1402,In_1346);
xor U1819 (N_1819,In_1954,In_1009);
and U1820 (N_1820,In_2072,In_445);
or U1821 (N_1821,In_493,In_1046);
nand U1822 (N_1822,In_1664,In_1909);
or U1823 (N_1823,In_2382,In_1023);
and U1824 (N_1824,In_601,In_375);
or U1825 (N_1825,In_2478,In_1590);
nor U1826 (N_1826,In_1850,In_735);
nand U1827 (N_1827,In_164,In_1384);
nor U1828 (N_1828,In_378,In_1848);
nand U1829 (N_1829,In_1988,In_1433);
and U1830 (N_1830,In_462,In_1476);
and U1831 (N_1831,In_730,In_635);
nor U1832 (N_1832,In_267,In_1236);
nor U1833 (N_1833,In_2246,In_2151);
xor U1834 (N_1834,In_2218,In_1946);
and U1835 (N_1835,In_2124,In_1112);
or U1836 (N_1836,In_78,In_1168);
and U1837 (N_1837,In_184,In_2349);
nand U1838 (N_1838,In_1548,In_18);
and U1839 (N_1839,In_2076,In_1591);
nor U1840 (N_1840,In_1479,In_1380);
nor U1841 (N_1841,In_217,In_1990);
or U1842 (N_1842,In_1068,In_575);
or U1843 (N_1843,In_1226,In_538);
nand U1844 (N_1844,In_1814,In_936);
nand U1845 (N_1845,In_464,In_1205);
nor U1846 (N_1846,In_212,In_587);
xor U1847 (N_1847,In_2244,In_407);
nor U1848 (N_1848,In_2351,In_194);
nand U1849 (N_1849,In_112,In_339);
nor U1850 (N_1850,In_1995,In_1635);
xor U1851 (N_1851,In_1892,In_916);
xor U1852 (N_1852,In_1458,In_1182);
nand U1853 (N_1853,In_2176,In_241);
nand U1854 (N_1854,In_2362,In_923);
xor U1855 (N_1855,In_1982,In_1777);
and U1856 (N_1856,In_536,In_1581);
nand U1857 (N_1857,In_2124,In_1002);
or U1858 (N_1858,In_2087,In_2241);
or U1859 (N_1859,In_377,In_332);
and U1860 (N_1860,In_1686,In_1615);
or U1861 (N_1861,In_1671,In_1802);
nor U1862 (N_1862,In_330,In_817);
nor U1863 (N_1863,In_784,In_390);
xor U1864 (N_1864,In_456,In_1514);
nand U1865 (N_1865,In_494,In_752);
nand U1866 (N_1866,In_851,In_2398);
and U1867 (N_1867,In_668,In_627);
nand U1868 (N_1868,In_1390,In_2065);
and U1869 (N_1869,In_1581,In_72);
or U1870 (N_1870,In_555,In_2005);
nand U1871 (N_1871,In_1169,In_429);
or U1872 (N_1872,In_345,In_2289);
xnor U1873 (N_1873,In_1579,In_718);
xor U1874 (N_1874,In_1449,In_605);
and U1875 (N_1875,In_1648,In_1777);
nor U1876 (N_1876,In_982,In_326);
xor U1877 (N_1877,In_1679,In_611);
nand U1878 (N_1878,In_1138,In_560);
and U1879 (N_1879,In_1404,In_1738);
xnor U1880 (N_1880,In_104,In_1532);
and U1881 (N_1881,In_326,In_642);
and U1882 (N_1882,In_666,In_1768);
nor U1883 (N_1883,In_662,In_608);
nor U1884 (N_1884,In_2245,In_993);
nor U1885 (N_1885,In_1382,In_1677);
or U1886 (N_1886,In_436,In_966);
and U1887 (N_1887,In_2325,In_1198);
or U1888 (N_1888,In_138,In_2107);
or U1889 (N_1889,In_68,In_2048);
xnor U1890 (N_1890,In_1616,In_1757);
nor U1891 (N_1891,In_1682,In_517);
nor U1892 (N_1892,In_1088,In_1886);
and U1893 (N_1893,In_1866,In_168);
and U1894 (N_1894,In_1928,In_2013);
xor U1895 (N_1895,In_925,In_2336);
nand U1896 (N_1896,In_2237,In_2150);
nand U1897 (N_1897,In_2104,In_1818);
nand U1898 (N_1898,In_946,In_775);
or U1899 (N_1899,In_1933,In_454);
and U1900 (N_1900,In_642,In_1566);
xnor U1901 (N_1901,In_483,In_2365);
or U1902 (N_1902,In_443,In_1103);
nand U1903 (N_1903,In_2435,In_830);
xnor U1904 (N_1904,In_673,In_2095);
and U1905 (N_1905,In_816,In_2129);
and U1906 (N_1906,In_1575,In_949);
nor U1907 (N_1907,In_780,In_1181);
nor U1908 (N_1908,In_1402,In_2488);
xor U1909 (N_1909,In_1863,In_5);
nor U1910 (N_1910,In_1969,In_227);
or U1911 (N_1911,In_2326,In_346);
and U1912 (N_1912,In_1098,In_587);
and U1913 (N_1913,In_320,In_2025);
nand U1914 (N_1914,In_110,In_604);
or U1915 (N_1915,In_1139,In_2260);
or U1916 (N_1916,In_1136,In_476);
nand U1917 (N_1917,In_1616,In_1742);
xor U1918 (N_1918,In_1695,In_2469);
and U1919 (N_1919,In_1283,In_2345);
or U1920 (N_1920,In_2304,In_126);
and U1921 (N_1921,In_121,In_1676);
nand U1922 (N_1922,In_420,In_1958);
nand U1923 (N_1923,In_595,In_1769);
nand U1924 (N_1924,In_285,In_1827);
and U1925 (N_1925,In_2453,In_1186);
and U1926 (N_1926,In_2471,In_919);
xor U1927 (N_1927,In_1696,In_144);
or U1928 (N_1928,In_1852,In_1554);
and U1929 (N_1929,In_386,In_1818);
or U1930 (N_1930,In_1821,In_1431);
or U1931 (N_1931,In_1286,In_336);
and U1932 (N_1932,In_2048,In_2353);
nand U1933 (N_1933,In_6,In_267);
xnor U1934 (N_1934,In_2244,In_1882);
or U1935 (N_1935,In_98,In_2095);
nand U1936 (N_1936,In_1699,In_765);
or U1937 (N_1937,In_2362,In_672);
or U1938 (N_1938,In_1002,In_2428);
and U1939 (N_1939,In_843,In_1977);
xnor U1940 (N_1940,In_2396,In_1417);
xnor U1941 (N_1941,In_2112,In_2273);
nand U1942 (N_1942,In_1276,In_907);
nand U1943 (N_1943,In_1173,In_1839);
xor U1944 (N_1944,In_2350,In_1650);
nand U1945 (N_1945,In_415,In_1642);
and U1946 (N_1946,In_23,In_2345);
and U1947 (N_1947,In_1027,In_1293);
nor U1948 (N_1948,In_1198,In_298);
nor U1949 (N_1949,In_499,In_1175);
nand U1950 (N_1950,In_1357,In_1489);
xnor U1951 (N_1951,In_1123,In_975);
nor U1952 (N_1952,In_2055,In_1770);
nor U1953 (N_1953,In_439,In_2325);
or U1954 (N_1954,In_304,In_89);
nand U1955 (N_1955,In_836,In_459);
nand U1956 (N_1956,In_266,In_2361);
or U1957 (N_1957,In_974,In_260);
nor U1958 (N_1958,In_2062,In_1406);
nand U1959 (N_1959,In_2102,In_1054);
and U1960 (N_1960,In_2316,In_154);
or U1961 (N_1961,In_1997,In_2355);
xor U1962 (N_1962,In_1628,In_1848);
xnor U1963 (N_1963,In_2078,In_577);
nor U1964 (N_1964,In_1890,In_2220);
nor U1965 (N_1965,In_2184,In_305);
nor U1966 (N_1966,In_605,In_280);
nand U1967 (N_1967,In_2213,In_1862);
and U1968 (N_1968,In_611,In_1093);
or U1969 (N_1969,In_2129,In_610);
and U1970 (N_1970,In_1435,In_276);
nand U1971 (N_1971,In_1930,In_853);
xor U1972 (N_1972,In_920,In_1370);
xnor U1973 (N_1973,In_360,In_1088);
or U1974 (N_1974,In_528,In_1241);
nand U1975 (N_1975,In_776,In_396);
and U1976 (N_1976,In_2318,In_721);
xor U1977 (N_1977,In_1131,In_235);
or U1978 (N_1978,In_1063,In_1332);
xor U1979 (N_1979,In_2188,In_2134);
nand U1980 (N_1980,In_765,In_865);
and U1981 (N_1981,In_972,In_891);
or U1982 (N_1982,In_1128,In_47);
nand U1983 (N_1983,In_2285,In_960);
and U1984 (N_1984,In_1652,In_440);
xor U1985 (N_1985,In_408,In_1353);
nand U1986 (N_1986,In_1450,In_852);
xor U1987 (N_1987,In_2078,In_377);
nor U1988 (N_1988,In_2435,In_1162);
or U1989 (N_1989,In_881,In_335);
nor U1990 (N_1990,In_1755,In_420);
nor U1991 (N_1991,In_728,In_197);
nand U1992 (N_1992,In_2408,In_2028);
nand U1993 (N_1993,In_1886,In_1522);
xnor U1994 (N_1994,In_1666,In_302);
or U1995 (N_1995,In_157,In_546);
or U1996 (N_1996,In_2372,In_2445);
nor U1997 (N_1997,In_438,In_2150);
nor U1998 (N_1998,In_1658,In_1602);
or U1999 (N_1999,In_1326,In_952);
and U2000 (N_2000,In_2138,In_1785);
and U2001 (N_2001,In_1211,In_375);
or U2002 (N_2002,In_2042,In_438);
nand U2003 (N_2003,In_2369,In_474);
and U2004 (N_2004,In_437,In_208);
or U2005 (N_2005,In_329,In_1294);
xor U2006 (N_2006,In_751,In_2349);
and U2007 (N_2007,In_2124,In_774);
or U2008 (N_2008,In_838,In_567);
xnor U2009 (N_2009,In_1982,In_68);
or U2010 (N_2010,In_839,In_308);
and U2011 (N_2011,In_1931,In_59);
or U2012 (N_2012,In_1832,In_124);
nand U2013 (N_2013,In_2388,In_582);
xor U2014 (N_2014,In_308,In_1931);
xor U2015 (N_2015,In_233,In_1116);
and U2016 (N_2016,In_1317,In_467);
nand U2017 (N_2017,In_2212,In_283);
and U2018 (N_2018,In_1775,In_1639);
nor U2019 (N_2019,In_666,In_1903);
nor U2020 (N_2020,In_861,In_2111);
or U2021 (N_2021,In_939,In_1603);
nand U2022 (N_2022,In_462,In_692);
nand U2023 (N_2023,In_1998,In_552);
nand U2024 (N_2024,In_464,In_1536);
or U2025 (N_2025,In_736,In_131);
and U2026 (N_2026,In_2092,In_2372);
xor U2027 (N_2027,In_2047,In_2312);
and U2028 (N_2028,In_2208,In_859);
or U2029 (N_2029,In_328,In_1403);
or U2030 (N_2030,In_90,In_135);
xnor U2031 (N_2031,In_922,In_1557);
nor U2032 (N_2032,In_1647,In_1144);
or U2033 (N_2033,In_1065,In_488);
xor U2034 (N_2034,In_969,In_1439);
xnor U2035 (N_2035,In_522,In_273);
and U2036 (N_2036,In_1342,In_891);
xnor U2037 (N_2037,In_872,In_2215);
nor U2038 (N_2038,In_2333,In_215);
nor U2039 (N_2039,In_213,In_2085);
and U2040 (N_2040,In_1377,In_1390);
xor U2041 (N_2041,In_1833,In_451);
and U2042 (N_2042,In_389,In_1352);
and U2043 (N_2043,In_1008,In_586);
nand U2044 (N_2044,In_2036,In_980);
or U2045 (N_2045,In_1140,In_513);
xor U2046 (N_2046,In_555,In_194);
nor U2047 (N_2047,In_1541,In_2368);
nand U2048 (N_2048,In_72,In_1309);
xor U2049 (N_2049,In_1344,In_83);
or U2050 (N_2050,In_1048,In_1550);
nand U2051 (N_2051,In_1562,In_774);
or U2052 (N_2052,In_805,In_1792);
or U2053 (N_2053,In_1823,In_178);
or U2054 (N_2054,In_2346,In_516);
xor U2055 (N_2055,In_1439,In_611);
nand U2056 (N_2056,In_627,In_1179);
xnor U2057 (N_2057,In_2345,In_1568);
nor U2058 (N_2058,In_206,In_1188);
nor U2059 (N_2059,In_181,In_66);
nand U2060 (N_2060,In_2187,In_1945);
or U2061 (N_2061,In_2422,In_1743);
xnor U2062 (N_2062,In_1394,In_457);
or U2063 (N_2063,In_869,In_1792);
or U2064 (N_2064,In_567,In_2494);
nor U2065 (N_2065,In_485,In_718);
or U2066 (N_2066,In_1495,In_947);
nor U2067 (N_2067,In_1168,In_1029);
or U2068 (N_2068,In_1927,In_91);
nand U2069 (N_2069,In_1899,In_1496);
and U2070 (N_2070,In_1834,In_1604);
and U2071 (N_2071,In_1812,In_2014);
and U2072 (N_2072,In_2359,In_1718);
nor U2073 (N_2073,In_1727,In_1059);
nand U2074 (N_2074,In_332,In_1750);
and U2075 (N_2075,In_2487,In_811);
and U2076 (N_2076,In_985,In_1131);
xor U2077 (N_2077,In_2048,In_2275);
and U2078 (N_2078,In_11,In_2240);
nor U2079 (N_2079,In_336,In_777);
nand U2080 (N_2080,In_147,In_1618);
or U2081 (N_2081,In_691,In_2171);
and U2082 (N_2082,In_1437,In_2285);
nor U2083 (N_2083,In_473,In_485);
and U2084 (N_2084,In_1998,In_1105);
xnor U2085 (N_2085,In_426,In_30);
xor U2086 (N_2086,In_978,In_1670);
xnor U2087 (N_2087,In_949,In_541);
xor U2088 (N_2088,In_554,In_1007);
xor U2089 (N_2089,In_2389,In_396);
nor U2090 (N_2090,In_2232,In_222);
xor U2091 (N_2091,In_404,In_938);
and U2092 (N_2092,In_387,In_1138);
nand U2093 (N_2093,In_1738,In_2300);
xnor U2094 (N_2094,In_1623,In_571);
and U2095 (N_2095,In_2093,In_394);
nand U2096 (N_2096,In_1920,In_1533);
nand U2097 (N_2097,In_130,In_2299);
or U2098 (N_2098,In_1932,In_2433);
nand U2099 (N_2099,In_2497,In_999);
or U2100 (N_2100,In_1068,In_1754);
nand U2101 (N_2101,In_1335,In_931);
and U2102 (N_2102,In_1886,In_1095);
nand U2103 (N_2103,In_1670,In_1178);
and U2104 (N_2104,In_4,In_924);
or U2105 (N_2105,In_1151,In_1726);
nand U2106 (N_2106,In_1382,In_1861);
nand U2107 (N_2107,In_1093,In_322);
or U2108 (N_2108,In_2081,In_237);
and U2109 (N_2109,In_175,In_338);
nor U2110 (N_2110,In_1962,In_1043);
nand U2111 (N_2111,In_2001,In_1843);
xor U2112 (N_2112,In_1485,In_485);
nand U2113 (N_2113,In_524,In_2162);
xor U2114 (N_2114,In_1694,In_161);
or U2115 (N_2115,In_1069,In_198);
and U2116 (N_2116,In_689,In_793);
or U2117 (N_2117,In_2209,In_1410);
nand U2118 (N_2118,In_2167,In_935);
nor U2119 (N_2119,In_1942,In_1665);
and U2120 (N_2120,In_2143,In_611);
nand U2121 (N_2121,In_1530,In_2140);
and U2122 (N_2122,In_2000,In_1663);
or U2123 (N_2123,In_109,In_1866);
nor U2124 (N_2124,In_1777,In_663);
xor U2125 (N_2125,In_1460,In_566);
nand U2126 (N_2126,In_835,In_717);
nor U2127 (N_2127,In_85,In_652);
nor U2128 (N_2128,In_705,In_2044);
and U2129 (N_2129,In_2390,In_1955);
or U2130 (N_2130,In_2438,In_1137);
nand U2131 (N_2131,In_849,In_1054);
or U2132 (N_2132,In_1461,In_1575);
nand U2133 (N_2133,In_2341,In_220);
nor U2134 (N_2134,In_1028,In_176);
and U2135 (N_2135,In_366,In_2045);
nand U2136 (N_2136,In_1740,In_607);
and U2137 (N_2137,In_1213,In_1931);
nand U2138 (N_2138,In_1334,In_688);
nand U2139 (N_2139,In_2251,In_2147);
xnor U2140 (N_2140,In_1040,In_2081);
xnor U2141 (N_2141,In_1586,In_2190);
xnor U2142 (N_2142,In_2246,In_2122);
nor U2143 (N_2143,In_1799,In_676);
or U2144 (N_2144,In_1987,In_736);
xor U2145 (N_2145,In_2387,In_1551);
nor U2146 (N_2146,In_1142,In_2231);
xor U2147 (N_2147,In_949,In_1920);
xnor U2148 (N_2148,In_1761,In_1428);
xor U2149 (N_2149,In_1208,In_2003);
xnor U2150 (N_2150,In_1262,In_236);
nor U2151 (N_2151,In_1279,In_1552);
xor U2152 (N_2152,In_2026,In_162);
xnor U2153 (N_2153,In_2378,In_920);
nor U2154 (N_2154,In_1319,In_1487);
nor U2155 (N_2155,In_175,In_1493);
or U2156 (N_2156,In_1605,In_1088);
and U2157 (N_2157,In_1105,In_1062);
nand U2158 (N_2158,In_624,In_120);
or U2159 (N_2159,In_2146,In_2002);
and U2160 (N_2160,In_1101,In_2061);
and U2161 (N_2161,In_1170,In_142);
or U2162 (N_2162,In_1142,In_1666);
xor U2163 (N_2163,In_831,In_803);
or U2164 (N_2164,In_1787,In_245);
and U2165 (N_2165,In_2450,In_2287);
nor U2166 (N_2166,In_834,In_1745);
xor U2167 (N_2167,In_1225,In_1936);
or U2168 (N_2168,In_580,In_1124);
xor U2169 (N_2169,In_844,In_1499);
xor U2170 (N_2170,In_352,In_217);
nand U2171 (N_2171,In_1247,In_1325);
xor U2172 (N_2172,In_1787,In_2121);
or U2173 (N_2173,In_1222,In_164);
or U2174 (N_2174,In_1502,In_1196);
or U2175 (N_2175,In_1283,In_510);
xor U2176 (N_2176,In_154,In_353);
nor U2177 (N_2177,In_1883,In_137);
or U2178 (N_2178,In_1954,In_141);
nor U2179 (N_2179,In_1626,In_572);
and U2180 (N_2180,In_1953,In_76);
nand U2181 (N_2181,In_427,In_355);
xor U2182 (N_2182,In_624,In_85);
and U2183 (N_2183,In_470,In_40);
or U2184 (N_2184,In_1819,In_90);
xor U2185 (N_2185,In_1461,In_576);
and U2186 (N_2186,In_1900,In_636);
nand U2187 (N_2187,In_1269,In_1617);
nand U2188 (N_2188,In_125,In_473);
nand U2189 (N_2189,In_1635,In_2467);
xnor U2190 (N_2190,In_1250,In_2229);
and U2191 (N_2191,In_1455,In_2119);
and U2192 (N_2192,In_1168,In_1670);
xnor U2193 (N_2193,In_471,In_1247);
xnor U2194 (N_2194,In_1737,In_1318);
nor U2195 (N_2195,In_1608,In_1478);
or U2196 (N_2196,In_656,In_1268);
and U2197 (N_2197,In_1591,In_2182);
and U2198 (N_2198,In_1714,In_353);
xnor U2199 (N_2199,In_2453,In_619);
nand U2200 (N_2200,In_473,In_202);
and U2201 (N_2201,In_461,In_648);
nor U2202 (N_2202,In_1811,In_1853);
and U2203 (N_2203,In_1040,In_909);
and U2204 (N_2204,In_517,In_968);
xor U2205 (N_2205,In_2212,In_1470);
and U2206 (N_2206,In_861,In_1920);
xnor U2207 (N_2207,In_621,In_781);
nand U2208 (N_2208,In_2132,In_207);
nand U2209 (N_2209,In_100,In_615);
nor U2210 (N_2210,In_1407,In_1023);
and U2211 (N_2211,In_1787,In_69);
nor U2212 (N_2212,In_796,In_1556);
and U2213 (N_2213,In_1583,In_1184);
nor U2214 (N_2214,In_657,In_2210);
nor U2215 (N_2215,In_2395,In_2283);
nand U2216 (N_2216,In_1620,In_705);
nand U2217 (N_2217,In_2024,In_988);
nor U2218 (N_2218,In_341,In_303);
xor U2219 (N_2219,In_481,In_432);
and U2220 (N_2220,In_638,In_1482);
nand U2221 (N_2221,In_2414,In_1388);
xnor U2222 (N_2222,In_1035,In_985);
nand U2223 (N_2223,In_2199,In_2002);
nand U2224 (N_2224,In_1206,In_355);
nor U2225 (N_2225,In_4,In_1360);
nand U2226 (N_2226,In_1785,In_1227);
xor U2227 (N_2227,In_1580,In_67);
nand U2228 (N_2228,In_2023,In_2476);
and U2229 (N_2229,In_263,In_1319);
nand U2230 (N_2230,In_1930,In_973);
xor U2231 (N_2231,In_2415,In_2298);
or U2232 (N_2232,In_2152,In_1960);
and U2233 (N_2233,In_1406,In_298);
or U2234 (N_2234,In_241,In_26);
nand U2235 (N_2235,In_885,In_1548);
and U2236 (N_2236,In_2065,In_621);
or U2237 (N_2237,In_706,In_693);
nor U2238 (N_2238,In_210,In_100);
or U2239 (N_2239,In_825,In_768);
and U2240 (N_2240,In_2000,In_1035);
nand U2241 (N_2241,In_908,In_753);
nand U2242 (N_2242,In_1625,In_2096);
nor U2243 (N_2243,In_2289,In_1576);
or U2244 (N_2244,In_195,In_91);
or U2245 (N_2245,In_1348,In_1560);
or U2246 (N_2246,In_760,In_1596);
xnor U2247 (N_2247,In_1741,In_2215);
xnor U2248 (N_2248,In_1017,In_912);
and U2249 (N_2249,In_1614,In_1383);
and U2250 (N_2250,In_1211,In_771);
and U2251 (N_2251,In_1710,In_1388);
xor U2252 (N_2252,In_522,In_805);
and U2253 (N_2253,In_2046,In_1636);
xor U2254 (N_2254,In_498,In_288);
nor U2255 (N_2255,In_400,In_421);
and U2256 (N_2256,In_918,In_1818);
or U2257 (N_2257,In_13,In_1864);
nand U2258 (N_2258,In_523,In_122);
and U2259 (N_2259,In_1635,In_1979);
and U2260 (N_2260,In_1768,In_548);
and U2261 (N_2261,In_2199,In_395);
nor U2262 (N_2262,In_1134,In_1915);
nand U2263 (N_2263,In_1264,In_496);
and U2264 (N_2264,In_464,In_527);
and U2265 (N_2265,In_2358,In_479);
xor U2266 (N_2266,In_938,In_1877);
or U2267 (N_2267,In_1211,In_1133);
xor U2268 (N_2268,In_749,In_764);
and U2269 (N_2269,In_1326,In_1574);
nor U2270 (N_2270,In_1165,In_626);
and U2271 (N_2271,In_1102,In_1819);
or U2272 (N_2272,In_63,In_2473);
nor U2273 (N_2273,In_540,In_1767);
and U2274 (N_2274,In_1895,In_1250);
xnor U2275 (N_2275,In_1591,In_753);
nor U2276 (N_2276,In_832,In_456);
nand U2277 (N_2277,In_73,In_1495);
nand U2278 (N_2278,In_1775,In_498);
nor U2279 (N_2279,In_675,In_797);
xnor U2280 (N_2280,In_1921,In_1375);
nand U2281 (N_2281,In_1814,In_849);
nor U2282 (N_2282,In_632,In_609);
or U2283 (N_2283,In_1662,In_349);
xor U2284 (N_2284,In_411,In_585);
nor U2285 (N_2285,In_798,In_6);
or U2286 (N_2286,In_851,In_1831);
or U2287 (N_2287,In_2306,In_2362);
or U2288 (N_2288,In_1215,In_261);
nand U2289 (N_2289,In_1316,In_367);
or U2290 (N_2290,In_2094,In_2048);
or U2291 (N_2291,In_1703,In_457);
xnor U2292 (N_2292,In_1867,In_2390);
xnor U2293 (N_2293,In_2295,In_1831);
xnor U2294 (N_2294,In_843,In_1181);
xor U2295 (N_2295,In_1339,In_1568);
nand U2296 (N_2296,In_1586,In_307);
nand U2297 (N_2297,In_1351,In_484);
and U2298 (N_2298,In_1797,In_1280);
nand U2299 (N_2299,In_1427,In_2319);
or U2300 (N_2300,In_1657,In_700);
and U2301 (N_2301,In_1664,In_351);
xor U2302 (N_2302,In_551,In_1927);
xnor U2303 (N_2303,In_299,In_1366);
and U2304 (N_2304,In_1108,In_848);
xor U2305 (N_2305,In_1583,In_1496);
nor U2306 (N_2306,In_1722,In_123);
or U2307 (N_2307,In_2350,In_1698);
or U2308 (N_2308,In_236,In_681);
xnor U2309 (N_2309,In_230,In_841);
nor U2310 (N_2310,In_1973,In_1185);
nand U2311 (N_2311,In_1589,In_150);
or U2312 (N_2312,In_949,In_273);
xor U2313 (N_2313,In_780,In_2099);
and U2314 (N_2314,In_2126,In_2464);
or U2315 (N_2315,In_1222,In_427);
and U2316 (N_2316,In_2014,In_348);
xnor U2317 (N_2317,In_782,In_1993);
nand U2318 (N_2318,In_1443,In_1738);
nand U2319 (N_2319,In_2069,In_577);
xor U2320 (N_2320,In_1931,In_1028);
nand U2321 (N_2321,In_2085,In_543);
nor U2322 (N_2322,In_2473,In_1073);
nor U2323 (N_2323,In_812,In_1307);
or U2324 (N_2324,In_793,In_634);
xnor U2325 (N_2325,In_972,In_2479);
or U2326 (N_2326,In_281,In_1600);
nand U2327 (N_2327,In_354,In_2022);
xor U2328 (N_2328,In_14,In_1880);
xor U2329 (N_2329,In_811,In_255);
xor U2330 (N_2330,In_1626,In_2487);
nand U2331 (N_2331,In_2175,In_1747);
or U2332 (N_2332,In_71,In_1938);
xor U2333 (N_2333,In_2497,In_1342);
nor U2334 (N_2334,In_1040,In_239);
nand U2335 (N_2335,In_1575,In_712);
and U2336 (N_2336,In_2373,In_2170);
nor U2337 (N_2337,In_1732,In_1923);
xnor U2338 (N_2338,In_1492,In_1475);
xor U2339 (N_2339,In_259,In_359);
or U2340 (N_2340,In_1960,In_861);
or U2341 (N_2341,In_932,In_402);
or U2342 (N_2342,In_164,In_1887);
and U2343 (N_2343,In_430,In_130);
nor U2344 (N_2344,In_1930,In_306);
xnor U2345 (N_2345,In_2455,In_653);
or U2346 (N_2346,In_935,In_2405);
xnor U2347 (N_2347,In_1724,In_325);
nand U2348 (N_2348,In_1913,In_2390);
or U2349 (N_2349,In_1103,In_950);
nor U2350 (N_2350,In_2144,In_900);
xor U2351 (N_2351,In_1422,In_338);
xor U2352 (N_2352,In_292,In_559);
nand U2353 (N_2353,In_536,In_2404);
nand U2354 (N_2354,In_774,In_2187);
nor U2355 (N_2355,In_291,In_2180);
xnor U2356 (N_2356,In_984,In_2021);
and U2357 (N_2357,In_1764,In_1163);
or U2358 (N_2358,In_815,In_1426);
nor U2359 (N_2359,In_1338,In_467);
nand U2360 (N_2360,In_1739,In_708);
and U2361 (N_2361,In_1300,In_1137);
nand U2362 (N_2362,In_115,In_492);
and U2363 (N_2363,In_1498,In_503);
xnor U2364 (N_2364,In_344,In_1645);
or U2365 (N_2365,In_1768,In_231);
or U2366 (N_2366,In_1555,In_1641);
xnor U2367 (N_2367,In_1103,In_130);
or U2368 (N_2368,In_479,In_1798);
nand U2369 (N_2369,In_1832,In_1805);
or U2370 (N_2370,In_2307,In_2384);
or U2371 (N_2371,In_1716,In_433);
and U2372 (N_2372,In_2312,In_162);
nor U2373 (N_2373,In_1368,In_1173);
nand U2374 (N_2374,In_2197,In_1217);
nand U2375 (N_2375,In_1043,In_1456);
or U2376 (N_2376,In_974,In_2411);
and U2377 (N_2377,In_327,In_2409);
and U2378 (N_2378,In_2393,In_1301);
and U2379 (N_2379,In_840,In_42);
nand U2380 (N_2380,In_34,In_2188);
and U2381 (N_2381,In_746,In_1254);
nor U2382 (N_2382,In_2444,In_967);
or U2383 (N_2383,In_1904,In_1545);
xor U2384 (N_2384,In_1762,In_2340);
and U2385 (N_2385,In_2026,In_2496);
nor U2386 (N_2386,In_1584,In_73);
nand U2387 (N_2387,In_1175,In_1727);
nand U2388 (N_2388,In_440,In_322);
nor U2389 (N_2389,In_1040,In_735);
and U2390 (N_2390,In_1256,In_2172);
xnor U2391 (N_2391,In_780,In_1036);
and U2392 (N_2392,In_152,In_185);
or U2393 (N_2393,In_755,In_1014);
or U2394 (N_2394,In_2035,In_528);
and U2395 (N_2395,In_12,In_1514);
nor U2396 (N_2396,In_1969,In_43);
xnor U2397 (N_2397,In_722,In_1669);
or U2398 (N_2398,In_1855,In_504);
nor U2399 (N_2399,In_1707,In_406);
and U2400 (N_2400,In_1807,In_1490);
nor U2401 (N_2401,In_2396,In_366);
nand U2402 (N_2402,In_1100,In_71);
xor U2403 (N_2403,In_1133,In_57);
and U2404 (N_2404,In_1148,In_468);
xnor U2405 (N_2405,In_2497,In_939);
xnor U2406 (N_2406,In_473,In_1242);
nor U2407 (N_2407,In_313,In_575);
xnor U2408 (N_2408,In_309,In_1420);
and U2409 (N_2409,In_1051,In_1998);
nor U2410 (N_2410,In_1996,In_953);
nand U2411 (N_2411,In_284,In_2317);
nand U2412 (N_2412,In_1508,In_816);
xor U2413 (N_2413,In_2172,In_1752);
and U2414 (N_2414,In_511,In_1922);
or U2415 (N_2415,In_54,In_340);
xor U2416 (N_2416,In_1144,In_2122);
or U2417 (N_2417,In_1674,In_130);
or U2418 (N_2418,In_1862,In_2428);
nand U2419 (N_2419,In_1127,In_1539);
xnor U2420 (N_2420,In_128,In_1745);
and U2421 (N_2421,In_2370,In_135);
nor U2422 (N_2422,In_2328,In_1137);
or U2423 (N_2423,In_618,In_677);
xnor U2424 (N_2424,In_1905,In_1629);
and U2425 (N_2425,In_441,In_1027);
nand U2426 (N_2426,In_1532,In_303);
nor U2427 (N_2427,In_1362,In_165);
xnor U2428 (N_2428,In_899,In_1047);
nor U2429 (N_2429,In_1794,In_2039);
nand U2430 (N_2430,In_1243,In_160);
or U2431 (N_2431,In_1518,In_836);
xnor U2432 (N_2432,In_403,In_2371);
nor U2433 (N_2433,In_1764,In_2211);
or U2434 (N_2434,In_1726,In_1317);
nor U2435 (N_2435,In_540,In_2486);
nor U2436 (N_2436,In_980,In_941);
and U2437 (N_2437,In_2220,In_739);
and U2438 (N_2438,In_902,In_1227);
xor U2439 (N_2439,In_831,In_1241);
and U2440 (N_2440,In_1258,In_1202);
or U2441 (N_2441,In_707,In_1542);
nor U2442 (N_2442,In_92,In_1803);
or U2443 (N_2443,In_398,In_1976);
and U2444 (N_2444,In_2023,In_294);
nor U2445 (N_2445,In_1167,In_1843);
nand U2446 (N_2446,In_1141,In_968);
or U2447 (N_2447,In_1314,In_739);
and U2448 (N_2448,In_1791,In_2417);
and U2449 (N_2449,In_2378,In_761);
nor U2450 (N_2450,In_361,In_945);
nor U2451 (N_2451,In_322,In_1185);
nor U2452 (N_2452,In_2007,In_2189);
or U2453 (N_2453,In_2306,In_2247);
xnor U2454 (N_2454,In_1344,In_2005);
nor U2455 (N_2455,In_565,In_1614);
or U2456 (N_2456,In_1772,In_1619);
and U2457 (N_2457,In_335,In_726);
or U2458 (N_2458,In_1785,In_1976);
nor U2459 (N_2459,In_1395,In_554);
xnor U2460 (N_2460,In_1779,In_19);
xor U2461 (N_2461,In_23,In_1214);
or U2462 (N_2462,In_1384,In_1164);
nand U2463 (N_2463,In_2414,In_117);
xnor U2464 (N_2464,In_460,In_1817);
xor U2465 (N_2465,In_126,In_1189);
nor U2466 (N_2466,In_2037,In_2483);
nor U2467 (N_2467,In_141,In_435);
or U2468 (N_2468,In_2477,In_1414);
nor U2469 (N_2469,In_411,In_2220);
nand U2470 (N_2470,In_2388,In_14);
or U2471 (N_2471,In_345,In_295);
xor U2472 (N_2472,In_1143,In_2063);
and U2473 (N_2473,In_2061,In_1293);
nand U2474 (N_2474,In_281,In_1594);
nand U2475 (N_2475,In_1680,In_1125);
or U2476 (N_2476,In_1368,In_477);
or U2477 (N_2477,In_550,In_2410);
nor U2478 (N_2478,In_1400,In_380);
xnor U2479 (N_2479,In_146,In_51);
and U2480 (N_2480,In_779,In_314);
nand U2481 (N_2481,In_989,In_1586);
and U2482 (N_2482,In_2037,In_2274);
nand U2483 (N_2483,In_2192,In_1925);
and U2484 (N_2484,In_2048,In_784);
xor U2485 (N_2485,In_1226,In_1693);
nor U2486 (N_2486,In_369,In_416);
xor U2487 (N_2487,In_1088,In_2069);
xor U2488 (N_2488,In_618,In_2179);
and U2489 (N_2489,In_2008,In_1212);
nand U2490 (N_2490,In_1533,In_2308);
or U2491 (N_2491,In_2451,In_494);
or U2492 (N_2492,In_678,In_165);
nand U2493 (N_2493,In_801,In_1933);
xor U2494 (N_2494,In_2121,In_1396);
and U2495 (N_2495,In_1117,In_1445);
nand U2496 (N_2496,In_1727,In_2209);
nor U2497 (N_2497,In_641,In_823);
or U2498 (N_2498,In_1181,In_245);
or U2499 (N_2499,In_2386,In_946);
or U2500 (N_2500,In_1553,In_1156);
nor U2501 (N_2501,In_1677,In_2434);
or U2502 (N_2502,In_1415,In_1827);
nor U2503 (N_2503,In_767,In_1433);
and U2504 (N_2504,In_1943,In_794);
nand U2505 (N_2505,In_10,In_1084);
xnor U2506 (N_2506,In_1147,In_1498);
nand U2507 (N_2507,In_1087,In_122);
nor U2508 (N_2508,In_1953,In_248);
nand U2509 (N_2509,In_730,In_1174);
or U2510 (N_2510,In_1164,In_1078);
nand U2511 (N_2511,In_2259,In_1977);
and U2512 (N_2512,In_1831,In_487);
and U2513 (N_2513,In_129,In_2373);
nor U2514 (N_2514,In_1805,In_1494);
nor U2515 (N_2515,In_1927,In_1150);
nand U2516 (N_2516,In_654,In_2299);
xnor U2517 (N_2517,In_716,In_876);
xnor U2518 (N_2518,In_1680,In_1780);
or U2519 (N_2519,In_199,In_1339);
nand U2520 (N_2520,In_2275,In_615);
or U2521 (N_2521,In_2363,In_2029);
nor U2522 (N_2522,In_2434,In_1811);
xor U2523 (N_2523,In_1680,In_1574);
nor U2524 (N_2524,In_1805,In_1243);
nand U2525 (N_2525,In_1895,In_226);
or U2526 (N_2526,In_1567,In_2198);
and U2527 (N_2527,In_1416,In_2025);
nor U2528 (N_2528,In_685,In_126);
xor U2529 (N_2529,In_175,In_2066);
xnor U2530 (N_2530,In_2169,In_923);
and U2531 (N_2531,In_386,In_2165);
nand U2532 (N_2532,In_809,In_1526);
xnor U2533 (N_2533,In_1688,In_1168);
xnor U2534 (N_2534,In_2426,In_871);
nand U2535 (N_2535,In_767,In_781);
or U2536 (N_2536,In_1745,In_1190);
and U2537 (N_2537,In_2252,In_896);
nand U2538 (N_2538,In_4,In_1645);
or U2539 (N_2539,In_37,In_791);
or U2540 (N_2540,In_103,In_761);
or U2541 (N_2541,In_2276,In_1527);
nor U2542 (N_2542,In_700,In_2197);
xor U2543 (N_2543,In_1249,In_450);
and U2544 (N_2544,In_886,In_737);
xnor U2545 (N_2545,In_2374,In_621);
xor U2546 (N_2546,In_385,In_635);
nand U2547 (N_2547,In_2103,In_2098);
and U2548 (N_2548,In_2049,In_1634);
and U2549 (N_2549,In_1022,In_1498);
nor U2550 (N_2550,In_166,In_164);
or U2551 (N_2551,In_242,In_1285);
nand U2552 (N_2552,In_932,In_1944);
xnor U2553 (N_2553,In_146,In_1617);
xor U2554 (N_2554,In_1677,In_1443);
nor U2555 (N_2555,In_1281,In_538);
xnor U2556 (N_2556,In_1555,In_588);
nand U2557 (N_2557,In_404,In_2221);
nand U2558 (N_2558,In_1529,In_2474);
nand U2559 (N_2559,In_740,In_2032);
nor U2560 (N_2560,In_1338,In_16);
nor U2561 (N_2561,In_2164,In_1685);
and U2562 (N_2562,In_1849,In_1226);
and U2563 (N_2563,In_1652,In_1637);
nand U2564 (N_2564,In_1239,In_1372);
nor U2565 (N_2565,In_1460,In_1164);
and U2566 (N_2566,In_92,In_773);
and U2567 (N_2567,In_2418,In_1644);
nand U2568 (N_2568,In_32,In_904);
xor U2569 (N_2569,In_510,In_839);
nor U2570 (N_2570,In_2448,In_2359);
nand U2571 (N_2571,In_2360,In_1959);
or U2572 (N_2572,In_161,In_1296);
nand U2573 (N_2573,In_1224,In_1262);
nand U2574 (N_2574,In_747,In_189);
nand U2575 (N_2575,In_2238,In_424);
and U2576 (N_2576,In_180,In_614);
or U2577 (N_2577,In_2374,In_1513);
and U2578 (N_2578,In_62,In_1374);
xnor U2579 (N_2579,In_2182,In_1897);
or U2580 (N_2580,In_1733,In_1654);
or U2581 (N_2581,In_1741,In_658);
or U2582 (N_2582,In_1337,In_597);
and U2583 (N_2583,In_2141,In_1945);
nor U2584 (N_2584,In_2476,In_940);
or U2585 (N_2585,In_416,In_1207);
nand U2586 (N_2586,In_2453,In_2135);
nor U2587 (N_2587,In_1972,In_2454);
or U2588 (N_2588,In_547,In_1740);
xnor U2589 (N_2589,In_1584,In_2144);
and U2590 (N_2590,In_699,In_214);
nor U2591 (N_2591,In_734,In_1679);
nand U2592 (N_2592,In_1693,In_1649);
xnor U2593 (N_2593,In_993,In_88);
nand U2594 (N_2594,In_532,In_1891);
nor U2595 (N_2595,In_2112,In_7);
nor U2596 (N_2596,In_1127,In_1630);
or U2597 (N_2597,In_1215,In_2418);
nor U2598 (N_2598,In_2041,In_1817);
or U2599 (N_2599,In_1894,In_1938);
nor U2600 (N_2600,In_2145,In_2080);
and U2601 (N_2601,In_765,In_522);
xnor U2602 (N_2602,In_1403,In_33);
and U2603 (N_2603,In_0,In_782);
nand U2604 (N_2604,In_1668,In_1402);
xnor U2605 (N_2605,In_288,In_2040);
nand U2606 (N_2606,In_1653,In_2268);
nand U2607 (N_2607,In_625,In_1772);
xnor U2608 (N_2608,In_2294,In_1366);
nand U2609 (N_2609,In_71,In_1230);
or U2610 (N_2610,In_1359,In_453);
and U2611 (N_2611,In_1528,In_883);
nand U2612 (N_2612,In_2222,In_1962);
or U2613 (N_2613,In_960,In_2254);
and U2614 (N_2614,In_1294,In_1847);
nand U2615 (N_2615,In_661,In_2366);
or U2616 (N_2616,In_1141,In_1527);
nor U2617 (N_2617,In_1231,In_1232);
nand U2618 (N_2618,In_1047,In_1071);
nor U2619 (N_2619,In_2376,In_1345);
and U2620 (N_2620,In_1177,In_499);
nor U2621 (N_2621,In_2308,In_378);
or U2622 (N_2622,In_2495,In_1470);
nor U2623 (N_2623,In_1061,In_1671);
nor U2624 (N_2624,In_931,In_1528);
and U2625 (N_2625,In_406,In_941);
nor U2626 (N_2626,In_2195,In_2468);
and U2627 (N_2627,In_1358,In_554);
xor U2628 (N_2628,In_1327,In_2190);
and U2629 (N_2629,In_746,In_355);
nand U2630 (N_2630,In_300,In_342);
or U2631 (N_2631,In_2199,In_536);
nand U2632 (N_2632,In_883,In_1982);
xor U2633 (N_2633,In_713,In_1059);
nand U2634 (N_2634,In_1843,In_1607);
nor U2635 (N_2635,In_825,In_184);
xor U2636 (N_2636,In_2061,In_34);
nor U2637 (N_2637,In_274,In_1149);
nand U2638 (N_2638,In_529,In_1980);
nor U2639 (N_2639,In_32,In_1527);
nor U2640 (N_2640,In_2272,In_262);
nand U2641 (N_2641,In_268,In_1637);
and U2642 (N_2642,In_5,In_1165);
and U2643 (N_2643,In_1380,In_1726);
or U2644 (N_2644,In_1508,In_2347);
nor U2645 (N_2645,In_1857,In_1193);
nand U2646 (N_2646,In_1505,In_2196);
and U2647 (N_2647,In_2464,In_641);
nor U2648 (N_2648,In_1799,In_1930);
xnor U2649 (N_2649,In_2294,In_189);
and U2650 (N_2650,In_936,In_207);
and U2651 (N_2651,In_819,In_438);
or U2652 (N_2652,In_1353,In_1228);
nor U2653 (N_2653,In_2391,In_744);
nand U2654 (N_2654,In_1437,In_858);
xnor U2655 (N_2655,In_2006,In_2150);
nand U2656 (N_2656,In_1870,In_741);
or U2657 (N_2657,In_1098,In_686);
nor U2658 (N_2658,In_2465,In_1969);
nand U2659 (N_2659,In_2138,In_2380);
and U2660 (N_2660,In_1052,In_516);
nand U2661 (N_2661,In_851,In_101);
xnor U2662 (N_2662,In_1455,In_71);
or U2663 (N_2663,In_1770,In_2148);
and U2664 (N_2664,In_1161,In_1166);
nand U2665 (N_2665,In_1604,In_181);
and U2666 (N_2666,In_166,In_470);
xnor U2667 (N_2667,In_252,In_2344);
or U2668 (N_2668,In_401,In_971);
or U2669 (N_2669,In_2413,In_2324);
or U2670 (N_2670,In_515,In_2444);
nand U2671 (N_2671,In_1146,In_1055);
nor U2672 (N_2672,In_193,In_1675);
nor U2673 (N_2673,In_816,In_1313);
and U2674 (N_2674,In_1714,In_1662);
xor U2675 (N_2675,In_2351,In_224);
nand U2676 (N_2676,In_2010,In_1711);
nand U2677 (N_2677,In_14,In_1670);
nor U2678 (N_2678,In_1311,In_2282);
nand U2679 (N_2679,In_652,In_1832);
xor U2680 (N_2680,In_1411,In_457);
and U2681 (N_2681,In_1040,In_1190);
xnor U2682 (N_2682,In_1875,In_854);
nor U2683 (N_2683,In_1082,In_1733);
and U2684 (N_2684,In_117,In_2032);
nand U2685 (N_2685,In_564,In_2234);
or U2686 (N_2686,In_1283,In_348);
nor U2687 (N_2687,In_599,In_2167);
or U2688 (N_2688,In_1101,In_2362);
or U2689 (N_2689,In_581,In_437);
xor U2690 (N_2690,In_701,In_713);
xor U2691 (N_2691,In_265,In_273);
or U2692 (N_2692,In_2063,In_80);
and U2693 (N_2693,In_2404,In_1948);
and U2694 (N_2694,In_2252,In_1022);
and U2695 (N_2695,In_1236,In_2042);
or U2696 (N_2696,In_2379,In_1151);
and U2697 (N_2697,In_1013,In_578);
nor U2698 (N_2698,In_2145,In_610);
nor U2699 (N_2699,In_129,In_1455);
and U2700 (N_2700,In_1894,In_96);
and U2701 (N_2701,In_180,In_1875);
xnor U2702 (N_2702,In_1918,In_1563);
xnor U2703 (N_2703,In_1562,In_193);
and U2704 (N_2704,In_1457,In_238);
xor U2705 (N_2705,In_488,In_1411);
or U2706 (N_2706,In_1659,In_2247);
xnor U2707 (N_2707,In_1556,In_991);
nor U2708 (N_2708,In_1813,In_1431);
or U2709 (N_2709,In_1746,In_2391);
nand U2710 (N_2710,In_2328,In_2122);
nand U2711 (N_2711,In_1441,In_1170);
xor U2712 (N_2712,In_279,In_1313);
nor U2713 (N_2713,In_1833,In_1249);
and U2714 (N_2714,In_2312,In_1933);
nor U2715 (N_2715,In_1799,In_228);
nand U2716 (N_2716,In_2279,In_2370);
or U2717 (N_2717,In_1609,In_1299);
xnor U2718 (N_2718,In_1272,In_2019);
nor U2719 (N_2719,In_1434,In_1777);
xnor U2720 (N_2720,In_1223,In_1047);
and U2721 (N_2721,In_831,In_1432);
or U2722 (N_2722,In_2351,In_289);
and U2723 (N_2723,In_2355,In_199);
nor U2724 (N_2724,In_437,In_1692);
or U2725 (N_2725,In_81,In_411);
xor U2726 (N_2726,In_99,In_2256);
nand U2727 (N_2727,In_2261,In_1761);
or U2728 (N_2728,In_216,In_2202);
or U2729 (N_2729,In_1197,In_1740);
xor U2730 (N_2730,In_297,In_1375);
xor U2731 (N_2731,In_83,In_958);
nor U2732 (N_2732,In_1900,In_1395);
or U2733 (N_2733,In_332,In_2264);
xor U2734 (N_2734,In_456,In_1703);
and U2735 (N_2735,In_377,In_1426);
nand U2736 (N_2736,In_1322,In_995);
nor U2737 (N_2737,In_1157,In_2419);
and U2738 (N_2738,In_2085,In_1563);
or U2739 (N_2739,In_529,In_2462);
nor U2740 (N_2740,In_1849,In_1135);
nand U2741 (N_2741,In_256,In_1161);
nor U2742 (N_2742,In_408,In_443);
xor U2743 (N_2743,In_1209,In_2153);
or U2744 (N_2744,In_596,In_2025);
nand U2745 (N_2745,In_1646,In_537);
or U2746 (N_2746,In_1329,In_2290);
and U2747 (N_2747,In_30,In_1540);
nor U2748 (N_2748,In_1907,In_176);
xnor U2749 (N_2749,In_1989,In_644);
xnor U2750 (N_2750,In_2450,In_57);
or U2751 (N_2751,In_2372,In_992);
nor U2752 (N_2752,In_648,In_1666);
nor U2753 (N_2753,In_1846,In_2479);
xor U2754 (N_2754,In_2105,In_864);
nand U2755 (N_2755,In_1504,In_2233);
or U2756 (N_2756,In_571,In_1830);
and U2757 (N_2757,In_832,In_1813);
xnor U2758 (N_2758,In_2211,In_1244);
or U2759 (N_2759,In_544,In_273);
nand U2760 (N_2760,In_889,In_142);
xor U2761 (N_2761,In_1890,In_1926);
xor U2762 (N_2762,In_400,In_1819);
nor U2763 (N_2763,In_2180,In_1840);
xnor U2764 (N_2764,In_670,In_1404);
or U2765 (N_2765,In_511,In_866);
nand U2766 (N_2766,In_310,In_356);
nor U2767 (N_2767,In_1638,In_39);
nand U2768 (N_2768,In_56,In_1438);
xnor U2769 (N_2769,In_2493,In_1695);
nand U2770 (N_2770,In_1953,In_392);
and U2771 (N_2771,In_972,In_188);
nor U2772 (N_2772,In_2330,In_1513);
xnor U2773 (N_2773,In_2208,In_1906);
nand U2774 (N_2774,In_680,In_512);
and U2775 (N_2775,In_129,In_36);
and U2776 (N_2776,In_1758,In_1658);
xnor U2777 (N_2777,In_1665,In_95);
and U2778 (N_2778,In_321,In_1562);
and U2779 (N_2779,In_1888,In_1510);
or U2780 (N_2780,In_200,In_312);
or U2781 (N_2781,In_1729,In_1870);
and U2782 (N_2782,In_2086,In_1975);
and U2783 (N_2783,In_1058,In_423);
or U2784 (N_2784,In_1762,In_1889);
nor U2785 (N_2785,In_391,In_2154);
and U2786 (N_2786,In_330,In_93);
and U2787 (N_2787,In_611,In_2298);
nand U2788 (N_2788,In_441,In_1991);
nor U2789 (N_2789,In_1615,In_2432);
nor U2790 (N_2790,In_2042,In_2198);
or U2791 (N_2791,In_131,In_1923);
and U2792 (N_2792,In_1024,In_2258);
nand U2793 (N_2793,In_1500,In_1884);
nor U2794 (N_2794,In_2429,In_1340);
and U2795 (N_2795,In_2298,In_2028);
nand U2796 (N_2796,In_2130,In_501);
xnor U2797 (N_2797,In_1035,In_1755);
or U2798 (N_2798,In_1022,In_1499);
and U2799 (N_2799,In_1061,In_465);
and U2800 (N_2800,In_335,In_594);
xor U2801 (N_2801,In_1395,In_1871);
or U2802 (N_2802,In_629,In_1322);
xor U2803 (N_2803,In_1477,In_2153);
xnor U2804 (N_2804,In_1302,In_2370);
nand U2805 (N_2805,In_1079,In_2256);
and U2806 (N_2806,In_2218,In_1151);
xor U2807 (N_2807,In_1541,In_2001);
nand U2808 (N_2808,In_383,In_330);
nor U2809 (N_2809,In_317,In_2218);
or U2810 (N_2810,In_524,In_2249);
and U2811 (N_2811,In_1490,In_911);
nand U2812 (N_2812,In_614,In_160);
nor U2813 (N_2813,In_645,In_450);
or U2814 (N_2814,In_1691,In_1107);
or U2815 (N_2815,In_1561,In_899);
xor U2816 (N_2816,In_385,In_527);
and U2817 (N_2817,In_2426,In_111);
nand U2818 (N_2818,In_1813,In_238);
or U2819 (N_2819,In_2350,In_789);
nor U2820 (N_2820,In_627,In_2034);
or U2821 (N_2821,In_1785,In_1898);
nor U2822 (N_2822,In_19,In_1911);
and U2823 (N_2823,In_1152,In_2123);
and U2824 (N_2824,In_89,In_1413);
and U2825 (N_2825,In_996,In_649);
and U2826 (N_2826,In_207,In_2210);
nor U2827 (N_2827,In_1662,In_1682);
or U2828 (N_2828,In_138,In_1428);
and U2829 (N_2829,In_132,In_677);
or U2830 (N_2830,In_52,In_1523);
or U2831 (N_2831,In_969,In_2136);
nand U2832 (N_2832,In_1316,In_1606);
nor U2833 (N_2833,In_2151,In_1952);
nor U2834 (N_2834,In_828,In_141);
or U2835 (N_2835,In_2109,In_1899);
nor U2836 (N_2836,In_692,In_937);
xor U2837 (N_2837,In_842,In_131);
and U2838 (N_2838,In_1206,In_2415);
and U2839 (N_2839,In_1165,In_896);
nand U2840 (N_2840,In_1252,In_199);
xor U2841 (N_2841,In_1817,In_2095);
and U2842 (N_2842,In_208,In_1829);
nor U2843 (N_2843,In_1987,In_786);
nor U2844 (N_2844,In_158,In_1869);
xnor U2845 (N_2845,In_2138,In_577);
nand U2846 (N_2846,In_1691,In_1748);
or U2847 (N_2847,In_36,In_1527);
or U2848 (N_2848,In_32,In_2123);
or U2849 (N_2849,In_769,In_275);
and U2850 (N_2850,In_1277,In_1194);
nand U2851 (N_2851,In_2195,In_2431);
or U2852 (N_2852,In_1148,In_2459);
nor U2853 (N_2853,In_998,In_559);
xor U2854 (N_2854,In_2321,In_1069);
nor U2855 (N_2855,In_1962,In_302);
nand U2856 (N_2856,In_1271,In_1947);
and U2857 (N_2857,In_1075,In_644);
or U2858 (N_2858,In_1825,In_1902);
or U2859 (N_2859,In_2390,In_1357);
xor U2860 (N_2860,In_599,In_747);
or U2861 (N_2861,In_776,In_2259);
xnor U2862 (N_2862,In_1143,In_284);
or U2863 (N_2863,In_436,In_1480);
nor U2864 (N_2864,In_2463,In_836);
and U2865 (N_2865,In_1377,In_361);
and U2866 (N_2866,In_1952,In_861);
xnor U2867 (N_2867,In_2133,In_1594);
nor U2868 (N_2868,In_573,In_1912);
nand U2869 (N_2869,In_892,In_2379);
xor U2870 (N_2870,In_41,In_1390);
or U2871 (N_2871,In_676,In_1903);
xor U2872 (N_2872,In_1362,In_2396);
xor U2873 (N_2873,In_741,In_977);
xnor U2874 (N_2874,In_1630,In_2310);
xnor U2875 (N_2875,In_1100,In_1393);
nand U2876 (N_2876,In_1392,In_2455);
nor U2877 (N_2877,In_2335,In_325);
xor U2878 (N_2878,In_2129,In_1852);
nor U2879 (N_2879,In_1922,In_2076);
and U2880 (N_2880,In_192,In_963);
nor U2881 (N_2881,In_2364,In_2417);
and U2882 (N_2882,In_956,In_769);
or U2883 (N_2883,In_1247,In_1223);
or U2884 (N_2884,In_2455,In_2051);
nand U2885 (N_2885,In_539,In_1733);
xnor U2886 (N_2886,In_974,In_869);
nor U2887 (N_2887,In_70,In_1915);
and U2888 (N_2888,In_546,In_1424);
nor U2889 (N_2889,In_847,In_316);
nor U2890 (N_2890,In_2377,In_1707);
or U2891 (N_2891,In_2170,In_1740);
xor U2892 (N_2892,In_472,In_2331);
and U2893 (N_2893,In_1172,In_229);
and U2894 (N_2894,In_2368,In_2206);
xor U2895 (N_2895,In_125,In_384);
or U2896 (N_2896,In_1207,In_1882);
or U2897 (N_2897,In_196,In_2222);
or U2898 (N_2898,In_144,In_835);
xor U2899 (N_2899,In_538,In_1546);
nor U2900 (N_2900,In_2379,In_1130);
xor U2901 (N_2901,In_1887,In_1536);
and U2902 (N_2902,In_1058,In_2420);
nand U2903 (N_2903,In_1802,In_361);
nor U2904 (N_2904,In_851,In_1788);
nor U2905 (N_2905,In_157,In_587);
and U2906 (N_2906,In_1934,In_2387);
nor U2907 (N_2907,In_501,In_814);
nor U2908 (N_2908,In_1408,In_2454);
nand U2909 (N_2909,In_340,In_661);
or U2910 (N_2910,In_773,In_180);
nor U2911 (N_2911,In_2434,In_1421);
and U2912 (N_2912,In_340,In_1547);
and U2913 (N_2913,In_934,In_949);
and U2914 (N_2914,In_916,In_1151);
nor U2915 (N_2915,In_1635,In_1203);
xor U2916 (N_2916,In_2380,In_223);
nand U2917 (N_2917,In_2330,In_2414);
or U2918 (N_2918,In_2394,In_1041);
nand U2919 (N_2919,In_1760,In_675);
nand U2920 (N_2920,In_2368,In_743);
nor U2921 (N_2921,In_743,In_917);
or U2922 (N_2922,In_459,In_809);
and U2923 (N_2923,In_1526,In_2025);
xnor U2924 (N_2924,In_48,In_1328);
nand U2925 (N_2925,In_51,In_1363);
or U2926 (N_2926,In_1240,In_1734);
nor U2927 (N_2927,In_690,In_1394);
xnor U2928 (N_2928,In_282,In_1360);
nand U2929 (N_2929,In_1708,In_2449);
nand U2930 (N_2930,In_1355,In_247);
nand U2931 (N_2931,In_1450,In_894);
or U2932 (N_2932,In_533,In_818);
nand U2933 (N_2933,In_1905,In_901);
nand U2934 (N_2934,In_463,In_913);
and U2935 (N_2935,In_2119,In_1542);
or U2936 (N_2936,In_359,In_1631);
or U2937 (N_2937,In_1019,In_299);
nor U2938 (N_2938,In_436,In_66);
and U2939 (N_2939,In_557,In_614);
xnor U2940 (N_2940,In_896,In_2375);
nand U2941 (N_2941,In_2297,In_457);
nand U2942 (N_2942,In_2344,In_1500);
nor U2943 (N_2943,In_1505,In_1180);
and U2944 (N_2944,In_134,In_1389);
or U2945 (N_2945,In_667,In_708);
or U2946 (N_2946,In_2132,In_62);
xnor U2947 (N_2947,In_1241,In_1407);
nor U2948 (N_2948,In_1930,In_1109);
nand U2949 (N_2949,In_1888,In_1318);
and U2950 (N_2950,In_898,In_437);
xor U2951 (N_2951,In_486,In_2355);
xor U2952 (N_2952,In_1182,In_101);
xor U2953 (N_2953,In_1094,In_908);
nand U2954 (N_2954,In_1070,In_678);
xnor U2955 (N_2955,In_2036,In_321);
and U2956 (N_2956,In_1881,In_2258);
and U2957 (N_2957,In_541,In_195);
and U2958 (N_2958,In_1515,In_2283);
xnor U2959 (N_2959,In_412,In_355);
xnor U2960 (N_2960,In_1633,In_1545);
nand U2961 (N_2961,In_1052,In_893);
nand U2962 (N_2962,In_1975,In_1896);
or U2963 (N_2963,In_1711,In_1973);
nor U2964 (N_2964,In_1192,In_1510);
and U2965 (N_2965,In_921,In_1247);
nor U2966 (N_2966,In_1369,In_1645);
xnor U2967 (N_2967,In_1678,In_1337);
nor U2968 (N_2968,In_245,In_1032);
nand U2969 (N_2969,In_413,In_1084);
or U2970 (N_2970,In_2145,In_2359);
xor U2971 (N_2971,In_2363,In_268);
nand U2972 (N_2972,In_1791,In_2241);
xnor U2973 (N_2973,In_150,In_964);
nor U2974 (N_2974,In_292,In_1194);
nor U2975 (N_2975,In_349,In_386);
nand U2976 (N_2976,In_885,In_1582);
and U2977 (N_2977,In_642,In_1814);
or U2978 (N_2978,In_2068,In_803);
and U2979 (N_2979,In_1777,In_1456);
nor U2980 (N_2980,In_1514,In_2419);
nor U2981 (N_2981,In_828,In_1140);
xor U2982 (N_2982,In_686,In_2308);
and U2983 (N_2983,In_137,In_1063);
xor U2984 (N_2984,In_82,In_73);
or U2985 (N_2985,In_1575,In_1686);
and U2986 (N_2986,In_1235,In_1863);
and U2987 (N_2987,In_332,In_721);
and U2988 (N_2988,In_712,In_1840);
nand U2989 (N_2989,In_2462,In_521);
nor U2990 (N_2990,In_1550,In_380);
xnor U2991 (N_2991,In_712,In_486);
and U2992 (N_2992,In_2069,In_590);
nand U2993 (N_2993,In_2149,In_24);
nand U2994 (N_2994,In_1198,In_2414);
xor U2995 (N_2995,In_1160,In_56);
nand U2996 (N_2996,In_1261,In_2472);
or U2997 (N_2997,In_2112,In_1153);
xnor U2998 (N_2998,In_1256,In_1171);
nor U2999 (N_2999,In_2078,In_2180);
and U3000 (N_3000,In_1190,In_1263);
nor U3001 (N_3001,In_2306,In_2195);
nor U3002 (N_3002,In_816,In_647);
and U3003 (N_3003,In_1891,In_220);
nand U3004 (N_3004,In_2392,In_93);
or U3005 (N_3005,In_1049,In_1669);
or U3006 (N_3006,In_1892,In_2427);
xnor U3007 (N_3007,In_2076,In_44);
or U3008 (N_3008,In_663,In_1175);
and U3009 (N_3009,In_267,In_1457);
and U3010 (N_3010,In_2028,In_2073);
or U3011 (N_3011,In_2276,In_261);
nand U3012 (N_3012,In_194,In_1159);
xnor U3013 (N_3013,In_639,In_458);
nor U3014 (N_3014,In_1119,In_1120);
nand U3015 (N_3015,In_1090,In_1326);
or U3016 (N_3016,In_227,In_1849);
nor U3017 (N_3017,In_1810,In_2263);
nor U3018 (N_3018,In_662,In_845);
nor U3019 (N_3019,In_1315,In_79);
nand U3020 (N_3020,In_708,In_1293);
xor U3021 (N_3021,In_404,In_256);
nor U3022 (N_3022,In_1385,In_1450);
nand U3023 (N_3023,In_890,In_2338);
nor U3024 (N_3024,In_422,In_1896);
xor U3025 (N_3025,In_357,In_602);
nand U3026 (N_3026,In_1275,In_1532);
or U3027 (N_3027,In_1882,In_1212);
or U3028 (N_3028,In_2207,In_2204);
nor U3029 (N_3029,In_25,In_1022);
and U3030 (N_3030,In_1027,In_1124);
and U3031 (N_3031,In_1075,In_1307);
nor U3032 (N_3032,In_2316,In_507);
xor U3033 (N_3033,In_1189,In_342);
xnor U3034 (N_3034,In_459,In_950);
xor U3035 (N_3035,In_1259,In_2239);
nor U3036 (N_3036,In_2137,In_880);
or U3037 (N_3037,In_830,In_924);
and U3038 (N_3038,In_762,In_321);
nor U3039 (N_3039,In_1728,In_490);
xor U3040 (N_3040,In_1076,In_2259);
nand U3041 (N_3041,In_2256,In_1407);
and U3042 (N_3042,In_1372,In_1574);
nand U3043 (N_3043,In_2366,In_1346);
nand U3044 (N_3044,In_593,In_595);
nand U3045 (N_3045,In_823,In_2497);
and U3046 (N_3046,In_5,In_1916);
nor U3047 (N_3047,In_232,In_2258);
nor U3048 (N_3048,In_938,In_1755);
and U3049 (N_3049,In_1119,In_1276);
or U3050 (N_3050,In_2040,In_74);
or U3051 (N_3051,In_1826,In_2434);
nor U3052 (N_3052,In_2097,In_1964);
or U3053 (N_3053,In_588,In_257);
nand U3054 (N_3054,In_952,In_2255);
or U3055 (N_3055,In_1738,In_885);
nor U3056 (N_3056,In_2489,In_516);
or U3057 (N_3057,In_1591,In_884);
nor U3058 (N_3058,In_1980,In_711);
nand U3059 (N_3059,In_428,In_2414);
or U3060 (N_3060,In_1341,In_1432);
xor U3061 (N_3061,In_2221,In_297);
nand U3062 (N_3062,In_403,In_1662);
or U3063 (N_3063,In_398,In_1724);
xnor U3064 (N_3064,In_2431,In_1767);
nand U3065 (N_3065,In_1182,In_1264);
xnor U3066 (N_3066,In_1813,In_387);
and U3067 (N_3067,In_1456,In_1577);
and U3068 (N_3068,In_2129,In_2087);
nand U3069 (N_3069,In_997,In_1834);
and U3070 (N_3070,In_1300,In_1356);
nand U3071 (N_3071,In_155,In_895);
or U3072 (N_3072,In_2282,In_114);
nor U3073 (N_3073,In_928,In_7);
xor U3074 (N_3074,In_183,In_635);
and U3075 (N_3075,In_1689,In_1069);
or U3076 (N_3076,In_2066,In_1593);
nand U3077 (N_3077,In_2416,In_392);
and U3078 (N_3078,In_1278,In_1494);
nand U3079 (N_3079,In_2330,In_1832);
xor U3080 (N_3080,In_464,In_557);
xor U3081 (N_3081,In_2343,In_571);
nand U3082 (N_3082,In_2344,In_1629);
xnor U3083 (N_3083,In_2323,In_756);
xor U3084 (N_3084,In_1400,In_1803);
and U3085 (N_3085,In_1010,In_130);
and U3086 (N_3086,In_1390,In_887);
nand U3087 (N_3087,In_306,In_642);
xnor U3088 (N_3088,In_539,In_2458);
nor U3089 (N_3089,In_2245,In_874);
nand U3090 (N_3090,In_50,In_412);
xnor U3091 (N_3091,In_1116,In_1959);
nor U3092 (N_3092,In_636,In_2106);
or U3093 (N_3093,In_155,In_1695);
or U3094 (N_3094,In_2345,In_588);
and U3095 (N_3095,In_1998,In_2312);
nand U3096 (N_3096,In_1114,In_2069);
nand U3097 (N_3097,In_1431,In_362);
xnor U3098 (N_3098,In_1907,In_2464);
nor U3099 (N_3099,In_1628,In_1775);
nor U3100 (N_3100,In_722,In_937);
and U3101 (N_3101,In_456,In_1596);
or U3102 (N_3102,In_2416,In_2195);
nor U3103 (N_3103,In_135,In_1146);
nor U3104 (N_3104,In_2034,In_252);
xnor U3105 (N_3105,In_385,In_889);
or U3106 (N_3106,In_2084,In_225);
nand U3107 (N_3107,In_2487,In_1930);
nor U3108 (N_3108,In_2126,In_1346);
nand U3109 (N_3109,In_468,In_742);
or U3110 (N_3110,In_1488,In_459);
and U3111 (N_3111,In_982,In_547);
nor U3112 (N_3112,In_436,In_134);
or U3113 (N_3113,In_2150,In_1772);
nand U3114 (N_3114,In_1689,In_2456);
xnor U3115 (N_3115,In_705,In_540);
and U3116 (N_3116,In_886,In_1247);
nand U3117 (N_3117,In_1113,In_434);
nor U3118 (N_3118,In_28,In_1383);
or U3119 (N_3119,In_0,In_712);
or U3120 (N_3120,In_1614,In_718);
xor U3121 (N_3121,In_838,In_1712);
nand U3122 (N_3122,In_2478,In_1729);
nand U3123 (N_3123,In_566,In_1093);
or U3124 (N_3124,In_932,In_1079);
and U3125 (N_3125,In_2451,In_368);
nor U3126 (N_3126,In_2447,In_2015);
or U3127 (N_3127,In_1447,In_2251);
xnor U3128 (N_3128,In_968,In_109);
or U3129 (N_3129,In_2,In_2057);
xor U3130 (N_3130,In_1645,In_784);
nand U3131 (N_3131,In_1053,In_2155);
nor U3132 (N_3132,In_1475,In_686);
nor U3133 (N_3133,In_1326,In_526);
nand U3134 (N_3134,In_385,In_1256);
nor U3135 (N_3135,In_752,In_1470);
and U3136 (N_3136,In_975,In_377);
nor U3137 (N_3137,In_2027,In_1012);
xor U3138 (N_3138,In_2396,In_872);
and U3139 (N_3139,In_561,In_1662);
xnor U3140 (N_3140,In_573,In_1304);
xnor U3141 (N_3141,In_95,In_1111);
and U3142 (N_3142,In_623,In_349);
or U3143 (N_3143,In_1644,In_984);
or U3144 (N_3144,In_1698,In_561);
nand U3145 (N_3145,In_2304,In_2188);
and U3146 (N_3146,In_2088,In_1027);
and U3147 (N_3147,In_840,In_2266);
nor U3148 (N_3148,In_1799,In_229);
nand U3149 (N_3149,In_1389,In_543);
or U3150 (N_3150,In_1180,In_1990);
and U3151 (N_3151,In_195,In_1237);
and U3152 (N_3152,In_1247,In_94);
nor U3153 (N_3153,In_1513,In_374);
nor U3154 (N_3154,In_1009,In_1853);
and U3155 (N_3155,In_138,In_2430);
or U3156 (N_3156,In_139,In_1272);
nand U3157 (N_3157,In_2222,In_1005);
or U3158 (N_3158,In_1321,In_1474);
nor U3159 (N_3159,In_1039,In_240);
or U3160 (N_3160,In_684,In_1153);
or U3161 (N_3161,In_1134,In_125);
or U3162 (N_3162,In_2396,In_2323);
nand U3163 (N_3163,In_725,In_1260);
nand U3164 (N_3164,In_223,In_2382);
nand U3165 (N_3165,In_25,In_342);
nor U3166 (N_3166,In_1725,In_1061);
or U3167 (N_3167,In_2130,In_1184);
nand U3168 (N_3168,In_208,In_2024);
nor U3169 (N_3169,In_2162,In_381);
and U3170 (N_3170,In_1019,In_529);
xor U3171 (N_3171,In_413,In_2417);
nor U3172 (N_3172,In_2311,In_94);
and U3173 (N_3173,In_1652,In_814);
or U3174 (N_3174,In_2061,In_587);
nor U3175 (N_3175,In_1565,In_1445);
nor U3176 (N_3176,In_1299,In_233);
and U3177 (N_3177,In_1194,In_1907);
xnor U3178 (N_3178,In_1052,In_294);
nor U3179 (N_3179,In_940,In_2071);
nand U3180 (N_3180,In_307,In_2092);
nor U3181 (N_3181,In_487,In_1885);
xor U3182 (N_3182,In_1740,In_906);
or U3183 (N_3183,In_1123,In_682);
nor U3184 (N_3184,In_855,In_2058);
nor U3185 (N_3185,In_2428,In_88);
xnor U3186 (N_3186,In_2229,In_1114);
nor U3187 (N_3187,In_1518,In_847);
and U3188 (N_3188,In_2263,In_1260);
xor U3189 (N_3189,In_1903,In_1799);
or U3190 (N_3190,In_2199,In_2197);
xor U3191 (N_3191,In_872,In_2152);
xor U3192 (N_3192,In_2395,In_874);
or U3193 (N_3193,In_629,In_2149);
nand U3194 (N_3194,In_400,In_1305);
or U3195 (N_3195,In_1740,In_358);
and U3196 (N_3196,In_477,In_1795);
xor U3197 (N_3197,In_2048,In_1730);
nand U3198 (N_3198,In_668,In_887);
nor U3199 (N_3199,In_237,In_2244);
nor U3200 (N_3200,In_1808,In_298);
and U3201 (N_3201,In_1851,In_195);
nor U3202 (N_3202,In_103,In_2132);
nand U3203 (N_3203,In_691,In_1755);
xor U3204 (N_3204,In_2489,In_443);
nor U3205 (N_3205,In_140,In_2495);
and U3206 (N_3206,In_1935,In_310);
or U3207 (N_3207,In_1291,In_2407);
and U3208 (N_3208,In_1337,In_2147);
nand U3209 (N_3209,In_648,In_266);
nor U3210 (N_3210,In_1273,In_586);
or U3211 (N_3211,In_2383,In_562);
nand U3212 (N_3212,In_670,In_1106);
xnor U3213 (N_3213,In_793,In_678);
and U3214 (N_3214,In_137,In_1362);
or U3215 (N_3215,In_191,In_1307);
xor U3216 (N_3216,In_270,In_278);
and U3217 (N_3217,In_237,In_489);
and U3218 (N_3218,In_2487,In_1373);
nand U3219 (N_3219,In_1566,In_650);
xnor U3220 (N_3220,In_106,In_849);
or U3221 (N_3221,In_2278,In_884);
or U3222 (N_3222,In_1056,In_505);
nor U3223 (N_3223,In_1619,In_1137);
nor U3224 (N_3224,In_1612,In_2120);
nand U3225 (N_3225,In_1197,In_1642);
or U3226 (N_3226,In_1316,In_33);
or U3227 (N_3227,In_524,In_1853);
nand U3228 (N_3228,In_1659,In_1547);
and U3229 (N_3229,In_2387,In_1493);
and U3230 (N_3230,In_1827,In_1229);
nor U3231 (N_3231,In_1717,In_883);
and U3232 (N_3232,In_901,In_1030);
nor U3233 (N_3233,In_1492,In_2192);
nor U3234 (N_3234,In_1858,In_711);
nor U3235 (N_3235,In_306,In_49);
xor U3236 (N_3236,In_1652,In_25);
nor U3237 (N_3237,In_180,In_2019);
nor U3238 (N_3238,In_332,In_1936);
nand U3239 (N_3239,In_1494,In_1217);
nand U3240 (N_3240,In_2352,In_819);
nand U3241 (N_3241,In_219,In_717);
nor U3242 (N_3242,In_66,In_371);
and U3243 (N_3243,In_360,In_1760);
nor U3244 (N_3244,In_1186,In_1829);
nor U3245 (N_3245,In_1071,In_2115);
nand U3246 (N_3246,In_764,In_554);
nand U3247 (N_3247,In_1494,In_167);
nand U3248 (N_3248,In_2224,In_1857);
nand U3249 (N_3249,In_856,In_2179);
or U3250 (N_3250,In_2221,In_1191);
xor U3251 (N_3251,In_1202,In_807);
xor U3252 (N_3252,In_1729,In_498);
and U3253 (N_3253,In_2378,In_1716);
nor U3254 (N_3254,In_2246,In_260);
and U3255 (N_3255,In_856,In_735);
nor U3256 (N_3256,In_643,In_992);
nand U3257 (N_3257,In_1416,In_301);
xor U3258 (N_3258,In_2063,In_2074);
nor U3259 (N_3259,In_657,In_452);
and U3260 (N_3260,In_2481,In_991);
or U3261 (N_3261,In_517,In_239);
or U3262 (N_3262,In_555,In_1473);
or U3263 (N_3263,In_1795,In_226);
or U3264 (N_3264,In_1444,In_420);
xnor U3265 (N_3265,In_513,In_1657);
nand U3266 (N_3266,In_1658,In_2277);
nand U3267 (N_3267,In_68,In_1711);
xor U3268 (N_3268,In_1580,In_942);
nand U3269 (N_3269,In_1687,In_450);
or U3270 (N_3270,In_2348,In_1291);
nor U3271 (N_3271,In_1628,In_822);
nor U3272 (N_3272,In_770,In_559);
nor U3273 (N_3273,In_182,In_2059);
xnor U3274 (N_3274,In_1915,In_1336);
or U3275 (N_3275,In_2466,In_1977);
or U3276 (N_3276,In_1645,In_1003);
and U3277 (N_3277,In_502,In_1848);
or U3278 (N_3278,In_1498,In_2283);
xor U3279 (N_3279,In_2363,In_256);
xnor U3280 (N_3280,In_217,In_705);
nand U3281 (N_3281,In_971,In_553);
and U3282 (N_3282,In_1164,In_323);
nor U3283 (N_3283,In_1509,In_2271);
xor U3284 (N_3284,In_1298,In_87);
xnor U3285 (N_3285,In_1177,In_1369);
or U3286 (N_3286,In_1453,In_2066);
and U3287 (N_3287,In_91,In_753);
xor U3288 (N_3288,In_106,In_1875);
and U3289 (N_3289,In_304,In_407);
nand U3290 (N_3290,In_2415,In_2159);
or U3291 (N_3291,In_2250,In_1580);
and U3292 (N_3292,In_1893,In_2472);
and U3293 (N_3293,In_1101,In_1256);
or U3294 (N_3294,In_1667,In_1119);
or U3295 (N_3295,In_1556,In_901);
nand U3296 (N_3296,In_1934,In_643);
xnor U3297 (N_3297,In_0,In_1671);
or U3298 (N_3298,In_1797,In_4);
nand U3299 (N_3299,In_594,In_777);
or U3300 (N_3300,In_467,In_60);
nand U3301 (N_3301,In_473,In_1398);
and U3302 (N_3302,In_1541,In_1728);
nand U3303 (N_3303,In_1930,In_1547);
xnor U3304 (N_3304,In_1644,In_220);
xor U3305 (N_3305,In_2248,In_1666);
xor U3306 (N_3306,In_1339,In_350);
xor U3307 (N_3307,In_2190,In_1681);
and U3308 (N_3308,In_582,In_1209);
xnor U3309 (N_3309,In_2228,In_2400);
xor U3310 (N_3310,In_1520,In_2016);
nor U3311 (N_3311,In_663,In_1224);
or U3312 (N_3312,In_1151,In_435);
and U3313 (N_3313,In_1340,In_249);
nor U3314 (N_3314,In_601,In_2302);
or U3315 (N_3315,In_1917,In_617);
xor U3316 (N_3316,In_1616,In_735);
or U3317 (N_3317,In_446,In_1088);
xnor U3318 (N_3318,In_696,In_1607);
and U3319 (N_3319,In_41,In_707);
nor U3320 (N_3320,In_8,In_2075);
and U3321 (N_3321,In_1219,In_2251);
and U3322 (N_3322,In_84,In_369);
and U3323 (N_3323,In_1129,In_1738);
and U3324 (N_3324,In_312,In_66);
xnor U3325 (N_3325,In_1222,In_30);
or U3326 (N_3326,In_2080,In_1786);
xnor U3327 (N_3327,In_1837,In_1629);
and U3328 (N_3328,In_1423,In_1446);
xor U3329 (N_3329,In_2022,In_1671);
nand U3330 (N_3330,In_1687,In_1215);
xnor U3331 (N_3331,In_16,In_1917);
and U3332 (N_3332,In_2266,In_1971);
and U3333 (N_3333,In_1041,In_1285);
nor U3334 (N_3334,In_42,In_1682);
or U3335 (N_3335,In_765,In_1449);
nand U3336 (N_3336,In_2401,In_86);
xor U3337 (N_3337,In_2463,In_237);
xor U3338 (N_3338,In_2403,In_2090);
xor U3339 (N_3339,In_1558,In_1701);
and U3340 (N_3340,In_2022,In_1218);
nor U3341 (N_3341,In_330,In_1160);
xor U3342 (N_3342,In_487,In_2179);
and U3343 (N_3343,In_1185,In_2110);
nand U3344 (N_3344,In_563,In_1726);
xor U3345 (N_3345,In_1989,In_2188);
nand U3346 (N_3346,In_1395,In_457);
and U3347 (N_3347,In_639,In_2047);
or U3348 (N_3348,In_1336,In_268);
xor U3349 (N_3349,In_2333,In_705);
xnor U3350 (N_3350,In_334,In_1966);
xnor U3351 (N_3351,In_1454,In_1288);
and U3352 (N_3352,In_1507,In_744);
nand U3353 (N_3353,In_310,In_262);
nor U3354 (N_3354,In_1359,In_749);
nand U3355 (N_3355,In_1432,In_1748);
nand U3356 (N_3356,In_2172,In_1292);
nand U3357 (N_3357,In_1215,In_2425);
or U3358 (N_3358,In_1234,In_1918);
xnor U3359 (N_3359,In_2392,In_1460);
nand U3360 (N_3360,In_2336,In_725);
or U3361 (N_3361,In_1131,In_1574);
nand U3362 (N_3362,In_1353,In_2221);
or U3363 (N_3363,In_1360,In_1371);
nor U3364 (N_3364,In_938,In_1901);
and U3365 (N_3365,In_470,In_27);
nand U3366 (N_3366,In_2162,In_579);
and U3367 (N_3367,In_670,In_541);
xnor U3368 (N_3368,In_1828,In_2038);
nor U3369 (N_3369,In_839,In_588);
xor U3370 (N_3370,In_1085,In_2367);
or U3371 (N_3371,In_2216,In_1091);
xnor U3372 (N_3372,In_1549,In_2033);
or U3373 (N_3373,In_1009,In_78);
nand U3374 (N_3374,In_2483,In_853);
nand U3375 (N_3375,In_1895,In_1465);
nand U3376 (N_3376,In_1809,In_1311);
nor U3377 (N_3377,In_1891,In_995);
and U3378 (N_3378,In_1758,In_163);
or U3379 (N_3379,In_2426,In_787);
or U3380 (N_3380,In_967,In_1405);
nand U3381 (N_3381,In_472,In_414);
nand U3382 (N_3382,In_51,In_1097);
nand U3383 (N_3383,In_386,In_1821);
xor U3384 (N_3384,In_402,In_2242);
or U3385 (N_3385,In_734,In_2324);
and U3386 (N_3386,In_1829,In_736);
nor U3387 (N_3387,In_1989,In_412);
nor U3388 (N_3388,In_1179,In_237);
xor U3389 (N_3389,In_1365,In_1280);
nand U3390 (N_3390,In_2290,In_813);
nand U3391 (N_3391,In_546,In_624);
and U3392 (N_3392,In_2216,In_583);
nor U3393 (N_3393,In_507,In_2103);
and U3394 (N_3394,In_767,In_1630);
nand U3395 (N_3395,In_1347,In_1183);
and U3396 (N_3396,In_1103,In_1247);
or U3397 (N_3397,In_1989,In_121);
nor U3398 (N_3398,In_162,In_1652);
and U3399 (N_3399,In_123,In_285);
nor U3400 (N_3400,In_485,In_1284);
xnor U3401 (N_3401,In_1250,In_1417);
or U3402 (N_3402,In_792,In_1192);
xor U3403 (N_3403,In_1831,In_590);
and U3404 (N_3404,In_186,In_2040);
xnor U3405 (N_3405,In_1020,In_104);
xor U3406 (N_3406,In_658,In_2008);
nor U3407 (N_3407,In_138,In_1735);
xnor U3408 (N_3408,In_1773,In_301);
or U3409 (N_3409,In_879,In_2233);
nand U3410 (N_3410,In_36,In_1911);
and U3411 (N_3411,In_1570,In_2342);
xnor U3412 (N_3412,In_662,In_1608);
nor U3413 (N_3413,In_642,In_1507);
xor U3414 (N_3414,In_1362,In_438);
or U3415 (N_3415,In_1844,In_1211);
xnor U3416 (N_3416,In_974,In_1285);
or U3417 (N_3417,In_1162,In_2363);
nor U3418 (N_3418,In_1972,In_2201);
nand U3419 (N_3419,In_175,In_352);
or U3420 (N_3420,In_2461,In_476);
nand U3421 (N_3421,In_2005,In_1956);
nand U3422 (N_3422,In_241,In_2187);
nand U3423 (N_3423,In_557,In_1908);
nand U3424 (N_3424,In_970,In_665);
or U3425 (N_3425,In_1180,In_1894);
xor U3426 (N_3426,In_1368,In_1280);
or U3427 (N_3427,In_964,In_548);
xor U3428 (N_3428,In_1890,In_2353);
or U3429 (N_3429,In_2215,In_1497);
xor U3430 (N_3430,In_1691,In_2262);
xnor U3431 (N_3431,In_1578,In_1882);
xor U3432 (N_3432,In_1082,In_303);
and U3433 (N_3433,In_32,In_1255);
nand U3434 (N_3434,In_2441,In_352);
nand U3435 (N_3435,In_2229,In_1118);
nand U3436 (N_3436,In_864,In_528);
nor U3437 (N_3437,In_1266,In_279);
and U3438 (N_3438,In_1070,In_1623);
xnor U3439 (N_3439,In_1877,In_264);
nor U3440 (N_3440,In_10,In_2430);
nand U3441 (N_3441,In_2175,In_1669);
nand U3442 (N_3442,In_2387,In_1601);
nor U3443 (N_3443,In_2313,In_7);
or U3444 (N_3444,In_307,In_2224);
nand U3445 (N_3445,In_2092,In_1669);
nor U3446 (N_3446,In_2309,In_1695);
or U3447 (N_3447,In_1556,In_91);
xor U3448 (N_3448,In_816,In_2258);
nand U3449 (N_3449,In_2217,In_1823);
or U3450 (N_3450,In_1593,In_81);
nand U3451 (N_3451,In_1059,In_2437);
nand U3452 (N_3452,In_1926,In_814);
xnor U3453 (N_3453,In_2283,In_1248);
nor U3454 (N_3454,In_519,In_1531);
nand U3455 (N_3455,In_2041,In_989);
xor U3456 (N_3456,In_67,In_1135);
nor U3457 (N_3457,In_522,In_2269);
or U3458 (N_3458,In_658,In_211);
nand U3459 (N_3459,In_1879,In_1107);
nand U3460 (N_3460,In_252,In_266);
and U3461 (N_3461,In_1803,In_2092);
or U3462 (N_3462,In_2078,In_954);
xnor U3463 (N_3463,In_1905,In_1577);
and U3464 (N_3464,In_842,In_1632);
and U3465 (N_3465,In_2443,In_1071);
nor U3466 (N_3466,In_2355,In_1486);
nand U3467 (N_3467,In_1647,In_953);
nand U3468 (N_3468,In_1095,In_262);
or U3469 (N_3469,In_705,In_933);
xnor U3470 (N_3470,In_670,In_1590);
xor U3471 (N_3471,In_2245,In_623);
or U3472 (N_3472,In_502,In_153);
nor U3473 (N_3473,In_2466,In_2201);
or U3474 (N_3474,In_297,In_1852);
nand U3475 (N_3475,In_907,In_2465);
xnor U3476 (N_3476,In_653,In_217);
nor U3477 (N_3477,In_732,In_721);
nand U3478 (N_3478,In_2014,In_533);
xnor U3479 (N_3479,In_702,In_512);
and U3480 (N_3480,In_315,In_2455);
nor U3481 (N_3481,In_1721,In_652);
and U3482 (N_3482,In_2134,In_219);
nor U3483 (N_3483,In_2045,In_2406);
nor U3484 (N_3484,In_1391,In_1013);
or U3485 (N_3485,In_37,In_92);
xnor U3486 (N_3486,In_1577,In_1655);
or U3487 (N_3487,In_1207,In_505);
nor U3488 (N_3488,In_643,In_2222);
or U3489 (N_3489,In_1453,In_2292);
nand U3490 (N_3490,In_1666,In_461);
nand U3491 (N_3491,In_569,In_1712);
nor U3492 (N_3492,In_1461,In_1111);
xor U3493 (N_3493,In_1011,In_2387);
and U3494 (N_3494,In_1839,In_114);
xor U3495 (N_3495,In_1216,In_2225);
or U3496 (N_3496,In_136,In_1150);
nand U3497 (N_3497,In_1360,In_1546);
or U3498 (N_3498,In_41,In_961);
nand U3499 (N_3499,In_219,In_591);
xnor U3500 (N_3500,In_815,In_517);
and U3501 (N_3501,In_932,In_2008);
nor U3502 (N_3502,In_2267,In_2410);
xnor U3503 (N_3503,In_595,In_1787);
and U3504 (N_3504,In_92,In_524);
nand U3505 (N_3505,In_1163,In_238);
nand U3506 (N_3506,In_82,In_1627);
nand U3507 (N_3507,In_204,In_1317);
nor U3508 (N_3508,In_1973,In_561);
and U3509 (N_3509,In_1430,In_1999);
nand U3510 (N_3510,In_94,In_502);
or U3511 (N_3511,In_1308,In_1480);
and U3512 (N_3512,In_2271,In_1066);
and U3513 (N_3513,In_105,In_919);
and U3514 (N_3514,In_1522,In_1734);
nor U3515 (N_3515,In_1961,In_1373);
nor U3516 (N_3516,In_517,In_2484);
or U3517 (N_3517,In_1208,In_1618);
or U3518 (N_3518,In_2207,In_2464);
nor U3519 (N_3519,In_1422,In_512);
or U3520 (N_3520,In_283,In_272);
xor U3521 (N_3521,In_246,In_2266);
and U3522 (N_3522,In_2367,In_1859);
or U3523 (N_3523,In_445,In_2452);
and U3524 (N_3524,In_1159,In_2384);
and U3525 (N_3525,In_113,In_2215);
and U3526 (N_3526,In_156,In_1107);
nand U3527 (N_3527,In_375,In_941);
nand U3528 (N_3528,In_2089,In_236);
nand U3529 (N_3529,In_1539,In_681);
nand U3530 (N_3530,In_1898,In_258);
or U3531 (N_3531,In_1532,In_1364);
xor U3532 (N_3532,In_110,In_138);
xor U3533 (N_3533,In_382,In_863);
nor U3534 (N_3534,In_1431,In_404);
or U3535 (N_3535,In_202,In_1397);
nor U3536 (N_3536,In_1862,In_192);
xnor U3537 (N_3537,In_566,In_2081);
xor U3538 (N_3538,In_926,In_1218);
xnor U3539 (N_3539,In_2277,In_1499);
xor U3540 (N_3540,In_269,In_1474);
or U3541 (N_3541,In_1162,In_2040);
and U3542 (N_3542,In_2466,In_566);
xor U3543 (N_3543,In_2020,In_1995);
or U3544 (N_3544,In_578,In_1824);
or U3545 (N_3545,In_176,In_1904);
nand U3546 (N_3546,In_2042,In_411);
and U3547 (N_3547,In_1956,In_375);
or U3548 (N_3548,In_701,In_928);
and U3549 (N_3549,In_681,In_1612);
xnor U3550 (N_3550,In_427,In_1177);
nor U3551 (N_3551,In_1783,In_2127);
and U3552 (N_3552,In_1102,In_2174);
and U3553 (N_3553,In_2425,In_424);
xnor U3554 (N_3554,In_863,In_701);
and U3555 (N_3555,In_276,In_989);
xnor U3556 (N_3556,In_349,In_999);
xor U3557 (N_3557,In_358,In_1258);
or U3558 (N_3558,In_749,In_1898);
or U3559 (N_3559,In_695,In_1605);
nand U3560 (N_3560,In_1601,In_1216);
nor U3561 (N_3561,In_1541,In_563);
nor U3562 (N_3562,In_1010,In_1846);
nor U3563 (N_3563,In_2022,In_2354);
nor U3564 (N_3564,In_2307,In_1593);
nor U3565 (N_3565,In_142,In_245);
xor U3566 (N_3566,In_415,In_462);
nand U3567 (N_3567,In_3,In_541);
nand U3568 (N_3568,In_2031,In_1138);
and U3569 (N_3569,In_2067,In_1947);
and U3570 (N_3570,In_1272,In_2470);
or U3571 (N_3571,In_1970,In_2343);
and U3572 (N_3572,In_108,In_914);
nand U3573 (N_3573,In_2435,In_967);
nor U3574 (N_3574,In_1926,In_1505);
or U3575 (N_3575,In_311,In_734);
and U3576 (N_3576,In_1612,In_1538);
nand U3577 (N_3577,In_2068,In_1772);
or U3578 (N_3578,In_751,In_2458);
nor U3579 (N_3579,In_1679,In_490);
xor U3580 (N_3580,In_361,In_66);
or U3581 (N_3581,In_1834,In_817);
and U3582 (N_3582,In_6,In_25);
nor U3583 (N_3583,In_1232,In_1615);
nand U3584 (N_3584,In_2488,In_1173);
nand U3585 (N_3585,In_1410,In_335);
and U3586 (N_3586,In_1805,In_1711);
nor U3587 (N_3587,In_198,In_1854);
or U3588 (N_3588,In_360,In_665);
or U3589 (N_3589,In_254,In_2201);
and U3590 (N_3590,In_2372,In_1663);
nand U3591 (N_3591,In_2030,In_522);
and U3592 (N_3592,In_1597,In_699);
xor U3593 (N_3593,In_886,In_1631);
or U3594 (N_3594,In_1544,In_1208);
nor U3595 (N_3595,In_1519,In_1674);
nand U3596 (N_3596,In_92,In_710);
and U3597 (N_3597,In_770,In_329);
or U3598 (N_3598,In_2126,In_156);
and U3599 (N_3599,In_381,In_2208);
nor U3600 (N_3600,In_1986,In_1454);
or U3601 (N_3601,In_859,In_1380);
nor U3602 (N_3602,In_818,In_1276);
and U3603 (N_3603,In_469,In_359);
nor U3604 (N_3604,In_2240,In_1159);
or U3605 (N_3605,In_1773,In_1892);
nand U3606 (N_3606,In_853,In_1622);
nand U3607 (N_3607,In_1306,In_2028);
and U3608 (N_3608,In_2145,In_423);
nor U3609 (N_3609,In_803,In_1016);
or U3610 (N_3610,In_1645,In_1835);
xor U3611 (N_3611,In_27,In_2214);
nand U3612 (N_3612,In_1686,In_1288);
and U3613 (N_3613,In_304,In_372);
xnor U3614 (N_3614,In_1609,In_2406);
and U3615 (N_3615,In_559,In_1982);
or U3616 (N_3616,In_415,In_1572);
xnor U3617 (N_3617,In_2275,In_459);
and U3618 (N_3618,In_2345,In_2237);
and U3619 (N_3619,In_2365,In_2128);
nand U3620 (N_3620,In_32,In_809);
and U3621 (N_3621,In_2024,In_2319);
nand U3622 (N_3622,In_2010,In_2278);
xor U3623 (N_3623,In_918,In_975);
and U3624 (N_3624,In_226,In_2332);
xnor U3625 (N_3625,In_1756,In_330);
and U3626 (N_3626,In_597,In_1256);
or U3627 (N_3627,In_2062,In_909);
nand U3628 (N_3628,In_1864,In_2462);
or U3629 (N_3629,In_1570,In_555);
or U3630 (N_3630,In_2254,In_1508);
xor U3631 (N_3631,In_342,In_96);
xor U3632 (N_3632,In_1920,In_1765);
or U3633 (N_3633,In_796,In_434);
xor U3634 (N_3634,In_1894,In_1290);
or U3635 (N_3635,In_2275,In_10);
xnor U3636 (N_3636,In_894,In_1352);
xor U3637 (N_3637,In_1944,In_1290);
and U3638 (N_3638,In_1442,In_751);
nor U3639 (N_3639,In_895,In_1041);
and U3640 (N_3640,In_1428,In_2120);
or U3641 (N_3641,In_2382,In_252);
xor U3642 (N_3642,In_875,In_458);
nand U3643 (N_3643,In_16,In_992);
or U3644 (N_3644,In_2112,In_2257);
xor U3645 (N_3645,In_1981,In_663);
xnor U3646 (N_3646,In_1517,In_258);
nor U3647 (N_3647,In_604,In_230);
and U3648 (N_3648,In_1689,In_931);
xor U3649 (N_3649,In_1638,In_346);
and U3650 (N_3650,In_2336,In_1216);
nor U3651 (N_3651,In_714,In_811);
nand U3652 (N_3652,In_604,In_1756);
xnor U3653 (N_3653,In_1128,In_1009);
nand U3654 (N_3654,In_1196,In_2209);
or U3655 (N_3655,In_377,In_2282);
and U3656 (N_3656,In_1018,In_2034);
or U3657 (N_3657,In_1288,In_1679);
or U3658 (N_3658,In_1625,In_1432);
and U3659 (N_3659,In_1990,In_981);
nand U3660 (N_3660,In_1143,In_1576);
nor U3661 (N_3661,In_2093,In_1054);
and U3662 (N_3662,In_1929,In_1020);
nor U3663 (N_3663,In_2253,In_1510);
nor U3664 (N_3664,In_1508,In_2195);
nor U3665 (N_3665,In_2179,In_2119);
xnor U3666 (N_3666,In_250,In_1643);
or U3667 (N_3667,In_582,In_876);
or U3668 (N_3668,In_1483,In_1926);
and U3669 (N_3669,In_1585,In_1757);
or U3670 (N_3670,In_2178,In_2005);
nor U3671 (N_3671,In_364,In_1114);
xnor U3672 (N_3672,In_1814,In_470);
and U3673 (N_3673,In_300,In_1521);
and U3674 (N_3674,In_897,In_418);
nand U3675 (N_3675,In_2071,In_12);
and U3676 (N_3676,In_339,In_2065);
or U3677 (N_3677,In_1940,In_934);
and U3678 (N_3678,In_1788,In_1775);
nor U3679 (N_3679,In_2288,In_2457);
nand U3680 (N_3680,In_1371,In_1353);
nand U3681 (N_3681,In_1117,In_856);
and U3682 (N_3682,In_177,In_2228);
or U3683 (N_3683,In_926,In_2432);
xor U3684 (N_3684,In_1538,In_1477);
nor U3685 (N_3685,In_59,In_370);
xnor U3686 (N_3686,In_1656,In_362);
and U3687 (N_3687,In_2149,In_1813);
and U3688 (N_3688,In_284,In_312);
and U3689 (N_3689,In_337,In_124);
or U3690 (N_3690,In_1874,In_1598);
nand U3691 (N_3691,In_1283,In_2283);
and U3692 (N_3692,In_1366,In_1567);
or U3693 (N_3693,In_1048,In_1042);
xor U3694 (N_3694,In_1494,In_2265);
nor U3695 (N_3695,In_654,In_1667);
or U3696 (N_3696,In_1013,In_2476);
or U3697 (N_3697,In_2498,In_2164);
and U3698 (N_3698,In_1821,In_1066);
xor U3699 (N_3699,In_352,In_187);
xnor U3700 (N_3700,In_2123,In_2254);
nor U3701 (N_3701,In_1494,In_238);
xnor U3702 (N_3702,In_1994,In_658);
or U3703 (N_3703,In_1719,In_1093);
nor U3704 (N_3704,In_1956,In_103);
xnor U3705 (N_3705,In_1515,In_1585);
nor U3706 (N_3706,In_2121,In_2196);
and U3707 (N_3707,In_534,In_753);
nand U3708 (N_3708,In_909,In_1877);
xor U3709 (N_3709,In_2186,In_1881);
or U3710 (N_3710,In_1982,In_335);
and U3711 (N_3711,In_634,In_754);
xor U3712 (N_3712,In_353,In_2311);
and U3713 (N_3713,In_2087,In_256);
nor U3714 (N_3714,In_392,In_1882);
nand U3715 (N_3715,In_2022,In_326);
and U3716 (N_3716,In_1066,In_1022);
xnor U3717 (N_3717,In_620,In_1080);
xnor U3718 (N_3718,In_1006,In_189);
or U3719 (N_3719,In_1418,In_1620);
xnor U3720 (N_3720,In_573,In_691);
or U3721 (N_3721,In_490,In_686);
nand U3722 (N_3722,In_346,In_1973);
xor U3723 (N_3723,In_2368,In_1246);
nand U3724 (N_3724,In_1518,In_742);
xnor U3725 (N_3725,In_2022,In_2326);
xnor U3726 (N_3726,In_887,In_653);
nor U3727 (N_3727,In_2430,In_767);
and U3728 (N_3728,In_1902,In_1439);
nand U3729 (N_3729,In_126,In_613);
nand U3730 (N_3730,In_207,In_2149);
nand U3731 (N_3731,In_2332,In_1074);
and U3732 (N_3732,In_875,In_593);
nand U3733 (N_3733,In_1177,In_516);
or U3734 (N_3734,In_776,In_861);
nor U3735 (N_3735,In_2428,In_1052);
and U3736 (N_3736,In_326,In_1249);
nand U3737 (N_3737,In_949,In_1131);
xnor U3738 (N_3738,In_829,In_256);
xor U3739 (N_3739,In_2187,In_2401);
nand U3740 (N_3740,In_1295,In_1098);
and U3741 (N_3741,In_2285,In_783);
and U3742 (N_3742,In_61,In_796);
nor U3743 (N_3743,In_204,In_1024);
nand U3744 (N_3744,In_694,In_1751);
and U3745 (N_3745,In_1641,In_432);
and U3746 (N_3746,In_1020,In_2249);
or U3747 (N_3747,In_1697,In_1132);
xor U3748 (N_3748,In_311,In_147);
and U3749 (N_3749,In_329,In_2201);
nand U3750 (N_3750,In_2119,In_1328);
xnor U3751 (N_3751,In_1527,In_2479);
and U3752 (N_3752,In_1514,In_1002);
nor U3753 (N_3753,In_1744,In_1590);
and U3754 (N_3754,In_82,In_906);
nor U3755 (N_3755,In_732,In_1686);
and U3756 (N_3756,In_1595,In_1693);
and U3757 (N_3757,In_901,In_2050);
and U3758 (N_3758,In_1496,In_531);
and U3759 (N_3759,In_2255,In_1635);
xor U3760 (N_3760,In_1942,In_1044);
nand U3761 (N_3761,In_731,In_1397);
nand U3762 (N_3762,In_1119,In_776);
nor U3763 (N_3763,In_2177,In_2103);
nor U3764 (N_3764,In_1479,In_537);
nor U3765 (N_3765,In_2119,In_138);
xor U3766 (N_3766,In_997,In_267);
nand U3767 (N_3767,In_1034,In_546);
nand U3768 (N_3768,In_1118,In_1377);
and U3769 (N_3769,In_1342,In_2286);
nor U3770 (N_3770,In_833,In_836);
nor U3771 (N_3771,In_911,In_1778);
nor U3772 (N_3772,In_649,In_261);
nor U3773 (N_3773,In_1119,In_939);
xor U3774 (N_3774,In_946,In_101);
or U3775 (N_3775,In_1109,In_2214);
and U3776 (N_3776,In_806,In_391);
and U3777 (N_3777,In_1261,In_1356);
xor U3778 (N_3778,In_1590,In_816);
or U3779 (N_3779,In_714,In_2256);
nand U3780 (N_3780,In_1256,In_472);
nand U3781 (N_3781,In_935,In_1616);
nand U3782 (N_3782,In_476,In_929);
nand U3783 (N_3783,In_1782,In_2030);
and U3784 (N_3784,In_1804,In_1995);
and U3785 (N_3785,In_1239,In_1193);
nor U3786 (N_3786,In_2051,In_2433);
nor U3787 (N_3787,In_51,In_198);
and U3788 (N_3788,In_592,In_2063);
or U3789 (N_3789,In_1360,In_1670);
or U3790 (N_3790,In_1589,In_1736);
or U3791 (N_3791,In_2342,In_187);
and U3792 (N_3792,In_261,In_1924);
xor U3793 (N_3793,In_2131,In_1541);
nand U3794 (N_3794,In_2273,In_1230);
xor U3795 (N_3795,In_1136,In_488);
xor U3796 (N_3796,In_193,In_2150);
xor U3797 (N_3797,In_2443,In_1626);
and U3798 (N_3798,In_2460,In_544);
or U3799 (N_3799,In_1800,In_579);
and U3800 (N_3800,In_665,In_1256);
and U3801 (N_3801,In_2052,In_2353);
xnor U3802 (N_3802,In_2087,In_2);
or U3803 (N_3803,In_555,In_1337);
nor U3804 (N_3804,In_479,In_785);
and U3805 (N_3805,In_1575,In_1992);
and U3806 (N_3806,In_997,In_2469);
or U3807 (N_3807,In_1873,In_1140);
nand U3808 (N_3808,In_1884,In_324);
xor U3809 (N_3809,In_655,In_1331);
xnor U3810 (N_3810,In_199,In_327);
or U3811 (N_3811,In_569,In_1829);
nand U3812 (N_3812,In_2156,In_1258);
nor U3813 (N_3813,In_163,In_2415);
and U3814 (N_3814,In_2439,In_431);
nand U3815 (N_3815,In_2024,In_2437);
nand U3816 (N_3816,In_2287,In_799);
xor U3817 (N_3817,In_1086,In_1195);
xor U3818 (N_3818,In_516,In_1837);
xor U3819 (N_3819,In_361,In_2305);
and U3820 (N_3820,In_1189,In_1521);
xnor U3821 (N_3821,In_2441,In_2363);
nand U3822 (N_3822,In_786,In_2051);
xnor U3823 (N_3823,In_90,In_1141);
nor U3824 (N_3824,In_1134,In_857);
nor U3825 (N_3825,In_1109,In_1446);
nor U3826 (N_3826,In_1514,In_328);
and U3827 (N_3827,In_789,In_1954);
and U3828 (N_3828,In_2290,In_1848);
or U3829 (N_3829,In_1849,In_925);
or U3830 (N_3830,In_2130,In_342);
nand U3831 (N_3831,In_1355,In_2318);
xnor U3832 (N_3832,In_381,In_1756);
xor U3833 (N_3833,In_67,In_468);
or U3834 (N_3834,In_2,In_1590);
or U3835 (N_3835,In_689,In_2459);
and U3836 (N_3836,In_2136,In_1486);
xnor U3837 (N_3837,In_1016,In_2390);
nor U3838 (N_3838,In_609,In_1987);
nand U3839 (N_3839,In_75,In_1040);
and U3840 (N_3840,In_2266,In_2151);
xnor U3841 (N_3841,In_2025,In_1753);
nand U3842 (N_3842,In_239,In_1763);
nand U3843 (N_3843,In_2040,In_1676);
nand U3844 (N_3844,In_2065,In_1036);
or U3845 (N_3845,In_1885,In_2181);
or U3846 (N_3846,In_2214,In_2351);
and U3847 (N_3847,In_2290,In_1743);
nor U3848 (N_3848,In_133,In_2121);
nand U3849 (N_3849,In_656,In_1712);
xor U3850 (N_3850,In_1095,In_2430);
xor U3851 (N_3851,In_91,In_1341);
or U3852 (N_3852,In_2185,In_13);
and U3853 (N_3853,In_656,In_1785);
nor U3854 (N_3854,In_1223,In_1511);
nor U3855 (N_3855,In_518,In_1954);
nor U3856 (N_3856,In_2253,In_187);
nor U3857 (N_3857,In_1857,In_1170);
nor U3858 (N_3858,In_629,In_1812);
nand U3859 (N_3859,In_243,In_76);
nor U3860 (N_3860,In_1814,In_245);
nor U3861 (N_3861,In_2028,In_1483);
or U3862 (N_3862,In_1476,In_559);
or U3863 (N_3863,In_1039,In_2106);
or U3864 (N_3864,In_1823,In_1396);
nand U3865 (N_3865,In_723,In_1661);
or U3866 (N_3866,In_203,In_1092);
and U3867 (N_3867,In_553,In_1383);
xnor U3868 (N_3868,In_2041,In_2081);
or U3869 (N_3869,In_182,In_1179);
and U3870 (N_3870,In_401,In_2354);
and U3871 (N_3871,In_327,In_624);
nand U3872 (N_3872,In_1412,In_604);
xor U3873 (N_3873,In_2247,In_1591);
and U3874 (N_3874,In_1109,In_1425);
nor U3875 (N_3875,In_1849,In_449);
xnor U3876 (N_3876,In_1410,In_1425);
nor U3877 (N_3877,In_835,In_1828);
or U3878 (N_3878,In_2270,In_1185);
or U3879 (N_3879,In_1305,In_1815);
xnor U3880 (N_3880,In_2116,In_130);
or U3881 (N_3881,In_745,In_239);
and U3882 (N_3882,In_904,In_1211);
xor U3883 (N_3883,In_1856,In_994);
or U3884 (N_3884,In_182,In_1607);
nor U3885 (N_3885,In_5,In_1356);
nor U3886 (N_3886,In_1601,In_29);
and U3887 (N_3887,In_558,In_2462);
xnor U3888 (N_3888,In_1025,In_1468);
xnor U3889 (N_3889,In_2397,In_2208);
nor U3890 (N_3890,In_212,In_937);
nand U3891 (N_3891,In_1872,In_740);
nand U3892 (N_3892,In_1256,In_2072);
nor U3893 (N_3893,In_298,In_816);
nor U3894 (N_3894,In_2088,In_113);
nand U3895 (N_3895,In_2363,In_1803);
or U3896 (N_3896,In_1287,In_1226);
xor U3897 (N_3897,In_1672,In_1764);
nand U3898 (N_3898,In_602,In_848);
xnor U3899 (N_3899,In_1983,In_1842);
nor U3900 (N_3900,In_1222,In_1243);
or U3901 (N_3901,In_1299,In_47);
nor U3902 (N_3902,In_2068,In_26);
nor U3903 (N_3903,In_1397,In_853);
xor U3904 (N_3904,In_2154,In_1768);
nand U3905 (N_3905,In_181,In_492);
xnor U3906 (N_3906,In_2180,In_1504);
xnor U3907 (N_3907,In_1940,In_1031);
and U3908 (N_3908,In_2169,In_2366);
and U3909 (N_3909,In_1345,In_1493);
nor U3910 (N_3910,In_1793,In_2039);
nor U3911 (N_3911,In_1242,In_217);
nand U3912 (N_3912,In_365,In_760);
nor U3913 (N_3913,In_744,In_725);
nor U3914 (N_3914,In_402,In_1394);
or U3915 (N_3915,In_2027,In_1405);
nor U3916 (N_3916,In_904,In_2246);
nand U3917 (N_3917,In_467,In_49);
or U3918 (N_3918,In_1673,In_131);
or U3919 (N_3919,In_2259,In_464);
nand U3920 (N_3920,In_608,In_1231);
or U3921 (N_3921,In_252,In_2465);
and U3922 (N_3922,In_160,In_1153);
nand U3923 (N_3923,In_1673,In_1581);
and U3924 (N_3924,In_653,In_445);
xor U3925 (N_3925,In_960,In_469);
xor U3926 (N_3926,In_2376,In_1635);
or U3927 (N_3927,In_1109,In_2301);
nand U3928 (N_3928,In_674,In_1608);
nor U3929 (N_3929,In_2017,In_442);
nor U3930 (N_3930,In_971,In_1861);
nor U3931 (N_3931,In_2164,In_314);
nand U3932 (N_3932,In_1795,In_1085);
or U3933 (N_3933,In_1680,In_2365);
and U3934 (N_3934,In_707,In_1942);
xnor U3935 (N_3935,In_885,In_840);
nor U3936 (N_3936,In_435,In_579);
and U3937 (N_3937,In_568,In_1462);
or U3938 (N_3938,In_1811,In_286);
and U3939 (N_3939,In_332,In_73);
xor U3940 (N_3940,In_842,In_1984);
and U3941 (N_3941,In_1178,In_2414);
and U3942 (N_3942,In_2490,In_1308);
and U3943 (N_3943,In_213,In_968);
nor U3944 (N_3944,In_2460,In_618);
nand U3945 (N_3945,In_615,In_201);
xnor U3946 (N_3946,In_757,In_2423);
nand U3947 (N_3947,In_838,In_1839);
or U3948 (N_3948,In_1802,In_1115);
or U3949 (N_3949,In_882,In_2267);
nand U3950 (N_3950,In_1950,In_38);
nor U3951 (N_3951,In_930,In_353);
nand U3952 (N_3952,In_2191,In_2097);
and U3953 (N_3953,In_1447,In_525);
and U3954 (N_3954,In_657,In_1803);
nor U3955 (N_3955,In_221,In_152);
and U3956 (N_3956,In_1576,In_680);
and U3957 (N_3957,In_795,In_1334);
nand U3958 (N_3958,In_2152,In_1402);
and U3959 (N_3959,In_1830,In_57);
or U3960 (N_3960,In_419,In_2458);
nor U3961 (N_3961,In_533,In_788);
or U3962 (N_3962,In_29,In_2395);
nand U3963 (N_3963,In_605,In_2281);
xnor U3964 (N_3964,In_2058,In_1622);
or U3965 (N_3965,In_2310,In_2473);
or U3966 (N_3966,In_2182,In_167);
nand U3967 (N_3967,In_1169,In_890);
nor U3968 (N_3968,In_1525,In_1407);
and U3969 (N_3969,In_1753,In_943);
or U3970 (N_3970,In_2445,In_447);
or U3971 (N_3971,In_2386,In_440);
xnor U3972 (N_3972,In_505,In_2081);
xor U3973 (N_3973,In_1395,In_638);
and U3974 (N_3974,In_564,In_678);
and U3975 (N_3975,In_809,In_2363);
or U3976 (N_3976,In_845,In_1165);
xnor U3977 (N_3977,In_1664,In_1183);
and U3978 (N_3978,In_610,In_2050);
nand U3979 (N_3979,In_1445,In_1400);
or U3980 (N_3980,In_524,In_1992);
and U3981 (N_3981,In_1526,In_1655);
nand U3982 (N_3982,In_561,In_2205);
nor U3983 (N_3983,In_125,In_745);
and U3984 (N_3984,In_2459,In_2272);
nand U3985 (N_3985,In_272,In_1408);
and U3986 (N_3986,In_2381,In_336);
nor U3987 (N_3987,In_909,In_829);
xor U3988 (N_3988,In_764,In_1422);
or U3989 (N_3989,In_1531,In_1398);
nand U3990 (N_3990,In_2071,In_1246);
nand U3991 (N_3991,In_2015,In_2281);
and U3992 (N_3992,In_368,In_915);
nor U3993 (N_3993,In_2188,In_4);
xnor U3994 (N_3994,In_2400,In_111);
xor U3995 (N_3995,In_977,In_445);
and U3996 (N_3996,In_2192,In_91);
and U3997 (N_3997,In_15,In_380);
xor U3998 (N_3998,In_1389,In_2290);
nor U3999 (N_3999,In_18,In_487);
nand U4000 (N_4000,In_657,In_1716);
nand U4001 (N_4001,In_2135,In_59);
and U4002 (N_4002,In_90,In_2359);
or U4003 (N_4003,In_2188,In_2492);
or U4004 (N_4004,In_1537,In_164);
and U4005 (N_4005,In_1705,In_1347);
and U4006 (N_4006,In_2239,In_1800);
nand U4007 (N_4007,In_1387,In_1576);
or U4008 (N_4008,In_2144,In_1693);
xor U4009 (N_4009,In_2285,In_656);
nand U4010 (N_4010,In_1466,In_1508);
and U4011 (N_4011,In_2195,In_1029);
xor U4012 (N_4012,In_231,In_1545);
nor U4013 (N_4013,In_772,In_81);
nor U4014 (N_4014,In_1415,In_2477);
and U4015 (N_4015,In_161,In_314);
xnor U4016 (N_4016,In_1982,In_877);
nand U4017 (N_4017,In_2435,In_1386);
and U4018 (N_4018,In_1973,In_1662);
xnor U4019 (N_4019,In_1749,In_904);
nand U4020 (N_4020,In_662,In_148);
and U4021 (N_4021,In_1884,In_279);
and U4022 (N_4022,In_2497,In_344);
xnor U4023 (N_4023,In_2205,In_384);
and U4024 (N_4024,In_434,In_2401);
nand U4025 (N_4025,In_2319,In_1732);
xor U4026 (N_4026,In_926,In_172);
nand U4027 (N_4027,In_2030,In_296);
nand U4028 (N_4028,In_1731,In_2266);
nand U4029 (N_4029,In_2453,In_536);
nor U4030 (N_4030,In_704,In_1106);
or U4031 (N_4031,In_2171,In_1985);
xnor U4032 (N_4032,In_1329,In_1699);
nand U4033 (N_4033,In_1541,In_1941);
nor U4034 (N_4034,In_812,In_748);
and U4035 (N_4035,In_1847,In_1685);
or U4036 (N_4036,In_1519,In_1852);
or U4037 (N_4037,In_1371,In_796);
nand U4038 (N_4038,In_1455,In_1648);
nor U4039 (N_4039,In_398,In_1617);
or U4040 (N_4040,In_1853,In_2150);
or U4041 (N_4041,In_493,In_1293);
xor U4042 (N_4042,In_1853,In_1655);
or U4043 (N_4043,In_104,In_810);
xor U4044 (N_4044,In_2417,In_1137);
nand U4045 (N_4045,In_73,In_1120);
nor U4046 (N_4046,In_159,In_877);
xnor U4047 (N_4047,In_1337,In_247);
and U4048 (N_4048,In_2366,In_2371);
and U4049 (N_4049,In_1505,In_331);
nand U4050 (N_4050,In_2025,In_29);
and U4051 (N_4051,In_551,In_1093);
or U4052 (N_4052,In_2003,In_1302);
xor U4053 (N_4053,In_163,In_323);
nor U4054 (N_4054,In_347,In_2400);
nand U4055 (N_4055,In_1236,In_1999);
or U4056 (N_4056,In_63,In_1697);
nor U4057 (N_4057,In_474,In_1109);
or U4058 (N_4058,In_2237,In_1620);
and U4059 (N_4059,In_698,In_674);
xor U4060 (N_4060,In_1,In_2354);
nand U4061 (N_4061,In_25,In_1883);
xnor U4062 (N_4062,In_1243,In_1958);
nand U4063 (N_4063,In_2218,In_1818);
and U4064 (N_4064,In_786,In_1386);
or U4065 (N_4065,In_2317,In_1989);
or U4066 (N_4066,In_1253,In_1277);
and U4067 (N_4067,In_264,In_62);
nor U4068 (N_4068,In_1580,In_1756);
xor U4069 (N_4069,In_1094,In_1839);
or U4070 (N_4070,In_393,In_1747);
or U4071 (N_4071,In_464,In_1321);
nand U4072 (N_4072,In_496,In_1148);
xnor U4073 (N_4073,In_1839,In_1124);
and U4074 (N_4074,In_45,In_2298);
nor U4075 (N_4075,In_1927,In_1264);
xor U4076 (N_4076,In_2066,In_2227);
and U4077 (N_4077,In_1354,In_1115);
and U4078 (N_4078,In_443,In_1475);
xnor U4079 (N_4079,In_1342,In_821);
nor U4080 (N_4080,In_2200,In_380);
or U4081 (N_4081,In_732,In_2041);
and U4082 (N_4082,In_721,In_2404);
and U4083 (N_4083,In_2424,In_2364);
and U4084 (N_4084,In_2276,In_1189);
nor U4085 (N_4085,In_1218,In_231);
and U4086 (N_4086,In_893,In_158);
xnor U4087 (N_4087,In_780,In_2247);
nand U4088 (N_4088,In_317,In_2481);
or U4089 (N_4089,In_874,In_2041);
nor U4090 (N_4090,In_1855,In_624);
nor U4091 (N_4091,In_482,In_1723);
or U4092 (N_4092,In_2321,In_726);
xnor U4093 (N_4093,In_1219,In_1456);
nor U4094 (N_4094,In_1296,In_379);
xnor U4095 (N_4095,In_1600,In_2436);
nor U4096 (N_4096,In_323,In_2016);
and U4097 (N_4097,In_1679,In_1393);
and U4098 (N_4098,In_823,In_2278);
nor U4099 (N_4099,In_361,In_1994);
or U4100 (N_4100,In_1340,In_904);
or U4101 (N_4101,In_1148,In_2131);
and U4102 (N_4102,In_2445,In_1064);
or U4103 (N_4103,In_436,In_879);
xor U4104 (N_4104,In_1944,In_229);
nor U4105 (N_4105,In_2485,In_1383);
xnor U4106 (N_4106,In_1362,In_2442);
or U4107 (N_4107,In_2367,In_2106);
xnor U4108 (N_4108,In_1286,In_327);
xnor U4109 (N_4109,In_663,In_415);
nor U4110 (N_4110,In_1233,In_2336);
nand U4111 (N_4111,In_342,In_2356);
nand U4112 (N_4112,In_1318,In_2455);
nand U4113 (N_4113,In_2278,In_1810);
nand U4114 (N_4114,In_1038,In_2077);
xor U4115 (N_4115,In_2295,In_35);
and U4116 (N_4116,In_1022,In_1195);
and U4117 (N_4117,In_2094,In_1973);
xnor U4118 (N_4118,In_1142,In_1126);
and U4119 (N_4119,In_1320,In_2375);
and U4120 (N_4120,In_2239,In_252);
xor U4121 (N_4121,In_843,In_107);
nand U4122 (N_4122,In_1909,In_664);
nand U4123 (N_4123,In_712,In_1317);
nor U4124 (N_4124,In_2122,In_2496);
nor U4125 (N_4125,In_95,In_304);
xor U4126 (N_4126,In_556,In_685);
xor U4127 (N_4127,In_2231,In_32);
xnor U4128 (N_4128,In_775,In_2210);
or U4129 (N_4129,In_1486,In_1037);
or U4130 (N_4130,In_1788,In_1341);
or U4131 (N_4131,In_2177,In_808);
xnor U4132 (N_4132,In_2023,In_531);
or U4133 (N_4133,In_1695,In_885);
nor U4134 (N_4134,In_1115,In_1319);
nand U4135 (N_4135,In_749,In_1688);
nand U4136 (N_4136,In_1174,In_261);
nand U4137 (N_4137,In_1523,In_870);
and U4138 (N_4138,In_2173,In_184);
or U4139 (N_4139,In_715,In_2309);
nand U4140 (N_4140,In_335,In_2133);
and U4141 (N_4141,In_2131,In_457);
or U4142 (N_4142,In_1626,In_2289);
and U4143 (N_4143,In_1700,In_1542);
nand U4144 (N_4144,In_1834,In_1054);
or U4145 (N_4145,In_96,In_1251);
or U4146 (N_4146,In_1057,In_2192);
nand U4147 (N_4147,In_468,In_453);
or U4148 (N_4148,In_1373,In_1333);
nor U4149 (N_4149,In_325,In_1768);
and U4150 (N_4150,In_2050,In_824);
and U4151 (N_4151,In_167,In_2354);
and U4152 (N_4152,In_617,In_1467);
or U4153 (N_4153,In_173,In_2389);
nor U4154 (N_4154,In_2226,In_1542);
nor U4155 (N_4155,In_2422,In_1370);
xor U4156 (N_4156,In_1026,In_1252);
xor U4157 (N_4157,In_2086,In_2438);
or U4158 (N_4158,In_2151,In_1375);
and U4159 (N_4159,In_1536,In_1922);
xnor U4160 (N_4160,In_2139,In_249);
or U4161 (N_4161,In_1454,In_1737);
nor U4162 (N_4162,In_515,In_1980);
xnor U4163 (N_4163,In_2267,In_1727);
xnor U4164 (N_4164,In_1346,In_1322);
nand U4165 (N_4165,In_432,In_192);
or U4166 (N_4166,In_1988,In_2244);
nand U4167 (N_4167,In_1442,In_1680);
xnor U4168 (N_4168,In_405,In_483);
or U4169 (N_4169,In_916,In_1298);
nor U4170 (N_4170,In_596,In_1843);
xnor U4171 (N_4171,In_420,In_885);
and U4172 (N_4172,In_1233,In_1348);
nor U4173 (N_4173,In_1536,In_1559);
or U4174 (N_4174,In_151,In_1240);
nor U4175 (N_4175,In_1992,In_2409);
nor U4176 (N_4176,In_2016,In_1529);
nand U4177 (N_4177,In_2023,In_2252);
xor U4178 (N_4178,In_1847,In_1865);
and U4179 (N_4179,In_948,In_244);
nand U4180 (N_4180,In_522,In_1833);
nor U4181 (N_4181,In_1090,In_561);
nand U4182 (N_4182,In_1164,In_25);
nor U4183 (N_4183,In_1041,In_2216);
or U4184 (N_4184,In_2481,In_2080);
nand U4185 (N_4185,In_643,In_473);
or U4186 (N_4186,In_2444,In_2006);
nand U4187 (N_4187,In_1516,In_2233);
nor U4188 (N_4188,In_1777,In_925);
xnor U4189 (N_4189,In_2120,In_1945);
and U4190 (N_4190,In_837,In_1249);
nor U4191 (N_4191,In_793,In_1984);
nor U4192 (N_4192,In_1938,In_43);
and U4193 (N_4193,In_945,In_1501);
xnor U4194 (N_4194,In_188,In_2019);
nor U4195 (N_4195,In_878,In_1768);
xnor U4196 (N_4196,In_6,In_873);
nand U4197 (N_4197,In_536,In_1069);
and U4198 (N_4198,In_2183,In_1683);
nand U4199 (N_4199,In_2144,In_2059);
xor U4200 (N_4200,In_997,In_689);
or U4201 (N_4201,In_1661,In_1653);
or U4202 (N_4202,In_1957,In_1612);
and U4203 (N_4203,In_1379,In_2284);
nor U4204 (N_4204,In_2190,In_2249);
nand U4205 (N_4205,In_649,In_2355);
nor U4206 (N_4206,In_684,In_208);
nand U4207 (N_4207,In_122,In_1832);
or U4208 (N_4208,In_2132,In_2401);
or U4209 (N_4209,In_338,In_1470);
xnor U4210 (N_4210,In_1783,In_2298);
xnor U4211 (N_4211,In_1440,In_1802);
and U4212 (N_4212,In_2029,In_937);
nor U4213 (N_4213,In_1788,In_2427);
nor U4214 (N_4214,In_289,In_642);
or U4215 (N_4215,In_1475,In_2052);
xnor U4216 (N_4216,In_44,In_1379);
xnor U4217 (N_4217,In_202,In_2090);
xnor U4218 (N_4218,In_1874,In_2229);
or U4219 (N_4219,In_20,In_292);
nor U4220 (N_4220,In_1650,In_867);
nor U4221 (N_4221,In_1200,In_2217);
nand U4222 (N_4222,In_1602,In_442);
nor U4223 (N_4223,In_206,In_201);
or U4224 (N_4224,In_1508,In_1008);
nand U4225 (N_4225,In_74,In_2185);
xor U4226 (N_4226,In_1290,In_1452);
and U4227 (N_4227,In_959,In_588);
nand U4228 (N_4228,In_484,In_1107);
nor U4229 (N_4229,In_313,In_714);
and U4230 (N_4230,In_894,In_35);
and U4231 (N_4231,In_282,In_1311);
nand U4232 (N_4232,In_223,In_1012);
xnor U4233 (N_4233,In_1479,In_78);
nor U4234 (N_4234,In_906,In_2082);
nor U4235 (N_4235,In_1846,In_791);
nor U4236 (N_4236,In_307,In_1939);
nor U4237 (N_4237,In_1760,In_190);
nor U4238 (N_4238,In_1031,In_1011);
or U4239 (N_4239,In_2208,In_2244);
nand U4240 (N_4240,In_1916,In_2474);
nand U4241 (N_4241,In_429,In_866);
and U4242 (N_4242,In_1276,In_1162);
or U4243 (N_4243,In_2405,In_1787);
or U4244 (N_4244,In_1363,In_1764);
and U4245 (N_4245,In_1387,In_2147);
and U4246 (N_4246,In_897,In_2459);
xnor U4247 (N_4247,In_297,In_1425);
nor U4248 (N_4248,In_1687,In_1751);
nor U4249 (N_4249,In_907,In_1846);
xor U4250 (N_4250,In_674,In_1394);
nor U4251 (N_4251,In_496,In_814);
and U4252 (N_4252,In_1501,In_2120);
and U4253 (N_4253,In_473,In_1186);
nand U4254 (N_4254,In_446,In_1977);
nor U4255 (N_4255,In_769,In_471);
nor U4256 (N_4256,In_2250,In_1675);
nand U4257 (N_4257,In_2076,In_1829);
and U4258 (N_4258,In_829,In_2137);
xor U4259 (N_4259,In_1356,In_1152);
nor U4260 (N_4260,In_1700,In_805);
xor U4261 (N_4261,In_106,In_416);
xor U4262 (N_4262,In_994,In_2427);
xor U4263 (N_4263,In_1105,In_534);
and U4264 (N_4264,In_466,In_676);
or U4265 (N_4265,In_364,In_2438);
nand U4266 (N_4266,In_175,In_2376);
xor U4267 (N_4267,In_2429,In_2424);
and U4268 (N_4268,In_1855,In_326);
nand U4269 (N_4269,In_1966,In_1901);
nand U4270 (N_4270,In_1414,In_346);
or U4271 (N_4271,In_2325,In_977);
xor U4272 (N_4272,In_1133,In_2193);
nand U4273 (N_4273,In_127,In_1043);
nand U4274 (N_4274,In_615,In_2);
or U4275 (N_4275,In_2373,In_710);
or U4276 (N_4276,In_26,In_1829);
nor U4277 (N_4277,In_1992,In_1201);
or U4278 (N_4278,In_673,In_2086);
nor U4279 (N_4279,In_136,In_694);
nor U4280 (N_4280,In_1567,In_2166);
nand U4281 (N_4281,In_301,In_1876);
nand U4282 (N_4282,In_1580,In_1117);
and U4283 (N_4283,In_506,In_1749);
and U4284 (N_4284,In_2221,In_2003);
xor U4285 (N_4285,In_2279,In_1280);
nor U4286 (N_4286,In_1691,In_36);
nor U4287 (N_4287,In_532,In_1613);
nor U4288 (N_4288,In_1386,In_1143);
nand U4289 (N_4289,In_1551,In_308);
xnor U4290 (N_4290,In_1029,In_853);
or U4291 (N_4291,In_477,In_2382);
xnor U4292 (N_4292,In_2465,In_484);
and U4293 (N_4293,In_970,In_315);
or U4294 (N_4294,In_1078,In_1361);
xor U4295 (N_4295,In_45,In_700);
nor U4296 (N_4296,In_517,In_253);
or U4297 (N_4297,In_2287,In_1801);
and U4298 (N_4298,In_2143,In_1365);
and U4299 (N_4299,In_944,In_674);
nor U4300 (N_4300,In_1315,In_413);
nor U4301 (N_4301,In_2001,In_193);
and U4302 (N_4302,In_1742,In_1768);
and U4303 (N_4303,In_1908,In_2243);
and U4304 (N_4304,In_1486,In_1673);
xnor U4305 (N_4305,In_998,In_1991);
nand U4306 (N_4306,In_1536,In_2434);
nand U4307 (N_4307,In_408,In_371);
xor U4308 (N_4308,In_1715,In_628);
or U4309 (N_4309,In_1818,In_1170);
and U4310 (N_4310,In_1310,In_1663);
or U4311 (N_4311,In_182,In_606);
nand U4312 (N_4312,In_992,In_1002);
nand U4313 (N_4313,In_1188,In_2033);
xor U4314 (N_4314,In_133,In_275);
nor U4315 (N_4315,In_1758,In_1226);
or U4316 (N_4316,In_1550,In_256);
nor U4317 (N_4317,In_466,In_2247);
or U4318 (N_4318,In_588,In_2095);
and U4319 (N_4319,In_263,In_438);
or U4320 (N_4320,In_56,In_288);
or U4321 (N_4321,In_167,In_867);
and U4322 (N_4322,In_1160,In_853);
nand U4323 (N_4323,In_2357,In_1820);
or U4324 (N_4324,In_991,In_2141);
xor U4325 (N_4325,In_804,In_1696);
nor U4326 (N_4326,In_435,In_915);
nand U4327 (N_4327,In_297,In_2229);
or U4328 (N_4328,In_1039,In_1229);
xor U4329 (N_4329,In_1974,In_1953);
nor U4330 (N_4330,In_179,In_1919);
nor U4331 (N_4331,In_2455,In_1095);
nand U4332 (N_4332,In_328,In_599);
and U4333 (N_4333,In_1548,In_1713);
nand U4334 (N_4334,In_2105,In_455);
nor U4335 (N_4335,In_1562,In_2286);
and U4336 (N_4336,In_2068,In_685);
nor U4337 (N_4337,In_2452,In_2461);
xnor U4338 (N_4338,In_83,In_1904);
nand U4339 (N_4339,In_373,In_2178);
nand U4340 (N_4340,In_759,In_702);
nor U4341 (N_4341,In_1784,In_82);
and U4342 (N_4342,In_900,In_400);
or U4343 (N_4343,In_1558,In_1060);
and U4344 (N_4344,In_958,In_486);
and U4345 (N_4345,In_653,In_263);
nand U4346 (N_4346,In_999,In_1862);
and U4347 (N_4347,In_379,In_1395);
nand U4348 (N_4348,In_2384,In_734);
xnor U4349 (N_4349,In_366,In_40);
nand U4350 (N_4350,In_2456,In_1580);
and U4351 (N_4351,In_174,In_1597);
nand U4352 (N_4352,In_578,In_2116);
xnor U4353 (N_4353,In_1466,In_310);
nor U4354 (N_4354,In_11,In_257);
nor U4355 (N_4355,In_1962,In_1992);
xor U4356 (N_4356,In_570,In_1613);
nand U4357 (N_4357,In_2440,In_732);
nand U4358 (N_4358,In_1555,In_1624);
and U4359 (N_4359,In_228,In_584);
and U4360 (N_4360,In_856,In_972);
nand U4361 (N_4361,In_308,In_2236);
nand U4362 (N_4362,In_2084,In_350);
or U4363 (N_4363,In_279,In_719);
nand U4364 (N_4364,In_356,In_1304);
nor U4365 (N_4365,In_1648,In_502);
nand U4366 (N_4366,In_2040,In_1863);
xor U4367 (N_4367,In_753,In_1789);
and U4368 (N_4368,In_612,In_517);
or U4369 (N_4369,In_445,In_123);
xor U4370 (N_4370,In_199,In_1156);
and U4371 (N_4371,In_504,In_1930);
xnor U4372 (N_4372,In_111,In_1351);
or U4373 (N_4373,In_510,In_1573);
or U4374 (N_4374,In_841,In_743);
nand U4375 (N_4375,In_966,In_1331);
nor U4376 (N_4376,In_1571,In_1935);
or U4377 (N_4377,In_1042,In_97);
xnor U4378 (N_4378,In_574,In_1341);
or U4379 (N_4379,In_624,In_2267);
nand U4380 (N_4380,In_2276,In_2054);
xnor U4381 (N_4381,In_65,In_2070);
or U4382 (N_4382,In_680,In_2440);
or U4383 (N_4383,In_420,In_942);
nor U4384 (N_4384,In_218,In_1533);
and U4385 (N_4385,In_2221,In_1336);
xor U4386 (N_4386,In_1892,In_1251);
or U4387 (N_4387,In_1764,In_918);
xnor U4388 (N_4388,In_218,In_2252);
and U4389 (N_4389,In_2489,In_2418);
or U4390 (N_4390,In_121,In_2135);
and U4391 (N_4391,In_1480,In_1284);
nand U4392 (N_4392,In_243,In_1895);
xor U4393 (N_4393,In_241,In_1968);
and U4394 (N_4394,In_2023,In_2126);
or U4395 (N_4395,In_2056,In_1862);
and U4396 (N_4396,In_376,In_280);
and U4397 (N_4397,In_2145,In_1619);
or U4398 (N_4398,In_2499,In_2333);
xor U4399 (N_4399,In_1717,In_2227);
or U4400 (N_4400,In_743,In_1594);
or U4401 (N_4401,In_2195,In_1329);
nor U4402 (N_4402,In_1104,In_493);
and U4403 (N_4403,In_2054,In_457);
xor U4404 (N_4404,In_986,In_1514);
nand U4405 (N_4405,In_2301,In_674);
and U4406 (N_4406,In_1907,In_534);
xor U4407 (N_4407,In_379,In_1717);
xnor U4408 (N_4408,In_516,In_1670);
and U4409 (N_4409,In_323,In_1542);
or U4410 (N_4410,In_999,In_1455);
xor U4411 (N_4411,In_527,In_516);
xor U4412 (N_4412,In_2195,In_325);
or U4413 (N_4413,In_1042,In_2464);
xnor U4414 (N_4414,In_998,In_1807);
nand U4415 (N_4415,In_2082,In_450);
nor U4416 (N_4416,In_1869,In_1561);
or U4417 (N_4417,In_1916,In_2405);
or U4418 (N_4418,In_822,In_442);
nand U4419 (N_4419,In_861,In_1251);
nand U4420 (N_4420,In_971,In_353);
xnor U4421 (N_4421,In_21,In_2209);
nand U4422 (N_4422,In_1234,In_2162);
nand U4423 (N_4423,In_2398,In_615);
or U4424 (N_4424,In_2121,In_776);
or U4425 (N_4425,In_1791,In_991);
or U4426 (N_4426,In_444,In_1630);
nor U4427 (N_4427,In_2300,In_2262);
xor U4428 (N_4428,In_854,In_1784);
and U4429 (N_4429,In_2018,In_1193);
and U4430 (N_4430,In_741,In_404);
nand U4431 (N_4431,In_26,In_1836);
nand U4432 (N_4432,In_2064,In_1330);
nor U4433 (N_4433,In_520,In_1481);
nand U4434 (N_4434,In_173,In_1782);
nand U4435 (N_4435,In_55,In_571);
nand U4436 (N_4436,In_894,In_1642);
or U4437 (N_4437,In_2377,In_184);
xnor U4438 (N_4438,In_2015,In_719);
or U4439 (N_4439,In_1937,In_2111);
nand U4440 (N_4440,In_1976,In_387);
nand U4441 (N_4441,In_1882,In_696);
or U4442 (N_4442,In_130,In_340);
nand U4443 (N_4443,In_1255,In_1295);
nor U4444 (N_4444,In_630,In_1520);
nor U4445 (N_4445,In_2476,In_915);
xor U4446 (N_4446,In_962,In_548);
and U4447 (N_4447,In_564,In_1507);
and U4448 (N_4448,In_82,In_904);
and U4449 (N_4449,In_493,In_1618);
nand U4450 (N_4450,In_320,In_195);
nand U4451 (N_4451,In_1322,In_1787);
or U4452 (N_4452,In_2406,In_1613);
or U4453 (N_4453,In_2338,In_2352);
or U4454 (N_4454,In_1035,In_1738);
xnor U4455 (N_4455,In_2413,In_1979);
and U4456 (N_4456,In_798,In_402);
nor U4457 (N_4457,In_2289,In_2021);
or U4458 (N_4458,In_1765,In_1160);
and U4459 (N_4459,In_1332,In_1515);
or U4460 (N_4460,In_2226,In_264);
or U4461 (N_4461,In_2210,In_2146);
or U4462 (N_4462,In_740,In_2075);
nand U4463 (N_4463,In_1918,In_279);
or U4464 (N_4464,In_2480,In_1620);
or U4465 (N_4465,In_2256,In_1457);
and U4466 (N_4466,In_1834,In_874);
or U4467 (N_4467,In_2367,In_266);
or U4468 (N_4468,In_1728,In_1278);
xnor U4469 (N_4469,In_1482,In_1642);
or U4470 (N_4470,In_2136,In_2284);
and U4471 (N_4471,In_2373,In_523);
or U4472 (N_4472,In_422,In_1294);
or U4473 (N_4473,In_1662,In_331);
and U4474 (N_4474,In_20,In_827);
or U4475 (N_4475,In_583,In_1426);
nand U4476 (N_4476,In_2095,In_332);
nand U4477 (N_4477,In_164,In_924);
nor U4478 (N_4478,In_459,In_2165);
xnor U4479 (N_4479,In_228,In_2162);
nor U4480 (N_4480,In_422,In_525);
nand U4481 (N_4481,In_554,In_1601);
nand U4482 (N_4482,In_1275,In_783);
or U4483 (N_4483,In_1905,In_13);
and U4484 (N_4484,In_1070,In_1071);
xor U4485 (N_4485,In_2319,In_2138);
or U4486 (N_4486,In_1122,In_1135);
or U4487 (N_4487,In_1544,In_1462);
nand U4488 (N_4488,In_2257,In_2430);
nand U4489 (N_4489,In_1297,In_234);
or U4490 (N_4490,In_1834,In_132);
xor U4491 (N_4491,In_2245,In_540);
or U4492 (N_4492,In_1782,In_664);
and U4493 (N_4493,In_625,In_1170);
xor U4494 (N_4494,In_598,In_429);
nand U4495 (N_4495,In_561,In_596);
nor U4496 (N_4496,In_485,In_1192);
nand U4497 (N_4497,In_452,In_900);
nor U4498 (N_4498,In_1603,In_853);
and U4499 (N_4499,In_1869,In_1780);
and U4500 (N_4500,In_121,In_2325);
nor U4501 (N_4501,In_132,In_1271);
nand U4502 (N_4502,In_1203,In_1969);
xnor U4503 (N_4503,In_635,In_1514);
nor U4504 (N_4504,In_1050,In_1816);
or U4505 (N_4505,In_2222,In_2297);
nor U4506 (N_4506,In_646,In_1938);
xnor U4507 (N_4507,In_2347,In_2080);
xor U4508 (N_4508,In_1514,In_1407);
or U4509 (N_4509,In_954,In_2217);
nor U4510 (N_4510,In_838,In_1954);
nand U4511 (N_4511,In_1221,In_731);
and U4512 (N_4512,In_488,In_1197);
xnor U4513 (N_4513,In_1536,In_1891);
xnor U4514 (N_4514,In_2272,In_2305);
nand U4515 (N_4515,In_1769,In_110);
or U4516 (N_4516,In_277,In_1145);
nand U4517 (N_4517,In_618,In_521);
nand U4518 (N_4518,In_243,In_1709);
or U4519 (N_4519,In_858,In_2101);
nand U4520 (N_4520,In_1849,In_908);
and U4521 (N_4521,In_1989,In_1243);
and U4522 (N_4522,In_2320,In_577);
nor U4523 (N_4523,In_522,In_1350);
nand U4524 (N_4524,In_1265,In_1752);
and U4525 (N_4525,In_1182,In_1481);
or U4526 (N_4526,In_797,In_564);
or U4527 (N_4527,In_1667,In_492);
nand U4528 (N_4528,In_579,In_858);
nor U4529 (N_4529,In_1351,In_311);
or U4530 (N_4530,In_1613,In_1130);
xor U4531 (N_4531,In_2081,In_27);
or U4532 (N_4532,In_1751,In_2284);
or U4533 (N_4533,In_27,In_1180);
or U4534 (N_4534,In_2232,In_358);
nor U4535 (N_4535,In_389,In_436);
nor U4536 (N_4536,In_734,In_1577);
and U4537 (N_4537,In_1761,In_660);
nor U4538 (N_4538,In_1169,In_95);
nand U4539 (N_4539,In_1651,In_2307);
xor U4540 (N_4540,In_732,In_110);
nand U4541 (N_4541,In_2229,In_1205);
or U4542 (N_4542,In_2382,In_626);
and U4543 (N_4543,In_588,In_2205);
xor U4544 (N_4544,In_1302,In_419);
and U4545 (N_4545,In_645,In_147);
nor U4546 (N_4546,In_1962,In_1660);
or U4547 (N_4547,In_2136,In_2370);
xnor U4548 (N_4548,In_813,In_2361);
xnor U4549 (N_4549,In_997,In_2461);
nand U4550 (N_4550,In_142,In_1562);
nor U4551 (N_4551,In_1190,In_1255);
and U4552 (N_4552,In_627,In_2223);
and U4553 (N_4553,In_1578,In_2063);
nand U4554 (N_4554,In_991,In_1460);
nor U4555 (N_4555,In_1376,In_1882);
xor U4556 (N_4556,In_387,In_2357);
xnor U4557 (N_4557,In_2196,In_807);
xnor U4558 (N_4558,In_1123,In_336);
nor U4559 (N_4559,In_1452,In_638);
and U4560 (N_4560,In_1749,In_1658);
nand U4561 (N_4561,In_2346,In_1639);
nor U4562 (N_4562,In_1979,In_551);
nand U4563 (N_4563,In_645,In_1962);
nor U4564 (N_4564,In_1281,In_527);
nand U4565 (N_4565,In_1584,In_1305);
and U4566 (N_4566,In_346,In_686);
or U4567 (N_4567,In_956,In_1279);
xnor U4568 (N_4568,In_1952,In_1285);
nor U4569 (N_4569,In_315,In_2228);
and U4570 (N_4570,In_1103,In_450);
or U4571 (N_4571,In_1804,In_790);
and U4572 (N_4572,In_2348,In_1563);
and U4573 (N_4573,In_1018,In_825);
or U4574 (N_4574,In_750,In_1509);
nand U4575 (N_4575,In_191,In_676);
xnor U4576 (N_4576,In_1804,In_1800);
xnor U4577 (N_4577,In_1277,In_1299);
nand U4578 (N_4578,In_322,In_140);
and U4579 (N_4579,In_130,In_1058);
or U4580 (N_4580,In_97,In_2147);
or U4581 (N_4581,In_48,In_2355);
nand U4582 (N_4582,In_1060,In_1555);
or U4583 (N_4583,In_1843,In_2211);
xor U4584 (N_4584,In_754,In_2171);
or U4585 (N_4585,In_307,In_939);
and U4586 (N_4586,In_1907,In_1326);
nor U4587 (N_4587,In_2450,In_2083);
xor U4588 (N_4588,In_482,In_2164);
or U4589 (N_4589,In_1943,In_1787);
nand U4590 (N_4590,In_1638,In_1969);
nand U4591 (N_4591,In_1202,In_1506);
or U4592 (N_4592,In_2115,In_1964);
nand U4593 (N_4593,In_2157,In_2000);
or U4594 (N_4594,In_1850,In_1537);
nand U4595 (N_4595,In_690,In_362);
nor U4596 (N_4596,In_62,In_1529);
nand U4597 (N_4597,In_822,In_1944);
nand U4598 (N_4598,In_2120,In_2273);
or U4599 (N_4599,In_801,In_1634);
xnor U4600 (N_4600,In_1086,In_1062);
and U4601 (N_4601,In_159,In_1225);
nand U4602 (N_4602,In_1245,In_761);
xnor U4603 (N_4603,In_61,In_2330);
and U4604 (N_4604,In_1349,In_2234);
or U4605 (N_4605,In_1869,In_1711);
and U4606 (N_4606,In_2454,In_922);
nand U4607 (N_4607,In_1145,In_876);
xor U4608 (N_4608,In_1788,In_329);
or U4609 (N_4609,In_2326,In_152);
nand U4610 (N_4610,In_853,In_1797);
nand U4611 (N_4611,In_1885,In_1729);
nor U4612 (N_4612,In_2382,In_81);
nor U4613 (N_4613,In_2036,In_1959);
and U4614 (N_4614,In_2136,In_2301);
and U4615 (N_4615,In_883,In_604);
nand U4616 (N_4616,In_1257,In_2494);
xor U4617 (N_4617,In_2170,In_847);
or U4618 (N_4618,In_311,In_2033);
or U4619 (N_4619,In_1757,In_2424);
nand U4620 (N_4620,In_343,In_2221);
or U4621 (N_4621,In_735,In_82);
xnor U4622 (N_4622,In_2326,In_979);
or U4623 (N_4623,In_740,In_1950);
nor U4624 (N_4624,In_1590,In_717);
nand U4625 (N_4625,In_761,In_2201);
nor U4626 (N_4626,In_975,In_2152);
or U4627 (N_4627,In_2221,In_226);
and U4628 (N_4628,In_2330,In_761);
xnor U4629 (N_4629,In_317,In_1343);
nor U4630 (N_4630,In_261,In_170);
nor U4631 (N_4631,In_107,In_2188);
xnor U4632 (N_4632,In_1886,In_1470);
and U4633 (N_4633,In_2281,In_480);
or U4634 (N_4634,In_2438,In_580);
and U4635 (N_4635,In_541,In_2083);
nand U4636 (N_4636,In_812,In_1383);
nand U4637 (N_4637,In_1098,In_128);
nand U4638 (N_4638,In_298,In_2395);
xnor U4639 (N_4639,In_669,In_481);
and U4640 (N_4640,In_1324,In_1402);
nand U4641 (N_4641,In_2435,In_1349);
or U4642 (N_4642,In_879,In_675);
or U4643 (N_4643,In_2250,In_537);
or U4644 (N_4644,In_441,In_573);
or U4645 (N_4645,In_2183,In_565);
nand U4646 (N_4646,In_848,In_691);
nor U4647 (N_4647,In_2342,In_1380);
and U4648 (N_4648,In_22,In_1112);
xnor U4649 (N_4649,In_1421,In_53);
nand U4650 (N_4650,In_2262,In_1390);
xor U4651 (N_4651,In_92,In_723);
or U4652 (N_4652,In_1279,In_2003);
nor U4653 (N_4653,In_27,In_82);
or U4654 (N_4654,In_320,In_2408);
or U4655 (N_4655,In_1322,In_1386);
or U4656 (N_4656,In_1727,In_766);
and U4657 (N_4657,In_1351,In_2209);
xor U4658 (N_4658,In_1627,In_2177);
nand U4659 (N_4659,In_812,In_1092);
or U4660 (N_4660,In_305,In_1308);
xor U4661 (N_4661,In_73,In_1791);
xnor U4662 (N_4662,In_44,In_266);
xnor U4663 (N_4663,In_899,In_1326);
and U4664 (N_4664,In_723,In_829);
and U4665 (N_4665,In_766,In_824);
nor U4666 (N_4666,In_1592,In_1132);
nand U4667 (N_4667,In_416,In_453);
xor U4668 (N_4668,In_393,In_2487);
and U4669 (N_4669,In_308,In_2482);
and U4670 (N_4670,In_1208,In_811);
xnor U4671 (N_4671,In_288,In_2070);
nor U4672 (N_4672,In_2049,In_654);
and U4673 (N_4673,In_357,In_21);
and U4674 (N_4674,In_1024,In_1069);
and U4675 (N_4675,In_1087,In_1003);
nand U4676 (N_4676,In_274,In_732);
nand U4677 (N_4677,In_65,In_2023);
or U4678 (N_4678,In_2073,In_1391);
nor U4679 (N_4679,In_1666,In_883);
nand U4680 (N_4680,In_2048,In_1616);
nand U4681 (N_4681,In_543,In_1070);
nor U4682 (N_4682,In_1692,In_122);
xor U4683 (N_4683,In_1540,In_1356);
or U4684 (N_4684,In_1077,In_405);
and U4685 (N_4685,In_2014,In_2113);
nand U4686 (N_4686,In_1301,In_1945);
and U4687 (N_4687,In_95,In_2224);
xnor U4688 (N_4688,In_2474,In_1184);
or U4689 (N_4689,In_1916,In_1404);
or U4690 (N_4690,In_2089,In_662);
and U4691 (N_4691,In_542,In_598);
nand U4692 (N_4692,In_2332,In_2004);
nor U4693 (N_4693,In_932,In_2092);
nor U4694 (N_4694,In_1660,In_353);
xor U4695 (N_4695,In_2158,In_1321);
nor U4696 (N_4696,In_125,In_553);
xnor U4697 (N_4697,In_499,In_1144);
nand U4698 (N_4698,In_831,In_2436);
xor U4699 (N_4699,In_2209,In_2028);
nand U4700 (N_4700,In_2444,In_624);
and U4701 (N_4701,In_1881,In_19);
nor U4702 (N_4702,In_1252,In_1872);
nor U4703 (N_4703,In_1862,In_1252);
nor U4704 (N_4704,In_1370,In_684);
nand U4705 (N_4705,In_2479,In_582);
or U4706 (N_4706,In_253,In_2452);
and U4707 (N_4707,In_293,In_2202);
or U4708 (N_4708,In_1930,In_1171);
nor U4709 (N_4709,In_1269,In_931);
xor U4710 (N_4710,In_186,In_1206);
nor U4711 (N_4711,In_1251,In_1109);
or U4712 (N_4712,In_1435,In_2155);
or U4713 (N_4713,In_2381,In_1358);
and U4714 (N_4714,In_1573,In_988);
or U4715 (N_4715,In_1851,In_1191);
nand U4716 (N_4716,In_2094,In_1478);
nor U4717 (N_4717,In_1236,In_2229);
nor U4718 (N_4718,In_413,In_1384);
nand U4719 (N_4719,In_482,In_1847);
or U4720 (N_4720,In_136,In_1901);
and U4721 (N_4721,In_1414,In_1304);
or U4722 (N_4722,In_18,In_47);
and U4723 (N_4723,In_934,In_1656);
nor U4724 (N_4724,In_329,In_1786);
nand U4725 (N_4725,In_2112,In_1619);
and U4726 (N_4726,In_919,In_1263);
nor U4727 (N_4727,In_2230,In_1328);
nor U4728 (N_4728,In_2092,In_1696);
xor U4729 (N_4729,In_2384,In_588);
or U4730 (N_4730,In_1288,In_155);
nor U4731 (N_4731,In_695,In_1457);
nand U4732 (N_4732,In_1190,In_1015);
xor U4733 (N_4733,In_1509,In_2256);
nor U4734 (N_4734,In_2269,In_313);
or U4735 (N_4735,In_32,In_463);
and U4736 (N_4736,In_1677,In_194);
nand U4737 (N_4737,In_1867,In_583);
nand U4738 (N_4738,In_1059,In_1122);
and U4739 (N_4739,In_1161,In_2462);
nand U4740 (N_4740,In_1196,In_1984);
xnor U4741 (N_4741,In_2303,In_1987);
or U4742 (N_4742,In_1731,In_1808);
and U4743 (N_4743,In_541,In_1885);
xnor U4744 (N_4744,In_2339,In_1937);
or U4745 (N_4745,In_179,In_2420);
xnor U4746 (N_4746,In_1618,In_394);
nor U4747 (N_4747,In_192,In_582);
and U4748 (N_4748,In_1746,In_2309);
nor U4749 (N_4749,In_1142,In_1078);
or U4750 (N_4750,In_1538,In_1102);
or U4751 (N_4751,In_1480,In_1619);
xor U4752 (N_4752,In_2106,In_444);
xnor U4753 (N_4753,In_1419,In_760);
nor U4754 (N_4754,In_1040,In_1181);
xor U4755 (N_4755,In_749,In_1635);
nand U4756 (N_4756,In_56,In_1790);
nand U4757 (N_4757,In_1703,In_75);
nor U4758 (N_4758,In_431,In_1613);
nand U4759 (N_4759,In_1758,In_317);
and U4760 (N_4760,In_1116,In_1242);
and U4761 (N_4761,In_1655,In_1616);
nor U4762 (N_4762,In_2089,In_15);
or U4763 (N_4763,In_2022,In_2440);
and U4764 (N_4764,In_1409,In_765);
or U4765 (N_4765,In_302,In_1983);
xor U4766 (N_4766,In_1867,In_2347);
nand U4767 (N_4767,In_2168,In_665);
nand U4768 (N_4768,In_425,In_342);
xnor U4769 (N_4769,In_966,In_2385);
and U4770 (N_4770,In_839,In_2404);
nand U4771 (N_4771,In_866,In_779);
nand U4772 (N_4772,In_1741,In_1351);
or U4773 (N_4773,In_2136,In_1379);
or U4774 (N_4774,In_2350,In_1296);
and U4775 (N_4775,In_1440,In_585);
xor U4776 (N_4776,In_1636,In_1206);
nand U4777 (N_4777,In_46,In_1420);
xor U4778 (N_4778,In_1907,In_1484);
nand U4779 (N_4779,In_2313,In_944);
xnor U4780 (N_4780,In_1644,In_2078);
xor U4781 (N_4781,In_1642,In_1287);
nand U4782 (N_4782,In_2195,In_945);
and U4783 (N_4783,In_1067,In_309);
nor U4784 (N_4784,In_2191,In_1631);
xnor U4785 (N_4785,In_2177,In_1145);
nor U4786 (N_4786,In_860,In_1991);
xnor U4787 (N_4787,In_489,In_163);
or U4788 (N_4788,In_114,In_1432);
and U4789 (N_4789,In_268,In_1105);
xnor U4790 (N_4790,In_1051,In_1116);
nor U4791 (N_4791,In_861,In_79);
and U4792 (N_4792,In_1337,In_2448);
nand U4793 (N_4793,In_1442,In_1900);
nor U4794 (N_4794,In_2096,In_2168);
xor U4795 (N_4795,In_410,In_1238);
xnor U4796 (N_4796,In_1906,In_1011);
xor U4797 (N_4797,In_588,In_1409);
or U4798 (N_4798,In_286,In_2314);
nor U4799 (N_4799,In_178,In_1113);
xnor U4800 (N_4800,In_751,In_1500);
nand U4801 (N_4801,In_614,In_1119);
nor U4802 (N_4802,In_82,In_2262);
nand U4803 (N_4803,In_801,In_708);
or U4804 (N_4804,In_176,In_2373);
nand U4805 (N_4805,In_38,In_2314);
and U4806 (N_4806,In_738,In_2384);
nand U4807 (N_4807,In_2374,In_492);
xnor U4808 (N_4808,In_1681,In_2464);
xnor U4809 (N_4809,In_283,In_1551);
xnor U4810 (N_4810,In_2205,In_810);
or U4811 (N_4811,In_1422,In_935);
nand U4812 (N_4812,In_2034,In_235);
and U4813 (N_4813,In_1740,In_1648);
and U4814 (N_4814,In_1565,In_1386);
xnor U4815 (N_4815,In_1075,In_1852);
xor U4816 (N_4816,In_1428,In_1465);
and U4817 (N_4817,In_341,In_593);
or U4818 (N_4818,In_384,In_559);
xor U4819 (N_4819,In_1574,In_1347);
nand U4820 (N_4820,In_495,In_514);
and U4821 (N_4821,In_2244,In_2031);
nand U4822 (N_4822,In_2005,In_948);
xnor U4823 (N_4823,In_852,In_754);
xnor U4824 (N_4824,In_1701,In_1871);
xnor U4825 (N_4825,In_790,In_2125);
xnor U4826 (N_4826,In_1549,In_1206);
or U4827 (N_4827,In_1282,In_1436);
xnor U4828 (N_4828,In_1984,In_1564);
and U4829 (N_4829,In_1888,In_613);
and U4830 (N_4830,In_2138,In_1109);
or U4831 (N_4831,In_2248,In_2145);
or U4832 (N_4832,In_2467,In_2313);
nand U4833 (N_4833,In_510,In_1190);
xnor U4834 (N_4834,In_2370,In_1304);
or U4835 (N_4835,In_2165,In_1653);
and U4836 (N_4836,In_798,In_1027);
nor U4837 (N_4837,In_2331,In_1252);
xnor U4838 (N_4838,In_781,In_1830);
or U4839 (N_4839,In_2163,In_196);
and U4840 (N_4840,In_2218,In_2463);
xor U4841 (N_4841,In_981,In_1306);
or U4842 (N_4842,In_841,In_2243);
and U4843 (N_4843,In_659,In_2261);
xor U4844 (N_4844,In_2360,In_2340);
nand U4845 (N_4845,In_2029,In_18);
and U4846 (N_4846,In_979,In_2257);
nand U4847 (N_4847,In_643,In_324);
or U4848 (N_4848,In_1109,In_1525);
or U4849 (N_4849,In_1057,In_2023);
and U4850 (N_4850,In_1162,In_1925);
nand U4851 (N_4851,In_1658,In_1308);
or U4852 (N_4852,In_1718,In_1984);
nor U4853 (N_4853,In_1128,In_1416);
nand U4854 (N_4854,In_1317,In_1614);
nand U4855 (N_4855,In_1654,In_2060);
xor U4856 (N_4856,In_1246,In_2444);
nor U4857 (N_4857,In_2060,In_2439);
or U4858 (N_4858,In_2080,In_51);
nor U4859 (N_4859,In_1590,In_2280);
xnor U4860 (N_4860,In_668,In_983);
nand U4861 (N_4861,In_1724,In_174);
nand U4862 (N_4862,In_709,In_1646);
and U4863 (N_4863,In_544,In_474);
nand U4864 (N_4864,In_485,In_1469);
and U4865 (N_4865,In_1557,In_1282);
xor U4866 (N_4866,In_719,In_1970);
nor U4867 (N_4867,In_79,In_737);
xnor U4868 (N_4868,In_1916,In_122);
and U4869 (N_4869,In_1480,In_1400);
or U4870 (N_4870,In_1726,In_909);
and U4871 (N_4871,In_631,In_2438);
nand U4872 (N_4872,In_832,In_690);
or U4873 (N_4873,In_1876,In_2304);
and U4874 (N_4874,In_1225,In_1519);
and U4875 (N_4875,In_456,In_1383);
nand U4876 (N_4876,In_1865,In_1338);
or U4877 (N_4877,In_752,In_1768);
or U4878 (N_4878,In_2315,In_295);
nand U4879 (N_4879,In_1521,In_853);
or U4880 (N_4880,In_2282,In_557);
nor U4881 (N_4881,In_1135,In_1578);
xnor U4882 (N_4882,In_1393,In_632);
xnor U4883 (N_4883,In_1425,In_305);
or U4884 (N_4884,In_1649,In_2297);
nand U4885 (N_4885,In_1329,In_1388);
or U4886 (N_4886,In_1807,In_588);
or U4887 (N_4887,In_1096,In_549);
xnor U4888 (N_4888,In_990,In_319);
or U4889 (N_4889,In_2349,In_573);
or U4890 (N_4890,In_1279,In_1095);
and U4891 (N_4891,In_2289,In_2310);
or U4892 (N_4892,In_1268,In_786);
and U4893 (N_4893,In_2490,In_1266);
xnor U4894 (N_4894,In_1595,In_90);
nand U4895 (N_4895,In_278,In_1579);
xnor U4896 (N_4896,In_724,In_1072);
and U4897 (N_4897,In_1375,In_790);
and U4898 (N_4898,In_1483,In_850);
or U4899 (N_4899,In_1573,In_1464);
or U4900 (N_4900,In_307,In_2019);
xnor U4901 (N_4901,In_2055,In_413);
or U4902 (N_4902,In_994,In_115);
and U4903 (N_4903,In_57,In_2148);
or U4904 (N_4904,In_525,In_1312);
nor U4905 (N_4905,In_1492,In_591);
and U4906 (N_4906,In_691,In_2178);
nor U4907 (N_4907,In_467,In_2376);
or U4908 (N_4908,In_1910,In_2181);
xor U4909 (N_4909,In_2083,In_657);
and U4910 (N_4910,In_502,In_487);
or U4911 (N_4911,In_189,In_588);
or U4912 (N_4912,In_1437,In_1159);
xor U4913 (N_4913,In_1887,In_1241);
nand U4914 (N_4914,In_2079,In_1726);
and U4915 (N_4915,In_721,In_219);
nand U4916 (N_4916,In_1508,In_607);
or U4917 (N_4917,In_2245,In_494);
nand U4918 (N_4918,In_422,In_848);
nand U4919 (N_4919,In_1712,In_1491);
nor U4920 (N_4920,In_1630,In_1201);
nand U4921 (N_4921,In_1920,In_1240);
or U4922 (N_4922,In_1290,In_1202);
or U4923 (N_4923,In_569,In_1724);
and U4924 (N_4924,In_149,In_15);
and U4925 (N_4925,In_575,In_1503);
or U4926 (N_4926,In_175,In_1385);
or U4927 (N_4927,In_526,In_1839);
nand U4928 (N_4928,In_1864,In_2137);
and U4929 (N_4929,In_705,In_1848);
nand U4930 (N_4930,In_1942,In_1603);
nor U4931 (N_4931,In_395,In_897);
and U4932 (N_4932,In_1622,In_1530);
nand U4933 (N_4933,In_2362,In_418);
nand U4934 (N_4934,In_2351,In_2280);
nand U4935 (N_4935,In_1202,In_245);
xor U4936 (N_4936,In_1351,In_1829);
xor U4937 (N_4937,In_1961,In_388);
or U4938 (N_4938,In_512,In_236);
xor U4939 (N_4939,In_2186,In_2079);
nor U4940 (N_4940,In_1779,In_2327);
and U4941 (N_4941,In_1868,In_608);
xnor U4942 (N_4942,In_1853,In_1867);
and U4943 (N_4943,In_2003,In_2389);
nor U4944 (N_4944,In_154,In_861);
nor U4945 (N_4945,In_1292,In_311);
nand U4946 (N_4946,In_1829,In_0);
or U4947 (N_4947,In_2468,In_813);
nand U4948 (N_4948,In_2402,In_127);
nand U4949 (N_4949,In_2450,In_85);
nor U4950 (N_4950,In_887,In_1549);
and U4951 (N_4951,In_691,In_320);
and U4952 (N_4952,In_1019,In_1063);
nor U4953 (N_4953,In_526,In_220);
or U4954 (N_4954,In_1132,In_397);
nor U4955 (N_4955,In_359,In_2170);
and U4956 (N_4956,In_723,In_1890);
nor U4957 (N_4957,In_1353,In_73);
nand U4958 (N_4958,In_962,In_236);
or U4959 (N_4959,In_1216,In_1621);
or U4960 (N_4960,In_628,In_1162);
xor U4961 (N_4961,In_1072,In_1803);
xor U4962 (N_4962,In_683,In_609);
xor U4963 (N_4963,In_953,In_1105);
nand U4964 (N_4964,In_494,In_1846);
nand U4965 (N_4965,In_787,In_2371);
and U4966 (N_4966,In_1263,In_2208);
and U4967 (N_4967,In_878,In_684);
xnor U4968 (N_4968,In_589,In_402);
or U4969 (N_4969,In_736,In_1178);
nand U4970 (N_4970,In_1470,In_1380);
and U4971 (N_4971,In_2206,In_539);
xor U4972 (N_4972,In_240,In_1211);
nand U4973 (N_4973,In_2243,In_2411);
or U4974 (N_4974,In_2061,In_2416);
nand U4975 (N_4975,In_125,In_1331);
or U4976 (N_4976,In_1707,In_2133);
and U4977 (N_4977,In_132,In_56);
nand U4978 (N_4978,In_1074,In_934);
and U4979 (N_4979,In_714,In_865);
xnor U4980 (N_4980,In_1026,In_1167);
nor U4981 (N_4981,In_218,In_669);
nand U4982 (N_4982,In_31,In_200);
nand U4983 (N_4983,In_2496,In_71);
and U4984 (N_4984,In_550,In_990);
nor U4985 (N_4985,In_2057,In_1413);
nand U4986 (N_4986,In_417,In_1481);
and U4987 (N_4987,In_2283,In_1545);
and U4988 (N_4988,In_2308,In_2162);
and U4989 (N_4989,In_2119,In_1781);
nor U4990 (N_4990,In_1663,In_33);
and U4991 (N_4991,In_1529,In_565);
or U4992 (N_4992,In_2184,In_904);
or U4993 (N_4993,In_1280,In_401);
xnor U4994 (N_4994,In_342,In_2401);
nand U4995 (N_4995,In_680,In_1787);
and U4996 (N_4996,In_1232,In_1990);
nor U4997 (N_4997,In_52,In_1869);
or U4998 (N_4998,In_1374,In_2057);
or U4999 (N_4999,In_1427,In_1470);
nand U5000 (N_5000,N_3005,N_1294);
xnor U5001 (N_5001,N_4120,N_1735);
nor U5002 (N_5002,N_3718,N_2549);
xor U5003 (N_5003,N_4500,N_576);
nor U5004 (N_5004,N_2073,N_592);
and U5005 (N_5005,N_2785,N_2929);
nor U5006 (N_5006,N_2240,N_157);
nor U5007 (N_5007,N_50,N_781);
and U5008 (N_5008,N_673,N_2668);
or U5009 (N_5009,N_35,N_4968);
and U5010 (N_5010,N_1141,N_2288);
xnor U5011 (N_5011,N_3224,N_1049);
and U5012 (N_5012,N_2617,N_4157);
nor U5013 (N_5013,N_1787,N_3086);
nand U5014 (N_5014,N_49,N_4245);
or U5015 (N_5015,N_3317,N_1944);
and U5016 (N_5016,N_1633,N_1919);
nand U5017 (N_5017,N_4634,N_2208);
and U5018 (N_5018,N_3945,N_688);
or U5019 (N_5019,N_1535,N_3211);
and U5020 (N_5020,N_1279,N_2249);
nand U5021 (N_5021,N_3199,N_3433);
nor U5022 (N_5022,N_907,N_2887);
nor U5023 (N_5023,N_1712,N_3238);
nand U5024 (N_5024,N_950,N_602);
xnor U5025 (N_5025,N_2421,N_2134);
and U5026 (N_5026,N_4626,N_4525);
nand U5027 (N_5027,N_2539,N_4970);
and U5028 (N_5028,N_4305,N_2512);
xor U5029 (N_5029,N_4855,N_3228);
nand U5030 (N_5030,N_4177,N_614);
and U5031 (N_5031,N_2868,N_4702);
and U5032 (N_5032,N_1488,N_2172);
xnor U5033 (N_5033,N_4668,N_2173);
xor U5034 (N_5034,N_2385,N_1589);
xor U5035 (N_5035,N_4567,N_3797);
nor U5036 (N_5036,N_1047,N_94);
or U5037 (N_5037,N_993,N_4040);
nor U5038 (N_5038,N_4102,N_2349);
nor U5039 (N_5039,N_2825,N_1737);
and U5040 (N_5040,N_4793,N_662);
or U5041 (N_5041,N_3287,N_288);
or U5042 (N_5042,N_423,N_4153);
nor U5043 (N_5043,N_2462,N_1318);
nor U5044 (N_5044,N_4255,N_4532);
nand U5045 (N_5045,N_2739,N_2057);
nand U5046 (N_5046,N_1845,N_3314);
nand U5047 (N_5047,N_2426,N_2020);
xor U5048 (N_5048,N_4029,N_635);
xnor U5049 (N_5049,N_3331,N_891);
nor U5050 (N_5050,N_1829,N_231);
nand U5051 (N_5051,N_3673,N_1676);
and U5052 (N_5052,N_4595,N_413);
nor U5053 (N_5053,N_1616,N_3665);
or U5054 (N_5054,N_1500,N_3133);
and U5055 (N_5055,N_1503,N_1766);
or U5056 (N_5056,N_1144,N_1809);
nand U5057 (N_5057,N_3707,N_73);
or U5058 (N_5058,N_3068,N_151);
nand U5059 (N_5059,N_1950,N_871);
and U5060 (N_5060,N_2720,N_646);
and U5061 (N_5061,N_4164,N_731);
or U5062 (N_5062,N_3070,N_2333);
xor U5063 (N_5063,N_3705,N_2370);
xor U5064 (N_5064,N_4172,N_902);
xnor U5065 (N_5065,N_1752,N_4267);
and U5066 (N_5066,N_2460,N_496);
xor U5067 (N_5067,N_2055,N_400);
or U5068 (N_5068,N_2448,N_2352);
nand U5069 (N_5069,N_3107,N_4328);
and U5070 (N_5070,N_2640,N_3468);
nor U5071 (N_5071,N_2604,N_4998);
xnor U5072 (N_5072,N_3594,N_2544);
nor U5073 (N_5073,N_184,N_1137);
nor U5074 (N_5074,N_2420,N_1369);
nand U5075 (N_5075,N_2557,N_3613);
and U5076 (N_5076,N_1962,N_4447);
or U5077 (N_5077,N_259,N_2775);
xor U5078 (N_5078,N_3431,N_1731);
nor U5079 (N_5079,N_1446,N_2965);
or U5080 (N_5080,N_973,N_3593);
nor U5081 (N_5081,N_86,N_1763);
or U5082 (N_5082,N_4508,N_2708);
or U5083 (N_5083,N_4332,N_4146);
nand U5084 (N_5084,N_970,N_1903);
nand U5085 (N_5085,N_4200,N_2568);
nor U5086 (N_5086,N_3580,N_440);
nand U5087 (N_5087,N_3637,N_2910);
nor U5088 (N_5088,N_818,N_3085);
nor U5089 (N_5089,N_1365,N_4147);
and U5090 (N_5090,N_1689,N_57);
or U5091 (N_5091,N_1352,N_1884);
xnor U5092 (N_5092,N_725,N_1484);
and U5093 (N_5093,N_997,N_3957);
or U5094 (N_5094,N_1439,N_4050);
or U5095 (N_5095,N_586,N_794);
or U5096 (N_5096,N_2966,N_1552);
or U5097 (N_5097,N_4167,N_2136);
nor U5098 (N_5098,N_715,N_642);
and U5099 (N_5099,N_4947,N_1240);
or U5100 (N_5100,N_358,N_4647);
nor U5101 (N_5101,N_4457,N_3024);
xor U5102 (N_5102,N_4183,N_4234);
xnor U5103 (N_5103,N_2669,N_3730);
nor U5104 (N_5104,N_2920,N_2443);
and U5105 (N_5105,N_3509,N_3448);
or U5106 (N_5106,N_1195,N_4360);
nand U5107 (N_5107,N_2735,N_2287);
nor U5108 (N_5108,N_3479,N_733);
xnor U5109 (N_5109,N_821,N_3130);
nand U5110 (N_5110,N_3377,N_2300);
nor U5111 (N_5111,N_2493,N_4939);
or U5112 (N_5112,N_4299,N_410);
nor U5113 (N_5113,N_1678,N_4176);
nand U5114 (N_5114,N_1066,N_4964);
or U5115 (N_5115,N_2991,N_2744);
nand U5116 (N_5116,N_3848,N_3217);
and U5117 (N_5117,N_2268,N_1349);
nand U5118 (N_5118,N_757,N_146);
and U5119 (N_5119,N_1860,N_738);
xor U5120 (N_5120,N_308,N_1476);
nor U5121 (N_5121,N_1409,N_4208);
nor U5122 (N_5122,N_1230,N_2859);
and U5123 (N_5123,N_2398,N_4302);
nor U5124 (N_5124,N_3060,N_718);
and U5125 (N_5125,N_2409,N_2573);
xor U5126 (N_5126,N_4364,N_1063);
or U5127 (N_5127,N_3305,N_4489);
and U5128 (N_5128,N_3033,N_3459);
nand U5129 (N_5129,N_4286,N_4722);
nand U5130 (N_5130,N_4707,N_4432);
xor U5131 (N_5131,N_1213,N_3345);
xnor U5132 (N_5132,N_2611,N_1284);
nor U5133 (N_5133,N_1605,N_4784);
and U5134 (N_5134,N_3408,N_4428);
and U5135 (N_5135,N_4058,N_3414);
nor U5136 (N_5136,N_4469,N_3943);
xnor U5137 (N_5137,N_2464,N_269);
or U5138 (N_5138,N_1339,N_1810);
nor U5139 (N_5139,N_3187,N_1592);
and U5140 (N_5140,N_3353,N_1899);
or U5141 (N_5141,N_765,N_2417);
or U5142 (N_5142,N_3854,N_986);
xor U5143 (N_5143,N_3726,N_778);
and U5144 (N_5144,N_2927,N_1783);
nor U5145 (N_5145,N_219,N_4435);
nand U5146 (N_5146,N_1558,N_4529);
or U5147 (N_5147,N_932,N_2272);
nand U5148 (N_5148,N_3778,N_3889);
or U5149 (N_5149,N_499,N_2908);
and U5150 (N_5150,N_1869,N_88);
nand U5151 (N_5151,N_2742,N_2362);
nand U5152 (N_5152,N_1383,N_1357);
nor U5153 (N_5153,N_4690,N_2657);
nor U5154 (N_5154,N_1874,N_2941);
xor U5155 (N_5155,N_3050,N_2283);
and U5156 (N_5156,N_3900,N_2909);
xor U5157 (N_5157,N_418,N_3527);
and U5158 (N_5158,N_1929,N_4315);
nand U5159 (N_5159,N_4069,N_1483);
nor U5160 (N_5160,N_3684,N_3375);
and U5161 (N_5161,N_1041,N_2151);
or U5162 (N_5162,N_600,N_2865);
nand U5163 (N_5163,N_516,N_3501);
nor U5164 (N_5164,N_3746,N_491);
nand U5165 (N_5165,N_3012,N_2676);
xor U5166 (N_5166,N_436,N_807);
nand U5167 (N_5167,N_4415,N_1867);
xnor U5168 (N_5168,N_3939,N_2995);
xnor U5169 (N_5169,N_2722,N_1090);
and U5170 (N_5170,N_2623,N_1842);
xnor U5171 (N_5171,N_1632,N_2156);
and U5172 (N_5172,N_434,N_3052);
and U5173 (N_5173,N_1539,N_1348);
and U5174 (N_5174,N_2394,N_849);
nand U5175 (N_5175,N_2190,N_3584);
nor U5176 (N_5176,N_952,N_553);
or U5177 (N_5177,N_3011,N_4561);
nor U5178 (N_5178,N_36,N_812);
nor U5179 (N_5179,N_1458,N_2595);
xor U5180 (N_5180,N_2508,N_4962);
xor U5181 (N_5181,N_3197,N_1186);
and U5182 (N_5182,N_4752,N_2846);
and U5183 (N_5183,N_3349,N_2691);
or U5184 (N_5184,N_3624,N_3007);
nand U5185 (N_5185,N_4761,N_4861);
xnor U5186 (N_5186,N_506,N_580);
or U5187 (N_5187,N_4699,N_4052);
and U5188 (N_5188,N_1868,N_4353);
and U5189 (N_5189,N_4995,N_1580);
xor U5190 (N_5190,N_1865,N_2457);
xor U5191 (N_5191,N_3833,N_3378);
and U5192 (N_5192,N_1894,N_533);
xor U5193 (N_5193,N_2752,N_4689);
nor U5194 (N_5194,N_1401,N_3789);
nand U5195 (N_5195,N_1119,N_1293);
or U5196 (N_5196,N_2751,N_1264);
nand U5197 (N_5197,N_4021,N_1720);
or U5198 (N_5198,N_3556,N_1126);
or U5199 (N_5199,N_574,N_3427);
and U5200 (N_5200,N_3505,N_3524);
and U5201 (N_5201,N_4000,N_4913);
xor U5202 (N_5202,N_1654,N_4279);
xor U5203 (N_5203,N_2475,N_4882);
or U5204 (N_5204,N_1344,N_2914);
and U5205 (N_5205,N_2890,N_3341);
nor U5206 (N_5206,N_2748,N_451);
and U5207 (N_5207,N_937,N_4204);
or U5208 (N_5208,N_540,N_485);
and U5209 (N_5209,N_1496,N_1966);
and U5210 (N_5210,N_3991,N_158);
or U5211 (N_5211,N_3037,N_1262);
nand U5212 (N_5212,N_1743,N_1407);
and U5213 (N_5213,N_664,N_2343);
or U5214 (N_5214,N_2149,N_1800);
nand U5215 (N_5215,N_579,N_1398);
or U5216 (N_5216,N_2561,N_2590);
nor U5217 (N_5217,N_2569,N_2145);
nand U5218 (N_5218,N_4898,N_3102);
or U5219 (N_5219,N_252,N_4413);
or U5220 (N_5220,N_1555,N_3255);
xor U5221 (N_5221,N_1643,N_2298);
nand U5222 (N_5222,N_647,N_3625);
or U5223 (N_5223,N_4398,N_1817);
nor U5224 (N_5224,N_3484,N_1405);
or U5225 (N_5225,N_3793,N_3763);
or U5226 (N_5226,N_4080,N_989);
nand U5227 (N_5227,N_1173,N_1825);
nor U5228 (N_5228,N_4874,N_724);
nor U5229 (N_5229,N_4277,N_4017);
or U5230 (N_5230,N_170,N_1104);
xnor U5231 (N_5231,N_2044,N_4454);
or U5232 (N_5232,N_3291,N_3764);
or U5233 (N_5233,N_3622,N_4909);
and U5234 (N_5234,N_1662,N_4822);
nor U5235 (N_5235,N_2442,N_2982);
and U5236 (N_5236,N_2052,N_3172);
or U5237 (N_5237,N_2094,N_813);
or U5238 (N_5238,N_4853,N_4892);
and U5239 (N_5239,N_4429,N_3589);
nand U5240 (N_5240,N_1515,N_3340);
nand U5241 (N_5241,N_1375,N_1755);
or U5242 (N_5242,N_1187,N_1621);
xnor U5243 (N_5243,N_1494,N_2819);
xor U5244 (N_5244,N_2229,N_946);
xnor U5245 (N_5245,N_3495,N_822);
nand U5246 (N_5246,N_3901,N_636);
nor U5247 (N_5247,N_919,N_466);
xnor U5248 (N_5248,N_4133,N_3652);
and U5249 (N_5249,N_357,N_2210);
or U5250 (N_5250,N_3771,N_483);
nand U5251 (N_5251,N_3947,N_4341);
or U5252 (N_5252,N_622,N_3091);
nand U5253 (N_5253,N_263,N_633);
nor U5254 (N_5254,N_3599,N_2245);
and U5255 (N_5255,N_1099,N_2345);
and U5256 (N_5256,N_530,N_2033);
nand U5257 (N_5257,N_3709,N_141);
nor U5258 (N_5258,N_4825,N_159);
nand U5259 (N_5259,N_603,N_1017);
nand U5260 (N_5260,N_3549,N_1431);
or U5261 (N_5261,N_4673,N_4691);
nand U5262 (N_5262,N_2554,N_1360);
nor U5263 (N_5263,N_3232,N_2692);
nor U5264 (N_5264,N_1329,N_2811);
or U5265 (N_5265,N_1132,N_3811);
and U5266 (N_5266,N_3319,N_2129);
or U5267 (N_5267,N_2350,N_367);
and U5268 (N_5268,N_3098,N_3710);
and U5269 (N_5269,N_1208,N_3541);
or U5270 (N_5270,N_113,N_4908);
xor U5271 (N_5271,N_3888,N_3571);
or U5272 (N_5272,N_3065,N_4151);
nor U5273 (N_5273,N_4110,N_3696);
nor U5274 (N_5274,N_3016,N_2894);
nor U5275 (N_5275,N_1200,N_2491);
or U5276 (N_5276,N_1928,N_4078);
or U5277 (N_5277,N_4845,N_2436);
xor U5278 (N_5278,N_3756,N_4785);
nand U5279 (N_5279,N_38,N_3032);
nor U5280 (N_5280,N_2912,N_843);
nand U5281 (N_5281,N_48,N_2826);
or U5282 (N_5282,N_44,N_599);
or U5283 (N_5283,N_4308,N_2030);
xor U5284 (N_5284,N_167,N_3055);
nor U5285 (N_5285,N_2897,N_3225);
nand U5286 (N_5286,N_3270,N_2200);
or U5287 (N_5287,N_4813,N_4384);
or U5288 (N_5288,N_1669,N_3678);
nor U5289 (N_5289,N_1337,N_2083);
and U5290 (N_5290,N_2183,N_2061);
nor U5291 (N_5291,N_4303,N_796);
and U5292 (N_5292,N_3181,N_2821);
xnor U5293 (N_5293,N_4246,N_1875);
nor U5294 (N_5294,N_4678,N_2278);
nand U5295 (N_5295,N_4307,N_2233);
xor U5296 (N_5296,N_4560,N_2516);
nand U5297 (N_5297,N_1688,N_3041);
nor U5298 (N_5298,N_445,N_2437);
nand U5299 (N_5299,N_2559,N_1718);
or U5300 (N_5300,N_3126,N_1523);
nand U5301 (N_5301,N_284,N_4141);
xor U5302 (N_5302,N_1659,N_0);
and U5303 (N_5303,N_3499,N_3231);
and U5304 (N_5304,N_3667,N_1699);
xnor U5305 (N_5305,N_751,N_4425);
or U5306 (N_5306,N_2483,N_1770);
nor U5307 (N_5307,N_2886,N_320);
and U5308 (N_5308,N_3140,N_2987);
nand U5309 (N_5309,N_2984,N_4282);
nor U5310 (N_5310,N_3972,N_1571);
nor U5311 (N_5311,N_4854,N_1276);
nor U5312 (N_5312,N_735,N_4731);
nand U5313 (N_5313,N_1641,N_2497);
nand U5314 (N_5314,N_4756,N_1105);
nand U5315 (N_5315,N_1316,N_2401);
or U5316 (N_5316,N_957,N_1573);
nor U5317 (N_5317,N_960,N_850);
xor U5318 (N_5318,N_3471,N_1858);
or U5319 (N_5319,N_1498,N_2614);
nor U5320 (N_5320,N_1493,N_3034);
nor U5321 (N_5321,N_2289,N_2851);
nand U5322 (N_5322,N_4348,N_2131);
nand U5323 (N_5323,N_111,N_248);
xor U5324 (N_5324,N_2893,N_2608);
nand U5325 (N_5325,N_4330,N_4217);
nand U5326 (N_5326,N_2209,N_3721);
or U5327 (N_5327,N_2205,N_2452);
nor U5328 (N_5328,N_4827,N_304);
nand U5329 (N_5329,N_3500,N_4240);
or U5330 (N_5330,N_1815,N_2400);
nand U5331 (N_5331,N_3203,N_2662);
and U5332 (N_5332,N_2137,N_1006);
nand U5333 (N_5333,N_1430,N_2902);
nor U5334 (N_5334,N_1368,N_3653);
nor U5335 (N_5335,N_1038,N_1345);
nor U5336 (N_5336,N_766,N_3765);
or U5337 (N_5337,N_562,N_1915);
nand U5338 (N_5338,N_3389,N_4796);
and U5339 (N_5339,N_1355,N_4739);
nor U5340 (N_5340,N_1435,N_4296);
nand U5341 (N_5341,N_108,N_1680);
or U5342 (N_5342,N_218,N_4966);
and U5343 (N_5343,N_2935,N_1436);
xor U5344 (N_5344,N_2189,N_2683);
or U5345 (N_5345,N_4830,N_2015);
and U5346 (N_5346,N_2678,N_2986);
or U5347 (N_5347,N_4852,N_3935);
nor U5348 (N_5348,N_360,N_255);
or U5349 (N_5349,N_3292,N_4883);
nor U5350 (N_5350,N_215,N_2024);
and U5351 (N_5351,N_1615,N_1984);
or U5352 (N_5352,N_2727,N_3142);
xor U5353 (N_5353,N_3151,N_2973);
nand U5354 (N_5354,N_2833,N_3585);
and U5355 (N_5355,N_3320,N_4973);
xnor U5356 (N_5356,N_2588,N_1789);
and U5357 (N_5357,N_4715,N_2251);
or U5358 (N_5358,N_1343,N_1275);
xor U5359 (N_5359,N_4817,N_2857);
and U5360 (N_5360,N_4035,N_183);
xor U5361 (N_5361,N_2327,N_4979);
xnor U5362 (N_5362,N_1855,N_3845);
xor U5363 (N_5363,N_4810,N_3831);
or U5364 (N_5364,N_1889,N_3394);
or U5365 (N_5365,N_526,N_2427);
and U5366 (N_5366,N_54,N_3761);
or U5367 (N_5367,N_1269,N_2123);
and U5368 (N_5368,N_234,N_1779);
or U5369 (N_5369,N_4503,N_4181);
xnor U5370 (N_5370,N_4137,N_1265);
nor U5371 (N_5371,N_119,N_3738);
nor U5372 (N_5372,N_250,N_1084);
or U5373 (N_5373,N_3374,N_4187);
xor U5374 (N_5374,N_1157,N_4642);
xor U5375 (N_5375,N_1522,N_223);
nand U5376 (N_5376,N_969,N_1131);
and U5377 (N_5377,N_4582,N_4911);
or U5378 (N_5378,N_4088,N_2509);
xor U5379 (N_5379,N_3640,N_4372);
xor U5380 (N_5380,N_3694,N_2037);
xor U5381 (N_5381,N_1051,N_3716);
nor U5382 (N_5382,N_1354,N_2999);
nor U5383 (N_5383,N_4732,N_3649);
or U5384 (N_5384,N_2853,N_4004);
and U5385 (N_5385,N_1241,N_251);
or U5386 (N_5386,N_4700,N_2194);
or U5387 (N_5387,N_3534,N_3259);
or U5388 (N_5388,N_1191,N_2356);
and U5389 (N_5389,N_4263,N_1347);
nor U5390 (N_5390,N_4007,N_1491);
or U5391 (N_5391,N_652,N_903);
xnor U5392 (N_5392,N_192,N_93);
and U5393 (N_5393,N_1513,N_4518);
xor U5394 (N_5394,N_4608,N_550);
xnor U5395 (N_5395,N_3141,N_3766);
nand U5396 (N_5396,N_3336,N_1952);
nand U5397 (N_5397,N_4178,N_3128);
and U5398 (N_5398,N_2757,N_2891);
or U5399 (N_5399,N_2503,N_165);
and U5400 (N_5400,N_3608,N_492);
nor U5401 (N_5401,N_2911,N_484);
xor U5402 (N_5402,N_131,N_4742);
or U5403 (N_5403,N_438,N_901);
nand U5404 (N_5404,N_3355,N_2571);
nor U5405 (N_5405,N_4087,N_887);
nor U5406 (N_5406,N_4190,N_2458);
xor U5407 (N_5407,N_963,N_462);
xor U5408 (N_5408,N_198,N_498);
or U5409 (N_5409,N_3516,N_3917);
or U5410 (N_5410,N_908,N_2788);
and U5411 (N_5411,N_3736,N_979);
xnor U5412 (N_5412,N_4904,N_3164);
nand U5413 (N_5413,N_282,N_836);
nand U5414 (N_5414,N_2117,N_2424);
nand U5415 (N_5415,N_137,N_426);
or U5416 (N_5416,N_2135,N_1774);
xor U5417 (N_5417,N_1989,N_4154);
nand U5418 (N_5418,N_2253,N_2499);
or U5419 (N_5419,N_4149,N_4340);
and U5420 (N_5420,N_2316,N_4477);
and U5421 (N_5421,N_1819,N_1864);
xor U5422 (N_5422,N_904,N_22);
nand U5423 (N_5423,N_4757,N_2876);
xnor U5424 (N_5424,N_4480,N_1035);
and U5425 (N_5425,N_4140,N_3268);
nand U5426 (N_5426,N_1486,N_81);
and U5427 (N_5427,N_107,N_4236);
or U5428 (N_5428,N_3077,N_1304);
and U5429 (N_5429,N_2848,N_3798);
nand U5430 (N_5430,N_4649,N_1679);
xnor U5431 (N_5431,N_182,N_1217);
or U5432 (N_5432,N_4888,N_214);
nand U5433 (N_5433,N_3117,N_2959);
xor U5434 (N_5434,N_1568,N_4060);
and U5435 (N_5435,N_1353,N_4651);
nand U5436 (N_5436,N_3207,N_2658);
nand U5437 (N_5437,N_4259,N_501);
xnor U5438 (N_5438,N_569,N_2505);
xor U5439 (N_5439,N_2585,N_4772);
and U5440 (N_5440,N_2084,N_3089);
nor U5441 (N_5441,N_2105,N_3338);
nor U5442 (N_5442,N_193,N_2337);
and U5443 (N_5443,N_639,N_4184);
and U5444 (N_5444,N_2671,N_4346);
nand U5445 (N_5445,N_3193,N_741);
and U5446 (N_5446,N_555,N_548);
xnor U5447 (N_5447,N_4894,N_2125);
or U5448 (N_5448,N_2925,N_645);
nor U5449 (N_5449,N_285,N_3734);
or U5450 (N_5450,N_1773,N_2867);
xnor U5451 (N_5451,N_938,N_3732);
and U5452 (N_5452,N_566,N_4925);
or U5453 (N_5453,N_3137,N_118);
or U5454 (N_5454,N_1070,N_628);
nand U5455 (N_5455,N_4490,N_1999);
nor U5456 (N_5456,N_1022,N_4963);
nand U5457 (N_5457,N_3583,N_1754);
nor U5458 (N_5458,N_2041,N_3620);
or U5459 (N_5459,N_3648,N_1273);
or U5460 (N_5460,N_3456,N_1146);
xnor U5461 (N_5461,N_1060,N_3256);
nor U5462 (N_5462,N_53,N_1777);
nand U5463 (N_5463,N_1061,N_3426);
nand U5464 (N_5464,N_4790,N_4958);
nor U5465 (N_5465,N_4540,N_611);
or U5466 (N_5466,N_816,N_2180);
nor U5467 (N_5467,N_776,N_1741);
or U5468 (N_5468,N_2005,N_3159);
xnor U5469 (N_5469,N_4129,N_2586);
xnor U5470 (N_5470,N_814,N_1167);
nand U5471 (N_5471,N_2254,N_1156);
and U5472 (N_5472,N_3868,N_4583);
xnor U5473 (N_5473,N_3,N_1802);
or U5474 (N_5474,N_4066,N_2746);
nor U5475 (N_5475,N_3597,N_1482);
xor U5476 (N_5476,N_1564,N_359);
or U5477 (N_5477,N_267,N_99);
and U5478 (N_5478,N_2017,N_3245);
or U5479 (N_5479,N_701,N_421);
xor U5480 (N_5480,N_2315,N_1531);
nor U5481 (N_5481,N_333,N_1581);
nor U5482 (N_5482,N_1882,N_3173);
nor U5483 (N_5483,N_1941,N_1795);
and U5484 (N_5484,N_2144,N_2526);
nand U5485 (N_5485,N_1601,N_1653);
nand U5486 (N_5486,N_705,N_4310);
xnor U5487 (N_5487,N_4418,N_4719);
xnor U5488 (N_5488,N_3985,N_175);
nand U5489 (N_5489,N_2074,N_3508);
nor U5490 (N_5490,N_3783,N_2332);
nand U5491 (N_5491,N_2150,N_309);
nor U5492 (N_5492,N_3576,N_1033);
nor U5493 (N_5493,N_139,N_4455);
and U5494 (N_5494,N_3916,N_361);
and U5495 (N_5495,N_3361,N_852);
or U5496 (N_5496,N_4268,N_2772);
and U5497 (N_5497,N_681,N_1728);
nor U5498 (N_5498,N_2672,N_2078);
nor U5499 (N_5499,N_444,N_4304);
nor U5500 (N_5500,N_1668,N_612);
nand U5501 (N_5501,N_64,N_3719);
and U5502 (N_5502,N_3729,N_3153);
or U5503 (N_5503,N_4048,N_1321);
or U5504 (N_5504,N_3101,N_3038);
nor U5505 (N_5505,N_4747,N_2781);
or U5506 (N_5506,N_189,N_1462);
nor U5507 (N_5507,N_4549,N_3445);
nor U5508 (N_5508,N_678,N_3298);
or U5509 (N_5509,N_2242,N_4917);
xor U5510 (N_5510,N_3990,N_867);
and U5511 (N_5511,N_2711,N_510);
xnor U5512 (N_5512,N_3112,N_3960);
or U5513 (N_5513,N_4256,N_1590);
and U5514 (N_5514,N_3602,N_621);
nand U5515 (N_5515,N_4230,N_2661);
nand U5516 (N_5516,N_3276,N_1);
xnor U5517 (N_5517,N_4528,N_3432);
and U5518 (N_5518,N_1297,N_162);
or U5519 (N_5519,N_3569,N_4414);
and U5520 (N_5520,N_1717,N_2587);
nand U5521 (N_5521,N_4682,N_1016);
xnor U5522 (N_5522,N_1872,N_889);
xnor U5523 (N_5523,N_3849,N_3940);
nand U5524 (N_5524,N_1546,N_2670);
xnor U5525 (N_5525,N_1071,N_1254);
and U5526 (N_5526,N_2800,N_1323);
and U5527 (N_5527,N_60,N_3056);
nand U5528 (N_5528,N_3266,N_1960);
xnor U5529 (N_5529,N_3806,N_3220);
or U5530 (N_5530,N_2884,N_3782);
nand U5531 (N_5531,N_3697,N_1412);
xnor U5532 (N_5532,N_2085,N_1670);
nand U5533 (N_5533,N_1640,N_3410);
or U5534 (N_5534,N_3030,N_855);
xnor U5535 (N_5535,N_4988,N_2184);
xnor U5536 (N_5536,N_1824,N_3277);
and U5537 (N_5537,N_4834,N_443);
xnor U5538 (N_5538,N_693,N_1079);
nand U5539 (N_5539,N_244,N_3421);
nand U5540 (N_5540,N_1931,N_297);
or U5541 (N_5541,N_1260,N_30);
xnor U5542 (N_5542,N_4708,N_3310);
and U5543 (N_5543,N_1388,N_4531);
and U5544 (N_5544,N_1821,N_293);
xor U5545 (N_5545,N_2960,N_1610);
xnor U5546 (N_5546,N_4461,N_2630);
or U5547 (N_5547,N_3727,N_1617);
nor U5548 (N_5548,N_2633,N_1268);
nor U5549 (N_5549,N_1549,N_605);
nor U5550 (N_5550,N_283,N_4569);
or U5551 (N_5551,N_2598,N_2562);
and U5552 (N_5552,N_2226,N_1925);
xor U5553 (N_5553,N_3706,N_2070);
nand U5554 (N_5554,N_981,N_692);
and U5555 (N_5555,N_1958,N_2294);
or U5556 (N_5556,N_2003,N_4795);
or U5557 (N_5557,N_1647,N_2329);
nor U5558 (N_5558,N_3989,N_16);
nor U5559 (N_5559,N_4127,N_2858);
and U5560 (N_5560,N_4780,N_1092);
xor U5561 (N_5561,N_4445,N_2904);
nor U5562 (N_5562,N_2270,N_1312);
nand U5563 (N_5563,N_253,N_683);
or U5564 (N_5564,N_4990,N_3994);
xor U5565 (N_5565,N_1205,N_3912);
or U5566 (N_5566,N_1381,N_4530);
or U5567 (N_5567,N_2713,N_4743);
or U5568 (N_5568,N_3937,N_872);
xor U5569 (N_5569,N_1953,N_2304);
nand U5570 (N_5570,N_3286,N_3906);
xor U5571 (N_5571,N_1856,N_3703);
xnor U5572 (N_5572,N_1198,N_1311);
nor U5573 (N_5573,N_2046,N_143);
or U5574 (N_5574,N_4485,N_2985);
nor U5575 (N_5575,N_1115,N_3485);
nand U5576 (N_5576,N_3708,N_4836);
or U5577 (N_5577,N_101,N_568);
nor U5578 (N_5578,N_4698,N_3659);
or U5579 (N_5579,N_4555,N_1608);
nor U5580 (N_5580,N_732,N_2297);
nand U5581 (N_5581,N_704,N_1994);
nand U5582 (N_5582,N_4287,N_430);
nor U5583 (N_5583,N_2108,N_2307);
nor U5584 (N_5584,N_3908,N_230);
or U5585 (N_5585,N_420,N_336);
or U5586 (N_5586,N_2416,N_1630);
xor U5587 (N_5587,N_1932,N_2244);
xnor U5588 (N_5588,N_3701,N_422);
xnor U5589 (N_5589,N_1300,N_2250);
or U5590 (N_5590,N_779,N_2168);
xor U5591 (N_5591,N_3322,N_4841);
xor U5592 (N_5592,N_3846,N_2445);
and U5593 (N_5593,N_846,N_4410);
nor U5594 (N_5594,N_1452,N_2092);
nor U5595 (N_5595,N_1603,N_1175);
nand U5596 (N_5596,N_1048,N_669);
xor U5597 (N_5597,N_1218,N_1912);
and U5598 (N_5598,N_2806,N_2048);
or U5599 (N_5599,N_1385,N_4937);
nor U5600 (N_5600,N_3817,N_3515);
nand U5601 (N_5601,N_4269,N_3984);
and U5602 (N_5602,N_1012,N_3385);
and U5603 (N_5603,N_399,N_2341);
nand U5604 (N_5604,N_4646,N_684);
nor U5605 (N_5605,N_4053,N_1973);
xor U5606 (N_5606,N_1171,N_494);
xnor U5607 (N_5607,N_2066,N_2883);
and U5608 (N_5608,N_1325,N_1182);
xnor U5609 (N_5609,N_2905,N_1504);
or U5610 (N_5610,N_3958,N_4194);
or U5611 (N_5611,N_949,N_1480);
and U5612 (N_5612,N_4902,N_4781);
xnor U5613 (N_5613,N_340,N_2504);
or U5614 (N_5614,N_2582,N_2090);
nor U5615 (N_5615,N_2476,N_857);
xnor U5616 (N_5616,N_4599,N_4537);
nor U5617 (N_5617,N_4311,N_4321);
and U5618 (N_5618,N_3246,N_3272);
xnor U5619 (N_5619,N_3879,N_3715);
or U5620 (N_5620,N_1584,N_648);
nand U5621 (N_5621,N_327,N_74);
nand U5622 (N_5622,N_3820,N_1358);
nor U5623 (N_5623,N_804,N_3631);
xor U5624 (N_5624,N_3574,N_1804);
and U5625 (N_5625,N_1701,N_4960);
nor U5626 (N_5626,N_3059,N_3400);
or U5627 (N_5627,N_1784,N_3253);
nand U5628 (N_5628,N_3334,N_3623);
and U5629 (N_5629,N_3636,N_3993);
nor U5630 (N_5630,N_2192,N_179);
xor U5631 (N_5631,N_1363,N_2069);
xor U5632 (N_5632,N_1082,N_3860);
nand U5633 (N_5633,N_125,N_3364);
nand U5634 (N_5634,N_3532,N_2023);
and U5635 (N_5635,N_4767,N_2952);
xnor U5636 (N_5636,N_1460,N_4203);
nand U5637 (N_5637,N_2575,N_1692);
nand U5638 (N_5638,N_3699,N_2885);
xnor U5639 (N_5639,N_4840,N_959);
nand U5640 (N_5640,N_3048,N_4659);
and U5641 (N_5641,N_2397,N_2933);
and U5642 (N_5642,N_893,N_3407);
xnor U5643 (N_5643,N_1467,N_295);
or U5644 (N_5644,N_4357,N_292);
or U5645 (N_5645,N_3911,N_4590);
and U5646 (N_5646,N_3184,N_4658);
xnor U5647 (N_5647,N_289,N_3567);
xnor U5648 (N_5648,N_3752,N_4452);
or U5649 (N_5649,N_1243,N_4930);
or U5650 (N_5650,N_1626,N_117);
nand U5651 (N_5651,N_4661,N_626);
nor U5652 (N_5652,N_3794,N_2399);
nor U5653 (N_5653,N_2308,N_4288);
and U5654 (N_5654,N_2430,N_1811);
or U5655 (N_5655,N_4893,N_875);
xor U5656 (N_5656,N_1253,N_2993);
nor U5657 (N_5657,N_2201,N_4620);
nor U5658 (N_5658,N_3372,N_4073);
or U5659 (N_5659,N_2647,N_3568);
xnor U5660 (N_5660,N_2639,N_1014);
nand U5661 (N_5661,N_926,N_4482);
and U5662 (N_5662,N_4056,N_4703);
nor U5663 (N_5663,N_768,N_3733);
and U5664 (N_5664,N_3064,N_190);
or U5665 (N_5665,N_1194,N_3808);
xnor U5666 (N_5666,N_1076,N_4270);
or U5667 (N_5667,N_1892,N_512);
xor U5668 (N_5668,N_2928,N_1145);
and U5669 (N_5669,N_1997,N_2195);
and U5670 (N_5670,N_1331,N_2596);
and U5671 (N_5671,N_4733,N_80);
or U5672 (N_5672,N_2875,N_1880);
nor U5673 (N_5673,N_2296,N_3088);
or U5674 (N_5674,N_2449,N_2794);
nor U5675 (N_5675,N_1080,N_2510);
and U5676 (N_5676,N_1127,N_3423);
or U5677 (N_5677,N_4272,N_3883);
xor U5678 (N_5678,N_3656,N_3210);
nor U5679 (N_5679,N_577,N_3113);
xor U5680 (N_5680,N_1991,N_1296);
nand U5681 (N_5681,N_4887,N_2551);
xnor U5682 (N_5682,N_2606,N_2964);
nor U5683 (N_5683,N_2310,N_2829);
xor U5684 (N_5684,N_172,N_4758);
nor U5685 (N_5685,N_4496,N_1807);
and U5686 (N_5686,N_711,N_7);
nand U5687 (N_5687,N_482,N_1089);
nor U5688 (N_5688,N_3424,N_2130);
or U5689 (N_5689,N_28,N_3995);
nand U5690 (N_5690,N_2651,N_1384);
xnor U5691 (N_5691,N_1843,N_1665);
or U5692 (N_5692,N_2900,N_4276);
and U5693 (N_5693,N_72,N_4944);
nor U5694 (N_5694,N_1666,N_452);
xnor U5695 (N_5695,N_706,N_3836);
xor U5696 (N_5696,N_2164,N_4094);
or U5697 (N_5697,N_3156,N_4005);
or U5698 (N_5698,N_3443,N_4097);
nand U5699 (N_5699,N_912,N_1270);
or U5700 (N_5700,N_539,N_4379);
or U5701 (N_5701,N_2275,N_1620);
nand U5702 (N_5702,N_3546,N_2519);
or U5703 (N_5703,N_4629,N_3283);
nand U5704 (N_5704,N_2313,N_1471);
or U5705 (N_5705,N_1634,N_2518);
xor U5706 (N_5706,N_4100,N_3302);
or U5707 (N_5707,N_161,N_290);
xnor U5708 (N_5708,N_1364,N_911);
nand U5709 (N_5709,N_4280,N_2635);
and U5710 (N_5710,N_1411,N_3106);
nor U5711 (N_5711,N_1403,N_2980);
nor U5712 (N_5712,N_1441,N_4885);
nor U5713 (N_5713,N_3942,N_3503);
or U5714 (N_5714,N_1158,N_4760);
xor U5715 (N_5715,N_2141,N_1543);
xnor U5716 (N_5716,N_1762,N_1002);
nor U5717 (N_5717,N_4063,N_266);
xnor U5718 (N_5718,N_3381,N_4936);
xnor U5719 (N_5719,N_2259,N_4507);
xor U5720 (N_5720,N_1551,N_2102);
nand U5721 (N_5721,N_264,N_2693);
or U5722 (N_5722,N_1204,N_4322);
xnor U5723 (N_5723,N_374,N_3208);
and U5724 (N_5724,N_4650,N_2255);
and U5725 (N_5725,N_4278,N_373);
nor U5726 (N_5726,N_556,N_1533);
nand U5727 (N_5727,N_384,N_3481);
nor U5728 (N_5728,N_1122,N_3042);
and U5729 (N_5729,N_1050,N_1968);
and U5730 (N_5730,N_4712,N_2841);
nand U5731 (N_5731,N_1820,N_164);
nor U5732 (N_5732,N_3775,N_785);
nand U5733 (N_5733,N_1287,N_4156);
and U5734 (N_5734,N_2677,N_4479);
xor U5735 (N_5735,N_2560,N_924);
and U5736 (N_5736,N_1308,N_3095);
xnor U5737 (N_5737,N_4906,N_1464);
or U5738 (N_5738,N_4736,N_4969);
xnor U5739 (N_5739,N_203,N_1516);
nand U5740 (N_5740,N_149,N_4597);
or U5741 (N_5741,N_4090,N_4921);
nand U5742 (N_5742,N_4041,N_930);
nor U5743 (N_5743,N_4763,N_3401);
xor U5744 (N_5744,N_1636,N_805);
nor U5745 (N_5745,N_4394,N_3455);
xor U5746 (N_5746,N_237,N_102);
nand U5747 (N_5747,N_3348,N_1598);
and U5748 (N_5748,N_2301,N_3542);
and U5749 (N_5749,N_712,N_3335);
xor U5750 (N_5750,N_2120,N_4714);
xnor U5751 (N_5751,N_769,N_1408);
nor U5752 (N_5752,N_3540,N_471);
or U5753 (N_5753,N_1901,N_4084);
nand U5754 (N_5754,N_3521,N_4257);
nor U5755 (N_5755,N_827,N_564);
xnor U5756 (N_5756,N_2687,N_3280);
xnor U5757 (N_5757,N_1098,N_1280);
nor U5758 (N_5758,N_2863,N_1075);
or U5759 (N_5759,N_4213,N_1009);
or U5760 (N_5760,N_3773,N_4550);
or U5761 (N_5761,N_1726,N_210);
and U5762 (N_5762,N_2407,N_2387);
and U5763 (N_5763,N_1920,N_1611);
nor U5764 (N_5764,N_2745,N_1771);
and U5765 (N_5765,N_3966,N_1225);
xnor U5766 (N_5766,N_3632,N_489);
xor U5767 (N_5767,N_2736,N_124);
or U5768 (N_5768,N_2634,N_1314);
xnor U5769 (N_5769,N_4705,N_3711);
and U5770 (N_5770,N_4375,N_79);
xnor U5771 (N_5771,N_2665,N_2236);
nor U5772 (N_5772,N_2059,N_1370);
nand U5773 (N_5773,N_4635,N_437);
nand U5774 (N_5774,N_4997,N_4249);
or U5775 (N_5775,N_181,N_1004);
xor U5776 (N_5776,N_98,N_2319);
nand U5777 (N_5777,N_2087,N_1147);
xnor U5778 (N_5778,N_4150,N_3129);
xor U5779 (N_5779,N_3670,N_4575);
and U5780 (N_5780,N_3642,N_459);
xor U5781 (N_5781,N_4333,N_62);
nand U5782 (N_5782,N_820,N_3158);
xor U5783 (N_5783,N_424,N_2112);
nand U5784 (N_5784,N_1768,N_235);
or U5785 (N_5785,N_4465,N_3530);
nor U5786 (N_5786,N_1687,N_4049);
nor U5787 (N_5787,N_3451,N_860);
or U5788 (N_5788,N_824,N_1532);
or U5789 (N_5789,N_3565,N_1796);
nand U5790 (N_5790,N_1000,N_3183);
or U5791 (N_5791,N_1209,N_4294);
xor U5792 (N_5792,N_3247,N_881);
or U5793 (N_5793,N_3190,N_2110);
nor U5794 (N_5794,N_2116,N_2740);
nand U5795 (N_5795,N_925,N_3533);
or U5796 (N_5796,N_4592,N_1719);
xor U5797 (N_5797,N_4437,N_1854);
nor U5798 (N_5798,N_610,N_1152);
nand U5799 (N_5799,N_640,N_4459);
and U5800 (N_5800,N_337,N_454);
and U5801 (N_5801,N_4724,N_2177);
nand U5802 (N_5802,N_4171,N_2178);
nor U5803 (N_5803,N_4602,N_1442);
or U5804 (N_5804,N_2515,N_2146);
xor U5805 (N_5805,N_1760,N_4614);
xnor U5806 (N_5806,N_3186,N_4493);
xnor U5807 (N_5807,N_3603,N_1993);
nor U5808 (N_5808,N_144,N_583);
and U5809 (N_5809,N_404,N_1561);
nor U5810 (N_5810,N_4667,N_1574);
or U5811 (N_5811,N_254,N_173);
nor U5812 (N_5812,N_247,N_2414);
or U5813 (N_5813,N_2167,N_4776);
and U5814 (N_5814,N_604,N_729);
and U5815 (N_5815,N_3893,N_3558);
nor U5816 (N_5816,N_4681,N_4679);
or U5817 (N_5817,N_2523,N_3512);
xnor U5818 (N_5818,N_401,N_1064);
nor U5819 (N_5819,N_3605,N_1136);
nor U5820 (N_5820,N_2759,N_1624);
nand U5821 (N_5821,N_4366,N_1715);
nand U5822 (N_5822,N_1303,N_4354);
and U5823 (N_5823,N_1798,N_551);
and U5824 (N_5824,N_3977,N_3791);
xnor U5825 (N_5825,N_1926,N_939);
xnor U5826 (N_5826,N_2717,N_1397);
and U5827 (N_5827,N_3309,N_4143);
nand U5828 (N_5828,N_537,N_3573);
or U5829 (N_5829,N_3827,N_4125);
nor U5830 (N_5830,N_847,N_4199);
and U5831 (N_5831,N_2248,N_1250);
nor U5832 (N_5832,N_1367,N_2455);
and U5833 (N_5833,N_4253,N_905);
xor U5834 (N_5834,N_3215,N_4421);
nand U5835 (N_5835,N_1736,N_3391);
nor U5836 (N_5836,N_2932,N_717);
xnor U5837 (N_5837,N_68,N_3976);
nor U5838 (N_5838,N_1424,N_4924);
or U5839 (N_5839,N_1326,N_2330);
nor U5840 (N_5840,N_4859,N_4922);
or U5841 (N_5841,N_265,N_1541);
xor U5842 (N_5842,N_4409,N_1081);
nand U5843 (N_5843,N_389,N_2942);
or U5844 (N_5844,N_128,N_123);
or U5845 (N_5845,N_3316,N_447);
nor U5846 (N_5846,N_596,N_1714);
nor U5847 (N_5847,N_1540,N_627);
nand U5848 (N_5848,N_207,N_1455);
xnor U5849 (N_5849,N_1765,N_2500);
and U5850 (N_5850,N_2958,N_744);
nand U5851 (N_5851,N_3000,N_4225);
or U5852 (N_5852,N_191,N_4219);
or U5853 (N_5853,N_4170,N_3923);
or U5854 (N_5854,N_4654,N_2957);
xor U5855 (N_5855,N_4709,N_1724);
xnor U5856 (N_5856,N_4506,N_1847);
or U5857 (N_5857,N_2592,N_1930);
nand U5858 (N_5858,N_4356,N_2224);
and U5859 (N_5859,N_201,N_2072);
nor U5860 (N_5860,N_2429,N_2615);
and U5861 (N_5861,N_4416,N_2354);
and U5862 (N_5862,N_2767,N_441);
or U5863 (N_5863,N_2381,N_2862);
and U5864 (N_5864,N_3273,N_4907);
or U5865 (N_5865,N_345,N_3288);
nand U5866 (N_5866,N_4672,N_651);
or U5867 (N_5867,N_4033,N_3837);
xnor U5868 (N_5868,N_4325,N_4860);
nor U5869 (N_5869,N_2380,N_3119);
and U5870 (N_5870,N_3903,N_3362);
nand U5871 (N_5871,N_4638,N_1895);
or U5872 (N_5872,N_567,N_1852);
nor U5873 (N_5873,N_2133,N_1619);
nor U5874 (N_5874,N_3413,N_3209);
or U5875 (N_5875,N_525,N_4959);
nand U5876 (N_5876,N_3163,N_4552);
nor U5877 (N_5877,N_1891,N_742);
xor U5878 (N_5878,N_2373,N_1333);
nor U5879 (N_5879,N_2186,N_379);
or U5880 (N_5880,N_4293,N_316);
and U5881 (N_5881,N_1708,N_3452);
and U5882 (N_5882,N_3563,N_2716);
and U5883 (N_5883,N_3380,N_3463);
nand U5884 (N_5884,N_11,N_4142);
nand U5885 (N_5885,N_1477,N_3502);
or U5886 (N_5886,N_4792,N_2545);
nand U5887 (N_5887,N_2601,N_3918);
xnor U5888 (N_5888,N_4300,N_1834);
and U5889 (N_5889,N_2943,N_3647);
nand U5890 (N_5890,N_1380,N_1164);
xor U5891 (N_5891,N_1172,N_3617);
nand U5892 (N_5892,N_1870,N_2919);
xor U5893 (N_5893,N_171,N_2285);
and U5894 (N_5894,N_677,N_966);
nand U5895 (N_5895,N_4108,N_4762);
xor U5896 (N_5896,N_3925,N_3963);
xnor U5897 (N_5897,N_783,N_4994);
and U5898 (N_5898,N_4516,N_3662);
and U5899 (N_5899,N_2784,N_2212);
xnor U5900 (N_5900,N_1913,N_4241);
or U5901 (N_5901,N_3528,N_3241);
xor U5902 (N_5902,N_660,N_800);
xor U5903 (N_5903,N_4621,N_1606);
nand U5904 (N_5904,N_2425,N_2969);
or U5905 (N_5905,N_4006,N_2008);
and U5906 (N_5906,N_29,N_1534);
nand U5907 (N_5907,N_2962,N_2303);
nor U5908 (N_5908,N_4669,N_4012);
nand U5909 (N_5909,N_4317,N_3606);
or U5910 (N_5910,N_2331,N_1227);
nand U5911 (N_5911,N_1188,N_2584);
or U5912 (N_5912,N_4789,N_2770);
and U5913 (N_5913,N_953,N_561);
nor U5914 (N_5914,N_4611,N_3796);
or U5915 (N_5915,N_2696,N_955);
nor U5916 (N_5916,N_3028,N_1585);
or U5917 (N_5917,N_4983,N_2550);
and U5918 (N_5918,N_274,N_810);
nand U5919 (N_5919,N_1239,N_25);
nor U5920 (N_5920,N_4226,N_3039);
nand U5921 (N_5921,N_1459,N_650);
or U5922 (N_5922,N_1097,N_4847);
nand U5923 (N_5923,N_2602,N_4092);
nand U5924 (N_5924,N_707,N_47);
xor U5925 (N_5925,N_2043,N_4568);
xnor U5926 (N_5926,N_3767,N_2139);
xnor U5927 (N_5927,N_1799,N_3109);
or U5928 (N_5928,N_4803,N_1042);
nand U5929 (N_5929,N_1947,N_4453);
nand U5930 (N_5930,N_3019,N_4918);
and U5931 (N_5931,N_3324,N_2395);
nor U5932 (N_5932,N_4533,N_1544);
nor U5933 (N_5933,N_3014,N_1374);
nor U5934 (N_5934,N_1445,N_1663);
or U5935 (N_5935,N_13,N_1463);
nor U5936 (N_5936,N_3366,N_4216);
nand U5937 (N_5937,N_3332,N_1943);
nor U5938 (N_5938,N_58,N_1394);
or U5939 (N_5939,N_3227,N_1631);
nand U5940 (N_5940,N_3723,N_2413);
and U5941 (N_5941,N_406,N_2626);
or U5942 (N_5942,N_2095,N_1248);
xor U5943 (N_5943,N_2036,N_1406);
nor U5944 (N_5944,N_67,N_3360);
nand U5945 (N_5945,N_4849,N_1271);
nand U5946 (N_5946,N_3198,N_341);
xor U5947 (N_5947,N_3054,N_4239);
and U5948 (N_5948,N_2377,N_37);
or U5949 (N_5949,N_3356,N_3904);
xnor U5950 (N_5950,N_3081,N_665);
nand U5951 (N_5951,N_845,N_3757);
or U5952 (N_5952,N_3639,N_4047);
and U5953 (N_5953,N_2923,N_4809);
or U5954 (N_5954,N_1220,N_4343);
or U5955 (N_5955,N_999,N_1444);
xor U5956 (N_5956,N_4591,N_4943);
nand U5957 (N_5957,N_2338,N_1219);
or U5958 (N_5958,N_1517,N_1972);
or U5959 (N_5959,N_2968,N_2809);
xor U5960 (N_5960,N_4064,N_947);
or U5961 (N_5961,N_1328,N_464);
xor U5962 (N_5962,N_2656,N_2147);
or U5963 (N_5963,N_425,N_3350);
and U5964 (N_5964,N_3930,N_4096);
nor U5965 (N_5965,N_3318,N_227);
and U5966 (N_5966,N_4024,N_3592);
and U5967 (N_5967,N_823,N_3777);
xor U5968 (N_5968,N_784,N_411);
nor U5969 (N_5969,N_965,N_1808);
or U5970 (N_5970,N_1961,N_3327);
nor U5971 (N_5971,N_1320,N_4987);
and U5972 (N_5972,N_2438,N_56);
nand U5973 (N_5973,N_513,N_1566);
or U5974 (N_5974,N_1948,N_2034);
nand U5975 (N_5975,N_1310,N_1429);
nor U5976 (N_5976,N_486,N_1577);
xor U5977 (N_5977,N_2305,N_3795);
or U5978 (N_5978,N_4061,N_4013);
xor U5979 (N_5979,N_1102,N_3406);
nand U5980 (N_5980,N_4083,N_2981);
and U5981 (N_5981,N_2064,N_819);
and U5982 (N_5982,N_229,N_4222);
xor U5983 (N_5983,N_3200,N_3477);
and U5984 (N_5984,N_1816,N_808);
xnor U5985 (N_5985,N_3453,N_205);
xnor U5986 (N_5986,N_1521,N_968);
and U5987 (N_5987,N_3430,N_4016);
xnor U5988 (N_5988,N_3127,N_2768);
xnor U5989 (N_5989,N_1981,N_4159);
xnor U5990 (N_5990,N_2393,N_2056);
xnor U5991 (N_5991,N_3790,N_3093);
or U5992 (N_5992,N_897,N_1481);
xnor U5993 (N_5993,N_2511,N_1898);
nor U5994 (N_5994,N_585,N_4524);
and U5995 (N_5995,N_2874,N_3638);
xnor U5996 (N_5996,N_906,N_1165);
and U5997 (N_5997,N_377,N_1565);
nor U5998 (N_5998,N_601,N_1393);
and U5999 (N_5999,N_1857,N_4950);
nor U6000 (N_6000,N_176,N_4631);
xor U6001 (N_6001,N_3743,N_3742);
and U6002 (N_6002,N_1995,N_4292);
and U6003 (N_6003,N_332,N_4051);
and U6004 (N_6004,N_2619,N_116);
nand U6005 (N_6005,N_2045,N_3123);
xor U6006 (N_6006,N_2625,N_3049);
nor U6007 (N_6007,N_3627,N_4754);
and U6008 (N_6008,N_3321,N_4209);
nand U6009 (N_6009,N_1742,N_2127);
nand U6010 (N_6010,N_1185,N_2060);
and U6011 (N_6011,N_1623,N_2282);
nor U6012 (N_6012,N_2921,N_3301);
nand U6013 (N_6013,N_4915,N_405);
nand U6014 (N_6014,N_589,N_3010);
nor U6015 (N_6015,N_2081,N_3328);
nand U6016 (N_6016,N_2664,N_4598);
nor U6017 (N_6017,N_2336,N_1656);
nand U6018 (N_6018,N_2079,N_4057);
and U6019 (N_6019,N_2627,N_133);
nor U6020 (N_6020,N_323,N_3799);
xor U6021 (N_6021,N_2089,N_2419);
and U6022 (N_6022,N_3671,N_3191);
and U6023 (N_6023,N_1114,N_4320);
and U6024 (N_6024,N_609,N_4929);
or U6025 (N_6025,N_3390,N_789);
nand U6026 (N_6026,N_1450,N_1479);
nor U6027 (N_6027,N_2175,N_1772);
nand U6028 (N_6028,N_1963,N_1591);
and U6029 (N_6029,N_1527,N_2378);
or U6030 (N_6030,N_348,N_233);
or U6031 (N_6031,N_4438,N_918);
nor U6032 (N_6032,N_433,N_2753);
and U6033 (N_6033,N_2295,N_4135);
and U6034 (N_6034,N_3907,N_1660);
xnor U6035 (N_6035,N_3895,N_3025);
nor U6036 (N_6036,N_3078,N_752);
nor U6037 (N_6037,N_4748,N_2738);
and U6038 (N_6038,N_2391,N_1143);
or U6039 (N_6039,N_4971,N_1106);
xnor U6040 (N_6040,N_4387,N_3842);
xnor U6041 (N_6041,N_1879,N_4373);
and U6042 (N_6042,N_412,N_3744);
or U6043 (N_6043,N_66,N_2281);
xor U6044 (N_6044,N_1996,N_1693);
or U6045 (N_6045,N_2555,N_3212);
nor U6046 (N_6046,N_4977,N_4008);
xor U6047 (N_6047,N_2140,N_4275);
and U6048 (N_6048,N_2375,N_1690);
or U6049 (N_6049,N_4381,N_2613);
xnor U6050 (N_6050,N_4713,N_1838);
nor U6051 (N_6051,N_2931,N_2487);
nor U6052 (N_6052,N_3175,N_4914);
nand U6053 (N_6053,N_3890,N_3566);
nor U6054 (N_6054,N_2731,N_759);
and U6055 (N_6055,N_2684,N_376);
xor U6056 (N_6056,N_4001,N_1612);
nand U6057 (N_6057,N_4534,N_2741);
or U6058 (N_6058,N_132,N_4586);
and U6059 (N_6059,N_593,N_1091);
nor U6060 (N_6060,N_3822,N_1245);
or U6061 (N_6061,N_538,N_3342);
and U6062 (N_6062,N_1902,N_3278);
or U6063 (N_6063,N_2463,N_4900);
or U6064 (N_6064,N_3022,N_3717);
nand U6065 (N_6065,N_279,N_4264);
xor U6066 (N_6066,N_84,N_4819);
or U6067 (N_6067,N_3760,N_3978);
nand U6068 (N_6068,N_3192,N_4116);
or U6069 (N_6069,N_990,N_1330);
nor U6070 (N_6070,N_4232,N_3221);
or U6071 (N_6071,N_2257,N_4483);
xor U6072 (N_6072,N_3040,N_188);
nor U6073 (N_6073,N_1392,N_3143);
nor U6074 (N_6074,N_1077,N_2062);
or U6075 (N_6075,N_2836,N_1507);
nand U6076 (N_6076,N_1244,N_2118);
nor U6077 (N_6077,N_3387,N_2027);
xor U6078 (N_6078,N_962,N_55);
or U6079 (N_6079,N_4835,N_3905);
and U6080 (N_6080,N_338,N_2335);
nor U6081 (N_6081,N_4640,N_1419);
nand U6082 (N_6082,N_1117,N_4201);
and U6083 (N_6083,N_1159,N_3824);
nand U6084 (N_6084,N_2945,N_870);
nand U6085 (N_6085,N_3260,N_2718);
xnor U6086 (N_6086,N_1600,N_4214);
or U6087 (N_6087,N_1794,N_1399);
or U6088 (N_6088,N_1992,N_2111);
nor U6089 (N_6089,N_1155,N_3932);
nand U6090 (N_6090,N_3866,N_4290);
xor U6091 (N_6091,N_1023,N_4837);
and U6092 (N_6092,N_1448,N_988);
nor U6093 (N_6093,N_4377,N_3069);
nor U6094 (N_6094,N_3776,N_2578);
nor U6095 (N_6095,N_3536,N_3725);
or U6096 (N_6096,N_4152,N_1342);
and U6097 (N_6097,N_2591,N_690);
nor U6098 (N_6098,N_2795,N_4347);
nand U6099 (N_6099,N_4940,N_2642);
nand U6100 (N_6100,N_61,N_3829);
and U6101 (N_6101,N_535,N_1519);
and U6102 (N_6102,N_2320,N_3974);
xor U6103 (N_6103,N_835,N_617);
or U6104 (N_6104,N_1327,N_3496);
nand U6105 (N_6105,N_571,N_4161);
nand U6106 (N_6106,N_1900,N_956);
nand U6107 (N_6107,N_4242,N_573);
and U6108 (N_6108,N_3480,N_3177);
xnor U6109 (N_6109,N_3861,N_1226);
nand U6110 (N_6110,N_4165,N_4865);
nor U6111 (N_6111,N_75,N_3856);
xnor U6112 (N_6112,N_2938,N_523);
xnor U6113 (N_6113,N_4215,N_3847);
and U6114 (N_6114,N_4798,N_1909);
and U6115 (N_6115,N_1658,N_644);
nand U6116 (N_6116,N_3672,N_365);
or U6117 (N_6117,N_3803,N_2996);
xor U6118 (N_6118,N_1286,N_2754);
or U6119 (N_6119,N_2050,N_3082);
and U6120 (N_6120,N_1231,N_3658);
xnor U6121 (N_6121,N_2527,N_2972);
nand U6122 (N_6122,N_1008,N_2970);
nand U6123 (N_6123,N_1965,N_4808);
and U6124 (N_6124,N_4337,N_4535);
xnor U6125 (N_6125,N_1319,N_3864);
nand U6126 (N_6126,N_3850,N_2828);
xnor U6127 (N_6127,N_4134,N_2506);
nor U6128 (N_6128,N_3058,N_3099);
xor U6129 (N_6129,N_1740,N_3493);
xnor U6130 (N_6130,N_3418,N_2871);
nor U6131 (N_6131,N_17,N_2453);
or U6132 (N_6132,N_1934,N_4812);
nor U6133 (N_6133,N_3595,N_4618);
nor U6134 (N_6134,N_2547,N_3741);
xor U6135 (N_6135,N_4580,N_2723);
and U6136 (N_6136,N_2889,N_4625);
and U6137 (N_6137,N_1637,N_3179);
or U6138 (N_6138,N_1570,N_1011);
xor U6139 (N_6139,N_493,N_3018);
nand U6140 (N_6140,N_2269,N_3229);
nand U6141 (N_6141,N_4949,N_4406);
or U6142 (N_6142,N_326,N_4107);
xnor U6143 (N_6143,N_4329,N_2279);
or U6144 (N_6144,N_299,N_286);
xnor U6145 (N_6145,N_1675,N_1396);
and U6146 (N_6146,N_4349,N_780);
and U6147 (N_6147,N_3486,N_3464);
xnor U6148 (N_6148,N_4020,N_2165);
nor U6149 (N_6149,N_674,N_246);
nand U6150 (N_6150,N_4974,N_350);
xor U6151 (N_6151,N_4440,N_3909);
and U6152 (N_6152,N_3919,N_2896);
xnor U6153 (N_6153,N_3559,N_2080);
or U6154 (N_6154,N_2435,N_3358);
nand U6155 (N_6155,N_1289,N_3239);
and U6156 (N_6156,N_4467,N_1756);
or U6157 (N_6157,N_4876,N_1193);
or U6158 (N_6158,N_1181,N_3669);
and U6159 (N_6159,N_504,N_4478);
xor U6160 (N_6160,N_3312,N_3975);
or U6161 (N_6161,N_1309,N_3740);
and U6162 (N_6162,N_4946,N_2918);
and U6163 (N_6163,N_1645,N_3873);
and U6164 (N_6164,N_3017,N_4831);
nor U6165 (N_6165,N_4657,N_4610);
xnor U6166 (N_6166,N_740,N_3053);
nor U6167 (N_6167,N_3061,N_3949);
or U6168 (N_6168,N_1514,N_4022);
or U6169 (N_6169,N_653,N_1672);
and U6170 (N_6170,N_343,N_18);
and U6171 (N_6171,N_3388,N_4471);
nand U6172 (N_6172,N_899,N_1629);
nor U6173 (N_6173,N_4768,N_2915);
nor U6174 (N_6174,N_3352,N_6);
nor U6175 (N_6175,N_2688,N_3577);
or U6176 (N_6176,N_3498,N_3347);
nor U6177 (N_6177,N_4821,N_1644);
nor U6178 (N_6178,N_4369,N_4870);
or U6179 (N_6179,N_3749,N_3118);
nand U6180 (N_6180,N_3539,N_1747);
nor U6181 (N_6181,N_1166,N_4744);
nand U6182 (N_6182,N_352,N_3751);
and U6183 (N_6183,N_4355,N_3382);
or U6184 (N_6184,N_4119,N_743);
xor U6185 (N_6185,N_1599,N_1918);
or U6186 (N_6186,N_2992,N_2252);
and U6187 (N_6187,N_238,N_689);
nor U6188 (N_6188,N_2715,N_4927);
nor U6189 (N_6189,N_409,N_2574);
xor U6190 (N_6190,N_2755,N_3306);
nand U6191 (N_6191,N_4746,N_3234);
and U6192 (N_6192,N_4481,N_4085);
xor U6193 (N_6193,N_1685,N_1988);
and U6194 (N_6194,N_1356,N_1970);
xnor U6195 (N_6195,N_4556,N_1251);
or U6196 (N_6196,N_3405,N_682);
nand U6197 (N_6197,N_2115,N_806);
or U6198 (N_6198,N_4023,N_1086);
nand U6199 (N_6199,N_1986,N_4701);
nand U6200 (N_6200,N_4985,N_40);
or U6201 (N_6201,N_2810,N_1935);
or U6202 (N_6202,N_4368,N_1639);
nor U6203 (N_6203,N_1118,N_3148);
xnor U6204 (N_6204,N_709,N_4032);
nor U6205 (N_6205,N_388,N_2222);
and U6206 (N_6206,N_1203,N_2655);
nand U6207 (N_6207,N_974,N_4301);
and U6208 (N_6208,N_1140,N_3931);
and U6209 (N_6209,N_3980,N_262);
nand U6210 (N_6210,N_2789,N_1052);
or U6211 (N_6211,N_2866,N_878);
and U6212 (N_6212,N_2719,N_105);
nor U6213 (N_6213,N_863,N_2489);
xnor U6214 (N_6214,N_1557,N_2470);
or U6215 (N_6215,N_3080,N_2359);
nand U6216 (N_6216,N_719,N_2564);
and U6217 (N_6217,N_3663,N_2747);
xor U6218 (N_6218,N_3415,N_4462);
xor U6219 (N_6219,N_3202,N_1100);
nor U6220 (N_6220,N_342,N_1094);
and U6221 (N_6221,N_480,N_97);
and U6222 (N_6222,N_2844,N_3284);
nor U6223 (N_6223,N_1916,N_1801);
nor U6224 (N_6224,N_2318,N_2622);
and U6225 (N_6225,N_4751,N_666);
and U6226 (N_6226,N_4188,N_3155);
nor U6227 (N_6227,N_1744,N_1292);
nand U6228 (N_6228,N_1526,N_1007);
and U6229 (N_6229,N_1556,N_2565);
xnor U6230 (N_6230,N_2049,N_1595);
xor U6231 (N_6231,N_4227,N_1252);
nor U6232 (N_6232,N_220,N_1906);
and U6233 (N_6233,N_51,N_42);
and U6234 (N_6234,N_900,N_78);
nand U6235 (N_6235,N_972,N_1713);
nor U6236 (N_6236,N_2983,N_2392);
nand U6237 (N_6237,N_31,N_1046);
xnor U6238 (N_6238,N_4765,N_1180);
or U6239 (N_6239,N_3428,N_3461);
or U6240 (N_6240,N_4185,N_4600);
or U6241 (N_6241,N_3094,N_449);
xnor U6242 (N_6242,N_1461,N_3047);
and U6243 (N_6243,N_2721,N_4896);
or U6244 (N_6244,N_1390,N_1501);
xor U6245 (N_6245,N_2104,N_1956);
xnor U6246 (N_6246,N_2121,N_588);
and U6247 (N_6247,N_3244,N_3548);
or U6248 (N_6248,N_3396,N_2971);
and U6249 (N_6249,N_1835,N_4680);
nor U6250 (N_6250,N_1283,N_381);
and U6251 (N_6251,N_4509,N_3472);
and U6252 (N_6252,N_1635,N_122);
or U6253 (N_6253,N_19,N_3437);
xnor U6254 (N_6254,N_1782,N_2076);
and U6255 (N_6255,N_4395,N_2843);
nand U6256 (N_6256,N_1613,N_2605);
or U6257 (N_6257,N_3641,N_4879);
nand U6258 (N_6258,N_1542,N_2792);
or U6259 (N_6259,N_1764,N_1111);
and U6260 (N_6260,N_1124,N_994);
nor U6261 (N_6261,N_4197,N_3237);
and U6262 (N_6262,N_2211,N_3138);
and U6263 (N_6263,N_4542,N_737);
xnor U6264 (N_6264,N_4539,N_3887);
and U6265 (N_6265,N_3609,N_402);
and U6266 (N_6266,N_1281,N_2143);
and U6267 (N_6267,N_1646,N_85);
nor U6268 (N_6268,N_3403,N_3913);
or U6269 (N_6269,N_3416,N_515);
or U6270 (N_6270,N_417,N_834);
nor U6271 (N_6271,N_2166,N_2361);
xor U6272 (N_6272,N_1413,N_2681);
xor U6273 (N_6273,N_2763,N_1029);
or U6274 (N_6274,N_2106,N_2382);
nor U6275 (N_6275,N_2852,N_3131);
nand U6276 (N_6276,N_4505,N_4026);
and U6277 (N_6277,N_4588,N_4433);
and U6278 (N_6278,N_3511,N_4570);
xnor U6279 (N_6279,N_3834,N_3629);
and U6280 (N_6280,N_4666,N_1582);
or U6281 (N_6281,N_2756,N_127);
and U6282 (N_6282,N_3786,N_1160);
or U6283 (N_6283,N_2013,N_4543);
nand U6284 (N_6284,N_1775,N_882);
or U6285 (N_6285,N_3997,N_1732);
and U6286 (N_6286,N_2760,N_811);
and U6287 (N_6287,N_1525,N_3470);
nor U6288 (N_6288,N_2873,N_1841);
xnor U6289 (N_6289,N_70,N_4067);
nand U6290 (N_6290,N_4393,N_2456);
nor U6291 (N_6291,N_3170,N_3588);
or U6292 (N_6292,N_3223,N_1839);
or U6293 (N_6293,N_4055,N_4526);
xor U6294 (N_6294,N_3001,N_509);
or U6295 (N_6295,N_2948,N_3365);
xor U6296 (N_6296,N_4195,N_2071);
or U6297 (N_6297,N_3680,N_46);
or U6298 (N_6298,N_1831,N_2998);
xor U6299 (N_6299,N_2007,N_2895);
or U6300 (N_6300,N_1341,N_4972);
xnor U6301 (N_6301,N_3043,N_2474);
and U6302 (N_6302,N_24,N_543);
xor U6303 (N_6303,N_522,N_3299);
or U6304 (N_6304,N_667,N_23);
nand U6305 (N_6305,N_3303,N_414);
nor U6306 (N_6306,N_521,N_4514);
nand U6307 (N_6307,N_2247,N_2906);
nor U6308 (N_6308,N_3435,N_4361);
or U6309 (N_6309,N_2907,N_1921);
xor U6310 (N_6310,N_2075,N_4205);
or U6311 (N_6311,N_2798,N_658);
nand U6312 (N_6312,N_1425,N_1651);
nand U6313 (N_6313,N_408,N_967);
xnor U6314 (N_6314,N_3630,N_136);
nand U6315 (N_6315,N_3878,N_3998);
xor U6316 (N_6316,N_2367,N_470);
nor U6317 (N_6317,N_841,N_3487);
xor U6318 (N_6318,N_4075,N_598);
nor U6319 (N_6319,N_275,N_3865);
nor U6320 (N_6320,N_672,N_4596);
and U6321 (N_6321,N_2239,N_2710);
or U6322 (N_6322,N_873,N_1511);
or U6323 (N_6323,N_2667,N_4574);
and U6324 (N_6324,N_169,N_2058);
or U6325 (N_6325,N_4934,N_4674);
nor U6326 (N_6326,N_3813,N_1379);
nand U6327 (N_6327,N_467,N_3643);
nor U6328 (N_6328,N_3823,N_1391);
nor U6329 (N_6329,N_3439,N_4002);
or U6330 (N_6330,N_4652,N_4686);
or U6331 (N_6331,N_4545,N_1088);
or U6332 (N_6332,N_4380,N_3304);
and U6333 (N_6333,N_557,N_1655);
nand U6334 (N_6334,N_2537,N_3178);
or U6335 (N_6335,N_2219,N_2371);
nand U6336 (N_6336,N_3859,N_4423);
and U6337 (N_6337,N_3780,N_1586);
and U6338 (N_6338,N_2363,N_2749);
and U6339 (N_6339,N_385,N_909);
xor U6340 (N_6340,N_3444,N_736);
xnor U6341 (N_6341,N_1258,N_278);
and U6342 (N_6342,N_2818,N_694);
nand U6343 (N_6343,N_2163,N_200);
or U6344 (N_6344,N_2685,N_3002);
nor U6345 (N_6345,N_2799,N_386);
xnor U6346 (N_6346,N_2877,N_2035);
nor U6347 (N_6347,N_2346,N_65);
xnor U6348 (N_6348,N_2976,N_3816);
nor U6349 (N_6349,N_1497,N_4121);
nor U6350 (N_6350,N_1107,N_4274);
nor U6351 (N_6351,N_4897,N_876);
nor U6352 (N_6352,N_4117,N_1138);
and U6353 (N_6353,N_4220,N_3136);
or U6354 (N_6354,N_378,N_4065);
and U6355 (N_6355,N_4899,N_3934);
or U6356 (N_6356,N_3447,N_481);
and U6357 (N_6357,N_457,N_1053);
or U6358 (N_6358,N_1814,N_4553);
and U6359 (N_6359,N_1416,N_1402);
nor U6360 (N_6360,N_3267,N_3863);
nor U6361 (N_6361,N_4019,N_3874);
or U6362 (N_6362,N_2324,N_3379);
xnor U6363 (N_6363,N_2679,N_2888);
or U6364 (N_6364,N_4086,N_2524);
nor U6365 (N_6365,N_572,N_3120);
nor U6366 (N_6366,N_3852,N_3973);
xor U6367 (N_6367,N_4933,N_4965);
xor U6368 (N_6368,N_3894,N_403);
nand U6369 (N_6369,N_4391,N_4519);
xnor U6370 (N_6370,N_319,N_3805);
nand U6371 (N_6371,N_4265,N_3844);
nand U6372 (N_6372,N_356,N_245);
xor U6373 (N_6373,N_4139,N_4345);
or U6374 (N_6374,N_3230,N_3491);
nor U6375 (N_6375,N_2899,N_2029);
nor U6376 (N_6376,N_1112,N_3274);
and U6377 (N_6377,N_4563,N_4794);
xor U6378 (N_6378,N_306,N_4044);
and U6379 (N_6379,N_2814,N_4511);
or U6380 (N_6380,N_270,N_1153);
nand U6381 (N_6381,N_4014,N_2631);
nor U6382 (N_6382,N_2142,N_4696);
xor U6383 (N_6383,N_4162,N_3114);
nand U6384 (N_6384,N_2138,N_1267);
nand U6385 (N_6385,N_2855,N_691);
and U6386 (N_6386,N_2603,N_1722);
and U6387 (N_6387,N_595,N_4938);
or U6388 (N_6388,N_2939,N_260);
or U6389 (N_6389,N_3031,N_2261);
and U6390 (N_6390,N_3724,N_2484);
nand U6391 (N_6391,N_3825,N_2579);
and U6392 (N_6392,N_1313,N_1478);
xor U6393 (N_6393,N_1998,N_3235);
and U6394 (N_6394,N_1681,N_3621);
nand U6395 (N_6395,N_920,N_4996);
and U6396 (N_6396,N_2930,N_2109);
xnor U6397 (N_6397,N_4474,N_3092);
or U6398 (N_6398,N_4071,N_3682);
or U6399 (N_6399,N_2599,N_1738);
or U6400 (N_6400,N_4843,N_941);
or U6401 (N_6401,N_197,N_3111);
or U6402 (N_6402,N_2831,N_305);
nand U6403 (N_6403,N_739,N_1614);
nand U6404 (N_6404,N_4426,N_213);
nor U6405 (N_6405,N_549,N_508);
nor U6406 (N_6406,N_1572,N_2486);
or U6407 (N_6407,N_216,N_3376);
and U6408 (N_6408,N_1447,N_978);
nand U6409 (N_6409,N_3490,N_3214);
nor U6410 (N_6410,N_1359,N_2126);
xor U6411 (N_6411,N_3507,N_2543);
and U6412 (N_6412,N_4193,N_1291);
nand U6413 (N_6413,N_4043,N_3083);
xnor U6414 (N_6414,N_3927,N_1954);
xor U6415 (N_6415,N_3090,N_82);
or U6416 (N_6416,N_1914,N_2522);
xnor U6417 (N_6417,N_1456,N_4495);
nand U6418 (N_6418,N_1982,N_2237);
xnor U6419 (N_6419,N_2193,N_2570);
xor U6420 (N_6420,N_3781,N_1969);
or U6421 (N_6421,N_3961,N_786);
xnor U6422 (N_6422,N_2004,N_1034);
nor U6423 (N_6423,N_2535,N_3285);
xnor U6424 (N_6424,N_4324,N_2955);
and U6425 (N_6425,N_2780,N_2408);
or U6426 (N_6426,N_699,N_1691);
and U6427 (N_6427,N_89,N_4926);
nor U6428 (N_6428,N_1575,N_4829);
and U6429 (N_6429,N_726,N_2014);
nor U6430 (N_6430,N_4838,N_866);
nand U6431 (N_6431,N_3149,N_1538);
and U6432 (N_6432,N_874,N_3195);
xnor U6433 (N_6433,N_4520,N_4912);
nand U6434 (N_6434,N_2433,N_4981);
nand U6435 (N_6435,N_3146,N_4494);
nand U6436 (N_6436,N_680,N_2702);
xnor U6437 (N_6437,N_1905,N_2949);
nor U6438 (N_6438,N_616,N_397);
nor U6439 (N_6439,N_1202,N_3204);
nand U6440 (N_6440,N_2864,N_1560);
nor U6441 (N_6441,N_2698,N_1274);
xor U6442 (N_6442,N_1302,N_4585);
xor U6443 (N_6443,N_4155,N_4370);
and U6444 (N_6444,N_4603,N_788);
or U6445 (N_6445,N_2368,N_3441);
and U6446 (N_6446,N_372,N_1506);
or U6447 (N_6447,N_3044,N_392);
nand U6448 (N_6448,N_4842,N_1927);
nor U6449 (N_6449,N_318,N_3176);
nand U6450 (N_6450,N_2428,N_4446);
xnor U6451 (N_6451,N_1266,N_4484);
or U6452 (N_6452,N_3411,N_4430);
nor U6453 (N_6453,N_3755,N_2967);
and U6454 (N_6454,N_4128,N_1417);
nor U6455 (N_6455,N_3655,N_685);
nand U6456 (N_6456,N_4581,N_2325);
xor U6457 (N_6457,N_2690,N_3027);
xor U6458 (N_6458,N_3774,N_2712);
or U6459 (N_6459,N_4734,N_4284);
or U6460 (N_6460,N_4189,N_1190);
or U6461 (N_6461,N_1723,N_4339);
nor U6462 (N_6462,N_2478,N_2440);
nor U6463 (N_6463,N_2323,N_1184);
and U6464 (N_6464,N_1438,N_2649);
or U6465 (N_6465,N_4468,N_4404);
nor U6466 (N_6466,N_3754,N_927);
nor U6467 (N_6467,N_4371,N_331);
or U6468 (N_6468,N_3531,N_4636);
nand U6469 (N_6469,N_4802,N_2148);
nor U6470 (N_6470,N_581,N_3722);
and U6471 (N_6471,N_528,N_3988);
and U6472 (N_6472,N_4576,N_2845);
nor U6473 (N_6473,N_679,N_321);
xor U6474 (N_6474,N_1044,N_1222);
nor U6475 (N_6475,N_453,N_976);
xnor U6476 (N_6476,N_2926,N_934);
and U6477 (N_6477,N_3970,N_1618);
nand U6478 (N_6478,N_1121,N_2097);
nor U6479 (N_6479,N_3243,N_2364);
nor U6480 (N_6480,N_825,N_1907);
or U6481 (N_6481,N_4335,N_2835);
nor U6482 (N_6482,N_3393,N_3693);
nor U6483 (N_6483,N_4191,N_3434);
nor U6484 (N_6484,N_4749,N_3293);
nand U6485 (N_6485,N_728,N_4473);
xnor U6486 (N_6486,N_2734,N_2648);
nor U6487 (N_6487,N_3279,N_4725);
nor U6488 (N_6488,N_4572,N_277);
xnor U6489 (N_6489,N_798,N_1346);
nand U6490 (N_6490,N_2217,N_1032);
nand U6491 (N_6491,N_3914,N_3023);
or U6492 (N_6492,N_1578,N_1139);
nor U6493 (N_6493,N_490,N_43);
or U6494 (N_6494,N_552,N_2158);
or U6495 (N_6495,N_3915,N_1933);
nand U6496 (N_6496,N_4081,N_2322);
nand U6497 (N_6497,N_2256,N_166);
or U6498 (N_6498,N_618,N_3368);
and U6499 (N_6499,N_3686,N_3544);
nand U6500 (N_6500,N_4644,N_982);
or U6501 (N_6501,N_1031,N_2978);
or U6502 (N_6502,N_1502,N_782);
and U6503 (N_6503,N_2286,N_4878);
and U6504 (N_6504,N_3679,N_829);
or U6505 (N_6505,N_2695,N_2309);
and U6506 (N_6506,N_921,N_638);
and U6507 (N_6507,N_3097,N_2082);
xnor U6508 (N_6508,N_4196,N_1757);
or U6509 (N_6509,N_3383,N_3323);
nor U6510 (N_6510,N_4173,N_3367);
xnor U6511 (N_6511,N_1524,N_3579);
nor U6512 (N_6512,N_4283,N_1295);
or U6513 (N_6513,N_570,N_4109);
or U6514 (N_6514,N_3687,N_2646);
or U6515 (N_6515,N_344,N_2446);
nor U6516 (N_6516,N_2461,N_1058);
nand U6517 (N_6517,N_2513,N_1123);
nand U6518 (N_6518,N_2450,N_1376);
xor U6519 (N_6519,N_4584,N_2861);
and U6520 (N_6520,N_1785,N_3004);
and U6521 (N_6521,N_767,N_3681);
nand U6522 (N_6522,N_3768,N_148);
or U6523 (N_6523,N_898,N_3398);
xor U6524 (N_6524,N_2053,N_4656);
nand U6525 (N_6525,N_479,N_3473);
nor U6526 (N_6526,N_856,N_1135);
or U6527 (N_6527,N_2903,N_4451);
nor U6528 (N_6528,N_4030,N_749);
nand U6529 (N_6529,N_3134,N_944);
or U6530 (N_6530,N_2012,N_1305);
xor U6531 (N_6531,N_1828,N_206);
xor U6532 (N_6532,N_3167,N_529);
nor U6533 (N_6533,N_2778,N_1729);
xor U6534 (N_6534,N_4991,N_4112);
and U6535 (N_6535,N_755,N_4606);
and U6536 (N_6536,N_226,N_883);
or U6537 (N_6537,N_3194,N_375);
nor U6538 (N_6538,N_3213,N_4769);
xor U6539 (N_6539,N_4856,N_2786);
nor U6540 (N_6540,N_2451,N_723);
nand U6541 (N_6541,N_3550,N_4441);
or U6542 (N_6542,N_3562,N_1373);
nor U6543 (N_6543,N_4782,N_4291);
nand U6544 (N_6544,N_708,N_4823);
or U6545 (N_6545,N_518,N_1010);
or U6546 (N_6546,N_2618,N_3254);
xor U6547 (N_6547,N_4497,N_1803);
or U6548 (N_6548,N_4037,N_1528);
nand U6549 (N_6549,N_1069,N_4862);
or U6550 (N_6550,N_3262,N_4243);
or U6551 (N_6551,N_3460,N_713);
and U6552 (N_6552,N_1940,N_4103);
nand U6553 (N_6553,N_730,N_1946);
or U6554 (N_6554,N_3983,N_3369);
nand U6555 (N_6555,N_3695,N_3992);
nand U6556 (N_6556,N_4074,N_3478);
nand U6557 (N_6557,N_110,N_2202);
or U6558 (N_6558,N_9,N_1682);
or U6559 (N_6559,N_559,N_429);
xor U6560 (N_6560,N_2152,N_3420);
or U6561 (N_6561,N_1769,N_140);
or U6562 (N_6562,N_3899,N_4717);
or U6563 (N_6563,N_3619,N_3664);
nor U6564 (N_6564,N_607,N_754);
nand U6565 (N_6565,N_2418,N_4571);
and U6566 (N_6566,N_4730,N_4131);
or U6567 (N_6567,N_984,N_668);
xnor U6568 (N_6568,N_100,N_363);
and U6569 (N_6569,N_4890,N_842);
and U6570 (N_6570,N_3750,N_2576);
xnor U6571 (N_6571,N_4788,N_2954);
or U6572 (N_6572,N_4986,N_4466);
xnor U6573 (N_6573,N_582,N_745);
nand U6574 (N_6574,N_4984,N_2386);
and U6575 (N_6575,N_3748,N_2675);
xor U6576 (N_6576,N_4062,N_2114);
nor U6577 (N_6577,N_4633,N_3731);
and U6578 (N_6578,N_2787,N_1246);
or U6579 (N_6579,N_936,N_2580);
and U6580 (N_6580,N_3121,N_2199);
nand U6581 (N_6581,N_4774,N_1664);
and U6582 (N_6582,N_3051,N_2624);
nor U6583 (N_6583,N_3257,N_302);
or U6584 (N_6584,N_3981,N_2934);
or U6585 (N_6585,N_4824,N_3971);
xor U6586 (N_6586,N_697,N_59);
or U6587 (N_6587,N_517,N_4460);
and U6588 (N_6588,N_3661,N_4612);
nor U6589 (N_6589,N_4235,N_4952);
nor U6590 (N_6590,N_1607,N_1813);
and U6591 (N_6591,N_427,N_1822);
or U6592 (N_6592,N_2870,N_3021);
nor U6593 (N_6593,N_4844,N_3404);
and U6594 (N_6594,N_416,N_3150);
xnor U6595 (N_6595,N_2155,N_2472);
or U6596 (N_6596,N_4687,N_4976);
and U6597 (N_6597,N_790,N_4352);
nor U6598 (N_6598,N_3482,N_4694);
nor U6599 (N_6599,N_2214,N_2068);
nand U6600 (N_6600,N_880,N_696);
or U6601 (N_6601,N_4412,N_2860);
nand U6602 (N_6602,N_565,N_145);
nand U6603 (N_6603,N_1951,N_3968);
nand U6604 (N_6604,N_1628,N_1018);
nand U6605 (N_6605,N_4615,N_1976);
xnor U6606 (N_6606,N_4815,N_931);
or U6607 (N_6607,N_272,N_4779);
xor U6608 (N_6608,N_4695,N_1978);
or U6609 (N_6609,N_3616,N_383);
nand U6610 (N_6610,N_2232,N_746);
nand U6611 (N_6611,N_792,N_4863);
xnor U6612 (N_6612,N_2936,N_12);
and U6613 (N_6613,N_2274,N_3442);
xnor U6614 (N_6614,N_1861,N_1851);
or U6615 (N_6615,N_2730,N_2824);
and U6616 (N_6616,N_2196,N_2961);
nor U6617 (N_6617,N_1832,N_3469);
nand U6618 (N_6618,N_2230,N_1020);
nor U6619 (N_6619,N_2849,N_2567);
and U6620 (N_6620,N_1212,N_69);
nor U6621 (N_6621,N_1255,N_186);
or U6622 (N_6622,N_2231,N_240);
nor U6623 (N_6623,N_4114,N_2816);
and U6624 (N_6624,N_1290,N_830);
nor U6625 (N_6625,N_2583,N_2454);
or U6626 (N_6626,N_1753,N_1627);
nor U6627 (N_6627,N_4297,N_4536);
nor U6628 (N_6628,N_3265,N_3921);
nor U6629 (N_6629,N_3125,N_536);
and U6630 (N_6630,N_2498,N_2728);
or U6631 (N_6631,N_793,N_1793);
and U6632 (N_6632,N_1550,N_4627);
nand U6633 (N_6633,N_1361,N_1043);
nor U6634 (N_6634,N_4251,N_3924);
or U6635 (N_6635,N_1695,N_3357);
nor U6636 (N_6636,N_3263,N_4180);
xor U6637 (N_6637,N_2529,N_346);
and U6638 (N_6638,N_3946,N_1470);
xnor U6639 (N_6639,N_3828,N_4522);
and U6640 (N_6640,N_1299,N_777);
nand U6641 (N_6641,N_301,N_3698);
or U6642 (N_6642,N_527,N_291);
xor U6643 (N_6643,N_2101,N_1924);
nor U6644 (N_6644,N_1893,N_4396);
or U6645 (N_6645,N_92,N_4070);
and U6646 (N_6646,N_4884,N_4697);
nand U6647 (N_6647,N_2019,N_3953);
and U6648 (N_6648,N_390,N_4710);
nand U6649 (N_6649,N_2813,N_2694);
or U6650 (N_6650,N_1288,N_2521);
or U6651 (N_6651,N_3547,N_2306);
and U6652 (N_6652,N_4258,N_2645);
nand U6653 (N_6653,N_4436,N_2553);
xnor U6654 (N_6654,N_2636,N_3096);
nor U6655 (N_6655,N_228,N_714);
and U6656 (N_6656,N_3475,N_1518);
and U6657 (N_6657,N_4920,N_1548);
nor U6658 (N_6658,N_3801,N_138);
and U6659 (N_6659,N_3154,N_90);
nand U6660 (N_6660,N_1877,N_3419);
and U6661 (N_6661,N_3115,N_396);
xor U6662 (N_6662,N_4544,N_1334);
and U6663 (N_6663,N_4807,N_1716);
nand U6664 (N_6664,N_1490,N_3326);
xnor U6665 (N_6665,N_4706,N_2340);
xor U6666 (N_6666,N_3206,N_4738);
nand U6667 (N_6667,N_4558,N_1028);
and U6668 (N_6668,N_606,N_4727);
xnor U6669 (N_6669,N_3891,N_4028);
and U6670 (N_6670,N_929,N_1983);
xor U6671 (N_6671,N_2632,N_8);
nor U6672 (N_6672,N_2842,N_1778);
nor U6673 (N_6673,N_619,N_4334);
nand U6674 (N_6674,N_1706,N_4186);
nor U6675 (N_6675,N_3219,N_3552);
or U6676 (N_6676,N_3645,N_655);
or U6677 (N_6677,N_3308,N_3087);
nand U6678 (N_6678,N_488,N_1317);
nand U6679 (N_6679,N_2779,N_2705);
nand U6680 (N_6680,N_4628,N_1453);
nor U6681 (N_6681,N_4554,N_4662);
xnor U6682 (N_6682,N_2495,N_3700);
nor U6683 (N_6683,N_2988,N_2707);
nand U6684 (N_6684,N_2577,N_3465);
nor U6685 (N_6685,N_608,N_476);
and U6686 (N_6686,N_802,N_1372);
or U6687 (N_6687,N_3450,N_2348);
or U6688 (N_6688,N_2011,N_4755);
xnor U6689 (N_6689,N_2822,N_2533);
and U6690 (N_6690,N_2447,N_91);
xnor U6691 (N_6691,N_3587,N_625);
nor U6692 (N_6692,N_2000,N_393);
and U6693 (N_6693,N_212,N_4113);
xnor U6694 (N_6694,N_448,N_3072);
xor U6695 (N_6695,N_3800,N_4759);
xor U6696 (N_6696,N_4723,N_1733);
and U6697 (N_6697,N_1563,N_2704);
nor U6698 (N_6698,N_3073,N_4692);
nand U6699 (N_6699,N_4210,N_2944);
nand U6700 (N_6700,N_4338,N_2917);
and U6701 (N_6701,N_2334,N_3006);
nor U6702 (N_6702,N_4791,N_3251);
nand U6703 (N_6703,N_3519,N_4336);
xnor U6704 (N_6704,N_1826,N_4198);
nor U6705 (N_6705,N_2612,N_4871);
nor U6706 (N_6706,N_2067,N_753);
xor U6707 (N_6707,N_2777,N_3922);
and U6708 (N_6708,N_832,N_3333);
and U6709 (N_6709,N_221,N_4501);
or U6710 (N_6710,N_4901,N_469);
nor U6711 (N_6711,N_3354,N_2989);
nor U6712 (N_6712,N_4886,N_2620);
and U6713 (N_6713,N_4718,N_3853);
nor U6714 (N_6714,N_3020,N_1183);
nor U6715 (N_6715,N_1067,N_439);
nand U6716 (N_6716,N_2726,N_380);
nand U6717 (N_6717,N_3036,N_14);
xor U6718 (N_6718,N_3633,N_3690);
nor U6719 (N_6719,N_4309,N_2001);
nor U6720 (N_6720,N_2750,N_2997);
nand U6721 (N_6721,N_1509,N_3591);
xor U6722 (N_6722,N_2922,N_1443);
xor U6723 (N_6723,N_2353,N_1015);
or U6724 (N_6724,N_3956,N_1134);
nor U6725 (N_6725,N_3871,N_4399);
nand U6726 (N_6726,N_4828,N_3784);
xnor U6727 (N_6727,N_4547,N_865);
or U6728 (N_6728,N_391,N_3772);
xnor U6729 (N_6729,N_460,N_307);
or U6730 (N_6730,N_916,N_3522);
nand U6731 (N_6731,N_3646,N_3578);
xnor U6732 (N_6732,N_1179,N_4122);
xnor U6733 (N_6733,N_2038,N_1238);
or U6734 (N_6734,N_2572,N_1846);
xnor U6735 (N_6735,N_4566,N_3440);
or U6736 (N_6736,N_4486,N_2469);
nand U6737 (N_6737,N_1449,N_2271);
nor U6738 (N_6738,N_4089,N_502);
nor U6739 (N_6739,N_1567,N_303);
nor U6740 (N_6740,N_1704,N_1967);
or U6741 (N_6741,N_3812,N_2022);
or U6742 (N_6742,N_2724,N_3282);
xor U6743 (N_6743,N_4562,N_2234);
or U6744 (N_6744,N_2847,N_1457);
nand U6745 (N_6745,N_1642,N_3841);
and U6746 (N_6746,N_3311,N_2235);
and U6747 (N_6747,N_3226,N_2994);
or U6748 (N_6748,N_4622,N_933);
nand U6749 (N_6749,N_32,N_4392);
nor U6750 (N_6750,N_2431,N_142);
nand U6751 (N_6751,N_4745,N_1336);
xnor U6752 (N_6752,N_4510,N_1579);
nor U6753 (N_6753,N_3537,N_2241);
or U6754 (N_6754,N_2977,N_1142);
nand U6755 (N_6755,N_4250,N_1395);
nand U6756 (N_6756,N_2880,N_1085);
nand U6757 (N_6757,N_4967,N_637);
xnor U6758 (N_6758,N_1721,N_1812);
and U6759 (N_6759,N_2402,N_2637);
xnor U6760 (N_6760,N_4464,N_1362);
nor U6761 (N_6761,N_3855,N_1110);
xor U6762 (N_6762,N_3660,N_3520);
xnor U6763 (N_6763,N_4192,N_3691);
xor U6764 (N_6764,N_4632,N_3169);
nor U6765 (N_6765,N_3862,N_2411);
nand U6766 (N_6766,N_1505,N_546);
xnor U6767 (N_6767,N_3205,N_3132);
or U6768 (N_6768,N_2088,N_208);
nor U6769 (N_6769,N_2132,N_3337);
and U6770 (N_6770,N_2171,N_3564);
nand U6771 (N_6771,N_1806,N_4054);
nand U6772 (N_6772,N_3882,N_1588);
nor U6773 (N_6773,N_1468,N_3290);
nor U6774 (N_6774,N_106,N_1001);
nand U6775 (N_6775,N_2556,N_1177);
nor U6776 (N_6776,N_310,N_2879);
nand U6777 (N_6777,N_1025,N_1223);
or U6778 (N_6778,N_1871,N_495);
or U6779 (N_6779,N_507,N_2160);
or U6780 (N_6780,N_1593,N_3555);
or U6781 (N_6781,N_3300,N_716);
and U6782 (N_6782,N_1256,N_4858);
xnor U6783 (N_6783,N_3969,N_3870);
or U6784 (N_6784,N_2990,N_3821);
nor U6785 (N_6785,N_3446,N_3135);
nand U6786 (N_6786,N_3810,N_1389);
or U6787 (N_6787,N_4298,N_1492);
xnor U6788 (N_6788,N_4932,N_1974);
xnor U6789 (N_6789,N_2593,N_87);
and U6790 (N_6790,N_2956,N_3116);
or U6791 (N_6791,N_2823,N_4385);
nand U6792 (N_6792,N_4961,N_34);
nand U6793 (N_6793,N_1873,N_2314);
xor U6794 (N_6794,N_3590,N_1428);
and U6795 (N_6795,N_4401,N_1261);
nand U6796 (N_6796,N_2365,N_1176);
and U6797 (N_6797,N_3554,N_4025);
nor U6798 (N_6798,N_39,N_3258);
nand U6799 (N_6799,N_695,N_1174);
and U6800 (N_6800,N_1797,N_2187);
nor U6801 (N_6801,N_2169,N_3804);
nor U6802 (N_6802,N_1150,N_1734);
nand U6803 (N_6803,N_3920,N_1415);
nand U6804 (N_6804,N_1917,N_1378);
xor U6805 (N_6805,N_4179,N_4491);
xnor U6806 (N_6806,N_1324,N_1939);
nand U6807 (N_6807,N_4869,N_4801);
and U6808 (N_6808,N_1101,N_4224);
or U6809 (N_6809,N_1377,N_826);
nand U6810 (N_6810,N_828,N_225);
and U6811 (N_6811,N_922,N_456);
xnor U6812 (N_6812,N_3395,N_4653);
nor U6813 (N_6813,N_3370,N_349);
xnor U6814 (N_6814,N_1472,N_154);
or U6815 (N_6815,N_1272,N_2773);
or U6816 (N_6816,N_382,N_2267);
nand U6817 (N_6817,N_1257,N_3174);
nor U6818 (N_6818,N_2963,N_1162);
nand U6819 (N_6819,N_4228,N_1206);
and U6820 (N_6820,N_4775,N_1512);
and U6821 (N_6821,N_1559,N_868);
nand U6822 (N_6822,N_4289,N_948);
nor U6823 (N_6823,N_4098,N_2480);
xnor U6824 (N_6824,N_3013,N_4787);
xnor U6825 (N_6825,N_2827,N_2534);
xnor U6826 (N_6826,N_1780,N_3139);
xnor U6827 (N_6827,N_3553,N_4773);
and U6828 (N_6828,N_649,N_1087);
xnor U6829 (N_6829,N_296,N_771);
nand U6830 (N_6830,N_4011,N_2542);
nor U6831 (N_6831,N_4848,N_4211);
or U6832 (N_6832,N_4499,N_1529);
or U6833 (N_6833,N_2546,N_178);
nand U6834 (N_6834,N_2054,N_268);
or U6835 (N_6835,N_2047,N_4750);
xor U6836 (N_6836,N_687,N_415);
or U6837 (N_6837,N_761,N_1211);
or U6838 (N_6838,N_661,N_1192);
nand U6839 (N_6839,N_1830,N_4982);
or U6840 (N_6840,N_1003,N_1696);
and U6841 (N_6841,N_4685,N_3145);
nand U6842 (N_6842,N_4641,N_1650);
nand U6843 (N_6843,N_2761,N_3965);
nor U6844 (N_6844,N_1036,N_879);
xor U6845 (N_6845,N_3506,N_3928);
xor U6846 (N_6846,N_3551,N_10);
nor U6847 (N_6847,N_2311,N_3297);
nand U6848 (N_6848,N_975,N_1237);
or U6849 (N_6849,N_104,N_1908);
nor U6850 (N_6850,N_542,N_2091);
nand U6851 (N_6851,N_1977,N_1671);
or U6852 (N_6852,N_2093,N_2638);
nor U6853 (N_6853,N_4244,N_3397);
or U6854 (N_6854,N_1711,N_2128);
nand U6855 (N_6855,N_1878,N_3770);
nor U6856 (N_6856,N_1849,N_4502);
and U6857 (N_6857,N_839,N_4072);
or U6858 (N_6858,N_2805,N_4463);
and U6859 (N_6859,N_2376,N_1263);
xnor U6860 (N_6860,N_851,N_4975);
and U6861 (N_6861,N_2221,N_4778);
or U6862 (N_6862,N_2762,N_1896);
nand U6863 (N_6863,N_4166,N_3339);
xnor U6864 (N_6864,N_4953,N_3607);
and U6865 (N_6865,N_1657,N_632);
xnor U6866 (N_6866,N_2468,N_2765);
and U6867 (N_6867,N_370,N_1942);
xnor U6868 (N_6868,N_3543,N_2227);
or U6869 (N_6869,N_4910,N_4104);
xor U6870 (N_6870,N_4663,N_3838);
nor U6871 (N_6871,N_2892,N_4342);
nand U6872 (N_6872,N_315,N_1707);
or U6873 (N_6873,N_4231,N_1788);
nand U6874 (N_6874,N_890,N_4031);
or U6875 (N_6875,N_2974,N_4816);
and U6876 (N_6876,N_4079,N_1862);
or U6877 (N_6877,N_3982,N_3896);
or U6878 (N_6878,N_1040,N_461);
nor U6879 (N_6879,N_3835,N_3386);
or U6880 (N_6880,N_41,N_1937);
nor U6881 (N_6881,N_914,N_774);
xor U6882 (N_6882,N_4704,N_4492);
nor U6883 (N_6883,N_4229,N_3668);
nor U6884 (N_6884,N_2372,N_1602);
nand U6885 (N_6885,N_109,N_4777);
nor U6886 (N_6886,N_5,N_2700);
nand U6887 (N_6887,N_134,N_1335);
xnor U6888 (N_6888,N_1890,N_4639);
nand U6889 (N_6889,N_3819,N_3497);
nor U6890 (N_6890,N_1709,N_3242);
and U6891 (N_6891,N_3289,N_2459);
and U6892 (N_6892,N_1576,N_1537);
and U6893 (N_6893,N_2025,N_475);
or U6894 (N_6894,N_1350,N_4587);
or U6895 (N_6895,N_4740,N_4541);
and U6896 (N_6896,N_3079,N_4880);
or U6897 (N_6897,N_27,N_1422);
or U6898 (N_6898,N_273,N_2220);
and U6899 (N_6899,N_4665,N_2010);
nand U6900 (N_6900,N_2039,N_4163);
or U6901 (N_6901,N_686,N_4383);
nor U6902 (N_6902,N_2709,N_505);
or U6903 (N_6903,N_155,N_1495);
nand U6904 (N_6904,N_3074,N_2488);
or U6905 (N_6905,N_2666,N_4130);
and U6906 (N_6906,N_3950,N_2065);
nand U6907 (N_6907,N_3067,N_951);
and U6908 (N_6908,N_4951,N_2532);
or U6909 (N_6909,N_554,N_4504);
nand U6910 (N_6910,N_3959,N_4145);
and U6911 (N_6911,N_4664,N_4693);
or U6912 (N_6912,N_1530,N_4578);
or U6913 (N_6913,N_4498,N_3666);
nor U6914 (N_6914,N_3462,N_347);
nor U6915 (N_6915,N_3063,N_2536);
nor U6916 (N_6916,N_656,N_2218);
and U6917 (N_6917,N_1945,N_3009);
and U6918 (N_6918,N_4512,N_1433);
or U6919 (N_6919,N_3944,N_4003);
or U6920 (N_6920,N_4916,N_1649);
or U6921 (N_6921,N_3315,N_2471);
or U6922 (N_6922,N_1229,N_3510);
and U6923 (N_6923,N_4,N_2358);
xnor U6924 (N_6924,N_3884,N_1957);
nor U6925 (N_6925,N_1307,N_1285);
and U6926 (N_6926,N_4386,N_4475);
or U6927 (N_6927,N_764,N_3575);
xnor U6928 (N_6928,N_3313,N_1859);
nor U6929 (N_6929,N_1759,N_801);
or U6930 (N_6930,N_853,N_4783);
nand U6931 (N_6931,N_4405,N_2924);
nand U6932 (N_6932,N_3651,N_478);
nand U6933 (N_6933,N_1298,N_1727);
xor U6934 (N_6934,N_629,N_3881);
or U6935 (N_6935,N_2122,N_4158);
nand U6936 (N_6936,N_1673,N_2758);
or U6937 (N_6937,N_3948,N_1949);
nor U6938 (N_6938,N_2434,N_862);
xnor U6939 (N_6939,N_2975,N_2124);
or U6940 (N_6940,N_3570,N_3222);
xnor U6941 (N_6941,N_563,N_520);
and U6942 (N_6942,N_276,N_4770);
nand U6943 (N_6943,N_4538,N_2817);
or U6944 (N_6944,N_3759,N_799);
and U6945 (N_6945,N_114,N_2157);
xnor U6946 (N_6946,N_2477,N_2764);
and U6947 (N_6947,N_298,N_3704);
nand U6948 (N_6948,N_1881,N_748);
nand U6949 (N_6949,N_1487,N_2594);
nor U6950 (N_6950,N_432,N_4551);
or U6951 (N_6951,N_2689,N_861);
xnor U6952 (N_6952,N_4557,N_2937);
or U6953 (N_6953,N_3124,N_758);
nor U6954 (N_6954,N_3483,N_3084);
or U6955 (N_6955,N_95,N_202);
nor U6956 (N_6956,N_463,N_3962);
and U6957 (N_6957,N_3739,N_468);
nor U6958 (N_6958,N_2815,N_1130);
and U6959 (N_6959,N_1776,N_2796);
nor U6960 (N_6960,N_3363,N_3075);
nand U6961 (N_6961,N_3152,N_848);
nand U6962 (N_6962,N_1196,N_3062);
or U6963 (N_6963,N_45,N_2940);
and U6964 (N_6964,N_884,N_1234);
or U6965 (N_6965,N_428,N_63);
nor U6966 (N_6966,N_2326,N_3538);
and U6967 (N_6967,N_2197,N_2769);
nand U6968 (N_6968,N_3185,N_1833);
or U6969 (N_6969,N_1710,N_4260);
xnor U6970 (N_6970,N_2804,N_2616);
or U6971 (N_6971,N_4408,N_3346);
nand U6972 (N_6972,N_1037,N_3425);
nor U6973 (N_6973,N_1351,N_4319);
and U6974 (N_6974,N_3171,N_641);
or U6975 (N_6975,N_2276,N_168);
or U6976 (N_6976,N_3954,N_958);
and U6977 (N_6977,N_2714,N_1700);
and U6978 (N_6978,N_2838,N_4683);
and U6979 (N_6979,N_2854,N_2776);
nor U6980 (N_6980,N_222,N_4797);
xnor U6981 (N_6981,N_4419,N_4957);
and U6982 (N_6982,N_4010,N_147);
or U6983 (N_6983,N_1536,N_4411);
nand U6984 (N_6984,N_2185,N_3264);
xnor U6985 (N_6985,N_3951,N_3676);
xor U6986 (N_6986,N_3728,N_2396);
nand U6987 (N_6987,N_3514,N_3967);
nand U6988 (N_6988,N_4488,N_2581);
or U6989 (N_6989,N_2530,N_3582);
nand U6990 (N_6990,N_2628,N_4814);
nand U6991 (N_6991,N_2548,N_1332);
or U6992 (N_6992,N_3941,N_910);
nor U6993 (N_6993,N_2479,N_3458);
nor U6994 (N_6994,N_395,N_324);
nor U6995 (N_6995,N_500,N_3180);
xor U6996 (N_6996,N_791,N_3688);
nor U6997 (N_6997,N_1322,N_2321);
nand U6998 (N_6998,N_1277,N_174);
or U6999 (N_6999,N_334,N_1168);
and U7000 (N_7000,N_1781,N_3938);
or U7001 (N_7001,N_2501,N_2021);
and U7002 (N_7002,N_4106,N_1065);
xnor U7003 (N_7003,N_4068,N_3271);
or U7004 (N_7004,N_317,N_2837);
nand U7005 (N_7005,N_150,N_1189);
nand U7006 (N_7006,N_4388,N_1625);
nor U7007 (N_7007,N_531,N_256);
nor U7008 (N_7008,N_4138,N_487);
nor U7009 (N_7009,N_1674,N_419);
nand U7010 (N_7010,N_2946,N_1648);
xnor U7011 (N_7011,N_1622,N_4034);
nand U7012 (N_7012,N_2771,N_1545);
xnor U7013 (N_7013,N_2383,N_4513);
or U7014 (N_7014,N_2840,N_980);
nor U7015 (N_7015,N_2441,N_330);
xor U7016 (N_7016,N_435,N_3634);
nand U7017 (N_7017,N_1739,N_257);
and U7018 (N_7018,N_4737,N_945);
or U7019 (N_7019,N_631,N_4111);
nand U7020 (N_7020,N_455,N_2766);
nor U7021 (N_7021,N_1382,N_1499);
and U7022 (N_7022,N_2589,N_4766);
and U7023 (N_7023,N_2467,N_3996);
xnor U7024 (N_7024,N_3399,N_2198);
nor U7025 (N_7025,N_3737,N_597);
nor U7026 (N_7026,N_803,N_1170);
xnor U7027 (N_7027,N_624,N_676);
xnor U7028 (N_7028,N_3402,N_2732);
and U7029 (N_7029,N_4928,N_4359);
xnor U7030 (N_7030,N_3650,N_3029);
xor U7031 (N_7031,N_2328,N_4919);
nor U7032 (N_7032,N_3182,N_2302);
and U7033 (N_7033,N_2032,N_4688);
or U7034 (N_7034,N_1338,N_4948);
and U7035 (N_7035,N_1959,N_2610);
nand U7036 (N_7036,N_2485,N_3144);
and U7037 (N_7037,N_840,N_1242);
and U7038 (N_7038,N_1233,N_858);
and U7039 (N_7039,N_4444,N_620);
and U7040 (N_7040,N_2558,N_1125);
and U7041 (N_7041,N_4839,N_362);
xnor U7042 (N_7042,N_3330,N_4800);
xor U7043 (N_7043,N_2379,N_671);
xor U7044 (N_7044,N_1083,N_3714);
xor U7045 (N_7045,N_634,N_364);
xnor U7046 (N_7046,N_4832,N_4799);
nor U7047 (N_7047,N_3601,N_3677);
xnor U7048 (N_7048,N_2808,N_271);
nor U7049 (N_7049,N_4613,N_4237);
or U7050 (N_7050,N_797,N_4316);
or U7051 (N_7051,N_2042,N_2410);
nand U7052 (N_7052,N_4935,N_2293);
xnor U7053 (N_7053,N_1420,N_2374);
nand U7054 (N_7054,N_2525,N_3104);
nand U7055 (N_7055,N_2538,N_3457);
nor U7056 (N_7056,N_1306,N_1301);
or U7057 (N_7057,N_4389,N_831);
xnor U7058 (N_7058,N_928,N_2803);
nor U7059 (N_7059,N_3892,N_844);
and U7060 (N_7060,N_4331,N_243);
nor U7061 (N_7061,N_4619,N_1030);
and U7062 (N_7062,N_1587,N_670);
and U7063 (N_7063,N_4218,N_998);
nor U7064 (N_7064,N_4857,N_734);
or U7065 (N_7065,N_643,N_4362);
nand U7066 (N_7066,N_3525,N_2228);
nor U7067 (N_7067,N_2113,N_1848);
nand U7068 (N_7068,N_2357,N_2609);
nor U7069 (N_7069,N_3936,N_503);
or U7070 (N_7070,N_2389,N_3792);
nand U7071 (N_7071,N_311,N_698);
xor U7072 (N_7072,N_4671,N_3269);
nor U7073 (N_7073,N_4573,N_4643);
xor U7074 (N_7074,N_2673,N_1985);
or U7075 (N_7075,N_4655,N_3108);
and U7076 (N_7076,N_2812,N_4515);
or U7077 (N_7077,N_3504,N_4577);
nand U7078 (N_7078,N_355,N_2790);
and U7079 (N_7079,N_3712,N_869);
nand U7080 (N_7080,N_2643,N_3839);
xor U7081 (N_7081,N_442,N_3745);
or U7082 (N_7082,N_4281,N_4400);
and U7083 (N_7083,N_544,N_1207);
and U7084 (N_7084,N_4818,N_4168);
or U7085 (N_7085,N_2423,N_3964);
or U7086 (N_7086,N_2473,N_4105);
or U7087 (N_7087,N_2182,N_2291);
or U7088 (N_7088,N_3307,N_3296);
or U7089 (N_7089,N_4579,N_4487);
nand U7090 (N_7090,N_2086,N_4450);
and U7091 (N_7091,N_3610,N_2077);
xnor U7092 (N_7092,N_112,N_3015);
nand U7093 (N_7093,N_519,N_1677);
xor U7094 (N_7094,N_4015,N_3910);
and U7095 (N_7095,N_4206,N_992);
xnor U7096 (N_7096,N_4403,N_3809);
nand U7097 (N_7097,N_4099,N_180);
and U7098 (N_7098,N_954,N_1510);
or U7099 (N_7099,N_120,N_351);
xnor U7100 (N_7100,N_3252,N_3066);
or U7101 (N_7101,N_1432,N_2607);
and U7102 (N_7102,N_4363,N_756);
or U7103 (N_7103,N_4931,N_322);
xnor U7104 (N_7104,N_3545,N_1340);
and U7105 (N_7105,N_3412,N_2502);
nand U7106 (N_7106,N_3843,N_3869);
or U7107 (N_7107,N_1108,N_2260);
nor U7108 (N_7108,N_4589,N_2388);
and U7109 (N_7109,N_3384,N_3851);
nand U7110 (N_7110,N_4605,N_532);
nand U7111 (N_7111,N_3201,N_187);
nor U7112 (N_7112,N_281,N_3886);
xor U7113 (N_7113,N_4039,N_1883);
or U7114 (N_7114,N_2170,N_3147);
and U7115 (N_7115,N_1748,N_4942);
and U7116 (N_7116,N_465,N_3248);
nor U7117 (N_7117,N_763,N_4729);
xor U7118 (N_7118,N_4833,N_2266);
nand U7119 (N_7119,N_3161,N_1236);
nand U7120 (N_7120,N_3929,N_1792);
nand U7121 (N_7121,N_4207,N_3103);
nand U7122 (N_7122,N_4378,N_3897);
xor U7123 (N_7123,N_4318,N_96);
xnor U7124 (N_7124,N_287,N_2432);
and U7125 (N_7125,N_770,N_1215);
and U7126 (N_7126,N_2188,N_3422);
or U7127 (N_7127,N_940,N_4182);
or U7128 (N_7128,N_885,N_760);
nor U7129 (N_7129,N_314,N_996);
nor U7130 (N_7130,N_3815,N_1282);
or U7131 (N_7131,N_4365,N_1922);
nand U7132 (N_7132,N_2916,N_4764);
or U7133 (N_7133,N_4313,N_578);
and U7134 (N_7134,N_4728,N_3122);
xnor U7135 (N_7135,N_474,N_3979);
xor U7136 (N_7136,N_369,N_1129);
or U7137 (N_7137,N_2881,N_1638);
or U7138 (N_7138,N_1154,N_864);
xnor U7139 (N_7139,N_838,N_3409);
or U7140 (N_7140,N_2223,N_2262);
nand U7141 (N_7141,N_2494,N_3785);
or U7142 (N_7142,N_4458,N_2213);
or U7143 (N_7143,N_2351,N_1149);
nand U7144 (N_7144,N_4670,N_837);
nor U7145 (N_7145,N_4238,N_83);
and U7146 (N_7146,N_1888,N_2520);
or U7147 (N_7147,N_4954,N_232);
xor U7148 (N_7148,N_3236,N_2264);
xnor U7149 (N_7149,N_329,N_2807);
nand U7150 (N_7150,N_663,N_995);
or U7151 (N_7151,N_3885,N_1024);
nand U7152 (N_7152,N_2832,N_1055);
nand U7153 (N_7153,N_3685,N_1583);
nor U7154 (N_7154,N_2107,N_4594);
or U7155 (N_7155,N_1437,N_2347);
or U7156 (N_7156,N_4548,N_3611);
and U7157 (N_7157,N_2181,N_2342);
and U7158 (N_7158,N_2405,N_1955);
nand U7159 (N_7159,N_2644,N_1366);
and U7160 (N_7160,N_917,N_3046);
nand U7161 (N_7161,N_1221,N_659);
nor U7162 (N_7162,N_3675,N_312);
nand U7163 (N_7163,N_1923,N_2098);
nor U7164 (N_7164,N_2481,N_52);
and U7165 (N_7165,N_71,N_2783);
nor U7166 (N_7166,N_4169,N_4811);
nand U7167 (N_7167,N_4174,N_2292);
nor U7168 (N_7168,N_4402,N_2439);
nor U7169 (N_7169,N_4826,N_3657);
or U7170 (N_7170,N_833,N_2154);
nor U7171 (N_7171,N_2466,N_4434);
xor U7172 (N_7172,N_76,N_1247);
nand U7173 (N_7173,N_795,N_280);
nor U7174 (N_7174,N_4367,N_1827);
and U7175 (N_7175,N_4350,N_1844);
nor U7176 (N_7176,N_398,N_156);
nand U7177 (N_7177,N_242,N_3436);
nand U7178 (N_7178,N_2006,N_964);
nand U7179 (N_7179,N_4806,N_1746);
or U7180 (N_7180,N_4864,N_4422);
nand U7181 (N_7181,N_4753,N_353);
nand U7182 (N_7182,N_3474,N_3826);
nor U7183 (N_7183,N_4407,N_450);
and U7184 (N_7184,N_3392,N_239);
xnor U7185 (N_7185,N_2566,N_2412);
nor U7186 (N_7186,N_2016,N_2002);
or U7187 (N_7187,N_1214,N_2465);
nand U7188 (N_7188,N_2737,N_2621);
and U7189 (N_7189,N_915,N_2317);
nor U7190 (N_7190,N_2204,N_2299);
xor U7191 (N_7191,N_2404,N_3614);
nor U7192 (N_7192,N_547,N_895);
xor U7193 (N_7193,N_1725,N_775);
xor U7194 (N_7194,N_3600,N_160);
nand U7195 (N_7195,N_152,N_4721);
or U7196 (N_7196,N_2444,N_313);
nand U7197 (N_7197,N_913,N_4624);
and U7198 (N_7198,N_4527,N_2782);
nand U7199 (N_7199,N_261,N_1749);
or U7200 (N_7200,N_3872,N_1652);
xnor U7201 (N_7201,N_328,N_2600);
nand U7202 (N_7202,N_2951,N_2629);
xor U7203 (N_7203,N_2360,N_3955);
nand U7204 (N_7204,N_1434,N_2686);
nor U7205 (N_7205,N_3832,N_2496);
xor U7206 (N_7206,N_300,N_1410);
nand U7207 (N_7207,N_26,N_1386);
or U7208 (N_7208,N_1095,N_3753);
nand U7209 (N_7209,N_209,N_497);
xnor U7210 (N_7210,N_4660,N_1767);
or U7211 (N_7211,N_3492,N_2743);
xor U7212 (N_7212,N_630,N_4955);
and U7213 (N_7213,N_3986,N_3476);
nand U7214 (N_7214,N_3999,N_4820);
nand U7215 (N_7215,N_2026,N_3596);
and U7216 (N_7216,N_1073,N_4875);
xnor U7217 (N_7217,N_394,N_4771);
xnor U7218 (N_7218,N_4804,N_541);
nor U7219 (N_7219,N_4095,N_1818);
nand U7220 (N_7220,N_1837,N_4675);
and U7221 (N_7221,N_2215,N_886);
or U7222 (N_7222,N_545,N_1163);
xor U7223 (N_7223,N_2191,N_20);
and U7224 (N_7224,N_511,N_4327);
and U7225 (N_7225,N_4027,N_3329);
or U7226 (N_7226,N_4358,N_472);
and U7227 (N_7227,N_2531,N_4420);
or U7228 (N_7228,N_2953,N_3275);
and U7229 (N_7229,N_1836,N_3467);
or U7230 (N_7230,N_3867,N_4637);
and U7231 (N_7231,N_4059,N_4564);
xnor U7232 (N_7232,N_1475,N_892);
xor U7233 (N_7233,N_3581,N_1554);
or U7234 (N_7234,N_4476,N_534);
or U7235 (N_7235,N_1686,N_3166);
or U7236 (N_7236,N_3689,N_3281);
nand U7237 (N_7237,N_2901,N_2031);
xor U7238 (N_7238,N_4233,N_2682);
and U7239 (N_7239,N_2490,N_3814);
nand U7240 (N_7240,N_3626,N_4521);
nand U7241 (N_7241,N_942,N_943);
and U7242 (N_7242,N_4891,N_1489);
xor U7243 (N_7243,N_3249,N_1853);
or U7244 (N_7244,N_2729,N_4630);
xnor U7245 (N_7245,N_2415,N_1045);
or U7246 (N_7246,N_4262,N_2153);
xor U7247 (N_7247,N_3026,N_2206);
nor U7248 (N_7248,N_961,N_3513);
nand U7249 (N_7249,N_4160,N_3489);
or U7250 (N_7250,N_772,N_1249);
xnor U7251 (N_7251,N_3371,N_2913);
nand U7252 (N_7252,N_1876,N_2162);
or U7253 (N_7253,N_1473,N_1866);
or U7254 (N_7254,N_4607,N_2652);
xnor U7255 (N_7255,N_1971,N_700);
and U7256 (N_7256,N_4101,N_1216);
and U7257 (N_7257,N_2216,N_3057);
and U7258 (N_7258,N_2791,N_710);
nor U7259 (N_7259,N_1454,N_2040);
or U7260 (N_7260,N_204,N_3218);
nor U7261 (N_7261,N_3523,N_2641);
nor U7262 (N_7262,N_3189,N_4978);
nand U7263 (N_7263,N_3233,N_211);
xor U7264 (N_7264,N_809,N_477);
or U7265 (N_7265,N_3612,N_2725);
xnor U7266 (N_7266,N_4676,N_747);
nor U7267 (N_7267,N_4266,N_3162);
xnor U7268 (N_7268,N_558,N_1980);
xnor U7269 (N_7269,N_3071,N_3429);
nand U7270 (N_7270,N_4593,N_2898);
nand U7271 (N_7271,N_3250,N_1151);
or U7272 (N_7272,N_1609,N_1667);
xor U7273 (N_7273,N_1169,N_3168);
or U7274 (N_7274,N_431,N_1451);
and U7275 (N_7275,N_3517,N_2339);
nor U7276 (N_7276,N_4046,N_1062);
nand U7277 (N_7277,N_177,N_4565);
nor U7278 (N_7278,N_4247,N_4866);
and U7279 (N_7279,N_3702,N_2422);
nand U7280 (N_7280,N_1520,N_3604);
nand U7281 (N_7281,N_888,N_3762);
or U7282 (N_7282,N_4980,N_3735);
or U7283 (N_7283,N_130,N_935);
nor U7284 (N_7284,N_987,N_4559);
nand U7285 (N_7285,N_1840,N_985);
and U7286 (N_7286,N_727,N_1021);
nor U7287 (N_7287,N_1786,N_3654);
nand U7288 (N_7288,N_2650,N_4941);
nand U7289 (N_7289,N_33,N_1547);
nor U7290 (N_7290,N_1228,N_3295);
xnor U7291 (N_7291,N_560,N_2552);
or U7292 (N_7292,N_3933,N_1019);
nand U7293 (N_7293,N_4711,N_194);
xor U7294 (N_7294,N_1005,N_407);
nand U7295 (N_7295,N_2733,N_587);
nand U7296 (N_7296,N_1414,N_163);
nor U7297 (N_7297,N_3351,N_4439);
or U7298 (N_7298,N_1201,N_1027);
or U7299 (N_7299,N_4449,N_2207);
nand U7300 (N_7300,N_2950,N_4009);
and U7301 (N_7301,N_1074,N_4424);
or U7302 (N_7302,N_1148,N_4735);
xor U7303 (N_7303,N_859,N_15);
xor U7304 (N_7304,N_1683,N_4677);
nor U7305 (N_7305,N_241,N_4252);
and U7306 (N_7306,N_2174,N_514);
nor U7307 (N_7307,N_623,N_3560);
nand U7308 (N_7308,N_4903,N_4431);
and U7309 (N_7309,N_3926,N_1440);
or U7310 (N_7310,N_4314,N_2355);
nand U7311 (N_7311,N_1790,N_3325);
and U7312 (N_7312,N_2280,N_1026);
nand U7313 (N_7313,N_3876,N_4741);
nand U7314 (N_7314,N_2540,N_2659);
nand U7315 (N_7315,N_4390,N_4132);
nand U7316 (N_7316,N_3875,N_4115);
nor U7317 (N_7317,N_2273,N_3830);
nor U7318 (N_7318,N_2099,N_1161);
xor U7319 (N_7319,N_3858,N_4374);
xnor U7320 (N_7320,N_4616,N_1232);
and U7321 (N_7321,N_1485,N_2369);
or U7322 (N_7322,N_3105,N_4042);
xor U7323 (N_7323,N_3635,N_3035);
or U7324 (N_7324,N_4443,N_1569);
and U7325 (N_7325,N_2258,N_2706);
nand U7326 (N_7326,N_923,N_1113);
or U7327 (N_7327,N_4323,N_2366);
xnor U7328 (N_7328,N_185,N_387);
and U7329 (N_7329,N_4523,N_217);
or U7330 (N_7330,N_2834,N_199);
xor U7331 (N_7331,N_1013,N_590);
or U7332 (N_7332,N_1421,N_4312);
or U7333 (N_7333,N_1093,N_4851);
and U7334 (N_7334,N_4850,N_815);
nand U7335 (N_7335,N_1823,N_3449);
xor U7336 (N_7336,N_1661,N_3100);
and U7337 (N_7337,N_4470,N_2028);
and U7338 (N_7338,N_4038,N_4726);
nand U7339 (N_7339,N_3747,N_584);
or U7340 (N_7340,N_2243,N_1103);
nand U7341 (N_7341,N_971,N_4448);
and U7342 (N_7342,N_2159,N_1745);
and U7343 (N_7343,N_654,N_4956);
nor U7344 (N_7344,N_4923,N_4076);
nand U7345 (N_7345,N_2660,N_1698);
nor U7346 (N_7346,N_129,N_2793);
xor U7347 (N_7347,N_3758,N_2063);
nand U7348 (N_7348,N_750,N_1427);
xnor U7349 (N_7349,N_1904,N_1224);
nand U7350 (N_7350,N_2284,N_4136);
or U7351 (N_7351,N_3692,N_4989);
xor U7352 (N_7352,N_1562,N_613);
or U7353 (N_7353,N_3644,N_4261);
and U7354 (N_7354,N_21,N_4684);
nor U7355 (N_7355,N_3494,N_591);
or U7356 (N_7356,N_4889,N_1975);
nand U7357 (N_7357,N_3160,N_2246);
and U7358 (N_7358,N_575,N_2390);
nor U7359 (N_7359,N_3674,N_3615);
nand U7360 (N_7360,N_2179,N_1199);
xor U7361 (N_7361,N_4517,N_2203);
nand U7362 (N_7362,N_3683,N_4351);
nand U7363 (N_7363,N_4212,N_4609);
or U7364 (N_7364,N_3987,N_2654);
nor U7365 (N_7365,N_4271,N_196);
and U7366 (N_7366,N_354,N_2701);
or U7367 (N_7367,N_1863,N_3769);
nor U7368 (N_7368,N_877,N_983);
and U7369 (N_7369,N_1469,N_3618);
or U7370 (N_7370,N_1116,N_2703);
nand U7371 (N_7371,N_3807,N_4472);
or U7372 (N_7372,N_339,N_2009);
nand U7373 (N_7373,N_2018,N_368);
xnor U7374 (N_7374,N_4045,N_773);
nor U7375 (N_7375,N_4716,N_2161);
and U7376 (N_7376,N_1096,N_4123);
and U7377 (N_7377,N_2653,N_2869);
xor U7378 (N_7378,N_1885,N_4306);
nor U7379 (N_7379,N_3518,N_3373);
or U7380 (N_7380,N_4082,N_4805);
and U7381 (N_7381,N_2878,N_3165);
and U7382 (N_7382,N_1886,N_77);
and U7383 (N_7383,N_762,N_896);
or U7384 (N_7384,N_2051,N_4223);
or U7385 (N_7385,N_1474,N_1750);
nor U7386 (N_7386,N_4905,N_1850);
nand U7387 (N_7387,N_4248,N_4118);
xor U7388 (N_7388,N_3466,N_3344);
or U7389 (N_7389,N_458,N_594);
or U7390 (N_7390,N_1120,N_2597);
nand U7391 (N_7391,N_4221,N_1109);
nor U7392 (N_7392,N_103,N_854);
and U7393 (N_7393,N_1466,N_4648);
xor U7394 (N_7394,N_249,N_1979);
xnor U7395 (N_7395,N_4295,N_3802);
or U7396 (N_7396,N_2699,N_4036);
nor U7397 (N_7397,N_3713,N_2563);
and U7398 (N_7398,N_4093,N_2663);
nor U7399 (N_7399,N_524,N_3561);
xnor U7400 (N_7400,N_1938,N_4846);
or U7401 (N_7401,N_2514,N_4417);
xnor U7402 (N_7402,N_1404,N_2406);
xnor U7403 (N_7403,N_703,N_3557);
nand U7404 (N_7404,N_3359,N_3840);
nand U7405 (N_7405,N_1805,N_4144);
nor U7406 (N_7406,N_2872,N_3779);
xnor U7407 (N_7407,N_2801,N_4993);
and U7408 (N_7408,N_4427,N_1068);
or U7409 (N_7409,N_1910,N_3535);
and U7410 (N_7410,N_1964,N_4881);
xnor U7411 (N_7411,N_1553,N_3438);
or U7412 (N_7412,N_3880,N_3003);
and U7413 (N_7413,N_1597,N_1911);
nand U7414 (N_7414,N_1694,N_325);
or U7415 (N_7415,N_2312,N_1056);
xor U7416 (N_7416,N_1604,N_2492);
or U7417 (N_7417,N_371,N_1702);
xnor U7418 (N_7418,N_2103,N_2290);
nor U7419 (N_7419,N_4873,N_2384);
or U7420 (N_7420,N_1210,N_3857);
and U7421 (N_7421,N_2100,N_1730);
xnor U7422 (N_7422,N_4091,N_787);
xnor U7423 (N_7423,N_153,N_2674);
or U7424 (N_7424,N_4617,N_1751);
xnor U7425 (N_7425,N_4867,N_2263);
or U7426 (N_7426,N_4877,N_3952);
nand U7427 (N_7427,N_4175,N_126);
xor U7428 (N_7428,N_2839,N_1705);
xnor U7429 (N_7429,N_4992,N_366);
nor U7430 (N_7430,N_2797,N_2856);
xor U7431 (N_7431,N_3417,N_991);
nor U7432 (N_7432,N_4623,N_4945);
nor U7433 (N_7433,N_4148,N_4326);
and U7434 (N_7434,N_2482,N_135);
nor U7435 (N_7435,N_4273,N_2);
nor U7436 (N_7436,N_3787,N_1133);
or U7437 (N_7437,N_4077,N_2507);
nand U7438 (N_7438,N_4397,N_675);
nor U7439 (N_7439,N_3628,N_4601);
and U7440 (N_7440,N_2176,N_2517);
nand U7441 (N_7441,N_1897,N_2225);
xnor U7442 (N_7442,N_4442,N_3902);
or U7443 (N_7443,N_3216,N_4999);
nand U7444 (N_7444,N_2882,N_335);
nor U7445 (N_7445,N_3261,N_2096);
or U7446 (N_7446,N_3598,N_473);
nor U7447 (N_7447,N_3877,N_1059);
or U7448 (N_7448,N_4456,N_3788);
nand U7449 (N_7449,N_2850,N_4786);
nor U7450 (N_7450,N_1936,N_2830);
nor U7451 (N_7451,N_1508,N_4872);
and U7452 (N_7452,N_2947,N_1423);
nor U7453 (N_7453,N_3157,N_2238);
xnor U7454 (N_7454,N_1703,N_1371);
nor U7455 (N_7455,N_657,N_2528);
nand U7456 (N_7456,N_1315,N_4604);
nand U7457 (N_7457,N_1197,N_4254);
and U7458 (N_7458,N_1178,N_3572);
xnor U7459 (N_7459,N_4202,N_3454);
or U7460 (N_7460,N_1278,N_4018);
xor U7461 (N_7461,N_1758,N_615);
nor U7462 (N_7462,N_3196,N_1426);
nor U7463 (N_7463,N_1887,N_1039);
nand U7464 (N_7464,N_3898,N_4126);
nand U7465 (N_7465,N_1128,N_195);
nand U7466 (N_7466,N_977,N_1400);
xor U7467 (N_7467,N_1697,N_1761);
and U7468 (N_7468,N_1078,N_1418);
xor U7469 (N_7469,N_894,N_3529);
or U7470 (N_7470,N_702,N_115);
xor U7471 (N_7471,N_4344,N_1054);
or U7472 (N_7472,N_3526,N_2277);
or U7473 (N_7473,N_3008,N_2820);
or U7474 (N_7474,N_236,N_3188);
nor U7475 (N_7475,N_4645,N_4285);
or U7476 (N_7476,N_3240,N_2774);
or U7477 (N_7477,N_121,N_1259);
and U7478 (N_7478,N_1235,N_4376);
nor U7479 (N_7479,N_2119,N_4382);
or U7480 (N_7480,N_4720,N_3294);
or U7481 (N_7481,N_3488,N_1072);
or U7482 (N_7482,N_1465,N_1594);
xnor U7483 (N_7483,N_446,N_4895);
and U7484 (N_7484,N_1684,N_4124);
nand U7485 (N_7485,N_2344,N_3720);
nor U7486 (N_7486,N_721,N_3045);
nor U7487 (N_7487,N_2979,N_3818);
nand U7488 (N_7488,N_2403,N_294);
nand U7489 (N_7489,N_2680,N_2541);
nand U7490 (N_7490,N_1057,N_258);
nand U7491 (N_7491,N_722,N_1987);
xnor U7492 (N_7492,N_2265,N_224);
or U7493 (N_7493,N_2802,N_3586);
nand U7494 (N_7494,N_1791,N_720);
nor U7495 (N_7495,N_3076,N_1596);
or U7496 (N_7496,N_4868,N_4546);
xor U7497 (N_7497,N_817,N_3110);
and U7498 (N_7498,N_1387,N_1990);
nor U7499 (N_7499,N_2697,N_3343);
xnor U7500 (N_7500,N_1269,N_480);
nor U7501 (N_7501,N_890,N_3679);
nor U7502 (N_7502,N_2004,N_2586);
nand U7503 (N_7503,N_236,N_4851);
nor U7504 (N_7504,N_3484,N_2435);
nand U7505 (N_7505,N_3033,N_2627);
and U7506 (N_7506,N_553,N_3146);
nand U7507 (N_7507,N_2773,N_3291);
or U7508 (N_7508,N_4850,N_4935);
nand U7509 (N_7509,N_1904,N_1295);
nand U7510 (N_7510,N_453,N_2285);
nor U7511 (N_7511,N_1514,N_535);
and U7512 (N_7512,N_1387,N_3626);
and U7513 (N_7513,N_2570,N_2128);
or U7514 (N_7514,N_4219,N_4265);
or U7515 (N_7515,N_1969,N_809);
xnor U7516 (N_7516,N_3749,N_1492);
or U7517 (N_7517,N_3500,N_949);
nor U7518 (N_7518,N_3002,N_2717);
xor U7519 (N_7519,N_289,N_3021);
nor U7520 (N_7520,N_4285,N_2776);
or U7521 (N_7521,N_87,N_3279);
or U7522 (N_7522,N_753,N_4429);
xor U7523 (N_7523,N_2507,N_4959);
or U7524 (N_7524,N_2507,N_4439);
xor U7525 (N_7525,N_2439,N_2450);
xnor U7526 (N_7526,N_41,N_4017);
nand U7527 (N_7527,N_3647,N_2243);
nand U7528 (N_7528,N_674,N_570);
xor U7529 (N_7529,N_2334,N_881);
xor U7530 (N_7530,N_2796,N_1742);
or U7531 (N_7531,N_3612,N_4961);
nor U7532 (N_7532,N_4469,N_2808);
or U7533 (N_7533,N_4878,N_73);
nor U7534 (N_7534,N_4501,N_3562);
or U7535 (N_7535,N_2721,N_2368);
nand U7536 (N_7536,N_1716,N_86);
or U7537 (N_7537,N_275,N_1199);
nand U7538 (N_7538,N_178,N_4120);
nand U7539 (N_7539,N_389,N_4626);
and U7540 (N_7540,N_876,N_895);
nor U7541 (N_7541,N_1856,N_865);
nand U7542 (N_7542,N_1571,N_4642);
and U7543 (N_7543,N_2206,N_4652);
nor U7544 (N_7544,N_1427,N_2672);
nand U7545 (N_7545,N_2710,N_2890);
nand U7546 (N_7546,N_4422,N_1652);
and U7547 (N_7547,N_2287,N_115);
xor U7548 (N_7548,N_1039,N_1766);
nand U7549 (N_7549,N_568,N_3521);
or U7550 (N_7550,N_1820,N_717);
or U7551 (N_7551,N_3080,N_473);
nor U7552 (N_7552,N_1524,N_1517);
nor U7553 (N_7553,N_4732,N_669);
nand U7554 (N_7554,N_2256,N_1456);
and U7555 (N_7555,N_203,N_4185);
nand U7556 (N_7556,N_494,N_1584);
nand U7557 (N_7557,N_4523,N_4862);
nor U7558 (N_7558,N_3545,N_1653);
nor U7559 (N_7559,N_1215,N_1578);
nor U7560 (N_7560,N_1583,N_2068);
and U7561 (N_7561,N_1485,N_373);
or U7562 (N_7562,N_2427,N_4249);
nand U7563 (N_7563,N_3428,N_4685);
nand U7564 (N_7564,N_896,N_2702);
or U7565 (N_7565,N_3432,N_4963);
nor U7566 (N_7566,N_2589,N_346);
nor U7567 (N_7567,N_3170,N_1776);
nand U7568 (N_7568,N_962,N_2700);
nor U7569 (N_7569,N_1370,N_3059);
nor U7570 (N_7570,N_3051,N_2508);
nor U7571 (N_7571,N_3836,N_1343);
and U7572 (N_7572,N_3467,N_4673);
and U7573 (N_7573,N_4477,N_1539);
and U7574 (N_7574,N_2448,N_14);
or U7575 (N_7575,N_3049,N_917);
nand U7576 (N_7576,N_3892,N_3790);
or U7577 (N_7577,N_569,N_1578);
nand U7578 (N_7578,N_3053,N_846);
nor U7579 (N_7579,N_480,N_986);
and U7580 (N_7580,N_379,N_3813);
and U7581 (N_7581,N_2212,N_3215);
nor U7582 (N_7582,N_2043,N_3285);
and U7583 (N_7583,N_1412,N_2564);
or U7584 (N_7584,N_2817,N_429);
nor U7585 (N_7585,N_391,N_1379);
xnor U7586 (N_7586,N_536,N_3314);
and U7587 (N_7587,N_796,N_3673);
and U7588 (N_7588,N_2228,N_3475);
and U7589 (N_7589,N_1069,N_3514);
xnor U7590 (N_7590,N_1382,N_1690);
nand U7591 (N_7591,N_1665,N_2123);
or U7592 (N_7592,N_4437,N_4260);
and U7593 (N_7593,N_2925,N_960);
xnor U7594 (N_7594,N_2531,N_2627);
or U7595 (N_7595,N_4483,N_4893);
nand U7596 (N_7596,N_4541,N_4192);
or U7597 (N_7597,N_1945,N_1322);
xnor U7598 (N_7598,N_1375,N_4920);
or U7599 (N_7599,N_4188,N_152);
or U7600 (N_7600,N_944,N_3981);
and U7601 (N_7601,N_3850,N_1293);
nor U7602 (N_7602,N_2651,N_800);
or U7603 (N_7603,N_555,N_2961);
or U7604 (N_7604,N_3687,N_1833);
and U7605 (N_7605,N_1763,N_2065);
xor U7606 (N_7606,N_973,N_2151);
and U7607 (N_7607,N_4763,N_4043);
xor U7608 (N_7608,N_4490,N_3523);
xnor U7609 (N_7609,N_276,N_1135);
or U7610 (N_7610,N_903,N_1562);
nor U7611 (N_7611,N_1035,N_199);
xnor U7612 (N_7612,N_4185,N_4308);
nand U7613 (N_7613,N_3710,N_4998);
nand U7614 (N_7614,N_1334,N_4638);
xor U7615 (N_7615,N_2154,N_3465);
nor U7616 (N_7616,N_55,N_2415);
and U7617 (N_7617,N_1442,N_697);
nor U7618 (N_7618,N_2488,N_4613);
or U7619 (N_7619,N_4898,N_1693);
nor U7620 (N_7620,N_1988,N_747);
or U7621 (N_7621,N_3426,N_1693);
nor U7622 (N_7622,N_1446,N_2198);
xnor U7623 (N_7623,N_1421,N_1435);
xor U7624 (N_7624,N_1596,N_3837);
nor U7625 (N_7625,N_1334,N_3455);
or U7626 (N_7626,N_2976,N_3975);
nand U7627 (N_7627,N_4626,N_324);
or U7628 (N_7628,N_3578,N_2483);
xnor U7629 (N_7629,N_2834,N_2022);
or U7630 (N_7630,N_1412,N_132);
xnor U7631 (N_7631,N_2402,N_3514);
xor U7632 (N_7632,N_1876,N_782);
xnor U7633 (N_7633,N_4702,N_2404);
or U7634 (N_7634,N_4671,N_789);
and U7635 (N_7635,N_512,N_1706);
or U7636 (N_7636,N_3906,N_1887);
and U7637 (N_7637,N_814,N_3266);
or U7638 (N_7638,N_3616,N_2327);
or U7639 (N_7639,N_577,N_3406);
nand U7640 (N_7640,N_2900,N_4720);
nand U7641 (N_7641,N_1521,N_183);
and U7642 (N_7642,N_3553,N_4623);
xnor U7643 (N_7643,N_3012,N_2753);
nand U7644 (N_7644,N_2569,N_2236);
nor U7645 (N_7645,N_2544,N_3450);
xor U7646 (N_7646,N_4722,N_4571);
and U7647 (N_7647,N_98,N_2834);
nand U7648 (N_7648,N_1129,N_1814);
nand U7649 (N_7649,N_3107,N_4466);
xor U7650 (N_7650,N_2226,N_3296);
xor U7651 (N_7651,N_851,N_3051);
or U7652 (N_7652,N_3577,N_150);
or U7653 (N_7653,N_4983,N_4589);
nor U7654 (N_7654,N_1992,N_276);
nor U7655 (N_7655,N_3508,N_3049);
nor U7656 (N_7656,N_2314,N_2594);
nand U7657 (N_7657,N_3322,N_1570);
nand U7658 (N_7658,N_50,N_1457);
and U7659 (N_7659,N_4977,N_1237);
nand U7660 (N_7660,N_1025,N_3297);
xor U7661 (N_7661,N_1562,N_4497);
nor U7662 (N_7662,N_3095,N_3743);
nor U7663 (N_7663,N_4963,N_341);
nor U7664 (N_7664,N_4056,N_2109);
and U7665 (N_7665,N_4444,N_1386);
and U7666 (N_7666,N_3513,N_3589);
nor U7667 (N_7667,N_3400,N_2936);
nand U7668 (N_7668,N_4573,N_1493);
and U7669 (N_7669,N_3023,N_4311);
or U7670 (N_7670,N_3939,N_3537);
xor U7671 (N_7671,N_2525,N_666);
or U7672 (N_7672,N_1260,N_1266);
or U7673 (N_7673,N_1356,N_1598);
or U7674 (N_7674,N_325,N_3291);
xor U7675 (N_7675,N_4363,N_2573);
or U7676 (N_7676,N_1684,N_4151);
and U7677 (N_7677,N_146,N_337);
or U7678 (N_7678,N_2582,N_1854);
nor U7679 (N_7679,N_4023,N_3921);
and U7680 (N_7680,N_902,N_3914);
nor U7681 (N_7681,N_2693,N_2500);
xor U7682 (N_7682,N_1535,N_4684);
xor U7683 (N_7683,N_3367,N_3701);
nand U7684 (N_7684,N_612,N_4538);
nand U7685 (N_7685,N_611,N_2177);
and U7686 (N_7686,N_1493,N_478);
xor U7687 (N_7687,N_3563,N_1051);
nor U7688 (N_7688,N_1014,N_1154);
nor U7689 (N_7689,N_3743,N_1365);
or U7690 (N_7690,N_1106,N_4102);
nand U7691 (N_7691,N_3273,N_1067);
nand U7692 (N_7692,N_511,N_3550);
xor U7693 (N_7693,N_2283,N_4704);
or U7694 (N_7694,N_1135,N_1295);
nand U7695 (N_7695,N_58,N_944);
xor U7696 (N_7696,N_1144,N_153);
nor U7697 (N_7697,N_3869,N_1973);
or U7698 (N_7698,N_2584,N_2488);
nor U7699 (N_7699,N_3862,N_4723);
or U7700 (N_7700,N_3595,N_2769);
nand U7701 (N_7701,N_2475,N_1766);
or U7702 (N_7702,N_2982,N_2382);
xnor U7703 (N_7703,N_2296,N_2146);
nor U7704 (N_7704,N_2790,N_1370);
and U7705 (N_7705,N_4651,N_2527);
xnor U7706 (N_7706,N_4741,N_1408);
xor U7707 (N_7707,N_4113,N_3112);
or U7708 (N_7708,N_2526,N_3946);
or U7709 (N_7709,N_1767,N_2303);
xnor U7710 (N_7710,N_3491,N_4618);
and U7711 (N_7711,N_408,N_1325);
nand U7712 (N_7712,N_2295,N_1144);
nor U7713 (N_7713,N_1232,N_2745);
xor U7714 (N_7714,N_888,N_3779);
nand U7715 (N_7715,N_4012,N_2528);
or U7716 (N_7716,N_2174,N_3115);
or U7717 (N_7717,N_2032,N_1986);
nor U7718 (N_7718,N_4325,N_459);
or U7719 (N_7719,N_3601,N_1296);
nor U7720 (N_7720,N_236,N_1856);
xnor U7721 (N_7721,N_3534,N_373);
nand U7722 (N_7722,N_975,N_2180);
xnor U7723 (N_7723,N_352,N_894);
nand U7724 (N_7724,N_911,N_1031);
xor U7725 (N_7725,N_2321,N_3625);
nor U7726 (N_7726,N_3017,N_3709);
nor U7727 (N_7727,N_1566,N_2555);
or U7728 (N_7728,N_1752,N_2571);
nor U7729 (N_7729,N_2904,N_3582);
and U7730 (N_7730,N_816,N_777);
nand U7731 (N_7731,N_4689,N_3971);
nand U7732 (N_7732,N_3765,N_2769);
or U7733 (N_7733,N_2496,N_3773);
and U7734 (N_7734,N_50,N_3856);
nor U7735 (N_7735,N_3214,N_3331);
and U7736 (N_7736,N_743,N_4830);
and U7737 (N_7737,N_4051,N_4223);
and U7738 (N_7738,N_401,N_412);
xnor U7739 (N_7739,N_421,N_496);
nand U7740 (N_7740,N_1191,N_3316);
xnor U7741 (N_7741,N_3522,N_4741);
nand U7742 (N_7742,N_4989,N_404);
or U7743 (N_7743,N_4192,N_1084);
and U7744 (N_7744,N_2397,N_3692);
xnor U7745 (N_7745,N_2769,N_693);
nand U7746 (N_7746,N_2919,N_4931);
nor U7747 (N_7747,N_1510,N_3362);
xor U7748 (N_7748,N_4913,N_1202);
and U7749 (N_7749,N_3575,N_1459);
xnor U7750 (N_7750,N_1672,N_4645);
nor U7751 (N_7751,N_1960,N_1801);
nor U7752 (N_7752,N_3243,N_3696);
and U7753 (N_7753,N_1740,N_260);
nand U7754 (N_7754,N_4029,N_2175);
and U7755 (N_7755,N_2788,N_3163);
xor U7756 (N_7756,N_4440,N_3270);
xor U7757 (N_7757,N_4688,N_4562);
or U7758 (N_7758,N_4181,N_3474);
and U7759 (N_7759,N_479,N_467);
xnor U7760 (N_7760,N_305,N_3120);
xor U7761 (N_7761,N_2396,N_4415);
or U7762 (N_7762,N_108,N_866);
xnor U7763 (N_7763,N_2524,N_1492);
and U7764 (N_7764,N_1855,N_2208);
nor U7765 (N_7765,N_3473,N_1419);
or U7766 (N_7766,N_758,N_4649);
or U7767 (N_7767,N_4611,N_2418);
or U7768 (N_7768,N_2830,N_241);
or U7769 (N_7769,N_3446,N_4023);
and U7770 (N_7770,N_2515,N_2028);
and U7771 (N_7771,N_201,N_3223);
xor U7772 (N_7772,N_2978,N_4236);
nor U7773 (N_7773,N_2678,N_3434);
nor U7774 (N_7774,N_2424,N_3511);
nand U7775 (N_7775,N_3663,N_172);
and U7776 (N_7776,N_1187,N_1981);
nand U7777 (N_7777,N_3135,N_1445);
nor U7778 (N_7778,N_1202,N_4007);
xnor U7779 (N_7779,N_4428,N_2907);
or U7780 (N_7780,N_3184,N_1484);
and U7781 (N_7781,N_2193,N_1234);
and U7782 (N_7782,N_3898,N_3566);
nand U7783 (N_7783,N_4551,N_4611);
and U7784 (N_7784,N_2658,N_3450);
and U7785 (N_7785,N_3477,N_2302);
nand U7786 (N_7786,N_3797,N_4590);
and U7787 (N_7787,N_3055,N_4425);
or U7788 (N_7788,N_1618,N_4445);
and U7789 (N_7789,N_448,N_1912);
or U7790 (N_7790,N_3548,N_1951);
or U7791 (N_7791,N_2738,N_2587);
xor U7792 (N_7792,N_1384,N_2275);
or U7793 (N_7793,N_1159,N_1403);
nand U7794 (N_7794,N_3593,N_2723);
nor U7795 (N_7795,N_2859,N_645);
nor U7796 (N_7796,N_4789,N_4176);
nand U7797 (N_7797,N_3691,N_2979);
nor U7798 (N_7798,N_4673,N_4281);
or U7799 (N_7799,N_1190,N_907);
nor U7800 (N_7800,N_3024,N_781);
nand U7801 (N_7801,N_4139,N_1551);
nor U7802 (N_7802,N_4951,N_3786);
and U7803 (N_7803,N_2538,N_277);
and U7804 (N_7804,N_1140,N_638);
and U7805 (N_7805,N_2944,N_4408);
or U7806 (N_7806,N_2171,N_4037);
xnor U7807 (N_7807,N_3589,N_2889);
and U7808 (N_7808,N_3570,N_4853);
nor U7809 (N_7809,N_4065,N_524);
and U7810 (N_7810,N_2783,N_3968);
nor U7811 (N_7811,N_2665,N_3052);
nand U7812 (N_7812,N_1068,N_2336);
and U7813 (N_7813,N_3196,N_2659);
or U7814 (N_7814,N_145,N_727);
nand U7815 (N_7815,N_4321,N_4053);
and U7816 (N_7816,N_2989,N_3069);
xnor U7817 (N_7817,N_2872,N_4962);
xnor U7818 (N_7818,N_1396,N_2856);
xor U7819 (N_7819,N_301,N_2803);
xnor U7820 (N_7820,N_3494,N_1379);
xnor U7821 (N_7821,N_4739,N_4316);
or U7822 (N_7822,N_2926,N_1750);
xor U7823 (N_7823,N_1711,N_3405);
and U7824 (N_7824,N_4941,N_3485);
nand U7825 (N_7825,N_54,N_3688);
nand U7826 (N_7826,N_3752,N_889);
nand U7827 (N_7827,N_2532,N_3771);
xnor U7828 (N_7828,N_1708,N_4748);
nand U7829 (N_7829,N_4731,N_1193);
nor U7830 (N_7830,N_835,N_145);
and U7831 (N_7831,N_4818,N_3528);
nor U7832 (N_7832,N_1854,N_3614);
nor U7833 (N_7833,N_3627,N_2766);
or U7834 (N_7834,N_4255,N_4);
and U7835 (N_7835,N_3002,N_3466);
and U7836 (N_7836,N_2001,N_4132);
or U7837 (N_7837,N_35,N_1462);
or U7838 (N_7838,N_3845,N_4218);
nand U7839 (N_7839,N_1798,N_4346);
and U7840 (N_7840,N_4223,N_686);
nor U7841 (N_7841,N_2271,N_829);
nand U7842 (N_7842,N_4476,N_3604);
and U7843 (N_7843,N_4657,N_3159);
nand U7844 (N_7844,N_218,N_1911);
nand U7845 (N_7845,N_2978,N_1868);
or U7846 (N_7846,N_3055,N_2890);
or U7847 (N_7847,N_534,N_644);
nand U7848 (N_7848,N_4543,N_1411);
nand U7849 (N_7849,N_2287,N_2319);
nand U7850 (N_7850,N_454,N_4681);
nor U7851 (N_7851,N_1853,N_331);
or U7852 (N_7852,N_1540,N_3446);
nand U7853 (N_7853,N_3516,N_747);
nand U7854 (N_7854,N_3604,N_4097);
xnor U7855 (N_7855,N_3330,N_4719);
xnor U7856 (N_7856,N_1228,N_1722);
nand U7857 (N_7857,N_810,N_533);
or U7858 (N_7858,N_3859,N_48);
nor U7859 (N_7859,N_4887,N_1837);
nand U7860 (N_7860,N_2778,N_1897);
and U7861 (N_7861,N_682,N_4010);
and U7862 (N_7862,N_2418,N_1527);
nor U7863 (N_7863,N_2999,N_2677);
nor U7864 (N_7864,N_4350,N_1827);
or U7865 (N_7865,N_4185,N_3911);
and U7866 (N_7866,N_3549,N_2356);
nand U7867 (N_7867,N_2182,N_1367);
or U7868 (N_7868,N_680,N_4349);
nand U7869 (N_7869,N_895,N_41);
nand U7870 (N_7870,N_2468,N_1697);
nand U7871 (N_7871,N_4269,N_2058);
and U7872 (N_7872,N_3977,N_1217);
nand U7873 (N_7873,N_2219,N_2682);
nor U7874 (N_7874,N_1821,N_306);
nand U7875 (N_7875,N_2318,N_1780);
nor U7876 (N_7876,N_2952,N_2367);
or U7877 (N_7877,N_3279,N_1686);
nor U7878 (N_7878,N_85,N_3017);
nand U7879 (N_7879,N_3284,N_1684);
xor U7880 (N_7880,N_3751,N_2473);
or U7881 (N_7881,N_2518,N_826);
nand U7882 (N_7882,N_3962,N_4835);
nor U7883 (N_7883,N_3031,N_891);
nand U7884 (N_7884,N_2566,N_3292);
and U7885 (N_7885,N_1609,N_4589);
or U7886 (N_7886,N_2652,N_4389);
or U7887 (N_7887,N_714,N_572);
xor U7888 (N_7888,N_1159,N_1952);
nand U7889 (N_7889,N_3094,N_3544);
or U7890 (N_7890,N_3296,N_1929);
xnor U7891 (N_7891,N_1322,N_285);
and U7892 (N_7892,N_2018,N_1965);
nor U7893 (N_7893,N_3981,N_3289);
nor U7894 (N_7894,N_955,N_4204);
xor U7895 (N_7895,N_1240,N_4142);
and U7896 (N_7896,N_4818,N_4825);
nand U7897 (N_7897,N_752,N_123);
nor U7898 (N_7898,N_1867,N_2908);
xnor U7899 (N_7899,N_105,N_2279);
and U7900 (N_7900,N_1130,N_3304);
nor U7901 (N_7901,N_679,N_636);
nand U7902 (N_7902,N_2025,N_1981);
nor U7903 (N_7903,N_301,N_4338);
nor U7904 (N_7904,N_4087,N_339);
nor U7905 (N_7905,N_4039,N_204);
or U7906 (N_7906,N_4470,N_3039);
nand U7907 (N_7907,N_4800,N_3243);
nor U7908 (N_7908,N_2374,N_404);
or U7909 (N_7909,N_2615,N_882);
or U7910 (N_7910,N_1602,N_3874);
nor U7911 (N_7911,N_4623,N_4439);
nand U7912 (N_7912,N_2254,N_2217);
and U7913 (N_7913,N_1748,N_1673);
nor U7914 (N_7914,N_3688,N_3895);
nor U7915 (N_7915,N_3881,N_2161);
nor U7916 (N_7916,N_4664,N_1293);
and U7917 (N_7917,N_4663,N_3360);
nand U7918 (N_7918,N_766,N_2620);
nand U7919 (N_7919,N_4506,N_4289);
xor U7920 (N_7920,N_2918,N_3010);
or U7921 (N_7921,N_545,N_3170);
and U7922 (N_7922,N_4264,N_2688);
nand U7923 (N_7923,N_4075,N_2008);
nand U7924 (N_7924,N_1619,N_1172);
nor U7925 (N_7925,N_1764,N_2948);
xor U7926 (N_7926,N_3939,N_1291);
or U7927 (N_7927,N_2692,N_1395);
or U7928 (N_7928,N_1154,N_4715);
nand U7929 (N_7929,N_753,N_4092);
nor U7930 (N_7930,N_2893,N_4357);
or U7931 (N_7931,N_2000,N_304);
or U7932 (N_7932,N_2251,N_2581);
nor U7933 (N_7933,N_1212,N_766);
xnor U7934 (N_7934,N_4277,N_2074);
and U7935 (N_7935,N_4897,N_3930);
and U7936 (N_7936,N_4223,N_3229);
nor U7937 (N_7937,N_682,N_1162);
nor U7938 (N_7938,N_1240,N_56);
and U7939 (N_7939,N_4611,N_729);
and U7940 (N_7940,N_731,N_4749);
xor U7941 (N_7941,N_1207,N_2481);
nor U7942 (N_7942,N_1837,N_2020);
nor U7943 (N_7943,N_3868,N_4030);
nand U7944 (N_7944,N_2251,N_4126);
nand U7945 (N_7945,N_455,N_2165);
nor U7946 (N_7946,N_2588,N_1211);
nor U7947 (N_7947,N_4002,N_2413);
xor U7948 (N_7948,N_4140,N_3131);
and U7949 (N_7949,N_717,N_3107);
xor U7950 (N_7950,N_3511,N_4527);
nor U7951 (N_7951,N_1665,N_4627);
and U7952 (N_7952,N_4972,N_4219);
xnor U7953 (N_7953,N_636,N_941);
nand U7954 (N_7954,N_4752,N_2925);
and U7955 (N_7955,N_3206,N_3582);
or U7956 (N_7956,N_3764,N_4866);
or U7957 (N_7957,N_1996,N_2215);
xor U7958 (N_7958,N_4833,N_4560);
nand U7959 (N_7959,N_2557,N_2221);
or U7960 (N_7960,N_3501,N_3319);
xor U7961 (N_7961,N_3243,N_3393);
or U7962 (N_7962,N_3394,N_3793);
or U7963 (N_7963,N_347,N_4263);
nand U7964 (N_7964,N_2935,N_4077);
and U7965 (N_7965,N_3070,N_4713);
or U7966 (N_7966,N_4142,N_355);
nand U7967 (N_7967,N_3591,N_2929);
xnor U7968 (N_7968,N_2386,N_3390);
or U7969 (N_7969,N_1837,N_261);
and U7970 (N_7970,N_3695,N_1300);
nor U7971 (N_7971,N_2534,N_4916);
nor U7972 (N_7972,N_3272,N_3442);
and U7973 (N_7973,N_4612,N_1140);
nor U7974 (N_7974,N_3443,N_3339);
nand U7975 (N_7975,N_447,N_597);
nand U7976 (N_7976,N_590,N_1984);
xor U7977 (N_7977,N_4555,N_4486);
or U7978 (N_7978,N_1653,N_4341);
and U7979 (N_7979,N_327,N_1037);
nand U7980 (N_7980,N_4043,N_1151);
nand U7981 (N_7981,N_26,N_4858);
xor U7982 (N_7982,N_1551,N_3814);
xor U7983 (N_7983,N_3697,N_2112);
nor U7984 (N_7984,N_4969,N_1816);
xor U7985 (N_7985,N_4245,N_2090);
xor U7986 (N_7986,N_3399,N_3763);
and U7987 (N_7987,N_2580,N_569);
nand U7988 (N_7988,N_1327,N_3266);
or U7989 (N_7989,N_4745,N_2502);
and U7990 (N_7990,N_327,N_3481);
or U7991 (N_7991,N_2213,N_1160);
or U7992 (N_7992,N_1782,N_2439);
nor U7993 (N_7993,N_332,N_1436);
or U7994 (N_7994,N_2418,N_4459);
or U7995 (N_7995,N_2442,N_2806);
nand U7996 (N_7996,N_4194,N_4077);
xor U7997 (N_7997,N_4094,N_2335);
xnor U7998 (N_7998,N_4921,N_1930);
nor U7999 (N_7999,N_241,N_3589);
or U8000 (N_8000,N_342,N_4106);
xnor U8001 (N_8001,N_4311,N_2968);
or U8002 (N_8002,N_2956,N_4021);
nor U8003 (N_8003,N_83,N_3006);
nor U8004 (N_8004,N_3463,N_248);
or U8005 (N_8005,N_2933,N_4557);
nand U8006 (N_8006,N_4924,N_4839);
xnor U8007 (N_8007,N_1249,N_1782);
or U8008 (N_8008,N_1410,N_478);
nand U8009 (N_8009,N_788,N_3284);
nor U8010 (N_8010,N_1762,N_4812);
and U8011 (N_8011,N_1826,N_1515);
nand U8012 (N_8012,N_1909,N_4304);
xor U8013 (N_8013,N_3011,N_4168);
or U8014 (N_8014,N_626,N_338);
or U8015 (N_8015,N_3983,N_1578);
or U8016 (N_8016,N_2912,N_4975);
nor U8017 (N_8017,N_1748,N_4767);
nor U8018 (N_8018,N_4560,N_4526);
xnor U8019 (N_8019,N_1570,N_3437);
nor U8020 (N_8020,N_4256,N_1791);
and U8021 (N_8021,N_4883,N_1452);
or U8022 (N_8022,N_2672,N_3092);
and U8023 (N_8023,N_1431,N_2001);
nand U8024 (N_8024,N_1318,N_3803);
nand U8025 (N_8025,N_2719,N_4132);
nor U8026 (N_8026,N_3559,N_1611);
nor U8027 (N_8027,N_2692,N_2769);
nor U8028 (N_8028,N_4343,N_2547);
nand U8029 (N_8029,N_4160,N_2782);
and U8030 (N_8030,N_2232,N_1739);
and U8031 (N_8031,N_2760,N_4519);
xor U8032 (N_8032,N_2507,N_630);
or U8033 (N_8033,N_1022,N_1444);
nand U8034 (N_8034,N_1053,N_1540);
or U8035 (N_8035,N_405,N_1768);
nand U8036 (N_8036,N_528,N_792);
nand U8037 (N_8037,N_3260,N_1626);
and U8038 (N_8038,N_2406,N_1282);
nor U8039 (N_8039,N_816,N_1762);
nor U8040 (N_8040,N_4931,N_3836);
nand U8041 (N_8041,N_1756,N_1963);
or U8042 (N_8042,N_1535,N_1962);
xnor U8043 (N_8043,N_461,N_1367);
xnor U8044 (N_8044,N_2200,N_698);
nand U8045 (N_8045,N_2864,N_2970);
and U8046 (N_8046,N_3492,N_970);
or U8047 (N_8047,N_433,N_1264);
xnor U8048 (N_8048,N_4808,N_4083);
and U8049 (N_8049,N_2518,N_2324);
nand U8050 (N_8050,N_438,N_4112);
nor U8051 (N_8051,N_1535,N_979);
and U8052 (N_8052,N_282,N_1160);
nor U8053 (N_8053,N_1234,N_4607);
nand U8054 (N_8054,N_4680,N_1500);
xor U8055 (N_8055,N_4250,N_3023);
nand U8056 (N_8056,N_4407,N_2878);
nor U8057 (N_8057,N_4844,N_4792);
nand U8058 (N_8058,N_4941,N_2929);
nor U8059 (N_8059,N_1965,N_4389);
nand U8060 (N_8060,N_3824,N_2492);
nand U8061 (N_8061,N_21,N_3223);
nand U8062 (N_8062,N_1776,N_2078);
nor U8063 (N_8063,N_2154,N_4984);
and U8064 (N_8064,N_4911,N_440);
xnor U8065 (N_8065,N_2984,N_1234);
nor U8066 (N_8066,N_1942,N_4144);
or U8067 (N_8067,N_4664,N_4320);
nor U8068 (N_8068,N_166,N_926);
and U8069 (N_8069,N_3802,N_4553);
and U8070 (N_8070,N_4019,N_449);
and U8071 (N_8071,N_2144,N_2856);
nor U8072 (N_8072,N_1975,N_3282);
and U8073 (N_8073,N_3752,N_883);
nand U8074 (N_8074,N_2807,N_4387);
and U8075 (N_8075,N_3541,N_3329);
xor U8076 (N_8076,N_2005,N_3457);
xor U8077 (N_8077,N_281,N_43);
nor U8078 (N_8078,N_3470,N_1061);
and U8079 (N_8079,N_4,N_2655);
or U8080 (N_8080,N_1673,N_4530);
nand U8081 (N_8081,N_2601,N_1141);
nand U8082 (N_8082,N_1186,N_853);
nand U8083 (N_8083,N_989,N_1373);
and U8084 (N_8084,N_1713,N_2208);
nand U8085 (N_8085,N_2333,N_3957);
nand U8086 (N_8086,N_4266,N_4118);
nor U8087 (N_8087,N_3672,N_115);
and U8088 (N_8088,N_4254,N_2495);
xor U8089 (N_8089,N_1611,N_2558);
xor U8090 (N_8090,N_1669,N_2705);
or U8091 (N_8091,N_385,N_3582);
nand U8092 (N_8092,N_3623,N_3308);
and U8093 (N_8093,N_2408,N_4534);
nand U8094 (N_8094,N_739,N_1967);
nand U8095 (N_8095,N_2428,N_4181);
xnor U8096 (N_8096,N_3195,N_761);
or U8097 (N_8097,N_4472,N_3188);
nand U8098 (N_8098,N_3194,N_1543);
nand U8099 (N_8099,N_4852,N_285);
nand U8100 (N_8100,N_988,N_63);
xor U8101 (N_8101,N_2372,N_2718);
or U8102 (N_8102,N_2631,N_4719);
nor U8103 (N_8103,N_1502,N_3695);
and U8104 (N_8104,N_781,N_4242);
xor U8105 (N_8105,N_11,N_97);
xnor U8106 (N_8106,N_655,N_4155);
nand U8107 (N_8107,N_3910,N_2819);
nor U8108 (N_8108,N_4036,N_2600);
or U8109 (N_8109,N_2766,N_668);
xor U8110 (N_8110,N_1286,N_3738);
xnor U8111 (N_8111,N_4477,N_1473);
xor U8112 (N_8112,N_3503,N_1807);
nor U8113 (N_8113,N_4415,N_2648);
or U8114 (N_8114,N_683,N_4605);
and U8115 (N_8115,N_918,N_4962);
or U8116 (N_8116,N_2757,N_3093);
nor U8117 (N_8117,N_4876,N_1473);
nor U8118 (N_8118,N_4078,N_1144);
nand U8119 (N_8119,N_2768,N_3075);
or U8120 (N_8120,N_968,N_1777);
and U8121 (N_8121,N_448,N_3130);
or U8122 (N_8122,N_211,N_696);
or U8123 (N_8123,N_2330,N_2168);
nand U8124 (N_8124,N_4799,N_541);
or U8125 (N_8125,N_996,N_3467);
xnor U8126 (N_8126,N_3309,N_2308);
nand U8127 (N_8127,N_4005,N_4713);
nand U8128 (N_8128,N_1371,N_2421);
nand U8129 (N_8129,N_959,N_2078);
xor U8130 (N_8130,N_3661,N_4594);
or U8131 (N_8131,N_3643,N_511);
nand U8132 (N_8132,N_2993,N_2326);
xnor U8133 (N_8133,N_3149,N_3314);
nor U8134 (N_8134,N_457,N_904);
or U8135 (N_8135,N_3247,N_11);
or U8136 (N_8136,N_930,N_1964);
nor U8137 (N_8137,N_2280,N_507);
or U8138 (N_8138,N_1433,N_1311);
nor U8139 (N_8139,N_3657,N_4000);
xor U8140 (N_8140,N_973,N_2666);
xor U8141 (N_8141,N_4594,N_2433);
nor U8142 (N_8142,N_1734,N_399);
and U8143 (N_8143,N_79,N_1381);
and U8144 (N_8144,N_3733,N_717);
or U8145 (N_8145,N_1738,N_592);
nand U8146 (N_8146,N_440,N_1242);
and U8147 (N_8147,N_4268,N_2743);
or U8148 (N_8148,N_4224,N_555);
nor U8149 (N_8149,N_4195,N_1377);
nand U8150 (N_8150,N_355,N_2327);
xnor U8151 (N_8151,N_3133,N_2888);
or U8152 (N_8152,N_4437,N_4173);
nand U8153 (N_8153,N_963,N_761);
or U8154 (N_8154,N_1204,N_1674);
nand U8155 (N_8155,N_2843,N_367);
xor U8156 (N_8156,N_4274,N_1855);
nor U8157 (N_8157,N_1999,N_2458);
and U8158 (N_8158,N_1340,N_4950);
nor U8159 (N_8159,N_3219,N_1354);
nand U8160 (N_8160,N_3664,N_4055);
and U8161 (N_8161,N_2034,N_2464);
or U8162 (N_8162,N_413,N_1080);
nand U8163 (N_8163,N_1784,N_4573);
or U8164 (N_8164,N_1253,N_2663);
nor U8165 (N_8165,N_780,N_4907);
and U8166 (N_8166,N_4496,N_904);
nor U8167 (N_8167,N_1251,N_1211);
or U8168 (N_8168,N_4716,N_1676);
nand U8169 (N_8169,N_3940,N_3799);
and U8170 (N_8170,N_527,N_2038);
xnor U8171 (N_8171,N_2918,N_1571);
and U8172 (N_8172,N_52,N_2936);
xnor U8173 (N_8173,N_4238,N_1339);
nor U8174 (N_8174,N_909,N_291);
or U8175 (N_8175,N_929,N_645);
xnor U8176 (N_8176,N_53,N_4481);
or U8177 (N_8177,N_2297,N_4725);
nand U8178 (N_8178,N_675,N_2352);
nor U8179 (N_8179,N_4705,N_2198);
or U8180 (N_8180,N_2523,N_4068);
and U8181 (N_8181,N_1459,N_1678);
or U8182 (N_8182,N_4029,N_4703);
and U8183 (N_8183,N_3035,N_4713);
nor U8184 (N_8184,N_1779,N_4250);
and U8185 (N_8185,N_505,N_750);
and U8186 (N_8186,N_2372,N_4888);
and U8187 (N_8187,N_2686,N_4946);
and U8188 (N_8188,N_3097,N_1897);
nor U8189 (N_8189,N_679,N_2944);
nor U8190 (N_8190,N_3086,N_1346);
and U8191 (N_8191,N_4885,N_3281);
or U8192 (N_8192,N_4608,N_440);
and U8193 (N_8193,N_3354,N_656);
and U8194 (N_8194,N_1314,N_3011);
or U8195 (N_8195,N_3193,N_3253);
nand U8196 (N_8196,N_4377,N_3846);
nor U8197 (N_8197,N_567,N_4100);
nor U8198 (N_8198,N_1540,N_3307);
nor U8199 (N_8199,N_2391,N_4727);
nor U8200 (N_8200,N_2476,N_2124);
and U8201 (N_8201,N_4164,N_1632);
xnor U8202 (N_8202,N_3329,N_3274);
nand U8203 (N_8203,N_2560,N_1584);
nand U8204 (N_8204,N_85,N_3598);
and U8205 (N_8205,N_338,N_694);
and U8206 (N_8206,N_780,N_2467);
nor U8207 (N_8207,N_1513,N_1425);
xor U8208 (N_8208,N_3236,N_4632);
nand U8209 (N_8209,N_3214,N_4084);
nor U8210 (N_8210,N_1466,N_2510);
and U8211 (N_8211,N_2001,N_3782);
xnor U8212 (N_8212,N_1496,N_1063);
or U8213 (N_8213,N_731,N_931);
and U8214 (N_8214,N_1682,N_1672);
and U8215 (N_8215,N_3661,N_331);
xnor U8216 (N_8216,N_2951,N_1801);
and U8217 (N_8217,N_2549,N_2920);
and U8218 (N_8218,N_3494,N_2172);
nor U8219 (N_8219,N_2317,N_464);
nor U8220 (N_8220,N_609,N_3424);
nor U8221 (N_8221,N_2259,N_1353);
and U8222 (N_8222,N_408,N_4350);
or U8223 (N_8223,N_3216,N_2990);
or U8224 (N_8224,N_612,N_4415);
or U8225 (N_8225,N_4260,N_3287);
and U8226 (N_8226,N_314,N_4175);
nand U8227 (N_8227,N_3102,N_3726);
xor U8228 (N_8228,N_4750,N_2241);
nand U8229 (N_8229,N_1480,N_2309);
nand U8230 (N_8230,N_2175,N_3207);
and U8231 (N_8231,N_2375,N_1822);
xnor U8232 (N_8232,N_4214,N_4395);
or U8233 (N_8233,N_3003,N_1085);
and U8234 (N_8234,N_4645,N_230);
nand U8235 (N_8235,N_2171,N_4970);
and U8236 (N_8236,N_3003,N_4248);
and U8237 (N_8237,N_4058,N_589);
nand U8238 (N_8238,N_2844,N_2920);
nor U8239 (N_8239,N_307,N_4155);
and U8240 (N_8240,N_4003,N_1768);
xor U8241 (N_8241,N_3755,N_2924);
xnor U8242 (N_8242,N_3111,N_3793);
and U8243 (N_8243,N_4856,N_1749);
or U8244 (N_8244,N_1218,N_2341);
nand U8245 (N_8245,N_464,N_1269);
nand U8246 (N_8246,N_2597,N_4636);
nand U8247 (N_8247,N_3497,N_2428);
and U8248 (N_8248,N_2772,N_2430);
or U8249 (N_8249,N_2050,N_1003);
xor U8250 (N_8250,N_339,N_3367);
xnor U8251 (N_8251,N_3020,N_1273);
nor U8252 (N_8252,N_3878,N_937);
and U8253 (N_8253,N_4740,N_655);
or U8254 (N_8254,N_4227,N_1922);
nand U8255 (N_8255,N_602,N_2144);
and U8256 (N_8256,N_3394,N_3151);
nor U8257 (N_8257,N_2949,N_2228);
nor U8258 (N_8258,N_1653,N_802);
or U8259 (N_8259,N_576,N_1210);
nand U8260 (N_8260,N_4882,N_335);
and U8261 (N_8261,N_1790,N_428);
nand U8262 (N_8262,N_1748,N_294);
xnor U8263 (N_8263,N_3665,N_297);
xor U8264 (N_8264,N_2076,N_508);
and U8265 (N_8265,N_3079,N_3356);
xnor U8266 (N_8266,N_2541,N_4245);
or U8267 (N_8267,N_308,N_972);
or U8268 (N_8268,N_3488,N_2982);
or U8269 (N_8269,N_87,N_1472);
xor U8270 (N_8270,N_45,N_1036);
xnor U8271 (N_8271,N_2048,N_2256);
and U8272 (N_8272,N_223,N_4623);
xnor U8273 (N_8273,N_2787,N_2169);
nor U8274 (N_8274,N_657,N_2703);
or U8275 (N_8275,N_3522,N_4259);
nand U8276 (N_8276,N_1266,N_2546);
or U8277 (N_8277,N_2598,N_1757);
xor U8278 (N_8278,N_1907,N_2384);
xor U8279 (N_8279,N_3945,N_83);
and U8280 (N_8280,N_3702,N_3511);
nand U8281 (N_8281,N_1472,N_4888);
xnor U8282 (N_8282,N_2275,N_4659);
nor U8283 (N_8283,N_188,N_2320);
xor U8284 (N_8284,N_870,N_1344);
nand U8285 (N_8285,N_3314,N_3227);
xor U8286 (N_8286,N_3692,N_4169);
xnor U8287 (N_8287,N_2793,N_4230);
or U8288 (N_8288,N_605,N_919);
and U8289 (N_8289,N_145,N_4016);
xor U8290 (N_8290,N_4081,N_3830);
or U8291 (N_8291,N_3255,N_455);
and U8292 (N_8292,N_4031,N_2241);
nand U8293 (N_8293,N_3569,N_3493);
and U8294 (N_8294,N_4091,N_4348);
nor U8295 (N_8295,N_2781,N_2465);
xor U8296 (N_8296,N_1760,N_1549);
and U8297 (N_8297,N_3455,N_3319);
nor U8298 (N_8298,N_112,N_856);
or U8299 (N_8299,N_3317,N_2029);
and U8300 (N_8300,N_1316,N_4481);
nand U8301 (N_8301,N_1295,N_4284);
xor U8302 (N_8302,N_4160,N_1396);
nand U8303 (N_8303,N_2606,N_845);
xor U8304 (N_8304,N_493,N_1942);
and U8305 (N_8305,N_1574,N_1760);
and U8306 (N_8306,N_2167,N_1863);
xor U8307 (N_8307,N_2974,N_566);
nand U8308 (N_8308,N_2451,N_791);
and U8309 (N_8309,N_3715,N_4972);
or U8310 (N_8310,N_1103,N_1746);
nor U8311 (N_8311,N_1042,N_4421);
nor U8312 (N_8312,N_3617,N_4851);
nand U8313 (N_8313,N_352,N_1440);
and U8314 (N_8314,N_3507,N_3898);
xnor U8315 (N_8315,N_1009,N_3761);
or U8316 (N_8316,N_497,N_1504);
nand U8317 (N_8317,N_4715,N_3960);
nor U8318 (N_8318,N_2805,N_1334);
and U8319 (N_8319,N_1320,N_1078);
xnor U8320 (N_8320,N_1804,N_2190);
and U8321 (N_8321,N_773,N_3436);
and U8322 (N_8322,N_4733,N_525);
or U8323 (N_8323,N_2868,N_18);
and U8324 (N_8324,N_1363,N_2456);
nor U8325 (N_8325,N_2787,N_3266);
nor U8326 (N_8326,N_793,N_3380);
or U8327 (N_8327,N_1360,N_3909);
and U8328 (N_8328,N_3621,N_4931);
and U8329 (N_8329,N_4695,N_545);
nand U8330 (N_8330,N_4448,N_4500);
nor U8331 (N_8331,N_4543,N_589);
nor U8332 (N_8332,N_2485,N_2434);
and U8333 (N_8333,N_3548,N_4539);
nor U8334 (N_8334,N_1926,N_2154);
nor U8335 (N_8335,N_1251,N_730);
nand U8336 (N_8336,N_4279,N_3402);
or U8337 (N_8337,N_3590,N_3503);
nor U8338 (N_8338,N_1977,N_3892);
nor U8339 (N_8339,N_760,N_594);
nand U8340 (N_8340,N_103,N_4537);
xor U8341 (N_8341,N_2493,N_2692);
xor U8342 (N_8342,N_3143,N_3896);
or U8343 (N_8343,N_3504,N_1315);
xor U8344 (N_8344,N_216,N_3314);
nor U8345 (N_8345,N_5,N_2375);
xor U8346 (N_8346,N_2258,N_2392);
or U8347 (N_8347,N_3716,N_4633);
xnor U8348 (N_8348,N_3140,N_1141);
and U8349 (N_8349,N_3012,N_2304);
nand U8350 (N_8350,N_3719,N_1656);
nand U8351 (N_8351,N_372,N_2713);
and U8352 (N_8352,N_4325,N_869);
and U8353 (N_8353,N_1711,N_105);
and U8354 (N_8354,N_4183,N_767);
or U8355 (N_8355,N_1196,N_1972);
or U8356 (N_8356,N_747,N_3072);
and U8357 (N_8357,N_3204,N_1559);
nand U8358 (N_8358,N_1753,N_3813);
or U8359 (N_8359,N_57,N_3035);
nor U8360 (N_8360,N_4130,N_2107);
nand U8361 (N_8361,N_4688,N_517);
and U8362 (N_8362,N_2885,N_4775);
nor U8363 (N_8363,N_28,N_1322);
nor U8364 (N_8364,N_952,N_266);
nand U8365 (N_8365,N_3135,N_4674);
and U8366 (N_8366,N_578,N_746);
nand U8367 (N_8367,N_551,N_4641);
nand U8368 (N_8368,N_662,N_140);
nand U8369 (N_8369,N_1121,N_4751);
or U8370 (N_8370,N_14,N_4006);
and U8371 (N_8371,N_2397,N_1604);
nor U8372 (N_8372,N_1128,N_3163);
nand U8373 (N_8373,N_1982,N_1354);
and U8374 (N_8374,N_867,N_2309);
nand U8375 (N_8375,N_2104,N_2253);
or U8376 (N_8376,N_569,N_4440);
nand U8377 (N_8377,N_4910,N_3524);
nor U8378 (N_8378,N_1878,N_3816);
nor U8379 (N_8379,N_3206,N_1367);
or U8380 (N_8380,N_3840,N_1385);
nand U8381 (N_8381,N_1864,N_2319);
and U8382 (N_8382,N_270,N_3651);
nand U8383 (N_8383,N_2301,N_4053);
nand U8384 (N_8384,N_3042,N_4258);
or U8385 (N_8385,N_659,N_92);
nor U8386 (N_8386,N_3079,N_3824);
nor U8387 (N_8387,N_2066,N_3834);
nor U8388 (N_8388,N_1559,N_310);
and U8389 (N_8389,N_3662,N_2689);
and U8390 (N_8390,N_440,N_2052);
and U8391 (N_8391,N_4886,N_2812);
nand U8392 (N_8392,N_4573,N_3057);
and U8393 (N_8393,N_4319,N_2381);
or U8394 (N_8394,N_500,N_893);
nand U8395 (N_8395,N_1341,N_2988);
nand U8396 (N_8396,N_1621,N_162);
nand U8397 (N_8397,N_969,N_898);
and U8398 (N_8398,N_1772,N_1681);
nor U8399 (N_8399,N_4426,N_3777);
and U8400 (N_8400,N_627,N_3556);
nand U8401 (N_8401,N_4050,N_4751);
xor U8402 (N_8402,N_1339,N_4661);
xor U8403 (N_8403,N_516,N_3724);
or U8404 (N_8404,N_4482,N_28);
nand U8405 (N_8405,N_3543,N_2668);
or U8406 (N_8406,N_2606,N_576);
nor U8407 (N_8407,N_3681,N_2101);
nand U8408 (N_8408,N_1348,N_3290);
nor U8409 (N_8409,N_36,N_974);
or U8410 (N_8410,N_3183,N_3187);
nor U8411 (N_8411,N_2163,N_1221);
or U8412 (N_8412,N_4959,N_600);
nor U8413 (N_8413,N_3922,N_206);
and U8414 (N_8414,N_35,N_3893);
nand U8415 (N_8415,N_881,N_2544);
nand U8416 (N_8416,N_4946,N_3134);
and U8417 (N_8417,N_4095,N_4920);
xor U8418 (N_8418,N_2686,N_2526);
or U8419 (N_8419,N_11,N_2310);
and U8420 (N_8420,N_2873,N_52);
xnor U8421 (N_8421,N_672,N_3694);
or U8422 (N_8422,N_3735,N_1894);
nand U8423 (N_8423,N_1395,N_3617);
nand U8424 (N_8424,N_579,N_749);
xnor U8425 (N_8425,N_4967,N_473);
and U8426 (N_8426,N_347,N_2746);
xnor U8427 (N_8427,N_2379,N_2476);
and U8428 (N_8428,N_4271,N_3819);
xnor U8429 (N_8429,N_2053,N_1631);
and U8430 (N_8430,N_246,N_300);
and U8431 (N_8431,N_872,N_4705);
xor U8432 (N_8432,N_4585,N_1362);
nand U8433 (N_8433,N_1030,N_1577);
xor U8434 (N_8434,N_190,N_3686);
nor U8435 (N_8435,N_4579,N_3168);
and U8436 (N_8436,N_2800,N_2273);
nand U8437 (N_8437,N_3262,N_1606);
and U8438 (N_8438,N_912,N_4502);
nor U8439 (N_8439,N_3375,N_1649);
nor U8440 (N_8440,N_3195,N_3529);
nor U8441 (N_8441,N_1919,N_3584);
and U8442 (N_8442,N_3950,N_436);
or U8443 (N_8443,N_4514,N_4833);
nand U8444 (N_8444,N_4295,N_4953);
or U8445 (N_8445,N_1386,N_2863);
or U8446 (N_8446,N_3073,N_1932);
and U8447 (N_8447,N_2064,N_3399);
nand U8448 (N_8448,N_2023,N_4098);
and U8449 (N_8449,N_90,N_846);
or U8450 (N_8450,N_376,N_362);
and U8451 (N_8451,N_2887,N_2029);
xnor U8452 (N_8452,N_4087,N_4470);
and U8453 (N_8453,N_475,N_1671);
or U8454 (N_8454,N_1355,N_2446);
nor U8455 (N_8455,N_2113,N_2798);
nand U8456 (N_8456,N_4555,N_1200);
nand U8457 (N_8457,N_4367,N_4817);
xnor U8458 (N_8458,N_1929,N_1237);
or U8459 (N_8459,N_4564,N_3159);
nand U8460 (N_8460,N_126,N_1406);
or U8461 (N_8461,N_285,N_4478);
and U8462 (N_8462,N_1708,N_1257);
nor U8463 (N_8463,N_4894,N_3124);
nor U8464 (N_8464,N_1568,N_2957);
and U8465 (N_8465,N_3352,N_765);
xnor U8466 (N_8466,N_1981,N_1367);
nand U8467 (N_8467,N_2977,N_4793);
or U8468 (N_8468,N_483,N_2859);
and U8469 (N_8469,N_1175,N_2421);
nor U8470 (N_8470,N_1069,N_1867);
or U8471 (N_8471,N_4242,N_3555);
nor U8472 (N_8472,N_1013,N_474);
nand U8473 (N_8473,N_2251,N_4273);
nor U8474 (N_8474,N_57,N_1610);
and U8475 (N_8475,N_3945,N_121);
or U8476 (N_8476,N_4153,N_3294);
or U8477 (N_8477,N_1350,N_305);
or U8478 (N_8478,N_2732,N_1372);
and U8479 (N_8479,N_3495,N_4203);
nor U8480 (N_8480,N_441,N_2302);
and U8481 (N_8481,N_1987,N_4583);
and U8482 (N_8482,N_1912,N_1692);
xor U8483 (N_8483,N_1244,N_2463);
or U8484 (N_8484,N_4464,N_4815);
and U8485 (N_8485,N_1452,N_1699);
xnor U8486 (N_8486,N_3825,N_696);
and U8487 (N_8487,N_2037,N_1846);
or U8488 (N_8488,N_2755,N_354);
or U8489 (N_8489,N_2129,N_3767);
and U8490 (N_8490,N_2866,N_2145);
xnor U8491 (N_8491,N_1544,N_2587);
and U8492 (N_8492,N_4399,N_2147);
xor U8493 (N_8493,N_4694,N_598);
and U8494 (N_8494,N_2342,N_8);
nand U8495 (N_8495,N_4116,N_3526);
nand U8496 (N_8496,N_2612,N_50);
nor U8497 (N_8497,N_4144,N_4948);
xor U8498 (N_8498,N_2497,N_4076);
xor U8499 (N_8499,N_2285,N_801);
xor U8500 (N_8500,N_1616,N_360);
or U8501 (N_8501,N_1167,N_4400);
and U8502 (N_8502,N_533,N_980);
nor U8503 (N_8503,N_4142,N_4005);
nor U8504 (N_8504,N_2080,N_4051);
or U8505 (N_8505,N_3561,N_1719);
or U8506 (N_8506,N_4731,N_2491);
nor U8507 (N_8507,N_674,N_3405);
nor U8508 (N_8508,N_73,N_2242);
or U8509 (N_8509,N_2336,N_2608);
nand U8510 (N_8510,N_4278,N_1841);
nand U8511 (N_8511,N_369,N_1688);
xor U8512 (N_8512,N_3531,N_522);
and U8513 (N_8513,N_2961,N_4073);
and U8514 (N_8514,N_4481,N_4657);
xnor U8515 (N_8515,N_3090,N_4806);
or U8516 (N_8516,N_3060,N_655);
nor U8517 (N_8517,N_4176,N_3578);
or U8518 (N_8518,N_285,N_1601);
and U8519 (N_8519,N_1889,N_2358);
or U8520 (N_8520,N_1842,N_20);
nand U8521 (N_8521,N_4499,N_590);
nor U8522 (N_8522,N_1866,N_3996);
nor U8523 (N_8523,N_2602,N_774);
nor U8524 (N_8524,N_4126,N_2898);
and U8525 (N_8525,N_4104,N_4990);
xor U8526 (N_8526,N_3832,N_4239);
or U8527 (N_8527,N_2896,N_3300);
xor U8528 (N_8528,N_4164,N_3381);
xor U8529 (N_8529,N_4232,N_2207);
and U8530 (N_8530,N_4399,N_292);
nor U8531 (N_8531,N_3348,N_3243);
xor U8532 (N_8532,N_1990,N_3981);
nor U8533 (N_8533,N_902,N_2153);
and U8534 (N_8534,N_2904,N_68);
and U8535 (N_8535,N_279,N_614);
xnor U8536 (N_8536,N_3102,N_1156);
nor U8537 (N_8537,N_2676,N_3228);
and U8538 (N_8538,N_3788,N_2530);
xnor U8539 (N_8539,N_3404,N_2662);
nand U8540 (N_8540,N_2409,N_4769);
xor U8541 (N_8541,N_971,N_4893);
and U8542 (N_8542,N_1148,N_3019);
or U8543 (N_8543,N_4325,N_3311);
nand U8544 (N_8544,N_4463,N_4506);
nor U8545 (N_8545,N_4332,N_2808);
xnor U8546 (N_8546,N_3255,N_4990);
and U8547 (N_8547,N_3529,N_3994);
or U8548 (N_8548,N_3410,N_664);
and U8549 (N_8549,N_3435,N_4344);
xor U8550 (N_8550,N_4108,N_2221);
and U8551 (N_8551,N_755,N_1232);
or U8552 (N_8552,N_4436,N_4092);
xnor U8553 (N_8553,N_4738,N_4014);
and U8554 (N_8554,N_837,N_2151);
xor U8555 (N_8555,N_4163,N_1454);
and U8556 (N_8556,N_3271,N_580);
xnor U8557 (N_8557,N_2203,N_4735);
nor U8558 (N_8558,N_1538,N_4913);
nor U8559 (N_8559,N_404,N_46);
nand U8560 (N_8560,N_4589,N_205);
or U8561 (N_8561,N_4366,N_579);
nand U8562 (N_8562,N_2811,N_4804);
xnor U8563 (N_8563,N_270,N_3168);
and U8564 (N_8564,N_2274,N_3722);
nor U8565 (N_8565,N_3178,N_427);
nor U8566 (N_8566,N_3074,N_2670);
or U8567 (N_8567,N_3340,N_256);
or U8568 (N_8568,N_4041,N_994);
and U8569 (N_8569,N_2721,N_3889);
or U8570 (N_8570,N_736,N_4870);
nand U8571 (N_8571,N_431,N_3382);
or U8572 (N_8572,N_2542,N_2963);
nand U8573 (N_8573,N_2787,N_2846);
and U8574 (N_8574,N_2441,N_3761);
nand U8575 (N_8575,N_2174,N_4382);
nand U8576 (N_8576,N_4509,N_3865);
nand U8577 (N_8577,N_4265,N_2484);
nor U8578 (N_8578,N_2770,N_3276);
nand U8579 (N_8579,N_2363,N_3012);
and U8580 (N_8580,N_3857,N_2839);
nand U8581 (N_8581,N_1065,N_3852);
and U8582 (N_8582,N_1096,N_2567);
nand U8583 (N_8583,N_2889,N_323);
nand U8584 (N_8584,N_4118,N_3021);
or U8585 (N_8585,N_2946,N_1386);
or U8586 (N_8586,N_1644,N_4016);
nor U8587 (N_8587,N_3476,N_2792);
nand U8588 (N_8588,N_1065,N_2536);
or U8589 (N_8589,N_4570,N_724);
nor U8590 (N_8590,N_3628,N_1498);
xnor U8591 (N_8591,N_2033,N_2385);
or U8592 (N_8592,N_4088,N_527);
nand U8593 (N_8593,N_3570,N_1912);
nand U8594 (N_8594,N_3774,N_468);
and U8595 (N_8595,N_889,N_3711);
nand U8596 (N_8596,N_3336,N_843);
or U8597 (N_8597,N_4845,N_2629);
nand U8598 (N_8598,N_4034,N_4953);
and U8599 (N_8599,N_1550,N_2039);
nor U8600 (N_8600,N_1655,N_93);
and U8601 (N_8601,N_833,N_1420);
nor U8602 (N_8602,N_1286,N_3506);
xor U8603 (N_8603,N_540,N_3240);
nor U8604 (N_8604,N_784,N_358);
nand U8605 (N_8605,N_1638,N_2527);
xor U8606 (N_8606,N_1130,N_1444);
and U8607 (N_8607,N_936,N_342);
and U8608 (N_8608,N_3214,N_2436);
or U8609 (N_8609,N_4793,N_1631);
xnor U8610 (N_8610,N_932,N_3392);
xnor U8611 (N_8611,N_4253,N_671);
and U8612 (N_8612,N_20,N_2447);
xnor U8613 (N_8613,N_4481,N_3474);
nor U8614 (N_8614,N_1744,N_24);
nand U8615 (N_8615,N_1507,N_4483);
and U8616 (N_8616,N_3014,N_2897);
or U8617 (N_8617,N_2980,N_680);
and U8618 (N_8618,N_4949,N_3);
and U8619 (N_8619,N_1750,N_4166);
nand U8620 (N_8620,N_901,N_1257);
or U8621 (N_8621,N_2316,N_1037);
nand U8622 (N_8622,N_2709,N_405);
and U8623 (N_8623,N_4239,N_1425);
and U8624 (N_8624,N_750,N_1728);
and U8625 (N_8625,N_4151,N_3603);
xnor U8626 (N_8626,N_3076,N_4541);
nor U8627 (N_8627,N_448,N_2498);
and U8628 (N_8628,N_3651,N_4339);
nand U8629 (N_8629,N_4764,N_3872);
xor U8630 (N_8630,N_2346,N_884);
and U8631 (N_8631,N_3636,N_1798);
xor U8632 (N_8632,N_2572,N_776);
or U8633 (N_8633,N_4403,N_259);
xor U8634 (N_8634,N_4400,N_3623);
and U8635 (N_8635,N_3624,N_4857);
nor U8636 (N_8636,N_1804,N_943);
or U8637 (N_8637,N_16,N_1364);
or U8638 (N_8638,N_1293,N_4795);
xnor U8639 (N_8639,N_2781,N_1904);
nand U8640 (N_8640,N_4192,N_3859);
nand U8641 (N_8641,N_1331,N_3975);
nor U8642 (N_8642,N_1580,N_2056);
xnor U8643 (N_8643,N_0,N_2436);
or U8644 (N_8644,N_4331,N_4399);
nor U8645 (N_8645,N_4688,N_129);
and U8646 (N_8646,N_1160,N_2238);
nand U8647 (N_8647,N_752,N_4332);
xnor U8648 (N_8648,N_1719,N_322);
xnor U8649 (N_8649,N_1585,N_3408);
or U8650 (N_8650,N_3343,N_839);
or U8651 (N_8651,N_3685,N_2924);
and U8652 (N_8652,N_273,N_3057);
and U8653 (N_8653,N_1983,N_3016);
nor U8654 (N_8654,N_2537,N_4334);
nor U8655 (N_8655,N_3852,N_4595);
nand U8656 (N_8656,N_3271,N_1527);
nand U8657 (N_8657,N_1305,N_3143);
nor U8658 (N_8658,N_1052,N_4792);
and U8659 (N_8659,N_2648,N_3573);
xor U8660 (N_8660,N_3107,N_3801);
nor U8661 (N_8661,N_4693,N_2711);
nand U8662 (N_8662,N_4824,N_4733);
or U8663 (N_8663,N_518,N_3894);
nor U8664 (N_8664,N_772,N_2526);
nand U8665 (N_8665,N_2728,N_3024);
nor U8666 (N_8666,N_2073,N_3058);
and U8667 (N_8667,N_785,N_4761);
xor U8668 (N_8668,N_4408,N_52);
nor U8669 (N_8669,N_3896,N_1115);
nand U8670 (N_8670,N_3984,N_2514);
or U8671 (N_8671,N_3126,N_3689);
or U8672 (N_8672,N_148,N_1077);
nor U8673 (N_8673,N_553,N_3414);
nand U8674 (N_8674,N_1735,N_3186);
or U8675 (N_8675,N_4492,N_1555);
xnor U8676 (N_8676,N_3000,N_4312);
and U8677 (N_8677,N_3924,N_3578);
xnor U8678 (N_8678,N_3023,N_1553);
nand U8679 (N_8679,N_1324,N_4323);
xnor U8680 (N_8680,N_3304,N_157);
or U8681 (N_8681,N_3615,N_3460);
xnor U8682 (N_8682,N_2401,N_1431);
and U8683 (N_8683,N_3334,N_3741);
and U8684 (N_8684,N_2641,N_352);
and U8685 (N_8685,N_4296,N_2821);
or U8686 (N_8686,N_2992,N_2030);
and U8687 (N_8687,N_4170,N_4992);
or U8688 (N_8688,N_2452,N_3527);
nand U8689 (N_8689,N_4168,N_3111);
or U8690 (N_8690,N_642,N_3235);
or U8691 (N_8691,N_4087,N_774);
and U8692 (N_8692,N_2244,N_258);
nand U8693 (N_8693,N_3547,N_10);
xnor U8694 (N_8694,N_1036,N_2481);
and U8695 (N_8695,N_4310,N_4820);
or U8696 (N_8696,N_560,N_1429);
or U8697 (N_8697,N_3564,N_466);
nand U8698 (N_8698,N_3412,N_2608);
or U8699 (N_8699,N_1452,N_1203);
or U8700 (N_8700,N_2978,N_4845);
and U8701 (N_8701,N_541,N_4963);
xnor U8702 (N_8702,N_2133,N_4950);
xnor U8703 (N_8703,N_3104,N_2349);
nor U8704 (N_8704,N_2473,N_4546);
or U8705 (N_8705,N_1640,N_3859);
xnor U8706 (N_8706,N_236,N_538);
or U8707 (N_8707,N_504,N_4431);
nand U8708 (N_8708,N_3738,N_4199);
xnor U8709 (N_8709,N_4225,N_2636);
or U8710 (N_8710,N_4905,N_375);
xor U8711 (N_8711,N_2925,N_956);
nor U8712 (N_8712,N_4462,N_4051);
or U8713 (N_8713,N_2462,N_2914);
and U8714 (N_8714,N_1923,N_4716);
nor U8715 (N_8715,N_4147,N_473);
nor U8716 (N_8716,N_2179,N_3766);
xor U8717 (N_8717,N_59,N_789);
nand U8718 (N_8718,N_1845,N_3785);
nor U8719 (N_8719,N_3185,N_2230);
xnor U8720 (N_8720,N_1479,N_4390);
and U8721 (N_8721,N_644,N_3830);
and U8722 (N_8722,N_3404,N_919);
nor U8723 (N_8723,N_4299,N_2200);
nor U8724 (N_8724,N_1471,N_3786);
or U8725 (N_8725,N_4943,N_3555);
xor U8726 (N_8726,N_2229,N_4497);
nor U8727 (N_8727,N_3697,N_3548);
and U8728 (N_8728,N_149,N_4819);
and U8729 (N_8729,N_2227,N_3892);
nand U8730 (N_8730,N_4038,N_3235);
or U8731 (N_8731,N_3899,N_627);
xor U8732 (N_8732,N_155,N_3359);
xnor U8733 (N_8733,N_4614,N_4870);
nor U8734 (N_8734,N_1539,N_203);
nand U8735 (N_8735,N_585,N_1369);
nor U8736 (N_8736,N_1689,N_2113);
or U8737 (N_8737,N_1397,N_2923);
nor U8738 (N_8738,N_2005,N_2075);
and U8739 (N_8739,N_549,N_1974);
and U8740 (N_8740,N_2178,N_2197);
xnor U8741 (N_8741,N_3119,N_4082);
nand U8742 (N_8742,N_84,N_44);
and U8743 (N_8743,N_3146,N_4473);
and U8744 (N_8744,N_2761,N_3813);
nor U8745 (N_8745,N_59,N_1758);
or U8746 (N_8746,N_3242,N_357);
and U8747 (N_8747,N_2886,N_2811);
xnor U8748 (N_8748,N_3982,N_3510);
nand U8749 (N_8749,N_950,N_1268);
xnor U8750 (N_8750,N_3980,N_4362);
nand U8751 (N_8751,N_3088,N_4150);
and U8752 (N_8752,N_576,N_4337);
nor U8753 (N_8753,N_3153,N_4362);
or U8754 (N_8754,N_35,N_1760);
and U8755 (N_8755,N_3906,N_226);
nor U8756 (N_8756,N_3685,N_1784);
nand U8757 (N_8757,N_1734,N_2688);
xor U8758 (N_8758,N_2719,N_610);
and U8759 (N_8759,N_4751,N_442);
and U8760 (N_8760,N_2440,N_3713);
nor U8761 (N_8761,N_1498,N_1030);
xor U8762 (N_8762,N_774,N_2575);
and U8763 (N_8763,N_54,N_1958);
xnor U8764 (N_8764,N_1453,N_2868);
nor U8765 (N_8765,N_185,N_4004);
xor U8766 (N_8766,N_551,N_1232);
nor U8767 (N_8767,N_1240,N_3020);
nor U8768 (N_8768,N_1885,N_3445);
or U8769 (N_8769,N_684,N_3549);
nor U8770 (N_8770,N_3808,N_3717);
nand U8771 (N_8771,N_4623,N_715);
or U8772 (N_8772,N_4292,N_4469);
and U8773 (N_8773,N_2246,N_3647);
nor U8774 (N_8774,N_2794,N_1263);
xnor U8775 (N_8775,N_973,N_3182);
or U8776 (N_8776,N_2311,N_4576);
and U8777 (N_8777,N_290,N_2044);
xor U8778 (N_8778,N_4113,N_3203);
nand U8779 (N_8779,N_4305,N_4973);
or U8780 (N_8780,N_8,N_1930);
or U8781 (N_8781,N_4521,N_196);
nand U8782 (N_8782,N_81,N_2421);
nand U8783 (N_8783,N_2226,N_3953);
nor U8784 (N_8784,N_4898,N_1423);
nand U8785 (N_8785,N_3726,N_549);
nor U8786 (N_8786,N_3125,N_4965);
and U8787 (N_8787,N_2554,N_3870);
and U8788 (N_8788,N_2521,N_2437);
and U8789 (N_8789,N_4590,N_452);
and U8790 (N_8790,N_4962,N_4383);
and U8791 (N_8791,N_840,N_3325);
xnor U8792 (N_8792,N_4908,N_809);
xor U8793 (N_8793,N_2110,N_1063);
xor U8794 (N_8794,N_3520,N_4760);
or U8795 (N_8795,N_4438,N_276);
nor U8796 (N_8796,N_815,N_972);
nand U8797 (N_8797,N_2898,N_1309);
xor U8798 (N_8798,N_1411,N_1712);
and U8799 (N_8799,N_77,N_2585);
xnor U8800 (N_8800,N_4988,N_2289);
xnor U8801 (N_8801,N_4646,N_480);
nand U8802 (N_8802,N_1173,N_3061);
and U8803 (N_8803,N_1104,N_1826);
nand U8804 (N_8804,N_196,N_2555);
xnor U8805 (N_8805,N_4007,N_4159);
nor U8806 (N_8806,N_2305,N_2312);
nor U8807 (N_8807,N_2347,N_1);
and U8808 (N_8808,N_941,N_3375);
nor U8809 (N_8809,N_368,N_4822);
nor U8810 (N_8810,N_4374,N_2636);
nand U8811 (N_8811,N_4042,N_1804);
nand U8812 (N_8812,N_669,N_2532);
or U8813 (N_8813,N_1997,N_4644);
nand U8814 (N_8814,N_1967,N_4082);
nor U8815 (N_8815,N_2776,N_655);
nand U8816 (N_8816,N_3116,N_1892);
nand U8817 (N_8817,N_236,N_3682);
xor U8818 (N_8818,N_2140,N_4252);
nand U8819 (N_8819,N_3433,N_325);
or U8820 (N_8820,N_3488,N_3588);
nor U8821 (N_8821,N_1459,N_244);
xnor U8822 (N_8822,N_4342,N_3276);
xor U8823 (N_8823,N_4947,N_4260);
nor U8824 (N_8824,N_4144,N_418);
and U8825 (N_8825,N_498,N_1988);
or U8826 (N_8826,N_3745,N_1119);
and U8827 (N_8827,N_2443,N_2028);
nor U8828 (N_8828,N_1144,N_1982);
and U8829 (N_8829,N_2091,N_3744);
and U8830 (N_8830,N_2948,N_3435);
nor U8831 (N_8831,N_2722,N_3011);
nor U8832 (N_8832,N_35,N_4017);
nand U8833 (N_8833,N_2396,N_3999);
xor U8834 (N_8834,N_3808,N_249);
and U8835 (N_8835,N_422,N_3032);
nand U8836 (N_8836,N_2612,N_2732);
nand U8837 (N_8837,N_2605,N_3519);
or U8838 (N_8838,N_3960,N_774);
or U8839 (N_8839,N_2870,N_3245);
xor U8840 (N_8840,N_4851,N_3976);
nor U8841 (N_8841,N_392,N_2454);
xnor U8842 (N_8842,N_1831,N_2129);
and U8843 (N_8843,N_4973,N_938);
and U8844 (N_8844,N_1302,N_2848);
xor U8845 (N_8845,N_1866,N_1477);
nand U8846 (N_8846,N_2528,N_2354);
or U8847 (N_8847,N_957,N_2712);
xnor U8848 (N_8848,N_2372,N_1944);
xnor U8849 (N_8849,N_4834,N_3895);
xor U8850 (N_8850,N_268,N_345);
and U8851 (N_8851,N_817,N_4678);
and U8852 (N_8852,N_4514,N_4719);
xor U8853 (N_8853,N_3312,N_2079);
and U8854 (N_8854,N_2652,N_3179);
or U8855 (N_8855,N_3480,N_4800);
nor U8856 (N_8856,N_1846,N_2434);
and U8857 (N_8857,N_2099,N_4936);
or U8858 (N_8858,N_2239,N_1844);
or U8859 (N_8859,N_1782,N_230);
nor U8860 (N_8860,N_2904,N_2078);
and U8861 (N_8861,N_2789,N_850);
xor U8862 (N_8862,N_4768,N_2590);
or U8863 (N_8863,N_4958,N_2787);
or U8864 (N_8864,N_1720,N_1754);
xor U8865 (N_8865,N_4872,N_447);
or U8866 (N_8866,N_2303,N_2154);
and U8867 (N_8867,N_3297,N_1222);
xor U8868 (N_8868,N_313,N_4918);
xor U8869 (N_8869,N_2913,N_1057);
and U8870 (N_8870,N_535,N_3430);
or U8871 (N_8871,N_2189,N_3798);
xnor U8872 (N_8872,N_845,N_73);
nor U8873 (N_8873,N_3137,N_4160);
nor U8874 (N_8874,N_4304,N_1782);
or U8875 (N_8875,N_1161,N_161);
xor U8876 (N_8876,N_4977,N_2816);
or U8877 (N_8877,N_1613,N_3611);
nand U8878 (N_8878,N_4178,N_4962);
or U8879 (N_8879,N_726,N_4903);
xor U8880 (N_8880,N_2962,N_319);
and U8881 (N_8881,N_2846,N_4442);
nor U8882 (N_8882,N_4536,N_1280);
nor U8883 (N_8883,N_3173,N_2865);
or U8884 (N_8884,N_2433,N_2615);
or U8885 (N_8885,N_4864,N_3198);
nand U8886 (N_8886,N_2036,N_1539);
nor U8887 (N_8887,N_217,N_1250);
nand U8888 (N_8888,N_997,N_3435);
nand U8889 (N_8889,N_959,N_2171);
nand U8890 (N_8890,N_791,N_454);
or U8891 (N_8891,N_2165,N_1017);
nor U8892 (N_8892,N_4347,N_3762);
and U8893 (N_8893,N_4689,N_4048);
or U8894 (N_8894,N_3599,N_886);
or U8895 (N_8895,N_925,N_1856);
nor U8896 (N_8896,N_4100,N_2209);
nor U8897 (N_8897,N_4273,N_3341);
or U8898 (N_8898,N_782,N_4669);
nor U8899 (N_8899,N_4691,N_845);
xor U8900 (N_8900,N_855,N_1606);
or U8901 (N_8901,N_4951,N_3668);
and U8902 (N_8902,N_982,N_4308);
nor U8903 (N_8903,N_3281,N_2437);
nor U8904 (N_8904,N_2997,N_4871);
xnor U8905 (N_8905,N_1430,N_124);
nor U8906 (N_8906,N_1483,N_4593);
xor U8907 (N_8907,N_246,N_2260);
and U8908 (N_8908,N_900,N_1656);
nor U8909 (N_8909,N_4988,N_2629);
nor U8910 (N_8910,N_3033,N_2372);
nand U8911 (N_8911,N_723,N_961);
and U8912 (N_8912,N_364,N_3201);
xor U8913 (N_8913,N_4618,N_4791);
nand U8914 (N_8914,N_4746,N_1816);
or U8915 (N_8915,N_1083,N_3890);
nor U8916 (N_8916,N_1819,N_3300);
nand U8917 (N_8917,N_588,N_2319);
nor U8918 (N_8918,N_426,N_3928);
nand U8919 (N_8919,N_4479,N_4373);
nand U8920 (N_8920,N_3505,N_4958);
and U8921 (N_8921,N_2130,N_2849);
or U8922 (N_8922,N_2956,N_4581);
and U8923 (N_8923,N_1182,N_2256);
and U8924 (N_8924,N_1626,N_4673);
nand U8925 (N_8925,N_4161,N_4417);
or U8926 (N_8926,N_2330,N_131);
nand U8927 (N_8927,N_226,N_4689);
and U8928 (N_8928,N_2396,N_4743);
and U8929 (N_8929,N_482,N_4074);
nand U8930 (N_8930,N_2270,N_2467);
and U8931 (N_8931,N_101,N_409);
nor U8932 (N_8932,N_2019,N_2754);
nand U8933 (N_8933,N_1218,N_574);
xnor U8934 (N_8934,N_500,N_4786);
and U8935 (N_8935,N_1993,N_1245);
nor U8936 (N_8936,N_1348,N_1267);
or U8937 (N_8937,N_1652,N_4033);
and U8938 (N_8938,N_4568,N_3301);
nand U8939 (N_8939,N_3160,N_4210);
nand U8940 (N_8940,N_2442,N_220);
and U8941 (N_8941,N_4973,N_1760);
nand U8942 (N_8942,N_3225,N_4198);
nor U8943 (N_8943,N_4056,N_1046);
or U8944 (N_8944,N_4143,N_4421);
nor U8945 (N_8945,N_3291,N_4688);
or U8946 (N_8946,N_2146,N_2976);
xor U8947 (N_8947,N_1285,N_1250);
nor U8948 (N_8948,N_1294,N_302);
nand U8949 (N_8949,N_1241,N_4476);
xnor U8950 (N_8950,N_1064,N_706);
nand U8951 (N_8951,N_1121,N_3468);
nor U8952 (N_8952,N_425,N_596);
nor U8953 (N_8953,N_952,N_660);
nor U8954 (N_8954,N_2929,N_1732);
and U8955 (N_8955,N_2662,N_2867);
or U8956 (N_8956,N_4158,N_3838);
and U8957 (N_8957,N_2975,N_4843);
nand U8958 (N_8958,N_1616,N_1881);
nand U8959 (N_8959,N_468,N_2905);
nand U8960 (N_8960,N_3406,N_4010);
nor U8961 (N_8961,N_911,N_707);
and U8962 (N_8962,N_4624,N_4379);
nor U8963 (N_8963,N_2585,N_2647);
and U8964 (N_8964,N_4804,N_1380);
xnor U8965 (N_8965,N_3761,N_1811);
or U8966 (N_8966,N_3160,N_1668);
nor U8967 (N_8967,N_3478,N_3992);
and U8968 (N_8968,N_4054,N_3594);
nand U8969 (N_8969,N_783,N_4509);
nor U8970 (N_8970,N_1178,N_1718);
and U8971 (N_8971,N_4307,N_1249);
nor U8972 (N_8972,N_2298,N_4955);
nor U8973 (N_8973,N_174,N_101);
or U8974 (N_8974,N_2751,N_846);
nand U8975 (N_8975,N_2585,N_631);
nor U8976 (N_8976,N_4893,N_3118);
nor U8977 (N_8977,N_2982,N_4312);
xor U8978 (N_8978,N_4187,N_1036);
nand U8979 (N_8979,N_4302,N_1739);
xnor U8980 (N_8980,N_4998,N_2403);
xnor U8981 (N_8981,N_2017,N_1287);
nor U8982 (N_8982,N_1808,N_1640);
or U8983 (N_8983,N_3311,N_4265);
xor U8984 (N_8984,N_2249,N_1416);
xnor U8985 (N_8985,N_2398,N_4981);
or U8986 (N_8986,N_225,N_406);
nor U8987 (N_8987,N_2849,N_4085);
xor U8988 (N_8988,N_664,N_2556);
and U8989 (N_8989,N_1449,N_2125);
xnor U8990 (N_8990,N_1041,N_640);
and U8991 (N_8991,N_338,N_3516);
and U8992 (N_8992,N_3009,N_226);
nand U8993 (N_8993,N_1578,N_2822);
or U8994 (N_8994,N_2655,N_1033);
nand U8995 (N_8995,N_1609,N_3136);
and U8996 (N_8996,N_2789,N_3923);
and U8997 (N_8997,N_4731,N_865);
nand U8998 (N_8998,N_3129,N_2393);
xor U8999 (N_8999,N_3141,N_1442);
xnor U9000 (N_9000,N_473,N_1915);
nand U9001 (N_9001,N_4755,N_1880);
nand U9002 (N_9002,N_1962,N_4873);
or U9003 (N_9003,N_1086,N_2271);
and U9004 (N_9004,N_2160,N_4021);
xor U9005 (N_9005,N_944,N_3674);
or U9006 (N_9006,N_2165,N_1952);
nor U9007 (N_9007,N_449,N_4322);
nand U9008 (N_9008,N_3342,N_3873);
or U9009 (N_9009,N_823,N_2754);
nand U9010 (N_9010,N_3761,N_4112);
and U9011 (N_9011,N_2957,N_4904);
nor U9012 (N_9012,N_1371,N_1154);
xnor U9013 (N_9013,N_720,N_1561);
nor U9014 (N_9014,N_158,N_155);
nor U9015 (N_9015,N_4762,N_4264);
nand U9016 (N_9016,N_3276,N_4697);
and U9017 (N_9017,N_4336,N_3932);
and U9018 (N_9018,N_1594,N_17);
nand U9019 (N_9019,N_2695,N_4373);
and U9020 (N_9020,N_3631,N_4313);
nor U9021 (N_9021,N_4413,N_3901);
or U9022 (N_9022,N_1874,N_3177);
or U9023 (N_9023,N_4678,N_4672);
nand U9024 (N_9024,N_3452,N_3674);
nand U9025 (N_9025,N_2703,N_486);
and U9026 (N_9026,N_594,N_129);
and U9027 (N_9027,N_4853,N_474);
or U9028 (N_9028,N_389,N_1568);
and U9029 (N_9029,N_1146,N_2912);
and U9030 (N_9030,N_870,N_4964);
and U9031 (N_9031,N_1487,N_3234);
or U9032 (N_9032,N_1390,N_1091);
xnor U9033 (N_9033,N_3598,N_4633);
nand U9034 (N_9034,N_4680,N_3983);
nor U9035 (N_9035,N_988,N_4641);
nand U9036 (N_9036,N_1702,N_1038);
xnor U9037 (N_9037,N_4083,N_4620);
xor U9038 (N_9038,N_447,N_3885);
and U9039 (N_9039,N_1765,N_3603);
or U9040 (N_9040,N_47,N_4287);
and U9041 (N_9041,N_3972,N_1052);
and U9042 (N_9042,N_745,N_674);
or U9043 (N_9043,N_3915,N_79);
and U9044 (N_9044,N_3397,N_1258);
nor U9045 (N_9045,N_1382,N_300);
or U9046 (N_9046,N_3410,N_99);
xor U9047 (N_9047,N_3640,N_4765);
and U9048 (N_9048,N_1868,N_4836);
and U9049 (N_9049,N_1993,N_4183);
xnor U9050 (N_9050,N_4833,N_4164);
or U9051 (N_9051,N_2871,N_1031);
and U9052 (N_9052,N_2234,N_374);
or U9053 (N_9053,N_2033,N_621);
and U9054 (N_9054,N_4262,N_4625);
or U9055 (N_9055,N_3266,N_1355);
and U9056 (N_9056,N_2909,N_2261);
nand U9057 (N_9057,N_643,N_1905);
and U9058 (N_9058,N_3093,N_2689);
and U9059 (N_9059,N_5,N_2623);
and U9060 (N_9060,N_3908,N_1873);
nor U9061 (N_9061,N_2467,N_2452);
xnor U9062 (N_9062,N_2620,N_542);
xnor U9063 (N_9063,N_2787,N_3073);
nand U9064 (N_9064,N_815,N_260);
and U9065 (N_9065,N_4720,N_3402);
nand U9066 (N_9066,N_498,N_4158);
or U9067 (N_9067,N_2594,N_3121);
and U9068 (N_9068,N_4922,N_1740);
and U9069 (N_9069,N_2840,N_3688);
nand U9070 (N_9070,N_3809,N_680);
or U9071 (N_9071,N_2943,N_463);
nor U9072 (N_9072,N_5,N_4088);
or U9073 (N_9073,N_3507,N_4390);
xor U9074 (N_9074,N_2455,N_3260);
nor U9075 (N_9075,N_1209,N_773);
and U9076 (N_9076,N_2452,N_4624);
nand U9077 (N_9077,N_698,N_1078);
nor U9078 (N_9078,N_2317,N_999);
or U9079 (N_9079,N_4497,N_2993);
and U9080 (N_9080,N_3241,N_4327);
nor U9081 (N_9081,N_3124,N_4099);
nor U9082 (N_9082,N_3732,N_3341);
nand U9083 (N_9083,N_3206,N_617);
xnor U9084 (N_9084,N_4473,N_3216);
nand U9085 (N_9085,N_2431,N_1870);
xnor U9086 (N_9086,N_3708,N_2505);
nor U9087 (N_9087,N_1143,N_4789);
nand U9088 (N_9088,N_3981,N_4196);
and U9089 (N_9089,N_422,N_341);
and U9090 (N_9090,N_1956,N_3513);
xnor U9091 (N_9091,N_1950,N_4350);
xor U9092 (N_9092,N_2067,N_684);
xor U9093 (N_9093,N_2295,N_1719);
or U9094 (N_9094,N_1748,N_1025);
xnor U9095 (N_9095,N_2780,N_1282);
nand U9096 (N_9096,N_1510,N_4721);
or U9097 (N_9097,N_3165,N_949);
and U9098 (N_9098,N_379,N_4327);
and U9099 (N_9099,N_3345,N_4572);
and U9100 (N_9100,N_4665,N_2093);
nand U9101 (N_9101,N_4498,N_965);
nor U9102 (N_9102,N_3490,N_2237);
nand U9103 (N_9103,N_4796,N_4165);
and U9104 (N_9104,N_620,N_70);
or U9105 (N_9105,N_508,N_2974);
nand U9106 (N_9106,N_3458,N_3029);
or U9107 (N_9107,N_757,N_3186);
nand U9108 (N_9108,N_2528,N_3131);
nor U9109 (N_9109,N_4120,N_3140);
and U9110 (N_9110,N_2020,N_4341);
xor U9111 (N_9111,N_3232,N_3462);
xor U9112 (N_9112,N_4959,N_4810);
nand U9113 (N_9113,N_3765,N_2828);
or U9114 (N_9114,N_1204,N_4311);
or U9115 (N_9115,N_2658,N_2256);
nor U9116 (N_9116,N_1426,N_924);
nor U9117 (N_9117,N_1902,N_2036);
xnor U9118 (N_9118,N_4608,N_2663);
and U9119 (N_9119,N_4203,N_1706);
or U9120 (N_9120,N_2271,N_1934);
nand U9121 (N_9121,N_3922,N_2407);
xor U9122 (N_9122,N_840,N_4174);
nor U9123 (N_9123,N_4035,N_4891);
xor U9124 (N_9124,N_2961,N_3955);
xnor U9125 (N_9125,N_1037,N_2716);
and U9126 (N_9126,N_2823,N_3220);
nor U9127 (N_9127,N_3206,N_1794);
xor U9128 (N_9128,N_4700,N_726);
xnor U9129 (N_9129,N_431,N_187);
xor U9130 (N_9130,N_3153,N_2775);
xnor U9131 (N_9131,N_352,N_2693);
and U9132 (N_9132,N_2589,N_4973);
nand U9133 (N_9133,N_4863,N_2923);
or U9134 (N_9134,N_4074,N_2275);
or U9135 (N_9135,N_3650,N_4359);
nand U9136 (N_9136,N_1041,N_452);
nor U9137 (N_9137,N_4464,N_4852);
xor U9138 (N_9138,N_1381,N_4446);
or U9139 (N_9139,N_313,N_3690);
xnor U9140 (N_9140,N_896,N_2462);
or U9141 (N_9141,N_4035,N_3724);
xnor U9142 (N_9142,N_4003,N_1055);
nand U9143 (N_9143,N_1428,N_3302);
xnor U9144 (N_9144,N_4136,N_2718);
nor U9145 (N_9145,N_4634,N_4877);
and U9146 (N_9146,N_495,N_1391);
nand U9147 (N_9147,N_1878,N_2618);
xnor U9148 (N_9148,N_1553,N_623);
and U9149 (N_9149,N_1788,N_4705);
and U9150 (N_9150,N_4711,N_2376);
nor U9151 (N_9151,N_2231,N_1463);
or U9152 (N_9152,N_3407,N_760);
or U9153 (N_9153,N_2939,N_101);
nand U9154 (N_9154,N_534,N_2273);
or U9155 (N_9155,N_1719,N_3944);
and U9156 (N_9156,N_349,N_3363);
and U9157 (N_9157,N_834,N_666);
xnor U9158 (N_9158,N_4561,N_2191);
or U9159 (N_9159,N_2954,N_3508);
and U9160 (N_9160,N_2601,N_1365);
xor U9161 (N_9161,N_4322,N_4430);
or U9162 (N_9162,N_835,N_3749);
xor U9163 (N_9163,N_2956,N_3792);
or U9164 (N_9164,N_1399,N_3593);
and U9165 (N_9165,N_539,N_593);
nor U9166 (N_9166,N_2347,N_530);
nand U9167 (N_9167,N_2902,N_3566);
and U9168 (N_9168,N_1696,N_3544);
xnor U9169 (N_9169,N_4217,N_851);
and U9170 (N_9170,N_3688,N_4282);
and U9171 (N_9171,N_4171,N_4871);
nand U9172 (N_9172,N_2283,N_2135);
and U9173 (N_9173,N_3184,N_1130);
or U9174 (N_9174,N_1142,N_2936);
nand U9175 (N_9175,N_470,N_916);
nand U9176 (N_9176,N_4101,N_212);
nand U9177 (N_9177,N_3971,N_2199);
nor U9178 (N_9178,N_4733,N_4042);
nand U9179 (N_9179,N_1094,N_2757);
nor U9180 (N_9180,N_1571,N_2838);
xor U9181 (N_9181,N_1223,N_985);
and U9182 (N_9182,N_1853,N_2049);
xnor U9183 (N_9183,N_147,N_1651);
nand U9184 (N_9184,N_4888,N_4921);
xor U9185 (N_9185,N_3895,N_3807);
xor U9186 (N_9186,N_4046,N_2416);
nand U9187 (N_9187,N_3453,N_1965);
or U9188 (N_9188,N_2098,N_762);
xnor U9189 (N_9189,N_3757,N_303);
and U9190 (N_9190,N_4579,N_1728);
nand U9191 (N_9191,N_2898,N_4375);
and U9192 (N_9192,N_455,N_2886);
xnor U9193 (N_9193,N_4654,N_1554);
xnor U9194 (N_9194,N_2450,N_2102);
nor U9195 (N_9195,N_3368,N_4818);
xnor U9196 (N_9196,N_726,N_3678);
nor U9197 (N_9197,N_2749,N_3995);
nor U9198 (N_9198,N_131,N_3672);
xor U9199 (N_9199,N_2504,N_4132);
xnor U9200 (N_9200,N_1876,N_1644);
and U9201 (N_9201,N_95,N_3791);
nor U9202 (N_9202,N_801,N_3394);
xor U9203 (N_9203,N_4576,N_450);
nand U9204 (N_9204,N_401,N_1625);
xor U9205 (N_9205,N_280,N_402);
or U9206 (N_9206,N_4019,N_4620);
nand U9207 (N_9207,N_2659,N_4864);
and U9208 (N_9208,N_4052,N_1778);
or U9209 (N_9209,N_1850,N_4750);
and U9210 (N_9210,N_4184,N_2696);
or U9211 (N_9211,N_2172,N_3796);
or U9212 (N_9212,N_938,N_4441);
xnor U9213 (N_9213,N_996,N_2023);
nand U9214 (N_9214,N_4665,N_1065);
and U9215 (N_9215,N_4359,N_2156);
and U9216 (N_9216,N_3319,N_855);
nor U9217 (N_9217,N_3894,N_3222);
nor U9218 (N_9218,N_3888,N_4263);
or U9219 (N_9219,N_691,N_1734);
or U9220 (N_9220,N_2930,N_3342);
or U9221 (N_9221,N_405,N_4543);
nand U9222 (N_9222,N_2160,N_2384);
nand U9223 (N_9223,N_778,N_1115);
nand U9224 (N_9224,N_3314,N_4430);
or U9225 (N_9225,N_1982,N_3877);
nor U9226 (N_9226,N_285,N_1145);
xnor U9227 (N_9227,N_4122,N_3856);
and U9228 (N_9228,N_3130,N_1749);
and U9229 (N_9229,N_1413,N_1003);
and U9230 (N_9230,N_3041,N_2267);
nand U9231 (N_9231,N_4386,N_3399);
and U9232 (N_9232,N_3209,N_4478);
xor U9233 (N_9233,N_129,N_4317);
xnor U9234 (N_9234,N_3182,N_2754);
nand U9235 (N_9235,N_3098,N_784);
nor U9236 (N_9236,N_3940,N_4396);
nand U9237 (N_9237,N_813,N_3540);
or U9238 (N_9238,N_3376,N_4410);
nand U9239 (N_9239,N_4785,N_2120);
xor U9240 (N_9240,N_3461,N_4594);
xnor U9241 (N_9241,N_376,N_1674);
nand U9242 (N_9242,N_2815,N_4963);
nor U9243 (N_9243,N_4010,N_1277);
nand U9244 (N_9244,N_2074,N_2976);
and U9245 (N_9245,N_3839,N_923);
xnor U9246 (N_9246,N_2337,N_2144);
xor U9247 (N_9247,N_458,N_537);
nor U9248 (N_9248,N_4005,N_791);
or U9249 (N_9249,N_2096,N_1151);
nand U9250 (N_9250,N_1363,N_3085);
xor U9251 (N_9251,N_2112,N_2132);
nand U9252 (N_9252,N_3420,N_3418);
nand U9253 (N_9253,N_1252,N_2837);
xor U9254 (N_9254,N_3125,N_985);
nor U9255 (N_9255,N_1432,N_3567);
xnor U9256 (N_9256,N_3690,N_2789);
or U9257 (N_9257,N_1955,N_3992);
xor U9258 (N_9258,N_3445,N_365);
or U9259 (N_9259,N_1825,N_2433);
xor U9260 (N_9260,N_2720,N_3725);
or U9261 (N_9261,N_1365,N_2812);
nand U9262 (N_9262,N_696,N_1136);
xnor U9263 (N_9263,N_2690,N_3139);
or U9264 (N_9264,N_3003,N_3048);
nor U9265 (N_9265,N_855,N_2736);
xnor U9266 (N_9266,N_4595,N_2196);
nand U9267 (N_9267,N_3081,N_4654);
nand U9268 (N_9268,N_1747,N_525);
or U9269 (N_9269,N_2462,N_1563);
nor U9270 (N_9270,N_436,N_873);
xor U9271 (N_9271,N_13,N_3944);
xnor U9272 (N_9272,N_404,N_1930);
and U9273 (N_9273,N_2976,N_2219);
nand U9274 (N_9274,N_3788,N_345);
nor U9275 (N_9275,N_3985,N_2861);
xor U9276 (N_9276,N_3277,N_2205);
nand U9277 (N_9277,N_4776,N_1194);
or U9278 (N_9278,N_4493,N_4950);
nand U9279 (N_9279,N_4090,N_3673);
or U9280 (N_9280,N_2040,N_3356);
nand U9281 (N_9281,N_2397,N_1695);
and U9282 (N_9282,N_3137,N_3000);
or U9283 (N_9283,N_3564,N_2160);
xnor U9284 (N_9284,N_2935,N_2580);
xor U9285 (N_9285,N_13,N_642);
xnor U9286 (N_9286,N_1357,N_1887);
nand U9287 (N_9287,N_755,N_4702);
nor U9288 (N_9288,N_1405,N_4206);
xnor U9289 (N_9289,N_1735,N_2260);
xor U9290 (N_9290,N_4946,N_3954);
nor U9291 (N_9291,N_3759,N_3489);
nand U9292 (N_9292,N_3090,N_947);
nand U9293 (N_9293,N_387,N_1041);
xnor U9294 (N_9294,N_3686,N_2304);
nor U9295 (N_9295,N_434,N_4482);
or U9296 (N_9296,N_4766,N_3787);
or U9297 (N_9297,N_2775,N_1548);
nand U9298 (N_9298,N_1203,N_3195);
nor U9299 (N_9299,N_2485,N_4162);
nor U9300 (N_9300,N_4669,N_2738);
and U9301 (N_9301,N_2369,N_3282);
and U9302 (N_9302,N_3781,N_4062);
xor U9303 (N_9303,N_2455,N_320);
xnor U9304 (N_9304,N_925,N_4655);
or U9305 (N_9305,N_4587,N_120);
nor U9306 (N_9306,N_3931,N_481);
xnor U9307 (N_9307,N_2550,N_2261);
or U9308 (N_9308,N_1196,N_2596);
and U9309 (N_9309,N_464,N_3679);
nor U9310 (N_9310,N_3349,N_814);
or U9311 (N_9311,N_4658,N_1830);
and U9312 (N_9312,N_4272,N_4997);
and U9313 (N_9313,N_2278,N_3619);
nand U9314 (N_9314,N_3682,N_2422);
and U9315 (N_9315,N_281,N_846);
and U9316 (N_9316,N_4482,N_4280);
nand U9317 (N_9317,N_3008,N_3864);
and U9318 (N_9318,N_2362,N_4468);
nor U9319 (N_9319,N_3601,N_9);
xor U9320 (N_9320,N_2127,N_1837);
and U9321 (N_9321,N_538,N_4573);
or U9322 (N_9322,N_1474,N_44);
nand U9323 (N_9323,N_4892,N_3517);
or U9324 (N_9324,N_716,N_3852);
or U9325 (N_9325,N_4454,N_1850);
nand U9326 (N_9326,N_4424,N_2250);
and U9327 (N_9327,N_4903,N_3174);
and U9328 (N_9328,N_2567,N_4805);
nand U9329 (N_9329,N_483,N_2520);
nor U9330 (N_9330,N_4484,N_1147);
xnor U9331 (N_9331,N_3996,N_1363);
nand U9332 (N_9332,N_185,N_2463);
xor U9333 (N_9333,N_13,N_1040);
nor U9334 (N_9334,N_3179,N_4641);
or U9335 (N_9335,N_2545,N_144);
or U9336 (N_9336,N_4671,N_1588);
xor U9337 (N_9337,N_152,N_1892);
nand U9338 (N_9338,N_4515,N_3388);
xnor U9339 (N_9339,N_3034,N_4166);
or U9340 (N_9340,N_4536,N_110);
xnor U9341 (N_9341,N_4084,N_3706);
nor U9342 (N_9342,N_1888,N_3030);
xnor U9343 (N_9343,N_1624,N_2918);
nor U9344 (N_9344,N_3260,N_4753);
nand U9345 (N_9345,N_1246,N_3833);
nand U9346 (N_9346,N_3695,N_2800);
nor U9347 (N_9347,N_734,N_336);
xnor U9348 (N_9348,N_2746,N_1272);
nor U9349 (N_9349,N_3306,N_829);
or U9350 (N_9350,N_4997,N_881);
and U9351 (N_9351,N_4423,N_687);
xnor U9352 (N_9352,N_4854,N_970);
and U9353 (N_9353,N_2043,N_36);
and U9354 (N_9354,N_3237,N_989);
or U9355 (N_9355,N_1063,N_2060);
nand U9356 (N_9356,N_3414,N_1712);
nor U9357 (N_9357,N_1902,N_411);
nor U9358 (N_9358,N_3056,N_2177);
xnor U9359 (N_9359,N_416,N_4209);
and U9360 (N_9360,N_3062,N_4267);
and U9361 (N_9361,N_2795,N_1583);
or U9362 (N_9362,N_746,N_3016);
and U9363 (N_9363,N_2511,N_847);
nand U9364 (N_9364,N_2247,N_1742);
or U9365 (N_9365,N_3127,N_2879);
xor U9366 (N_9366,N_1800,N_2088);
xor U9367 (N_9367,N_356,N_2440);
or U9368 (N_9368,N_2870,N_2776);
nand U9369 (N_9369,N_1703,N_2065);
nor U9370 (N_9370,N_783,N_1029);
nand U9371 (N_9371,N_4709,N_1728);
and U9372 (N_9372,N_183,N_3643);
and U9373 (N_9373,N_324,N_4844);
or U9374 (N_9374,N_3563,N_4537);
and U9375 (N_9375,N_824,N_1281);
nand U9376 (N_9376,N_598,N_4167);
nand U9377 (N_9377,N_4268,N_1248);
xnor U9378 (N_9378,N_2099,N_1387);
and U9379 (N_9379,N_4488,N_3750);
or U9380 (N_9380,N_203,N_3352);
nand U9381 (N_9381,N_1182,N_3039);
xnor U9382 (N_9382,N_732,N_3575);
nand U9383 (N_9383,N_470,N_2385);
nor U9384 (N_9384,N_1864,N_940);
or U9385 (N_9385,N_3399,N_1129);
xor U9386 (N_9386,N_1030,N_568);
xor U9387 (N_9387,N_590,N_2130);
or U9388 (N_9388,N_2300,N_68);
or U9389 (N_9389,N_3485,N_4333);
nor U9390 (N_9390,N_3726,N_3716);
xor U9391 (N_9391,N_586,N_4010);
xor U9392 (N_9392,N_4640,N_2832);
or U9393 (N_9393,N_3386,N_1662);
nand U9394 (N_9394,N_2488,N_2580);
and U9395 (N_9395,N_361,N_4540);
nand U9396 (N_9396,N_3676,N_3858);
or U9397 (N_9397,N_427,N_626);
and U9398 (N_9398,N_605,N_3790);
nand U9399 (N_9399,N_2257,N_225);
or U9400 (N_9400,N_4446,N_4117);
or U9401 (N_9401,N_3337,N_2518);
nand U9402 (N_9402,N_2413,N_2650);
nand U9403 (N_9403,N_508,N_3362);
nand U9404 (N_9404,N_3863,N_1452);
nor U9405 (N_9405,N_400,N_4706);
or U9406 (N_9406,N_166,N_1545);
or U9407 (N_9407,N_1502,N_1785);
nand U9408 (N_9408,N_2613,N_275);
nand U9409 (N_9409,N_2833,N_1064);
nor U9410 (N_9410,N_2306,N_4818);
nand U9411 (N_9411,N_2334,N_3650);
xor U9412 (N_9412,N_3026,N_138);
xor U9413 (N_9413,N_3478,N_348);
or U9414 (N_9414,N_1212,N_2277);
or U9415 (N_9415,N_538,N_3596);
nand U9416 (N_9416,N_1559,N_184);
nand U9417 (N_9417,N_1675,N_3875);
nand U9418 (N_9418,N_1415,N_2476);
or U9419 (N_9419,N_593,N_615);
or U9420 (N_9420,N_4010,N_2702);
nor U9421 (N_9421,N_3556,N_838);
and U9422 (N_9422,N_4090,N_80);
nor U9423 (N_9423,N_2014,N_1301);
xor U9424 (N_9424,N_1386,N_2949);
nor U9425 (N_9425,N_462,N_2368);
and U9426 (N_9426,N_2658,N_3420);
nand U9427 (N_9427,N_4108,N_4029);
or U9428 (N_9428,N_2076,N_4514);
nand U9429 (N_9429,N_2366,N_851);
nand U9430 (N_9430,N_3576,N_3720);
xnor U9431 (N_9431,N_3641,N_717);
xor U9432 (N_9432,N_3292,N_4650);
nor U9433 (N_9433,N_4956,N_2026);
and U9434 (N_9434,N_2975,N_3055);
xnor U9435 (N_9435,N_2789,N_707);
and U9436 (N_9436,N_3848,N_1757);
and U9437 (N_9437,N_3888,N_3355);
xnor U9438 (N_9438,N_3508,N_408);
or U9439 (N_9439,N_3545,N_2364);
or U9440 (N_9440,N_1466,N_4300);
or U9441 (N_9441,N_492,N_802);
nand U9442 (N_9442,N_1178,N_2066);
nand U9443 (N_9443,N_2275,N_2615);
and U9444 (N_9444,N_329,N_496);
nor U9445 (N_9445,N_1890,N_1286);
or U9446 (N_9446,N_4315,N_4927);
nand U9447 (N_9447,N_2823,N_771);
or U9448 (N_9448,N_2998,N_3030);
xor U9449 (N_9449,N_4297,N_3606);
xor U9450 (N_9450,N_945,N_4094);
and U9451 (N_9451,N_781,N_373);
and U9452 (N_9452,N_4509,N_757);
xor U9453 (N_9453,N_4445,N_4047);
or U9454 (N_9454,N_3071,N_1124);
nand U9455 (N_9455,N_4399,N_385);
nor U9456 (N_9456,N_4156,N_629);
nor U9457 (N_9457,N_1918,N_2211);
and U9458 (N_9458,N_1878,N_3137);
nor U9459 (N_9459,N_4975,N_362);
nand U9460 (N_9460,N_431,N_388);
or U9461 (N_9461,N_4955,N_3507);
nand U9462 (N_9462,N_4603,N_3175);
nand U9463 (N_9463,N_95,N_1043);
nand U9464 (N_9464,N_1660,N_4078);
nor U9465 (N_9465,N_676,N_1108);
and U9466 (N_9466,N_3557,N_750);
xnor U9467 (N_9467,N_2867,N_1756);
and U9468 (N_9468,N_3996,N_3387);
or U9469 (N_9469,N_2413,N_4894);
nor U9470 (N_9470,N_2292,N_1323);
and U9471 (N_9471,N_2140,N_33);
and U9472 (N_9472,N_880,N_3090);
nor U9473 (N_9473,N_4863,N_4374);
or U9474 (N_9474,N_2783,N_2504);
nand U9475 (N_9475,N_215,N_4866);
nor U9476 (N_9476,N_4213,N_2047);
nand U9477 (N_9477,N_4846,N_726);
xor U9478 (N_9478,N_3024,N_4713);
or U9479 (N_9479,N_2344,N_4143);
nand U9480 (N_9480,N_2957,N_3634);
or U9481 (N_9481,N_48,N_1219);
nand U9482 (N_9482,N_4265,N_1903);
and U9483 (N_9483,N_442,N_4071);
xor U9484 (N_9484,N_3460,N_580);
xor U9485 (N_9485,N_2532,N_3769);
xnor U9486 (N_9486,N_2514,N_3268);
nor U9487 (N_9487,N_2152,N_3268);
and U9488 (N_9488,N_3269,N_2857);
or U9489 (N_9489,N_2404,N_1242);
nor U9490 (N_9490,N_3894,N_1683);
nor U9491 (N_9491,N_114,N_3800);
and U9492 (N_9492,N_342,N_857);
and U9493 (N_9493,N_126,N_493);
or U9494 (N_9494,N_3654,N_3082);
xor U9495 (N_9495,N_752,N_4983);
or U9496 (N_9496,N_2503,N_2614);
nor U9497 (N_9497,N_1974,N_163);
xor U9498 (N_9498,N_692,N_209);
xor U9499 (N_9499,N_31,N_3603);
nand U9500 (N_9500,N_2863,N_1483);
and U9501 (N_9501,N_2138,N_2754);
or U9502 (N_9502,N_4926,N_3311);
xor U9503 (N_9503,N_4049,N_1613);
nor U9504 (N_9504,N_3313,N_119);
xnor U9505 (N_9505,N_257,N_4016);
and U9506 (N_9506,N_4390,N_4234);
nor U9507 (N_9507,N_177,N_485);
and U9508 (N_9508,N_1690,N_1402);
or U9509 (N_9509,N_789,N_3142);
and U9510 (N_9510,N_4720,N_3881);
and U9511 (N_9511,N_1228,N_2453);
xnor U9512 (N_9512,N_3477,N_3781);
nor U9513 (N_9513,N_336,N_394);
or U9514 (N_9514,N_981,N_2004);
xor U9515 (N_9515,N_4935,N_798);
xnor U9516 (N_9516,N_1180,N_4769);
or U9517 (N_9517,N_178,N_4210);
nand U9518 (N_9518,N_2801,N_2497);
nand U9519 (N_9519,N_3282,N_1359);
xor U9520 (N_9520,N_3435,N_1851);
or U9521 (N_9521,N_137,N_365);
nor U9522 (N_9522,N_1275,N_1621);
xor U9523 (N_9523,N_4153,N_88);
nand U9524 (N_9524,N_3119,N_841);
nand U9525 (N_9525,N_817,N_3374);
or U9526 (N_9526,N_4113,N_2749);
nor U9527 (N_9527,N_3841,N_625);
nor U9528 (N_9528,N_3523,N_1808);
or U9529 (N_9529,N_1110,N_539);
and U9530 (N_9530,N_752,N_2741);
xnor U9531 (N_9531,N_1909,N_1782);
and U9532 (N_9532,N_1479,N_3198);
and U9533 (N_9533,N_2768,N_4142);
xor U9534 (N_9534,N_1607,N_2135);
nand U9535 (N_9535,N_4016,N_3225);
and U9536 (N_9536,N_285,N_2761);
xor U9537 (N_9537,N_814,N_4198);
and U9538 (N_9538,N_2891,N_1274);
nand U9539 (N_9539,N_4531,N_4949);
nand U9540 (N_9540,N_3543,N_948);
nand U9541 (N_9541,N_1892,N_3752);
and U9542 (N_9542,N_1331,N_3347);
and U9543 (N_9543,N_3384,N_2632);
and U9544 (N_9544,N_3143,N_129);
or U9545 (N_9545,N_3585,N_2642);
and U9546 (N_9546,N_232,N_1034);
nor U9547 (N_9547,N_1805,N_20);
nor U9548 (N_9548,N_3742,N_4500);
nand U9549 (N_9549,N_777,N_3703);
and U9550 (N_9550,N_4032,N_4099);
or U9551 (N_9551,N_2261,N_2911);
xnor U9552 (N_9552,N_141,N_757);
or U9553 (N_9553,N_1162,N_3554);
or U9554 (N_9554,N_2657,N_1280);
or U9555 (N_9555,N_2032,N_383);
xor U9556 (N_9556,N_2119,N_1227);
nor U9557 (N_9557,N_2256,N_2903);
and U9558 (N_9558,N_2591,N_2630);
nand U9559 (N_9559,N_3153,N_4733);
nor U9560 (N_9560,N_142,N_3207);
xnor U9561 (N_9561,N_880,N_4489);
and U9562 (N_9562,N_2572,N_4984);
or U9563 (N_9563,N_4690,N_1142);
nor U9564 (N_9564,N_52,N_4791);
or U9565 (N_9565,N_2988,N_332);
and U9566 (N_9566,N_2730,N_2023);
and U9567 (N_9567,N_3060,N_2697);
or U9568 (N_9568,N_4314,N_1850);
nand U9569 (N_9569,N_3369,N_117);
or U9570 (N_9570,N_34,N_780);
nor U9571 (N_9571,N_1440,N_1759);
or U9572 (N_9572,N_381,N_2396);
or U9573 (N_9573,N_841,N_455);
nor U9574 (N_9574,N_4548,N_3267);
xnor U9575 (N_9575,N_1949,N_60);
and U9576 (N_9576,N_1853,N_3633);
and U9577 (N_9577,N_3898,N_266);
nand U9578 (N_9578,N_1809,N_2631);
xnor U9579 (N_9579,N_1057,N_4853);
xnor U9580 (N_9580,N_4523,N_2897);
xor U9581 (N_9581,N_3071,N_2473);
nor U9582 (N_9582,N_1457,N_1041);
xnor U9583 (N_9583,N_313,N_2349);
nor U9584 (N_9584,N_4749,N_4842);
or U9585 (N_9585,N_3363,N_1636);
xor U9586 (N_9586,N_3690,N_2173);
nand U9587 (N_9587,N_2547,N_58);
and U9588 (N_9588,N_1087,N_851);
or U9589 (N_9589,N_3235,N_4830);
and U9590 (N_9590,N_4655,N_2156);
and U9591 (N_9591,N_446,N_3859);
xor U9592 (N_9592,N_214,N_3661);
and U9593 (N_9593,N_1468,N_3264);
or U9594 (N_9594,N_2659,N_2350);
xnor U9595 (N_9595,N_4521,N_620);
nand U9596 (N_9596,N_527,N_2103);
and U9597 (N_9597,N_1875,N_4720);
or U9598 (N_9598,N_3468,N_3625);
nand U9599 (N_9599,N_1443,N_2604);
and U9600 (N_9600,N_3955,N_3917);
xor U9601 (N_9601,N_2738,N_1712);
or U9602 (N_9602,N_2135,N_2337);
and U9603 (N_9603,N_4002,N_4858);
and U9604 (N_9604,N_4450,N_806);
and U9605 (N_9605,N_1183,N_3089);
or U9606 (N_9606,N_1296,N_266);
xor U9607 (N_9607,N_1837,N_1998);
or U9608 (N_9608,N_4661,N_4444);
and U9609 (N_9609,N_3273,N_1119);
or U9610 (N_9610,N_4302,N_2184);
and U9611 (N_9611,N_2382,N_2256);
xor U9612 (N_9612,N_1459,N_4070);
xor U9613 (N_9613,N_3309,N_3079);
xnor U9614 (N_9614,N_4354,N_2795);
xnor U9615 (N_9615,N_3389,N_3459);
nand U9616 (N_9616,N_2532,N_2452);
xnor U9617 (N_9617,N_2751,N_4516);
xor U9618 (N_9618,N_661,N_1766);
nor U9619 (N_9619,N_376,N_2871);
and U9620 (N_9620,N_906,N_1786);
xor U9621 (N_9621,N_655,N_2858);
and U9622 (N_9622,N_3635,N_1337);
nor U9623 (N_9623,N_1014,N_4912);
xnor U9624 (N_9624,N_4933,N_3501);
and U9625 (N_9625,N_4472,N_4764);
and U9626 (N_9626,N_3577,N_1405);
xnor U9627 (N_9627,N_369,N_2503);
or U9628 (N_9628,N_1683,N_69);
and U9629 (N_9629,N_3490,N_942);
nand U9630 (N_9630,N_381,N_3311);
xor U9631 (N_9631,N_1419,N_3387);
or U9632 (N_9632,N_3553,N_4177);
nor U9633 (N_9633,N_59,N_540);
nand U9634 (N_9634,N_4263,N_121);
xor U9635 (N_9635,N_4667,N_3111);
nand U9636 (N_9636,N_3779,N_2846);
and U9637 (N_9637,N_2161,N_4285);
or U9638 (N_9638,N_2387,N_2840);
or U9639 (N_9639,N_4869,N_3505);
and U9640 (N_9640,N_495,N_3422);
xor U9641 (N_9641,N_2864,N_2954);
nor U9642 (N_9642,N_2148,N_4559);
and U9643 (N_9643,N_2940,N_2026);
nor U9644 (N_9644,N_902,N_1420);
xor U9645 (N_9645,N_3609,N_1484);
xor U9646 (N_9646,N_1800,N_972);
and U9647 (N_9647,N_560,N_3965);
nor U9648 (N_9648,N_4024,N_2531);
and U9649 (N_9649,N_426,N_4324);
xnor U9650 (N_9650,N_4616,N_2315);
nand U9651 (N_9651,N_2714,N_1511);
or U9652 (N_9652,N_625,N_1850);
and U9653 (N_9653,N_2898,N_2661);
and U9654 (N_9654,N_559,N_3238);
or U9655 (N_9655,N_88,N_2985);
and U9656 (N_9656,N_3453,N_4636);
and U9657 (N_9657,N_4316,N_3546);
nand U9658 (N_9658,N_1676,N_3026);
and U9659 (N_9659,N_1386,N_2650);
or U9660 (N_9660,N_3999,N_4230);
xor U9661 (N_9661,N_2974,N_62);
or U9662 (N_9662,N_2362,N_3869);
nor U9663 (N_9663,N_1080,N_3355);
nor U9664 (N_9664,N_1056,N_4537);
and U9665 (N_9665,N_2653,N_2726);
xor U9666 (N_9666,N_770,N_1429);
nand U9667 (N_9667,N_1824,N_3686);
nand U9668 (N_9668,N_2815,N_491);
nand U9669 (N_9669,N_2299,N_793);
or U9670 (N_9670,N_3930,N_2244);
nor U9671 (N_9671,N_2455,N_2584);
nand U9672 (N_9672,N_4809,N_1921);
and U9673 (N_9673,N_4143,N_3037);
or U9674 (N_9674,N_2534,N_3021);
xnor U9675 (N_9675,N_3757,N_4923);
or U9676 (N_9676,N_820,N_1683);
nor U9677 (N_9677,N_205,N_2739);
xor U9678 (N_9678,N_66,N_2872);
xor U9679 (N_9679,N_2646,N_1863);
or U9680 (N_9680,N_1016,N_1507);
nor U9681 (N_9681,N_1354,N_4005);
nor U9682 (N_9682,N_4075,N_4848);
and U9683 (N_9683,N_3620,N_903);
xnor U9684 (N_9684,N_335,N_607);
and U9685 (N_9685,N_933,N_108);
xor U9686 (N_9686,N_2703,N_2956);
or U9687 (N_9687,N_1451,N_3061);
nor U9688 (N_9688,N_3019,N_1483);
xor U9689 (N_9689,N_2224,N_1936);
and U9690 (N_9690,N_3133,N_3289);
nor U9691 (N_9691,N_931,N_2692);
and U9692 (N_9692,N_4766,N_2841);
xor U9693 (N_9693,N_742,N_1522);
xor U9694 (N_9694,N_522,N_2117);
nor U9695 (N_9695,N_1934,N_198);
or U9696 (N_9696,N_3849,N_1526);
nor U9697 (N_9697,N_1253,N_870);
xor U9698 (N_9698,N_3464,N_2148);
xnor U9699 (N_9699,N_2189,N_3059);
xor U9700 (N_9700,N_684,N_1824);
nand U9701 (N_9701,N_804,N_4716);
nand U9702 (N_9702,N_4813,N_1296);
and U9703 (N_9703,N_4482,N_228);
and U9704 (N_9704,N_4776,N_3575);
nand U9705 (N_9705,N_2681,N_451);
nor U9706 (N_9706,N_1079,N_3150);
xnor U9707 (N_9707,N_1062,N_707);
and U9708 (N_9708,N_1973,N_2674);
and U9709 (N_9709,N_3619,N_1216);
nor U9710 (N_9710,N_4306,N_884);
xnor U9711 (N_9711,N_3710,N_2392);
xnor U9712 (N_9712,N_739,N_4705);
nand U9713 (N_9713,N_155,N_1232);
and U9714 (N_9714,N_764,N_3015);
and U9715 (N_9715,N_4862,N_4766);
xnor U9716 (N_9716,N_1410,N_4629);
and U9717 (N_9717,N_3280,N_4067);
or U9718 (N_9718,N_2618,N_3862);
nand U9719 (N_9719,N_1257,N_4257);
xnor U9720 (N_9720,N_3473,N_1928);
or U9721 (N_9721,N_2172,N_3150);
nand U9722 (N_9722,N_1925,N_3373);
and U9723 (N_9723,N_2588,N_377);
and U9724 (N_9724,N_4852,N_3200);
nor U9725 (N_9725,N_839,N_3323);
xnor U9726 (N_9726,N_749,N_2794);
and U9727 (N_9727,N_1124,N_3436);
or U9728 (N_9728,N_2014,N_4654);
xor U9729 (N_9729,N_2807,N_19);
or U9730 (N_9730,N_3857,N_239);
nand U9731 (N_9731,N_1088,N_3811);
nand U9732 (N_9732,N_1312,N_3817);
nand U9733 (N_9733,N_1058,N_3153);
nand U9734 (N_9734,N_144,N_3445);
nor U9735 (N_9735,N_16,N_1298);
nand U9736 (N_9736,N_4956,N_2541);
xnor U9737 (N_9737,N_1077,N_940);
nor U9738 (N_9738,N_461,N_3669);
or U9739 (N_9739,N_1405,N_2734);
or U9740 (N_9740,N_4375,N_768);
nor U9741 (N_9741,N_4231,N_4359);
and U9742 (N_9742,N_4366,N_4132);
and U9743 (N_9743,N_4304,N_3280);
nor U9744 (N_9744,N_2036,N_2527);
xor U9745 (N_9745,N_3256,N_3509);
nor U9746 (N_9746,N_3515,N_3169);
or U9747 (N_9747,N_4279,N_1741);
xor U9748 (N_9748,N_3178,N_466);
nand U9749 (N_9749,N_1931,N_1661);
xor U9750 (N_9750,N_2936,N_1676);
nand U9751 (N_9751,N_4057,N_4852);
xnor U9752 (N_9752,N_340,N_3080);
nor U9753 (N_9753,N_1751,N_3335);
and U9754 (N_9754,N_3391,N_3255);
and U9755 (N_9755,N_1726,N_4546);
or U9756 (N_9756,N_3794,N_3664);
nor U9757 (N_9757,N_4065,N_1307);
nand U9758 (N_9758,N_45,N_3849);
and U9759 (N_9759,N_4846,N_4427);
xnor U9760 (N_9760,N_1430,N_264);
or U9761 (N_9761,N_1584,N_2397);
or U9762 (N_9762,N_4607,N_3334);
xor U9763 (N_9763,N_1098,N_2759);
xnor U9764 (N_9764,N_814,N_4240);
xor U9765 (N_9765,N_21,N_4614);
xor U9766 (N_9766,N_3011,N_1103);
xor U9767 (N_9767,N_1216,N_3299);
or U9768 (N_9768,N_1531,N_3081);
or U9769 (N_9769,N_2533,N_1544);
nand U9770 (N_9770,N_2977,N_4622);
nor U9771 (N_9771,N_2523,N_4513);
xor U9772 (N_9772,N_3754,N_644);
xor U9773 (N_9773,N_1626,N_4781);
or U9774 (N_9774,N_1465,N_1248);
xor U9775 (N_9775,N_3511,N_3600);
nor U9776 (N_9776,N_1947,N_3566);
or U9777 (N_9777,N_2562,N_570);
nand U9778 (N_9778,N_3208,N_968);
nor U9779 (N_9779,N_2069,N_2911);
nor U9780 (N_9780,N_1259,N_3603);
and U9781 (N_9781,N_2967,N_689);
or U9782 (N_9782,N_1465,N_647);
nor U9783 (N_9783,N_798,N_3967);
nor U9784 (N_9784,N_2012,N_1663);
nand U9785 (N_9785,N_1642,N_684);
xor U9786 (N_9786,N_4007,N_461);
xnor U9787 (N_9787,N_1783,N_1153);
or U9788 (N_9788,N_801,N_3321);
xnor U9789 (N_9789,N_3778,N_3569);
nand U9790 (N_9790,N_1533,N_4083);
and U9791 (N_9791,N_499,N_4345);
and U9792 (N_9792,N_692,N_3389);
nor U9793 (N_9793,N_3124,N_2984);
or U9794 (N_9794,N_2025,N_2495);
or U9795 (N_9795,N_1670,N_1021);
and U9796 (N_9796,N_3753,N_1190);
xor U9797 (N_9797,N_21,N_4572);
xor U9798 (N_9798,N_2581,N_103);
xnor U9799 (N_9799,N_800,N_625);
xnor U9800 (N_9800,N_3263,N_2141);
nor U9801 (N_9801,N_2001,N_1609);
or U9802 (N_9802,N_1434,N_2290);
xor U9803 (N_9803,N_2530,N_2856);
and U9804 (N_9804,N_4618,N_1634);
or U9805 (N_9805,N_4419,N_4045);
xor U9806 (N_9806,N_225,N_2754);
nand U9807 (N_9807,N_3512,N_1161);
nor U9808 (N_9808,N_3275,N_1689);
and U9809 (N_9809,N_63,N_2731);
or U9810 (N_9810,N_1834,N_1932);
nor U9811 (N_9811,N_949,N_3247);
nor U9812 (N_9812,N_3749,N_2758);
or U9813 (N_9813,N_3542,N_1110);
nor U9814 (N_9814,N_4370,N_3375);
xor U9815 (N_9815,N_1264,N_4957);
or U9816 (N_9816,N_1857,N_3836);
xnor U9817 (N_9817,N_1155,N_4734);
and U9818 (N_9818,N_2664,N_4407);
or U9819 (N_9819,N_2095,N_2002);
nand U9820 (N_9820,N_1897,N_1482);
and U9821 (N_9821,N_3184,N_336);
and U9822 (N_9822,N_748,N_838);
nor U9823 (N_9823,N_221,N_2895);
nand U9824 (N_9824,N_3857,N_4015);
nor U9825 (N_9825,N_2797,N_2531);
and U9826 (N_9826,N_1473,N_1532);
or U9827 (N_9827,N_2955,N_770);
and U9828 (N_9828,N_317,N_24);
xor U9829 (N_9829,N_782,N_3247);
nand U9830 (N_9830,N_4217,N_554);
nand U9831 (N_9831,N_78,N_3518);
xor U9832 (N_9832,N_3584,N_2934);
and U9833 (N_9833,N_2335,N_3764);
and U9834 (N_9834,N_73,N_4454);
nor U9835 (N_9835,N_2198,N_4116);
nand U9836 (N_9836,N_4103,N_2713);
and U9837 (N_9837,N_142,N_728);
nor U9838 (N_9838,N_776,N_3208);
and U9839 (N_9839,N_2096,N_4779);
or U9840 (N_9840,N_243,N_264);
xnor U9841 (N_9841,N_861,N_1333);
or U9842 (N_9842,N_753,N_2283);
xnor U9843 (N_9843,N_2296,N_359);
and U9844 (N_9844,N_1126,N_4887);
nand U9845 (N_9845,N_645,N_2007);
nor U9846 (N_9846,N_1803,N_4423);
or U9847 (N_9847,N_1103,N_4923);
nor U9848 (N_9848,N_3727,N_4478);
and U9849 (N_9849,N_3534,N_2005);
or U9850 (N_9850,N_3432,N_4718);
nor U9851 (N_9851,N_4152,N_3899);
nand U9852 (N_9852,N_1122,N_676);
nand U9853 (N_9853,N_2902,N_609);
and U9854 (N_9854,N_962,N_2047);
and U9855 (N_9855,N_3620,N_182);
xor U9856 (N_9856,N_4221,N_1537);
or U9857 (N_9857,N_3795,N_4907);
nand U9858 (N_9858,N_3273,N_4202);
nand U9859 (N_9859,N_2891,N_3362);
and U9860 (N_9860,N_4978,N_1124);
nor U9861 (N_9861,N_1909,N_3379);
xor U9862 (N_9862,N_4627,N_158);
or U9863 (N_9863,N_4913,N_1176);
and U9864 (N_9864,N_2955,N_4748);
nor U9865 (N_9865,N_1797,N_3520);
or U9866 (N_9866,N_1941,N_1811);
or U9867 (N_9867,N_476,N_1249);
nor U9868 (N_9868,N_885,N_169);
xor U9869 (N_9869,N_3069,N_1382);
and U9870 (N_9870,N_3861,N_3006);
and U9871 (N_9871,N_4757,N_4536);
or U9872 (N_9872,N_4225,N_4299);
xor U9873 (N_9873,N_4750,N_2396);
nor U9874 (N_9874,N_3358,N_2754);
nand U9875 (N_9875,N_4473,N_2681);
nand U9876 (N_9876,N_4757,N_3623);
nand U9877 (N_9877,N_3652,N_4217);
nor U9878 (N_9878,N_4655,N_707);
and U9879 (N_9879,N_3114,N_2203);
and U9880 (N_9880,N_1276,N_2057);
and U9881 (N_9881,N_1649,N_4653);
or U9882 (N_9882,N_3489,N_705);
xnor U9883 (N_9883,N_2499,N_2261);
nand U9884 (N_9884,N_1704,N_541);
xnor U9885 (N_9885,N_1746,N_220);
xnor U9886 (N_9886,N_1801,N_2359);
xnor U9887 (N_9887,N_4138,N_2250);
or U9888 (N_9888,N_1369,N_1907);
xor U9889 (N_9889,N_3685,N_692);
nand U9890 (N_9890,N_1029,N_1132);
xnor U9891 (N_9891,N_1160,N_3946);
nand U9892 (N_9892,N_3224,N_3272);
xnor U9893 (N_9893,N_4692,N_4408);
xor U9894 (N_9894,N_358,N_15);
xor U9895 (N_9895,N_917,N_4200);
or U9896 (N_9896,N_2612,N_238);
or U9897 (N_9897,N_2885,N_552);
nor U9898 (N_9898,N_893,N_1489);
and U9899 (N_9899,N_4616,N_4776);
and U9900 (N_9900,N_1373,N_239);
xor U9901 (N_9901,N_361,N_2059);
and U9902 (N_9902,N_522,N_1176);
nand U9903 (N_9903,N_4458,N_1513);
or U9904 (N_9904,N_4491,N_4010);
xor U9905 (N_9905,N_3640,N_4609);
or U9906 (N_9906,N_129,N_3616);
xor U9907 (N_9907,N_9,N_1381);
nand U9908 (N_9908,N_62,N_4002);
or U9909 (N_9909,N_4257,N_726);
and U9910 (N_9910,N_3100,N_2373);
nand U9911 (N_9911,N_4175,N_37);
xnor U9912 (N_9912,N_1166,N_3574);
and U9913 (N_9913,N_444,N_3307);
nor U9914 (N_9914,N_88,N_626);
xnor U9915 (N_9915,N_85,N_530);
or U9916 (N_9916,N_2948,N_2846);
and U9917 (N_9917,N_4969,N_1668);
nor U9918 (N_9918,N_3626,N_3602);
and U9919 (N_9919,N_3441,N_4322);
xor U9920 (N_9920,N_3405,N_792);
xnor U9921 (N_9921,N_801,N_1533);
or U9922 (N_9922,N_4242,N_3154);
and U9923 (N_9923,N_3037,N_2708);
nor U9924 (N_9924,N_3744,N_1709);
and U9925 (N_9925,N_3349,N_1788);
nand U9926 (N_9926,N_3675,N_4075);
nand U9927 (N_9927,N_4203,N_282);
xnor U9928 (N_9928,N_4275,N_2778);
xnor U9929 (N_9929,N_4590,N_4531);
nand U9930 (N_9930,N_4700,N_4444);
xor U9931 (N_9931,N_2762,N_2362);
nand U9932 (N_9932,N_4177,N_1781);
nand U9933 (N_9933,N_70,N_542);
nand U9934 (N_9934,N_358,N_2800);
nand U9935 (N_9935,N_2534,N_654);
nand U9936 (N_9936,N_1852,N_1578);
xor U9937 (N_9937,N_4230,N_1325);
xnor U9938 (N_9938,N_1636,N_962);
nand U9939 (N_9939,N_2412,N_4939);
nor U9940 (N_9940,N_3846,N_4684);
and U9941 (N_9941,N_396,N_230);
xnor U9942 (N_9942,N_4219,N_3024);
xnor U9943 (N_9943,N_2935,N_3650);
and U9944 (N_9944,N_4517,N_4281);
or U9945 (N_9945,N_4478,N_3332);
nor U9946 (N_9946,N_4735,N_1201);
nor U9947 (N_9947,N_3778,N_1149);
and U9948 (N_9948,N_292,N_4384);
or U9949 (N_9949,N_4031,N_2945);
xor U9950 (N_9950,N_1116,N_2492);
or U9951 (N_9951,N_4171,N_761);
or U9952 (N_9952,N_4783,N_129);
nor U9953 (N_9953,N_3557,N_2262);
nor U9954 (N_9954,N_1946,N_858);
or U9955 (N_9955,N_4789,N_2067);
nand U9956 (N_9956,N_2651,N_939);
xnor U9957 (N_9957,N_1919,N_1624);
nand U9958 (N_9958,N_3971,N_3907);
and U9959 (N_9959,N_4172,N_3050);
nor U9960 (N_9960,N_1376,N_2327);
nor U9961 (N_9961,N_649,N_4711);
xor U9962 (N_9962,N_1588,N_82);
or U9963 (N_9963,N_3935,N_1302);
nand U9964 (N_9964,N_1002,N_2764);
or U9965 (N_9965,N_2237,N_1801);
nand U9966 (N_9966,N_3529,N_4044);
and U9967 (N_9967,N_1040,N_4648);
nand U9968 (N_9968,N_3298,N_2012);
or U9969 (N_9969,N_3372,N_1067);
nand U9970 (N_9970,N_231,N_4777);
nand U9971 (N_9971,N_4610,N_2296);
and U9972 (N_9972,N_2347,N_287);
or U9973 (N_9973,N_3704,N_3277);
xnor U9974 (N_9974,N_2981,N_150);
xor U9975 (N_9975,N_2600,N_257);
nand U9976 (N_9976,N_3749,N_2679);
xor U9977 (N_9977,N_4459,N_4666);
or U9978 (N_9978,N_3962,N_2049);
and U9979 (N_9979,N_4879,N_71);
nand U9980 (N_9980,N_4507,N_1818);
nor U9981 (N_9981,N_2068,N_3145);
xor U9982 (N_9982,N_316,N_2842);
nor U9983 (N_9983,N_846,N_2630);
and U9984 (N_9984,N_3714,N_3394);
or U9985 (N_9985,N_3027,N_1660);
or U9986 (N_9986,N_2238,N_1647);
or U9987 (N_9987,N_1913,N_2092);
nor U9988 (N_9988,N_3123,N_1372);
nand U9989 (N_9989,N_561,N_1664);
and U9990 (N_9990,N_741,N_3488);
nor U9991 (N_9991,N_4762,N_4874);
nor U9992 (N_9992,N_3654,N_3114);
xnor U9993 (N_9993,N_1682,N_4825);
nand U9994 (N_9994,N_123,N_1993);
nor U9995 (N_9995,N_241,N_3862);
nor U9996 (N_9996,N_3492,N_3132);
and U9997 (N_9997,N_387,N_2438);
or U9998 (N_9998,N_1544,N_581);
nand U9999 (N_9999,N_2514,N_2654);
and U10000 (N_10000,N_9140,N_5244);
xnor U10001 (N_10001,N_7325,N_7700);
xnor U10002 (N_10002,N_5104,N_9774);
nand U10003 (N_10003,N_9717,N_9341);
and U10004 (N_10004,N_9370,N_8498);
and U10005 (N_10005,N_7677,N_5179);
nor U10006 (N_10006,N_5435,N_6639);
nand U10007 (N_10007,N_9889,N_8805);
and U10008 (N_10008,N_7217,N_9356);
and U10009 (N_10009,N_7293,N_9649);
nand U10010 (N_10010,N_5547,N_6300);
or U10011 (N_10011,N_6720,N_8535);
and U10012 (N_10012,N_7762,N_5243);
xnor U10013 (N_10013,N_5726,N_5503);
nand U10014 (N_10014,N_8036,N_8879);
nor U10015 (N_10015,N_8105,N_6058);
and U10016 (N_10016,N_9667,N_9837);
nor U10017 (N_10017,N_8560,N_5755);
nand U10018 (N_10018,N_7574,N_9778);
nor U10019 (N_10019,N_6550,N_5568);
nand U10020 (N_10020,N_7551,N_8334);
nand U10021 (N_10021,N_8602,N_6282);
nand U10022 (N_10022,N_7246,N_6296);
and U10023 (N_10023,N_5810,N_8723);
xor U10024 (N_10024,N_7037,N_9284);
nor U10025 (N_10025,N_8218,N_7532);
nand U10026 (N_10026,N_9292,N_9611);
xnor U10027 (N_10027,N_7719,N_9076);
and U10028 (N_10028,N_5937,N_8040);
nor U10029 (N_10029,N_5446,N_9217);
xor U10030 (N_10030,N_9849,N_7054);
nor U10031 (N_10031,N_8320,N_8383);
nor U10032 (N_10032,N_5680,N_8719);
nand U10033 (N_10033,N_9555,N_8623);
or U10034 (N_10034,N_9218,N_8944);
nand U10035 (N_10035,N_5079,N_7711);
xnor U10036 (N_10036,N_6878,N_6760);
or U10037 (N_10037,N_9927,N_6496);
xnor U10038 (N_10038,N_6194,N_9050);
and U10039 (N_10039,N_5606,N_5721);
xor U10040 (N_10040,N_7896,N_9124);
nand U10041 (N_10041,N_5310,N_6561);
xnor U10042 (N_10042,N_7140,N_7233);
xnor U10043 (N_10043,N_8314,N_9808);
nand U10044 (N_10044,N_5252,N_5672);
and U10045 (N_10045,N_8143,N_5671);
and U10046 (N_10046,N_5954,N_9977);
nand U10047 (N_10047,N_6601,N_6684);
xor U10048 (N_10048,N_6184,N_5231);
or U10049 (N_10049,N_5015,N_8999);
or U10050 (N_10050,N_9576,N_5081);
nor U10051 (N_10051,N_5058,N_6543);
nor U10052 (N_10052,N_9883,N_5363);
or U10053 (N_10053,N_5515,N_8791);
or U10054 (N_10054,N_6341,N_5922);
nand U10055 (N_10055,N_5343,N_6822);
nand U10056 (N_10056,N_9418,N_7210);
xnor U10057 (N_10057,N_7484,N_9701);
or U10058 (N_10058,N_5913,N_9027);
xnor U10059 (N_10059,N_7148,N_5450);
and U10060 (N_10060,N_6798,N_9036);
xnor U10061 (N_10061,N_6059,N_8172);
and U10062 (N_10062,N_9473,N_6213);
xnor U10063 (N_10063,N_6144,N_9268);
nand U10064 (N_10064,N_8123,N_7174);
nand U10065 (N_10065,N_9968,N_8896);
and U10066 (N_10066,N_9622,N_6612);
xor U10067 (N_10067,N_5313,N_7726);
and U10068 (N_10068,N_5185,N_7330);
nand U10069 (N_10069,N_6066,N_6412);
and U10070 (N_10070,N_5200,N_9914);
nand U10071 (N_10071,N_6558,N_5351);
and U10072 (N_10072,N_8043,N_6273);
xnor U10073 (N_10073,N_7682,N_9035);
and U10074 (N_10074,N_7007,N_5425);
or U10075 (N_10075,N_6071,N_5305);
xor U10076 (N_10076,N_9643,N_5824);
xor U10077 (N_10077,N_8090,N_9945);
and U10078 (N_10078,N_7195,N_9197);
xnor U10079 (N_10079,N_9413,N_5308);
and U10080 (N_10080,N_7722,N_8850);
nor U10081 (N_10081,N_7687,N_6335);
nand U10082 (N_10082,N_7613,N_5155);
nor U10083 (N_10083,N_8539,N_6329);
and U10084 (N_10084,N_7640,N_8661);
nand U10085 (N_10085,N_6706,N_6969);
and U10086 (N_10086,N_9167,N_9624);
nor U10087 (N_10087,N_7855,N_5137);
or U10088 (N_10088,N_9790,N_5384);
and U10089 (N_10089,N_5697,N_6976);
and U10090 (N_10090,N_9032,N_7566);
or U10091 (N_10091,N_7845,N_5784);
xnor U10092 (N_10092,N_8670,N_8596);
nor U10093 (N_10093,N_5072,N_9346);
xnor U10094 (N_10094,N_8772,N_8900);
or U10095 (N_10095,N_7492,N_5283);
and U10096 (N_10096,N_8159,N_5530);
or U10097 (N_10097,N_9738,N_7983);
or U10098 (N_10098,N_5742,N_7692);
or U10099 (N_10099,N_5345,N_8754);
xor U10100 (N_10100,N_6418,N_5447);
xnor U10101 (N_10101,N_8681,N_8308);
or U10102 (N_10102,N_9533,N_8426);
and U10103 (N_10103,N_9182,N_6010);
or U10104 (N_10104,N_5952,N_5579);
nor U10105 (N_10105,N_5796,N_9496);
and U10106 (N_10106,N_5717,N_6046);
nand U10107 (N_10107,N_6032,N_8996);
xnor U10108 (N_10108,N_9761,N_7130);
or U10109 (N_10109,N_6247,N_5999);
nand U10110 (N_10110,N_7906,N_7922);
xnor U10111 (N_10111,N_6348,N_9144);
nand U10112 (N_10112,N_9491,N_6655);
nor U10113 (N_10113,N_7443,N_5986);
and U10114 (N_10114,N_7810,N_7841);
xnor U10115 (N_10115,N_8825,N_5273);
nand U10116 (N_10116,N_9386,N_6591);
and U10117 (N_10117,N_7609,N_7717);
nand U10118 (N_10118,N_5086,N_8787);
and U10119 (N_10119,N_9985,N_7177);
nor U10120 (N_10120,N_6987,N_7043);
xor U10121 (N_10121,N_6697,N_6669);
and U10122 (N_10122,N_6468,N_6605);
nor U10123 (N_10123,N_5330,N_5929);
or U10124 (N_10124,N_8213,N_5379);
and U10125 (N_10125,N_5370,N_6693);
or U10126 (N_10126,N_7286,N_5059);
xor U10127 (N_10127,N_8046,N_9823);
nor U10128 (N_10128,N_6417,N_9949);
xnor U10129 (N_10129,N_5840,N_8522);
nand U10130 (N_10130,N_9507,N_5764);
nor U10131 (N_10131,N_5553,N_7314);
or U10132 (N_10132,N_6364,N_6179);
or U10133 (N_10133,N_6648,N_7990);
and U10134 (N_10134,N_5967,N_8229);
and U10135 (N_10135,N_7065,N_6527);
or U10136 (N_10136,N_7310,N_6872);
nand U10137 (N_10137,N_9753,N_6033);
nand U10138 (N_10138,N_7989,N_5092);
nor U10139 (N_10139,N_6708,N_9007);
nor U10140 (N_10140,N_9759,N_5766);
or U10141 (N_10141,N_6952,N_6338);
xor U10142 (N_10142,N_9591,N_7049);
or U10143 (N_10143,N_5266,N_8193);
and U10144 (N_10144,N_5600,N_5293);
nor U10145 (N_10145,N_5117,N_9002);
xnor U10146 (N_10146,N_7051,N_7159);
xnor U10147 (N_10147,N_7373,N_9063);
or U10148 (N_10148,N_6299,N_8385);
or U10149 (N_10149,N_8017,N_5780);
nand U10150 (N_10150,N_7555,N_9150);
nand U10151 (N_10151,N_7880,N_9899);
nand U10152 (N_10152,N_5382,N_8400);
nor U10153 (N_10153,N_8110,N_9443);
nor U10154 (N_10154,N_7781,N_6890);
nor U10155 (N_10155,N_8547,N_9869);
xor U10156 (N_10156,N_7721,N_5501);
nand U10157 (N_10157,N_6419,N_5955);
nor U10158 (N_10158,N_7926,N_5067);
and U10159 (N_10159,N_7077,N_6420);
and U10160 (N_10160,N_8666,N_8746);
or U10161 (N_10161,N_7006,N_8037);
xnor U10162 (N_10162,N_6228,N_5626);
xnor U10163 (N_10163,N_5202,N_9805);
nand U10164 (N_10164,N_6112,N_9669);
xor U10165 (N_10165,N_8161,N_5258);
xor U10166 (N_10166,N_8093,N_7501);
nor U10167 (N_10167,N_6559,N_6676);
nor U10168 (N_10168,N_8868,N_6089);
nand U10169 (N_10169,N_9239,N_5846);
nor U10170 (N_10170,N_7885,N_8472);
nor U10171 (N_10171,N_5208,N_8116);
and U10172 (N_10172,N_9707,N_5710);
nand U10173 (N_10173,N_7339,N_7671);
xnor U10174 (N_10174,N_9569,N_6451);
or U10175 (N_10175,N_5031,N_6493);
or U10176 (N_10176,N_5168,N_7596);
or U10177 (N_10177,N_6238,N_6689);
xor U10178 (N_10178,N_5436,N_6305);
nand U10179 (N_10179,N_8339,N_5933);
xnor U10180 (N_10180,N_7081,N_8827);
nand U10181 (N_10181,N_9506,N_9594);
nor U10182 (N_10182,N_9402,N_5335);
and U10183 (N_10183,N_6776,N_6941);
nand U10184 (N_10184,N_9721,N_6195);
nand U10185 (N_10185,N_7122,N_9118);
nor U10186 (N_10186,N_5131,N_9361);
xnor U10187 (N_10187,N_8653,N_8733);
or U10188 (N_10188,N_9605,N_5281);
and U10189 (N_10189,N_9991,N_6544);
xor U10190 (N_10190,N_7748,N_6777);
or U10191 (N_10191,N_7564,N_6534);
and U10192 (N_10192,N_9562,N_9152);
xnor U10193 (N_10193,N_8290,N_7331);
or U10194 (N_10194,N_5508,N_9151);
xnor U10195 (N_10195,N_6389,N_5704);
nand U10196 (N_10196,N_9842,N_5254);
and U10197 (N_10197,N_7289,N_7123);
or U10198 (N_10198,N_8469,N_8075);
nor U10199 (N_10199,N_6778,N_5338);
nor U10200 (N_10200,N_7674,N_6026);
xor U10201 (N_10201,N_9368,N_9585);
xnor U10202 (N_10202,N_5355,N_8209);
nand U10203 (N_10203,N_7363,N_6846);
nand U10204 (N_10204,N_8373,N_9091);
nor U10205 (N_10205,N_5950,N_7543);
or U10206 (N_10206,N_9971,N_7228);
or U10207 (N_10207,N_7418,N_9828);
or U10208 (N_10208,N_8346,N_8702);
nor U10209 (N_10209,N_5132,N_5905);
nand U10210 (N_10210,N_8651,N_6506);
and U10211 (N_10211,N_7452,N_9427);
and U10212 (N_10212,N_9107,N_9254);
nand U10213 (N_10213,N_5235,N_6276);
xor U10214 (N_10214,N_6542,N_6198);
nand U10215 (N_10215,N_8758,N_6710);
xor U10216 (N_10216,N_7147,N_5918);
nor U10217 (N_10217,N_8050,N_7980);
or U10218 (N_10218,N_9094,N_5904);
and U10219 (N_10219,N_6260,N_6268);
nand U10220 (N_10220,N_7761,N_8318);
or U10221 (N_10221,N_6652,N_8398);
and U10222 (N_10222,N_7535,N_6408);
or U10223 (N_10223,N_8028,N_9532);
or U10224 (N_10224,N_5242,N_6790);
and U10225 (N_10225,N_5720,N_6239);
and U10226 (N_10226,N_5312,N_7815);
or U10227 (N_10227,N_8080,N_9604);
nor U10228 (N_10228,N_9924,N_5669);
nand U10229 (N_10229,N_8327,N_8674);
and U10230 (N_10230,N_7798,N_8949);
nor U10231 (N_10231,N_8904,N_8935);
or U10232 (N_10232,N_8298,N_6472);
or U10233 (N_10233,N_5674,N_9044);
xnor U10234 (N_10234,N_6568,N_9796);
and U10235 (N_10235,N_5653,N_7992);
nand U10236 (N_10236,N_5945,N_9983);
or U10237 (N_10237,N_5139,N_5045);
and U10238 (N_10238,N_5576,N_7852);
and U10239 (N_10239,N_9069,N_7486);
xnor U10240 (N_10240,N_7627,N_7539);
nor U10241 (N_10241,N_7426,N_9235);
or U10242 (N_10242,N_5125,N_6193);
nor U10243 (N_10243,N_8158,N_9674);
or U10244 (N_10244,N_7457,N_8676);
xnor U10245 (N_10245,N_7215,N_7356);
xor U10246 (N_10246,N_9189,N_7480);
or U10247 (N_10247,N_9620,N_7662);
and U10248 (N_10248,N_7981,N_8911);
nor U10249 (N_10249,N_8087,N_7139);
nor U10250 (N_10250,N_9952,N_6812);
or U10251 (N_10251,N_6843,N_7739);
nand U10252 (N_10252,N_5221,N_7197);
or U10253 (N_10253,N_9918,N_7872);
or U10254 (N_10254,N_7207,N_9619);
nand U10255 (N_10255,N_7519,N_9739);
nor U10256 (N_10256,N_7379,N_8088);
nand U10257 (N_10257,N_6853,N_6093);
or U10258 (N_10258,N_6003,N_9166);
nand U10259 (N_10259,N_9158,N_9033);
xnor U10260 (N_10260,N_8541,N_7828);
and U10261 (N_10261,N_6111,N_6234);
or U10262 (N_10262,N_5691,N_6682);
nor U10263 (N_10263,N_9087,N_7375);
or U10264 (N_10264,N_6683,N_5364);
nand U10265 (N_10265,N_5633,N_8204);
nand U10266 (N_10266,N_6448,N_6369);
nand U10267 (N_10267,N_9464,N_7227);
nor U10268 (N_10268,N_5619,N_5218);
nor U10269 (N_10269,N_5286,N_5033);
xnor U10270 (N_10270,N_7685,N_8291);
nand U10271 (N_10271,N_5227,N_8014);
nand U10272 (N_10272,N_8362,N_9508);
xor U10273 (N_10273,N_9040,N_7984);
nor U10274 (N_10274,N_7715,N_9610);
nor U10275 (N_10275,N_9621,N_8288);
xor U10276 (N_10276,N_5407,N_6021);
nor U10277 (N_10277,N_5692,N_9375);
xor U10278 (N_10278,N_5687,N_6883);
xnor U10279 (N_10279,N_9019,N_8214);
nor U10280 (N_10280,N_7237,N_7038);
xor U10281 (N_10281,N_5361,N_7534);
or U10282 (N_10282,N_7076,N_5152);
and U10283 (N_10283,N_8439,N_6154);
or U10284 (N_10284,N_8713,N_5206);
nor U10285 (N_10285,N_9929,N_6699);
nor U10286 (N_10286,N_6162,N_7902);
nor U10287 (N_10287,N_8920,N_6113);
or U10288 (N_10288,N_8937,N_6881);
or U10289 (N_10289,N_8113,N_9729);
and U10290 (N_10290,N_9200,N_9559);
xnor U10291 (N_10291,N_6063,N_7580);
and U10292 (N_10292,N_7658,N_7202);
nor U10293 (N_10293,N_7821,N_7239);
and U10294 (N_10294,N_5620,N_6159);
xor U10295 (N_10295,N_8260,N_6197);
and U10296 (N_10296,N_8358,N_6083);
or U10297 (N_10297,N_7069,N_7308);
nand U10298 (N_10298,N_8106,N_5426);
nor U10299 (N_10299,N_8610,N_8870);
or U10300 (N_10300,N_6042,N_9744);
and U10301 (N_10301,N_6965,N_7728);
nor U10302 (N_10302,N_6114,N_9793);
nor U10303 (N_10303,N_9066,N_7449);
xor U10304 (N_10304,N_6874,N_6138);
or U10305 (N_10305,N_7268,N_5142);
and U10306 (N_10306,N_5270,N_8003);
or U10307 (N_10307,N_9811,N_6929);
or U10308 (N_10308,N_5781,N_6907);
xnor U10309 (N_10309,N_5114,N_7583);
nand U10310 (N_10310,N_8634,N_6469);
xnor U10311 (N_10311,N_6914,N_5932);
or U10312 (N_10312,N_6330,N_6137);
nand U10313 (N_10313,N_6986,N_5972);
nand U10314 (N_10314,N_7929,N_7313);
nand U10315 (N_10315,N_5782,N_8203);
nor U10316 (N_10316,N_8978,N_6370);
xnor U10317 (N_10317,N_5554,N_8828);
xor U10318 (N_10318,N_8155,N_7988);
nand U10319 (N_10319,N_8202,N_5850);
or U10320 (N_10320,N_8379,N_5275);
xnor U10321 (N_10321,N_8961,N_5462);
nor U10322 (N_10322,N_6366,N_9908);
and U10323 (N_10323,N_7579,N_9279);
nand U10324 (N_10324,N_6600,N_8264);
or U10325 (N_10325,N_7940,N_8943);
xor U10326 (N_10326,N_6319,N_8683);
nand U10327 (N_10327,N_8923,N_9468);
and U10328 (N_10328,N_5538,N_6110);
nand U10329 (N_10329,N_6386,N_7327);
and U10330 (N_10330,N_6920,N_9110);
xor U10331 (N_10331,N_7141,N_7342);
nand U10332 (N_10332,N_8335,N_6255);
xor U10333 (N_10333,N_9926,N_8410);
nor U10334 (N_10334,N_8729,N_6022);
xnor U10335 (N_10335,N_8420,N_8391);
nor U10336 (N_10336,N_7707,N_8559);
or U10337 (N_10337,N_8607,N_9972);
xor U10338 (N_10338,N_7219,N_5920);
or U10339 (N_10339,N_9981,N_9592);
nor U10340 (N_10340,N_9111,N_9075);
nand U10341 (N_10341,N_5891,N_5673);
xnor U10342 (N_10342,N_9462,N_7150);
nand U10343 (N_10343,N_6813,N_5853);
xor U10344 (N_10344,N_5344,N_6779);
or U10345 (N_10345,N_7320,N_7364);
or U10346 (N_10346,N_9130,N_5414);
or U10347 (N_10347,N_6148,N_8514);
xnor U10348 (N_10348,N_7475,N_8639);
and U10349 (N_10349,N_7332,N_9873);
and U10350 (N_10350,N_6579,N_7655);
or U10351 (N_10351,N_6025,N_7478);
xnor U10352 (N_10352,N_8876,N_8459);
xnor U10353 (N_10353,N_5613,N_7878);
xor U10354 (N_10354,N_5614,N_8842);
and U10355 (N_10355,N_6806,N_9851);
nand U10356 (N_10356,N_7011,N_7424);
and U10357 (N_10357,N_9997,N_8914);
nand U10358 (N_10358,N_6819,N_8768);
or U10359 (N_10359,N_6035,N_7820);
or U10360 (N_10360,N_8412,N_9113);
nor U10361 (N_10361,N_9333,N_6272);
nand U10362 (N_10362,N_8760,N_8219);
and U10363 (N_10363,N_5480,N_7198);
and U10364 (N_10364,N_5951,N_7436);
nand U10365 (N_10365,N_5875,N_6796);
and U10366 (N_10366,N_6845,N_5439);
nand U10367 (N_10367,N_9905,N_8771);
xor U10368 (N_10368,N_5819,N_6313);
nor U10369 (N_10369,N_9871,N_9568);
xor U10370 (N_10370,N_5468,N_8767);
or U10371 (N_10371,N_5839,N_7680);
and U10372 (N_10372,N_8424,N_5042);
nand U10373 (N_10373,N_7455,N_8886);
and U10374 (N_10374,N_8047,N_6804);
or U10375 (N_10375,N_7255,N_9574);
xnor U10376 (N_10376,N_6721,N_6916);
and U10377 (N_10377,N_5109,N_9098);
nand U10378 (N_10378,N_9727,N_5616);
nor U10379 (N_10379,N_7216,N_6808);
and U10380 (N_10380,N_5993,N_7001);
nand U10381 (N_10381,N_6133,N_6264);
or U10382 (N_10382,N_6507,N_7132);
nand U10383 (N_10383,N_7511,N_6135);
nand U10384 (N_10384,N_5184,N_6342);
xor U10385 (N_10385,N_7252,N_5842);
nor U10386 (N_10386,N_8257,N_9999);
nand U10387 (N_10387,N_9834,N_5337);
nand U10388 (N_10388,N_9628,N_6118);
or U10389 (N_10389,N_8130,N_7098);
nand U10390 (N_10390,N_8009,N_5274);
xnor U10391 (N_10391,N_7686,N_9434);
and U10392 (N_10392,N_7072,N_9688);
nand U10393 (N_10393,N_7738,N_9515);
xor U10394 (N_10394,N_6663,N_8192);
nor U10395 (N_10395,N_6908,N_8153);
or U10396 (N_10396,N_7577,N_7846);
and U10397 (N_10397,N_6438,N_9982);
and U10398 (N_10398,N_5946,N_7502);
nand U10399 (N_10399,N_6337,N_8108);
nor U10400 (N_10400,N_6487,N_5838);
nor U10401 (N_10401,N_9765,N_9121);
or U10402 (N_10402,N_9271,N_7747);
nor U10403 (N_10403,N_9665,N_5588);
xor U10404 (N_10404,N_5910,N_5165);
xnor U10405 (N_10405,N_7059,N_6423);
nor U10406 (N_10406,N_6831,N_5474);
nand U10407 (N_10407,N_6623,N_7256);
xnor U10408 (N_10408,N_6485,N_9081);
and U10409 (N_10409,N_6678,N_5814);
nand U10410 (N_10410,N_5097,N_5392);
and U10411 (N_10411,N_6927,N_9852);
nand U10412 (N_10412,N_6424,N_6641);
nor U10413 (N_10413,N_6219,N_7595);
xnor U10414 (N_10414,N_7930,N_5238);
or U10415 (N_10415,N_5422,N_7319);
nand U10416 (N_10416,N_6943,N_6352);
xor U10417 (N_10417,N_9504,N_5065);
nor U10418 (N_10418,N_9369,N_9973);
and U10419 (N_10419,N_6728,N_6607);
or U10420 (N_10420,N_9954,N_7023);
or U10421 (N_10421,N_6156,N_6246);
nor U10422 (N_10422,N_8671,N_6414);
nand U10423 (N_10423,N_5297,N_5349);
and U10424 (N_10424,N_7553,N_9021);
xor U10425 (N_10425,N_7193,N_6374);
or U10426 (N_10426,N_5592,N_9786);
nand U10427 (N_10427,N_6894,N_9332);
and U10428 (N_10428,N_9781,N_7889);
or U10429 (N_10429,N_9513,N_9678);
xor U10430 (N_10430,N_9691,N_7050);
or U10431 (N_10431,N_8934,N_7542);
nand U10432 (N_10432,N_5973,N_6763);
xnor U10433 (N_10433,N_7209,N_8727);
nor U10434 (N_10434,N_7611,N_8215);
nor U10435 (N_10435,N_8965,N_9273);
and U10436 (N_10436,N_5759,N_9303);
nand U10437 (N_10437,N_6099,N_9560);
nor U10438 (N_10438,N_8603,N_9455);
and U10439 (N_10439,N_8715,N_7030);
nand U10440 (N_10440,N_8809,N_5844);
and U10441 (N_10441,N_9409,N_5374);
or U10442 (N_10442,N_9011,N_7961);
xnor U10443 (N_10443,N_6501,N_9960);
xnor U10444 (N_10444,N_5415,N_8109);
xor U10445 (N_10445,N_7768,N_6407);
or U10446 (N_10446,N_9399,N_8121);
and U10447 (N_10447,N_6000,N_6539);
or U10448 (N_10448,N_5860,N_9536);
xnor U10449 (N_10449,N_7340,N_7755);
xor U10450 (N_10450,N_5226,N_7575);
and U10451 (N_10451,N_6869,N_8798);
xor U10452 (N_10452,N_5404,N_9380);
and U10453 (N_10453,N_8761,N_9718);
or U10454 (N_10454,N_9047,N_7103);
nand U10455 (N_10455,N_8018,N_6257);
or U10456 (N_10456,N_7782,N_8399);
nor U10457 (N_10457,N_5959,N_5602);
nor U10458 (N_10458,N_5713,N_8856);
xnor U10459 (N_10459,N_5173,N_8826);
nand U10460 (N_10460,N_7318,N_6750);
nand U10461 (N_10461,N_9055,N_8170);
and U10462 (N_10462,N_9459,N_7537);
nand U10463 (N_10463,N_7143,N_9447);
nand U10464 (N_10464,N_8840,N_7751);
nor U10465 (N_10465,N_8354,N_8992);
nor U10466 (N_10466,N_6218,N_6082);
nor U10467 (N_10467,N_7413,N_7649);
nand U10468 (N_10468,N_9350,N_6158);
xor U10469 (N_10469,N_8749,N_8578);
or U10470 (N_10470,N_5004,N_8632);
and U10471 (N_10471,N_9116,N_7249);
xnor U10472 (N_10472,N_8079,N_5490);
and U10473 (N_10473,N_9408,N_6049);
xnor U10474 (N_10474,N_6754,N_8259);
or U10475 (N_10475,N_5189,N_9294);
nand U10476 (N_10476,N_9431,N_5285);
or U10477 (N_10477,N_6857,N_8951);
nor U10478 (N_10478,N_6209,N_8571);
xor U10479 (N_10479,N_8368,N_6540);
nor U10480 (N_10480,N_5751,N_9785);
and U10481 (N_10481,N_8872,N_6404);
nor U10482 (N_10482,N_8630,N_7860);
nor U10483 (N_10483,N_9485,N_8356);
nor U10484 (N_10484,N_7718,N_6453);
xnor U10485 (N_10485,N_6513,N_9256);
and U10486 (N_10486,N_6731,N_5385);
xnor U10487 (N_10487,N_5528,N_5787);
and U10488 (N_10488,N_6698,N_8077);
and U10489 (N_10489,N_6562,N_8680);
nor U10490 (N_10490,N_9607,N_8044);
or U10491 (N_10491,N_5980,N_9192);
nor U10492 (N_10492,N_8757,N_9710);
and U10493 (N_10493,N_9245,N_5212);
nor U10494 (N_10494,N_7934,N_6304);
or U10495 (N_10495,N_6422,N_5460);
xor U10496 (N_10496,N_5837,N_7593);
and U10497 (N_10497,N_6211,N_6288);
and U10498 (N_10498,N_9843,N_5400);
and U10499 (N_10499,N_9797,N_8190);
or U10500 (N_10500,N_7172,N_5129);
and U10501 (N_10501,N_8223,N_5365);
nor U10502 (N_10502,N_8654,N_6031);
nor U10503 (N_10503,N_6512,N_9043);
nand U10504 (N_10504,N_6541,N_6517);
or U10505 (N_10505,N_5712,N_8917);
xor U10506 (N_10506,N_8664,N_7073);
nor U10507 (N_10507,N_7294,N_8021);
nand U10508 (N_10508,N_8059,N_8705);
or U10509 (N_10509,N_5979,N_9195);
nor U10510 (N_10510,N_7476,N_9948);
nand U10511 (N_10511,N_6859,N_8307);
nor U10512 (N_10512,N_7315,N_8744);
nor U10513 (N_10513,N_6130,N_5166);
nand U10514 (N_10514,N_6855,N_8407);
xnor U10515 (N_10515,N_6797,N_9037);
or U10516 (N_10516,N_6477,N_7759);
or U10517 (N_10517,N_5484,N_9696);
and U10518 (N_10518,N_9474,N_8660);
nand U10519 (N_10519,N_6709,N_7411);
or U10520 (N_10520,N_7624,N_9330);
nand U10521 (N_10521,N_9086,N_6510);
xor U10522 (N_10522,N_7033,N_8126);
or U10523 (N_10523,N_9731,N_7530);
and U10524 (N_10524,N_8102,N_7213);
or U10525 (N_10525,N_9514,N_6473);
or U10526 (N_10526,N_9147,N_7185);
nor U10527 (N_10527,N_6884,N_5334);
nor U10528 (N_10528,N_5482,N_5995);
nand U10529 (N_10529,N_6931,N_8704);
nand U10530 (N_10530,N_9656,N_8641);
nor U10531 (N_10531,N_9358,N_6972);
and U10532 (N_10532,N_6749,N_5569);
and U10533 (N_10533,N_8445,N_5123);
nor U10534 (N_10534,N_6688,N_6410);
nand U10535 (N_10535,N_7279,N_5873);
or U10536 (N_10536,N_7716,N_7941);
nor U10537 (N_10537,N_6454,N_8765);
xnor U10538 (N_10538,N_6018,N_8444);
and U10539 (N_10539,N_5373,N_5047);
nor U10540 (N_10540,N_5359,N_7620);
nor U10541 (N_10541,N_8145,N_7301);
nand U10542 (N_10542,N_5336,N_8751);
nand U10543 (N_10543,N_8952,N_9961);
and U10544 (N_10544,N_8716,N_5790);
or U10545 (N_10545,N_8330,N_6899);
or U10546 (N_10546,N_7376,N_5229);
nor U10547 (N_10547,N_9417,N_5603);
or U10548 (N_10548,N_6322,N_9735);
xor U10549 (N_10549,N_5635,N_9694);
and U10550 (N_10550,N_6619,N_9290);
nor U10551 (N_10551,N_6200,N_6391);
xnor U10552 (N_10552,N_5369,N_5188);
xor U10553 (N_10553,N_8898,N_8277);
and U10554 (N_10554,N_8374,N_5828);
and U10555 (N_10555,N_5282,N_9482);
nand U10556 (N_10556,N_8406,N_7380);
nand U10557 (N_10557,N_6462,N_7154);
and U10558 (N_10558,N_8313,N_6556);
and U10559 (N_10559,N_9220,N_8555);
nand U10560 (N_10560,N_9039,N_5427);
nand U10561 (N_10561,N_8703,N_5170);
and U10562 (N_10562,N_7538,N_7312);
or U10563 (N_10563,N_5325,N_6898);
or U10564 (N_10564,N_5121,N_9411);
nor U10565 (N_10565,N_7055,N_7608);
nor U10566 (N_10566,N_8169,N_9787);
nand U10567 (N_10567,N_6552,N_6172);
and U10568 (N_10568,N_6910,N_7993);
nand U10569 (N_10569,N_8493,N_9699);
nor U10570 (N_10570,N_7731,N_5140);
nor U10571 (N_10571,N_7190,N_7879);
or U10572 (N_10572,N_5022,N_5307);
and U10573 (N_10573,N_8084,N_7456);
and U10574 (N_10574,N_5505,N_7094);
and U10575 (N_10575,N_7244,N_9481);
nand U10576 (N_10576,N_6079,N_7295);
or U10577 (N_10577,N_8901,N_6719);
nand U10578 (N_10578,N_7546,N_5239);
xnor U10579 (N_10579,N_5423,N_5763);
nand U10580 (N_10580,N_6834,N_5329);
nand U10581 (N_10581,N_7181,N_7157);
and U10582 (N_10582,N_7222,N_6889);
and U10583 (N_10583,N_9329,N_7839);
and U10584 (N_10584,N_7901,N_6954);
or U10585 (N_10585,N_9572,N_7625);
nor U10586 (N_10586,N_8986,N_8333);
and U10587 (N_10587,N_8636,N_8199);
xnor U10588 (N_10588,N_6962,N_8332);
nor U10589 (N_10589,N_7212,N_9861);
and U10590 (N_10590,N_5269,N_6767);
and U10591 (N_10591,N_8415,N_5339);
nand U10592 (N_10592,N_5948,N_9917);
nor U10593 (N_10593,N_8769,N_5417);
or U10594 (N_10594,N_8178,N_7998);
nand U10595 (N_10595,N_8554,N_6178);
or U10596 (N_10596,N_9545,N_5476);
and U10597 (N_10597,N_5883,N_9794);
and U10598 (N_10598,N_5906,N_6223);
xor U10599 (N_10599,N_9149,N_8913);
or U10600 (N_10600,N_8450,N_9813);
nor U10601 (N_10601,N_9030,N_7515);
nor U10602 (N_10602,N_9275,N_7155);
xnor U10603 (N_10603,N_7699,N_6640);
xor U10604 (N_10604,N_6087,N_9114);
xor U10605 (N_10605,N_6181,N_6755);
or U10606 (N_10606,N_6494,N_9704);
nand U10607 (N_10607,N_7734,N_8243);
nand U10608 (N_10608,N_6180,N_9008);
nor U10609 (N_10609,N_8942,N_9103);
nor U10610 (N_10610,N_7243,N_8567);
xnor U10611 (N_10611,N_5657,N_8743);
nand U10612 (N_10612,N_6516,N_5309);
nand U10613 (N_10613,N_7034,N_6939);
xor U10614 (N_10614,N_7186,N_7652);
and U10615 (N_10615,N_9955,N_8501);
or U10616 (N_10616,N_5529,N_5797);
xor U10617 (N_10617,N_7266,N_8883);
xor U10618 (N_10618,N_7736,N_9631);
and U10619 (N_10619,N_9307,N_5138);
or U10620 (N_10620,N_8388,N_9698);
nor U10621 (N_10621,N_8885,N_5362);
nor U10622 (N_10622,N_5144,N_6631);
or U10623 (N_10623,N_5675,N_5527);
nor U10624 (N_10624,N_9426,N_9864);
or U10625 (N_10625,N_6405,N_7936);
or U10626 (N_10626,N_8564,N_5639);
and U10627 (N_10627,N_8546,N_6944);
xnor U10628 (N_10628,N_6717,N_9071);
and U10629 (N_10629,N_5861,N_6932);
xnor U10630 (N_10630,N_7638,N_6897);
nand U10631 (N_10631,N_7277,N_9858);
xor U10632 (N_10632,N_5960,N_6862);
or U10633 (N_10633,N_9203,N_8480);
or U10634 (N_10634,N_6281,N_5605);
or U10635 (N_10635,N_9551,N_5074);
nor U10636 (N_10636,N_6634,N_8588);
and U10637 (N_10637,N_8100,N_8119);
nor U10638 (N_10638,N_8361,N_9684);
xnor U10639 (N_10639,N_9742,N_9895);
nand U10640 (N_10640,N_6788,N_6549);
nor U10641 (N_10641,N_7021,N_8366);
nand U10642 (N_10642,N_6732,N_8927);
nand U10643 (N_10643,N_6323,N_7387);
xnor U10644 (N_10644,N_6729,N_6701);
nor U10645 (N_10645,N_8177,N_5798);
nand U10646 (N_10646,N_8538,N_5536);
nand U10647 (N_10647,N_7900,N_8941);
nor U10648 (N_10648,N_5191,N_6252);
and U10649 (N_10649,N_9109,N_6436);
and U10650 (N_10650,N_9975,N_8403);
nand U10651 (N_10651,N_7806,N_7965);
nor U10652 (N_10652,N_5424,N_9172);
xnor U10653 (N_10653,N_7124,N_5509);
and U10654 (N_10654,N_5767,N_8637);
and U10655 (N_10655,N_5690,N_9073);
nand U10656 (N_10656,N_8494,N_9053);
xnor U10657 (N_10657,N_7158,N_6563);
xor U10658 (N_10658,N_9237,N_6102);
xor U10659 (N_10659,N_5570,N_5851);
xnor U10660 (N_10660,N_7651,N_6661);
nand U10661 (N_10661,N_9106,N_9831);
xnor U10662 (N_10662,N_5898,N_5214);
nand U10663 (N_10663,N_9176,N_9424);
and U10664 (N_10664,N_6886,N_7703);
and U10665 (N_10665,N_8506,N_9963);
nand U10666 (N_10666,N_7758,N_6217);
or U10667 (N_10667,N_7985,N_8505);
nor U10668 (N_10668,N_6011,N_9088);
or U10669 (N_10669,N_9856,N_5066);
and U10670 (N_10670,N_9383,N_9221);
or U10671 (N_10671,N_6891,N_9486);
xor U10672 (N_10672,N_7881,N_6362);
and U10673 (N_10673,N_7614,N_8718);
and U10674 (N_10674,N_8150,N_7180);
or U10675 (N_10675,N_6587,N_6350);
xnor U10676 (N_10676,N_8766,N_7560);
nor U10677 (N_10677,N_8797,N_5778);
and U10678 (N_10678,N_7785,N_6278);
nand U10679 (N_10679,N_5150,N_8249);
or U10680 (N_10680,N_9493,N_5560);
nor U10681 (N_10681,N_6360,N_5161);
xor U10682 (N_10682,N_8070,N_9223);
nand U10683 (N_10683,N_7271,N_6240);
and U10684 (N_10684,N_9163,N_7442);
xnor U10685 (N_10685,N_8222,N_6290);
xor U10686 (N_10686,N_7105,N_8305);
and U10687 (N_10687,N_6249,N_7788);
xnor U10688 (N_10688,N_5183,N_7962);
xor U10689 (N_10689,N_5575,N_8271);
and U10690 (N_10690,N_9844,N_5013);
xnor U10691 (N_10691,N_9538,N_7152);
nor U10692 (N_10692,N_5511,N_6491);
xor U10693 (N_10693,N_7783,N_8245);
or U10694 (N_10694,N_7078,N_5630);
and U10695 (N_10695,N_8053,N_9228);
nand U10696 (N_10696,N_5655,N_7462);
xor U10697 (N_10697,N_5085,N_8551);
nand U10698 (N_10698,N_5924,N_7628);
nand U10699 (N_10699,N_5256,N_8936);
nand U10700 (N_10700,N_7948,N_8974);
nand U10701 (N_10701,N_5643,N_5459);
or U10702 (N_10702,N_5652,N_9138);
or U10703 (N_10703,N_5938,N_9250);
nand U10704 (N_10704,N_9675,N_5561);
nand U10705 (N_10705,N_5342,N_7026);
nor U10706 (N_10706,N_7794,N_6870);
nand U10707 (N_10707,N_8819,N_7569);
or U10708 (N_10708,N_5805,N_8436);
xnor U10709 (N_10709,N_8144,N_9525);
xnor U10710 (N_10710,N_5931,N_8336);
nor U10711 (N_10711,N_9097,N_5391);
nor U10712 (N_10712,N_8924,N_6489);
and U10713 (N_10713,N_8728,N_7377);
nor U10714 (N_10714,N_5926,N_7949);
and U10715 (N_10715,N_7861,N_6615);
or U10716 (N_10716,N_7374,N_8807);
and U10717 (N_10717,N_6928,N_9549);
nand U10718 (N_10718,N_5823,N_8954);
nor U10719 (N_10719,N_8474,N_7787);
xor U10720 (N_10720,N_9338,N_6484);
nor U10721 (N_10721,N_9100,N_6800);
nor U10722 (N_10722,N_6847,N_7109);
and U10723 (N_10723,N_6202,N_6444);
nand U10724 (N_10724,N_5915,N_9441);
or U10725 (N_10725,N_9465,N_7865);
nor U10726 (N_10726,N_8137,N_7485);
nand U10727 (N_10727,N_6435,N_7823);
or U10728 (N_10728,N_7924,N_7849);
or U10729 (N_10729,N_7388,N_8830);
and U10730 (N_10730,N_6747,N_5091);
xnor U10731 (N_10731,N_9986,N_6244);
nand U10732 (N_10732,N_7836,N_9226);
or U10733 (N_10733,N_6315,N_7317);
nand U10734 (N_10734,N_8508,N_9644);
nand U10735 (N_10735,N_7533,N_8753);
nand U10736 (N_10736,N_7838,N_5581);
xnor U10737 (N_10737,N_8979,N_5358);
nand U10738 (N_10738,N_7029,N_9886);
xnor U10739 (N_10739,N_6746,N_5812);
and U10740 (N_10740,N_6280,N_6519);
or U10741 (N_10741,N_8299,N_9677);
or U10742 (N_10742,N_8629,N_7058);
nand U10743 (N_10743,N_7260,N_5868);
or U10744 (N_10744,N_6151,N_9524);
xnor U10745 (N_10745,N_9365,N_9535);
nor U10746 (N_10746,N_8832,N_6647);
nor U10747 (N_10747,N_9372,N_5923);
or U10748 (N_10748,N_8972,N_9741);
xor U10749 (N_10749,N_9489,N_8185);
nor U10750 (N_10750,N_6694,N_5368);
or U10751 (N_10751,N_9324,N_5454);
and U10752 (N_10752,N_8266,N_5549);
xor U10753 (N_10753,N_6019,N_5147);
or U10754 (N_10754,N_7943,N_8065);
or U10755 (N_10755,N_8489,N_5865);
xnor U10756 (N_10756,N_7567,N_6525);
nand U10757 (N_10757,N_8814,N_6455);
xor U10758 (N_10758,N_7042,N_5591);
or U10759 (N_10759,N_7278,N_6027);
and U10760 (N_10760,N_8789,N_6302);
xnor U10761 (N_10761,N_5215,N_6922);
or U10762 (N_10762,N_6745,N_7771);
and U10763 (N_10763,N_7329,N_8987);
or U10764 (N_10764,N_5052,N_7954);
or U10765 (N_10765,N_5716,N_8933);
xnor U10766 (N_10766,N_6505,N_6328);
nor U10767 (N_10767,N_8734,N_9587);
xnor U10768 (N_10768,N_6344,N_9444);
or U10769 (N_10769,N_5204,N_5062);
nand U10770 (N_10770,N_8658,N_6654);
nor U10771 (N_10771,N_8540,N_5888);
or U10772 (N_10772,N_7590,N_9956);
and U10773 (N_10773,N_5071,N_5877);
nor U10774 (N_10774,N_5120,N_6157);
or U10775 (N_10775,N_5677,N_6936);
nand U10776 (N_10776,N_7028,N_8994);
and U10777 (N_10777,N_9672,N_9728);
nor U10778 (N_10778,N_7696,N_6136);
or U10779 (N_10779,N_7518,N_5241);
xor U10780 (N_10780,N_5233,N_6815);
xor U10781 (N_10781,N_9344,N_7250);
and U10782 (N_10782,N_9909,N_5176);
nor U10783 (N_10783,N_8454,N_9714);
xor U10784 (N_10784,N_7650,N_5118);
and U10785 (N_10785,N_6271,N_5248);
or U10786 (N_10786,N_5314,N_8962);
xor U10787 (N_10787,N_9052,N_9184);
xnor U10788 (N_10788,N_5897,N_9820);
nand U10789 (N_10789,N_9580,N_9101);
or U10790 (N_10790,N_5133,N_5957);
and U10791 (N_10791,N_8829,N_6961);
nand U10792 (N_10792,N_7931,N_6638);
and U10793 (N_10793,N_6514,N_9457);
or U10794 (N_10794,N_5665,N_8775);
or U10795 (N_10795,N_6604,N_6382);
nand U10796 (N_10796,N_5863,N_6691);
nand U10797 (N_10797,N_7153,N_8304);
or U10798 (N_10798,N_7637,N_6925);
nor U10799 (N_10799,N_9809,N_7408);
and U10800 (N_10800,N_8524,N_5731);
and U10801 (N_10801,N_9054,N_9913);
xnor U10802 (N_10802,N_6664,N_7789);
or U10803 (N_10803,N_6397,N_9498);
and U10804 (N_10804,N_5163,N_9249);
nand U10805 (N_10805,N_8384,N_5808);
xnor U10806 (N_10806,N_6440,N_8125);
and U10807 (N_10807,N_5956,N_7473);
nor U10808 (N_10808,N_5776,N_6388);
nand U10809 (N_10809,N_7619,N_6164);
or U10810 (N_10810,N_8644,N_7083);
xnor U10811 (N_10811,N_8176,N_8895);
xnor U10812 (N_10812,N_9132,N_5696);
and U10813 (N_10813,N_8887,N_6564);
xnor U10814 (N_10814,N_5803,N_5947);
and U10815 (N_10815,N_7868,N_7334);
nor U10816 (N_10816,N_9171,N_5815);
and U10817 (N_10817,N_5537,N_8975);
nor U10818 (N_10818,N_8709,N_6065);
or U10819 (N_10819,N_8609,N_8747);
and U10820 (N_10820,N_5693,N_6990);
nor U10821 (N_10821,N_6764,N_8915);
or U10822 (N_10822,N_5240,N_9616);
or U10823 (N_10823,N_8287,N_9045);
nand U10824 (N_10824,N_5260,N_8843);
xor U10825 (N_10825,N_6835,N_6817);
nand U10826 (N_10826,N_9763,N_6443);
xnor U10827 (N_10827,N_7261,N_7406);
nand U10828 (N_10828,N_6230,N_7382);
or U10829 (N_10829,N_7745,N_5078);
or U10830 (N_10830,N_9776,N_6971);
nor U10831 (N_10831,N_7765,N_5444);
or U10832 (N_10832,N_6518,N_6700);
xnor U10833 (N_10833,N_7809,N_7585);
and U10834 (N_10834,N_6805,N_9134);
or U10835 (N_10835,N_8448,N_8783);
nand U10836 (N_10836,N_6610,N_8558);
and U10837 (N_10837,N_6463,N_9178);
and U10838 (N_10838,N_5002,N_7587);
nand U10839 (N_10839,N_7523,N_7498);
or U10840 (N_10840,N_9661,N_6609);
xnor U10841 (N_10841,N_5090,N_6756);
and U10842 (N_10842,N_9756,N_8656);
nand U10843 (N_10843,N_5752,N_7335);
xor U10844 (N_10844,N_7888,N_8928);
and U10845 (N_10845,N_6786,N_7933);
xor U10846 (N_10846,N_5563,N_6727);
and U10847 (N_10847,N_6060,N_5927);
or U10848 (N_10848,N_6055,N_7866);
nor U10849 (N_10849,N_5445,N_7349);
nor U10850 (N_10850,N_9404,N_5465);
xor U10851 (N_10851,N_8411,N_7814);
nand U10852 (N_10852,N_7737,N_7091);
nand U10853 (N_10853,N_8066,N_8795);
nand U10854 (N_10854,N_5437,N_5748);
nand U10855 (N_10855,N_9174,N_8292);
nor U10856 (N_10856,N_9433,N_9407);
xnor U10857 (N_10857,N_9164,N_9752);
or U10858 (N_10858,N_7003,N_6237);
xor U10859 (N_10859,N_8246,N_5831);
and U10860 (N_10860,N_8349,N_9912);
and U10861 (N_10861,N_8230,N_5982);
nor U10862 (N_10862,N_5095,N_9502);
or U10863 (N_10863,N_9216,N_8133);
xnor U10864 (N_10864,N_9499,N_8953);
nor U10865 (N_10865,N_6978,N_5936);
or U10866 (N_10866,N_6858,N_7673);
or U10867 (N_10867,N_9868,N_9180);
xor U10868 (N_10868,N_6013,N_5615);
and U10869 (N_10869,N_5662,N_7779);
or U10870 (N_10870,N_9242,N_5276);
nor U10871 (N_10871,N_9597,N_9183);
and U10872 (N_10872,N_6325,N_8880);
nor U10873 (N_10873,N_7581,N_8437);
or U10874 (N_10874,N_8774,N_6773);
and U10875 (N_10875,N_7705,N_7477);
nand U10876 (N_10876,N_9769,N_9452);
xnor U10877 (N_10877,N_8601,N_6332);
nand U10878 (N_10878,N_9980,N_9722);
nand U10879 (N_10879,N_8056,N_8241);
and U10880 (N_10880,N_7048,N_5193);
nand U10881 (N_10881,N_6759,N_9543);
xnor U10882 (N_10882,N_7853,N_7269);
nor U10883 (N_10883,N_7096,N_7600);
or U10884 (N_10884,N_9398,N_6442);
and U10885 (N_10885,N_6298,N_7032);
nor U10886 (N_10886,N_6127,N_6232);
nand U10887 (N_10887,N_9315,N_9321);
nor U10888 (N_10888,N_5289,N_6285);
nor U10889 (N_10889,N_5048,N_6716);
nor U10890 (N_10890,N_7947,N_8672);
nor U10891 (N_10891,N_5222,N_8174);
nor U10892 (N_10892,N_5154,N_8717);
nand U10893 (N_10893,N_7063,N_5027);
nand U10894 (N_10894,N_8735,N_7272);
or U10895 (N_10895,N_9117,N_8622);
and U10896 (N_10896,N_8503,N_9161);
nor U10897 (N_10897,N_8069,N_5049);
xor U10898 (N_10898,N_6974,N_9373);
nor U10899 (N_10899,N_5968,N_9629);
nor U10900 (N_10900,N_8950,N_7871);
xnor U10901 (N_10901,N_9453,N_6836);
and U10902 (N_10902,N_6303,N_5502);
and U10903 (N_10903,N_5667,N_7357);
nand U10904 (N_10904,N_8720,N_6365);
nand U10905 (N_10905,N_7875,N_6128);
nand U10906 (N_10906,N_9013,N_6679);
and U10907 (N_10907,N_9824,N_6394);
and U10908 (N_10908,N_6346,N_8892);
nand U10909 (N_10909,N_5747,N_7392);
xnor U10910 (N_10910,N_7276,N_9788);
nor U10911 (N_10911,N_8557,N_7618);
nand U10912 (N_10912,N_9327,N_6385);
or U10913 (N_10913,N_8708,N_6051);
or U10914 (N_10914,N_7253,N_5040);
xor U10915 (N_10915,N_7766,N_8086);
and U10916 (N_10916,N_6545,N_6888);
nand U10917 (N_10917,N_9206,N_9495);
and U10918 (N_10918,N_6356,N_8580);
nor U10919 (N_10919,N_9458,N_8355);
nor U10920 (N_10920,N_7945,N_9286);
nor U10921 (N_10921,N_7689,N_6347);
nand U10922 (N_10922,N_8468,N_9780);
nor U10923 (N_10923,N_5698,N_8062);
and U10924 (N_10924,N_8128,N_8154);
or U10925 (N_10925,N_7826,N_9009);
nand U10926 (N_10926,N_7090,N_7119);
xor U10927 (N_10927,N_8310,N_5609);
nor U10928 (N_10928,N_8615,N_5544);
nor U10929 (N_10929,N_6840,N_9702);
nor U10930 (N_10930,N_7039,N_7052);
and U10931 (N_10931,N_9845,N_5418);
nand U10932 (N_10932,N_6175,N_6673);
nand U10933 (N_10933,N_7086,N_8451);
and U10934 (N_10934,N_8919,N_9065);
and U10935 (N_10935,N_7369,N_5997);
or U10936 (N_10936,N_8225,N_7396);
xnor U10937 (N_10937,N_7670,N_8893);
nand U10938 (N_10938,N_7162,N_6774);
or U10939 (N_10939,N_8512,N_9799);
nand U10940 (N_10940,N_8326,N_8206);
nand U10941 (N_10941,N_9724,N_8724);
nor U10942 (N_10942,N_8160,N_9253);
xnor U10943 (N_10943,N_7088,N_6188);
nand U10944 (N_10944,N_9342,N_8115);
or U10945 (N_10945,N_7115,N_8135);
nand U10946 (N_10946,N_8035,N_9806);
xor U10947 (N_10947,N_6095,N_7446);
xor U10948 (N_10948,N_5775,N_6837);
nor U10949 (N_10949,N_9170,N_8897);
nand U10950 (N_10950,N_8697,N_8482);
or U10951 (N_10951,N_6084,N_9772);
or U10952 (N_10952,N_7194,N_5135);
or U10953 (N_10953,N_9782,N_5021);
nor U10954 (N_10954,N_9833,N_6129);
xor U10955 (N_10955,N_9881,N_9123);
nand U10956 (N_10956,N_8293,N_6399);
and U10957 (N_10957,N_5506,N_5562);
nor U10958 (N_10958,N_7371,N_6270);
nor U10959 (N_10959,N_9128,N_6014);
nand U10960 (N_10960,N_7835,N_6809);
or U10961 (N_10961,N_8008,N_6696);
and U10962 (N_10962,N_5535,N_7967);
or U10963 (N_10963,N_7187,N_5295);
or U10964 (N_10964,N_5854,N_9596);
xor U10965 (N_10965,N_5498,N_5788);
or U10966 (N_10966,N_8101,N_5278);
nor U10967 (N_10967,N_9085,N_9475);
nand U10968 (N_10968,N_6383,N_8139);
and U10969 (N_10969,N_5902,N_7824);
xor U10970 (N_10970,N_5199,N_5794);
nand U10971 (N_10971,N_5694,N_6169);
or U10972 (N_10972,N_9821,N_5146);
nor U10973 (N_10973,N_8273,N_6945);
nor U10974 (N_10974,N_5622,N_7712);
and U10975 (N_10975,N_6119,N_8509);
and U10976 (N_10976,N_5128,N_5878);
nand U10977 (N_10977,N_5375,N_5008);
xnor U10978 (N_10978,N_6980,N_5247);
nand U10979 (N_10979,N_9509,N_9815);
or U10980 (N_10980,N_6548,N_5940);
nand U10981 (N_10981,N_9503,N_8184);
and U10982 (N_10982,N_8531,N_5727);
nand U10983 (N_10983,N_6901,N_7904);
or U10984 (N_10984,N_5319,N_8956);
nor U10985 (N_10985,N_9935,N_9841);
or U10986 (N_10986,N_8847,N_6792);
nand U10987 (N_10987,N_7461,N_6185);
nand U10988 (N_10988,N_8903,N_9314);
or U10989 (N_10989,N_7621,N_5848);
xnor U10990 (N_10990,N_7087,N_6363);
xor U10991 (N_10991,N_9943,N_7075);
nand U10992 (N_10992,N_8586,N_5003);
xnor U10993 (N_10993,N_6625,N_5834);
or U10994 (N_10994,N_5514,N_7893);
and U10995 (N_10995,N_9803,N_6160);
xor U10996 (N_10996,N_5750,N_5835);
nor U10997 (N_10997,N_6460,N_5896);
nor U10998 (N_10998,N_8256,N_7976);
xnor U10999 (N_10999,N_5487,N_6635);
nor U11000 (N_11000,N_9260,N_8269);
or U11001 (N_11001,N_8669,N_7528);
or U11002 (N_11002,N_5327,N_7144);
xnor U11003 (N_11003,N_9214,N_7173);
nor U11004 (N_11004,N_6153,N_5291);
and U11005 (N_11005,N_8060,N_6795);
nor U11006 (N_11006,N_6293,N_6205);
xnor U11007 (N_11007,N_7170,N_8649);
xor U11008 (N_11008,N_9004,N_7370);
nor U11009 (N_11009,N_9488,N_7005);
nand U11010 (N_11010,N_6821,N_7683);
and U11011 (N_11011,N_7797,N_8862);
nor U11012 (N_11012,N_9241,N_5205);
xnor U11013 (N_11013,N_6361,N_5688);
nor U11014 (N_11014,N_7648,N_8834);
xnor U11015 (N_11015,N_7676,N_9438);
xor U11016 (N_11016,N_5586,N_5709);
nor U11017 (N_11017,N_7573,N_9829);
or U11018 (N_11018,N_7235,N_9892);
nor U11019 (N_11019,N_6658,N_5271);
or U11020 (N_11020,N_5489,N_7106);
or U11021 (N_11021,N_6504,N_9614);
nand U11022 (N_11022,N_7729,N_6499);
or U11023 (N_11023,N_8605,N_9822);
nor U11024 (N_11024,N_9915,N_8208);
nand U11025 (N_11025,N_7599,N_9354);
xnor U11026 (N_11026,N_8838,N_8585);
nand U11027 (N_11027,N_7642,N_6450);
nor U11028 (N_11028,N_5151,N_8263);
xnor U11029 (N_11029,N_9328,N_5801);
and U11030 (N_11030,N_9190,N_7604);
xor U11031 (N_11031,N_5890,N_5397);
nand U11032 (N_11032,N_7986,N_5792);
and U11033 (N_11033,N_9919,N_9470);
or U11034 (N_11034,N_9353,N_9859);
nor U11035 (N_11035,N_6339,N_6286);
xor U11036 (N_11036,N_9931,N_5328);
nor U11037 (N_11037,N_7512,N_7508);
nand U11038 (N_11038,N_9251,N_9818);
and U11039 (N_11039,N_6630,N_8367);
and U11040 (N_11040,N_6166,N_7453);
nor U11041 (N_11041,N_6043,N_9396);
nor U11042 (N_11042,N_6467,N_8659);
nand U11043 (N_11043,N_8057,N_8548);
xor U11044 (N_11044,N_9625,N_5348);
xnor U11045 (N_11045,N_5971,N_9689);
nor U11046 (N_11046,N_9084,N_7167);
and U11047 (N_11047,N_6571,N_6478);
xnor U11048 (N_11048,N_9090,N_7634);
and U11049 (N_11049,N_7830,N_6334);
xnor U11050 (N_11050,N_8316,N_6037);
nor U11051 (N_11051,N_5477,N_6572);
and U11052 (N_11052,N_8258,N_5882);
xor U11053 (N_11053,N_7448,N_7421);
or U11054 (N_11054,N_7404,N_7230);
xor U11055 (N_11055,N_7321,N_5580);
nand U11056 (N_11056,N_5827,N_5725);
nor U11057 (N_11057,N_8803,N_6547);
nor U11058 (N_11058,N_5322,N_7360);
and U11059 (N_11059,N_7772,N_8908);
xnor U11060 (N_11060,N_5879,N_8486);
nor U11061 (N_11061,N_5866,N_9283);
nand U11062 (N_11062,N_6783,N_7163);
nor U11063 (N_11063,N_9264,N_9719);
nor U11064 (N_11064,N_7341,N_6149);
nand U11065 (N_11065,N_7358,N_7089);
nor U11066 (N_11066,N_5287,N_8675);
or U11067 (N_11067,N_7336,N_7359);
or U11068 (N_11068,N_8321,N_8005);
and U11069 (N_11069,N_9745,N_9310);
xor U11070 (N_11070,N_5552,N_8267);
or U11071 (N_11071,N_6902,N_8240);
or U11072 (N_11072,N_7175,N_7381);
nor U11073 (N_11073,N_7920,N_5649);
and U11074 (N_11074,N_6887,N_5557);
nand U11075 (N_11075,N_7740,N_6236);
nor U11076 (N_11076,N_5634,N_5525);
and U11077 (N_11077,N_9074,N_5521);
nand U11078 (N_11078,N_5761,N_8833);
nand U11079 (N_11079,N_6632,N_8589);
or U11080 (N_11080,N_9898,N_7311);
xor U11081 (N_11081,N_5921,N_7229);
nor U11082 (N_11082,N_5666,N_9897);
and U11083 (N_11083,N_5668,N_9384);
xnor U11084 (N_11084,N_5884,N_8960);
nor U11085 (N_11085,N_7641,N_5555);
xnor U11086 (N_11086,N_9202,N_5096);
and U11087 (N_11087,N_7944,N_6098);
and U11088 (N_11088,N_9879,N_5316);
xnor U11089 (N_11089,N_7220,N_6447);
xor U11090 (N_11090,N_9517,N_8191);
and U11091 (N_11091,N_7630,N_8284);
and U11092 (N_11092,N_8348,N_9713);
and U11093 (N_11093,N_6827,N_6581);
nand U11094 (N_11094,N_9348,N_5760);
nand U11095 (N_11095,N_8606,N_8997);
nor U11096 (N_11096,N_8076,N_5236);
nor U11097 (N_11097,N_6956,N_7639);
nand U11098 (N_11098,N_8732,N_6367);
xor U11099 (N_11099,N_5057,N_9602);
and U11100 (N_11100,N_7270,N_9477);
nor U11101 (N_11101,N_7892,N_5565);
and U11102 (N_11102,N_6642,N_5809);
nand U11103 (N_11103,N_8912,N_8315);
xnor U11104 (N_11104,N_8875,N_8976);
xor U11105 (N_11105,N_7496,N_8810);
nor U11106 (N_11106,N_8311,N_7623);
nor U11107 (N_11107,N_5159,N_7353);
nand U11108 (N_11108,N_6002,N_8816);
xor U11109 (N_11109,N_7012,N_5041);
nand U11110 (N_11110,N_6101,N_8635);
nand U11111 (N_11111,N_7505,N_9018);
and U11112 (N_11112,N_8959,N_7710);
nand U11113 (N_11113,N_9142,N_7919);
and U11114 (N_11114,N_7306,N_6432);
xnor U11115 (N_11115,N_5670,N_7136);
nand U11116 (N_11116,N_7576,N_9345);
xor U11117 (N_11117,N_5250,N_9558);
nand U11118 (N_11118,N_7701,N_8425);
and U11119 (N_11119,N_9529,N_9996);
nand U11120 (N_11120,N_8802,N_7403);
nand U11121 (N_11121,N_7264,N_6301);
nor U11122 (N_11122,N_8010,N_8570);
nor U11123 (N_11123,N_6911,N_9725);
nor U11124 (N_11124,N_9412,N_8165);
and U11125 (N_11125,N_5543,N_9789);
nor U11126 (N_11126,N_8067,N_9238);
and U11127 (N_11127,N_6998,N_6483);
nor U11128 (N_11128,N_9400,N_6957);
or U11129 (N_11129,N_8642,N_9658);
nor U11130 (N_11130,N_8796,N_5578);
xnor U11131 (N_11131,N_6052,N_9308);
or U11132 (N_11132,N_8376,N_7390);
nand U11133 (N_11133,N_7660,N_7568);
xor U11134 (N_11134,N_7467,N_7345);
and U11135 (N_11135,N_7489,N_7389);
and U11136 (N_11136,N_8527,N_5182);
or U11137 (N_11137,N_7445,N_8650);
and U11138 (N_11138,N_8595,N_8417);
or U11139 (N_11139,N_9938,N_8396);
nor U11140 (N_11140,N_6758,N_5100);
nand U11141 (N_11141,N_5534,N_9623);
nor U11142 (N_11142,N_9654,N_6893);
xor U11143 (N_11143,N_8921,N_8136);
or U11144 (N_11144,N_6524,N_6766);
nand U11145 (N_11145,N_9131,N_6081);
and U11146 (N_11146,N_8731,N_6429);
and U11147 (N_11147,N_9022,N_7401);
nor U11148 (N_11148,N_7245,N_7224);
or U11149 (N_11149,N_5771,N_6126);
nand U11150 (N_11150,N_9059,N_7251);
xor U11151 (N_11151,N_8073,N_8331);
and U11152 (N_11152,N_7425,N_8932);
or U11153 (N_11153,N_8631,N_8435);
xor U11154 (N_11154,N_5268,N_8902);
or U11155 (N_11155,N_8025,N_6498);
and U11156 (N_11156,N_8616,N_8848);
and U11157 (N_11157,N_6086,N_8369);
and U11158 (N_11158,N_9890,N_6622);
or U11159 (N_11159,N_6871,N_5101);
nand U11160 (N_11160,N_8528,N_7292);
nor U11161 (N_11161,N_9957,N_8667);
and U11162 (N_11162,N_6187,N_6844);
and U11163 (N_11163,N_9299,N_7420);
nand U11164 (N_11164,N_8502,N_8483);
nand U11165 (N_11165,N_9720,N_7840);
nand U11166 (N_11166,N_7819,N_7679);
or U11167 (N_11167,N_5491,N_8007);
nor U11168 (N_11168,N_9651,N_6393);
xor U11169 (N_11169,N_7238,N_9848);
nand U11170 (N_11170,N_6015,N_6569);
and U11171 (N_11171,N_9274,N_7914);
xor U11172 (N_11172,N_5907,N_9119);
nand U11173 (N_11173,N_7594,N_8811);
nor U11174 (N_11174,N_5353,N_6896);
xnor U11175 (N_11175,N_6643,N_9668);
and U11176 (N_11176,N_8780,N_9690);
nor U11177 (N_11177,N_5585,N_6626);
xor U11178 (N_11178,N_8054,N_9089);
and U11179 (N_11179,N_9432,N_9415);
and U11180 (N_11180,N_6267,N_8693);
xnor U11181 (N_11181,N_6933,N_5061);
nor U11182 (N_11182,N_6040,N_9942);
nand U11183 (N_11183,N_8465,N_6636);
and U11184 (N_11184,N_6775,N_6078);
nand U11185 (N_11185,N_6981,N_5681);
nor U11186 (N_11186,N_5718,N_7833);
or U11187 (N_11187,N_8283,N_9079);
and U11188 (N_11188,N_9288,N_6324);
nand U11189 (N_11189,N_8640,N_6284);
or U11190 (N_11190,N_5942,N_6885);
or U11191 (N_11191,N_6618,N_9751);
nor U11192 (N_11192,N_8869,N_9920);
and U11193 (N_11193,N_6253,N_7767);
nor U11194 (N_11194,N_7168,N_9685);
and U11195 (N_11195,N_6005,N_8359);
and U11196 (N_11196,N_7964,N_7859);
or U11197 (N_11197,N_5964,N_8759);
and U11198 (N_11198,N_8357,N_6165);
nand U11199 (N_11199,N_9145,N_5641);
xnor U11200 (N_11200,N_6791,N_9583);
nor U11201 (N_11201,N_5175,N_7085);
nand U11202 (N_11202,N_5377,N_7142);
xnor U11203 (N_11203,N_6183,N_9225);
xnor U11204 (N_11204,N_6863,N_6220);
nand U11205 (N_11205,N_8823,N_9068);
and U11206 (N_11206,N_5601,N_7957);
nor U11207 (N_11207,N_9775,N_6254);
xnor U11208 (N_11208,N_7795,N_6586);
and U11209 (N_11209,N_9736,N_7385);
nand U11210 (N_11210,N_7829,N_6152);
and U11211 (N_11211,N_5500,N_9600);
and U11212 (N_11212,N_6999,N_8682);
or U11213 (N_11213,N_5141,N_8236);
nor U11214 (N_11214,N_6670,N_5974);
and U11215 (N_11215,N_6667,N_8984);
nor U11216 (N_11216,N_7774,N_8416);
and U11217 (N_11217,N_6814,N_8244);
and U11218 (N_11218,N_8991,N_8476);
nor U11219 (N_11219,N_9599,N_5371);
and U11220 (N_11220,N_7714,N_7120);
xnor U11221 (N_11221,N_8146,N_8591);
or U11222 (N_11222,N_9941,N_9877);
and U11223 (N_11223,N_9367,N_7562);
nor U11224 (N_11224,N_5467,N_7430);
xor U11225 (N_11225,N_7908,N_8026);
nand U11226 (N_11226,N_5770,N_9049);
or U11227 (N_11227,N_5006,N_8216);
and U11228 (N_11228,N_5034,N_6452);
xor U11229 (N_11229,N_7066,N_7657);
nor U11230 (N_11230,N_6380,N_5545);
xor U11231 (N_11231,N_8201,N_6321);
and U11232 (N_11232,N_6580,N_7082);
or U11233 (N_11233,N_7481,N_9179);
or U11234 (N_11234,N_8863,N_8081);
or U11235 (N_11235,N_6091,N_8866);
nor U11236 (N_11236,N_9887,N_5475);
nor U11237 (N_11237,N_9343,N_6913);
xnor U11238 (N_11238,N_7516,N_8894);
xnor U11239 (N_11239,N_8490,N_6105);
and U11240 (N_11240,N_9198,N_9102);
xnor U11241 (N_11241,N_7956,N_5108);
xor U11242 (N_11242,N_9992,N_5401);
and U11243 (N_11243,N_8652,N_9472);
nand U11244 (N_11244,N_5899,N_6824);
nand U11245 (N_11245,N_5919,N_6387);
xnor U11246 (N_11246,N_9641,N_8300);
nand U11247 (N_11247,N_8846,N_5419);
xor U11248 (N_11248,N_8748,N_7419);
and U11249 (N_11249,N_6307,N_7832);
nand U11250 (N_11250,N_6573,N_5211);
and U11251 (N_11251,N_8668,N_7149);
and U11252 (N_11252,N_7666,N_7013);
xnor U11253 (N_11253,N_9479,N_7208);
nand U11254 (N_11254,N_9331,N_9835);
or U11255 (N_11255,N_8289,N_7817);
xnor U11256 (N_11256,N_9449,N_9478);
and U11257 (N_11257,N_6816,N_7778);
nand U11258 (N_11258,N_5855,N_7950);
and U11259 (N_11259,N_9233,N_8082);
or U11260 (N_11260,N_8285,N_6403);
and U11261 (N_11261,N_8168,N_9974);
nor U11262 (N_11262,N_7018,N_6147);
xor U11263 (N_11263,N_8945,N_9244);
or U11264 (N_11264,N_9846,N_5969);
and U11265 (N_11265,N_5346,N_9839);
nand U11266 (N_11266,N_5055,N_8166);
and U11267 (N_11267,N_8612,N_7047);
nor U11268 (N_11268,N_7891,N_6937);
xnor U11269 (N_11269,N_6946,N_7723);
nand U11270 (N_11270,N_5988,N_8582);
and U11271 (N_11271,N_9057,N_6449);
nand U11272 (N_11272,N_9642,N_7366);
or U11273 (N_11273,N_6206,N_8012);
nand U11274 (N_11274,N_5023,N_7882);
and U11275 (N_11275,N_5106,N_6533);
or U11276 (N_11276,N_6214,N_9095);
and U11277 (N_11277,N_6575,N_7285);
nand U11278 (N_11278,N_5659,N_9322);
and U11279 (N_11279,N_9435,N_8877);
nand U11280 (N_11280,N_7146,N_6964);
and U11281 (N_11281,N_8520,N_5513);
nor U11282 (N_11282,N_7730,N_8092);
xor U11283 (N_11283,N_9617,N_7851);
xnor U11284 (N_11284,N_5372,N_8598);
nor U11285 (N_11285,N_8171,N_5259);
nor U11286 (N_11286,N_6912,N_6333);
and U11287 (N_11287,N_8700,N_7970);
nand U11288 (N_11288,N_5225,N_5196);
nand U11289 (N_11289,N_6398,N_8181);
xnor U11290 (N_11290,N_7597,N_6415);
or U11291 (N_11291,N_7509,N_6690);
nor U11292 (N_11292,N_8852,N_7067);
and U11293 (N_11293,N_5395,N_7869);
nor U11294 (N_11294,N_8404,N_6090);
and U11295 (N_11295,N_5201,N_7290);
or U11296 (N_11296,N_9884,N_5664);
nand U11297 (N_11297,N_6125,N_6208);
xor U11298 (N_11298,N_5255,N_8804);
and U11299 (N_11299,N_6793,N_8340);
nor U11300 (N_11300,N_8536,N_5507);
nor U11301 (N_11301,N_7525,N_9900);
and U11302 (N_11302,N_9627,N_6588);
nand U11303 (N_11303,N_7811,N_6603);
or U11304 (N_11304,N_5094,N_7111);
or U11305 (N_11305,N_5901,N_6637);
and U11306 (N_11306,N_7524,N_7211);
nand U11307 (N_11307,N_9885,N_8446);
or U11308 (N_11308,N_6926,N_9573);
nand U11309 (N_11309,N_6007,N_9921);
nand U11310 (N_11310,N_8534,N_8344);
and U11311 (N_11311,N_7757,N_9715);
or U11312 (N_11312,N_5001,N_9456);
or U11313 (N_11313,N_8419,N_7937);
xor U11314 (N_11314,N_7746,N_9466);
nand U11315 (N_11315,N_6376,N_5009);
nor U11316 (N_11316,N_7514,N_5473);
nor U11317 (N_11317,N_6752,N_6583);
nor U11318 (N_11318,N_7084,N_6409);
or U11319 (N_11319,N_9902,N_8428);
nor U11320 (N_11320,N_6983,N_8303);
nor U11321 (N_11321,N_7070,N_7112);
nor U11322 (N_11322,N_8806,N_9265);
and U11323 (N_11323,N_5646,N_6103);
nand U11324 (N_11324,N_9812,N_9270);
nand U11325 (N_11325,N_6215,N_8363);
nor U11326 (N_11326,N_7024,N_5157);
xor U11327 (N_11327,N_5623,N_9766);
nand U11328 (N_11328,N_6283,N_7544);
or U11329 (N_11329,N_8985,N_6530);
nor U11330 (N_11330,N_6751,N_9768);
nor U11331 (N_11331,N_9564,N_9437);
xor U11332 (N_11332,N_5642,N_8562);
nor U11333 (N_11333,N_8141,N_8722);
xnor U11334 (N_11334,N_6292,N_5611);
nor U11335 (N_11335,N_7969,N_5181);
or U11336 (N_11336,N_5583,N_8068);
nor U11337 (N_11337,N_6291,N_6866);
nand U11338 (N_11338,N_8272,N_5046);
or U11339 (N_11339,N_6526,N_8899);
or U11340 (N_11340,N_9819,N_7550);
or U11341 (N_11341,N_5463,N_5216);
nand U11342 (N_11342,N_9108,N_5682);
and U11343 (N_11343,N_5976,N_7400);
nor U11344 (N_11344,N_5708,N_9347);
nand U11345 (N_11345,N_6879,N_9236);
or U11346 (N_11346,N_9133,N_9067);
or U11347 (N_11347,N_8392,N_6704);
xor U11348 (N_11348,N_7221,N_6396);
and U11349 (N_11349,N_9248,N_9154);
and U11350 (N_11350,N_7200,N_8205);
and U11351 (N_11351,N_6616,N_9355);
and U11352 (N_11352,N_7678,N_9006);
xnor U11353 (N_11353,N_5702,N_9657);
or U11354 (N_11354,N_7133,N_8248);
and U11355 (N_11355,N_9212,N_5724);
or U11356 (N_11356,N_5676,N_6951);
or U11357 (N_11357,N_9038,N_8792);
nor U11358 (N_11358,N_9565,N_6839);
nor U11359 (N_11359,N_5388,N_6057);
nand U11360 (N_11360,N_8328,N_7520);
nand U11361 (N_11361,N_8873,N_6650);
and U11362 (N_11362,N_5360,N_5531);
xnor U11363 (N_11363,N_5386,N_8302);
nor U11364 (N_11364,N_7526,N_9547);
xor U11365 (N_11365,N_6199,N_9122);
and U11366 (N_11366,N_8955,N_9734);
nor U11367 (N_11367,N_8523,N_6938);
xnor U11368 (N_11368,N_5987,N_8799);
nor U11369 (N_11369,N_5025,N_7118);
nand U11370 (N_11370,N_8982,N_9663);
and U11371 (N_11371,N_7071,N_7825);
nor U11372 (N_11372,N_6277,N_9364);
and U11373 (N_11373,N_8319,N_9687);
nor U11374 (N_11374,N_6073,N_7060);
nor U11375 (N_11375,N_5765,N_6724);
nor U11376 (N_11376,N_9523,N_8237);
nor U11377 (N_11377,N_8473,N_7344);
or U11378 (N_11378,N_6308,N_5556);
or U11379 (N_11379,N_5864,N_5485);
and U11380 (N_11380,N_7691,N_6876);
or U11381 (N_11381,N_8387,N_8198);
and U11382 (N_11382,N_9126,N_9874);
and U11383 (N_11383,N_9500,N_6074);
nor U11384 (N_11384,N_8971,N_7101);
nand U11385 (N_11385,N_5466,N_6108);
and U11386 (N_11386,N_5093,N_7008);
nor U11387 (N_11387,N_6316,N_8120);
nand U11388 (N_11388,N_6787,N_8691);
nand U11389 (N_11389,N_5160,N_7046);
nor U11390 (N_11390,N_7169,N_6250);
or U11391 (N_11391,N_9278,N_6413);
xor U11392 (N_11392,N_9653,N_5410);
or U11393 (N_11393,N_8164,N_5341);
xor U11394 (N_11394,N_9012,N_9552);
nor U11395 (N_11395,N_7080,N_9450);
or U11396 (N_11396,N_9634,N_8381);
nor U11397 (N_11397,N_5257,N_7409);
nor U11398 (N_11398,N_9934,N_9187);
nor U11399 (N_11399,N_5136,N_7975);
nor U11400 (N_11400,N_7191,N_6892);
and U11401 (N_11401,N_8714,N_6439);
nand U11402 (N_11402,N_6666,N_8309);
or U11403 (N_11403,N_9723,N_7262);
or U11404 (N_11404,N_5494,N_9635);
and U11405 (N_11405,N_7432,N_7102);
or U11406 (N_11406,N_9058,N_8794);
and U11407 (N_11407,N_6994,N_5857);
xnor U11408 (N_11408,N_7834,N_6400);
xnor U11409 (N_11409,N_8657,N_5793);
nand U11410 (N_11410,N_5517,N_7928);
xnor U11411 (N_11411,N_9589,N_6985);
or U11412 (N_11412,N_9638,N_6225);
nor U11413 (N_11413,N_7602,N_6712);
or U11414 (N_11414,N_8750,N_6551);
nor U11415 (N_11415,N_5280,N_6832);
nand U11416 (N_11416,N_6646,N_5115);
nand U11417 (N_11417,N_9598,N_9366);
or U11418 (N_11418,N_8857,N_9853);
nand U11419 (N_11419,N_9740,N_7495);
and U11420 (N_11420,N_6041,N_5584);
nor U11421 (N_11421,N_5456,N_6780);
or U11422 (N_11422,N_6340,N_7704);
nand U11423 (N_11423,N_5632,N_9771);
xor U11424 (N_11424,N_5845,N_7459);
nor U11425 (N_11425,N_5991,N_5451);
and U11426 (N_11426,N_6411,N_8413);
and U11427 (N_11427,N_9673,N_8122);
and U11428 (N_11428,N_8432,N_7632);
nor U11429 (N_11429,N_6614,N_8207);
xnor U11430 (N_11430,N_7463,N_9146);
or U11431 (N_11431,N_6163,N_7474);
or U11432 (N_11432,N_6258,N_7773);
nor U11433 (N_11433,N_5962,N_8022);
xor U11434 (N_11434,N_7612,N_5441);
nand U11435 (N_11435,N_5703,N_5599);
nand U11436 (N_11436,N_5566,N_5618);
or U11437 (N_11437,N_6466,N_5740);
or U11438 (N_11438,N_6995,N_8529);
and U11439 (N_11439,N_9403,N_6170);
and U11440 (N_11440,N_9754,N_9711);
or U11441 (N_11441,N_5186,N_6279);
nor U11442 (N_11442,N_5777,N_8200);
or U11443 (N_11443,N_7226,N_7108);
xnor U11444 (N_11444,N_7874,N_8556);
nor U11445 (N_11445,N_9855,N_9222);
nor U11446 (N_11446,N_5457,N_8495);
or U11447 (N_11447,N_6492,N_8189);
nand U11448 (N_11448,N_5440,N_5914);
nor U11449 (N_11449,N_6918,N_7592);
or U11450 (N_11450,N_7622,N_5024);
nor U11451 (N_11451,N_7415,N_7843);
nor U11452 (N_11452,N_8422,N_5228);
nand U11453 (N_11453,N_9246,N_9201);
or U11454 (N_11454,N_8253,N_6606);
xor U11455 (N_11455,N_7973,N_9816);
nand U11456 (N_11456,N_5393,N_5434);
or U11457 (N_11457,N_8818,N_8441);
or U11458 (N_11458,N_7663,N_9911);
or U11459 (N_11459,N_9420,N_5746);
or U11460 (N_11460,N_9041,N_5939);
nand U11461 (N_11461,N_7110,N_7354);
nand U11462 (N_11462,N_6851,N_7725);
nor U11463 (N_11463,N_5869,N_9847);
nand U11464 (N_11464,N_9497,N_5856);
nor U11465 (N_11465,N_8983,N_7996);
nor U11466 (N_11466,N_8579,N_8665);
nand U11467 (N_11467,N_8427,N_7653);
and U11468 (N_11468,N_8861,N_8294);
nand U11469 (N_11469,N_5647,N_9219);
nand U11470 (N_11470,N_9141,N_8061);
and U11471 (N_11471,N_6967,N_6117);
nor U11472 (N_11472,N_7092,N_9159);
nand U11473 (N_11473,N_7935,N_7372);
or U11474 (N_11474,N_8491,N_8710);
or U11475 (N_11475,N_7598,N_8778);
xnor U11476 (N_11476,N_8859,N_5277);
xor U11477 (N_11477,N_6210,N_5429);
nand U11478 (N_11478,N_8970,N_7727);
xor U11479 (N_11479,N_9483,N_8196);
nor U11480 (N_11480,N_9959,N_5625);
xnor U11481 (N_11481,N_7348,N_7297);
nand U11482 (N_11482,N_9650,N_5082);
xnor U11483 (N_11483,N_5994,N_5261);
xnor U11484 (N_11484,N_7428,N_8779);
nor U11485 (N_11485,N_6592,N_7801);
nor U11486 (N_11486,N_9304,N_7966);
nand U11487 (N_11487,N_6075,N_7503);
nand U11488 (N_11488,N_6651,N_6097);
xor U11489 (N_11489,N_9227,N_8513);
nand U11490 (N_11490,N_9061,N_8091);
xnor U11491 (N_11491,N_6242,N_5403);
and U11492 (N_11492,N_7241,N_9064);
nor U11493 (N_11493,N_7283,N_5686);
or U11494 (N_11494,N_8574,N_9866);
xor U11495 (N_11495,N_8167,N_8004);
nor U11496 (N_11496,N_7464,N_6145);
and U11497 (N_11497,N_6743,N_5488);
or U11498 (N_11498,N_9893,N_9660);
nor U11499 (N_11499,N_8566,N_8865);
nand U11500 (N_11500,N_5084,N_9764);
or U11501 (N_11501,N_5190,N_9410);
xor U11502 (N_11502,N_5651,N_9860);
and U11503 (N_11503,N_9810,N_5449);
nor U11504 (N_11504,N_7695,N_9906);
xor U11505 (N_11505,N_9175,N_9312);
nor U11506 (N_11506,N_5663,N_7113);
nand U11507 (N_11507,N_6392,N_5064);
or U11508 (N_11508,N_9838,N_9325);
nor U11509 (N_11509,N_6828,N_9894);
and U11510 (N_11510,N_9416,N_7259);
or U11511 (N_11511,N_5885,N_9072);
or U11512 (N_11512,N_7760,N_6203);
nor U11513 (N_11513,N_9393,N_7258);
nand U11514 (N_11514,N_7923,N_6590);
and U11515 (N_11515,N_8390,N_7338);
xor U11516 (N_11516,N_7412,N_7960);
nor U11517 (N_11517,N_6982,N_7164);
or U11518 (N_11518,N_9683,N_5209);
nor U11519 (N_11519,N_5925,N_8210);
xnor U11520 (N_11520,N_5332,N_7804);
nand U11521 (N_11521,N_5743,N_5112);
or U11522 (N_11522,N_7205,N_9378);
and U11523 (N_11523,N_6736,N_8064);
and U11524 (N_11524,N_8864,N_7646);
nor U11525 (N_11525,N_5504,N_9255);
or U11526 (N_11526,N_8517,N_5880);
nor U11527 (N_11527,N_5908,N_8048);
xnor U11528 (N_11528,N_7522,N_9467);
nor U11529 (N_11529,N_5390,N_8351);
nor U11530 (N_11530,N_6248,N_6535);
and U11531 (N_11531,N_7968,N_5210);
xor U11532 (N_11532,N_8147,N_8039);
nand U11533 (N_11533,N_5874,N_7504);
nand U11534 (N_11534,N_9232,N_6107);
nand U11535 (N_11535,N_9005,N_5245);
xnor U11536 (N_11536,N_6349,N_9757);
nor U11537 (N_11537,N_9933,N_7398);
or U11538 (N_11538,N_8497,N_7754);
xor U11539 (N_11539,N_7847,N_7247);
and U11540 (N_11540,N_8232,N_5598);
xor U11541 (N_11541,N_9586,N_7410);
nand U11542 (N_11542,N_5087,N_8338);
and U11543 (N_11543,N_7352,N_6991);
and U11544 (N_11544,N_8099,N_6695);
or U11545 (N_11545,N_7458,N_9231);
xor U11546 (N_11546,N_6056,N_8777);
xnor U11547 (N_11547,N_8074,N_7234);
or U11548 (N_11548,N_7218,N_7131);
or U11549 (N_11549,N_6585,N_7025);
or U11550 (N_11550,N_9646,N_9743);
xnor U11551 (N_11551,N_9857,N_6702);
xor U11552 (N_11552,N_6132,N_9211);
and U11553 (N_11553,N_5051,N_6865);
or U11554 (N_11554,N_6297,N_9901);
nor U11555 (N_11555,N_7578,N_6314);
nand U11556 (N_11556,N_8095,N_9995);
xnor U11557 (N_11557,N_8447,N_9682);
or U11558 (N_11558,N_5567,N_7667);
or U11559 (N_11559,N_8255,N_8694);
nor U11560 (N_11560,N_8006,N_5177);
and U11561 (N_11561,N_9695,N_9460);
or U11562 (N_11562,N_7203,N_9916);
nand U11563 (N_11563,N_6004,N_5533);
or U11564 (N_11564,N_9891,N_9655);
xor U11565 (N_11565,N_6481,N_8822);
nand U11566 (N_11566,N_5749,N_6923);
nor U11567 (N_11567,N_6801,N_9177);
and U11568 (N_11568,N_7494,N_8071);
nand U11569 (N_11569,N_8163,N_9210);
nand U11570 (N_11570,N_6096,N_5903);
nand U11571 (N_11571,N_9519,N_9469);
nand U11572 (N_11572,N_6825,N_9511);
xnor U11573 (N_11573,N_5399,N_9471);
nor U11574 (N_11574,N_5590,N_7441);
and U11575 (N_11575,N_6917,N_6577);
and U11576 (N_11576,N_9773,N_6123);
nor U11577 (N_11577,N_6992,N_5826);
or U11578 (N_11578,N_5558,N_9907);
nor U11579 (N_11579,N_8963,N_8679);
nor U11580 (N_11580,N_6560,N_6345);
nor U11581 (N_11581,N_8499,N_6711);
or U11582 (N_11582,N_6554,N_6849);
and U11583 (N_11583,N_8633,N_8922);
and U11584 (N_11584,N_7280,N_7661);
or U11585 (N_11585,N_7958,N_9984);
xor U11586 (N_11586,N_7254,N_9534);
or U11587 (N_11587,N_5195,N_6799);
or U11588 (N_11588,N_5617,N_8841);
xnor U11589 (N_11589,N_8350,N_7036);
nor U11590 (N_11590,N_7827,N_8180);
and U11591 (N_11591,N_7895,N_8471);
or U11592 (N_11592,N_6538,N_6053);
xor U11593 (N_11593,N_6427,N_9422);
or U11594 (N_11594,N_8698,N_6653);
xor U11595 (N_11595,N_9153,N_7010);
and U11596 (N_11596,N_8874,N_8542);
nor U11597 (N_11597,N_6645,N_5413);
nand U11598 (N_11598,N_5492,N_7854);
xor U11599 (N_11599,N_6955,N_8926);
nand U11600 (N_11600,N_6685,N_8614);
nor U11601 (N_11601,N_8686,N_6748);
or U11602 (N_11602,N_9526,N_8104);
nand U11603 (N_11603,N_5572,N_5039);
nor U11604 (N_11604,N_7822,N_6377);
xor U11605 (N_11605,N_6384,N_9136);
nor U11606 (N_11606,N_7299,N_7899);
nor U11607 (N_11607,N_7536,N_8790);
or U11608 (N_11608,N_8042,N_7805);
or U11609 (N_11609,N_8695,N_6621);
nand U11610 (N_11610,N_9339,N_6486);
nor U11611 (N_11611,N_7422,N_8565);
xor U11612 (N_11612,N_6979,N_5102);
nand U11613 (N_11613,N_8378,N_5683);
xnor U11614 (N_11614,N_8023,N_6660);
or U11615 (N_11615,N_5871,N_8235);
or U11616 (N_11616,N_9337,N_7151);
or U11617 (N_11617,N_7884,N_9612);
or U11618 (N_11618,N_6471,N_6351);
nor U11619 (N_11619,N_8988,N_5577);
xor U11620 (N_11620,N_5380,N_8443);
or U11621 (N_11621,N_7982,N_9394);
xnor U11622 (N_11622,N_6295,N_5965);
or U11623 (N_11623,N_9439,N_8226);
nand U11624 (N_11624,N_5394,N_8500);
nor U11625 (N_11625,N_5324,N_9419);
and U11626 (N_11626,N_5540,N_8916);
and U11627 (N_11627,N_6665,N_9204);
and U11628 (N_11628,N_8853,N_7780);
nor U11629 (N_11629,N_5320,N_7720);
nor U11630 (N_11630,N_5786,N_6088);
or U11631 (N_11631,N_9414,N_9259);
xor U11632 (N_11632,N_6509,N_8024);
xnor U11633 (N_11633,N_5153,N_9112);
nand U11634 (N_11634,N_7898,N_8643);
xnor U11635 (N_11635,N_7842,N_8041);
or U11636 (N_11636,N_8234,N_6289);
nor U11637 (N_11637,N_9923,N_8375);
nand U11638 (N_11638,N_5249,N_5043);
xnor U11639 (N_11639,N_7529,N_9708);
xnor U11640 (N_11640,N_7199,N_5089);
nand U11641 (N_11641,N_8756,N_7971);
nand U11642 (N_11642,N_8129,N_9446);
nor U11643 (N_11643,N_6613,N_8663);
or U11644 (N_11644,N_6714,N_5867);
xor U11645 (N_11645,N_5356,N_6080);
nor U11646 (N_11646,N_7472,N_5497);
xnor U11647 (N_11647,N_6318,N_6842);
nor U11648 (N_11648,N_9015,N_6115);
nand U11649 (N_11649,N_9990,N_7552);
and U11650 (N_11650,N_7343,N_7913);
xnor U11651 (N_11651,N_8434,N_8429);
and U11652 (N_11652,N_6529,N_8837);
or U11653 (N_11653,N_6017,N_8835);
and U11654 (N_11654,N_9451,N_8433);
nand U11655 (N_11655,N_6598,N_9693);
and U11656 (N_11656,N_9640,N_6602);
nand U11657 (N_11657,N_9939,N_8739);
and U11658 (N_11658,N_8812,N_6723);
nand U11659 (N_11659,N_9531,N_5220);
and U11660 (N_11660,N_6692,N_5719);
nand U11661 (N_11661,N_5730,N_6973);
nor U11662 (N_11662,N_8599,N_5636);
or U11663 (N_11663,N_6479,N_9390);
xnor U11664 (N_11664,N_8341,N_9726);
and U11665 (N_11665,N_5124,N_8831);
and U11666 (N_11666,N_6576,N_7903);
xnor U11667 (N_11667,N_7346,N_5296);
and U11668 (N_11668,N_9209,N_9584);
xnor U11669 (N_11669,N_6343,N_8402);
nor U11670 (N_11670,N_5267,N_5442);
nor U11671 (N_11671,N_9487,N_9539);
nor U11672 (N_11672,N_8577,N_5518);
nand U11673 (N_11673,N_7793,N_9647);
nor U11674 (N_11674,N_9609,N_6106);
and U11675 (N_11675,N_5321,N_8583);
nor U11676 (N_11676,N_6761,N_5158);
nand U11677 (N_11677,N_8297,N_7513);
nand U11678 (N_11678,N_6446,N_7304);
nand U11679 (N_11679,N_5739,N_6109);
xor U11680 (N_11680,N_8414,N_7668);
and U11681 (N_11681,N_6226,N_7921);
and U11682 (N_11682,N_8781,N_6566);
or U11683 (N_11683,N_6062,N_6861);
and U11684 (N_11684,N_8242,N_6877);
and U11685 (N_11685,N_6633,N_9652);
or U11686 (N_11686,N_8270,N_6935);
nor U11687 (N_11687,N_6668,N_6850);
or U11688 (N_11688,N_7812,N_6251);
nand U11689 (N_11689,N_7427,N_7669);
nor U11690 (N_11690,N_6557,N_7912);
and U11691 (N_11691,N_8993,N_5207);
or U11692 (N_11692,N_8228,N_8611);
and U11693 (N_11693,N_8386,N_8763);
or U11694 (N_11694,N_6934,N_9034);
or U11695 (N_11695,N_6794,N_8543);
nand U11696 (N_11696,N_8030,N_9267);
xor U11697 (N_11697,N_5306,N_8224);
xnor U11698 (N_11698,N_8370,N_5486);
nand U11699 (N_11699,N_6177,N_6045);
and U11700 (N_11700,N_5900,N_6735);
nor U11701 (N_11701,N_6522,N_7302);
nor U11702 (N_11702,N_8487,N_5300);
nand U11703 (N_11703,N_9804,N_7166);
or U11704 (N_11704,N_5779,N_6359);
and U11705 (N_11705,N_6627,N_5522);
xor U11706 (N_11706,N_5597,N_5192);
or U11707 (N_11707,N_7064,N_8380);
or U11708 (N_11708,N_7753,N_9406);
or U11709 (N_11709,N_9550,N_5876);
and U11710 (N_11710,N_5701,N_9791);
nor U11711 (N_11711,N_6167,N_6594);
nor U11712 (N_11712,N_7192,N_5829);
or U11713 (N_11713,N_6833,N_9266);
xnor U11714 (N_11714,N_6567,N_8453);
or U11715 (N_11715,N_7470,N_8127);
nor U11716 (N_11716,N_9381,N_9363);
nand U11717 (N_11717,N_8737,N_8784);
nor U11718 (N_11718,N_9092,N_5262);
or U11719 (N_11719,N_7770,N_5126);
or U11720 (N_11720,N_6737,N_9872);
or U11721 (N_11721,N_7298,N_5825);
xnor U11722 (N_11722,N_6770,N_5858);
xor U11723 (N_11723,N_7201,N_7497);
nand U11724 (N_11724,N_8250,N_5934);
and U11725 (N_11725,N_5098,N_6726);
nor U11726 (N_11726,N_9277,N_7507);
or U11727 (N_11727,N_5629,N_5604);
xor U11728 (N_11728,N_9950,N_9196);
nand U11729 (N_11729,N_6596,N_8552);
and U11730 (N_11730,N_9162,N_8323);
nor U11731 (N_11731,N_7979,N_9993);
or U11732 (N_11732,N_6231,N_7764);
xor U11733 (N_11733,N_6707,N_8114);
xnor U11734 (N_11734,N_7894,N_9965);
nand U11735 (N_11735,N_6437,N_6644);
and U11736 (N_11736,N_8389,N_7326);
and U11737 (N_11737,N_8627,N_6659);
or U11738 (N_11738,N_7236,N_6320);
nor U11739 (N_11739,N_8440,N_9080);
and U11740 (N_11740,N_8409,N_9155);
and U11741 (N_11741,N_5194,N_9296);
and U11742 (N_11742,N_7883,N_6742);
xor U11743 (N_11743,N_9349,N_6327);
xor U11744 (N_11744,N_5800,N_5405);
nand U11745 (N_11745,N_5378,N_6265);
or U11746 (N_11746,N_6378,N_9554);
nand U11747 (N_11747,N_7125,N_8212);
or U11748 (N_11748,N_6216,N_6036);
nor U11749 (N_11749,N_5499,N_5548);
nand U11750 (N_11750,N_8072,N_8329);
nor U11751 (N_11751,N_8545,N_9461);
or U11752 (N_11752,N_6068,N_6875);
or U11753 (N_11753,N_9173,N_5512);
nor U11754 (N_11754,N_6503,N_8112);
and U11755 (N_11755,N_9989,N_8312);
nor U11756 (N_11756,N_6482,N_7189);
xor U11757 (N_11757,N_8600,N_9000);
nand U11758 (N_11758,N_5811,N_7916);
or U11759 (N_11759,N_7517,N_5029);
and U11760 (N_11760,N_8526,N_8488);
nor U11761 (N_11761,N_7565,N_8182);
and U11762 (N_11762,N_5302,N_9563);
xnor U11763 (N_11763,N_6122,N_6039);
nand U11764 (N_11764,N_6671,N_7863);
xnor U11765 (N_11765,N_7709,N_9323);
xnor U11766 (N_11766,N_9994,N_7654);
nand U11767 (N_11767,N_7694,N_6139);
nand U11768 (N_11768,N_5785,N_5149);
nand U11769 (N_11769,N_8372,N_9800);
or U11770 (N_11770,N_6173,N_8786);
or U11771 (N_11771,N_9666,N_7601);
nand U11772 (N_11772,N_7232,N_7910);
and U11773 (N_11773,N_7027,N_9297);
nor U11774 (N_11774,N_5949,N_8608);
nor U11775 (N_11775,N_6263,N_7431);
or U11776 (N_11776,N_8587,N_9928);
xnor U11777 (N_11777,N_5791,N_9522);
nand U11778 (N_11778,N_9882,N_6458);
xnor U11779 (N_11779,N_7572,N_8477);
or U11780 (N_11780,N_6950,N_5053);
or U11781 (N_11781,N_9826,N_6963);
or U11782 (N_11782,N_6262,N_6930);
nand U11783 (N_11783,N_6906,N_7905);
nand U11784 (N_11784,N_5331,N_8624);
nor U11785 (N_11785,N_8518,N_9680);
xnor U11786 (N_11786,N_7204,N_8274);
and U11787 (N_11787,N_8038,N_8157);
and U11788 (N_11788,N_5263,N_9188);
nor U11789 (N_11789,N_7263,N_9662);
xnor U11790 (N_11790,N_9023,N_6476);
or U11791 (N_11791,N_9025,N_7756);
and U11792 (N_11792,N_8461,N_7816);
and U11793 (N_11793,N_9639,N_5318);
or U11794 (N_11794,N_5119,N_5654);
nand U11795 (N_11795,N_5799,N_9777);
nor U11796 (N_11796,N_5383,N_8931);
nand U11797 (N_11797,N_9016,N_9213);
nand U11798 (N_11798,N_8740,N_8966);
xnor U11799 (N_11799,N_9230,N_9156);
nand U11800 (N_11800,N_6781,N_8421);
nor U11801 (N_11801,N_8844,N_9243);
or U11802 (N_11802,N_7242,N_6895);
nor U11803 (N_11803,N_8946,N_8980);
nor U11804 (N_11804,N_5723,N_6523);
or U11805 (N_11805,N_8342,N_6072);
nand U11806 (N_11806,N_7952,N_7972);
nand U11807 (N_11807,N_7775,N_7368);
or U11808 (N_11808,N_9234,N_6317);
and U11809 (N_11809,N_7616,N_8969);
nand U11810 (N_11810,N_5772,N_9207);
nand U11811 (N_11811,N_8909,N_9582);
nand U11812 (N_11812,N_9351,N_7095);
xor U11813 (N_11813,N_6880,N_7864);
or U11814 (N_11814,N_7437,N_8345);
xor U11815 (N_11815,N_9463,N_7796);
or U11816 (N_11816,N_5807,N_5758);
nor U11817 (N_11817,N_7741,N_9395);
xor U11818 (N_11818,N_6807,N_5452);
and U11819 (N_11819,N_9046,N_8981);
xnor U11820 (N_11820,N_5011,N_7022);
nand U11821 (N_11821,N_8525,N_9405);
and U11822 (N_11822,N_5326,N_9700);
nand U11823 (N_11823,N_7035,N_6739);
or U11824 (N_11824,N_8773,N_8301);
xor U11825 (N_11825,N_9590,N_9630);
nor U11826 (N_11826,N_6753,N_8890);
xnor U11827 (N_11827,N_7510,N_7466);
and U11828 (N_11828,N_7549,N_9319);
xnor U11829 (N_11829,N_8521,N_8132);
nor U11830 (N_11830,N_5038,N_5836);
and U11831 (N_11831,N_5366,N_9280);
xor U11832 (N_11832,N_5817,N_5172);
nor U11833 (N_11833,N_6970,N_8019);
or U11834 (N_11834,N_6312,N_6241);
nor U11835 (N_11835,N_7570,N_6546);
and U11836 (N_11836,N_8282,N_9979);
nor U11837 (N_11837,N_7558,N_9686);
nor U11838 (N_11838,N_8800,N_5822);
nand U11839 (N_11839,N_8278,N_9276);
or U11840 (N_11840,N_6465,N_5164);
nand U11841 (N_11841,N_7857,N_8337);
or U11842 (N_11842,N_9017,N_7056);
nand U11843 (N_11843,N_9096,N_8239);
and U11844 (N_11844,N_7161,N_5431);
nor U11845 (N_11845,N_5012,N_5122);
nand U11846 (N_11846,N_7763,N_5069);
xnor U11847 (N_11847,N_6873,N_8467);
or U11848 (N_11848,N_9031,N_6854);
xnor U11849 (N_11849,N_8238,N_5107);
nand U11850 (N_11850,N_8124,N_9546);
xor U11851 (N_11851,N_6221,N_6085);
xor U11852 (N_11852,N_7040,N_8032);
nand U11853 (N_11853,N_7015,N_6023);
nand U11854 (N_11854,N_7540,N_8324);
nor U11855 (N_11855,N_5736,N_5063);
nand U11856 (N_11856,N_7693,N_8175);
and U11857 (N_11857,N_6744,N_5894);
nor U11858 (N_11858,N_6502,N_7790);
nor U11859 (N_11859,N_6903,N_7636);
nor U11860 (N_11860,N_8617,N_7062);
and U11861 (N_11861,N_9252,N_5970);
xnor U11862 (N_11862,N_8138,N_7777);
nand U11863 (N_11863,N_8118,N_9827);
or U11864 (N_11864,N_5010,N_9801);
xor U11865 (N_11865,N_5187,N_9732);
and U11866 (N_11866,N_7450,N_5162);
and U11867 (N_11867,N_5493,N_7488);
or U11868 (N_11868,N_9953,N_9964);
xor U11869 (N_11869,N_7732,N_8706);
nand U11870 (N_11870,N_8687,N_9951);
nor U11871 (N_11871,N_7041,N_7724);
or U11872 (N_11872,N_6006,N_9863);
and U11873 (N_11873,N_8925,N_9792);
nand U11874 (N_11874,N_8918,N_5644);
or U11875 (N_11875,N_9240,N_8013);
nor U11876 (N_11876,N_6818,N_8233);
or U11877 (N_11877,N_7223,N_5909);
nor U11878 (N_11878,N_8801,N_8572);
or U11879 (N_11879,N_7061,N_7708);
nand U11880 (N_11880,N_6012,N_6020);
xor U11881 (N_11881,N_6222,N_8492);
nand U11882 (N_11882,N_7750,N_6182);
nand U11883 (N_11883,N_9969,N_7044);
nand U11884 (N_11884,N_5707,N_8544);
and U11885 (N_11885,N_5631,N_8891);
or U11886 (N_11886,N_8423,N_6584);
or U11887 (N_11887,N_9770,N_9588);
nor U11888 (N_11888,N_9060,N_5075);
nand U11889 (N_11889,N_9608,N_6715);
and U11890 (N_11890,N_8645,N_7176);
nor U11891 (N_11891,N_9316,N_6975);
nand U11892 (N_11892,N_6555,N_7460);
nand U11893 (N_11893,N_9548,N_9903);
nor U11894 (N_11894,N_9193,N_6028);
nor U11895 (N_11895,N_8948,N_9181);
nand U11896 (N_11896,N_5443,N_7547);
nor U11897 (N_11897,N_5290,N_9618);
xnor U11898 (N_11898,N_8878,N_6029);
nor U11899 (N_11899,N_9516,N_6989);
nor U11900 (N_11900,N_8195,N_5943);
xnor U11901 (N_11901,N_6988,N_5870);
or U11902 (N_11902,N_7561,N_6064);
xor U11903 (N_11903,N_6457,N_8906);
or U11904 (N_11904,N_6841,N_6882);
or U11905 (N_11905,N_5816,N_7784);
nor U11906 (N_11906,N_8725,N_7545);
nor U11907 (N_11907,N_6578,N_5981);
xor U11908 (N_11908,N_6769,N_9830);
nand U11909 (N_11909,N_7391,N_8098);
nand U11910 (N_11910,N_7307,N_5323);
nor U11911 (N_11911,N_9749,N_9932);
xor U11912 (N_11912,N_7997,N_7287);
or U11913 (N_11913,N_9374,N_7324);
or U11914 (N_11914,N_6856,N_7959);
nor U11915 (N_11915,N_5729,N_9505);
xor U11916 (N_11916,N_8179,N_8360);
xor U11917 (N_11917,N_7020,N_6624);
xnor U11918 (N_11918,N_5559,N_9291);
xnor U11919 (N_11919,N_9510,N_7617);
nand U11920 (N_11920,N_7897,N_7240);
xnor U11921 (N_11921,N_6495,N_6977);
nand U11922 (N_11922,N_7362,N_8625);
nor U11923 (N_11923,N_6030,N_5076);
and U11924 (N_11924,N_7862,N_7557);
xor U11925 (N_11925,N_6480,N_7288);
or U11926 (N_11926,N_9148,N_5408);
nor U11927 (N_11927,N_7351,N_5180);
and U11928 (N_11928,N_8466,N_8516);
nand U11929 (N_11929,N_9867,N_8220);
and U11930 (N_11930,N_5054,N_5458);
and U11931 (N_11931,N_8286,N_5733);
and U11932 (N_11932,N_7803,N_9802);
nor U11933 (N_11933,N_5711,N_7791);
xor U11934 (N_11934,N_9160,N_7690);
and U11935 (N_11935,N_6649,N_8117);
nand U11936 (N_11936,N_6121,N_8618);
and U11937 (N_11937,N_6919,N_8576);
nor U11938 (N_11938,N_8484,N_6433);
or U11939 (N_11939,N_5237,N_7610);
xor U11940 (N_11940,N_7355,N_5060);
and U11941 (N_11941,N_9836,N_5895);
nor U11942 (N_11942,N_7114,N_9318);
or U11943 (N_11943,N_6038,N_7743);
and U11944 (N_11944,N_7196,N_8854);
nand U11945 (N_11945,N_5352,N_7407);
nand U11946 (N_11946,N_9925,N_9748);
xnor U11947 (N_11947,N_5469,N_7586);
nor U11948 (N_11948,N_5037,N_5843);
xor U11949 (N_11949,N_7554,N_8762);
or U11950 (N_11950,N_6703,N_6357);
and U11951 (N_11951,N_7675,N_9706);
xnor U11952 (N_11952,N_8989,N_7493);
nand U11953 (N_11953,N_6765,N_5111);
xnor U11954 (N_11954,N_7591,N_7145);
or U11955 (N_11955,N_5068,N_6048);
nand U11956 (N_11956,N_8431,N_6949);
and U11957 (N_11957,N_9946,N_8712);
or U11958 (N_11958,N_5859,N_5830);
nor U11959 (N_11959,N_9165,N_6993);
nand U11960 (N_11960,N_6740,N_9357);
nand U11961 (N_11961,N_5143,N_8377);
xor U11962 (N_11962,N_8638,N_7656);
nor U11963 (N_11963,N_8045,N_9850);
nor U11964 (N_11964,N_6582,N_9272);
and U11965 (N_11965,N_8027,N_7316);
and U11966 (N_11966,N_6134,N_8162);
and U11967 (N_11967,N_5134,N_9298);
or U11968 (N_11968,N_9733,N_7079);
nor U11969 (N_11969,N_7469,N_8785);
nand U11970 (N_11970,N_9566,N_5471);
and U11971 (N_11971,N_7367,N_5756);
xor U11972 (N_11972,N_5833,N_9257);
or U11973 (N_11973,N_5016,N_6368);
xnor U11974 (N_11974,N_6243,N_7165);
and U11975 (N_11975,N_7347,N_7800);
or U11976 (N_11976,N_5019,N_5495);
xnor U11977 (N_11977,N_7397,N_6984);
xor U11978 (N_11978,N_6722,N_9703);
nand U11979 (N_11979,N_9825,N_9289);
nand U11980 (N_11980,N_6190,N_9480);
and U11981 (N_11981,N_8860,N_7742);
and U11982 (N_11982,N_8871,N_6070);
xnor U11983 (N_11983,N_7953,N_6675);
or U11984 (N_11984,N_5171,N_5953);
nor U11985 (N_11985,N_5984,N_9139);
or U11986 (N_11986,N_6904,N_6421);
and U11987 (N_11987,N_7735,N_9208);
xor U11988 (N_11988,N_5832,N_5113);
and U11989 (N_11989,N_7440,N_6434);
and U11990 (N_11990,N_5354,N_8511);
nand U11991 (N_11991,N_6705,N_9440);
or U11992 (N_11992,N_6826,N_8131);
and U11993 (N_11993,N_6508,N_7322);
xor U11994 (N_11994,N_7521,N_5930);
nand U11995 (N_11995,N_8755,N_8418);
and U11996 (N_11996,N_7405,N_6942);
or U11997 (N_11997,N_5077,N_8889);
nand U11998 (N_11998,N_7386,N_6269);
nor U11999 (N_11999,N_7291,N_5156);
nand U12000 (N_12000,N_9922,N_9888);
nand U12001 (N_12001,N_7393,N_9783);
xnor U12002 (N_12002,N_7946,N_7858);
xnor U12003 (N_12003,N_5881,N_8907);
nor U12004 (N_12004,N_6120,N_5411);
and U12005 (N_12005,N_7938,N_8584);
or U12006 (N_12006,N_9681,N_8507);
or U12007 (N_12007,N_7664,N_6092);
or U12008 (N_12008,N_6966,N_6810);
xnor U12009 (N_12009,N_8382,N_7274);
xor U12010 (N_12010,N_7126,N_7444);
xnor U12011 (N_12011,N_6171,N_7004);
xor U12012 (N_12012,N_9577,N_9335);
and U12013 (N_12013,N_7454,N_5734);
xor U12014 (N_12014,N_6067,N_8888);
nand U12015 (N_12015,N_6061,N_5928);
or U12016 (N_12016,N_8397,N_6373);
nand U12017 (N_12017,N_7995,N_5412);
and U12018 (N_12018,N_8156,N_9758);
nor U12019 (N_12019,N_5571,N_8655);
nor U12020 (N_12020,N_7702,N_5887);
or U12021 (N_12021,N_6713,N_6459);
and U12022 (N_12022,N_9633,N_5990);
and U12023 (N_12023,N_7991,N_7479);
xnor U12024 (N_12024,N_6968,N_5638);
or U12025 (N_12025,N_6948,N_8194);
and U12026 (N_12026,N_9317,N_7927);
nor U12027 (N_12027,N_7813,N_5564);
xnor U12028 (N_12028,N_5056,N_6909);
nand U12029 (N_12029,N_7121,N_7856);
or U12030 (N_12030,N_6116,N_8628);
nor U12031 (N_12031,N_6077,N_9454);
nand U12032 (N_12032,N_7876,N_8620);
nor U12033 (N_12033,N_6757,N_9129);
and U12034 (N_12034,N_8140,N_6953);
nand U12035 (N_12035,N_8673,N_9854);
nor U12036 (N_12036,N_7128,N_6001);
and U12037 (N_12037,N_9282,N_7267);
and U12038 (N_12038,N_6686,N_6597);
xnor U12039 (N_12039,N_9125,N_5741);
nand U12040 (N_12040,N_6142,N_5532);
or U12041 (N_12041,N_5802,N_9352);
nand U12042 (N_12042,N_5398,N_6629);
and U12043 (N_12043,N_5912,N_6662);
and U12044 (N_12044,N_5722,N_5315);
and U12045 (N_12045,N_8371,N_6718);
and U12046 (N_12046,N_9798,N_5685);
or U12047 (N_12047,N_5774,N_8002);
nor U12048 (N_12048,N_7807,N_9527);
nor U12049 (N_12049,N_9676,N_6531);
xor U12050 (N_12050,N_6274,N_5594);
and U12051 (N_12051,N_5044,N_7416);
nor U12052 (N_12052,N_8813,N_5288);
xor U12053 (N_12053,N_5587,N_6191);
or U12054 (N_12054,N_6176,N_5127);
or U12055 (N_12055,N_8782,N_7031);
nand U12056 (N_12056,N_8254,N_9494);
or U12057 (N_12057,N_6672,N_8839);
nand U12058 (N_12058,N_9712,N_6528);
and U12059 (N_12059,N_8187,N_5496);
or U12060 (N_12060,N_5637,N_9185);
nand U12061 (N_12061,N_6537,N_6358);
xnor U12062 (N_12062,N_6959,N_5596);
or U12063 (N_12063,N_9430,N_5017);
xnor U12064 (N_12064,N_5700,N_5050);
or U12065 (N_12065,N_8343,N_8770);
nor U12066 (N_12066,N_9261,N_8322);
or U12067 (N_12067,N_5893,N_9521);
or U12068 (N_12068,N_5251,N_5645);
or U12069 (N_12069,N_6868,N_7877);
or U12070 (N_12070,N_9692,N_9553);
and U12071 (N_12071,N_7134,N_7265);
nand U12072 (N_12072,N_5148,N_8569);
and U12073 (N_12073,N_8646,N_9709);
and U12074 (N_12074,N_6474,N_5841);
nor U12075 (N_12075,N_5757,N_7633);
nand U12076 (N_12076,N_7541,N_5347);
nand U12077 (N_12077,N_6536,N_7068);
nor U12078 (N_12078,N_7870,N_9978);
nor U12079 (N_12079,N_5317,N_5818);
nor U12080 (N_12080,N_9976,N_7053);
and U12081 (N_12081,N_7099,N_5640);
nor U12082 (N_12082,N_7117,N_7433);
nor U12083 (N_12083,N_9143,N_7588);
nand U12084 (N_12084,N_8481,N_5624);
nand U12085 (N_12085,N_9048,N_9750);
xor U12086 (N_12086,N_5265,N_5099);
or U12087 (N_12087,N_9382,N_8845);
xnor U12088 (N_12088,N_5032,N_7850);
nor U12089 (N_12089,N_9293,N_8103);
xnor U12090 (N_12090,N_7399,N_8394);
or U12091 (N_12091,N_6124,N_8678);
nor U12092 (N_12092,N_7955,N_9632);
nand U12093 (N_12093,N_5650,N_8280);
nand U12094 (N_12094,N_7171,N_7471);
and U12095 (N_12095,N_7837,N_6050);
and U12096 (N_12096,N_9336,N_8034);
nand U12097 (N_12097,N_8929,N_5847);
xor U12098 (N_12098,N_8456,N_8685);
and U12099 (N_12099,N_7017,N_9528);
or U12100 (N_12100,N_7447,N_7603);
nand U12101 (N_12101,N_9099,N_6069);
xnor U12102 (N_12102,N_9157,N_9579);
nor U12103 (N_12103,N_5298,N_6789);
nor U12104 (N_12104,N_6475,N_6189);
and U12105 (N_12105,N_9024,N_8967);
nand U12106 (N_12106,N_8083,N_7867);
nor U12107 (N_12107,N_5608,N_8449);
nand U12108 (N_12108,N_5483,N_6287);
and U12109 (N_12109,N_8947,N_7500);
and U12110 (N_12110,N_6461,N_6677);
or U12111 (N_12111,N_6730,N_5977);
xnor U12112 (N_12112,N_8452,N_7188);
or U12113 (N_12113,N_8281,N_9083);
nor U12114 (N_12114,N_9093,N_6076);
nor U12115 (N_12115,N_8188,N_8408);
nor U12116 (N_12116,N_7786,N_6608);
xor U12117 (N_12117,N_9281,N_7160);
nand U12118 (N_12118,N_5524,N_5715);
nand U12119 (N_12119,N_9944,N_8726);
or U12120 (N_12120,N_8268,N_7361);
xnor U12121 (N_12121,N_5705,N_8858);
and U12122 (N_12122,N_7184,N_5333);
and U12123 (N_12123,N_7589,N_7014);
and U12124 (N_12124,N_7925,N_7665);
nand U12125 (N_12125,N_8519,N_6224);
xor U12126 (N_12126,N_7248,N_5966);
and U12127 (N_12127,N_8247,N_8742);
xor U12128 (N_12128,N_5519,N_5728);
and U12129 (N_12129,N_9870,N_9570);
and U12130 (N_12130,N_6310,N_9762);
and U12131 (N_12131,N_6830,N_7423);
nor U12132 (N_12132,N_5516,N_6803);
or U12133 (N_12133,N_7365,N_5550);
or U12134 (N_12134,N_8968,N_5178);
nand U12135 (N_12135,N_5589,N_8111);
xnor U12136 (N_12136,N_6570,N_6741);
nand U12137 (N_12137,N_8353,N_8824);
xor U12138 (N_12138,N_7584,N_5246);
and U12139 (N_12139,N_6947,N_7886);
xor U12140 (N_12140,N_6212,N_9105);
and U12141 (N_12141,N_7792,N_7571);
xor U12142 (N_12142,N_8097,N_6426);
or U12143 (N_12143,N_7644,N_8939);
nand U12144 (N_12144,N_9379,N_9664);
nor U12145 (N_12145,N_7337,N_6390);
nor U12146 (N_12146,N_5357,N_5985);
nor U12147 (N_12147,N_5174,N_7939);
and U12148 (N_12148,N_9595,N_9056);
xor U12149 (N_12149,N_9215,N_8964);
xnor U12150 (N_12150,N_8306,N_8793);
nor U12151 (N_12151,N_5448,N_6511);
xnor U12152 (N_12152,N_9671,N_7808);
xor U12153 (N_12153,N_5014,N_6900);
and U12154 (N_12154,N_5197,N_5607);
nand U12155 (N_12155,N_6802,N_6515);
nor U12156 (N_12156,N_8227,N_6628);
or U12157 (N_12157,N_8515,N_7548);
nor U12158 (N_12158,N_5367,N_6940);
and U12159 (N_12159,N_6532,N_9737);
xor U12160 (N_12160,N_8721,N_9603);
nor U12161 (N_12161,N_5080,N_8478);
nor U12162 (N_12162,N_7776,N_6864);
nor U12163 (N_12163,N_9512,N_9601);
xor U12164 (N_12164,N_9593,N_5478);
and U12165 (N_12165,N_5464,N_7116);
or U12166 (N_12166,N_7706,N_9305);
and U12167 (N_12167,N_9360,N_7384);
or U12168 (N_12168,N_7487,N_6331);
or U12169 (N_12169,N_7225,N_6687);
and U12170 (N_12170,N_8279,N_6245);
or U12171 (N_12171,N_5961,N_6416);
and U12172 (N_12172,N_8479,N_5975);
and U12173 (N_12173,N_9648,N_8613);
nand U12174 (N_12174,N_9832,N_5167);
nand U12175 (N_12175,N_6905,N_5409);
xor U12176 (N_12176,N_5510,N_6402);
or U12177 (N_12177,N_7435,N_9541);
and U12178 (N_12178,N_9287,N_6997);
nor U12179 (N_12179,N_7394,N_9062);
or U12180 (N_12180,N_9575,N_8052);
or U12181 (N_12181,N_8504,N_8910);
xor U12182 (N_12182,N_9026,N_7887);
nand U12183 (N_12183,N_5593,N_6738);
or U12184 (N_12184,N_7659,N_5745);
nand U12185 (N_12185,N_9387,N_5732);
and U12186 (N_12186,N_6867,N_5628);
xnor U12187 (N_12187,N_7491,N_8430);
and U12188 (N_12188,N_9078,N_7323);
nor U12189 (N_12189,N_8347,N_5773);
or U12190 (N_12190,N_9385,N_5301);
xor U12191 (N_12191,N_9490,N_9730);
nand U12192 (N_12192,N_8186,N_6565);
nor U12193 (N_12193,N_6309,N_9442);
nand U12194 (N_12194,N_9767,N_5582);
nand U12195 (N_12195,N_6574,N_9910);
xor U12196 (N_12196,N_8049,N_8251);
xnor U12197 (N_12197,N_8938,N_8276);
nor U12198 (N_12198,N_9966,N_5026);
and U12199 (N_12199,N_5889,N_8078);
and U12200 (N_12200,N_6379,N_9501);
xor U12201 (N_12201,N_5304,N_9285);
nand U12202 (N_12202,N_6762,N_7932);
xor U12203 (N_12203,N_5088,N_5916);
nand U12204 (N_12204,N_6143,N_6820);
or U12205 (N_12205,N_6771,N_9556);
or U12206 (N_12206,N_9010,N_8151);
or U12207 (N_12207,N_7179,N_6229);
nand U12208 (N_12208,N_5648,N_5546);
nand U12209 (N_12209,N_9626,N_7178);
nor U12210 (N_12210,N_7074,N_7744);
or U12211 (N_12211,N_6054,N_9224);
or U12212 (N_12212,N_5892,N_5656);
and U12213 (N_12213,N_9998,N_6430);
nor U12214 (N_12214,N_9779,N_8592);
or U12215 (N_12215,N_5917,N_9705);
or U12216 (N_12216,N_7911,N_5253);
nor U12217 (N_12217,N_9205,N_9476);
and U12218 (N_12218,N_8836,N_8325);
xor U12219 (N_12219,N_7019,N_8464);
or U12220 (N_12220,N_7305,N_9389);
nor U12221 (N_12221,N_5935,N_7606);
nand U12222 (N_12222,N_8851,N_9077);
or U12223 (N_12223,N_9295,N_9613);
xor U12224 (N_12224,N_9747,N_5783);
xor U12225 (N_12225,N_7629,N_5294);
nor U12226 (N_12226,N_8217,N_8096);
or U12227 (N_12227,N_9104,N_5070);
xnor U12228 (N_12228,N_9615,N_5232);
nand U12229 (N_12229,N_8568,N_5978);
and U12230 (N_12230,N_6395,N_5416);
xnor U12231 (N_12231,N_9716,N_8134);
or U12232 (N_12232,N_8881,N_8882);
and U12233 (N_12233,N_8884,N_8821);
and U12234 (N_12234,N_8553,N_6024);
nand U12235 (N_12235,N_6611,N_8648);
or U12236 (N_12236,N_6146,N_8211);
nor U12237 (N_12237,N_5272,N_6034);
and U12238 (N_12238,N_7977,N_5453);
nand U12239 (N_12239,N_7802,N_6355);
and U12240 (N_12240,N_8957,N_8626);
nand U12241 (N_12241,N_7978,N_9326);
nor U12242 (N_12242,N_7275,N_7698);
nor U12243 (N_12243,N_6009,N_7527);
nor U12244 (N_12244,N_8930,N_7907);
and U12245 (N_12245,N_6681,N_8730);
or U12246 (N_12246,N_6996,N_8815);
nor U12247 (N_12247,N_8055,N_7499);
and U12248 (N_12248,N_9359,N_8849);
nor U12249 (N_12249,N_9340,N_5030);
and U12250 (N_12250,N_7752,N_8530);
nor U12251 (N_12251,N_7483,N_5116);
xnor U12252 (N_12252,N_9263,N_5661);
and U12253 (N_12253,N_5852,N_8262);
and U12254 (N_12254,N_9936,N_9904);
or U12255 (N_12255,N_6306,N_5911);
xnor U12256 (N_12256,N_5714,N_9962);
nand U12257 (N_12257,N_7490,N_7350);
and U12258 (N_12258,N_5103,N_6406);
and U12259 (N_12259,N_6431,N_6354);
nor U12260 (N_12260,N_5789,N_7915);
nand U12261 (N_12261,N_5813,N_9817);
nor U12262 (N_12262,N_5689,N_7104);
nand U12263 (N_12263,N_8692,N_9967);
nand U12264 (N_12264,N_7378,N_6371);
nor U12265 (N_12265,N_7093,N_5284);
xor U12266 (N_12266,N_7333,N_5886);
nand U12267 (N_12267,N_8958,N_9169);
xnor U12268 (N_12268,N_7468,N_7987);
and U12269 (N_12269,N_9970,N_5230);
or U12270 (N_12270,N_7688,N_6924);
or U12271 (N_12271,N_8550,N_8020);
xor U12272 (N_12272,N_5523,N_8058);
or U12273 (N_12273,N_9581,N_6680);
nor U12274 (N_12274,N_6100,N_6372);
or U12275 (N_12275,N_8684,N_9930);
xnor U12276 (N_12276,N_8496,N_5234);
nand U12277 (N_12277,N_5983,N_8738);
and U12278 (N_12278,N_8690,N_7643);
or U12279 (N_12279,N_9199,N_5944);
or U12280 (N_12280,N_5806,N_5989);
and U12281 (N_12281,N_9391,N_6311);
and U12282 (N_12282,N_5110,N_6008);
xnor U12283 (N_12283,N_6811,N_9042);
or U12284 (N_12284,N_7107,N_9334);
nand U12285 (N_12285,N_8867,N_6326);
or U12286 (N_12286,N_5430,N_8462);
nand U12287 (N_12287,N_8647,N_5821);
nand U12288 (N_12288,N_9606,N_9637);
xnor U12289 (N_12289,N_8973,N_9636);
nand U12290 (N_12290,N_7951,N_5520);
nand U12291 (N_12291,N_8031,N_5438);
nor U12292 (N_12292,N_7016,N_6734);
or U12293 (N_12293,N_5472,N_6829);
and U12294 (N_12294,N_9262,N_8677);
or U12295 (N_12295,N_6259,N_6823);
nand U12296 (N_12296,N_5303,N_5551);
nor U12297 (N_12297,N_8173,N_5428);
or U12298 (N_12298,N_8463,N_6456);
nand U12299 (N_12299,N_6785,N_9020);
xnor U12300 (N_12300,N_7631,N_5073);
or U12301 (N_12301,N_7303,N_9229);
nor U12302 (N_12302,N_7206,N_7009);
nand U12303 (N_12303,N_8688,N_8689);
nor U12304 (N_12304,N_5461,N_5573);
nor U12305 (N_12305,N_7909,N_6141);
nand U12306 (N_12306,N_6464,N_8107);
nor U12307 (N_12307,N_5035,N_6852);
nor U12308 (N_12308,N_8152,N_7873);
nand U12309 (N_12309,N_8063,N_9186);
nand U12310 (N_12310,N_8016,N_9401);
or U12311 (N_12311,N_7769,N_6235);
nand U12312 (N_12312,N_6227,N_8998);
nor U12313 (N_12313,N_7328,N_5036);
nor U12314 (N_12314,N_8696,N_5744);
or U12315 (N_12315,N_5996,N_8736);
xor U12316 (N_12316,N_5706,N_7918);
nor U12317 (N_12317,N_7414,N_8455);
and U12318 (N_12318,N_8711,N_5433);
or U12319 (N_12319,N_9428,N_5735);
nor U12320 (N_12320,N_6782,N_6733);
nand U12321 (N_12321,N_8593,N_6168);
nor U12322 (N_12322,N_8581,N_9313);
and U12323 (N_12323,N_8015,N_7963);
xnor U12324 (N_12324,N_8590,N_9320);
xnor U12325 (N_12325,N_7300,N_8995);
or U12326 (N_12326,N_6204,N_8352);
or U12327 (N_12327,N_5402,N_8364);
nand U12328 (N_12328,N_8699,N_5574);
or U12329 (N_12329,N_6488,N_9876);
and U12330 (N_12330,N_9127,N_8460);
or U12331 (N_12331,N_6860,N_8011);
nor U12332 (N_12332,N_8000,N_5738);
nand U12333 (N_12333,N_5083,N_7137);
nand U12334 (N_12334,N_6470,N_5820);
nand U12335 (N_12335,N_7451,N_5998);
nor U12336 (N_12336,N_6915,N_6275);
or U12337 (N_12337,N_8977,N_8470);
nand U12338 (N_12338,N_8457,N_8808);
xnor U12339 (N_12339,N_6958,N_8295);
and U12340 (N_12340,N_9247,N_8033);
nor U12341 (N_12341,N_5481,N_5406);
nor U12342 (N_12342,N_8051,N_7999);
nand U12343 (N_12343,N_6140,N_6261);
nand U12344 (N_12344,N_6192,N_6186);
or U12345 (N_12345,N_9362,N_5350);
nor U12346 (N_12346,N_6599,N_7917);
xnor U12347 (N_12347,N_8707,N_5020);
nor U12348 (N_12348,N_6520,N_8475);
xor U12349 (N_12349,N_9371,N_6155);
xnor U12350 (N_12350,N_5299,N_9300);
or U12351 (N_12351,N_6174,N_6294);
xnor U12352 (N_12352,N_7395,N_6595);
nor U12353 (N_12353,N_7183,N_6441);
xor U12354 (N_12354,N_6161,N_7282);
or U12355 (N_12355,N_5612,N_6150);
or U12356 (N_12356,N_6233,N_5595);
nand U12357 (N_12357,N_7582,N_5684);
nand U12358 (N_12358,N_7482,N_9377);
nand U12359 (N_12359,N_7182,N_9492);
or U12360 (N_12360,N_8405,N_8231);
xor U12361 (N_12361,N_7799,N_9578);
or U12362 (N_12362,N_9880,N_9544);
or U12363 (N_12363,N_9014,N_7135);
or U12364 (N_12364,N_8764,N_7156);
and U12365 (N_12365,N_7231,N_8533);
xnor U12366 (N_12366,N_9814,N_8604);
nor U12367 (N_12367,N_6266,N_7417);
xor U12368 (N_12368,N_5219,N_6656);
xor U12369 (N_12369,N_8094,N_8183);
nor U12370 (N_12370,N_5420,N_5660);
nor U12371 (N_12371,N_7531,N_8252);
nand U12372 (N_12372,N_6336,N_9392);
and U12373 (N_12373,N_8401,N_6196);
and U12374 (N_12374,N_6256,N_5145);
and U12375 (N_12375,N_9542,N_9530);
or U12376 (N_12376,N_6428,N_5872);
or U12377 (N_12377,N_9958,N_5762);
nand U12378 (N_12378,N_6784,N_8621);
nor U12379 (N_12379,N_8549,N_9878);
nor U12380 (N_12380,N_8741,N_8275);
xor U12381 (N_12381,N_9484,N_9003);
and U12382 (N_12382,N_9376,N_9302);
xnor U12383 (N_12383,N_7559,N_5539);
nand U12384 (N_12384,N_6094,N_5963);
nand U12385 (N_12385,N_8990,N_7127);
xor U12386 (N_12386,N_7281,N_6131);
or U12387 (N_12387,N_6381,N_6521);
and U12388 (N_12388,N_5470,N_9670);
nor U12389 (N_12389,N_5610,N_8393);
nand U12390 (N_12390,N_9001,N_7434);
xnor U12391 (N_12391,N_7402,N_7713);
and U12392 (N_12392,N_6490,N_9082);
xnor U12393 (N_12393,N_9135,N_9306);
nor U12394 (N_12394,N_8619,N_5541);
nand U12395 (N_12395,N_5542,N_5007);
nand U12396 (N_12396,N_8752,N_9115);
and U12397 (N_12397,N_9520,N_6657);
nand U12398 (N_12398,N_8817,N_9445);
xor U12399 (N_12399,N_9070,N_9865);
or U12400 (N_12400,N_9947,N_6425);
or U12401 (N_12401,N_8940,N_9258);
nor U12402 (N_12402,N_7097,N_9051);
or U12403 (N_12403,N_8149,N_6497);
xor U12404 (N_12404,N_7749,N_9436);
xor U12405 (N_12405,N_8148,N_8510);
or U12406 (N_12406,N_6848,N_7002);
and U12407 (N_12407,N_5678,N_9168);
or U12408 (N_12408,N_5795,N_5396);
nor U12409 (N_12409,N_5526,N_8788);
or U12410 (N_12410,N_6768,N_7645);
nand U12411 (N_12411,N_7848,N_6772);
xnor U12412 (N_12412,N_5292,N_8458);
xor U12413 (N_12413,N_9029,N_7045);
or U12414 (N_12414,N_8395,N_5223);
nand U12415 (N_12415,N_8485,N_5005);
and U12416 (N_12416,N_7438,N_7890);
xnor U12417 (N_12417,N_9987,N_5737);
or U12418 (N_12418,N_5105,N_7273);
nand U12419 (N_12419,N_7296,N_8221);
and U12420 (N_12420,N_9988,N_9561);
and U12421 (N_12421,N_8261,N_6725);
and U12422 (N_12422,N_5754,N_9397);
nor U12423 (N_12423,N_5992,N_5279);
nor U12424 (N_12424,N_6553,N_8142);
nand U12425 (N_12425,N_7697,N_8365);
nand U12426 (N_12426,N_9645,N_9537);
nand U12427 (N_12427,N_5387,N_6016);
and U12428 (N_12428,N_8573,N_8001);
and U12429 (N_12429,N_8442,N_5376);
nand U12430 (N_12430,N_8438,N_5421);
nor U12431 (N_12431,N_5198,N_9421);
xor U12432 (N_12432,N_7615,N_8575);
nand U12433 (N_12433,N_7607,N_5769);
nand U12434 (N_12434,N_5311,N_7000);
xor U12435 (N_12435,N_8296,N_5018);
nand U12436 (N_12436,N_9784,N_5000);
nor U12437 (N_12437,N_9840,N_8085);
and U12438 (N_12438,N_9429,N_6838);
xor U12439 (N_12439,N_5941,N_8662);
nand U12440 (N_12440,N_6620,N_9309);
nor U12441 (N_12441,N_9697,N_6353);
nor U12442 (N_12442,N_6047,N_9896);
nor U12443 (N_12443,N_5340,N_7465);
nand U12444 (N_12444,N_9807,N_5217);
and U12445 (N_12445,N_7257,N_8265);
xnor U12446 (N_12446,N_7974,N_5658);
nand U12447 (N_12447,N_7309,N_6375);
nor U12448 (N_12448,N_8594,N_6104);
xnor U12449 (N_12449,N_5849,N_8561);
nor U12450 (N_12450,N_7506,N_7129);
xnor U12451 (N_12451,N_5753,N_5768);
nor U12452 (N_12452,N_7818,N_8597);
xor U12453 (N_12453,N_6617,N_8197);
nand U12454 (N_12454,N_5679,N_5862);
nand U12455 (N_12455,N_5804,N_5381);
nor U12456 (N_12456,N_9448,N_6674);
xor U12457 (N_12457,N_9269,N_9423);
xnor U12458 (N_12458,N_7138,N_6207);
nor U12459 (N_12459,N_8089,N_5130);
nor U12460 (N_12460,N_7383,N_9940);
xor U12461 (N_12461,N_9557,N_5621);
nor U12462 (N_12462,N_5224,N_7214);
nor U12463 (N_12463,N_7647,N_7563);
nor U12464 (N_12464,N_6921,N_5699);
xor U12465 (N_12465,N_9425,N_7605);
xnor U12466 (N_12466,N_8532,N_7684);
nor U12467 (N_12467,N_6593,N_9137);
xnor U12468 (N_12468,N_7439,N_7635);
nor U12469 (N_12469,N_9120,N_6500);
xnor U12470 (N_12470,N_8855,N_7942);
or U12471 (N_12471,N_9191,N_9301);
nor U12472 (N_12472,N_7284,N_6960);
and U12473 (N_12473,N_9679,N_9937);
and U12474 (N_12474,N_6044,N_5627);
nand U12475 (N_12475,N_9795,N_6401);
and U12476 (N_12476,N_8820,N_9518);
nand U12477 (N_12477,N_9875,N_7844);
nor U12478 (N_12478,N_9571,N_7994);
xnor U12479 (N_12479,N_8563,N_6445);
nand U12480 (N_12480,N_5264,N_8701);
xnor U12481 (N_12481,N_8317,N_6201);
xnor U12482 (N_12482,N_9746,N_7429);
nor U12483 (N_12483,N_5479,N_9028);
nand U12484 (N_12484,N_5432,N_7831);
nand U12485 (N_12485,N_9540,N_6589);
xor U12486 (N_12486,N_8537,N_7681);
and U12487 (N_12487,N_5455,N_9760);
and U12488 (N_12488,N_5389,N_9862);
and U12489 (N_12489,N_7057,N_5028);
nor U12490 (N_12490,N_9388,N_5958);
nand U12491 (N_12491,N_9659,N_7100);
nand U12492 (N_12492,N_9755,N_7733);
xor U12493 (N_12493,N_7556,N_5695);
xor U12494 (N_12494,N_8905,N_8776);
and U12495 (N_12495,N_7626,N_8745);
and U12496 (N_12496,N_7672,N_9311);
or U12497 (N_12497,N_9567,N_5203);
nor U12498 (N_12498,N_9194,N_5213);
or U12499 (N_12499,N_8029,N_5169);
xor U12500 (N_12500,N_5317,N_9601);
or U12501 (N_12501,N_7804,N_5767);
or U12502 (N_12502,N_5163,N_6398);
or U12503 (N_12503,N_9634,N_9524);
and U12504 (N_12504,N_7220,N_8861);
and U12505 (N_12505,N_9572,N_9746);
xor U12506 (N_12506,N_6552,N_7449);
xor U12507 (N_12507,N_6393,N_5149);
or U12508 (N_12508,N_8714,N_8174);
and U12509 (N_12509,N_6491,N_9498);
or U12510 (N_12510,N_7908,N_6875);
and U12511 (N_12511,N_8045,N_9370);
or U12512 (N_12512,N_5068,N_9799);
and U12513 (N_12513,N_8586,N_9021);
nand U12514 (N_12514,N_7669,N_7038);
nor U12515 (N_12515,N_8079,N_9251);
or U12516 (N_12516,N_6826,N_8889);
and U12517 (N_12517,N_9515,N_6740);
xor U12518 (N_12518,N_7775,N_9436);
xor U12519 (N_12519,N_8753,N_7316);
or U12520 (N_12520,N_5891,N_6561);
and U12521 (N_12521,N_5640,N_8441);
and U12522 (N_12522,N_6632,N_7791);
nor U12523 (N_12523,N_9578,N_9124);
xor U12524 (N_12524,N_6227,N_9350);
nand U12525 (N_12525,N_9944,N_5359);
xnor U12526 (N_12526,N_5846,N_7982);
nand U12527 (N_12527,N_5580,N_8544);
nor U12528 (N_12528,N_9900,N_5094);
nor U12529 (N_12529,N_8201,N_6281);
nor U12530 (N_12530,N_5777,N_6437);
and U12531 (N_12531,N_9434,N_6046);
or U12532 (N_12532,N_8430,N_9554);
nand U12533 (N_12533,N_8293,N_5200);
or U12534 (N_12534,N_6476,N_7356);
nand U12535 (N_12535,N_8895,N_7055);
nand U12536 (N_12536,N_8578,N_9035);
and U12537 (N_12537,N_5819,N_5698);
nor U12538 (N_12538,N_9226,N_9865);
or U12539 (N_12539,N_7025,N_7692);
or U12540 (N_12540,N_8135,N_6889);
and U12541 (N_12541,N_8487,N_8898);
nor U12542 (N_12542,N_9830,N_8991);
nand U12543 (N_12543,N_6929,N_8187);
or U12544 (N_12544,N_8082,N_6125);
or U12545 (N_12545,N_9091,N_8081);
nor U12546 (N_12546,N_5130,N_9524);
xor U12547 (N_12547,N_5587,N_6928);
xnor U12548 (N_12548,N_6938,N_6604);
xnor U12549 (N_12549,N_6852,N_5552);
and U12550 (N_12550,N_6554,N_7101);
xnor U12551 (N_12551,N_8276,N_8226);
xnor U12552 (N_12552,N_9077,N_9377);
nor U12553 (N_12553,N_7039,N_6223);
nand U12554 (N_12554,N_5010,N_5300);
and U12555 (N_12555,N_7229,N_8107);
nand U12556 (N_12556,N_6962,N_9289);
nor U12557 (N_12557,N_8515,N_7648);
nand U12558 (N_12558,N_9444,N_5040);
and U12559 (N_12559,N_9729,N_9861);
or U12560 (N_12560,N_8553,N_9102);
or U12561 (N_12561,N_7756,N_8641);
and U12562 (N_12562,N_6328,N_8222);
nand U12563 (N_12563,N_6931,N_9685);
or U12564 (N_12564,N_8431,N_8205);
nor U12565 (N_12565,N_6116,N_6261);
or U12566 (N_12566,N_8853,N_9790);
and U12567 (N_12567,N_9300,N_5914);
nand U12568 (N_12568,N_5980,N_7833);
and U12569 (N_12569,N_7880,N_6283);
nor U12570 (N_12570,N_5752,N_8289);
xor U12571 (N_12571,N_8325,N_9539);
nor U12572 (N_12572,N_9578,N_6246);
or U12573 (N_12573,N_9646,N_9192);
xor U12574 (N_12574,N_6270,N_9921);
nor U12575 (N_12575,N_7961,N_5531);
nand U12576 (N_12576,N_6923,N_9468);
xnor U12577 (N_12577,N_7494,N_8072);
nor U12578 (N_12578,N_5502,N_6610);
nor U12579 (N_12579,N_8133,N_6958);
nand U12580 (N_12580,N_7909,N_5025);
or U12581 (N_12581,N_5424,N_6670);
or U12582 (N_12582,N_5120,N_5785);
nor U12583 (N_12583,N_8275,N_9076);
and U12584 (N_12584,N_9524,N_5173);
nand U12585 (N_12585,N_8009,N_7378);
nand U12586 (N_12586,N_9332,N_6104);
and U12587 (N_12587,N_9796,N_9125);
nand U12588 (N_12588,N_8413,N_6907);
xor U12589 (N_12589,N_7693,N_5096);
and U12590 (N_12590,N_7216,N_8375);
or U12591 (N_12591,N_5065,N_8475);
xor U12592 (N_12592,N_9252,N_7095);
or U12593 (N_12593,N_5036,N_7266);
xnor U12594 (N_12594,N_9731,N_5353);
nand U12595 (N_12595,N_8781,N_9227);
nand U12596 (N_12596,N_6827,N_7796);
xnor U12597 (N_12597,N_9936,N_9125);
and U12598 (N_12598,N_9035,N_6891);
nand U12599 (N_12599,N_9693,N_5721);
nor U12600 (N_12600,N_5690,N_5938);
and U12601 (N_12601,N_7387,N_5431);
or U12602 (N_12602,N_9702,N_6524);
xnor U12603 (N_12603,N_8184,N_9517);
or U12604 (N_12604,N_5442,N_5578);
or U12605 (N_12605,N_6781,N_7568);
or U12606 (N_12606,N_8797,N_7442);
xnor U12607 (N_12607,N_6395,N_8065);
nand U12608 (N_12608,N_5434,N_5473);
nor U12609 (N_12609,N_7142,N_6512);
or U12610 (N_12610,N_8271,N_9071);
nor U12611 (N_12611,N_9375,N_8242);
nand U12612 (N_12612,N_6097,N_6181);
xor U12613 (N_12613,N_5999,N_6999);
and U12614 (N_12614,N_5278,N_8803);
or U12615 (N_12615,N_8688,N_7859);
or U12616 (N_12616,N_9262,N_6923);
xor U12617 (N_12617,N_8507,N_9662);
nor U12618 (N_12618,N_6039,N_8849);
nand U12619 (N_12619,N_5620,N_6792);
or U12620 (N_12620,N_8486,N_8627);
nand U12621 (N_12621,N_5747,N_5066);
nand U12622 (N_12622,N_5489,N_6975);
and U12623 (N_12623,N_5918,N_9147);
xor U12624 (N_12624,N_8998,N_9100);
nor U12625 (N_12625,N_7236,N_6117);
nor U12626 (N_12626,N_5391,N_6017);
or U12627 (N_12627,N_5190,N_7342);
and U12628 (N_12628,N_6354,N_6443);
xnor U12629 (N_12629,N_6248,N_8861);
or U12630 (N_12630,N_5237,N_8935);
or U12631 (N_12631,N_6868,N_8911);
xor U12632 (N_12632,N_6998,N_8988);
nor U12633 (N_12633,N_7828,N_8877);
and U12634 (N_12634,N_9064,N_6546);
nor U12635 (N_12635,N_8504,N_6285);
nor U12636 (N_12636,N_6949,N_8574);
xnor U12637 (N_12637,N_5726,N_8627);
and U12638 (N_12638,N_5877,N_9536);
and U12639 (N_12639,N_7311,N_7050);
nand U12640 (N_12640,N_9977,N_6620);
and U12641 (N_12641,N_8310,N_8661);
nor U12642 (N_12642,N_8606,N_5172);
or U12643 (N_12643,N_5715,N_5097);
nor U12644 (N_12644,N_7443,N_7353);
nor U12645 (N_12645,N_7674,N_8917);
nor U12646 (N_12646,N_6882,N_9856);
and U12647 (N_12647,N_5991,N_9398);
nand U12648 (N_12648,N_6297,N_7078);
and U12649 (N_12649,N_9590,N_9749);
nor U12650 (N_12650,N_5872,N_7775);
xnor U12651 (N_12651,N_6545,N_5152);
and U12652 (N_12652,N_9564,N_5165);
xnor U12653 (N_12653,N_6336,N_6290);
nand U12654 (N_12654,N_7838,N_8423);
or U12655 (N_12655,N_7232,N_7854);
or U12656 (N_12656,N_9631,N_7528);
nor U12657 (N_12657,N_6452,N_5512);
xor U12658 (N_12658,N_8628,N_7090);
or U12659 (N_12659,N_8384,N_5960);
and U12660 (N_12660,N_5047,N_7384);
xnor U12661 (N_12661,N_5350,N_9586);
nor U12662 (N_12662,N_5685,N_5942);
nor U12663 (N_12663,N_5127,N_5654);
nor U12664 (N_12664,N_5818,N_5079);
xor U12665 (N_12665,N_8695,N_6685);
or U12666 (N_12666,N_8828,N_8940);
nand U12667 (N_12667,N_8547,N_7146);
nand U12668 (N_12668,N_6962,N_6145);
nand U12669 (N_12669,N_9445,N_7717);
nor U12670 (N_12670,N_7960,N_8227);
nor U12671 (N_12671,N_7700,N_9565);
or U12672 (N_12672,N_9978,N_8834);
nor U12673 (N_12673,N_6964,N_8128);
nor U12674 (N_12674,N_9803,N_9902);
xnor U12675 (N_12675,N_7320,N_8166);
nor U12676 (N_12676,N_8388,N_9672);
and U12677 (N_12677,N_6154,N_9065);
nor U12678 (N_12678,N_5104,N_5609);
or U12679 (N_12679,N_7098,N_6806);
nor U12680 (N_12680,N_7706,N_5935);
xor U12681 (N_12681,N_9557,N_6069);
nand U12682 (N_12682,N_7618,N_5079);
nand U12683 (N_12683,N_6537,N_5652);
and U12684 (N_12684,N_8683,N_8311);
nand U12685 (N_12685,N_8437,N_8794);
and U12686 (N_12686,N_9718,N_8989);
xnor U12687 (N_12687,N_7655,N_6325);
nand U12688 (N_12688,N_5105,N_5164);
nor U12689 (N_12689,N_9970,N_8353);
nor U12690 (N_12690,N_6305,N_5033);
xor U12691 (N_12691,N_6318,N_6896);
or U12692 (N_12692,N_8254,N_6826);
or U12693 (N_12693,N_9891,N_9773);
and U12694 (N_12694,N_7453,N_9561);
nor U12695 (N_12695,N_6123,N_5847);
xnor U12696 (N_12696,N_5578,N_8971);
nand U12697 (N_12697,N_8992,N_8475);
xnor U12698 (N_12698,N_5543,N_6961);
or U12699 (N_12699,N_5520,N_5400);
or U12700 (N_12700,N_7087,N_8522);
or U12701 (N_12701,N_7119,N_9836);
nor U12702 (N_12702,N_7011,N_8123);
and U12703 (N_12703,N_8369,N_7820);
or U12704 (N_12704,N_9292,N_7250);
nand U12705 (N_12705,N_7735,N_8896);
nand U12706 (N_12706,N_9814,N_7251);
or U12707 (N_12707,N_5820,N_7568);
xor U12708 (N_12708,N_5625,N_6218);
xnor U12709 (N_12709,N_9683,N_5278);
and U12710 (N_12710,N_6946,N_8069);
xor U12711 (N_12711,N_9621,N_9480);
nor U12712 (N_12712,N_6315,N_5101);
nand U12713 (N_12713,N_7845,N_8171);
and U12714 (N_12714,N_5688,N_6270);
or U12715 (N_12715,N_7910,N_7779);
nand U12716 (N_12716,N_6674,N_7372);
or U12717 (N_12717,N_7182,N_9620);
or U12718 (N_12718,N_8596,N_9958);
or U12719 (N_12719,N_9970,N_9879);
or U12720 (N_12720,N_6390,N_8953);
nor U12721 (N_12721,N_5069,N_5226);
or U12722 (N_12722,N_8299,N_5683);
or U12723 (N_12723,N_7146,N_6820);
and U12724 (N_12724,N_9046,N_7642);
xor U12725 (N_12725,N_9909,N_8234);
xor U12726 (N_12726,N_6190,N_6403);
and U12727 (N_12727,N_7376,N_8701);
nor U12728 (N_12728,N_9512,N_7860);
and U12729 (N_12729,N_5675,N_9797);
or U12730 (N_12730,N_8029,N_6817);
or U12731 (N_12731,N_9201,N_8544);
nand U12732 (N_12732,N_9389,N_6958);
nor U12733 (N_12733,N_7314,N_9810);
and U12734 (N_12734,N_9617,N_5185);
xnor U12735 (N_12735,N_6824,N_5725);
nor U12736 (N_12736,N_8885,N_8875);
or U12737 (N_12737,N_6655,N_8838);
nor U12738 (N_12738,N_8753,N_7575);
xor U12739 (N_12739,N_5726,N_6742);
and U12740 (N_12740,N_7685,N_6968);
xnor U12741 (N_12741,N_9505,N_9634);
and U12742 (N_12742,N_7715,N_6309);
and U12743 (N_12743,N_7837,N_7743);
nor U12744 (N_12744,N_8157,N_7196);
xor U12745 (N_12745,N_5698,N_9708);
and U12746 (N_12746,N_5885,N_8745);
xnor U12747 (N_12747,N_8086,N_7460);
or U12748 (N_12748,N_6838,N_9836);
nor U12749 (N_12749,N_8295,N_8534);
or U12750 (N_12750,N_5307,N_8257);
nor U12751 (N_12751,N_6579,N_6507);
and U12752 (N_12752,N_7117,N_8559);
nor U12753 (N_12753,N_6350,N_5168);
nor U12754 (N_12754,N_9020,N_5934);
or U12755 (N_12755,N_7222,N_9356);
xor U12756 (N_12756,N_9059,N_6499);
or U12757 (N_12757,N_6036,N_6233);
nand U12758 (N_12758,N_5036,N_9631);
nand U12759 (N_12759,N_5717,N_9048);
xor U12760 (N_12760,N_5872,N_6959);
or U12761 (N_12761,N_8956,N_5847);
xnor U12762 (N_12762,N_9137,N_6174);
or U12763 (N_12763,N_6382,N_6867);
nor U12764 (N_12764,N_6939,N_7379);
or U12765 (N_12765,N_5236,N_9525);
nor U12766 (N_12766,N_6721,N_7179);
nor U12767 (N_12767,N_8170,N_5737);
and U12768 (N_12768,N_7811,N_9222);
xnor U12769 (N_12769,N_6003,N_8864);
and U12770 (N_12770,N_5097,N_6629);
or U12771 (N_12771,N_8684,N_5784);
or U12772 (N_12772,N_9658,N_8636);
xor U12773 (N_12773,N_5247,N_8637);
nand U12774 (N_12774,N_6194,N_8282);
nand U12775 (N_12775,N_7107,N_7267);
and U12776 (N_12776,N_8409,N_7482);
xor U12777 (N_12777,N_8406,N_6023);
xnor U12778 (N_12778,N_7539,N_8689);
and U12779 (N_12779,N_8787,N_8163);
or U12780 (N_12780,N_5392,N_9271);
nor U12781 (N_12781,N_9374,N_7733);
nor U12782 (N_12782,N_5786,N_6389);
or U12783 (N_12783,N_7113,N_5821);
nand U12784 (N_12784,N_5184,N_5982);
and U12785 (N_12785,N_8975,N_8245);
nand U12786 (N_12786,N_9428,N_6868);
xor U12787 (N_12787,N_9680,N_5755);
nor U12788 (N_12788,N_6371,N_9457);
xor U12789 (N_12789,N_7727,N_6811);
nor U12790 (N_12790,N_8785,N_9949);
nor U12791 (N_12791,N_6223,N_9632);
and U12792 (N_12792,N_9289,N_7104);
or U12793 (N_12793,N_6619,N_7743);
nor U12794 (N_12794,N_6385,N_5388);
nor U12795 (N_12795,N_5265,N_9394);
nor U12796 (N_12796,N_5868,N_5387);
and U12797 (N_12797,N_9099,N_9911);
or U12798 (N_12798,N_6002,N_7331);
xor U12799 (N_12799,N_6324,N_6323);
nor U12800 (N_12800,N_6304,N_6934);
nand U12801 (N_12801,N_9995,N_5915);
and U12802 (N_12802,N_5655,N_8811);
nor U12803 (N_12803,N_8336,N_9351);
or U12804 (N_12804,N_7006,N_8625);
nand U12805 (N_12805,N_6487,N_9417);
nor U12806 (N_12806,N_6034,N_9732);
xnor U12807 (N_12807,N_6529,N_9624);
or U12808 (N_12808,N_9620,N_6377);
xor U12809 (N_12809,N_8019,N_7113);
xor U12810 (N_12810,N_6156,N_7728);
and U12811 (N_12811,N_7711,N_7336);
or U12812 (N_12812,N_6513,N_9103);
xor U12813 (N_12813,N_9092,N_8803);
nand U12814 (N_12814,N_6894,N_6294);
nor U12815 (N_12815,N_8347,N_6890);
xnor U12816 (N_12816,N_9157,N_8607);
nand U12817 (N_12817,N_8244,N_8327);
or U12818 (N_12818,N_9017,N_5012);
or U12819 (N_12819,N_6937,N_9125);
nand U12820 (N_12820,N_7025,N_8243);
xor U12821 (N_12821,N_6426,N_9463);
or U12822 (N_12822,N_9195,N_5592);
and U12823 (N_12823,N_8011,N_7861);
or U12824 (N_12824,N_9344,N_8448);
nand U12825 (N_12825,N_6355,N_7573);
xnor U12826 (N_12826,N_9658,N_5301);
nor U12827 (N_12827,N_8306,N_5355);
xnor U12828 (N_12828,N_5428,N_8982);
nand U12829 (N_12829,N_5509,N_8160);
and U12830 (N_12830,N_6022,N_7480);
nor U12831 (N_12831,N_6430,N_5332);
and U12832 (N_12832,N_6025,N_5415);
nand U12833 (N_12833,N_7380,N_7743);
and U12834 (N_12834,N_7545,N_8894);
nand U12835 (N_12835,N_6045,N_6613);
or U12836 (N_12836,N_7253,N_5672);
xnor U12837 (N_12837,N_9524,N_7366);
or U12838 (N_12838,N_7414,N_7593);
and U12839 (N_12839,N_6389,N_5529);
or U12840 (N_12840,N_8078,N_6031);
or U12841 (N_12841,N_9282,N_9905);
xor U12842 (N_12842,N_7328,N_6208);
or U12843 (N_12843,N_8005,N_8294);
nor U12844 (N_12844,N_9739,N_8425);
nand U12845 (N_12845,N_6605,N_7452);
nand U12846 (N_12846,N_6305,N_5725);
nor U12847 (N_12847,N_9390,N_8634);
or U12848 (N_12848,N_7549,N_9592);
nand U12849 (N_12849,N_8098,N_6727);
and U12850 (N_12850,N_9708,N_7727);
or U12851 (N_12851,N_9717,N_9634);
xor U12852 (N_12852,N_5783,N_6786);
nand U12853 (N_12853,N_7964,N_6444);
or U12854 (N_12854,N_7637,N_5718);
and U12855 (N_12855,N_7960,N_5220);
nor U12856 (N_12856,N_9434,N_8910);
nand U12857 (N_12857,N_9429,N_7852);
and U12858 (N_12858,N_9266,N_8822);
xor U12859 (N_12859,N_6823,N_7466);
or U12860 (N_12860,N_7296,N_9464);
nand U12861 (N_12861,N_9322,N_5751);
nand U12862 (N_12862,N_9372,N_6403);
or U12863 (N_12863,N_8929,N_7556);
or U12864 (N_12864,N_7366,N_6849);
nand U12865 (N_12865,N_6514,N_9711);
or U12866 (N_12866,N_6202,N_5496);
and U12867 (N_12867,N_5201,N_6364);
xnor U12868 (N_12868,N_5652,N_8098);
nor U12869 (N_12869,N_9177,N_5258);
nor U12870 (N_12870,N_5321,N_5947);
nand U12871 (N_12871,N_6423,N_5289);
and U12872 (N_12872,N_6142,N_7875);
or U12873 (N_12873,N_8036,N_6043);
xnor U12874 (N_12874,N_9199,N_6105);
or U12875 (N_12875,N_5659,N_6355);
and U12876 (N_12876,N_6997,N_5823);
xnor U12877 (N_12877,N_6039,N_5713);
nor U12878 (N_12878,N_7676,N_9684);
xor U12879 (N_12879,N_6525,N_5603);
xnor U12880 (N_12880,N_6757,N_6446);
nand U12881 (N_12881,N_9214,N_7864);
nand U12882 (N_12882,N_7137,N_7184);
nand U12883 (N_12883,N_8279,N_7321);
nor U12884 (N_12884,N_8379,N_9688);
and U12885 (N_12885,N_6374,N_5673);
and U12886 (N_12886,N_5355,N_6673);
and U12887 (N_12887,N_6832,N_6036);
nand U12888 (N_12888,N_6925,N_8457);
and U12889 (N_12889,N_8776,N_8660);
nand U12890 (N_12890,N_8191,N_7680);
xor U12891 (N_12891,N_7403,N_5272);
xor U12892 (N_12892,N_5075,N_8322);
nor U12893 (N_12893,N_8394,N_8773);
nand U12894 (N_12894,N_7044,N_6930);
nor U12895 (N_12895,N_8915,N_8164);
xnor U12896 (N_12896,N_6177,N_6331);
and U12897 (N_12897,N_8535,N_7583);
and U12898 (N_12898,N_7530,N_9985);
and U12899 (N_12899,N_5965,N_5705);
nand U12900 (N_12900,N_9921,N_7793);
xor U12901 (N_12901,N_5280,N_7236);
nor U12902 (N_12902,N_9300,N_5560);
or U12903 (N_12903,N_9495,N_5752);
nand U12904 (N_12904,N_5502,N_7763);
and U12905 (N_12905,N_6707,N_8418);
and U12906 (N_12906,N_7600,N_7552);
or U12907 (N_12907,N_8991,N_6729);
nand U12908 (N_12908,N_8344,N_8449);
nor U12909 (N_12909,N_7751,N_8964);
xor U12910 (N_12910,N_5777,N_6305);
xnor U12911 (N_12911,N_5496,N_8541);
or U12912 (N_12912,N_7573,N_6454);
and U12913 (N_12913,N_7972,N_9297);
nand U12914 (N_12914,N_8981,N_6106);
xnor U12915 (N_12915,N_6686,N_9970);
xor U12916 (N_12916,N_9396,N_6468);
xnor U12917 (N_12917,N_7275,N_8284);
and U12918 (N_12918,N_9976,N_5581);
or U12919 (N_12919,N_5253,N_7518);
and U12920 (N_12920,N_8572,N_7387);
or U12921 (N_12921,N_7395,N_6115);
or U12922 (N_12922,N_5730,N_5548);
xor U12923 (N_12923,N_7422,N_7560);
or U12924 (N_12924,N_7048,N_6641);
nor U12925 (N_12925,N_9826,N_9615);
or U12926 (N_12926,N_8822,N_9263);
xor U12927 (N_12927,N_8078,N_7542);
nand U12928 (N_12928,N_5264,N_7723);
nor U12929 (N_12929,N_5673,N_5912);
and U12930 (N_12930,N_8134,N_9396);
and U12931 (N_12931,N_7913,N_7850);
and U12932 (N_12932,N_9744,N_5278);
and U12933 (N_12933,N_9830,N_6773);
nor U12934 (N_12934,N_8925,N_7276);
and U12935 (N_12935,N_7876,N_7340);
xor U12936 (N_12936,N_6986,N_7131);
nand U12937 (N_12937,N_8553,N_6299);
or U12938 (N_12938,N_6517,N_5856);
and U12939 (N_12939,N_8471,N_6619);
nor U12940 (N_12940,N_8973,N_9338);
nand U12941 (N_12941,N_9535,N_5096);
nor U12942 (N_12942,N_8723,N_9875);
and U12943 (N_12943,N_7308,N_9449);
and U12944 (N_12944,N_9410,N_9314);
xnor U12945 (N_12945,N_8880,N_6983);
and U12946 (N_12946,N_6904,N_6998);
or U12947 (N_12947,N_9854,N_7234);
xor U12948 (N_12948,N_6461,N_5533);
xor U12949 (N_12949,N_6962,N_6124);
or U12950 (N_12950,N_9311,N_5476);
xor U12951 (N_12951,N_8995,N_7821);
xnor U12952 (N_12952,N_5519,N_7722);
nand U12953 (N_12953,N_8653,N_9056);
nand U12954 (N_12954,N_6771,N_5098);
or U12955 (N_12955,N_7701,N_5934);
or U12956 (N_12956,N_5820,N_6041);
and U12957 (N_12957,N_9675,N_9028);
xor U12958 (N_12958,N_5409,N_8715);
xnor U12959 (N_12959,N_8473,N_6726);
and U12960 (N_12960,N_9184,N_6201);
and U12961 (N_12961,N_6206,N_8475);
and U12962 (N_12962,N_7970,N_6090);
nor U12963 (N_12963,N_5060,N_5597);
and U12964 (N_12964,N_5181,N_6302);
nor U12965 (N_12965,N_5102,N_8717);
nand U12966 (N_12966,N_7777,N_7751);
xor U12967 (N_12967,N_5954,N_8423);
xnor U12968 (N_12968,N_8589,N_9924);
and U12969 (N_12969,N_7751,N_6124);
or U12970 (N_12970,N_6526,N_5540);
xor U12971 (N_12971,N_5082,N_9099);
nor U12972 (N_12972,N_9510,N_9699);
nand U12973 (N_12973,N_5844,N_9100);
and U12974 (N_12974,N_7308,N_9977);
nor U12975 (N_12975,N_8240,N_8797);
nor U12976 (N_12976,N_8381,N_5062);
nor U12977 (N_12977,N_6968,N_7058);
and U12978 (N_12978,N_7020,N_8252);
nand U12979 (N_12979,N_6284,N_7268);
nor U12980 (N_12980,N_7944,N_5292);
or U12981 (N_12981,N_5266,N_9059);
nor U12982 (N_12982,N_9589,N_9082);
xor U12983 (N_12983,N_5386,N_8073);
xnor U12984 (N_12984,N_8086,N_9293);
and U12985 (N_12985,N_5378,N_7084);
nor U12986 (N_12986,N_7186,N_5397);
nand U12987 (N_12987,N_7669,N_6978);
xnor U12988 (N_12988,N_5722,N_9838);
nor U12989 (N_12989,N_6336,N_9061);
or U12990 (N_12990,N_5311,N_7084);
or U12991 (N_12991,N_6161,N_5884);
or U12992 (N_12992,N_7674,N_7191);
and U12993 (N_12993,N_8002,N_9741);
nand U12994 (N_12994,N_5552,N_5494);
nand U12995 (N_12995,N_8192,N_7140);
and U12996 (N_12996,N_8463,N_8701);
nand U12997 (N_12997,N_5186,N_7443);
nor U12998 (N_12998,N_7723,N_5643);
and U12999 (N_12999,N_6162,N_8088);
or U13000 (N_13000,N_6616,N_5872);
and U13001 (N_13001,N_8355,N_8891);
or U13002 (N_13002,N_7610,N_9403);
nor U13003 (N_13003,N_7982,N_7218);
nand U13004 (N_13004,N_5149,N_6023);
nor U13005 (N_13005,N_9193,N_5975);
and U13006 (N_13006,N_7939,N_5700);
xor U13007 (N_13007,N_6321,N_8410);
xnor U13008 (N_13008,N_7572,N_7205);
nor U13009 (N_13009,N_7993,N_6515);
nand U13010 (N_13010,N_9678,N_6250);
xor U13011 (N_13011,N_7745,N_6239);
nor U13012 (N_13012,N_8306,N_7087);
or U13013 (N_13013,N_6221,N_8486);
or U13014 (N_13014,N_5692,N_7708);
xor U13015 (N_13015,N_8501,N_6023);
or U13016 (N_13016,N_5396,N_9438);
nor U13017 (N_13017,N_9746,N_6863);
or U13018 (N_13018,N_6211,N_7448);
and U13019 (N_13019,N_7703,N_6128);
or U13020 (N_13020,N_8963,N_7756);
xor U13021 (N_13021,N_5096,N_5272);
and U13022 (N_13022,N_6436,N_6224);
or U13023 (N_13023,N_6682,N_6445);
nand U13024 (N_13024,N_7420,N_8141);
and U13025 (N_13025,N_9494,N_7768);
nor U13026 (N_13026,N_7317,N_6562);
and U13027 (N_13027,N_9371,N_7962);
xnor U13028 (N_13028,N_6559,N_5798);
nand U13029 (N_13029,N_8144,N_7529);
nor U13030 (N_13030,N_9510,N_9330);
xor U13031 (N_13031,N_6640,N_9138);
and U13032 (N_13032,N_7340,N_5157);
nand U13033 (N_13033,N_7991,N_6876);
and U13034 (N_13034,N_9106,N_6028);
and U13035 (N_13035,N_9767,N_5095);
xor U13036 (N_13036,N_5281,N_6604);
and U13037 (N_13037,N_9272,N_8265);
nor U13038 (N_13038,N_6471,N_7065);
nor U13039 (N_13039,N_9183,N_9209);
nand U13040 (N_13040,N_9801,N_7297);
and U13041 (N_13041,N_7645,N_5121);
nand U13042 (N_13042,N_5337,N_8197);
xor U13043 (N_13043,N_7430,N_7550);
or U13044 (N_13044,N_6396,N_6367);
nor U13045 (N_13045,N_9674,N_9767);
and U13046 (N_13046,N_7782,N_6085);
nor U13047 (N_13047,N_9785,N_5937);
nand U13048 (N_13048,N_9255,N_8341);
or U13049 (N_13049,N_5367,N_7442);
nand U13050 (N_13050,N_7128,N_8848);
or U13051 (N_13051,N_7145,N_9596);
nor U13052 (N_13052,N_6300,N_6408);
xnor U13053 (N_13053,N_5229,N_5417);
xor U13054 (N_13054,N_8939,N_8724);
nor U13055 (N_13055,N_5001,N_8434);
xor U13056 (N_13056,N_8377,N_7792);
and U13057 (N_13057,N_5244,N_8890);
xnor U13058 (N_13058,N_5117,N_9782);
nor U13059 (N_13059,N_6459,N_8543);
or U13060 (N_13060,N_6316,N_5358);
nand U13061 (N_13061,N_9575,N_8015);
and U13062 (N_13062,N_5304,N_5493);
or U13063 (N_13063,N_8067,N_7679);
xnor U13064 (N_13064,N_7474,N_7141);
or U13065 (N_13065,N_9607,N_5391);
xnor U13066 (N_13066,N_7990,N_7889);
or U13067 (N_13067,N_9955,N_8028);
or U13068 (N_13068,N_9793,N_8489);
nand U13069 (N_13069,N_7803,N_5573);
or U13070 (N_13070,N_8760,N_5216);
xor U13071 (N_13071,N_8330,N_5844);
or U13072 (N_13072,N_6581,N_8824);
and U13073 (N_13073,N_5662,N_9435);
xnor U13074 (N_13074,N_5995,N_9287);
and U13075 (N_13075,N_6177,N_6535);
nand U13076 (N_13076,N_5032,N_9272);
xnor U13077 (N_13077,N_6615,N_6654);
and U13078 (N_13078,N_5237,N_6857);
and U13079 (N_13079,N_6167,N_6788);
and U13080 (N_13080,N_8964,N_5820);
and U13081 (N_13081,N_8485,N_7551);
nand U13082 (N_13082,N_8597,N_9572);
xnor U13083 (N_13083,N_8201,N_5437);
nor U13084 (N_13084,N_5373,N_9193);
xnor U13085 (N_13085,N_6223,N_8413);
or U13086 (N_13086,N_7912,N_9479);
or U13087 (N_13087,N_8721,N_6080);
nor U13088 (N_13088,N_8008,N_8084);
nand U13089 (N_13089,N_6011,N_8907);
nor U13090 (N_13090,N_9347,N_6801);
xnor U13091 (N_13091,N_9146,N_8287);
or U13092 (N_13092,N_7081,N_9240);
xor U13093 (N_13093,N_8387,N_6976);
xor U13094 (N_13094,N_7492,N_5713);
nor U13095 (N_13095,N_7102,N_6430);
nand U13096 (N_13096,N_7117,N_7035);
nor U13097 (N_13097,N_6208,N_5012);
nor U13098 (N_13098,N_7786,N_9157);
xnor U13099 (N_13099,N_9747,N_8480);
nand U13100 (N_13100,N_8119,N_5231);
nor U13101 (N_13101,N_8209,N_8962);
nor U13102 (N_13102,N_5184,N_7030);
or U13103 (N_13103,N_5891,N_8258);
nand U13104 (N_13104,N_8965,N_8971);
nand U13105 (N_13105,N_5627,N_5707);
and U13106 (N_13106,N_9583,N_8910);
and U13107 (N_13107,N_9399,N_5069);
or U13108 (N_13108,N_9690,N_8829);
xnor U13109 (N_13109,N_5163,N_5017);
xnor U13110 (N_13110,N_8653,N_8403);
or U13111 (N_13111,N_5977,N_7099);
nand U13112 (N_13112,N_9928,N_9367);
and U13113 (N_13113,N_8555,N_8750);
or U13114 (N_13114,N_5611,N_7048);
nand U13115 (N_13115,N_9183,N_9459);
nand U13116 (N_13116,N_7104,N_9000);
xnor U13117 (N_13117,N_8312,N_7063);
nor U13118 (N_13118,N_9910,N_8120);
xnor U13119 (N_13119,N_5959,N_6568);
xor U13120 (N_13120,N_5480,N_5827);
nor U13121 (N_13121,N_8380,N_5245);
nor U13122 (N_13122,N_5979,N_8707);
xnor U13123 (N_13123,N_7456,N_9581);
xor U13124 (N_13124,N_6881,N_8969);
and U13125 (N_13125,N_5548,N_9948);
nand U13126 (N_13126,N_5271,N_8124);
and U13127 (N_13127,N_7016,N_7030);
nor U13128 (N_13128,N_7845,N_7490);
nor U13129 (N_13129,N_6496,N_7627);
xnor U13130 (N_13130,N_9793,N_6715);
nor U13131 (N_13131,N_9827,N_9535);
nand U13132 (N_13132,N_6520,N_7503);
or U13133 (N_13133,N_8998,N_6935);
nor U13134 (N_13134,N_5924,N_8599);
and U13135 (N_13135,N_7029,N_8810);
nand U13136 (N_13136,N_5662,N_6000);
nor U13137 (N_13137,N_7620,N_9075);
xor U13138 (N_13138,N_8650,N_6516);
and U13139 (N_13139,N_6447,N_7971);
nor U13140 (N_13140,N_5732,N_9951);
xor U13141 (N_13141,N_6947,N_5941);
or U13142 (N_13142,N_6566,N_5323);
and U13143 (N_13143,N_8479,N_5165);
and U13144 (N_13144,N_7123,N_5544);
or U13145 (N_13145,N_5148,N_5030);
nor U13146 (N_13146,N_9409,N_9594);
or U13147 (N_13147,N_8049,N_7816);
or U13148 (N_13148,N_6801,N_9999);
nand U13149 (N_13149,N_9304,N_7523);
nand U13150 (N_13150,N_7184,N_9847);
nor U13151 (N_13151,N_7138,N_5307);
or U13152 (N_13152,N_6571,N_7435);
or U13153 (N_13153,N_9523,N_7548);
xnor U13154 (N_13154,N_5566,N_8701);
nand U13155 (N_13155,N_6321,N_9498);
and U13156 (N_13156,N_9187,N_8682);
or U13157 (N_13157,N_6445,N_9184);
nor U13158 (N_13158,N_6942,N_7098);
or U13159 (N_13159,N_6237,N_6645);
nor U13160 (N_13160,N_6217,N_9881);
nand U13161 (N_13161,N_6641,N_8965);
xnor U13162 (N_13162,N_9254,N_5036);
nand U13163 (N_13163,N_8959,N_7151);
or U13164 (N_13164,N_6699,N_7977);
nor U13165 (N_13165,N_9602,N_5207);
nand U13166 (N_13166,N_8215,N_8918);
and U13167 (N_13167,N_7170,N_8208);
and U13168 (N_13168,N_8149,N_5312);
nand U13169 (N_13169,N_5766,N_9791);
xor U13170 (N_13170,N_8326,N_5352);
nor U13171 (N_13171,N_7704,N_7506);
and U13172 (N_13172,N_5292,N_7428);
nor U13173 (N_13173,N_7248,N_9977);
nor U13174 (N_13174,N_9219,N_7235);
nand U13175 (N_13175,N_6364,N_5572);
xor U13176 (N_13176,N_7213,N_5464);
nand U13177 (N_13177,N_9619,N_6782);
nand U13178 (N_13178,N_8621,N_7156);
xor U13179 (N_13179,N_5473,N_7060);
nor U13180 (N_13180,N_9768,N_7734);
nand U13181 (N_13181,N_5432,N_6978);
xnor U13182 (N_13182,N_5941,N_7732);
or U13183 (N_13183,N_5771,N_8992);
xor U13184 (N_13184,N_5617,N_5535);
nand U13185 (N_13185,N_9363,N_6318);
or U13186 (N_13186,N_7784,N_8763);
and U13187 (N_13187,N_6339,N_6057);
and U13188 (N_13188,N_9697,N_6279);
xnor U13189 (N_13189,N_7083,N_5309);
or U13190 (N_13190,N_6181,N_5212);
xor U13191 (N_13191,N_6826,N_8270);
nand U13192 (N_13192,N_5502,N_7596);
or U13193 (N_13193,N_6442,N_8002);
or U13194 (N_13194,N_7471,N_8574);
nor U13195 (N_13195,N_5993,N_9835);
xnor U13196 (N_13196,N_5082,N_7440);
or U13197 (N_13197,N_7122,N_9327);
nand U13198 (N_13198,N_6118,N_8431);
xor U13199 (N_13199,N_5548,N_6882);
or U13200 (N_13200,N_8120,N_9946);
and U13201 (N_13201,N_5661,N_6488);
xor U13202 (N_13202,N_9196,N_5259);
xor U13203 (N_13203,N_5916,N_8821);
or U13204 (N_13204,N_5166,N_7266);
nand U13205 (N_13205,N_8603,N_7289);
nor U13206 (N_13206,N_8879,N_9734);
and U13207 (N_13207,N_7374,N_7359);
and U13208 (N_13208,N_8370,N_8410);
nand U13209 (N_13209,N_7091,N_7146);
and U13210 (N_13210,N_8226,N_6222);
nand U13211 (N_13211,N_8243,N_7259);
nand U13212 (N_13212,N_7298,N_8306);
nor U13213 (N_13213,N_6086,N_7062);
nor U13214 (N_13214,N_9340,N_5475);
xor U13215 (N_13215,N_5664,N_6666);
nand U13216 (N_13216,N_6433,N_7219);
nor U13217 (N_13217,N_6434,N_5321);
and U13218 (N_13218,N_6872,N_9993);
nand U13219 (N_13219,N_6213,N_6646);
and U13220 (N_13220,N_5886,N_9888);
xnor U13221 (N_13221,N_9931,N_5608);
nor U13222 (N_13222,N_5404,N_5781);
and U13223 (N_13223,N_7917,N_5090);
xor U13224 (N_13224,N_7267,N_9674);
nand U13225 (N_13225,N_5654,N_8646);
or U13226 (N_13226,N_9179,N_8213);
and U13227 (N_13227,N_9895,N_9632);
or U13228 (N_13228,N_6762,N_5611);
nand U13229 (N_13229,N_5165,N_8980);
nor U13230 (N_13230,N_5725,N_7535);
xor U13231 (N_13231,N_7180,N_8939);
nor U13232 (N_13232,N_6159,N_6712);
nand U13233 (N_13233,N_5528,N_9379);
and U13234 (N_13234,N_7445,N_8571);
or U13235 (N_13235,N_9872,N_5688);
or U13236 (N_13236,N_5566,N_8400);
or U13237 (N_13237,N_6340,N_8002);
xor U13238 (N_13238,N_7484,N_6394);
nor U13239 (N_13239,N_9170,N_8668);
nand U13240 (N_13240,N_7138,N_9280);
and U13241 (N_13241,N_5347,N_9895);
or U13242 (N_13242,N_8169,N_8447);
xor U13243 (N_13243,N_7028,N_5172);
nor U13244 (N_13244,N_6118,N_8171);
nor U13245 (N_13245,N_7408,N_9230);
and U13246 (N_13246,N_6638,N_5110);
and U13247 (N_13247,N_6002,N_5989);
nand U13248 (N_13248,N_7302,N_9779);
and U13249 (N_13249,N_7582,N_8615);
and U13250 (N_13250,N_5167,N_8054);
nand U13251 (N_13251,N_6533,N_8195);
xor U13252 (N_13252,N_7950,N_6826);
xnor U13253 (N_13253,N_5816,N_9699);
or U13254 (N_13254,N_9636,N_6905);
nand U13255 (N_13255,N_7359,N_5223);
nand U13256 (N_13256,N_6810,N_6958);
xnor U13257 (N_13257,N_8115,N_8425);
or U13258 (N_13258,N_6488,N_8646);
xor U13259 (N_13259,N_9753,N_5672);
or U13260 (N_13260,N_8307,N_6803);
and U13261 (N_13261,N_8039,N_7558);
nand U13262 (N_13262,N_8577,N_8451);
xnor U13263 (N_13263,N_9377,N_7849);
and U13264 (N_13264,N_7782,N_8156);
and U13265 (N_13265,N_6250,N_5805);
or U13266 (N_13266,N_5734,N_8194);
or U13267 (N_13267,N_7977,N_6338);
nor U13268 (N_13268,N_9613,N_8364);
or U13269 (N_13269,N_8250,N_6394);
nor U13270 (N_13270,N_6778,N_5106);
or U13271 (N_13271,N_7670,N_6421);
or U13272 (N_13272,N_6454,N_5308);
and U13273 (N_13273,N_6546,N_7499);
nand U13274 (N_13274,N_5610,N_5260);
xnor U13275 (N_13275,N_5348,N_9766);
or U13276 (N_13276,N_9042,N_7758);
and U13277 (N_13277,N_8317,N_8252);
nor U13278 (N_13278,N_9480,N_7284);
nor U13279 (N_13279,N_9276,N_8119);
or U13280 (N_13280,N_8026,N_7076);
nand U13281 (N_13281,N_9504,N_6539);
nor U13282 (N_13282,N_7335,N_5454);
nand U13283 (N_13283,N_8547,N_7016);
xor U13284 (N_13284,N_6430,N_6534);
or U13285 (N_13285,N_8449,N_5069);
nor U13286 (N_13286,N_6247,N_6900);
nor U13287 (N_13287,N_8786,N_7094);
nand U13288 (N_13288,N_6344,N_9664);
or U13289 (N_13289,N_5942,N_6314);
or U13290 (N_13290,N_9370,N_8236);
nor U13291 (N_13291,N_9254,N_8926);
and U13292 (N_13292,N_9370,N_7057);
nor U13293 (N_13293,N_7867,N_7691);
xnor U13294 (N_13294,N_9366,N_7007);
nand U13295 (N_13295,N_6997,N_8753);
nor U13296 (N_13296,N_5963,N_5399);
xnor U13297 (N_13297,N_6085,N_9599);
or U13298 (N_13298,N_9475,N_6369);
and U13299 (N_13299,N_9359,N_9673);
xor U13300 (N_13300,N_8889,N_6567);
xor U13301 (N_13301,N_6885,N_6899);
nand U13302 (N_13302,N_5291,N_8756);
xnor U13303 (N_13303,N_5462,N_6771);
or U13304 (N_13304,N_7930,N_6336);
and U13305 (N_13305,N_7169,N_7820);
nor U13306 (N_13306,N_6395,N_5647);
nand U13307 (N_13307,N_6076,N_6848);
nor U13308 (N_13308,N_9102,N_7646);
or U13309 (N_13309,N_7360,N_5956);
nand U13310 (N_13310,N_7192,N_7692);
and U13311 (N_13311,N_8690,N_5038);
nand U13312 (N_13312,N_7434,N_5510);
xnor U13313 (N_13313,N_7857,N_6924);
or U13314 (N_13314,N_9072,N_8533);
and U13315 (N_13315,N_9401,N_6802);
nand U13316 (N_13316,N_7514,N_9098);
nand U13317 (N_13317,N_7759,N_9267);
or U13318 (N_13318,N_7428,N_8100);
xnor U13319 (N_13319,N_9521,N_8316);
or U13320 (N_13320,N_6642,N_8444);
nand U13321 (N_13321,N_9285,N_7551);
or U13322 (N_13322,N_8695,N_7123);
and U13323 (N_13323,N_6313,N_5152);
nand U13324 (N_13324,N_6106,N_6311);
xnor U13325 (N_13325,N_5293,N_8676);
and U13326 (N_13326,N_7907,N_6656);
or U13327 (N_13327,N_6445,N_5292);
nor U13328 (N_13328,N_6533,N_7078);
or U13329 (N_13329,N_8757,N_9214);
xnor U13330 (N_13330,N_8855,N_5167);
nand U13331 (N_13331,N_5154,N_9376);
nand U13332 (N_13332,N_7967,N_5663);
or U13333 (N_13333,N_7971,N_7936);
nand U13334 (N_13334,N_8058,N_7906);
and U13335 (N_13335,N_9206,N_9778);
xnor U13336 (N_13336,N_8444,N_8636);
nand U13337 (N_13337,N_9089,N_8958);
xor U13338 (N_13338,N_5386,N_5895);
and U13339 (N_13339,N_7825,N_5107);
nand U13340 (N_13340,N_7696,N_5628);
xnor U13341 (N_13341,N_5856,N_9708);
nand U13342 (N_13342,N_8533,N_5684);
or U13343 (N_13343,N_6405,N_7696);
xnor U13344 (N_13344,N_9426,N_8408);
nor U13345 (N_13345,N_6912,N_7042);
and U13346 (N_13346,N_9277,N_9805);
or U13347 (N_13347,N_9735,N_5917);
nand U13348 (N_13348,N_7408,N_8063);
xnor U13349 (N_13349,N_5201,N_9398);
and U13350 (N_13350,N_5296,N_5699);
and U13351 (N_13351,N_5071,N_5629);
nor U13352 (N_13352,N_5346,N_5445);
and U13353 (N_13353,N_6196,N_5863);
nand U13354 (N_13354,N_5501,N_8940);
nor U13355 (N_13355,N_7604,N_6013);
xor U13356 (N_13356,N_8415,N_5641);
xor U13357 (N_13357,N_8724,N_7620);
nor U13358 (N_13358,N_9212,N_6533);
nand U13359 (N_13359,N_6215,N_8218);
nand U13360 (N_13360,N_5448,N_9502);
xor U13361 (N_13361,N_5280,N_8372);
or U13362 (N_13362,N_9570,N_7040);
or U13363 (N_13363,N_9159,N_6542);
nor U13364 (N_13364,N_7049,N_8297);
nor U13365 (N_13365,N_6099,N_7243);
xnor U13366 (N_13366,N_9542,N_6837);
and U13367 (N_13367,N_7629,N_6772);
and U13368 (N_13368,N_6562,N_7406);
and U13369 (N_13369,N_5720,N_9128);
and U13370 (N_13370,N_5247,N_7110);
nor U13371 (N_13371,N_6110,N_9640);
or U13372 (N_13372,N_7528,N_5739);
and U13373 (N_13373,N_7583,N_5810);
nand U13374 (N_13374,N_6462,N_6820);
nand U13375 (N_13375,N_9268,N_5677);
and U13376 (N_13376,N_9792,N_6440);
xnor U13377 (N_13377,N_7399,N_7799);
or U13378 (N_13378,N_5163,N_6293);
nor U13379 (N_13379,N_9885,N_6882);
and U13380 (N_13380,N_6254,N_8999);
and U13381 (N_13381,N_9562,N_5005);
nor U13382 (N_13382,N_8741,N_6988);
nor U13383 (N_13383,N_7282,N_9454);
nand U13384 (N_13384,N_7717,N_7311);
nand U13385 (N_13385,N_6335,N_5871);
or U13386 (N_13386,N_7636,N_7234);
and U13387 (N_13387,N_7945,N_5458);
nor U13388 (N_13388,N_5410,N_5136);
nor U13389 (N_13389,N_7864,N_6699);
xnor U13390 (N_13390,N_5199,N_6529);
and U13391 (N_13391,N_5076,N_5297);
xnor U13392 (N_13392,N_9049,N_7586);
xnor U13393 (N_13393,N_7329,N_7088);
xor U13394 (N_13394,N_8417,N_7927);
and U13395 (N_13395,N_7763,N_7307);
nand U13396 (N_13396,N_5265,N_9108);
xnor U13397 (N_13397,N_5122,N_5900);
xor U13398 (N_13398,N_6326,N_5991);
and U13399 (N_13399,N_9936,N_6280);
nand U13400 (N_13400,N_5681,N_9830);
nand U13401 (N_13401,N_8255,N_5281);
nor U13402 (N_13402,N_7651,N_5147);
xnor U13403 (N_13403,N_7358,N_9587);
xor U13404 (N_13404,N_7850,N_5476);
nor U13405 (N_13405,N_8607,N_8754);
nor U13406 (N_13406,N_7287,N_5502);
and U13407 (N_13407,N_7766,N_9532);
xnor U13408 (N_13408,N_5842,N_6198);
and U13409 (N_13409,N_8161,N_5586);
xnor U13410 (N_13410,N_9654,N_9888);
nand U13411 (N_13411,N_9325,N_9939);
or U13412 (N_13412,N_9668,N_5627);
nor U13413 (N_13413,N_5011,N_8117);
nor U13414 (N_13414,N_8595,N_5990);
or U13415 (N_13415,N_7459,N_7924);
nand U13416 (N_13416,N_8593,N_8208);
nor U13417 (N_13417,N_6226,N_8834);
xnor U13418 (N_13418,N_7692,N_7724);
nand U13419 (N_13419,N_6988,N_7462);
nand U13420 (N_13420,N_7248,N_5023);
or U13421 (N_13421,N_9531,N_7290);
nand U13422 (N_13422,N_7966,N_8350);
xor U13423 (N_13423,N_5194,N_5698);
and U13424 (N_13424,N_8649,N_7602);
or U13425 (N_13425,N_6932,N_7484);
xnor U13426 (N_13426,N_7258,N_9592);
nand U13427 (N_13427,N_6979,N_5489);
xor U13428 (N_13428,N_7113,N_6786);
and U13429 (N_13429,N_7227,N_8354);
and U13430 (N_13430,N_7070,N_9488);
or U13431 (N_13431,N_6440,N_6292);
nand U13432 (N_13432,N_8830,N_8081);
xor U13433 (N_13433,N_7426,N_7152);
or U13434 (N_13434,N_5517,N_9372);
or U13435 (N_13435,N_9306,N_6329);
nand U13436 (N_13436,N_6134,N_5403);
or U13437 (N_13437,N_7720,N_9546);
or U13438 (N_13438,N_7934,N_8855);
nand U13439 (N_13439,N_9659,N_6443);
xnor U13440 (N_13440,N_7204,N_9840);
or U13441 (N_13441,N_7312,N_9951);
nand U13442 (N_13442,N_8507,N_8581);
nor U13443 (N_13443,N_9887,N_8256);
xor U13444 (N_13444,N_7499,N_9436);
or U13445 (N_13445,N_7700,N_7346);
and U13446 (N_13446,N_7665,N_7609);
nand U13447 (N_13447,N_7785,N_6460);
and U13448 (N_13448,N_9133,N_9893);
nand U13449 (N_13449,N_8388,N_8854);
and U13450 (N_13450,N_8098,N_8927);
nand U13451 (N_13451,N_8727,N_5175);
or U13452 (N_13452,N_5147,N_8839);
and U13453 (N_13453,N_5674,N_9280);
nand U13454 (N_13454,N_7669,N_6676);
or U13455 (N_13455,N_7112,N_7737);
nand U13456 (N_13456,N_6333,N_7882);
nor U13457 (N_13457,N_5538,N_7744);
or U13458 (N_13458,N_5015,N_8844);
or U13459 (N_13459,N_8526,N_7727);
or U13460 (N_13460,N_8115,N_5443);
nor U13461 (N_13461,N_5851,N_9074);
nor U13462 (N_13462,N_8544,N_6184);
or U13463 (N_13463,N_9593,N_9799);
or U13464 (N_13464,N_7973,N_9553);
or U13465 (N_13465,N_9595,N_6884);
xnor U13466 (N_13466,N_6691,N_5743);
xor U13467 (N_13467,N_5233,N_6675);
nand U13468 (N_13468,N_5642,N_6378);
and U13469 (N_13469,N_9090,N_5432);
nor U13470 (N_13470,N_5221,N_6507);
nor U13471 (N_13471,N_8507,N_5318);
nand U13472 (N_13472,N_7741,N_6039);
nand U13473 (N_13473,N_6195,N_5707);
nor U13474 (N_13474,N_7954,N_5694);
nand U13475 (N_13475,N_6290,N_8757);
xor U13476 (N_13476,N_7566,N_7537);
xnor U13477 (N_13477,N_5737,N_7322);
nand U13478 (N_13478,N_5292,N_6806);
or U13479 (N_13479,N_8169,N_5824);
xor U13480 (N_13480,N_8422,N_8893);
nor U13481 (N_13481,N_5609,N_7808);
xor U13482 (N_13482,N_8742,N_7332);
or U13483 (N_13483,N_5736,N_9164);
xnor U13484 (N_13484,N_5165,N_6278);
xnor U13485 (N_13485,N_7371,N_9434);
xor U13486 (N_13486,N_6878,N_5304);
nand U13487 (N_13487,N_5904,N_8055);
and U13488 (N_13488,N_5880,N_9167);
xnor U13489 (N_13489,N_6124,N_7260);
nor U13490 (N_13490,N_7685,N_7312);
or U13491 (N_13491,N_6849,N_8348);
or U13492 (N_13492,N_7877,N_7531);
nor U13493 (N_13493,N_5104,N_9818);
or U13494 (N_13494,N_5547,N_5586);
nand U13495 (N_13495,N_7345,N_8664);
nand U13496 (N_13496,N_7797,N_7064);
or U13497 (N_13497,N_8491,N_9704);
xor U13498 (N_13498,N_7474,N_7812);
xnor U13499 (N_13499,N_5089,N_9087);
nand U13500 (N_13500,N_8727,N_7146);
and U13501 (N_13501,N_8692,N_6642);
xor U13502 (N_13502,N_9221,N_8262);
or U13503 (N_13503,N_8754,N_9946);
and U13504 (N_13504,N_8725,N_6951);
or U13505 (N_13505,N_6714,N_9568);
nand U13506 (N_13506,N_8225,N_6416);
nor U13507 (N_13507,N_9422,N_8218);
or U13508 (N_13508,N_7427,N_5528);
or U13509 (N_13509,N_6633,N_9551);
nor U13510 (N_13510,N_9548,N_9527);
nand U13511 (N_13511,N_7279,N_9904);
xor U13512 (N_13512,N_5488,N_9859);
and U13513 (N_13513,N_9112,N_9509);
nand U13514 (N_13514,N_6938,N_9218);
xor U13515 (N_13515,N_8146,N_9126);
or U13516 (N_13516,N_7314,N_6063);
nor U13517 (N_13517,N_6229,N_7080);
nor U13518 (N_13518,N_9249,N_6901);
xnor U13519 (N_13519,N_6866,N_9387);
nand U13520 (N_13520,N_9272,N_6745);
xnor U13521 (N_13521,N_6096,N_6932);
nand U13522 (N_13522,N_5945,N_6981);
and U13523 (N_13523,N_9134,N_9625);
or U13524 (N_13524,N_9859,N_9403);
nand U13525 (N_13525,N_5280,N_9106);
xnor U13526 (N_13526,N_8064,N_5994);
xor U13527 (N_13527,N_5829,N_7898);
or U13528 (N_13528,N_7113,N_9922);
and U13529 (N_13529,N_5871,N_5742);
nand U13530 (N_13530,N_9262,N_6440);
xor U13531 (N_13531,N_5547,N_7733);
or U13532 (N_13532,N_5524,N_9478);
and U13533 (N_13533,N_9005,N_6317);
and U13534 (N_13534,N_6400,N_7288);
xor U13535 (N_13535,N_6352,N_8751);
nand U13536 (N_13536,N_8194,N_7402);
nor U13537 (N_13537,N_8091,N_7586);
or U13538 (N_13538,N_8339,N_5969);
and U13539 (N_13539,N_6865,N_9453);
or U13540 (N_13540,N_8152,N_7034);
and U13541 (N_13541,N_7405,N_9610);
or U13542 (N_13542,N_7397,N_6618);
and U13543 (N_13543,N_5582,N_9635);
nor U13544 (N_13544,N_5771,N_5988);
and U13545 (N_13545,N_8280,N_5914);
nor U13546 (N_13546,N_7447,N_6372);
nor U13547 (N_13547,N_8423,N_9571);
nand U13548 (N_13548,N_8876,N_6837);
xor U13549 (N_13549,N_9145,N_6906);
or U13550 (N_13550,N_8220,N_7956);
and U13551 (N_13551,N_6498,N_5622);
xor U13552 (N_13552,N_8071,N_7167);
and U13553 (N_13553,N_6537,N_9864);
and U13554 (N_13554,N_7062,N_5995);
nand U13555 (N_13555,N_5695,N_9778);
and U13556 (N_13556,N_7672,N_8567);
xnor U13557 (N_13557,N_9173,N_8937);
nor U13558 (N_13558,N_5917,N_5129);
nand U13559 (N_13559,N_8278,N_6374);
or U13560 (N_13560,N_9041,N_8047);
xor U13561 (N_13561,N_8812,N_7521);
and U13562 (N_13562,N_6514,N_9114);
xnor U13563 (N_13563,N_5182,N_7731);
and U13564 (N_13564,N_8986,N_6295);
or U13565 (N_13565,N_6626,N_9204);
or U13566 (N_13566,N_8964,N_5205);
xnor U13567 (N_13567,N_7652,N_7450);
nor U13568 (N_13568,N_5302,N_6690);
or U13569 (N_13569,N_5478,N_8927);
or U13570 (N_13570,N_6019,N_6963);
xor U13571 (N_13571,N_5444,N_5056);
nor U13572 (N_13572,N_5698,N_9858);
nor U13573 (N_13573,N_9384,N_9059);
nand U13574 (N_13574,N_8956,N_6775);
nand U13575 (N_13575,N_6825,N_7582);
nand U13576 (N_13576,N_9003,N_8030);
nand U13577 (N_13577,N_7500,N_7728);
and U13578 (N_13578,N_5592,N_6625);
nand U13579 (N_13579,N_8173,N_9097);
xor U13580 (N_13580,N_5749,N_8925);
nand U13581 (N_13581,N_5395,N_6289);
nor U13582 (N_13582,N_6719,N_7087);
and U13583 (N_13583,N_5794,N_5029);
or U13584 (N_13584,N_9461,N_6656);
nand U13585 (N_13585,N_7018,N_8375);
xor U13586 (N_13586,N_6349,N_9084);
and U13587 (N_13587,N_5737,N_5524);
or U13588 (N_13588,N_7386,N_9827);
or U13589 (N_13589,N_6420,N_8664);
nor U13590 (N_13590,N_5822,N_9487);
nor U13591 (N_13591,N_8092,N_7467);
and U13592 (N_13592,N_7446,N_8571);
or U13593 (N_13593,N_8321,N_7321);
xor U13594 (N_13594,N_5409,N_7156);
or U13595 (N_13595,N_5243,N_8422);
and U13596 (N_13596,N_9534,N_6428);
nor U13597 (N_13597,N_8116,N_9305);
and U13598 (N_13598,N_6919,N_9107);
nand U13599 (N_13599,N_7127,N_9773);
nand U13600 (N_13600,N_8156,N_6251);
xor U13601 (N_13601,N_6426,N_6689);
nor U13602 (N_13602,N_5133,N_6787);
and U13603 (N_13603,N_9110,N_5285);
nand U13604 (N_13604,N_8537,N_8914);
nand U13605 (N_13605,N_7689,N_9305);
nand U13606 (N_13606,N_6665,N_6801);
nand U13607 (N_13607,N_6273,N_5905);
xor U13608 (N_13608,N_9698,N_7831);
nor U13609 (N_13609,N_6105,N_5087);
nand U13610 (N_13610,N_8209,N_9190);
nand U13611 (N_13611,N_7743,N_9401);
nand U13612 (N_13612,N_7283,N_6300);
nand U13613 (N_13613,N_8788,N_9054);
or U13614 (N_13614,N_5138,N_8347);
xnor U13615 (N_13615,N_9130,N_9297);
and U13616 (N_13616,N_5024,N_5204);
or U13617 (N_13617,N_7845,N_6412);
or U13618 (N_13618,N_5705,N_7156);
xnor U13619 (N_13619,N_7340,N_8048);
and U13620 (N_13620,N_5814,N_7934);
nand U13621 (N_13621,N_6708,N_5039);
or U13622 (N_13622,N_8178,N_5303);
xnor U13623 (N_13623,N_9907,N_6244);
or U13624 (N_13624,N_5772,N_5428);
xnor U13625 (N_13625,N_6126,N_5680);
and U13626 (N_13626,N_8113,N_6304);
and U13627 (N_13627,N_8922,N_9851);
or U13628 (N_13628,N_7526,N_5444);
or U13629 (N_13629,N_7517,N_7542);
nand U13630 (N_13630,N_8932,N_8797);
nand U13631 (N_13631,N_5730,N_6980);
xnor U13632 (N_13632,N_5141,N_6780);
nor U13633 (N_13633,N_5723,N_8609);
nor U13634 (N_13634,N_9757,N_9812);
nor U13635 (N_13635,N_6304,N_7912);
nor U13636 (N_13636,N_8595,N_6262);
nor U13637 (N_13637,N_9784,N_7696);
xnor U13638 (N_13638,N_7861,N_8302);
and U13639 (N_13639,N_5283,N_7001);
nor U13640 (N_13640,N_5926,N_7406);
nand U13641 (N_13641,N_6429,N_9969);
and U13642 (N_13642,N_5089,N_9196);
nor U13643 (N_13643,N_9097,N_8842);
and U13644 (N_13644,N_5414,N_6463);
and U13645 (N_13645,N_8011,N_9345);
nand U13646 (N_13646,N_6731,N_9742);
and U13647 (N_13647,N_7781,N_8128);
nor U13648 (N_13648,N_9849,N_9758);
and U13649 (N_13649,N_7461,N_9807);
and U13650 (N_13650,N_8855,N_9666);
and U13651 (N_13651,N_7142,N_6225);
nand U13652 (N_13652,N_7656,N_8758);
and U13653 (N_13653,N_9294,N_5633);
or U13654 (N_13654,N_9141,N_5746);
nand U13655 (N_13655,N_7636,N_6292);
xnor U13656 (N_13656,N_9303,N_8427);
nand U13657 (N_13657,N_5247,N_5962);
nand U13658 (N_13658,N_5866,N_9106);
xor U13659 (N_13659,N_9422,N_8590);
xnor U13660 (N_13660,N_5244,N_7128);
nand U13661 (N_13661,N_8821,N_8738);
xnor U13662 (N_13662,N_8541,N_8032);
and U13663 (N_13663,N_9456,N_7640);
xor U13664 (N_13664,N_8583,N_8909);
xor U13665 (N_13665,N_9851,N_8014);
nor U13666 (N_13666,N_7259,N_6124);
and U13667 (N_13667,N_6492,N_6349);
nand U13668 (N_13668,N_8310,N_8079);
nor U13669 (N_13669,N_9191,N_8765);
and U13670 (N_13670,N_9020,N_5595);
xor U13671 (N_13671,N_9912,N_5912);
nor U13672 (N_13672,N_9004,N_5527);
nand U13673 (N_13673,N_6907,N_6950);
nand U13674 (N_13674,N_9834,N_7170);
nand U13675 (N_13675,N_7444,N_9867);
nor U13676 (N_13676,N_8156,N_8491);
or U13677 (N_13677,N_5118,N_5380);
nand U13678 (N_13678,N_8294,N_9037);
nand U13679 (N_13679,N_6605,N_9938);
nor U13680 (N_13680,N_9446,N_5771);
nand U13681 (N_13681,N_7935,N_5760);
xor U13682 (N_13682,N_6159,N_6586);
and U13683 (N_13683,N_5707,N_8720);
or U13684 (N_13684,N_8106,N_6009);
xnor U13685 (N_13685,N_9266,N_5532);
and U13686 (N_13686,N_8956,N_6722);
nand U13687 (N_13687,N_8770,N_6152);
xor U13688 (N_13688,N_7417,N_7725);
xnor U13689 (N_13689,N_6507,N_9129);
nand U13690 (N_13690,N_7115,N_8623);
nor U13691 (N_13691,N_5150,N_7999);
nor U13692 (N_13692,N_6663,N_8174);
xnor U13693 (N_13693,N_5137,N_6964);
or U13694 (N_13694,N_6398,N_9137);
or U13695 (N_13695,N_5106,N_8977);
or U13696 (N_13696,N_8255,N_8257);
nand U13697 (N_13697,N_8388,N_7815);
and U13698 (N_13698,N_5041,N_6838);
nand U13699 (N_13699,N_6937,N_6767);
or U13700 (N_13700,N_8632,N_5245);
nand U13701 (N_13701,N_5052,N_7764);
nor U13702 (N_13702,N_7671,N_5224);
xnor U13703 (N_13703,N_7599,N_8665);
and U13704 (N_13704,N_9359,N_8035);
xor U13705 (N_13705,N_8338,N_9064);
xnor U13706 (N_13706,N_9404,N_9729);
nand U13707 (N_13707,N_5792,N_7740);
or U13708 (N_13708,N_8752,N_6704);
nand U13709 (N_13709,N_6652,N_9950);
xnor U13710 (N_13710,N_6736,N_8147);
nand U13711 (N_13711,N_7369,N_6533);
and U13712 (N_13712,N_6978,N_5594);
and U13713 (N_13713,N_7632,N_6150);
or U13714 (N_13714,N_9792,N_8941);
nor U13715 (N_13715,N_6804,N_7897);
and U13716 (N_13716,N_7318,N_6840);
nand U13717 (N_13717,N_8230,N_8760);
nor U13718 (N_13718,N_8389,N_8513);
or U13719 (N_13719,N_9480,N_8775);
nand U13720 (N_13720,N_7940,N_6074);
nor U13721 (N_13721,N_6112,N_5577);
nor U13722 (N_13722,N_6156,N_5327);
xor U13723 (N_13723,N_8041,N_9249);
xor U13724 (N_13724,N_5951,N_9764);
and U13725 (N_13725,N_7284,N_7799);
nor U13726 (N_13726,N_5699,N_7945);
nor U13727 (N_13727,N_9077,N_9804);
and U13728 (N_13728,N_8184,N_6493);
nand U13729 (N_13729,N_8394,N_8869);
and U13730 (N_13730,N_7312,N_5358);
nand U13731 (N_13731,N_6038,N_7180);
nand U13732 (N_13732,N_8423,N_5759);
nand U13733 (N_13733,N_5246,N_5660);
nor U13734 (N_13734,N_8915,N_5722);
nand U13735 (N_13735,N_7242,N_9952);
or U13736 (N_13736,N_7136,N_5125);
nand U13737 (N_13737,N_5603,N_6092);
nand U13738 (N_13738,N_5403,N_8899);
or U13739 (N_13739,N_6715,N_7569);
or U13740 (N_13740,N_6636,N_6044);
and U13741 (N_13741,N_6631,N_9296);
nand U13742 (N_13742,N_9845,N_6970);
nor U13743 (N_13743,N_9938,N_8126);
nand U13744 (N_13744,N_5688,N_9073);
and U13745 (N_13745,N_9150,N_7038);
nor U13746 (N_13746,N_5874,N_8896);
xnor U13747 (N_13747,N_7386,N_8624);
nand U13748 (N_13748,N_5439,N_6067);
or U13749 (N_13749,N_6554,N_5783);
nand U13750 (N_13750,N_9623,N_9795);
nor U13751 (N_13751,N_9167,N_9195);
nand U13752 (N_13752,N_6155,N_7000);
or U13753 (N_13753,N_7198,N_7873);
or U13754 (N_13754,N_8291,N_5491);
and U13755 (N_13755,N_8364,N_7869);
and U13756 (N_13756,N_8477,N_8625);
or U13757 (N_13757,N_6727,N_8008);
and U13758 (N_13758,N_8619,N_9140);
and U13759 (N_13759,N_5584,N_9902);
or U13760 (N_13760,N_8268,N_6299);
or U13761 (N_13761,N_7351,N_6147);
nand U13762 (N_13762,N_5585,N_7697);
nand U13763 (N_13763,N_5853,N_7329);
nand U13764 (N_13764,N_6499,N_6816);
nand U13765 (N_13765,N_7915,N_8776);
nand U13766 (N_13766,N_9737,N_7024);
xnor U13767 (N_13767,N_5852,N_6302);
xnor U13768 (N_13768,N_8972,N_6061);
nand U13769 (N_13769,N_6926,N_8223);
nor U13770 (N_13770,N_9795,N_8815);
or U13771 (N_13771,N_6520,N_9233);
xnor U13772 (N_13772,N_8671,N_7980);
xnor U13773 (N_13773,N_8304,N_5004);
xor U13774 (N_13774,N_7345,N_8258);
and U13775 (N_13775,N_6743,N_9590);
and U13776 (N_13776,N_6590,N_7833);
and U13777 (N_13777,N_8970,N_6755);
xor U13778 (N_13778,N_8980,N_9543);
xor U13779 (N_13779,N_8760,N_8677);
nand U13780 (N_13780,N_9610,N_8282);
nor U13781 (N_13781,N_9254,N_5696);
and U13782 (N_13782,N_8131,N_7044);
xnor U13783 (N_13783,N_8794,N_7622);
nand U13784 (N_13784,N_9498,N_6365);
nand U13785 (N_13785,N_7931,N_9743);
or U13786 (N_13786,N_5457,N_7649);
or U13787 (N_13787,N_7080,N_7651);
nand U13788 (N_13788,N_8816,N_6729);
and U13789 (N_13789,N_9565,N_9283);
xnor U13790 (N_13790,N_6506,N_9269);
or U13791 (N_13791,N_8434,N_7492);
and U13792 (N_13792,N_9046,N_9911);
xnor U13793 (N_13793,N_8097,N_8736);
nand U13794 (N_13794,N_5220,N_9125);
xnor U13795 (N_13795,N_8424,N_5782);
and U13796 (N_13796,N_7552,N_5010);
and U13797 (N_13797,N_6393,N_8830);
nor U13798 (N_13798,N_7702,N_6573);
nand U13799 (N_13799,N_9053,N_5446);
nor U13800 (N_13800,N_9728,N_9837);
xor U13801 (N_13801,N_8765,N_9310);
nand U13802 (N_13802,N_5922,N_9892);
xnor U13803 (N_13803,N_7961,N_7703);
and U13804 (N_13804,N_5152,N_6871);
nand U13805 (N_13805,N_8503,N_8052);
and U13806 (N_13806,N_9011,N_6630);
nand U13807 (N_13807,N_5442,N_8168);
nor U13808 (N_13808,N_8826,N_9188);
or U13809 (N_13809,N_9729,N_7060);
nand U13810 (N_13810,N_6745,N_9876);
xor U13811 (N_13811,N_5502,N_9818);
nand U13812 (N_13812,N_7665,N_6313);
or U13813 (N_13813,N_8689,N_7545);
or U13814 (N_13814,N_7650,N_6461);
nor U13815 (N_13815,N_8079,N_8795);
or U13816 (N_13816,N_9416,N_7267);
and U13817 (N_13817,N_6912,N_6409);
xor U13818 (N_13818,N_5152,N_8031);
xnor U13819 (N_13819,N_5646,N_9151);
and U13820 (N_13820,N_6728,N_8579);
nor U13821 (N_13821,N_7542,N_5093);
nor U13822 (N_13822,N_5281,N_5049);
and U13823 (N_13823,N_9381,N_7034);
or U13824 (N_13824,N_7319,N_9301);
nor U13825 (N_13825,N_9529,N_6642);
nor U13826 (N_13826,N_8915,N_5796);
or U13827 (N_13827,N_8374,N_9146);
or U13828 (N_13828,N_5493,N_5890);
and U13829 (N_13829,N_8880,N_7336);
nand U13830 (N_13830,N_6758,N_6488);
nand U13831 (N_13831,N_8987,N_5840);
or U13832 (N_13832,N_6284,N_6453);
and U13833 (N_13833,N_5967,N_6905);
or U13834 (N_13834,N_5511,N_5076);
xnor U13835 (N_13835,N_6801,N_7773);
nand U13836 (N_13836,N_6172,N_7219);
nand U13837 (N_13837,N_6934,N_8388);
nor U13838 (N_13838,N_5254,N_6404);
xor U13839 (N_13839,N_5256,N_8120);
xor U13840 (N_13840,N_7943,N_8517);
nand U13841 (N_13841,N_8771,N_8973);
and U13842 (N_13842,N_8712,N_6230);
nand U13843 (N_13843,N_8483,N_8453);
and U13844 (N_13844,N_7649,N_6352);
and U13845 (N_13845,N_9212,N_6607);
nor U13846 (N_13846,N_5217,N_7018);
nor U13847 (N_13847,N_7427,N_8281);
xnor U13848 (N_13848,N_8732,N_8342);
nand U13849 (N_13849,N_5769,N_7652);
xor U13850 (N_13850,N_8866,N_8542);
nor U13851 (N_13851,N_5217,N_7080);
and U13852 (N_13852,N_9924,N_8140);
nand U13853 (N_13853,N_5241,N_8817);
and U13854 (N_13854,N_6870,N_8625);
and U13855 (N_13855,N_8972,N_9295);
nand U13856 (N_13856,N_9546,N_6386);
and U13857 (N_13857,N_5665,N_9966);
xor U13858 (N_13858,N_9651,N_7917);
nor U13859 (N_13859,N_7762,N_6395);
and U13860 (N_13860,N_8794,N_7037);
nor U13861 (N_13861,N_6551,N_7648);
xnor U13862 (N_13862,N_8482,N_5887);
and U13863 (N_13863,N_8626,N_5789);
or U13864 (N_13864,N_8110,N_5287);
or U13865 (N_13865,N_7181,N_8240);
and U13866 (N_13866,N_7683,N_7333);
and U13867 (N_13867,N_5918,N_9389);
nand U13868 (N_13868,N_5056,N_8305);
nor U13869 (N_13869,N_5497,N_6462);
or U13870 (N_13870,N_9305,N_7658);
nand U13871 (N_13871,N_8177,N_5476);
and U13872 (N_13872,N_6992,N_8208);
nor U13873 (N_13873,N_7331,N_5898);
and U13874 (N_13874,N_8993,N_9186);
or U13875 (N_13875,N_9183,N_9273);
xor U13876 (N_13876,N_8274,N_8958);
or U13877 (N_13877,N_6358,N_9946);
and U13878 (N_13878,N_9771,N_5309);
or U13879 (N_13879,N_5234,N_9010);
or U13880 (N_13880,N_9533,N_5339);
nor U13881 (N_13881,N_9261,N_6975);
xnor U13882 (N_13882,N_5253,N_7669);
or U13883 (N_13883,N_6351,N_6506);
xor U13884 (N_13884,N_7090,N_6194);
xor U13885 (N_13885,N_5149,N_9560);
and U13886 (N_13886,N_5529,N_5179);
and U13887 (N_13887,N_8914,N_9006);
xor U13888 (N_13888,N_9528,N_7330);
and U13889 (N_13889,N_8103,N_6190);
nor U13890 (N_13890,N_8581,N_9924);
or U13891 (N_13891,N_7638,N_5174);
or U13892 (N_13892,N_6277,N_6270);
nor U13893 (N_13893,N_5840,N_8414);
or U13894 (N_13894,N_7467,N_6035);
or U13895 (N_13895,N_9330,N_6085);
or U13896 (N_13896,N_6064,N_5227);
and U13897 (N_13897,N_7114,N_8336);
nand U13898 (N_13898,N_9857,N_9158);
nor U13899 (N_13899,N_7776,N_5268);
nor U13900 (N_13900,N_5653,N_5599);
or U13901 (N_13901,N_9191,N_6986);
nand U13902 (N_13902,N_8431,N_8633);
nand U13903 (N_13903,N_5472,N_8700);
or U13904 (N_13904,N_7879,N_7044);
xor U13905 (N_13905,N_5079,N_9339);
and U13906 (N_13906,N_5431,N_7874);
or U13907 (N_13907,N_5017,N_5924);
and U13908 (N_13908,N_8568,N_8376);
or U13909 (N_13909,N_8392,N_6330);
xnor U13910 (N_13910,N_5812,N_7222);
or U13911 (N_13911,N_5897,N_6263);
or U13912 (N_13912,N_5879,N_5217);
or U13913 (N_13913,N_6172,N_5436);
nor U13914 (N_13914,N_8349,N_8966);
and U13915 (N_13915,N_8602,N_7328);
or U13916 (N_13916,N_8653,N_6933);
or U13917 (N_13917,N_9208,N_8357);
nor U13918 (N_13918,N_6160,N_7591);
and U13919 (N_13919,N_5802,N_9854);
nand U13920 (N_13920,N_9610,N_5796);
and U13921 (N_13921,N_5156,N_6680);
nand U13922 (N_13922,N_9889,N_6798);
and U13923 (N_13923,N_8268,N_8401);
nand U13924 (N_13924,N_8642,N_6861);
nor U13925 (N_13925,N_8115,N_9914);
or U13926 (N_13926,N_9399,N_9973);
xnor U13927 (N_13927,N_6994,N_6287);
or U13928 (N_13928,N_9390,N_5962);
and U13929 (N_13929,N_7249,N_6160);
nor U13930 (N_13930,N_7896,N_9115);
nor U13931 (N_13931,N_6802,N_6818);
xnor U13932 (N_13932,N_8841,N_6637);
nand U13933 (N_13933,N_5209,N_5387);
or U13934 (N_13934,N_7930,N_8500);
or U13935 (N_13935,N_9459,N_9938);
nor U13936 (N_13936,N_9703,N_5976);
nand U13937 (N_13937,N_7896,N_7196);
nand U13938 (N_13938,N_7068,N_6232);
and U13939 (N_13939,N_6609,N_9254);
or U13940 (N_13940,N_6097,N_9525);
nand U13941 (N_13941,N_8304,N_6337);
xor U13942 (N_13942,N_7677,N_6778);
xor U13943 (N_13943,N_7961,N_7909);
and U13944 (N_13944,N_7072,N_7925);
and U13945 (N_13945,N_6585,N_6947);
nor U13946 (N_13946,N_7227,N_7195);
nand U13947 (N_13947,N_5519,N_5543);
and U13948 (N_13948,N_7418,N_9749);
and U13949 (N_13949,N_7939,N_9004);
nand U13950 (N_13950,N_5867,N_7699);
xor U13951 (N_13951,N_5412,N_9008);
nor U13952 (N_13952,N_9316,N_6710);
and U13953 (N_13953,N_6551,N_5235);
or U13954 (N_13954,N_7260,N_6760);
and U13955 (N_13955,N_5115,N_8981);
or U13956 (N_13956,N_6448,N_7712);
or U13957 (N_13957,N_7762,N_5130);
nor U13958 (N_13958,N_8148,N_9194);
or U13959 (N_13959,N_7851,N_8002);
nor U13960 (N_13960,N_7772,N_6268);
and U13961 (N_13961,N_6761,N_8584);
and U13962 (N_13962,N_6055,N_5067);
nor U13963 (N_13963,N_5424,N_5827);
nand U13964 (N_13964,N_6010,N_7711);
xor U13965 (N_13965,N_5633,N_6942);
nand U13966 (N_13966,N_9086,N_9479);
or U13967 (N_13967,N_9704,N_6945);
nand U13968 (N_13968,N_8575,N_5899);
nor U13969 (N_13969,N_8445,N_6082);
xor U13970 (N_13970,N_7032,N_6302);
xnor U13971 (N_13971,N_9017,N_5655);
nor U13972 (N_13972,N_8108,N_8006);
or U13973 (N_13973,N_5255,N_5256);
nand U13974 (N_13974,N_5604,N_5785);
nand U13975 (N_13975,N_7623,N_6632);
nor U13976 (N_13976,N_8884,N_6848);
or U13977 (N_13977,N_5297,N_7059);
and U13978 (N_13978,N_8606,N_9213);
xor U13979 (N_13979,N_5022,N_7804);
or U13980 (N_13980,N_6278,N_6610);
or U13981 (N_13981,N_8711,N_6062);
and U13982 (N_13982,N_9641,N_6646);
xor U13983 (N_13983,N_6778,N_7286);
xor U13984 (N_13984,N_8425,N_9335);
and U13985 (N_13985,N_7760,N_7875);
xnor U13986 (N_13986,N_8018,N_9598);
nor U13987 (N_13987,N_8448,N_6584);
xnor U13988 (N_13988,N_7197,N_6425);
xor U13989 (N_13989,N_7033,N_7518);
or U13990 (N_13990,N_9672,N_8210);
nor U13991 (N_13991,N_7324,N_9123);
xor U13992 (N_13992,N_6873,N_7769);
nor U13993 (N_13993,N_7498,N_8352);
and U13994 (N_13994,N_9909,N_8640);
xor U13995 (N_13995,N_6048,N_6763);
or U13996 (N_13996,N_5519,N_5447);
xnor U13997 (N_13997,N_6344,N_9481);
nor U13998 (N_13998,N_7102,N_9913);
xnor U13999 (N_13999,N_5424,N_6680);
nand U14000 (N_14000,N_9738,N_5988);
xnor U14001 (N_14001,N_5489,N_8444);
and U14002 (N_14002,N_5566,N_8938);
nor U14003 (N_14003,N_8607,N_5861);
xnor U14004 (N_14004,N_6760,N_8062);
nor U14005 (N_14005,N_9003,N_6171);
and U14006 (N_14006,N_6185,N_6259);
xor U14007 (N_14007,N_9989,N_6184);
nor U14008 (N_14008,N_5168,N_7749);
nand U14009 (N_14009,N_8586,N_6508);
nand U14010 (N_14010,N_9672,N_6995);
xnor U14011 (N_14011,N_8125,N_7301);
nor U14012 (N_14012,N_7987,N_7033);
xnor U14013 (N_14013,N_7918,N_8963);
or U14014 (N_14014,N_9162,N_8817);
or U14015 (N_14015,N_8090,N_9189);
or U14016 (N_14016,N_8657,N_5094);
xor U14017 (N_14017,N_5738,N_8203);
nor U14018 (N_14018,N_8240,N_9738);
nand U14019 (N_14019,N_5354,N_7887);
and U14020 (N_14020,N_7119,N_7352);
and U14021 (N_14021,N_6393,N_5699);
or U14022 (N_14022,N_8223,N_8893);
or U14023 (N_14023,N_6037,N_8146);
nand U14024 (N_14024,N_9763,N_7752);
xnor U14025 (N_14025,N_7927,N_5573);
or U14026 (N_14026,N_6868,N_9678);
or U14027 (N_14027,N_9830,N_5314);
nand U14028 (N_14028,N_5793,N_6411);
nor U14029 (N_14029,N_7221,N_7167);
and U14030 (N_14030,N_8582,N_9955);
nor U14031 (N_14031,N_5034,N_8168);
xor U14032 (N_14032,N_7970,N_6108);
nand U14033 (N_14033,N_7533,N_9697);
xnor U14034 (N_14034,N_5380,N_8905);
nand U14035 (N_14035,N_5053,N_6841);
and U14036 (N_14036,N_8535,N_6726);
or U14037 (N_14037,N_8189,N_6892);
or U14038 (N_14038,N_8612,N_8909);
or U14039 (N_14039,N_8017,N_7594);
nand U14040 (N_14040,N_5675,N_5414);
and U14041 (N_14041,N_8446,N_8226);
nand U14042 (N_14042,N_9220,N_5298);
or U14043 (N_14043,N_7828,N_8123);
xor U14044 (N_14044,N_8262,N_6155);
nor U14045 (N_14045,N_9866,N_9023);
and U14046 (N_14046,N_6257,N_6957);
and U14047 (N_14047,N_7773,N_8926);
and U14048 (N_14048,N_7069,N_6305);
or U14049 (N_14049,N_9258,N_7811);
or U14050 (N_14050,N_6151,N_9935);
nor U14051 (N_14051,N_5183,N_8869);
or U14052 (N_14052,N_9920,N_6561);
nor U14053 (N_14053,N_7510,N_6934);
xor U14054 (N_14054,N_8799,N_8113);
xnor U14055 (N_14055,N_5907,N_8134);
xnor U14056 (N_14056,N_5710,N_7547);
nor U14057 (N_14057,N_5058,N_7080);
xnor U14058 (N_14058,N_9075,N_5135);
and U14059 (N_14059,N_6890,N_8897);
nor U14060 (N_14060,N_9226,N_9509);
and U14061 (N_14061,N_5670,N_7183);
xnor U14062 (N_14062,N_7011,N_8992);
nor U14063 (N_14063,N_8594,N_5110);
nand U14064 (N_14064,N_9600,N_8071);
xor U14065 (N_14065,N_6752,N_6468);
xor U14066 (N_14066,N_7178,N_7798);
xor U14067 (N_14067,N_5131,N_5447);
xnor U14068 (N_14068,N_7397,N_9566);
nand U14069 (N_14069,N_8152,N_8636);
nor U14070 (N_14070,N_7259,N_6022);
nand U14071 (N_14071,N_7948,N_8222);
xor U14072 (N_14072,N_6714,N_7282);
xor U14073 (N_14073,N_5474,N_9986);
nor U14074 (N_14074,N_5212,N_6775);
and U14075 (N_14075,N_7882,N_9109);
xor U14076 (N_14076,N_6380,N_5328);
nand U14077 (N_14077,N_5060,N_6786);
xor U14078 (N_14078,N_5814,N_5621);
and U14079 (N_14079,N_6810,N_7051);
nand U14080 (N_14080,N_8332,N_9999);
xor U14081 (N_14081,N_6170,N_6311);
or U14082 (N_14082,N_5373,N_5630);
xor U14083 (N_14083,N_7500,N_6351);
xnor U14084 (N_14084,N_8646,N_8387);
and U14085 (N_14085,N_6172,N_6990);
xnor U14086 (N_14086,N_8422,N_9881);
xnor U14087 (N_14087,N_7563,N_7704);
nand U14088 (N_14088,N_8257,N_5610);
or U14089 (N_14089,N_7884,N_5235);
nand U14090 (N_14090,N_6158,N_8300);
nor U14091 (N_14091,N_5695,N_6720);
nand U14092 (N_14092,N_5010,N_9891);
or U14093 (N_14093,N_9244,N_9574);
and U14094 (N_14094,N_8880,N_9252);
xnor U14095 (N_14095,N_8990,N_6917);
and U14096 (N_14096,N_5500,N_9279);
and U14097 (N_14097,N_8158,N_9806);
or U14098 (N_14098,N_8072,N_6824);
and U14099 (N_14099,N_8306,N_7608);
nand U14100 (N_14100,N_8830,N_7198);
nor U14101 (N_14101,N_7826,N_9234);
or U14102 (N_14102,N_6629,N_9294);
xor U14103 (N_14103,N_5756,N_5180);
nand U14104 (N_14104,N_7688,N_9233);
or U14105 (N_14105,N_9219,N_5626);
xnor U14106 (N_14106,N_5940,N_6826);
or U14107 (N_14107,N_5764,N_8008);
or U14108 (N_14108,N_9435,N_6891);
nand U14109 (N_14109,N_8531,N_8285);
nor U14110 (N_14110,N_5147,N_8571);
and U14111 (N_14111,N_6015,N_7877);
xor U14112 (N_14112,N_8227,N_7827);
nor U14113 (N_14113,N_7803,N_5625);
xnor U14114 (N_14114,N_6982,N_8211);
and U14115 (N_14115,N_6527,N_7183);
and U14116 (N_14116,N_6524,N_6472);
xnor U14117 (N_14117,N_5079,N_6138);
and U14118 (N_14118,N_7127,N_5779);
or U14119 (N_14119,N_5751,N_5802);
or U14120 (N_14120,N_7102,N_5047);
and U14121 (N_14121,N_8233,N_9689);
and U14122 (N_14122,N_7190,N_7760);
and U14123 (N_14123,N_8422,N_6221);
xnor U14124 (N_14124,N_6604,N_8413);
nand U14125 (N_14125,N_7560,N_5589);
or U14126 (N_14126,N_5094,N_5130);
or U14127 (N_14127,N_7291,N_5812);
or U14128 (N_14128,N_6621,N_6409);
nor U14129 (N_14129,N_6032,N_8635);
nor U14130 (N_14130,N_6429,N_6814);
or U14131 (N_14131,N_7183,N_5347);
nand U14132 (N_14132,N_8839,N_9281);
nor U14133 (N_14133,N_6118,N_7861);
nor U14134 (N_14134,N_9467,N_5218);
nor U14135 (N_14135,N_9136,N_7191);
and U14136 (N_14136,N_5285,N_6632);
and U14137 (N_14137,N_7186,N_9467);
and U14138 (N_14138,N_8988,N_6209);
or U14139 (N_14139,N_5419,N_8604);
xor U14140 (N_14140,N_8791,N_9593);
and U14141 (N_14141,N_8417,N_9517);
nor U14142 (N_14142,N_9131,N_9838);
nor U14143 (N_14143,N_7116,N_5429);
xor U14144 (N_14144,N_7608,N_6931);
or U14145 (N_14145,N_6461,N_8130);
nand U14146 (N_14146,N_7673,N_8478);
nand U14147 (N_14147,N_5587,N_5640);
nand U14148 (N_14148,N_6291,N_6916);
xnor U14149 (N_14149,N_8910,N_8747);
xnor U14150 (N_14150,N_5795,N_9002);
and U14151 (N_14151,N_5654,N_7421);
or U14152 (N_14152,N_6897,N_8452);
xnor U14153 (N_14153,N_8139,N_5625);
or U14154 (N_14154,N_5083,N_7903);
nand U14155 (N_14155,N_5895,N_5602);
nor U14156 (N_14156,N_7144,N_6003);
nor U14157 (N_14157,N_9646,N_9279);
xnor U14158 (N_14158,N_8342,N_9539);
nand U14159 (N_14159,N_8261,N_7437);
and U14160 (N_14160,N_8750,N_6678);
nor U14161 (N_14161,N_5023,N_5166);
nor U14162 (N_14162,N_7202,N_8049);
nand U14163 (N_14163,N_7764,N_7592);
nand U14164 (N_14164,N_7521,N_9486);
and U14165 (N_14165,N_5741,N_5256);
nand U14166 (N_14166,N_5781,N_9323);
or U14167 (N_14167,N_6255,N_9489);
and U14168 (N_14168,N_6934,N_9226);
xnor U14169 (N_14169,N_7602,N_7832);
or U14170 (N_14170,N_7622,N_6566);
nand U14171 (N_14171,N_5077,N_9569);
nor U14172 (N_14172,N_8329,N_6137);
xnor U14173 (N_14173,N_8821,N_7982);
or U14174 (N_14174,N_5407,N_8746);
and U14175 (N_14175,N_7207,N_6794);
nand U14176 (N_14176,N_5547,N_8176);
nand U14177 (N_14177,N_9469,N_6766);
and U14178 (N_14178,N_7120,N_7746);
nor U14179 (N_14179,N_9221,N_7998);
and U14180 (N_14180,N_8152,N_9925);
nor U14181 (N_14181,N_8132,N_6702);
or U14182 (N_14182,N_8083,N_8071);
nor U14183 (N_14183,N_5490,N_5491);
or U14184 (N_14184,N_5468,N_8344);
xnor U14185 (N_14185,N_8098,N_5260);
and U14186 (N_14186,N_5133,N_5334);
nor U14187 (N_14187,N_8378,N_7933);
nand U14188 (N_14188,N_7230,N_9880);
nand U14189 (N_14189,N_6165,N_9289);
nand U14190 (N_14190,N_5600,N_8399);
xnor U14191 (N_14191,N_6328,N_5970);
and U14192 (N_14192,N_9688,N_8013);
or U14193 (N_14193,N_5347,N_9677);
and U14194 (N_14194,N_8956,N_9101);
and U14195 (N_14195,N_8228,N_6697);
and U14196 (N_14196,N_7053,N_6562);
xor U14197 (N_14197,N_7427,N_6454);
nor U14198 (N_14198,N_9401,N_7947);
nand U14199 (N_14199,N_8429,N_9881);
xnor U14200 (N_14200,N_5251,N_5952);
nand U14201 (N_14201,N_5362,N_8854);
or U14202 (N_14202,N_8729,N_6721);
nor U14203 (N_14203,N_7679,N_6943);
or U14204 (N_14204,N_8597,N_9753);
or U14205 (N_14205,N_5019,N_9733);
nand U14206 (N_14206,N_5254,N_5983);
nor U14207 (N_14207,N_8837,N_6160);
nor U14208 (N_14208,N_9801,N_6138);
nor U14209 (N_14209,N_5537,N_5881);
or U14210 (N_14210,N_5199,N_7999);
and U14211 (N_14211,N_9120,N_5135);
or U14212 (N_14212,N_7259,N_9282);
or U14213 (N_14213,N_7980,N_6133);
and U14214 (N_14214,N_5644,N_5208);
nand U14215 (N_14215,N_6487,N_5088);
or U14216 (N_14216,N_5359,N_7337);
xor U14217 (N_14217,N_9144,N_9833);
and U14218 (N_14218,N_5728,N_8286);
or U14219 (N_14219,N_5333,N_8210);
nor U14220 (N_14220,N_9019,N_5328);
xnor U14221 (N_14221,N_8856,N_9170);
nand U14222 (N_14222,N_5184,N_5474);
nor U14223 (N_14223,N_6055,N_6312);
xnor U14224 (N_14224,N_9145,N_8692);
and U14225 (N_14225,N_9609,N_7291);
or U14226 (N_14226,N_5661,N_7815);
xnor U14227 (N_14227,N_7712,N_9769);
xnor U14228 (N_14228,N_6644,N_5374);
nor U14229 (N_14229,N_5706,N_7837);
nor U14230 (N_14230,N_9932,N_8587);
xor U14231 (N_14231,N_8956,N_6790);
or U14232 (N_14232,N_8143,N_6153);
nor U14233 (N_14233,N_5172,N_6865);
and U14234 (N_14234,N_8310,N_8730);
and U14235 (N_14235,N_5760,N_8175);
xor U14236 (N_14236,N_8627,N_7801);
xor U14237 (N_14237,N_5957,N_9991);
nand U14238 (N_14238,N_5391,N_5049);
nand U14239 (N_14239,N_6449,N_6720);
nor U14240 (N_14240,N_8304,N_7375);
and U14241 (N_14241,N_5523,N_9003);
xor U14242 (N_14242,N_8667,N_7474);
and U14243 (N_14243,N_6576,N_7626);
nor U14244 (N_14244,N_9880,N_6110);
nand U14245 (N_14245,N_8440,N_8916);
nand U14246 (N_14246,N_5273,N_9790);
xor U14247 (N_14247,N_9137,N_6787);
nor U14248 (N_14248,N_9772,N_8559);
xnor U14249 (N_14249,N_8012,N_6010);
xnor U14250 (N_14250,N_8112,N_7274);
nand U14251 (N_14251,N_7544,N_7419);
xor U14252 (N_14252,N_5139,N_5003);
or U14253 (N_14253,N_5849,N_7567);
nor U14254 (N_14254,N_5102,N_7024);
or U14255 (N_14255,N_7610,N_6797);
or U14256 (N_14256,N_7296,N_8381);
nor U14257 (N_14257,N_9835,N_5254);
or U14258 (N_14258,N_5685,N_9904);
or U14259 (N_14259,N_5103,N_9192);
xor U14260 (N_14260,N_6166,N_6165);
and U14261 (N_14261,N_5718,N_8476);
and U14262 (N_14262,N_6668,N_5450);
nand U14263 (N_14263,N_6817,N_8870);
and U14264 (N_14264,N_6104,N_8535);
and U14265 (N_14265,N_8574,N_6086);
nand U14266 (N_14266,N_8428,N_5621);
nand U14267 (N_14267,N_5182,N_6909);
xnor U14268 (N_14268,N_6890,N_6015);
or U14269 (N_14269,N_7799,N_8356);
xor U14270 (N_14270,N_7940,N_8788);
xor U14271 (N_14271,N_9015,N_9677);
xnor U14272 (N_14272,N_9468,N_7650);
xnor U14273 (N_14273,N_7295,N_6474);
or U14274 (N_14274,N_5334,N_6293);
or U14275 (N_14275,N_9024,N_5380);
and U14276 (N_14276,N_6873,N_8952);
or U14277 (N_14277,N_8661,N_8037);
nor U14278 (N_14278,N_5342,N_7366);
nor U14279 (N_14279,N_7258,N_6508);
nor U14280 (N_14280,N_7059,N_6814);
xnor U14281 (N_14281,N_7474,N_8629);
or U14282 (N_14282,N_9354,N_7060);
or U14283 (N_14283,N_6266,N_8400);
nand U14284 (N_14284,N_6749,N_6743);
nor U14285 (N_14285,N_5103,N_5238);
nand U14286 (N_14286,N_9282,N_7457);
nand U14287 (N_14287,N_9030,N_5626);
nor U14288 (N_14288,N_5071,N_6473);
nand U14289 (N_14289,N_6653,N_7532);
and U14290 (N_14290,N_5440,N_8815);
and U14291 (N_14291,N_7897,N_6503);
and U14292 (N_14292,N_8306,N_6057);
nand U14293 (N_14293,N_9923,N_7985);
or U14294 (N_14294,N_9794,N_9223);
and U14295 (N_14295,N_5818,N_8251);
and U14296 (N_14296,N_9518,N_9407);
xnor U14297 (N_14297,N_8825,N_7885);
and U14298 (N_14298,N_7492,N_6532);
nand U14299 (N_14299,N_8658,N_9475);
nand U14300 (N_14300,N_8785,N_9423);
nor U14301 (N_14301,N_8487,N_8287);
or U14302 (N_14302,N_7157,N_5197);
and U14303 (N_14303,N_8349,N_5879);
or U14304 (N_14304,N_5702,N_7003);
xnor U14305 (N_14305,N_8464,N_5592);
or U14306 (N_14306,N_9950,N_9021);
xor U14307 (N_14307,N_7794,N_9512);
and U14308 (N_14308,N_7215,N_9155);
and U14309 (N_14309,N_5310,N_6559);
and U14310 (N_14310,N_6613,N_8990);
xnor U14311 (N_14311,N_7460,N_5510);
and U14312 (N_14312,N_5754,N_9715);
or U14313 (N_14313,N_9225,N_6388);
or U14314 (N_14314,N_8337,N_6198);
nor U14315 (N_14315,N_8602,N_8144);
or U14316 (N_14316,N_6336,N_9114);
xor U14317 (N_14317,N_5641,N_6960);
and U14318 (N_14318,N_5162,N_9746);
and U14319 (N_14319,N_7573,N_8917);
xor U14320 (N_14320,N_5600,N_9815);
or U14321 (N_14321,N_8322,N_8646);
or U14322 (N_14322,N_5456,N_7765);
and U14323 (N_14323,N_7795,N_5403);
xnor U14324 (N_14324,N_7664,N_6405);
and U14325 (N_14325,N_8263,N_9287);
or U14326 (N_14326,N_8226,N_9308);
xnor U14327 (N_14327,N_5360,N_8180);
or U14328 (N_14328,N_9922,N_9087);
or U14329 (N_14329,N_5749,N_7681);
xor U14330 (N_14330,N_8478,N_7338);
xor U14331 (N_14331,N_5401,N_6416);
and U14332 (N_14332,N_5505,N_5066);
nand U14333 (N_14333,N_8582,N_7692);
nor U14334 (N_14334,N_6290,N_7419);
nor U14335 (N_14335,N_7614,N_8798);
and U14336 (N_14336,N_8620,N_8072);
nand U14337 (N_14337,N_8599,N_5761);
xor U14338 (N_14338,N_7028,N_6662);
and U14339 (N_14339,N_7580,N_9688);
or U14340 (N_14340,N_8816,N_7291);
nand U14341 (N_14341,N_9930,N_6882);
and U14342 (N_14342,N_9789,N_7748);
xor U14343 (N_14343,N_9258,N_8478);
or U14344 (N_14344,N_9995,N_8998);
and U14345 (N_14345,N_6536,N_9544);
or U14346 (N_14346,N_7640,N_9994);
xor U14347 (N_14347,N_7990,N_8654);
nor U14348 (N_14348,N_8184,N_8975);
and U14349 (N_14349,N_9032,N_5460);
nor U14350 (N_14350,N_7256,N_6100);
and U14351 (N_14351,N_5598,N_5896);
nand U14352 (N_14352,N_8307,N_5985);
xnor U14353 (N_14353,N_6457,N_6562);
or U14354 (N_14354,N_5399,N_8352);
nor U14355 (N_14355,N_7731,N_8230);
nor U14356 (N_14356,N_9402,N_9542);
xor U14357 (N_14357,N_5241,N_9430);
nor U14358 (N_14358,N_8963,N_5904);
xor U14359 (N_14359,N_7506,N_5479);
xnor U14360 (N_14360,N_7903,N_7253);
xor U14361 (N_14361,N_9561,N_8637);
or U14362 (N_14362,N_6155,N_7097);
xor U14363 (N_14363,N_6363,N_9048);
xor U14364 (N_14364,N_5021,N_7423);
or U14365 (N_14365,N_5903,N_5007);
nor U14366 (N_14366,N_5721,N_9109);
nor U14367 (N_14367,N_8565,N_8673);
nand U14368 (N_14368,N_7799,N_5135);
xnor U14369 (N_14369,N_5910,N_7228);
nor U14370 (N_14370,N_9499,N_5526);
nor U14371 (N_14371,N_9588,N_5002);
nor U14372 (N_14372,N_8148,N_5469);
and U14373 (N_14373,N_7887,N_7503);
and U14374 (N_14374,N_5345,N_7127);
nor U14375 (N_14375,N_9396,N_7093);
nand U14376 (N_14376,N_5600,N_8921);
or U14377 (N_14377,N_7239,N_5204);
nor U14378 (N_14378,N_5524,N_5759);
nand U14379 (N_14379,N_9842,N_7597);
nand U14380 (N_14380,N_9527,N_9818);
and U14381 (N_14381,N_7516,N_6603);
or U14382 (N_14382,N_9004,N_7232);
nand U14383 (N_14383,N_7284,N_5641);
nand U14384 (N_14384,N_7443,N_6689);
or U14385 (N_14385,N_8539,N_7901);
and U14386 (N_14386,N_7407,N_7801);
nand U14387 (N_14387,N_6746,N_5740);
nand U14388 (N_14388,N_8138,N_5402);
xor U14389 (N_14389,N_6540,N_6584);
nand U14390 (N_14390,N_9254,N_6181);
nor U14391 (N_14391,N_6200,N_8905);
xor U14392 (N_14392,N_9691,N_8069);
or U14393 (N_14393,N_5930,N_9466);
nor U14394 (N_14394,N_8457,N_9980);
and U14395 (N_14395,N_7522,N_6046);
and U14396 (N_14396,N_9646,N_8075);
nor U14397 (N_14397,N_9605,N_6531);
and U14398 (N_14398,N_6522,N_8920);
or U14399 (N_14399,N_8872,N_7731);
and U14400 (N_14400,N_9010,N_7668);
nand U14401 (N_14401,N_9711,N_8984);
or U14402 (N_14402,N_7848,N_8914);
or U14403 (N_14403,N_5805,N_8240);
xnor U14404 (N_14404,N_9259,N_6780);
xnor U14405 (N_14405,N_8513,N_7703);
or U14406 (N_14406,N_8582,N_5597);
or U14407 (N_14407,N_9852,N_7996);
xnor U14408 (N_14408,N_8724,N_6428);
xnor U14409 (N_14409,N_5731,N_8354);
or U14410 (N_14410,N_8208,N_8437);
or U14411 (N_14411,N_6271,N_5641);
xnor U14412 (N_14412,N_5699,N_8067);
xnor U14413 (N_14413,N_5250,N_5678);
and U14414 (N_14414,N_9935,N_6186);
nor U14415 (N_14415,N_6214,N_8308);
nand U14416 (N_14416,N_5952,N_7822);
nand U14417 (N_14417,N_9000,N_9736);
nand U14418 (N_14418,N_7890,N_5804);
or U14419 (N_14419,N_8393,N_5446);
nor U14420 (N_14420,N_9288,N_6954);
nor U14421 (N_14421,N_6094,N_9852);
nor U14422 (N_14422,N_9526,N_9441);
or U14423 (N_14423,N_8274,N_8162);
or U14424 (N_14424,N_6589,N_6894);
xnor U14425 (N_14425,N_7486,N_8856);
nand U14426 (N_14426,N_6499,N_6011);
xnor U14427 (N_14427,N_7072,N_9002);
or U14428 (N_14428,N_9569,N_8678);
or U14429 (N_14429,N_8721,N_9724);
and U14430 (N_14430,N_8261,N_7673);
or U14431 (N_14431,N_5273,N_9443);
nor U14432 (N_14432,N_6609,N_7543);
or U14433 (N_14433,N_5054,N_5924);
xor U14434 (N_14434,N_6089,N_8779);
nand U14435 (N_14435,N_7691,N_8659);
xor U14436 (N_14436,N_5550,N_7016);
or U14437 (N_14437,N_8304,N_9187);
nand U14438 (N_14438,N_5845,N_8459);
nand U14439 (N_14439,N_5606,N_8881);
and U14440 (N_14440,N_6248,N_6990);
and U14441 (N_14441,N_9217,N_6564);
nand U14442 (N_14442,N_5942,N_8497);
nor U14443 (N_14443,N_6763,N_6170);
xor U14444 (N_14444,N_8533,N_6978);
or U14445 (N_14445,N_6064,N_8256);
nand U14446 (N_14446,N_6380,N_5747);
xor U14447 (N_14447,N_5690,N_5237);
xnor U14448 (N_14448,N_6043,N_5197);
and U14449 (N_14449,N_8065,N_6032);
nor U14450 (N_14450,N_9260,N_8774);
xnor U14451 (N_14451,N_8325,N_5438);
xnor U14452 (N_14452,N_5085,N_9757);
nand U14453 (N_14453,N_7286,N_7155);
xnor U14454 (N_14454,N_5853,N_9260);
nand U14455 (N_14455,N_5892,N_6245);
xnor U14456 (N_14456,N_8035,N_5891);
nor U14457 (N_14457,N_6936,N_5186);
nor U14458 (N_14458,N_7446,N_7986);
nand U14459 (N_14459,N_6225,N_9736);
or U14460 (N_14460,N_5850,N_8292);
or U14461 (N_14461,N_5469,N_6126);
nand U14462 (N_14462,N_8689,N_8148);
or U14463 (N_14463,N_5599,N_7803);
xor U14464 (N_14464,N_5158,N_7893);
and U14465 (N_14465,N_9223,N_6486);
nand U14466 (N_14466,N_6492,N_9035);
nand U14467 (N_14467,N_8247,N_5586);
or U14468 (N_14468,N_7522,N_7587);
nor U14469 (N_14469,N_5332,N_8918);
nor U14470 (N_14470,N_7321,N_6231);
nor U14471 (N_14471,N_6276,N_6480);
xor U14472 (N_14472,N_7879,N_6017);
or U14473 (N_14473,N_8868,N_5724);
or U14474 (N_14474,N_6586,N_8325);
or U14475 (N_14475,N_5844,N_5567);
xnor U14476 (N_14476,N_8070,N_7976);
and U14477 (N_14477,N_5035,N_6663);
xor U14478 (N_14478,N_8895,N_8130);
nor U14479 (N_14479,N_6989,N_6239);
nand U14480 (N_14480,N_8259,N_6693);
or U14481 (N_14481,N_7964,N_7644);
xnor U14482 (N_14482,N_9148,N_6404);
or U14483 (N_14483,N_8090,N_8727);
and U14484 (N_14484,N_8507,N_9365);
and U14485 (N_14485,N_8893,N_7582);
nand U14486 (N_14486,N_8742,N_9923);
and U14487 (N_14487,N_5409,N_6437);
nor U14488 (N_14488,N_5487,N_5575);
or U14489 (N_14489,N_9473,N_5215);
xnor U14490 (N_14490,N_6787,N_7111);
nand U14491 (N_14491,N_7605,N_5579);
and U14492 (N_14492,N_9017,N_7906);
and U14493 (N_14493,N_7972,N_9544);
and U14494 (N_14494,N_5596,N_6436);
nand U14495 (N_14495,N_6772,N_9654);
and U14496 (N_14496,N_8342,N_9706);
nand U14497 (N_14497,N_6118,N_9962);
nor U14498 (N_14498,N_5444,N_6992);
nand U14499 (N_14499,N_5335,N_8828);
and U14500 (N_14500,N_8996,N_6812);
xor U14501 (N_14501,N_8091,N_8658);
or U14502 (N_14502,N_8575,N_6416);
xor U14503 (N_14503,N_9376,N_8238);
nand U14504 (N_14504,N_5546,N_5575);
xor U14505 (N_14505,N_8720,N_8330);
or U14506 (N_14506,N_7158,N_9983);
nor U14507 (N_14507,N_8161,N_5036);
xor U14508 (N_14508,N_9335,N_5021);
and U14509 (N_14509,N_6188,N_8774);
and U14510 (N_14510,N_6136,N_9143);
xor U14511 (N_14511,N_5213,N_9111);
or U14512 (N_14512,N_5928,N_6582);
nand U14513 (N_14513,N_8155,N_8245);
or U14514 (N_14514,N_8024,N_6511);
and U14515 (N_14515,N_9165,N_7947);
xnor U14516 (N_14516,N_9619,N_9177);
or U14517 (N_14517,N_7368,N_5265);
or U14518 (N_14518,N_9490,N_8183);
nor U14519 (N_14519,N_7229,N_6165);
nor U14520 (N_14520,N_6773,N_5772);
and U14521 (N_14521,N_7835,N_5573);
and U14522 (N_14522,N_9832,N_5635);
nor U14523 (N_14523,N_9317,N_7967);
or U14524 (N_14524,N_9877,N_7604);
nor U14525 (N_14525,N_7329,N_6924);
xor U14526 (N_14526,N_9702,N_9643);
or U14527 (N_14527,N_6785,N_9113);
and U14528 (N_14528,N_5501,N_7970);
and U14529 (N_14529,N_5059,N_5646);
nand U14530 (N_14530,N_8635,N_8479);
and U14531 (N_14531,N_8298,N_7100);
and U14532 (N_14532,N_8038,N_9549);
nor U14533 (N_14533,N_6703,N_5160);
and U14534 (N_14534,N_9572,N_7052);
and U14535 (N_14535,N_6180,N_8165);
nand U14536 (N_14536,N_5458,N_7260);
nor U14537 (N_14537,N_9292,N_9882);
and U14538 (N_14538,N_7273,N_7180);
or U14539 (N_14539,N_9644,N_9132);
nand U14540 (N_14540,N_5716,N_5591);
or U14541 (N_14541,N_9007,N_7742);
and U14542 (N_14542,N_5276,N_9284);
xnor U14543 (N_14543,N_7812,N_6791);
xnor U14544 (N_14544,N_9196,N_7389);
and U14545 (N_14545,N_5825,N_8570);
and U14546 (N_14546,N_7867,N_5036);
or U14547 (N_14547,N_9314,N_8266);
xnor U14548 (N_14548,N_9572,N_8068);
and U14549 (N_14549,N_6826,N_7831);
nor U14550 (N_14550,N_8209,N_7016);
or U14551 (N_14551,N_9611,N_8872);
and U14552 (N_14552,N_7343,N_8746);
xor U14553 (N_14553,N_9891,N_6501);
and U14554 (N_14554,N_7735,N_7830);
or U14555 (N_14555,N_9646,N_8248);
xnor U14556 (N_14556,N_6419,N_6900);
xor U14557 (N_14557,N_7841,N_9476);
nand U14558 (N_14558,N_8593,N_8992);
nand U14559 (N_14559,N_8293,N_5733);
and U14560 (N_14560,N_6276,N_6851);
or U14561 (N_14561,N_6117,N_7202);
nor U14562 (N_14562,N_9302,N_6539);
xnor U14563 (N_14563,N_5039,N_6131);
or U14564 (N_14564,N_8554,N_8825);
and U14565 (N_14565,N_5791,N_6671);
and U14566 (N_14566,N_7452,N_5408);
and U14567 (N_14567,N_5369,N_5924);
or U14568 (N_14568,N_9761,N_9885);
xor U14569 (N_14569,N_7596,N_7152);
or U14570 (N_14570,N_6095,N_7067);
xor U14571 (N_14571,N_5156,N_7925);
or U14572 (N_14572,N_5209,N_5133);
nor U14573 (N_14573,N_9143,N_9346);
xor U14574 (N_14574,N_7345,N_5181);
and U14575 (N_14575,N_6894,N_7227);
or U14576 (N_14576,N_6971,N_5151);
nand U14577 (N_14577,N_9294,N_7785);
nor U14578 (N_14578,N_8240,N_9441);
nor U14579 (N_14579,N_6962,N_7935);
nor U14580 (N_14580,N_7197,N_6265);
nor U14581 (N_14581,N_8792,N_6038);
xor U14582 (N_14582,N_7027,N_7551);
and U14583 (N_14583,N_8727,N_9389);
xnor U14584 (N_14584,N_9284,N_9334);
and U14585 (N_14585,N_7631,N_5007);
xnor U14586 (N_14586,N_6600,N_6680);
and U14587 (N_14587,N_7373,N_9066);
nand U14588 (N_14588,N_7356,N_8616);
and U14589 (N_14589,N_6198,N_6764);
and U14590 (N_14590,N_7081,N_5858);
xnor U14591 (N_14591,N_9977,N_7793);
xor U14592 (N_14592,N_7491,N_8722);
or U14593 (N_14593,N_6881,N_9608);
or U14594 (N_14594,N_6874,N_5127);
or U14595 (N_14595,N_8267,N_8848);
xor U14596 (N_14596,N_8196,N_9579);
nor U14597 (N_14597,N_7748,N_7723);
or U14598 (N_14598,N_8124,N_8711);
or U14599 (N_14599,N_6589,N_5715);
nor U14600 (N_14600,N_8819,N_6174);
nor U14601 (N_14601,N_5105,N_8978);
or U14602 (N_14602,N_8159,N_7456);
and U14603 (N_14603,N_6310,N_5514);
nand U14604 (N_14604,N_7645,N_9348);
or U14605 (N_14605,N_5663,N_6592);
nand U14606 (N_14606,N_6321,N_9350);
nand U14607 (N_14607,N_8928,N_7100);
xor U14608 (N_14608,N_5134,N_7376);
nand U14609 (N_14609,N_5166,N_7985);
and U14610 (N_14610,N_9782,N_9257);
nand U14611 (N_14611,N_9179,N_8004);
nand U14612 (N_14612,N_9367,N_5363);
or U14613 (N_14613,N_8626,N_7487);
or U14614 (N_14614,N_9812,N_5051);
or U14615 (N_14615,N_9488,N_5706);
xor U14616 (N_14616,N_6009,N_9162);
and U14617 (N_14617,N_8665,N_5567);
nor U14618 (N_14618,N_5634,N_5617);
or U14619 (N_14619,N_5765,N_9392);
nand U14620 (N_14620,N_5217,N_7206);
and U14621 (N_14621,N_9689,N_9519);
xor U14622 (N_14622,N_7250,N_9874);
nand U14623 (N_14623,N_7109,N_6004);
and U14624 (N_14624,N_6456,N_6895);
nand U14625 (N_14625,N_6714,N_7515);
or U14626 (N_14626,N_9406,N_5070);
or U14627 (N_14627,N_5713,N_5589);
nor U14628 (N_14628,N_8027,N_7121);
nor U14629 (N_14629,N_8049,N_8608);
nand U14630 (N_14630,N_7046,N_9683);
or U14631 (N_14631,N_7345,N_7098);
or U14632 (N_14632,N_6072,N_6318);
and U14633 (N_14633,N_8654,N_5333);
nor U14634 (N_14634,N_6258,N_5285);
and U14635 (N_14635,N_6057,N_8402);
nor U14636 (N_14636,N_6547,N_7017);
xor U14637 (N_14637,N_5818,N_6930);
nor U14638 (N_14638,N_8778,N_9553);
nor U14639 (N_14639,N_7567,N_8330);
and U14640 (N_14640,N_5578,N_8102);
xnor U14641 (N_14641,N_7231,N_9094);
and U14642 (N_14642,N_8563,N_5626);
or U14643 (N_14643,N_5598,N_8512);
and U14644 (N_14644,N_9284,N_8174);
or U14645 (N_14645,N_5048,N_8174);
or U14646 (N_14646,N_8348,N_5500);
xnor U14647 (N_14647,N_7470,N_6873);
nor U14648 (N_14648,N_9729,N_8263);
and U14649 (N_14649,N_8929,N_5360);
or U14650 (N_14650,N_7586,N_7180);
nand U14651 (N_14651,N_7087,N_8097);
nor U14652 (N_14652,N_8018,N_9486);
nand U14653 (N_14653,N_6479,N_6981);
nand U14654 (N_14654,N_6894,N_7910);
xor U14655 (N_14655,N_9674,N_8538);
nor U14656 (N_14656,N_6111,N_5595);
nor U14657 (N_14657,N_9910,N_6446);
xor U14658 (N_14658,N_7555,N_5949);
nor U14659 (N_14659,N_7554,N_9394);
nand U14660 (N_14660,N_6652,N_8520);
and U14661 (N_14661,N_5828,N_7490);
and U14662 (N_14662,N_7846,N_6703);
nor U14663 (N_14663,N_6471,N_9171);
or U14664 (N_14664,N_5259,N_8117);
and U14665 (N_14665,N_5020,N_9219);
or U14666 (N_14666,N_7739,N_6719);
and U14667 (N_14667,N_6040,N_6929);
and U14668 (N_14668,N_5343,N_6219);
nand U14669 (N_14669,N_9383,N_9400);
nand U14670 (N_14670,N_6065,N_6490);
nor U14671 (N_14671,N_7066,N_9531);
xor U14672 (N_14672,N_7849,N_9692);
or U14673 (N_14673,N_7809,N_6749);
nand U14674 (N_14674,N_8147,N_9715);
and U14675 (N_14675,N_7957,N_9413);
nor U14676 (N_14676,N_7464,N_8281);
or U14677 (N_14677,N_9449,N_6396);
nor U14678 (N_14678,N_9445,N_7559);
nand U14679 (N_14679,N_5138,N_6539);
xnor U14680 (N_14680,N_6135,N_6676);
and U14681 (N_14681,N_6236,N_5416);
xor U14682 (N_14682,N_7294,N_5507);
or U14683 (N_14683,N_5834,N_6319);
or U14684 (N_14684,N_9476,N_5714);
nor U14685 (N_14685,N_6104,N_9392);
nor U14686 (N_14686,N_7719,N_7020);
nand U14687 (N_14687,N_5849,N_9772);
and U14688 (N_14688,N_8185,N_6598);
nand U14689 (N_14689,N_7205,N_7416);
xor U14690 (N_14690,N_7854,N_7319);
xor U14691 (N_14691,N_5856,N_9527);
or U14692 (N_14692,N_7493,N_9035);
nand U14693 (N_14693,N_5478,N_5741);
nor U14694 (N_14694,N_8396,N_6629);
and U14695 (N_14695,N_7914,N_5575);
or U14696 (N_14696,N_6331,N_6008);
nand U14697 (N_14697,N_9869,N_7648);
nand U14698 (N_14698,N_9442,N_9553);
nor U14699 (N_14699,N_8914,N_9385);
nand U14700 (N_14700,N_7047,N_9750);
nand U14701 (N_14701,N_9513,N_8025);
nand U14702 (N_14702,N_7064,N_9596);
nor U14703 (N_14703,N_9097,N_6121);
nand U14704 (N_14704,N_8814,N_8205);
or U14705 (N_14705,N_6244,N_5650);
and U14706 (N_14706,N_5247,N_7921);
nand U14707 (N_14707,N_5515,N_8694);
or U14708 (N_14708,N_5735,N_6449);
and U14709 (N_14709,N_8034,N_6921);
nor U14710 (N_14710,N_5903,N_9063);
nand U14711 (N_14711,N_8478,N_6786);
nand U14712 (N_14712,N_8731,N_9418);
nand U14713 (N_14713,N_8967,N_9266);
xor U14714 (N_14714,N_6923,N_6403);
nor U14715 (N_14715,N_6505,N_5268);
or U14716 (N_14716,N_5031,N_8409);
or U14717 (N_14717,N_9411,N_7481);
nand U14718 (N_14718,N_6853,N_7380);
nor U14719 (N_14719,N_7057,N_7938);
nand U14720 (N_14720,N_6228,N_8053);
xnor U14721 (N_14721,N_7058,N_6739);
nor U14722 (N_14722,N_5717,N_6775);
xnor U14723 (N_14723,N_6010,N_5897);
or U14724 (N_14724,N_8750,N_6976);
and U14725 (N_14725,N_8592,N_7647);
nand U14726 (N_14726,N_6549,N_6444);
and U14727 (N_14727,N_9046,N_5278);
nor U14728 (N_14728,N_5987,N_8576);
nand U14729 (N_14729,N_7611,N_6555);
nand U14730 (N_14730,N_8272,N_7790);
and U14731 (N_14731,N_6988,N_5807);
xnor U14732 (N_14732,N_9706,N_9476);
nor U14733 (N_14733,N_7449,N_6486);
nor U14734 (N_14734,N_9131,N_6146);
xor U14735 (N_14735,N_7449,N_5207);
nor U14736 (N_14736,N_9899,N_7420);
or U14737 (N_14737,N_7165,N_6678);
and U14738 (N_14738,N_7727,N_7902);
and U14739 (N_14739,N_5942,N_5548);
nor U14740 (N_14740,N_7632,N_7412);
or U14741 (N_14741,N_7620,N_8065);
and U14742 (N_14742,N_6605,N_8638);
nor U14743 (N_14743,N_7398,N_8563);
xnor U14744 (N_14744,N_6448,N_6602);
xor U14745 (N_14745,N_9685,N_8381);
and U14746 (N_14746,N_7264,N_9173);
and U14747 (N_14747,N_5154,N_8422);
nand U14748 (N_14748,N_6358,N_5727);
nand U14749 (N_14749,N_6158,N_7568);
and U14750 (N_14750,N_8781,N_8340);
nor U14751 (N_14751,N_8916,N_6534);
nand U14752 (N_14752,N_6194,N_8566);
nor U14753 (N_14753,N_9605,N_9609);
nor U14754 (N_14754,N_9713,N_6228);
nor U14755 (N_14755,N_6642,N_5863);
and U14756 (N_14756,N_6541,N_7617);
nand U14757 (N_14757,N_7876,N_6502);
xnor U14758 (N_14758,N_6979,N_9630);
nand U14759 (N_14759,N_8895,N_5494);
nand U14760 (N_14760,N_6344,N_7674);
and U14761 (N_14761,N_9108,N_8842);
xnor U14762 (N_14762,N_7666,N_6109);
nand U14763 (N_14763,N_7804,N_6092);
and U14764 (N_14764,N_7487,N_7423);
and U14765 (N_14765,N_7126,N_8868);
xnor U14766 (N_14766,N_9794,N_8193);
xor U14767 (N_14767,N_5999,N_6123);
nand U14768 (N_14768,N_6677,N_6354);
nand U14769 (N_14769,N_7549,N_8879);
and U14770 (N_14770,N_6907,N_7760);
nor U14771 (N_14771,N_9943,N_7270);
xnor U14772 (N_14772,N_7517,N_9141);
and U14773 (N_14773,N_6026,N_6524);
or U14774 (N_14774,N_5897,N_5845);
xor U14775 (N_14775,N_7529,N_5586);
or U14776 (N_14776,N_8636,N_6854);
and U14777 (N_14777,N_9940,N_7824);
xor U14778 (N_14778,N_6709,N_6487);
or U14779 (N_14779,N_9073,N_5230);
nand U14780 (N_14780,N_7953,N_7496);
nor U14781 (N_14781,N_6906,N_7231);
and U14782 (N_14782,N_6055,N_6704);
nor U14783 (N_14783,N_7774,N_6492);
and U14784 (N_14784,N_7515,N_6721);
xnor U14785 (N_14785,N_5759,N_5614);
nor U14786 (N_14786,N_7587,N_9474);
or U14787 (N_14787,N_8624,N_5640);
xor U14788 (N_14788,N_6178,N_9404);
and U14789 (N_14789,N_8771,N_8895);
or U14790 (N_14790,N_8838,N_5517);
xnor U14791 (N_14791,N_5210,N_6481);
or U14792 (N_14792,N_9665,N_7473);
and U14793 (N_14793,N_9250,N_9846);
and U14794 (N_14794,N_6460,N_6504);
nor U14795 (N_14795,N_6980,N_8464);
nor U14796 (N_14796,N_5989,N_7982);
nor U14797 (N_14797,N_7168,N_5660);
nor U14798 (N_14798,N_5194,N_8304);
xnor U14799 (N_14799,N_9178,N_9657);
or U14800 (N_14800,N_9617,N_7125);
xnor U14801 (N_14801,N_9918,N_5451);
or U14802 (N_14802,N_9562,N_8220);
nand U14803 (N_14803,N_6057,N_8255);
xnor U14804 (N_14804,N_5801,N_6983);
nand U14805 (N_14805,N_6195,N_6061);
or U14806 (N_14806,N_8214,N_7644);
nand U14807 (N_14807,N_7898,N_6301);
xor U14808 (N_14808,N_7973,N_8964);
nor U14809 (N_14809,N_8012,N_5661);
and U14810 (N_14810,N_8584,N_6872);
nand U14811 (N_14811,N_8943,N_9236);
and U14812 (N_14812,N_9883,N_5518);
nor U14813 (N_14813,N_5365,N_9986);
and U14814 (N_14814,N_6923,N_9034);
nand U14815 (N_14815,N_9475,N_7394);
nand U14816 (N_14816,N_8705,N_5805);
or U14817 (N_14817,N_5849,N_9515);
nand U14818 (N_14818,N_6803,N_7056);
nand U14819 (N_14819,N_7403,N_6740);
xnor U14820 (N_14820,N_6930,N_8782);
and U14821 (N_14821,N_5290,N_8271);
and U14822 (N_14822,N_7564,N_9483);
and U14823 (N_14823,N_7052,N_8129);
nor U14824 (N_14824,N_6937,N_6312);
or U14825 (N_14825,N_9410,N_7629);
nand U14826 (N_14826,N_5269,N_6107);
and U14827 (N_14827,N_5650,N_5829);
xor U14828 (N_14828,N_5685,N_5195);
or U14829 (N_14829,N_8855,N_5036);
xnor U14830 (N_14830,N_6405,N_6259);
or U14831 (N_14831,N_6194,N_7228);
xor U14832 (N_14832,N_7645,N_6697);
or U14833 (N_14833,N_8219,N_5533);
nor U14834 (N_14834,N_5643,N_7490);
and U14835 (N_14835,N_5978,N_7998);
xnor U14836 (N_14836,N_5913,N_6643);
nor U14837 (N_14837,N_5709,N_5259);
xor U14838 (N_14838,N_5568,N_5823);
and U14839 (N_14839,N_8567,N_9056);
xnor U14840 (N_14840,N_7239,N_7060);
xnor U14841 (N_14841,N_7071,N_8275);
nand U14842 (N_14842,N_9465,N_7944);
nand U14843 (N_14843,N_6901,N_8118);
and U14844 (N_14844,N_6274,N_7818);
xor U14845 (N_14845,N_9896,N_6618);
or U14846 (N_14846,N_7208,N_7615);
nor U14847 (N_14847,N_5180,N_6847);
and U14848 (N_14848,N_9155,N_8146);
xnor U14849 (N_14849,N_7157,N_7843);
nor U14850 (N_14850,N_7625,N_6253);
nor U14851 (N_14851,N_9725,N_6112);
nand U14852 (N_14852,N_6242,N_5970);
or U14853 (N_14853,N_8174,N_9010);
or U14854 (N_14854,N_6411,N_8236);
nand U14855 (N_14855,N_5177,N_6046);
and U14856 (N_14856,N_5872,N_7513);
or U14857 (N_14857,N_9642,N_6918);
xor U14858 (N_14858,N_6242,N_9935);
nor U14859 (N_14859,N_6951,N_7401);
xor U14860 (N_14860,N_9029,N_5764);
xor U14861 (N_14861,N_6241,N_6651);
nand U14862 (N_14862,N_9962,N_7800);
nor U14863 (N_14863,N_5072,N_6139);
and U14864 (N_14864,N_9136,N_8105);
and U14865 (N_14865,N_5437,N_7260);
or U14866 (N_14866,N_9597,N_6590);
nand U14867 (N_14867,N_5681,N_7343);
or U14868 (N_14868,N_6685,N_8110);
or U14869 (N_14869,N_9298,N_9471);
or U14870 (N_14870,N_9841,N_6352);
nor U14871 (N_14871,N_7887,N_5899);
or U14872 (N_14872,N_7138,N_6627);
or U14873 (N_14873,N_9940,N_9309);
nor U14874 (N_14874,N_6285,N_8154);
and U14875 (N_14875,N_6888,N_5194);
and U14876 (N_14876,N_8965,N_5306);
and U14877 (N_14877,N_9024,N_8630);
nand U14878 (N_14878,N_6532,N_9671);
nor U14879 (N_14879,N_8907,N_8419);
nand U14880 (N_14880,N_7740,N_7624);
and U14881 (N_14881,N_5036,N_7293);
and U14882 (N_14882,N_5755,N_9951);
nor U14883 (N_14883,N_5490,N_8270);
nand U14884 (N_14884,N_7029,N_5422);
xor U14885 (N_14885,N_7504,N_8837);
nand U14886 (N_14886,N_9114,N_6548);
and U14887 (N_14887,N_9357,N_7302);
xnor U14888 (N_14888,N_8343,N_9448);
xor U14889 (N_14889,N_9772,N_7575);
xnor U14890 (N_14890,N_6177,N_5128);
xnor U14891 (N_14891,N_8807,N_6327);
nand U14892 (N_14892,N_5298,N_6086);
nor U14893 (N_14893,N_9121,N_8562);
nor U14894 (N_14894,N_6945,N_5372);
nor U14895 (N_14895,N_8023,N_8929);
and U14896 (N_14896,N_5972,N_9749);
or U14897 (N_14897,N_7777,N_8860);
xnor U14898 (N_14898,N_7876,N_6492);
or U14899 (N_14899,N_8811,N_6082);
and U14900 (N_14900,N_5989,N_9931);
and U14901 (N_14901,N_7336,N_5633);
nand U14902 (N_14902,N_5481,N_5291);
nor U14903 (N_14903,N_6585,N_5479);
xnor U14904 (N_14904,N_6627,N_6303);
and U14905 (N_14905,N_6867,N_6318);
nor U14906 (N_14906,N_6029,N_5357);
xnor U14907 (N_14907,N_9295,N_6532);
or U14908 (N_14908,N_8790,N_9269);
or U14909 (N_14909,N_7077,N_5686);
and U14910 (N_14910,N_6778,N_7776);
nor U14911 (N_14911,N_7012,N_9200);
nand U14912 (N_14912,N_5114,N_5449);
nand U14913 (N_14913,N_8038,N_9163);
nor U14914 (N_14914,N_9864,N_5442);
nand U14915 (N_14915,N_6991,N_6313);
or U14916 (N_14916,N_9763,N_9792);
and U14917 (N_14917,N_6880,N_5328);
or U14918 (N_14918,N_9969,N_6311);
nor U14919 (N_14919,N_7861,N_6718);
and U14920 (N_14920,N_7088,N_7406);
xor U14921 (N_14921,N_5177,N_5843);
and U14922 (N_14922,N_6182,N_5033);
or U14923 (N_14923,N_9536,N_7492);
xor U14924 (N_14924,N_7382,N_7363);
nand U14925 (N_14925,N_7302,N_7818);
nand U14926 (N_14926,N_7444,N_9118);
xnor U14927 (N_14927,N_5565,N_7933);
xnor U14928 (N_14928,N_6534,N_6443);
and U14929 (N_14929,N_9636,N_9583);
or U14930 (N_14930,N_6551,N_6632);
xor U14931 (N_14931,N_5420,N_5010);
or U14932 (N_14932,N_8526,N_8715);
xor U14933 (N_14933,N_5849,N_7938);
nor U14934 (N_14934,N_8185,N_9647);
nand U14935 (N_14935,N_8983,N_8617);
nand U14936 (N_14936,N_9282,N_7149);
xor U14937 (N_14937,N_8100,N_5537);
and U14938 (N_14938,N_6510,N_8840);
or U14939 (N_14939,N_5242,N_6472);
and U14940 (N_14940,N_7376,N_7540);
nor U14941 (N_14941,N_9331,N_9134);
and U14942 (N_14942,N_6406,N_8258);
and U14943 (N_14943,N_6295,N_8675);
and U14944 (N_14944,N_9196,N_6500);
or U14945 (N_14945,N_6576,N_5525);
nand U14946 (N_14946,N_7384,N_9369);
xnor U14947 (N_14947,N_7841,N_6431);
and U14948 (N_14948,N_7987,N_8553);
nor U14949 (N_14949,N_6709,N_5998);
xnor U14950 (N_14950,N_9555,N_5077);
nor U14951 (N_14951,N_9398,N_9005);
and U14952 (N_14952,N_5916,N_7326);
or U14953 (N_14953,N_9247,N_7341);
xnor U14954 (N_14954,N_6878,N_8252);
nor U14955 (N_14955,N_9702,N_5456);
and U14956 (N_14956,N_8563,N_8280);
or U14957 (N_14957,N_6112,N_9688);
nor U14958 (N_14958,N_7961,N_7185);
or U14959 (N_14959,N_6783,N_8045);
xor U14960 (N_14960,N_9393,N_5796);
xor U14961 (N_14961,N_7247,N_6285);
nand U14962 (N_14962,N_8998,N_5973);
nand U14963 (N_14963,N_9520,N_6570);
and U14964 (N_14964,N_5159,N_5038);
xor U14965 (N_14965,N_5889,N_7227);
nand U14966 (N_14966,N_8695,N_8143);
or U14967 (N_14967,N_7513,N_8525);
nor U14968 (N_14968,N_8900,N_7143);
xnor U14969 (N_14969,N_6324,N_6282);
nand U14970 (N_14970,N_6464,N_7138);
xnor U14971 (N_14971,N_9635,N_7357);
and U14972 (N_14972,N_8156,N_8633);
nand U14973 (N_14973,N_6550,N_5002);
xnor U14974 (N_14974,N_8509,N_6239);
nor U14975 (N_14975,N_7510,N_6619);
nand U14976 (N_14976,N_5279,N_9666);
or U14977 (N_14977,N_9858,N_5506);
xnor U14978 (N_14978,N_8319,N_5906);
and U14979 (N_14979,N_9558,N_8404);
and U14980 (N_14980,N_7107,N_9046);
and U14981 (N_14981,N_6198,N_8834);
nand U14982 (N_14982,N_5658,N_6389);
nor U14983 (N_14983,N_5122,N_8290);
nand U14984 (N_14984,N_8782,N_9012);
nor U14985 (N_14985,N_6465,N_5629);
nand U14986 (N_14986,N_5005,N_6280);
nor U14987 (N_14987,N_9511,N_5501);
and U14988 (N_14988,N_8046,N_8752);
xnor U14989 (N_14989,N_8172,N_5347);
nand U14990 (N_14990,N_6585,N_9869);
xor U14991 (N_14991,N_5798,N_9076);
xnor U14992 (N_14992,N_6104,N_5090);
xor U14993 (N_14993,N_7326,N_5478);
or U14994 (N_14994,N_8073,N_9823);
xor U14995 (N_14995,N_6847,N_8444);
nand U14996 (N_14996,N_7388,N_5062);
or U14997 (N_14997,N_6903,N_9768);
nand U14998 (N_14998,N_7444,N_6085);
and U14999 (N_14999,N_5526,N_8532);
and U15000 (N_15000,N_10890,N_11168);
and U15001 (N_15001,N_10129,N_10491);
and U15002 (N_15002,N_12853,N_14355);
and U15003 (N_15003,N_11274,N_13339);
nor U15004 (N_15004,N_12696,N_14100);
nand U15005 (N_15005,N_11703,N_10564);
xor U15006 (N_15006,N_10644,N_11591);
and U15007 (N_15007,N_11898,N_13288);
and U15008 (N_15008,N_14103,N_11905);
and U15009 (N_15009,N_12588,N_13388);
xor U15010 (N_15010,N_13332,N_12985);
or U15011 (N_15011,N_12287,N_14839);
nand U15012 (N_15012,N_14901,N_13928);
nand U15013 (N_15013,N_14395,N_12187);
xnor U15014 (N_15014,N_13913,N_13156);
nor U15015 (N_15015,N_14855,N_11345);
nor U15016 (N_15016,N_14835,N_13852);
nand U15017 (N_15017,N_14825,N_12317);
or U15018 (N_15018,N_14184,N_12977);
nor U15019 (N_15019,N_11137,N_10228);
xor U15020 (N_15020,N_13746,N_12153);
xor U15021 (N_15021,N_14612,N_10670);
or U15022 (N_15022,N_12382,N_10076);
or U15023 (N_15023,N_14974,N_12273);
and U15024 (N_15024,N_10763,N_14125);
xor U15025 (N_15025,N_11681,N_13540);
or U15026 (N_15026,N_13801,N_11027);
nand U15027 (N_15027,N_12099,N_10908);
or U15028 (N_15028,N_10771,N_11235);
nor U15029 (N_15029,N_14389,N_13935);
or U15030 (N_15030,N_14004,N_10579);
xor U15031 (N_15031,N_11881,N_10474);
or U15032 (N_15032,N_14200,N_11590);
and U15033 (N_15033,N_11577,N_14412);
nand U15034 (N_15034,N_14164,N_11192);
nor U15035 (N_15035,N_13849,N_14179);
and U15036 (N_15036,N_14312,N_11428);
xnor U15037 (N_15037,N_10599,N_12201);
or U15038 (N_15038,N_14665,N_13412);
nand U15039 (N_15039,N_13790,N_11349);
nor U15040 (N_15040,N_11822,N_11042);
and U15041 (N_15041,N_12510,N_13863);
xnor U15042 (N_15042,N_10745,N_14322);
nand U15043 (N_15043,N_14463,N_12930);
or U15044 (N_15044,N_12028,N_12620);
nor U15045 (N_15045,N_12193,N_10959);
and U15046 (N_15046,N_10071,N_13755);
nand U15047 (N_15047,N_10351,N_10999);
nand U15048 (N_15048,N_14811,N_10854);
xnor U15049 (N_15049,N_11105,N_13101);
and U15050 (N_15050,N_12136,N_11947);
or U15051 (N_15051,N_13393,N_11074);
nor U15052 (N_15052,N_13542,N_12227);
nor U15053 (N_15053,N_13291,N_14746);
xnor U15054 (N_15054,N_10832,N_10981);
and U15055 (N_15055,N_10399,N_14566);
nand U15056 (N_15056,N_11626,N_10460);
xnor U15057 (N_15057,N_14510,N_14236);
and U15058 (N_15058,N_11280,N_10609);
nor U15059 (N_15059,N_12018,N_12892);
xnor U15060 (N_15060,N_11330,N_12882);
and U15061 (N_15061,N_10493,N_14625);
or U15062 (N_15062,N_11773,N_11987);
xor U15063 (N_15063,N_11298,N_10398);
or U15064 (N_15064,N_14961,N_11009);
nor U15065 (N_15065,N_11524,N_10873);
or U15066 (N_15066,N_14754,N_11210);
xor U15067 (N_15067,N_14884,N_13691);
and U15068 (N_15068,N_14187,N_11996);
nand U15069 (N_15069,N_13279,N_10938);
and U15070 (N_15070,N_14947,N_14186);
or U15071 (N_15071,N_11112,N_13494);
xnor U15072 (N_15072,N_13606,N_12726);
or U15073 (N_15073,N_13251,N_12377);
nand U15074 (N_15074,N_11799,N_13953);
nand U15075 (N_15075,N_11225,N_10161);
or U15076 (N_15076,N_13845,N_13985);
nand U15077 (N_15077,N_14420,N_11648);
nor U15078 (N_15078,N_14789,N_12810);
and U15079 (N_15079,N_14304,N_11698);
nor U15080 (N_15080,N_12668,N_11529);
xor U15081 (N_15081,N_13757,N_13577);
xor U15082 (N_15082,N_13824,N_14558);
xnor U15083 (N_15083,N_11587,N_11823);
and U15084 (N_15084,N_12570,N_14969);
nand U15085 (N_15085,N_10887,N_13711);
nor U15086 (N_15086,N_11747,N_14272);
xor U15087 (N_15087,N_13196,N_12016);
or U15088 (N_15088,N_14020,N_11020);
nand U15089 (N_15089,N_10503,N_12653);
nor U15090 (N_15090,N_13965,N_12222);
or U15091 (N_15091,N_12071,N_10544);
or U15092 (N_15092,N_12143,N_14454);
nand U15093 (N_15093,N_11082,N_10377);
nor U15094 (N_15094,N_14050,N_13854);
or U15095 (N_15095,N_14199,N_14807);
and U15096 (N_15096,N_10526,N_11408);
nor U15097 (N_15097,N_13313,N_10356);
nor U15098 (N_15098,N_12861,N_14728);
or U15099 (N_15099,N_13995,N_14702);
xor U15100 (N_15100,N_11402,N_12006);
or U15101 (N_15101,N_10422,N_11813);
and U15102 (N_15102,N_14241,N_12519);
nor U15103 (N_15103,N_11502,N_10857);
nand U15104 (N_15104,N_13017,N_14290);
nand U15105 (N_15105,N_14551,N_10812);
xnor U15106 (N_15106,N_10569,N_14271);
and U15107 (N_15107,N_11017,N_13302);
or U15108 (N_15108,N_13166,N_13910);
nand U15109 (N_15109,N_10344,N_13117);
or U15110 (N_15110,N_10679,N_13743);
and U15111 (N_15111,N_11907,N_11752);
or U15112 (N_15112,N_11778,N_10404);
and U15113 (N_15113,N_11391,N_10492);
or U15114 (N_15114,N_11169,N_14623);
nor U15115 (N_15115,N_11625,N_14792);
and U15116 (N_15116,N_12772,N_12847);
nand U15117 (N_15117,N_12060,N_11195);
or U15118 (N_15118,N_14921,N_10719);
nand U15119 (N_15119,N_13792,N_11885);
or U15120 (N_15120,N_12399,N_13823);
and U15121 (N_15121,N_10490,N_11367);
nor U15122 (N_15122,N_11796,N_11198);
or U15123 (N_15123,N_10989,N_13246);
or U15124 (N_15124,N_10225,N_14973);
xnor U15125 (N_15125,N_13038,N_12723);
nand U15126 (N_15126,N_12697,N_12009);
and U15127 (N_15127,N_12218,N_14010);
or U15128 (N_15128,N_14818,N_14868);
or U15129 (N_15129,N_12967,N_14779);
nor U15130 (N_15130,N_13178,N_10608);
or U15131 (N_15131,N_12657,N_11908);
xnor U15132 (N_15132,N_12206,N_14413);
nor U15133 (N_15133,N_10316,N_14924);
and U15134 (N_15134,N_13931,N_12237);
xor U15135 (N_15135,N_10355,N_14597);
xor U15136 (N_15136,N_11872,N_13908);
and U15137 (N_15137,N_10520,N_14022);
nand U15138 (N_15138,N_13026,N_14165);
xor U15139 (N_15139,N_14861,N_13582);
nand U15140 (N_15140,N_14756,N_11955);
nor U15141 (N_15141,N_13205,N_14846);
or U15142 (N_15142,N_14958,N_10242);
nand U15143 (N_15143,N_14114,N_11787);
nor U15144 (N_15144,N_11161,N_14274);
and U15145 (N_15145,N_10597,N_11394);
and U15146 (N_15146,N_13872,N_11542);
nand U15147 (N_15147,N_14488,N_13079);
nand U15148 (N_15148,N_14039,N_11411);
and U15149 (N_15149,N_13547,N_11535);
and U15150 (N_15150,N_13530,N_10525);
xnor U15151 (N_15151,N_13610,N_13467);
or U15152 (N_15152,N_12103,N_12675);
and U15153 (N_15153,N_13780,N_12763);
nand U15154 (N_15154,N_14742,N_11779);
nand U15155 (N_15155,N_10993,N_10434);
nor U15156 (N_15156,N_14099,N_11170);
nor U15157 (N_15157,N_14966,N_10409);
or U15158 (N_15158,N_12358,N_14279);
and U15159 (N_15159,N_12621,N_12761);
and U15160 (N_15160,N_11713,N_10953);
nand U15161 (N_15161,N_13713,N_13364);
and U15162 (N_15162,N_14822,N_12050);
nand U15163 (N_15163,N_12512,N_13053);
xnor U15164 (N_15164,N_12903,N_12068);
nor U15165 (N_15165,N_14492,N_11433);
or U15166 (N_15166,N_12446,N_14733);
nor U15167 (N_15167,N_11951,N_14790);
nand U15168 (N_15168,N_10028,N_14823);
xor U15169 (N_15169,N_12066,N_11550);
or U15170 (N_15170,N_11935,N_13643);
nor U15171 (N_15171,N_11891,N_10038);
nor U15172 (N_15172,N_13732,N_14208);
and U15173 (N_15173,N_10524,N_14242);
xnor U15174 (N_15174,N_10172,N_13640);
nor U15175 (N_15175,N_10996,N_10963);
nor U15176 (N_15176,N_12596,N_13659);
and U15177 (N_15177,N_11911,N_12662);
nand U15178 (N_15178,N_11448,N_13876);
or U15179 (N_15179,N_14520,N_14331);
xnor U15180 (N_15180,N_10137,N_14261);
nor U15181 (N_15181,N_11196,N_10813);
nor U15182 (N_15182,N_12665,N_13575);
nand U15183 (N_15183,N_11293,N_10466);
or U15184 (N_15184,N_10612,N_14554);
nor U15185 (N_15185,N_13857,N_12768);
or U15186 (N_15186,N_13973,N_13075);
xor U15187 (N_15187,N_12632,N_12753);
and U15188 (N_15188,N_11051,N_11346);
and U15189 (N_15189,N_10838,N_11836);
and U15190 (N_15190,N_13744,N_14719);
or U15191 (N_15191,N_14951,N_12958);
nor U15192 (N_15192,N_14535,N_11821);
nor U15193 (N_15193,N_10653,N_10333);
nor U15194 (N_15194,N_12047,N_12441);
and U15195 (N_15195,N_14222,N_11273);
xor U15196 (N_15196,N_14810,N_13923);
nand U15197 (N_15197,N_10619,N_10104);
nand U15198 (N_15198,N_12634,N_10322);
nor U15199 (N_15199,N_13626,N_14156);
and U15200 (N_15200,N_13955,N_10009);
and U15201 (N_15201,N_13325,N_12594);
xnor U15202 (N_15202,N_14078,N_12085);
nor U15203 (N_15203,N_11446,N_11283);
and U15204 (N_15204,N_12230,N_11233);
or U15205 (N_15205,N_10811,N_14243);
nand U15206 (N_15206,N_11518,N_11543);
nor U15207 (N_15207,N_12927,N_12804);
and U15208 (N_15208,N_13937,N_10014);
nand U15209 (N_15209,N_12395,N_11862);
and U15210 (N_15210,N_11879,N_11797);
and U15211 (N_15211,N_14086,N_10227);
nor U15212 (N_15212,N_11066,N_11732);
nand U15213 (N_15213,N_14018,N_11528);
xnor U15214 (N_15214,N_14649,N_12426);
xor U15215 (N_15215,N_10097,N_10907);
xnor U15216 (N_15216,N_11204,N_10588);
and U15217 (N_15217,N_11904,N_12267);
xnor U15218 (N_15218,N_13678,N_11175);
and U15219 (N_15219,N_12158,N_14584);
nor U15220 (N_15220,N_13440,N_10786);
nand U15221 (N_15221,N_10144,N_13232);
xor U15222 (N_15222,N_14531,N_13457);
nor U15223 (N_15223,N_13092,N_12817);
nor U15224 (N_15224,N_11647,N_13508);
nor U15225 (N_15225,N_12531,N_13980);
xor U15226 (N_15226,N_11269,N_13007);
or U15227 (N_15227,N_14066,N_12687);
and U15228 (N_15228,N_10478,N_12171);
and U15229 (N_15229,N_13051,N_11310);
or U15230 (N_15230,N_13870,N_12339);
nand U15231 (N_15231,N_11101,N_13129);
or U15232 (N_15232,N_10665,N_13450);
or U15233 (N_15233,N_10827,N_13550);
xnor U15234 (N_15234,N_14246,N_13903);
or U15235 (N_15235,N_10070,N_10461);
xor U15236 (N_15236,N_14077,N_13239);
nand U15237 (N_15237,N_14490,N_13906);
or U15238 (N_15238,N_10513,N_13182);
nor U15239 (N_15239,N_10185,N_12776);
or U15240 (N_15240,N_10123,N_10850);
xnor U15241 (N_15241,N_13386,N_14440);
nor U15242 (N_15242,N_14294,N_11685);
and U15243 (N_15243,N_11827,N_13921);
xor U15244 (N_15244,N_14647,N_11021);
or U15245 (N_15245,N_14211,N_11574);
nand U15246 (N_15246,N_10934,N_12915);
and U15247 (N_15247,N_11934,N_13829);
and U15248 (N_15248,N_11748,N_13059);
xnor U15249 (N_15249,N_11200,N_14918);
or U15250 (N_15250,N_13174,N_12253);
and U15251 (N_15251,N_11475,N_12294);
nand U15252 (N_15252,N_10842,N_14135);
or U15253 (N_15253,N_14579,N_14328);
nand U15254 (N_15254,N_13396,N_14615);
nor U15255 (N_15255,N_10671,N_13802);
nor U15256 (N_15256,N_10848,N_13796);
nor U15257 (N_15257,N_12767,N_12053);
xor U15258 (N_15258,N_12030,N_10234);
nor U15259 (N_15259,N_11389,N_13617);
and U15260 (N_15260,N_12003,N_12369);
or U15261 (N_15261,N_10237,N_10015);
and U15262 (N_15262,N_11876,N_11084);
and U15263 (N_15263,N_11945,N_14538);
or U15264 (N_15264,N_11994,N_13602);
xnor U15265 (N_15265,N_13573,N_11387);
and U15266 (N_15266,N_11831,N_12386);
nand U15267 (N_15267,N_12014,N_13869);
nor U15268 (N_15268,N_12284,N_11995);
or U15269 (N_15269,N_12376,N_12820);
and U15270 (N_15270,N_14939,N_11039);
nand U15271 (N_15271,N_13400,N_14934);
nand U15272 (N_15272,N_10688,N_12194);
nor U15273 (N_15273,N_14124,N_14275);
nand U15274 (N_15274,N_13131,N_10566);
nand U15275 (N_15275,N_12134,N_12209);
nand U15276 (N_15276,N_12859,N_10919);
nand U15277 (N_15277,N_12522,N_14512);
and U15278 (N_15278,N_10115,N_14590);
and U15279 (N_15279,N_12315,N_11494);
nand U15280 (N_15280,N_11437,N_14363);
xnor U15281 (N_15281,N_11211,N_11948);
and U15282 (N_15282,N_12914,N_13428);
xor U15283 (N_15283,N_14627,N_11899);
or U15284 (N_15284,N_12770,N_10949);
nor U15285 (N_15285,N_11867,N_12409);
nand U15286 (N_15286,N_14332,N_13716);
nor U15287 (N_15287,N_10371,N_11554);
and U15288 (N_15288,N_14968,N_14094);
nor U15289 (N_15289,N_10977,N_10477);
or U15290 (N_15290,N_11260,N_11354);
and U15291 (N_15291,N_14051,N_12102);
nand U15292 (N_15292,N_11179,N_10107);
xnor U15293 (N_15293,N_14672,N_13814);
xor U15294 (N_15294,N_12351,N_14170);
or U15295 (N_15295,N_11024,N_10820);
and U15296 (N_15296,N_12058,N_11497);
and U15297 (N_15297,N_14106,N_14108);
and U15298 (N_15298,N_13500,N_11142);
nor U15299 (N_15299,N_14244,N_14803);
xor U15300 (N_15300,N_13645,N_11505);
nand U15301 (N_15301,N_11108,N_14817);
and U15302 (N_15302,N_12801,N_12159);
nand U15303 (N_15303,N_13693,N_10204);
nor U15304 (N_15304,N_12962,N_13469);
xor U15305 (N_15305,N_10086,N_11672);
xnor U15306 (N_15306,N_13779,N_13430);
or U15307 (N_15307,N_10370,N_11359);
nand U15308 (N_15308,N_10946,N_10906);
xnor U15309 (N_15309,N_11058,N_10924);
nand U15310 (N_15310,N_12556,N_14879);
nand U15311 (N_15311,N_14740,N_12544);
nand U15312 (N_15312,N_13664,N_14012);
or U15313 (N_15313,N_10146,N_11686);
nand U15314 (N_15314,N_13464,N_14898);
nor U15315 (N_15315,N_14626,N_13218);
nor U15316 (N_15316,N_10205,N_10726);
nand U15317 (N_15317,N_11229,N_10681);
nor U15318 (N_15318,N_13614,N_10715);
xnor U15319 (N_15319,N_10802,N_13384);
nand U15320 (N_15320,N_12721,N_13193);
nor U15321 (N_15321,N_10869,N_14635);
nand U15322 (N_15322,N_13072,N_11807);
and U15323 (N_15323,N_14808,N_10375);
nand U15324 (N_15324,N_10241,N_12146);
or U15325 (N_15325,N_14029,N_10625);
nand U15326 (N_15326,N_12895,N_12566);
or U15327 (N_15327,N_10950,N_11660);
nor U15328 (N_15328,N_11256,N_10522);
or U15329 (N_15329,N_13127,N_11463);
or U15330 (N_15330,N_12021,N_13673);
xor U15331 (N_15331,N_10743,N_12345);
nor U15332 (N_15332,N_13326,N_11631);
nand U15333 (N_15333,N_10804,N_12337);
nor U15334 (N_15334,N_14878,N_14226);
and U15335 (N_15335,N_10277,N_14643);
xor U15336 (N_15336,N_10308,N_12031);
and U15337 (N_15337,N_13515,N_13939);
or U15338 (N_15338,N_10990,N_10047);
nand U15339 (N_15339,N_14037,N_14893);
nand U15340 (N_15340,N_12682,N_10892);
nand U15341 (N_15341,N_10354,N_14362);
or U15342 (N_15342,N_11580,N_11268);
or U15343 (N_15343,N_14709,N_11644);
or U15344 (N_15344,N_13266,N_14347);
nand U15345 (N_15345,N_11091,N_14644);
or U15346 (N_15346,N_12563,N_11215);
and U15347 (N_15347,N_14320,N_10660);
xnor U15348 (N_15348,N_13157,N_11567);
or U15349 (N_15349,N_10282,N_10378);
nand U15350 (N_15350,N_11767,N_11308);
nand U15351 (N_15351,N_13137,N_13704);
nand U15352 (N_15352,N_10352,N_13605);
and U15353 (N_15353,N_14085,N_12952);
nor U15354 (N_15354,N_12212,N_10488);
xor U15355 (N_15355,N_11783,N_11014);
and U15356 (N_15356,N_11209,N_11599);
nor U15357 (N_15357,N_13663,N_13418);
nor U15358 (N_15358,N_10512,N_14483);
nor U15359 (N_15359,N_14888,N_14428);
nand U15360 (N_15360,N_11362,N_11057);
or U15361 (N_15361,N_10575,N_12636);
and U15362 (N_15362,N_12991,N_11632);
xor U15363 (N_15363,N_11637,N_10170);
nand U15364 (N_15364,N_11061,N_10785);
and U15365 (N_15365,N_11674,N_13882);
nor U15366 (N_15366,N_12789,N_10002);
and U15367 (N_15367,N_13782,N_13046);
and U15368 (N_15368,N_11399,N_10332);
nor U15369 (N_15369,N_11976,N_13783);
xnor U15370 (N_15370,N_13571,N_14757);
xor U15371 (N_15371,N_13126,N_10223);
nand U15372 (N_15372,N_10814,N_10750);
xnor U15373 (N_15373,N_13098,N_10889);
nand U15374 (N_15374,N_12600,N_11653);
xnor U15375 (N_15375,N_11495,N_10915);
xor U15376 (N_15376,N_11062,N_11249);
xnor U15377 (N_15377,N_12683,N_12762);
nand U15378 (N_15378,N_14234,N_10806);
or U15379 (N_15379,N_10835,N_10433);
or U15380 (N_15380,N_14769,N_12108);
nand U15381 (N_15381,N_10256,N_14035);
and U15382 (N_15382,N_10032,N_11693);
xor U15383 (N_15383,N_12354,N_14120);
or U15384 (N_15384,N_12453,N_13918);
xnor U15385 (N_15385,N_10614,N_11670);
and U15386 (N_15386,N_12281,N_12260);
xor U15387 (N_15387,N_10067,N_11849);
xor U15388 (N_15388,N_12638,N_12299);
nor U15389 (N_15389,N_10531,N_13358);
and U15390 (N_15390,N_12224,N_10418);
xnor U15391 (N_15391,N_13555,N_12878);
and U15392 (N_15392,N_11459,N_13682);
or U15393 (N_15393,N_11522,N_12603);
and U15394 (N_15394,N_11984,N_11913);
nor U15395 (N_15395,N_14256,N_14448);
or U15396 (N_15396,N_11716,N_11578);
nand U15397 (N_15397,N_12593,N_12525);
xnor U15398 (N_15398,N_10279,N_11323);
xor U15399 (N_15399,N_12474,N_11294);
or U15400 (N_15400,N_13034,N_12123);
or U15401 (N_15401,N_10031,N_13551);
xor U15402 (N_15402,N_11028,N_11737);
nor U15403 (N_15403,N_11194,N_10878);
and U15404 (N_15404,N_11230,N_13425);
nor U15405 (N_15405,N_13108,N_11617);
or U15406 (N_15406,N_10446,N_13185);
xor U15407 (N_15407,N_13198,N_12518);
xnor U15408 (N_15408,N_13187,N_13609);
nand U15409 (N_15409,N_13039,N_13214);
xnor U15410 (N_15410,N_14980,N_10468);
nor U15411 (N_15411,N_12523,N_14705);
or U15412 (N_15412,N_13324,N_10039);
nand U15413 (N_15413,N_14444,N_13121);
nand U15414 (N_15414,N_14959,N_14730);
and U15415 (N_15415,N_12320,N_10438);
xnor U15416 (N_15416,N_13770,N_13360);
xnor U15417 (N_15417,N_10935,N_11544);
nand U15418 (N_15418,N_10909,N_12313);
nor U15419 (N_15419,N_14307,N_11639);
and U15420 (N_15420,N_10809,N_11299);
xor U15421 (N_15421,N_12084,N_13216);
xnor U15422 (N_15422,N_12349,N_13806);
and U15423 (N_15423,N_10649,N_10068);
nand U15424 (N_15424,N_14121,N_12027);
nor U15425 (N_15425,N_14062,N_13105);
or U15426 (N_15426,N_11743,N_12661);
xnor U15427 (N_15427,N_10437,N_10323);
xor U15428 (N_15428,N_14585,N_12631);
nand U15429 (N_15429,N_12907,N_13728);
xnor U15430 (N_15430,N_11817,N_14345);
xnor U15431 (N_15431,N_13145,N_13502);
xor U15432 (N_15432,N_14912,N_11010);
nand U15433 (N_15433,N_10300,N_12778);
or U15434 (N_15434,N_13085,N_14940);
and U15435 (N_15435,N_11700,N_13911);
or U15436 (N_15436,N_12165,N_10700);
nand U15437 (N_15437,N_13647,N_11243);
and U15438 (N_15438,N_10948,N_13426);
nand U15439 (N_15439,N_12160,N_13492);
nand U15440 (N_15440,N_14727,N_14801);
and U15441 (N_15441,N_13730,N_11974);
nor U15442 (N_15442,N_13712,N_11106);
nor U15443 (N_15443,N_13777,N_11739);
nand U15444 (N_15444,N_11164,N_13518);
nor U15445 (N_15445,N_13851,N_11485);
nor U15446 (N_15446,N_10886,N_10947);
nand U15447 (N_15447,N_14080,N_11139);
nor U15448 (N_15448,N_13723,N_11180);
or U15449 (N_15449,N_14827,N_11711);
nor U15450 (N_15450,N_12981,N_13454);
nand U15451 (N_15451,N_14296,N_13089);
nand U15452 (N_15452,N_12984,N_14301);
nand U15453 (N_15453,N_13272,N_10233);
nor U15454 (N_15454,N_13195,N_10105);
nor U15455 (N_15455,N_10991,N_12787);
xnor U15456 (N_15456,N_11707,N_14661);
xor U15457 (N_15457,N_14161,N_10696);
and U15458 (N_15458,N_14930,N_13527);
or U15459 (N_15459,N_14550,N_12296);
or U15460 (N_15460,N_10313,N_11889);
xnor U15461 (N_15461,N_13052,N_13970);
nor U15462 (N_15462,N_14498,N_12711);
and U15463 (N_15463,N_12151,N_11113);
nand U15464 (N_15464,N_10291,N_10273);
nand U15465 (N_15465,N_10090,N_10007);
and U15466 (N_15466,N_12608,N_11441);
xor U15467 (N_15467,N_14315,N_10113);
nor U15468 (N_15468,N_11348,N_14507);
and U15469 (N_15469,N_13112,N_13574);
nand U15470 (N_15470,N_12969,N_14183);
xnor U15471 (N_15471,N_13057,N_11745);
or U15472 (N_15472,N_11072,N_10834);
xnor U15473 (N_15473,N_11213,N_11146);
or U15474 (N_15474,N_11172,N_10630);
and U15475 (N_15475,N_13576,N_10944);
xnor U15476 (N_15476,N_10846,N_11094);
nor U15477 (N_15477,N_13686,N_11104);
xor U15478 (N_15478,N_14314,N_10383);
nand U15479 (N_15479,N_13275,N_12479);
or U15480 (N_15480,N_14616,N_10479);
or U15481 (N_15481,N_11070,N_10703);
xnor U15482 (N_15482,N_12994,N_10853);
or U15483 (N_15483,N_12655,N_13894);
and U15484 (N_15484,N_14139,N_14259);
and U15485 (N_15485,N_10782,N_11890);
and U15486 (N_15486,N_14043,N_14101);
or U15487 (N_15487,N_14680,N_10151);
or U15488 (N_15488,N_12759,N_10552);
or U15489 (N_15489,N_11383,N_12249);
or U15490 (N_15490,N_12901,N_10183);
and U15491 (N_15491,N_12642,N_13465);
nor U15492 (N_15492,N_12393,N_11259);
and U15493 (N_15493,N_12814,N_13307);
and U15494 (N_15494,N_10866,N_10917);
nand U15495 (N_15495,N_11270,N_13679);
or U15496 (N_15496,N_13041,N_11052);
nor U15497 (N_15497,N_14799,N_13560);
or U15498 (N_15498,N_14945,N_12756);
or U15499 (N_15499,N_13093,N_14411);
nand U15500 (N_15500,N_14583,N_11532);
nand U15501 (N_15501,N_10845,N_10672);
nor U15502 (N_15502,N_13971,N_10535);
xor U15503 (N_15503,N_13926,N_14175);
or U15504 (N_15504,N_14608,N_11596);
and U15505 (N_15505,N_11563,N_13062);
nor U15506 (N_15506,N_11740,N_12571);
nor U15507 (N_15507,N_11709,N_12127);
nand U15508 (N_15508,N_10611,N_12986);
and U15509 (N_15509,N_12270,N_10243);
nor U15510 (N_15510,N_11873,N_11880);
and U15511 (N_15511,N_12365,N_10843);
nor U15512 (N_15512,N_14813,N_11012);
nand U15513 (N_15513,N_13424,N_12064);
nor U15514 (N_15514,N_10135,N_10983);
or U15515 (N_15515,N_12690,N_12139);
nand U15516 (N_15516,N_12918,N_11598);
nand U15517 (N_15517,N_13957,N_11906);
or U15518 (N_15518,N_12162,N_13567);
nor U15519 (N_15519,N_12420,N_14783);
and U15520 (N_15520,N_11895,N_10473);
and U15521 (N_15521,N_10132,N_14456);
nand U15522 (N_15522,N_14515,N_12564);
or U15523 (N_15523,N_14176,N_14344);
xnor U15524 (N_15524,N_10263,N_12397);
and U15525 (N_15525,N_13173,N_11185);
and U15526 (N_15526,N_14300,N_14092);
nor U15527 (N_15527,N_10261,N_10922);
or U15528 (N_15528,N_10037,N_12589);
or U15529 (N_15529,N_10211,N_11786);
nor U15530 (N_15530,N_12775,N_14047);
nor U15531 (N_15531,N_14151,N_11334);
or U15532 (N_15532,N_11583,N_10624);
nor U15533 (N_15533,N_13714,N_13963);
or U15534 (N_15534,N_11205,N_12025);
nand U15535 (N_15535,N_12602,N_11156);
and U15536 (N_15536,N_11808,N_10913);
xor U15537 (N_15537,N_13701,N_12572);
xnor U15538 (N_15538,N_14254,N_14063);
xor U15539 (N_15539,N_13071,N_14014);
nand U15540 (N_15540,N_11943,N_14860);
and U15541 (N_15541,N_10134,N_14026);
nor U15542 (N_15542,N_10087,N_12063);
nor U15543 (N_15543,N_13634,N_14977);
and U15544 (N_15544,N_14916,N_11620);
or U15545 (N_15545,N_14330,N_11171);
nor U15546 (N_15546,N_10483,N_11450);
nand U15547 (N_15547,N_13201,N_13032);
nor U15548 (N_15548,N_12457,N_13528);
xor U15549 (N_15549,N_10860,N_14381);
or U15550 (N_15550,N_11627,N_10631);
xnor U15551 (N_15551,N_14819,N_12943);
nand U15552 (N_15552,N_11386,N_14423);
nand U15553 (N_15553,N_11398,N_12342);
or U15554 (N_15554,N_14724,N_13738);
xnor U15555 (N_15555,N_10453,N_11536);
and U15556 (N_15556,N_10365,N_10634);
or U15557 (N_15557,N_13022,N_12243);
xor U15558 (N_15558,N_13376,N_11182);
xor U15559 (N_15559,N_14178,N_13858);
and U15560 (N_15560,N_10742,N_12040);
nand U15561 (N_15561,N_14418,N_11667);
or U15562 (N_15562,N_10506,N_13417);
and U15563 (N_15563,N_11593,N_13049);
nand U15564 (N_15564,N_11602,N_14873);
xnor U15565 (N_15565,N_13264,N_10602);
and U15566 (N_15566,N_12248,N_11250);
nand U15567 (N_15567,N_14911,N_14194);
nand U15568 (N_15568,N_11937,N_14858);
xnor U15569 (N_15569,N_14229,N_11393);
nand U15570 (N_15570,N_12163,N_14083);
nand U15571 (N_15571,N_11616,N_13600);
nand U15572 (N_15572,N_12953,N_11140);
nand U15573 (N_15573,N_12802,N_10166);
nand U15574 (N_15574,N_13000,N_10545);
xor U15575 (N_15575,N_12874,N_10560);
nand U15576 (N_15576,N_10231,N_14468);
nor U15577 (N_15577,N_14614,N_14875);
and U15578 (N_15578,N_11344,N_11312);
nand U15579 (N_15579,N_12798,N_13345);
nand U15580 (N_15580,N_10517,N_11311);
or U15581 (N_15581,N_13661,N_10289);
nand U15582 (N_15582,N_10109,N_13964);
nor U15583 (N_15583,N_14794,N_11636);
xnor U15584 (N_15584,N_10080,N_14948);
nor U15585 (N_15585,N_13631,N_14793);
xor U15586 (N_15586,N_13353,N_14563);
xor U15587 (N_15587,N_10708,N_13742);
nand U15588 (N_15588,N_10484,N_11412);
xor U15589 (N_15589,N_12920,N_12852);
xor U15590 (N_15590,N_13884,N_14761);
nor U15591 (N_15591,N_13319,N_10432);
nand U15592 (N_15592,N_14408,N_12039);
nor U15593 (N_15593,N_10317,N_11365);
and U15594 (N_15594,N_14791,N_12092);
nor U15595 (N_15595,N_11130,N_13086);
xor U15596 (N_15596,N_11922,N_14671);
xnor U15597 (N_15597,N_10056,N_12482);
nand U15598 (N_15598,N_13717,N_12332);
nand U15599 (N_15599,N_10540,N_11555);
or U15600 (N_15600,N_11151,N_12835);
and U15601 (N_15601,N_13091,N_12720);
xnor U15602 (N_15602,N_14666,N_10841);
xnor U15603 (N_15603,N_14699,N_14067);
and U15604 (N_15604,N_12262,N_12880);
nand U15605 (N_15605,N_14712,N_12983);
xor U15606 (N_15606,N_13826,N_14502);
and U15607 (N_15607,N_12982,N_10741);
nand U15608 (N_15608,N_10435,N_13483);
nor U15609 (N_15609,N_11238,N_11496);
nor U15610 (N_15610,N_14053,N_11417);
and U15611 (N_15611,N_13204,N_11109);
xnor U15612 (N_15612,N_13950,N_13544);
nand U15613 (N_15613,N_12444,N_10368);
and U15614 (N_15614,N_13297,N_11766);
and U15615 (N_15615,N_11375,N_12390);
or U15616 (N_15616,N_13866,N_14409);
nor U15617 (N_15617,N_13370,N_12938);
xnor U15618 (N_15618,N_10927,N_12656);
nor U15619 (N_15619,N_13317,N_13154);
nand U15620 (N_15620,N_14361,N_12843);
or U15621 (N_15621,N_12364,N_14005);
nand U15622 (N_15622,N_11966,N_13165);
nand U15623 (N_15623,N_11267,N_10783);
xor U15624 (N_15624,N_13481,N_12725);
nor U15625 (N_15625,N_14310,N_11040);
and U15626 (N_15626,N_11347,N_12356);
xnor U15627 (N_15627,N_10412,N_12333);
or U15628 (N_15628,N_12578,N_10362);
nor U15629 (N_15629,N_13294,N_12757);
or U15630 (N_15630,N_12933,N_12330);
nand U15631 (N_15631,N_13657,N_14576);
or U15632 (N_15632,N_13652,N_14581);
nor U15633 (N_15633,N_13238,N_14676);
nand U15634 (N_15634,N_12256,N_14009);
nor U15635 (N_15635,N_13520,N_13504);
nor U15636 (N_15636,N_13538,N_13367);
or U15637 (N_15637,N_10639,N_10456);
and U15638 (N_15638,N_13257,N_14286);
nor U15639 (N_15639,N_14530,N_12863);
nand U15640 (N_15640,N_13128,N_10896);
nor U15641 (N_15641,N_10645,N_11442);
nor U15642 (N_15642,N_14452,N_14768);
and U15643 (N_15643,N_11790,N_10334);
nand U15644 (N_15644,N_14559,N_12537);
and U15645 (N_15645,N_11534,N_10632);
nor U15646 (N_15646,N_10298,N_14484);
xnor U15647 (N_15647,N_14985,N_13410);
and U15648 (N_15648,N_11447,N_13260);
or U15649 (N_15649,N_11990,N_13003);
nor U15650 (N_15650,N_11078,N_12072);
nand U15651 (N_15651,N_12693,N_10425);
and U15652 (N_15652,N_11443,N_10003);
and U15653 (N_15653,N_13978,N_10629);
or U15654 (N_15654,N_13381,N_13074);
xor U15655 (N_15655,N_12704,N_13161);
or U15656 (N_15656,N_12926,N_11946);
and U15657 (N_15657,N_10607,N_14205);
and U15658 (N_15658,N_13996,N_13066);
xnor U15659 (N_15659,N_12238,N_10350);
xnor U15660 (N_15660,N_10385,N_11710);
xor U15661 (N_15661,N_13284,N_13282);
nor U15662 (N_15662,N_12674,N_12079);
xor U15663 (N_15663,N_11638,N_10034);
xor U15664 (N_15664,N_13660,N_11197);
nand U15665 (N_15665,N_12509,N_12780);
nor U15666 (N_15666,N_12875,N_14192);
xor U15667 (N_15667,N_11425,N_11510);
or U15668 (N_15668,N_14759,N_10798);
nor U15669 (N_15669,N_10312,N_14473);
and U15670 (N_15670,N_12401,N_10059);
xnor U15671 (N_15671,N_13027,N_13490);
and U15672 (N_15672,N_12271,N_10442);
or U15673 (N_15673,N_14311,N_13694);
nand U15674 (N_15674,N_12293,N_14459);
and U15675 (N_15675,N_14857,N_13612);
xor U15676 (N_15676,N_10212,N_11227);
nor U15677 (N_15677,N_13152,N_12934);
xor U15678 (N_15678,N_12876,N_12504);
or U15679 (N_15679,N_13194,N_10390);
xnor U15680 (N_15680,N_12404,N_12144);
nor U15681 (N_15681,N_14131,N_11662);
and U15682 (N_15682,N_13229,N_10085);
nand U15683 (N_15683,N_12106,N_12443);
and U15684 (N_15684,N_12119,N_12747);
xor U15685 (N_15685,N_14787,N_10548);
nor U15686 (N_15686,N_13561,N_10250);
nand U15687 (N_15687,N_13569,N_10257);
xnor U15688 (N_15688,N_11665,N_14197);
or U15689 (N_15689,N_12815,N_10236);
nand U15690 (N_15690,N_14737,N_13476);
nand U15691 (N_15691,N_13021,N_11287);
nand U15692 (N_15692,N_13477,N_14582);
nor U15693 (N_15693,N_13925,N_14201);
and U15694 (N_15694,N_12362,N_13443);
nand U15695 (N_15695,N_14654,N_14965);
nor U15696 (N_15696,N_11325,N_13821);
or U15697 (N_15697,N_13503,N_10040);
and U15698 (N_15698,N_14588,N_13151);
nor U15699 (N_15699,N_13975,N_13707);
nor U15700 (N_15700,N_11942,N_14276);
nor U15701 (N_15701,N_13342,N_13290);
nor U15702 (N_15702,N_11055,N_13615);
or U15703 (N_15703,N_13281,N_12381);
xor U15704 (N_15704,N_14885,N_13025);
nor U15705 (N_15705,N_11277,N_14046);
or U15706 (N_15706,N_14527,N_14941);
and U15707 (N_15707,N_13639,N_11297);
xnor U15708 (N_15708,N_10576,N_12301);
and U15709 (N_15709,N_12429,N_13169);
nor U15710 (N_15710,N_11607,N_11460);
nor U15711 (N_15711,N_11993,N_10527);
or U15712 (N_15712,N_11374,N_14074);
nand U15713 (N_15713,N_12825,N_10449);
and U15714 (N_15714,N_12633,N_13365);
nand U15715 (N_15715,N_10692,N_11870);
nand U15716 (N_15716,N_11785,N_13511);
xor U15717 (N_15717,N_11338,N_14831);
or U15718 (N_15718,N_13983,N_10581);
nor U15719 (N_15719,N_11264,N_14734);
nor U15720 (N_15720,N_12508,N_14052);
or U15721 (N_15721,N_14372,N_11390);
or U15722 (N_15722,N_14567,N_11173);
and U15723 (N_15723,N_11924,N_11585);
and U15724 (N_15724,N_11687,N_12118);
nand U15725 (N_15725,N_11789,N_12302);
or U15726 (N_15726,N_11541,N_11473);
or U15727 (N_15727,N_13164,N_10397);
and U15728 (N_15728,N_12115,N_14346);
nor U15729 (N_15729,N_14265,N_12379);
or U15730 (N_15730,N_11328,N_11276);
and U15731 (N_15731,N_11537,N_12442);
and U15732 (N_15732,N_14638,N_11657);
or U15733 (N_15733,N_14667,N_11701);
nor U15734 (N_15734,N_10815,N_13273);
xnor U15735 (N_15735,N_14040,N_13484);
or U15736 (N_15736,N_11640,N_12722);
nor U15737 (N_15737,N_14357,N_13439);
nand U15738 (N_15738,N_14690,N_12517);
nor U15739 (N_15739,N_10102,N_14772);
xor U15740 (N_15740,N_11568,N_13804);
nand U15741 (N_15741,N_12129,N_13380);
and U15742 (N_15742,N_13116,N_13228);
nor U15743 (N_15743,N_10661,N_12254);
or U15744 (N_15744,N_12405,N_12740);
xor U15745 (N_15745,N_12710,N_11444);
xnor U15746 (N_15746,N_13453,N_14150);
and U15747 (N_15747,N_13922,N_14539);
and U15748 (N_15748,N_14038,N_12558);
nor U15749 (N_15749,N_10571,N_14399);
nand U15750 (N_15750,N_11088,N_11438);
nor U15751 (N_15751,N_10388,N_12413);
nor U15752 (N_15752,N_10954,N_11571);
or U15753 (N_15753,N_10379,N_12462);
or U15754 (N_15754,N_11728,N_13058);
nor U15755 (N_15755,N_12785,N_12430);
nand U15756 (N_15756,N_10448,N_10810);
xnor U15757 (N_15757,N_14283,N_14564);
and U15758 (N_15758,N_11038,N_13749);
nor U15759 (N_15759,N_11045,N_12456);
or U15760 (N_15760,N_12142,N_13990);
and U15761 (N_15761,N_10117,N_10532);
and U15762 (N_15762,N_10682,N_12526);
or U15763 (N_15763,N_10894,N_11986);
nand U15764 (N_15764,N_12830,N_11096);
or U15765 (N_15765,N_11549,N_11917);
and U15766 (N_15766,N_11474,N_11335);
xor U15767 (N_15767,N_14436,N_10697);
nor U15768 (N_15768,N_13668,N_10622);
and U15769 (N_15769,N_13488,N_14401);
xor U15770 (N_15770,N_13915,N_13084);
or U15771 (N_15771,N_14317,N_12794);
or U15772 (N_15772,N_12013,N_10680);
xnor U15773 (N_15773,N_10646,N_10060);
or U15774 (N_15774,N_13919,N_10683);
nand U15775 (N_15775,N_13096,N_14747);
xor U15776 (N_15776,N_14669,N_12649);
and U15777 (N_15777,N_14142,N_13343);
nor U15778 (N_15778,N_12325,N_10885);
xor U15779 (N_15779,N_10604,N_10833);
nand U15780 (N_15780,N_13721,N_11231);
and U15781 (N_15781,N_14489,N_10839);
nand U15782 (N_15782,N_12468,N_11970);
xor U15783 (N_15783,N_13844,N_10327);
and U15784 (N_15784,N_11257,N_13012);
nand U15785 (N_15785,N_12035,N_14557);
and U15786 (N_15786,N_12261,N_13125);
xnor U15787 (N_15787,N_12779,N_10746);
nand U15788 (N_15788,N_13192,N_10248);
or U15789 (N_15789,N_14162,N_12061);
nand U15790 (N_15790,N_12929,N_13674);
nor U15791 (N_15791,N_12966,N_13138);
nand U15792 (N_15792,N_12091,N_13883);
nand U15793 (N_15793,N_11341,N_14511);
xnor U15794 (N_15794,N_10124,N_10647);
or U15795 (N_15795,N_12475,N_14519);
and U15796 (N_15796,N_10255,N_13722);
xnor U15797 (N_15797,N_10307,N_14720);
xor U15798 (N_15798,N_14890,N_12378);
or U15799 (N_15799,N_11242,N_13636);
and U15800 (N_15800,N_10942,N_10775);
nand U15801 (N_15801,N_12731,N_12157);
nand U15802 (N_15802,N_10143,N_13466);
nand U15803 (N_15803,N_12105,N_13408);
and U15804 (N_15804,N_12615,N_14805);
nor U15805 (N_15805,N_12684,N_11581);
nor U15806 (N_15806,N_12221,N_10764);
nor U15807 (N_15807,N_10902,N_14508);
or U15808 (N_15808,N_13650,N_10973);
or U15809 (N_15809,N_12306,N_14954);
nor U15810 (N_15810,N_12792,N_14001);
xnor U15811 (N_15811,N_13987,N_11645);
nor U15812 (N_15812,N_13988,N_13951);
and U15813 (N_15813,N_12669,N_14650);
nor U15814 (N_15814,N_10069,N_14698);
nand U15815 (N_15815,N_12304,N_14111);
nor U15816 (N_15816,N_11768,N_13373);
nand U15817 (N_15817,N_11162,N_11999);
and U15818 (N_15818,N_10208,N_11396);
nor U15819 (N_15819,N_12219,N_10995);
nand U15820 (N_15820,N_11461,N_12207);
or U15821 (N_15821,N_12891,N_10347);
or U15822 (N_15822,N_12235,N_14877);
nand U15823 (N_15823,N_10416,N_12829);
and U15824 (N_15824,N_12045,N_11265);
and U15825 (N_15825,N_13653,N_14091);
nor U15826 (N_15826,N_12856,N_14560);
or U15827 (N_15827,N_10911,N_12463);
nor U15828 (N_15828,N_12997,N_12972);
xor U15829 (N_15829,N_14611,N_14068);
and U15830 (N_15830,N_13522,N_13377);
nand U15831 (N_15831,N_14853,N_10555);
or U15832 (N_15832,N_14738,N_13321);
nand U15833 (N_15833,N_12609,N_12643);
nand U15834 (N_15834,N_11314,N_12467);
or U15835 (N_15835,N_11646,N_10213);
xnor U15836 (N_15836,N_14425,N_13581);
nor U15837 (N_15837,N_12070,N_12244);
or U15838 (N_15838,N_10755,N_10216);
nand U15839 (N_15839,N_11718,N_13186);
nand U15840 (N_15840,N_11750,N_13620);
and U15841 (N_15841,N_12275,N_10314);
nand U15842 (N_15842,N_10956,N_12884);
xnor U15843 (N_15843,N_14849,N_11041);
xnor U15844 (N_15844,N_12911,N_11824);
or U15845 (N_15845,N_10793,N_12745);
xnor U15846 (N_15846,N_14485,N_13947);
and U15847 (N_15847,N_12750,N_13836);
and U15848 (N_15848,N_10536,N_13753);
and U15849 (N_15849,N_13235,N_14662);
nand U15850 (N_15850,N_14814,N_10043);
or U15851 (N_15851,N_14174,N_13961);
nor U15852 (N_15852,N_10339,N_11501);
or U15853 (N_15853,N_14798,N_11649);
xor U15854 (N_15854,N_14477,N_12231);
and U15855 (N_15855,N_10148,N_11973);
or U15856 (N_15856,N_14367,N_13532);
nor U15857 (N_15857,N_14044,N_14700);
and U15858 (N_15858,N_14933,N_11121);
nand U15859 (N_15859,N_12671,N_13967);
or U15860 (N_15860,N_10041,N_13399);
nor U15861 (N_15861,N_10796,N_12581);
xnor U15862 (N_15862,N_11527,N_12488);
or U15863 (N_15863,N_13215,N_14618);
and U15864 (N_15864,N_12751,N_12434);
or U15865 (N_15865,N_10518,N_14209);
nand U15866 (N_15866,N_13748,N_11663);
xnor U15867 (N_15867,N_12871,N_10229);
xnor U15868 (N_15868,N_14910,N_10001);
or U15869 (N_15869,N_13740,N_11628);
nor U15870 (N_15870,N_13040,N_13189);
nand U15871 (N_15871,N_11791,N_11049);
nor U15872 (N_15872,N_14393,N_10182);
xnor U15873 (N_15873,N_12297,N_10452);
or U15874 (N_15874,N_13822,N_13874);
xor U15875 (N_15875,N_14703,N_11792);
and U15876 (N_15876,N_12738,N_14932);
xnor U15877 (N_15877,N_11606,N_13395);
or U15878 (N_15878,N_10064,N_12384);
xor U15879 (N_15879,N_10405,N_12819);
nand U15880 (N_15880,N_11306,N_14926);
nor U15881 (N_15881,N_12694,N_12312);
nor U15882 (N_15882,N_13593,N_11559);
or U15883 (N_15883,N_13506,N_11184);
and U15884 (N_15884,N_13363,N_11129);
nand U15885 (N_15885,N_10266,N_10297);
nor U15886 (N_15886,N_12732,N_11025);
or U15887 (N_15887,N_12950,N_11351);
or U15888 (N_15888,N_13684,N_10200);
and U15889 (N_15889,N_10974,N_14715);
nor U15890 (N_15890,N_10559,N_13197);
nand U15891 (N_15891,N_11439,N_12605);
xor U15892 (N_15892,N_10530,N_12389);
nor U15893 (N_15893,N_12473,N_14392);
nor U15894 (N_15894,N_10901,N_14118);
nand U15895 (N_15895,N_14633,N_11959);
or U15896 (N_15896,N_10738,N_14809);
nor U15897 (N_15897,N_12528,N_13242);
and U15898 (N_15898,N_13767,N_12580);
nand U15899 (N_15899,N_10711,N_14223);
or U15900 (N_15900,N_12700,N_13879);
and U15901 (N_15901,N_14258,N_14528);
nor U15902 (N_15902,N_10240,N_12109);
nor U15903 (N_15903,N_11635,N_12140);
xnor U15904 (N_15904,N_13762,N_11586);
and U15905 (N_15905,N_12278,N_13579);
nand U15906 (N_15906,N_11315,N_10824);
nand U15907 (N_15907,N_10510,N_11037);
and U15908 (N_15908,N_11893,N_11694);
nand U15909 (N_15909,N_13316,N_13795);
nand U15910 (N_15910,N_13033,N_13943);
nand U15911 (N_15911,N_11029,N_12276);
xor U15912 (N_15912,N_11643,N_13029);
nor U15913 (N_15913,N_12904,N_14735);
and U15914 (N_15914,N_10230,N_11920);
xnor U15915 (N_15915,N_12536,N_12503);
nand U15916 (N_15916,N_13607,N_11634);
or U15917 (N_15917,N_11176,N_14177);
or U15918 (N_15918,N_13509,N_14758);
or U15919 (N_15919,N_14049,N_14978);
nor U15920 (N_15920,N_10072,N_14388);
and U15921 (N_15921,N_13226,N_14424);
or U15922 (N_15922,N_14543,N_13143);
nor U15923 (N_15923,N_13885,N_13054);
xor U15924 (N_15924,N_11526,N_11671);
or U15925 (N_15925,N_14847,N_10736);
and U15926 (N_15926,N_10740,N_13761);
nand U15927 (N_15927,N_12425,N_14675);
xnor U15928 (N_15928,N_14632,N_13314);
and U15929 (N_15929,N_12513,N_13283);
and U15930 (N_15930,N_10689,N_10819);
nand U15931 (N_15931,N_14562,N_13747);
nor U15932 (N_15932,N_14069,N_11856);
nand U15933 (N_15933,N_13006,N_14693);
xor U15934 (N_15934,N_12818,N_14826);
nor U15935 (N_15935,N_13525,N_13447);
xor U15936 (N_15936,N_10693,N_13590);
nand U15937 (N_15937,N_10463,N_14386);
or U15938 (N_15938,N_13383,N_14682);
nor U15939 (N_15939,N_13766,N_14655);
or U15940 (N_15940,N_14864,N_13240);
nand U15941 (N_15941,N_14545,N_13306);
and U15942 (N_15942,N_14285,N_13162);
and U15943 (N_15943,N_13513,N_11777);
xnor U15944 (N_15944,N_11720,N_14800);
and U15945 (N_15945,N_12452,N_10423);
or U15946 (N_15946,N_13351,N_12834);
nand U15947 (N_15947,N_11688,N_14711);
and U15948 (N_15948,N_13907,N_14619);
nor U15949 (N_15949,N_12412,N_14899);
or U15950 (N_15950,N_12141,N_11730);
nand U15951 (N_15951,N_14645,N_12511);
nand U15952 (N_15952,N_10724,N_13920);
xnor U15953 (N_15953,N_10932,N_14922);
xnor U15954 (N_15954,N_14887,N_12619);
or U15955 (N_15955,N_10210,N_12624);
or U15956 (N_15956,N_11882,N_10863);
nand U15957 (N_15957,N_13394,N_10986);
and U15958 (N_15958,N_10926,N_11421);
or U15959 (N_15959,N_12188,N_14555);
xnor U15960 (N_15960,N_11244,N_10471);
nand U15961 (N_15961,N_11759,N_14677);
nand U15962 (N_15962,N_12319,N_11449);
nor U15963 (N_15963,N_12112,N_13683);
nor U15964 (N_15964,N_13862,N_11814);
xor U15965 (N_15965,N_11888,N_13419);
nand U15966 (N_15966,N_10357,N_13989);
xor U15967 (N_15967,N_10128,N_11572);
nand U15968 (N_15968,N_14821,N_13946);
xnor U15969 (N_15969,N_11794,N_12960);
and U15970 (N_15970,N_12599,N_13685);
nor U15971 (N_15971,N_14663,N_11749);
or U15972 (N_15972,N_13778,N_13553);
and U15973 (N_15973,N_14353,N_10284);
xor U15974 (N_15974,N_14224,N_10816);
xnor U15975 (N_15975,N_14387,N_12601);
or U15976 (N_15976,N_14321,N_10467);
or U15977 (N_15977,N_14042,N_11582);
xor U15978 (N_15978,N_11538,N_12200);
or U15979 (N_15979,N_14907,N_11358);
nor U15980 (N_15980,N_13962,N_12514);
nand U15981 (N_15981,N_12083,N_14514);
nand U15982 (N_15982,N_14696,N_12749);
or U15983 (N_15983,N_11962,N_14105);
and U15984 (N_15984,N_10852,N_12323);
and U15985 (N_15985,N_12240,N_10095);
or U15986 (N_15986,N_13142,N_10421);
or U15987 (N_15987,N_13315,N_14305);
nor U15988 (N_15988,N_13270,N_13592);
xor U15989 (N_15989,N_11714,N_10500);
and U15990 (N_15990,N_12993,N_14030);
and U15991 (N_15991,N_10595,N_13736);
xor U15992 (N_15992,N_10324,N_11486);
nor U15993 (N_15993,N_10396,N_14904);
and U15994 (N_15994,N_10675,N_14881);
xor U15995 (N_15995,N_13496,N_10089);
or U15996 (N_15996,N_13403,N_11220);
xnor U15997 (N_15997,N_12951,N_11914);
nand U15998 (N_15998,N_13878,N_11507);
nand U15999 (N_15999,N_13741,N_10340);
nand U16000 (N_16000,N_11552,N_13611);
nand U16001 (N_16001,N_12587,N_13065);
and U16002 (N_16002,N_12677,N_12411);
nand U16003 (N_16003,N_11818,N_13433);
xor U16004 (N_16004,N_12046,N_13563);
nor U16005 (N_16005,N_10780,N_13793);
nand U16006 (N_16006,N_10861,N_14741);
nand U16007 (N_16007,N_13088,N_14636);
and U16008 (N_16008,N_11721,N_13048);
and U16009 (N_16009,N_11622,N_13109);
xnor U16010 (N_16010,N_12550,N_14048);
nand U16011 (N_16011,N_11487,N_12202);
nor U16012 (N_16012,N_11329,N_10206);
nor U16013 (N_16013,N_13299,N_13241);
nor U16014 (N_16014,N_10881,N_13848);
xor U16015 (N_16015,N_14964,N_11304);
nor U16016 (N_16016,N_12082,N_13799);
or U16017 (N_16017,N_14404,N_10019);
and U16018 (N_16018,N_11690,N_10061);
and U16019 (N_16019,N_13638,N_12073);
nor U16020 (N_16020,N_14358,N_11059);
and U16021 (N_16021,N_10893,N_11679);
xnor U16022 (N_16022,N_10348,N_10870);
or U16023 (N_16023,N_11423,N_10615);
nor U16024 (N_16024,N_12607,N_10648);
or U16025 (N_16025,N_13094,N_14497);
xor U16026 (N_16026,N_11083,N_10010);
and U16027 (N_16027,N_14288,N_14829);
nand U16028 (N_16028,N_11208,N_12868);
xnor U16029 (N_16029,N_11776,N_11434);
or U16030 (N_16030,N_11704,N_12673);
xor U16031 (N_16031,N_11798,N_11819);
xnor U16032 (N_16032,N_13107,N_12712);
nand U16033 (N_16033,N_13234,N_14574);
and U16034 (N_16034,N_12357,N_12236);
or U16035 (N_16035,N_14495,N_11573);
xnor U16036 (N_16036,N_13005,N_13830);
or U16037 (N_16037,N_13422,N_10757);
nand U16038 (N_16038,N_14573,N_12569);
xnor U16039 (N_16039,N_14471,N_10712);
and U16040 (N_16040,N_13018,N_11503);
nand U16041 (N_16041,N_14837,N_11868);
nand U16042 (N_16042,N_14494,N_13549);
nand U16043 (N_16043,N_10856,N_10358);
nor U16044 (N_16044,N_11981,N_13475);
or U16045 (N_16045,N_10864,N_11212);
and U16046 (N_16046,N_11609,N_12480);
and U16047 (N_16047,N_11432,N_13427);
nand U16048 (N_16048,N_11327,N_14664);
and U16049 (N_16049,N_10694,N_11138);
nor U16050 (N_16050,N_10657,N_14334);
nor U16051 (N_16051,N_10543,N_14057);
xor U16052 (N_16052,N_11127,N_13147);
or U16053 (N_16053,N_11682,N_13348);
or U16054 (N_16054,N_12809,N_13635);
xor U16055 (N_16055,N_11302,N_12579);
xor U16056 (N_16056,N_14461,N_14110);
nor U16057 (N_16057,N_10539,N_10221);
or U16058 (N_16058,N_12945,N_12407);
nand U16059 (N_16059,N_13649,N_12786);
and U16060 (N_16060,N_12257,N_14132);
and U16061 (N_16061,N_13482,N_14834);
xor U16062 (N_16062,N_14141,N_12626);
or U16063 (N_16063,N_14991,N_13060);
nand U16064 (N_16064,N_10879,N_13261);
or U16065 (N_16065,N_13303,N_13362);
nor U16066 (N_16066,N_10101,N_14937);
nand U16067 (N_16067,N_12752,N_11958);
nor U16068 (N_16068,N_10495,N_10568);
or U16069 (N_16069,N_12081,N_12890);
nand U16070 (N_16070,N_14023,N_14402);
and U16071 (N_16071,N_12341,N_10082);
nand U16072 (N_16072,N_13227,N_11060);
or U16073 (N_16073,N_13945,N_10193);
nor U16074 (N_16074,N_10523,N_13665);
xor U16075 (N_16075,N_11562,N_10320);
or U16076 (N_16076,N_12765,N_12707);
or U16077 (N_16077,N_12182,N_13865);
nand U16078 (N_16078,N_14716,N_14438);
and U16079 (N_16079,N_13670,N_14430);
xor U16080 (N_16080,N_13914,N_11144);
and U16081 (N_16081,N_14123,N_10868);
and U16082 (N_16082,N_13120,N_13016);
nor U16083 (N_16083,N_12346,N_13347);
and U16084 (N_16084,N_10669,N_10055);
and U16085 (N_16085,N_13859,N_14364);
or U16086 (N_16086,N_14784,N_13263);
or U16087 (N_16087,N_10778,N_10713);
or U16088 (N_16088,N_12855,N_13566);
or U16089 (N_16089,N_14979,N_13545);
nand U16090 (N_16090,N_11132,N_12595);
nand U16091 (N_16091,N_10195,N_11377);
nand U16092 (N_16092,N_10136,N_10659);
xnor U16093 (N_16093,N_13666,N_10295);
or U16094 (N_16094,N_14373,N_10603);
xnor U16095 (N_16095,N_14277,N_10033);
or U16096 (N_16096,N_14056,N_12255);
nand U16097 (N_16097,N_14348,N_11470);
nor U16098 (N_16098,N_14460,N_14065);
nor U16099 (N_16099,N_11678,N_14739);
xor U16100 (N_16100,N_10556,N_12155);
xnor U16101 (N_16101,N_10194,N_11850);
nor U16102 (N_16102,N_14339,N_12741);
xor U16103 (N_16103,N_14475,N_12999);
xnor U16104 (N_16104,N_10781,N_13429);
and U16105 (N_16105,N_13423,N_11073);
nand U16106 (N_16106,N_13539,N_11727);
and U16107 (N_16107,N_12561,N_12098);
nand U16108 (N_16108,N_13258,N_12625);
xnor U16109 (N_16109,N_10278,N_14917);
nor U16110 (N_16110,N_13587,N_13231);
xnor U16111 (N_16111,N_13023,N_11491);
or U16112 (N_16112,N_12265,N_13768);
nand U16113 (N_16113,N_11284,N_14854);
nor U16114 (N_16114,N_14743,N_14687);
and U16115 (N_16115,N_10005,N_13774);
xnor U16116 (N_16116,N_12392,N_10218);
and U16117 (N_16117,N_11608,N_14565);
nand U16118 (N_16118,N_14601,N_13835);
or U16119 (N_16119,N_10222,N_12527);
or U16120 (N_16120,N_10426,N_11940);
nand U16121 (N_16121,N_13681,N_10826);
and U16122 (N_16122,N_14500,N_11004);
nor U16123 (N_16123,N_11805,N_10960);
nor U16124 (N_16124,N_12164,N_10419);
or U16125 (N_16125,N_12652,N_11166);
xnor U16126 (N_16126,N_14232,N_14996);
nand U16127 (N_16127,N_13389,N_14060);
nand U16128 (N_16128,N_11366,N_13269);
and U16129 (N_16129,N_11481,N_14185);
nand U16130 (N_16130,N_13222,N_11406);
nand U16131 (N_16131,N_14045,N_12663);
xnor U16132 (N_16132,N_12344,N_13042);
nand U16133 (N_16133,N_11771,N_10551);
xor U16134 (N_16134,N_13013,N_14433);
xnor U16135 (N_16135,N_14678,N_11969);
nor U16136 (N_16136,N_13839,N_13411);
xor U16137 (N_16137,N_13431,N_12754);
nor U16138 (N_16138,N_11630,N_10858);
xnor U16139 (N_16139,N_11553,N_10720);
xor U16140 (N_16140,N_12172,N_13864);
xnor U16141 (N_16141,N_12485,N_10401);
xnor U16142 (N_16142,N_12881,N_13909);
nand U16143 (N_16143,N_10965,N_14729);
xor U16144 (N_16144,N_10709,N_14231);
or U16145 (N_16145,N_12777,N_11949);
or U16146 (N_16146,N_13966,N_14482);
nand U16147 (N_16147,N_10801,N_13180);
and U16148 (N_16148,N_10972,N_11430);
nor U16149 (N_16149,N_14651,N_11504);
nand U16150 (N_16150,N_12870,N_11471);
xnor U16151 (N_16151,N_13134,N_12490);
nand U16152 (N_16152,N_13210,N_12806);
nand U16153 (N_16153,N_11246,N_11651);
nand U16154 (N_16154,N_13754,N_11854);
or U16155 (N_16155,N_12858,N_12795);
nand U16156 (N_16156,N_10925,N_12264);
or U16157 (N_16157,N_14400,N_11464);
or U16158 (N_16158,N_14215,N_14518);
nand U16159 (N_16159,N_14405,N_11466);
and U16160 (N_16160,N_14993,N_11985);
and U16161 (N_16161,N_12813,N_12388);
and U16162 (N_16162,N_10088,N_10905);
nor U16163 (N_16163,N_13847,N_14872);
xnor U16164 (N_16164,N_13499,N_14147);
or U16165 (N_16165,N_12782,N_14499);
xor U16166 (N_16166,N_13267,N_11355);
or U16167 (N_16167,N_14340,N_12438);
nor U16168 (N_16168,N_13346,N_10876);
nor U16169 (N_16169,N_14845,N_13371);
and U16170 (N_16170,N_13637,N_11237);
nor U16171 (N_16171,N_10302,N_10976);
nand U16172 (N_16172,N_14990,N_11291);
nand U16173 (N_16173,N_14031,N_10169);
nand U16174 (N_16174,N_14710,N_11415);
or U16175 (N_16175,N_12568,N_12622);
or U16176 (N_16176,N_10577,N_11005);
or U16177 (N_16177,N_13497,N_10025);
or U16178 (N_16178,N_11677,N_11489);
xor U16179 (N_16179,N_14975,N_11765);
xor U16180 (N_16180,N_10058,N_14504);
and U16181 (N_16181,N_13068,N_14280);
and U16182 (N_16182,N_12258,N_13070);
or U16183 (N_16183,N_10338,N_11624);
nand U16184 (N_16184,N_11188,N_11054);
and U16185 (N_16185,N_10967,N_14778);
or U16186 (N_16186,N_11980,N_12310);
nor U16187 (N_16187,N_13752,N_14414);
nor U16188 (N_16188,N_11153,N_11705);
xor U16189 (N_16189,N_14396,N_14656);
xnor U16190 (N_16190,N_14824,N_13568);
nor U16191 (N_16191,N_11296,N_14920);
nand U16192 (N_16192,N_10580,N_13616);
and U16193 (N_16193,N_11659,N_12078);
or U16194 (N_16194,N_14841,N_12549);
and U16195 (N_16195,N_13808,N_14082);
xor U16196 (N_16196,N_14694,N_14812);
nand U16197 (N_16197,N_11251,N_10553);
and U16198 (N_16198,N_13135,N_10275);
nor U16199 (N_16199,N_13809,N_10751);
and U16200 (N_16200,N_13415,N_14081);
nand U16201 (N_16201,N_13318,N_11364);
xnor U16202 (N_16202,N_13486,N_10096);
nand U16203 (N_16203,N_13604,N_10966);
nor U16204 (N_16204,N_13993,N_13595);
or U16205 (N_16205,N_12470,N_13441);
or U16206 (N_16206,N_14981,N_14534);
and U16207 (N_16207,N_14642,N_14248);
xnor U16208 (N_16208,N_14383,N_11963);
and U16209 (N_16209,N_10147,N_10420);
and U16210 (N_16210,N_12447,N_13554);
xor U16211 (N_16211,N_14251,N_14587);
nor U16212 (N_16212,N_11281,N_12042);
xnor U16213 (N_16213,N_10904,N_11566);
or U16214 (N_16214,N_12575,N_11370);
or U16215 (N_16215,N_10714,N_12427);
xor U16216 (N_16216,N_13729,N_13507);
xor U16217 (N_16217,N_12002,N_10328);
nor U16218 (N_16218,N_14905,N_10847);
and U16219 (N_16219,N_10093,N_10249);
nor U16220 (N_16220,N_13200,N_11143);
nand U16221 (N_16221,N_13245,N_14610);
or U16222 (N_16222,N_13557,N_11240);
or U16223 (N_16223,N_11128,N_12591);
and U16224 (N_16224,N_12996,N_11453);
xnor U16225 (N_16225,N_11499,N_12702);
xnor U16226 (N_16226,N_12340,N_13406);
or U16227 (N_16227,N_13259,N_13435);
and U16228 (N_16228,N_11515,N_14752);
and U16229 (N_16229,N_12385,N_10578);
and U16230 (N_16230,N_13292,N_10601);
and U16231 (N_16231,N_12574,N_14173);
and U16232 (N_16232,N_12680,N_10285);
nand U16233 (N_16233,N_14714,N_13271);
xnor U16234 (N_16234,N_11925,N_10733);
nand U16235 (N_16235,N_11254,N_12897);
nand U16236 (N_16236,N_11989,N_12627);
and U16237 (N_16237,N_11684,N_10541);
nor U16238 (N_16238,N_10519,N_11222);
nor U16239 (N_16239,N_13463,N_12418);
or U16240 (N_16240,N_14206,N_12548);
nand U16241 (N_16241,N_11729,N_14166);
or U16242 (N_16242,N_14028,N_12487);
xnor U16243 (N_16243,N_10664,N_12363);
or U16244 (N_16244,N_10260,N_12057);
xor U16245 (N_16245,N_12493,N_12748);
xor U16246 (N_16246,N_10855,N_11380);
nor U16247 (N_16247,N_14575,N_11285);
or U16248 (N_16248,N_13662,N_14323);
nand U16249 (N_16249,N_11189,N_10769);
nor U16250 (N_16250,N_12318,N_12826);
or U16251 (N_16251,N_12259,N_13168);
nand U16252 (N_16252,N_12706,N_12954);
and U16253 (N_16253,N_10690,N_10883);
xnor U16254 (N_16254,N_11478,N_10299);
or U16255 (N_16255,N_11699,N_11451);
nand U16256 (N_16256,N_14375,N_12744);
and U16257 (N_16257,N_13253,N_14453);
xor U16258 (N_16258,N_11742,N_12848);
or U16259 (N_16259,N_10791,N_11508);
or U16260 (N_16260,N_14128,N_12460);
nor U16261 (N_16261,N_10618,N_11397);
xor U16262 (N_16262,N_11462,N_12583);
nand U16263 (N_16263,N_13414,N_11523);
nand U16264 (N_16264,N_11455,N_11784);
xnor U16265 (N_16265,N_13584,N_12737);
xor U16266 (N_16266,N_14944,N_11236);
nand U16267 (N_16267,N_12854,N_14773);
xor U16268 (N_16268,N_11067,N_12554);
or U16269 (N_16269,N_11271,N_11519);
xnor U16270 (N_16270,N_12507,N_11764);
and U16271 (N_16271,N_13873,N_13455);
and U16272 (N_16272,N_12869,N_13929);
or U16273 (N_16273,N_14263,N_11741);
or U16274 (N_16274,N_10224,N_12011);
xnor U16275 (N_16275,N_12557,N_14352);
and U16276 (N_16276,N_14949,N_10329);
xnor U16277 (N_16277,N_11427,N_10402);
and U16278 (N_16278,N_14416,N_10219);
or U16279 (N_16279,N_10979,N_11431);
nor U16280 (N_16280,N_12001,N_13892);
nor U16281 (N_16281,N_14568,N_11506);
nand U16282 (N_16282,N_14148,N_14443);
nand U16283 (N_16283,N_13082,N_10048);
nor U16284 (N_16284,N_10596,N_12505);
nand U16285 (N_16285,N_12867,N_11360);
and U16286 (N_16286,N_14159,N_10381);
and U16287 (N_16287,N_14763,N_10044);
or U16288 (N_16288,N_11134,N_12010);
nor U16289 (N_16289,N_13798,N_10267);
xor U16290 (N_16290,N_13438,N_10605);
and U16291 (N_16291,N_13256,N_11343);
and U16292 (N_16292,N_10156,N_13898);
nand U16293 (N_16293,N_10728,N_10120);
xnor U16294 (N_16294,N_12893,N_12524);
and U16295 (N_16295,N_10589,N_10191);
nand U16296 (N_16296,N_11855,N_13737);
or U16297 (N_16297,N_12597,N_14697);
or U16298 (N_16298,N_10112,N_12562);
nor U16299 (N_16299,N_10023,N_13789);
or U16300 (N_16300,N_14365,N_13608);
xnor U16301 (N_16301,N_12213,N_12629);
nor U16302 (N_16302,N_11102,N_10941);
and U16303 (N_16303,N_10181,N_13123);
or U16304 (N_16304,N_12150,N_14270);
and U16305 (N_16305,N_13680,N_14797);
nor U16306 (N_16306,N_14624,N_12167);
and U16307 (N_16307,N_12336,N_12251);
nand U16308 (N_16308,N_11158,N_12906);
nand U16309 (N_16309,N_12555,N_14117);
xor U16310 (N_16310,N_14419,N_13936);
or U16311 (N_16311,N_12350,N_14838);
nor U16312 (N_16312,N_13881,N_13148);
and U16313 (N_16313,N_10464,N_13958);
or U16314 (N_16314,N_13230,N_12128);
xor U16315 (N_16315,N_13090,N_11498);
nand U16316 (N_16316,N_13999,N_13887);
nand U16317 (N_16317,N_13113,N_11857);
nand U16318 (N_16318,N_13177,N_12483);
nor U16319 (N_16319,N_13011,N_14153);
xnor U16320 (N_16320,N_12215,N_11658);
and U16321 (N_16321,N_10198,N_11086);
nor U16322 (N_16322,N_13491,N_14592);
and U16323 (N_16323,N_10465,N_14093);
nor U16324 (N_16324,N_13160,N_14354);
nor U16325 (N_16325,N_10598,N_12181);
and U16326 (N_16326,N_14657,N_11248);
and U16327 (N_16327,N_12831,N_11859);
and U16328 (N_16328,N_11114,N_10767);
xnor U16329 (N_16329,N_11400,N_12170);
or U16330 (N_16330,N_12743,N_11087);
nor U16331 (N_16331,N_11384,N_10737);
nand U16332 (N_16332,N_10424,N_14537);
xor U16333 (N_16333,N_14225,N_11843);
and U16334 (N_16334,N_13473,N_10756);
nand U16335 (N_16335,N_10662,N_13019);
xnor U16336 (N_16336,N_11352,N_14992);
xnor U16337 (N_16337,N_10969,N_14011);
and U16338 (N_16338,N_11300,N_12466);
nand U16339 (N_16339,N_11992,N_12449);
nand U16340 (N_16340,N_11339,N_12935);
xnor U16341 (N_16341,N_11641,N_13498);
or U16342 (N_16342,N_10971,N_14866);
nand U16343 (N_16343,N_12087,N_12790);
and U16344 (N_16344,N_12004,N_13891);
nand U16345 (N_16345,N_13361,N_12298);
nand U16346 (N_16346,N_12845,N_11372);
xnor U16347 (N_16347,N_10066,N_12069);
or U16348 (N_16348,N_12149,N_11968);
nor U16349 (N_16349,N_11960,N_13119);
or U16350 (N_16350,N_11147,N_13448);
nor U16351 (N_16351,N_10480,N_12189);
nor U16352 (N_16352,N_13700,N_14541);
nor U16353 (N_16353,N_13114,N_12905);
and U16354 (N_16354,N_11932,N_14235);
and U16355 (N_16355,N_13558,N_13122);
xnor U16356 (N_16356,N_14929,N_11829);
nand U16357 (N_16357,N_14673,N_13401);
xnor U16358 (N_16358,N_10214,N_11774);
and U16359 (N_16359,N_10616,N_12928);
nand U16360 (N_16360,N_11116,N_10447);
xnor U16361 (N_16361,N_10702,N_14599);
or U16362 (N_16362,N_10800,N_10945);
and U16363 (N_16363,N_12924,N_12501);
nor U16364 (N_16364,N_12210,N_12423);
nand U16365 (N_16365,N_10762,N_11695);
or U16366 (N_16366,N_10024,N_10013);
nor U16367 (N_16367,N_12807,N_11181);
or U16368 (N_16368,N_10859,N_13630);
xnor U16369 (N_16369,N_11775,N_14869);
or U16370 (N_16370,N_10862,N_11997);
or U16371 (N_16371,N_13432,N_12923);
xor U16372 (N_16372,N_13268,N_12664);
nor U16373 (N_16373,N_13434,N_12439);
nand U16374 (N_16374,N_13710,N_10196);
xnor U16375 (N_16375,N_13327,N_12862);
nor U16376 (N_16376,N_12547,N_11961);
nand U16377 (N_16377,N_11708,N_14437);
nor U16378 (N_16378,N_11007,N_11077);
nand U16379 (N_16379,N_10158,N_11452);
nor U16380 (N_16380,N_13543,N_12849);
and U16381 (N_16381,N_13050,N_10875);
xnor U16382 (N_16382,N_12059,N_11221);
xor U16383 (N_16383,N_13405,N_14679);
nor U16384 (N_16384,N_13896,N_13301);
or U16385 (N_16385,N_13899,N_14016);
xor U16386 (N_16386,N_13044,N_11145);
xor U16387 (N_16387,N_10542,N_12691);
and U16388 (N_16388,N_13901,N_11610);
nand U16389 (N_16389,N_14842,N_12247);
nand U16390 (N_16390,N_11050,N_14297);
or U16391 (N_16391,N_12729,N_10652);
nand U16392 (N_16392,N_13875,N_13472);
nor U16393 (N_16393,N_13378,N_10360);
and U16394 (N_16394,N_10765,N_11201);
nand U16395 (N_16395,N_12478,N_10021);
nor U16396 (N_16396,N_11735,N_12530);
nand U16397 (N_16397,N_13601,N_13095);
xor U16398 (N_16398,N_13596,N_12560);
nand U16399 (N_16399,N_10244,N_10797);
nor U16400 (N_16400,N_10270,N_12432);
and U16401 (N_16401,N_13167,N_12500);
or U16402 (N_16402,N_11719,N_10472);
nand U16403 (N_16403,N_11289,N_11722);
nand U16404 (N_16404,N_14828,N_13344);
nand U16405 (N_16405,N_11834,N_12486);
or U16406 (N_16406,N_11884,N_14871);
and U16407 (N_16407,N_14517,N_12335);
nor U16408 (N_16408,N_11938,N_10103);
xnor U16409 (N_16409,N_10880,N_13860);
nor U16410 (N_16410,N_10415,N_11324);
or U16411 (N_16411,N_12948,N_10174);
xor U16412 (N_16412,N_10768,N_10636);
and U16413 (N_16413,N_11875,N_12539);
nand U16414 (N_16414,N_12094,N_13183);
or U16415 (N_16415,N_10035,N_13521);
nand U16416 (N_16416,N_12623,N_11691);
nand U16417 (N_16417,N_11933,N_10656);
xnor U16418 (N_16418,N_13702,N_13817);
nor U16419 (N_16419,N_10386,N_12532);
xnor U16420 (N_16420,N_12166,N_11998);
nor U16421 (N_16421,N_14487,N_10975);
or U16422 (N_16422,N_12639,N_11692);
nor U16423 (N_16423,N_12980,N_14341);
nand U16424 (N_16424,N_12970,N_11844);
xor U16425 (N_16425,N_12448,N_10301);
nand U16426 (N_16426,N_11095,N_12048);
xor U16427 (N_16427,N_12062,N_14070);
nor U16428 (N_16428,N_14639,N_11736);
xnor U16429 (N_16429,N_14914,N_11309);
nand U16430 (N_16430,N_13320,N_13902);
nor U16431 (N_16431,N_12309,N_10084);
nor U16432 (N_16432,N_13733,N_10469);
and U16433 (N_16433,N_10900,N_11262);
nor U16434 (N_16434,N_14145,N_11755);
and U16435 (N_16435,N_12799,N_10754);
nand U16436 (N_16436,N_13155,N_14883);
nand U16437 (N_16437,N_13981,N_10345);
or U16438 (N_16438,N_14369,N_12886);
nor U16439 (N_16439,N_13149,N_14302);
nor U16440 (N_16440,N_11846,N_10287);
nor U16441 (N_16441,N_11676,N_10410);
nor U16442 (N_16442,N_12516,N_13675);
xnor U16443 (N_16443,N_14203,N_13206);
nor U16444 (N_16444,N_10706,N_10899);
or U16445 (N_16445,N_10936,N_12708);
or U16446 (N_16446,N_14324,N_10130);
and U16447 (N_16447,N_12421,N_11103);
nand U16448 (N_16448,N_11016,N_10160);
nor U16449 (N_16449,N_13526,N_10554);
nor U16450 (N_16450,N_12783,N_13103);
or U16451 (N_16451,N_10970,N_13944);
nor U16452 (N_16452,N_14214,N_10335);
or U16453 (N_16453,N_10583,N_14874);
or U16454 (N_16454,N_13739,N_13133);
nor U16455 (N_16455,N_10574,N_10760);
and U16456 (N_16456,N_13461,N_12971);
xnor U16457 (N_16457,N_12051,N_14267);
nand U16458 (N_16458,N_13517,N_14513);
xnor U16459 (N_16459,N_14863,N_11576);
and U16460 (N_16460,N_13250,N_14268);
nor U16461 (N_16461,N_14204,N_14181);
and U16462 (N_16462,N_11548,N_13289);
or U16463 (N_16463,N_13512,N_14506);
xnor U16464 (N_16464,N_10620,N_14927);
nor U16465 (N_16465,N_13073,N_12192);
nand U16466 (N_16466,N_12973,N_11619);
nand U16467 (N_16467,N_14168,N_10655);
nand U16468 (N_16468,N_14189,N_14157);
nand U16469 (N_16469,N_10190,N_14207);
nor U16470 (N_16470,N_13221,N_11493);
and U16471 (N_16471,N_10716,N_13175);
and U16472 (N_16472,N_13794,N_10414);
and U16473 (N_16473,N_12808,N_13087);
and U16474 (N_16474,N_12839,N_14474);
nand U16475 (N_16475,N_11157,N_13402);
xor U16476 (N_16476,N_12024,N_10874);
or U16477 (N_16477,N_10565,N_14152);
or U16478 (N_16478,N_11860,N_14273);
and U16479 (N_16479,N_13010,N_13623);
nor U16480 (N_16480,N_12152,N_12481);
or U16481 (N_16481,N_14718,N_12110);
xnor U16482 (N_16482,N_10054,N_12328);
nand U16483 (N_16483,N_13390,N_14600);
xnor U16484 (N_16484,N_14137,N_14163);
nor U16485 (N_16485,N_14775,N_12559);
nor U16486 (N_16486,N_10254,N_13199);
nor U16487 (N_16487,N_14188,N_10052);
or U16488 (N_16488,N_14006,N_14986);
nor U16489 (N_16489,N_12403,N_13756);
and U16490 (N_16490,N_14281,N_14138);
and U16491 (N_16491,N_13356,N_11053);
and U16492 (N_16492,N_10226,N_14556);
and U16493 (N_16493,N_13219,N_14548);
xnor U16494 (N_16494,N_10725,N_14000);
or U16495 (N_16495,N_12022,N_14295);
or U16496 (N_16496,N_10286,N_11126);
nor U16497 (N_16497,N_14493,N_14867);
xnor U16498 (N_16498,N_10012,N_10450);
and U16499 (N_16499,N_11407,N_11357);
xor U16500 (N_16500,N_11458,N_10393);
or U16501 (N_16501,N_13104,N_11492);
or U16502 (N_16502,N_14202,N_14900);
and U16503 (N_16503,N_14041,N_11479);
xnor U16504 (N_16504,N_13759,N_11013);
or U16505 (N_16505,N_14198,N_12909);
and U16506 (N_16506,N_14479,N_13905);
nor U16507 (N_16507,N_11866,N_11032);
xnor U16508 (N_16508,N_12727,N_12533);
or U16509 (N_16509,N_13861,N_10411);
xnor U16510 (N_16510,N_11253,N_12667);
or U16511 (N_16511,N_10199,N_10376);
or U16512 (N_16512,N_13565,N_12990);
and U16513 (N_16513,N_11044,N_10572);
and U16514 (N_16514,N_12122,N_12373);
or U16515 (N_16515,N_11165,N_12788);
nand U16516 (N_16516,N_14003,N_11152);
nand U16517 (N_16517,N_14491,N_12266);
and U16518 (N_16518,N_13420,N_12311);
and U16519 (N_16519,N_12239,N_10515);
or U16520 (N_16520,N_12036,N_14480);
and U16521 (N_16521,N_13202,N_13045);
xor U16522 (N_16522,N_12228,N_14252);
or U16523 (N_16523,N_14337,N_12670);
and U16524 (N_16524,N_11371,N_10635);
xor U16525 (N_16525,N_11754,N_13487);
nand U16526 (N_16526,N_12234,N_10739);
and U16527 (N_16527,N_14247,N_10486);
and U16528 (N_16528,N_13628,N_12431);
nand U16529 (N_16529,N_12422,N_14552);
nand U16530 (N_16530,N_14501,N_10296);
or U16531 (N_16531,N_11615,N_12225);
or U16532 (N_16532,N_14158,N_13385);
nor U16533 (N_16533,N_13243,N_13265);
xor U16534 (N_16534,N_14536,N_13009);
and U16535 (N_16535,N_13474,N_13594);
nor U16536 (N_16536,N_10509,N_13726);
and U16537 (N_16537,N_10188,N_13311);
nand U16538 (N_16538,N_11445,N_11896);
nand U16539 (N_16539,N_13280,N_14707);
xor U16540 (N_16540,N_10427,N_14689);
nand U16541 (N_16541,N_14891,N_14370);
nor U16542 (N_16542,N_11019,N_14329);
and U16543 (N_16543,N_14540,N_14844);
nor U16544 (N_16544,N_12650,N_14704);
nand U16545 (N_16545,N_12132,N_12865);
and U16546 (N_16546,N_13969,N_14848);
or U16547 (N_16547,N_14144,N_11605);
or U16548 (N_16548,N_12850,N_10955);
nand U16549 (N_16549,N_10730,N_10094);
xor U16550 (N_16550,N_12387,N_14338);
nor U16551 (N_16551,N_14999,N_10168);
or U16552 (N_16552,N_13416,N_13462);
or U16553 (N_16553,N_13274,N_14836);
nor U16554 (N_16554,N_12359,N_14349);
nor U16555 (N_16555,N_12124,N_12565);
xnor U16556 (N_16556,N_12964,N_11683);
nand U16557 (N_16557,N_10593,N_13237);
or U16558 (N_16558,N_14021,N_10829);
nor U16559 (N_16559,N_11036,N_11595);
xor U16560 (N_16560,N_10872,N_11006);
xor U16561 (N_16561,N_13828,N_13669);
or U16562 (N_16562,N_12534,N_14027);
nor U16563 (N_16563,N_12374,N_12322);
nand U16564 (N_16564,N_14995,N_12492);
and U16565 (N_16565,N_12308,N_11133);
nor U16566 (N_16566,N_10114,N_11245);
nor U16567 (N_16567,N_11724,N_14249);
and U16568 (N_16568,N_10462,N_12613);
nand U16569 (N_16569,N_12280,N_12502);
and U16570 (N_16570,N_14571,N_13535);
and U16571 (N_16571,N_12699,N_10026);
nor U16572 (N_16572,N_14782,N_13564);
nor U16573 (N_16573,N_11547,N_10481);
or U16574 (N_16574,N_10538,N_11612);
xor U16575 (N_16575,N_14859,N_11333);
or U16576 (N_16576,N_12077,N_14856);
xor U16577 (N_16577,N_14002,N_10723);
xnor U16578 (N_16578,N_11403,N_13629);
or U16579 (N_16579,N_14033,N_10920);
or U16580 (N_16580,N_10201,N_11930);
and U16581 (N_16581,N_11816,N_11804);
or U16582 (N_16582,N_14299,N_14465);
nor U16583 (N_16583,N_10470,N_11575);
and U16584 (N_16584,N_14603,N_12730);
nor U16585 (N_16585,N_11802,N_13330);
nor U16586 (N_16586,N_14843,N_12008);
nand U16587 (N_16587,N_11001,N_14195);
and U16588 (N_16588,N_10431,N_12734);
and U16589 (N_16589,N_10321,N_14721);
nor U16590 (N_16590,N_12283,N_12860);
nand U16591 (N_16591,N_14998,N_12303);
or U16592 (N_16592,N_12713,N_13930);
or U16593 (N_16593,N_13516,N_14054);
and U16594 (N_16594,N_11216,N_11689);
xnor U16595 (N_16595,N_11217,N_13392);
nor U16596 (N_16596,N_12646,N_11047);
or U16597 (N_16597,N_12842,N_13583);
xnor U16598 (N_16598,N_13942,N_11909);
nand U16599 (N_16599,N_13020,N_10006);
or U16600 (N_16600,N_14313,N_13533);
or U16601 (N_16601,N_11342,N_13954);
and U16602 (N_16602,N_14641,N_10561);
nand U16603 (N_16603,N_11178,N_14935);
xor U16604 (N_16604,N_11611,N_11190);
nand U16605 (N_16605,N_12097,N_13459);
xor U16606 (N_16606,N_13352,N_14755);
or U16607 (N_16607,N_10476,N_13225);
xor U16608 (N_16608,N_14421,N_13262);
nor U16609 (N_16609,N_14572,N_12567);
or U16610 (N_16610,N_12116,N_13641);
nand U16611 (N_16611,N_14731,N_12101);
xnor U16612 (N_16612,N_13354,N_11513);
and U16613 (N_16613,N_12148,N_11313);
or U16614 (N_16614,N_11845,N_14717);
nor U16615 (N_16615,N_13322,N_10823);
and U16616 (N_16616,N_13773,N_13893);
or U16617 (N_16617,N_10770,N_12822);
and U16618 (N_16618,N_10734,N_10537);
nor U16619 (N_16619,N_11404,N_10408);
and U16620 (N_16620,N_14928,N_11465);
nor U16621 (N_16621,N_12489,N_11564);
xor U16622 (N_16622,N_11600,N_10436);
and U16623 (N_16623,N_11874,N_13632);
xor U16624 (N_16624,N_12879,N_11744);
nor U16625 (N_16625,N_11751,N_14196);
or U16626 (N_16626,N_13938,N_14686);
xnor U16627 (N_16627,N_10678,N_14316);
nor U16628 (N_16628,N_13493,N_13233);
or U16629 (N_16629,N_11048,N_11467);
or U16630 (N_16630,N_14660,N_14748);
or U16631 (N_16631,N_12104,N_12495);
nor U16632 (N_16632,N_12034,N_13819);
and U16633 (N_16633,N_13927,N_13534);
xor U16634 (N_16634,N_14435,N_14171);
nand U16635 (N_16635,N_13111,N_12666);
nand U16636 (N_16636,N_10268,N_11454);
nand U16637 (N_16637,N_12113,N_12499);
nand U16638 (N_16638,N_13788,N_12908);
nor U16639 (N_16639,N_11878,N_12921);
xor U16640 (N_16640,N_14336,N_10805);
xnor U16641 (N_16641,N_11967,N_11159);
nor U16642 (N_16642,N_12250,N_10867);
and U16643 (N_16643,N_14781,N_10508);
xor U16644 (N_16644,N_13834,N_10487);
xor U16645 (N_16645,N_10384,N_11320);
or U16646 (N_16646,N_13842,N_14071);
and U16647 (N_16647,N_10803,N_10744);
xor U16648 (N_16648,N_10142,N_14284);
and U16649 (N_16649,N_14631,N_14122);
nand U16650 (N_16650,N_10957,N_12540);
nor U16651 (N_16651,N_12245,N_13578);
and U16652 (N_16652,N_14221,N_11160);
nor U16653 (N_16653,N_10623,N_10594);
or U16654 (N_16654,N_12959,N_13211);
nand U16655 (N_16655,N_11500,N_11883);
nand U16656 (N_16656,N_13803,N_10016);
nand U16657 (N_16657,N_11099,N_14476);
nand U16658 (N_16658,N_11135,N_12156);
nor U16659 (N_16659,N_13531,N_13548);
xnor U16660 (N_16660,N_10417,N_11621);
nor U16661 (N_16661,N_11929,N_12827);
nand U16662 (N_16662,N_14744,N_14457);
xor U16663 (N_16663,N_13825,N_12998);
or U16664 (N_16664,N_10049,N_13478);
xor U16665 (N_16665,N_12216,N_12659);
nor U16666 (N_16666,N_12223,N_11757);
nor U16667 (N_16667,N_11892,N_13331);
nand U16668 (N_16668,N_13760,N_12226);
or U16669 (N_16669,N_10366,N_11738);
xor U16670 (N_16670,N_14266,N_13734);
nor U16671 (N_16671,N_12174,N_13035);
or U16672 (N_16672,N_12458,N_12837);
nor U16673 (N_16673,N_13546,N_12437);
nand U16674 (N_16674,N_14431,N_14652);
and U16675 (N_16675,N_11964,N_12805);
or U16676 (N_16676,N_12366,N_14984);
nor U16677 (N_16677,N_11668,N_12714);
and U16678 (N_16678,N_10710,N_13276);
nand U16679 (N_16679,N_12100,N_14681);
nand U16680 (N_16680,N_10189,N_14470);
nor U16681 (N_16681,N_13846,N_14936);
and U16682 (N_16682,N_10840,N_13644);
nor U16683 (N_16683,N_10073,N_12285);
or U16684 (N_16684,N_12902,N_10985);
nor U16685 (N_16685,N_10318,N_11991);
and U16686 (N_16686,N_10050,N_11780);
xor U16687 (N_16687,N_10162,N_13374);
and U16688 (N_16688,N_14777,N_11795);
nand U16689 (N_16689,N_11781,N_13471);
or U16690 (N_16690,N_11075,N_13357);
xor U16691 (N_16691,N_13991,N_14970);
or U16692 (N_16692,N_14509,N_13624);
nor U16693 (N_16693,N_12840,N_14034);
and U16694 (N_16694,N_11123,N_14598);
or U16695 (N_16695,N_12436,N_13791);
nand U16696 (N_16696,N_12917,N_13097);
nand U16697 (N_16697,N_13750,N_11186);
nand U16698 (N_16698,N_10083,N_11655);
nor U16699 (N_16699,N_10550,N_13769);
nand U16700 (N_16700,N_14445,N_12758);
xor U16701 (N_16701,N_14621,N_14391);
nand U16702 (N_16702,N_11149,N_12535);
nor U16703 (N_16703,N_13304,N_14982);
nor U16704 (N_16704,N_14227,N_11241);
nand U16705 (N_16705,N_11915,N_13719);
nor U16706 (N_16706,N_10074,N_14880);
and U16707 (N_16707,N_13179,N_11809);
or U16708 (N_16708,N_12074,N_10546);
or U16709 (N_16709,N_10444,N_13409);
xnor U16710 (N_16710,N_11918,N_10392);
and U16711 (N_16711,N_13369,N_12348);
or U16712 (N_16712,N_12942,N_10283);
or U16713 (N_16713,N_14976,N_11440);
xor U16714 (N_16714,N_14064,N_13974);
nand U16715 (N_16715,N_10139,N_14190);
nand U16716 (N_16716,N_10341,N_14061);
xor U16717 (N_16717,N_11604,N_10772);
and U16718 (N_16718,N_12269,N_11317);
or U16719 (N_16719,N_14764,N_13001);
or U16720 (N_16720,N_10184,N_14228);
or U16721 (N_16721,N_14629,N_13247);
nand U16722 (N_16722,N_11416,N_11385);
nor U16723 (N_16723,N_14524,N_11530);
and U16724 (N_16724,N_10516,N_12286);
xnor U16725 (N_16725,N_10252,N_11833);
nand U16726 (N_16726,N_10600,N_13100);
or U16727 (N_16727,N_10330,N_11944);
nand U16728 (N_16728,N_10674,N_10000);
and U16729 (N_16729,N_14032,N_13368);
and U16730 (N_16730,N_10643,N_13904);
nand U16731 (N_16731,N_14432,N_13136);
or U16732 (N_16732,N_11422,N_14343);
nand U16733 (N_16733,N_10497,N_14478);
xor U16734 (N_16734,N_14983,N_13407);
nand U16735 (N_16735,N_10929,N_10884);
or U16736 (N_16736,N_12017,N_13688);
and U16737 (N_16737,N_14762,N_13170);
nor U16738 (N_16738,N_10008,N_11840);
nor U16739 (N_16739,N_14406,N_10940);
xor U16740 (N_16740,N_14237,N_11826);
nand U16741 (N_16741,N_14802,N_10119);
nand U16742 (N_16742,N_14260,N_13917);
or U16743 (N_16743,N_13456,N_10591);
xor U16744 (N_16744,N_14646,N_11279);
nor U16745 (N_16745,N_12169,N_10818);
or U16746 (N_16746,N_13977,N_13949);
or U16747 (N_16747,N_13708,N_10877);
or U16748 (N_16748,N_12800,N_14327);
xnor U16749 (N_16749,N_11187,N_10165);
nand U16750 (N_16750,N_11076,N_13671);
and U16751 (N_16751,N_11793,N_13868);
and U16752 (N_16752,N_11218,N_11545);
nor U16753 (N_16753,N_11956,N_12211);
and U16754 (N_16754,N_12899,N_12161);
nand U16755 (N_16755,N_10822,N_10923);
or U16756 (N_16756,N_11319,N_14458);
or U16757 (N_16757,N_10288,N_13880);
or U16758 (N_16758,N_14182,N_13436);
nand U16759 (N_16759,N_13055,N_12037);
nand U16760 (N_16760,N_12701,N_13099);
xor U16761 (N_16761,N_12987,N_11043);
nand U16762 (N_16762,N_12968,N_12672);
or U16763 (N_16763,N_11979,N_14684);
xor U16764 (N_16764,N_12793,N_10749);
nor U16765 (N_16765,N_14143,N_11203);
nor U16766 (N_16766,N_12361,N_10584);
and U16767 (N_16767,N_11753,N_10511);
xnor U16768 (N_16768,N_10042,N_14774);
nor U16769 (N_16769,N_13718,N_13699);
nor U16770 (N_16770,N_13598,N_12370);
xnor U16771 (N_16771,N_14602,N_11782);
nand U16772 (N_16772,N_10459,N_12232);
nand U16773 (N_16773,N_13572,N_10501);
and U16774 (N_16774,N_12120,N_11064);
nand U16775 (N_16775,N_12912,N_10361);
nand U16776 (N_16776,N_12020,N_10173);
xnor U16777 (N_16777,N_11864,N_12866);
and U16778 (N_16778,N_13115,N_13150);
xnor U16779 (N_16779,N_11034,N_13248);
nand U16780 (N_16780,N_12679,N_11603);
or U16781 (N_16781,N_14753,N_11561);
or U16782 (N_16782,N_10202,N_11601);
nor U16783 (N_16783,N_14931,N_13340);
nand U16784 (N_16784,N_13856,N_10239);
xnor U16785 (N_16785,N_14385,N_10152);
nor U16786 (N_16786,N_13064,N_11435);
xor U16787 (N_16787,N_12114,N_12992);
and U16788 (N_16788,N_11120,N_12198);
nor U16789 (N_16789,N_12538,N_14708);
or U16790 (N_16790,N_13334,N_14876);
nor U16791 (N_16791,N_11266,N_12491);
or U16792 (N_16792,N_12836,N_14820);
nor U16793 (N_16793,N_10549,N_12086);
nor U16794 (N_16794,N_12469,N_13785);
nor U16795 (N_16795,N_14429,N_10610);
nand U16796 (N_16796,N_10502,N_13855);
and U16797 (N_16797,N_10914,N_13672);
nor U16798 (N_16798,N_11337,N_12300);
nand U16799 (N_16799,N_11978,N_13523);
or U16800 (N_16800,N_11912,N_10369);
and U16801 (N_16801,N_10994,N_12183);
or U16802 (N_16802,N_13654,N_12289);
nor U16803 (N_16803,N_13080,N_14586);
nand U16804 (N_16804,N_11977,N_14439);
and U16805 (N_16805,N_12963,N_10081);
and U16806 (N_16806,N_13585,N_14816);
nand U16807 (N_16807,N_14955,N_11511);
nand U16808 (N_16808,N_14467,N_12305);
nor U16809 (N_16809,N_13820,N_14542);
xnor U16810 (N_16810,N_13213,N_12272);
and U16811 (N_16811,N_11726,N_14292);
nand U16812 (N_16812,N_10303,N_11828);
nand U16813 (N_16813,N_13556,N_13697);
nand U16814 (N_16814,N_14289,N_13295);
nand U16815 (N_16815,N_11373,N_14126);
or U16816 (N_16816,N_13589,N_13689);
or U16817 (N_16817,N_12012,N_12433);
nor U16818 (N_16818,N_11290,N_11232);
or U16819 (N_16819,N_10498,N_10215);
or U16820 (N_16820,N_13818,N_10613);
or U16821 (N_16821,N_12107,N_13445);
or U16822 (N_16822,N_14076,N_11810);
nor U16823 (N_16823,N_14987,N_12979);
and U16824 (N_16824,N_14087,N_11558);
or U16825 (N_16825,N_10167,N_12736);
and U16826 (N_16826,N_14216,N_11292);
xnor U16827 (N_16827,N_11926,N_13867);
nand U16828 (N_16828,N_10962,N_11835);
and U16829 (N_16829,N_12604,N_14262);
xnor U16830 (N_16830,N_11080,N_11675);
xor U16831 (N_16831,N_12380,N_14306);
or U16832 (N_16832,N_10247,N_12989);
and U16833 (N_16833,N_12408,N_10343);
xor U16834 (N_16834,N_14257,N_13603);
and U16835 (N_16835,N_10178,N_12197);
xnor U16836 (N_16836,N_13570,N_10246);
nand U16837 (N_16837,N_13763,N_14892);
xnor U16838 (N_16838,N_12331,N_10099);
nor U16839 (N_16839,N_10717,N_13805);
and U16840 (N_16840,N_14895,N_13912);
nor U16841 (N_16841,N_11680,N_14134);
nand U16842 (N_16842,N_14496,N_10363);
xor U16843 (N_16843,N_13994,N_12367);
xnor U16844 (N_16844,N_12307,N_12368);
xor U16845 (N_16845,N_11941,N_11223);
xor U16846 (N_16846,N_10331,N_11000);
and U16847 (N_16847,N_12910,N_11031);
nand U16848 (N_16848,N_11429,N_10011);
or U16849 (N_16849,N_12026,N_12461);
or U16850 (N_16850,N_14455,N_13249);
nor U16851 (N_16851,N_13158,N_12383);
nor U16852 (N_16852,N_12598,N_12796);
nand U16853 (N_16853,N_13191,N_10888);
nor U16854 (N_16854,N_10022,N_11551);
and U16855 (N_16855,N_12375,N_12764);
xor U16856 (N_16856,N_11413,N_12416);
xor U16857 (N_16857,N_14503,N_13004);
or U16858 (N_16858,N_13296,N_10691);
xor U16859 (N_16859,N_13833,N_12324);
and U16860 (N_16860,N_12414,N_10175);
and U16861 (N_16861,N_11409,N_11806);
and U16862 (N_16862,N_13382,N_12791);
nand U16863 (N_16863,N_14218,N_10830);
or U16864 (N_16864,N_11071,N_13047);
nand U16865 (N_16865,N_13078,N_13622);
or U16866 (N_16866,N_11322,N_13633);
nand U16867 (N_16867,N_14942,N_14366);
or U16868 (N_16868,N_14561,N_14193);
or U16869 (N_16869,N_12618,N_14233);
nor U16870 (N_16870,N_11579,N_11512);
xor U16871 (N_16871,N_14723,N_12419);
and U16872 (N_16872,N_12220,N_14591);
and U16873 (N_16873,N_13286,N_10663);
xnor U16874 (N_16874,N_10091,N_10590);
or U16875 (N_16875,N_10533,N_13207);
xor U16876 (N_16876,N_11788,N_14376);
or U16877 (N_16877,N_11654,N_11642);
or U16878 (N_16878,N_11263,N_13591);
nand U16879 (N_16879,N_11472,N_11483);
or U16880 (N_16880,N_12396,N_14569);
and U16881 (N_16881,N_11613,N_14726);
nor U16882 (N_16882,N_13451,N_12947);
nand U16883 (N_16883,N_11381,N_10898);
nand U16884 (N_16884,N_14019,N_14167);
xor U16885 (N_16885,N_11830,N_11026);
nor U16886 (N_16886,N_12647,N_13141);
nand U16887 (N_16887,N_11531,N_13037);
nor U16888 (N_16888,N_12000,N_13437);
and U16889 (N_16889,N_10958,N_11923);
and U16890 (N_16890,N_12126,N_10364);
and U16891 (N_16891,N_13900,N_10698);
and U16892 (N_16892,N_11723,N_11533);
and U16893 (N_16893,N_14136,N_14308);
xnor U16894 (N_16894,N_12521,N_10931);
or U16895 (N_16895,N_11871,N_10051);
nor U16896 (N_16896,N_10573,N_11379);
nand U16897 (N_16897,N_13387,N_14441);
nor U16898 (N_16898,N_10180,N_10346);
or U16899 (N_16899,N_12614,N_12263);
nor U16900 (N_16900,N_10557,N_11023);
and U16901 (N_16901,N_14943,N_14523);
xor U16902 (N_16902,N_14079,N_10186);
nand U16903 (N_16903,N_14674,N_14648);
nand U16904 (N_16904,N_12117,N_10638);
and U16905 (N_16905,N_12584,N_11163);
nand U16906 (N_16906,N_11068,N_11887);
nand U16907 (N_16907,N_10633,N_10164);
or U16908 (N_16908,N_13203,N_14701);
nor U16909 (N_16909,N_14832,N_11897);
and U16910 (N_16910,N_10217,N_13036);
and U16911 (N_16911,N_10776,N_14852);
and U16912 (N_16912,N_12347,N_14397);
nand U16913 (N_16913,N_12922,N_10668);
xnor U16914 (N_16914,N_14830,N_10372);
xor U16915 (N_16915,N_11517,N_12660);
or U16916 (N_16916,N_11090,N_13599);
or U16917 (N_16917,N_10897,N_13397);
and U16918 (N_16918,N_10534,N_14988);
nor U16919 (N_16919,N_12641,N_12944);
nor U16920 (N_16920,N_12498,N_14169);
and U16921 (N_16921,N_14770,N_12080);
nand U16922 (N_16922,N_11247,N_13217);
nand U16923 (N_16923,N_10430,N_12168);
nand U16924 (N_16924,N_13941,N_13063);
xnor U16925 (N_16925,N_10294,N_10171);
xor U16926 (N_16926,N_14384,N_12925);
nor U16927 (N_16927,N_14862,N_13391);
or U16928 (N_16928,N_13968,N_12719);
nand U16929 (N_16929,N_13698,N_14685);
nor U16930 (N_16930,N_11763,N_13163);
and U16931 (N_16931,N_11332,N_13776);
or U16932 (N_16932,N_12177,N_10930);
and U16933 (N_16933,N_12424,N_14593);
nand U16934 (N_16934,N_12494,N_13853);
or U16935 (N_16935,N_13252,N_14594);
or U16936 (N_16936,N_12932,N_10980);
and U16937 (N_16937,N_10098,N_13338);
or U16938 (N_16938,N_10787,N_10027);
nand U16939 (N_16939,N_14360,N_14109);
xnor U16940 (N_16940,N_13960,N_13110);
and U16941 (N_16941,N_10395,N_13328);
and U16942 (N_16942,N_14025,N_11100);
and U16943 (N_16943,N_12931,N_12716);
xor U16944 (N_16944,N_11065,N_14925);
nor U16945 (N_16945,N_13656,N_10336);
nand U16946 (N_16946,N_12093,N_12290);
and U16947 (N_16947,N_11177,N_10641);
or U16948 (N_16948,N_10514,N_13480);
nand U16949 (N_16949,N_13479,N_13758);
nand U16950 (N_16950,N_11988,N_10903);
nor U16951 (N_16951,N_14607,N_14442);
xor U16952 (N_16952,N_13588,N_14950);
and U16953 (N_16953,N_13355,N_11815);
and U16954 (N_16954,N_12658,N_14213);
xor U16955 (N_16955,N_13460,N_14785);
nand U16956 (N_16956,N_10831,N_10382);
nand U16957 (N_16957,N_14750,N_13959);
nand U16958 (N_16958,N_11124,N_10063);
nor U16959 (N_16959,N_13524,N_14447);
and U16960 (N_16960,N_12033,N_13690);
and U16961 (N_16961,N_12616,N_10265);
and U16962 (N_16962,N_10759,N_14544);
or U16963 (N_16963,N_14154,N_11224);
nand U16964 (N_16964,N_12956,N_11769);
or U16965 (N_16965,N_11770,N_14250);
and U16966 (N_16966,N_10030,N_10701);
nand U16967 (N_16967,N_11858,N_12090);
xor U16968 (N_16968,N_14659,N_12338);
or U16969 (N_16969,N_11760,N_12246);
and U16970 (N_16970,N_14894,N_13727);
and U16971 (N_16971,N_11480,N_12546);
or U16972 (N_16972,N_10367,N_13172);
and U16973 (N_16973,N_13298,N_12896);
xor U16974 (N_16974,N_14546,N_12135);
nand U16975 (N_16975,N_11525,N_10004);
and U16976 (N_16976,N_14771,N_14434);
xor U16977 (N_16977,N_11853,N_10131);
and U16978 (N_16978,N_13775,N_10774);
and U16979 (N_16979,N_11477,N_12125);
xor U16980 (N_16980,N_10621,N_10108);
nor U16981 (N_16981,N_11839,N_10952);
or U16982 (N_16982,N_13952,N_14130);
or U16983 (N_16983,N_14688,N_14449);
nand U16984 (N_16984,N_14318,N_12617);
or U16985 (N_16985,N_13812,N_11520);
or U16986 (N_16986,N_12585,N_11136);
nand U16987 (N_16987,N_10727,N_11886);
and U16988 (N_16988,N_14112,N_13715);
or U16989 (N_16989,N_10100,N_14119);
and U16990 (N_16990,N_12889,N_10062);
nand U16991 (N_16991,N_14617,N_13933);
or U16992 (N_16992,N_10238,N_12329);
nor U16993 (N_16993,N_13786,N_12553);
nand U16994 (N_16994,N_14903,N_12454);
or U16995 (N_16995,N_10380,N_10865);
nand U16996 (N_16996,N_11275,N_13932);
nand U16997 (N_16997,N_11092,N_11482);
nor U16998 (N_16998,N_10916,N_12610);
xnor U16999 (N_16999,N_14691,N_14578);
xnor U17000 (N_17000,N_11081,N_11851);
xor U17001 (N_17001,N_12205,N_14505);
nor U17002 (N_17002,N_11369,N_12440);
and U17003 (N_17003,N_13285,N_10455);
or U17004 (N_17004,N_12611,N_14469);
or U17005 (N_17005,N_14780,N_12846);
and U17006 (N_17006,N_11761,N_11669);
or U17007 (N_17007,N_14804,N_10758);
nand U17008 (N_17008,N_13176,N_12314);
xor U17009 (N_17009,N_13787,N_10695);
nor U17010 (N_17010,N_10274,N_10018);
nand U17011 (N_17011,N_10485,N_12703);
or U17012 (N_17012,N_14595,N_10685);
nor U17013 (N_17013,N_13972,N_14351);
nand U17014 (N_17014,N_12885,N_13444);
or U17015 (N_17015,N_11063,N_14751);
and U17016 (N_17016,N_10642,N_14415);
or U17017 (N_17017,N_10253,N_14620);
nor U17018 (N_17018,N_12900,N_12406);
nand U17019 (N_17019,N_12864,N_11812);
or U17020 (N_17020,N_11046,N_12709);
xor U17021 (N_17021,N_10045,N_12410);
nand U17022 (N_17022,N_13118,N_11971);
or U17023 (N_17023,N_13349,N_11436);
nor U17024 (N_17024,N_11556,N_10496);
and U17025 (N_17025,N_10747,N_10271);
xor U17026 (N_17026,N_11258,N_12833);
nand U17027 (N_17027,N_14073,N_11772);
xnor U17028 (N_17028,N_14298,N_14570);
nand U17029 (N_17029,N_12586,N_14481);
nor U17030 (N_17030,N_14962,N_13337);
xnor U17031 (N_17031,N_12771,N_11861);
or U17032 (N_17032,N_13529,N_11557);
xor U17033 (N_17033,N_12936,N_10795);
nor U17034 (N_17034,N_14017,N_10851);
nor U17035 (N_17035,N_14653,N_13841);
nor U17036 (N_17036,N_11008,N_10507);
nor U17037 (N_17037,N_12295,N_11115);
xnor U17038 (N_17038,N_10570,N_10984);
xnor U17039 (N_17039,N_10176,N_11382);
nor U17040 (N_17040,N_10046,N_11661);
xnor U17041 (N_17041,N_10585,N_13597);
nand U17042 (N_17042,N_12766,N_12506);
xor U17043 (N_17043,N_12450,N_14796);
nand U17044 (N_17044,N_10150,N_10235);
or U17045 (N_17045,N_10837,N_13924);
and U17046 (N_17046,N_10828,N_11863);
and U17047 (N_17047,N_11174,N_11910);
or U17048 (N_17048,N_13703,N_14706);
xor U17049 (N_17049,N_10403,N_12606);
nor U17050 (N_17050,N_12543,N_12678);
nand U17051 (N_17051,N_10258,N_13986);
nor U17052 (N_17052,N_13030,N_13692);
and U17053 (N_17053,N_14129,N_12178);
xnor U17054 (N_17054,N_13705,N_12742);
or U17055 (N_17055,N_11252,N_10110);
nand U17056 (N_17056,N_10269,N_14450);
xnor U17057 (N_17057,N_11847,N_10304);
nor U17058 (N_17058,N_11521,N_13305);
nand U17059 (N_17059,N_14850,N_12872);
xnor U17060 (N_17060,N_11565,N_10558);
xnor U17061 (N_17061,N_10567,N_11758);
nor U17062 (N_17062,N_10943,N_11842);
or U17063 (N_17063,N_13287,N_14378);
nor U17064 (N_17064,N_13886,N_10209);
and U17065 (N_17065,N_12888,N_11356);
nor U17066 (N_17066,N_10627,N_13130);
nand U17067 (N_17067,N_13720,N_13293);
or U17068 (N_17068,N_12577,N_10475);
nand U17069 (N_17069,N_14282,N_12032);
and U17070 (N_17070,N_10154,N_14604);
and U17071 (N_17071,N_10731,N_11484);
and U17072 (N_17072,N_10494,N_12179);
xor U17073 (N_17073,N_10290,N_13813);
xor U17074 (N_17074,N_11756,N_14919);
and U17075 (N_17075,N_10029,N_11921);
or U17076 (N_17076,N_11902,N_14776);
nand U17077 (N_17077,N_11623,N_12055);
xor U17078 (N_17078,N_13731,N_14767);
xor U17079 (N_17079,N_13024,N_14240);
nor U17080 (N_17080,N_14766,N_11206);
and U17081 (N_17081,N_14090,N_12640);
or U17082 (N_17082,N_13871,N_12803);
and U17083 (N_17083,N_12229,N_11336);
nor U17084 (N_17084,N_10667,N_13254);
or U17085 (N_17085,N_11982,N_14683);
or U17086 (N_17086,N_12644,N_14833);
xnor U17087 (N_17087,N_12203,N_11110);
and U17088 (N_17088,N_10978,N_11916);
and U17089 (N_17089,N_14172,N_14462);
or U17090 (N_17090,N_10792,N_12769);
or U17091 (N_17091,N_12291,N_10203);
xnor U17092 (N_17092,N_14269,N_12451);
and U17093 (N_17093,N_10784,N_10704);
nor U17094 (N_17094,N_13831,N_14013);
and U17095 (N_17095,N_14466,N_13807);
and U17096 (N_17096,N_12630,N_12484);
nor U17097 (N_17097,N_14547,N_10586);
and U17098 (N_17098,N_11800,N_13255);
nor U17099 (N_17099,N_10197,N_11202);
or U17100 (N_17100,N_12542,N_13725);
nand U17101 (N_17101,N_14359,N_13696);
nor U17102 (N_17102,N_11592,N_13677);
and U17103 (N_17103,N_11594,N_14897);
nand U17104 (N_17104,N_11003,N_14149);
or U17105 (N_17105,N_13081,N_12838);
or U17106 (N_17106,N_13797,N_11901);
nor U17107 (N_17107,N_12190,N_10319);
or U17108 (N_17108,N_10106,N_11476);
nor U17109 (N_17109,N_11614,N_13278);
or U17110 (N_17110,N_10677,N_11107);
nor U17111 (N_17111,N_10825,N_10133);
nand U17112 (N_17112,N_10111,N_11629);
nand U17113 (N_17113,N_11056,N_14245);
or U17114 (N_17114,N_13208,N_14851);
or U17115 (N_17115,N_14160,N_14577);
nor U17116 (N_17116,N_10272,N_11957);
nor U17117 (N_17117,N_13840,N_13470);
nand U17118 (N_17118,N_13341,N_11468);
nor U17119 (N_17119,N_12241,N_12180);
nand U17120 (N_17120,N_11018,N_11361);
nand U17121 (N_17121,N_13209,N_12044);
nand U17122 (N_17122,N_10562,N_13948);
nor U17123 (N_17123,N_12173,N_10116);
xor U17124 (N_17124,N_14350,N_10264);
or U17125 (N_17125,N_12832,N_13446);
xnor U17126 (N_17126,N_11118,N_10628);
nor U17127 (N_17127,N_10077,N_12873);
nor U17128 (N_17128,N_11239,N_12343);
or U17129 (N_17129,N_11696,N_11877);
and U17130 (N_17130,N_11426,N_13329);
nor U17131 (N_17131,N_12121,N_10337);
nor U17132 (N_17132,N_12961,N_12955);
and U17133 (N_17133,N_14486,N_13541);
nand U17134 (N_17134,N_10407,N_11469);
xor U17135 (N_17135,N_10157,N_11983);
and U17136 (N_17136,N_12654,N_13724);
or U17137 (N_17137,N_13379,N_12685);
xnor U17138 (N_17138,N_14230,N_11702);
or U17139 (N_17139,N_10637,N_12988);
nor U17140 (N_17140,N_10718,N_13889);
nand U17141 (N_17141,N_14410,N_13800);
or U17142 (N_17142,N_13236,N_12326);
and U17143 (N_17143,N_14786,N_13655);
nor U17144 (N_17144,N_14840,N_10640);
xnor U17145 (N_17145,N_13619,N_14180);
and U17146 (N_17146,N_11928,N_13811);
nor U17147 (N_17147,N_10292,N_10849);
nor U17148 (N_17148,N_11597,N_11085);
or U17149 (N_17149,N_10928,N_13827);
xnor U17150 (N_17150,N_14896,N_14255);
xnor U17151 (N_17151,N_11633,N_10722);
or U17152 (N_17152,N_14102,N_14865);
or U17153 (N_17153,N_14426,N_11350);
xor U17154 (N_17154,N_11457,N_13667);
xor U17155 (N_17155,N_10309,N_13139);
and U17156 (N_17156,N_13745,N_11488);
and U17157 (N_17157,N_14333,N_10457);
and U17158 (N_17158,N_12724,N_14637);
nand U17159 (N_17159,N_11848,N_13413);
nor U17160 (N_17160,N_14521,N_12005);
and U17161 (N_17161,N_11363,N_11069);
or U17162 (N_17162,N_10752,N_13061);
nand U17163 (N_17163,N_14745,N_14446);
nand U17164 (N_17164,N_11125,N_12096);
xor U17165 (N_17165,N_11002,N_10259);
xor U17166 (N_17166,N_14953,N_11376);
and U17167 (N_17167,N_10149,N_12651);
and U17168 (N_17168,N_14913,N_11368);
nor U17169 (N_17169,N_14253,N_10968);
nand U17170 (N_17170,N_10748,N_13153);
nor U17171 (N_17171,N_14394,N_11927);
nor U17172 (N_17172,N_11589,N_10140);
and U17173 (N_17173,N_12728,N_10789);
xnor U17174 (N_17174,N_11865,N_10921);
nand U17175 (N_17175,N_13676,N_12145);
or U17176 (N_17176,N_13772,N_13212);
nor U17177 (N_17177,N_11255,N_14526);
nor U17178 (N_17178,N_12052,N_13890);
nand U17179 (N_17179,N_14113,N_10871);
xor U17180 (N_17180,N_10582,N_10992);
xor U17181 (N_17181,N_14722,N_12471);
xor U17182 (N_17182,N_12049,N_13312);
nor U17183 (N_17183,N_10489,N_13277);
and U17184 (N_17184,N_13837,N_11030);
nor U17185 (N_17185,N_14390,N_12268);
nor U17186 (N_17186,N_14606,N_12371);
nor U17187 (N_17187,N_11954,N_12828);
nor U17188 (N_17188,N_12233,N_12797);
nand U17189 (N_17189,N_10939,N_10891);
nor U17190 (N_17190,N_12698,N_13350);
or U17191 (N_17191,N_14634,N_14377);
nor U17192 (N_17192,N_12746,N_13485);
xnor U17193 (N_17193,N_12065,N_14960);
or U17194 (N_17194,N_12208,N_13056);
nor U17195 (N_17195,N_13618,N_11936);
and U17196 (N_17196,N_14107,N_11340);
nand U17197 (N_17197,N_14089,N_13997);
and U17198 (N_17198,N_11931,N_10138);
and U17199 (N_17199,N_11410,N_14765);
and U17200 (N_17200,N_10141,N_13132);
and U17201 (N_17201,N_12974,N_12015);
nand U17202 (N_17202,N_10529,N_13621);
nand U17203 (N_17203,N_12352,N_12147);
nand U17204 (N_17204,N_13706,N_14630);
nand U17205 (N_17205,N_10910,N_12476);
or U17206 (N_17206,N_10078,N_10729);
and U17207 (N_17207,N_12465,N_10735);
or U17208 (N_17208,N_14815,N_11307);
and U17209 (N_17209,N_12355,N_11939);
xnor U17210 (N_17210,N_11234,N_11734);
xor U17211 (N_17211,N_11618,N_13015);
nor U17212 (N_17212,N_10311,N_10125);
nor U17213 (N_17213,N_11318,N_10315);
or U17214 (N_17214,N_10145,N_12898);
and U17215 (N_17215,N_10617,N_14309);
and U17216 (N_17216,N_12946,N_11717);
nand U17217 (N_17217,N_13562,N_14133);
xor U17218 (N_17218,N_10406,N_10895);
and U17219 (N_17219,N_12545,N_10654);
and U17220 (N_17220,N_11953,N_10118);
and U17221 (N_17221,N_10773,N_12811);
nor U17222 (N_17222,N_12877,N_13613);
nor U17223 (N_17223,N_13843,N_12138);
nand U17224 (N_17224,N_12676,N_13449);
nor U17225 (N_17225,N_12883,N_12089);
xnor U17226 (N_17226,N_13336,N_14451);
or U17227 (N_17227,N_10912,N_11035);
nand U17228 (N_17228,N_11516,N_12242);
or U17229 (N_17229,N_12784,N_12894);
nand U17230 (N_17230,N_10482,N_11712);
nor U17231 (N_17231,N_12645,N_14407);
nand U17232 (N_17232,N_13895,N_10262);
or U17233 (N_17233,N_12582,N_10163);
nor U17234 (N_17234,N_11288,N_12372);
nand U17235 (N_17235,N_14522,N_12688);
xnor U17236 (N_17236,N_13181,N_11199);
nand U17237 (N_17237,N_10454,N_13519);
and U17238 (N_17238,N_11540,N_11869);
and U17239 (N_17239,N_10179,N_14529);
nand U17240 (N_17240,N_10686,N_13495);
xnor U17241 (N_17241,N_10982,N_13372);
nand U17242 (N_17242,N_14882,N_11832);
or U17243 (N_17243,N_11119,N_10707);
nor U17244 (N_17244,N_13442,N_14788);
xnor U17245 (N_17245,N_11418,N_11539);
nor U17246 (N_17246,N_13695,N_13687);
nand U17247 (N_17247,N_12857,N_14589);
or U17248 (N_17248,N_12019,N_11652);
and U17249 (N_17249,N_12576,N_11353);
xnor U17250 (N_17250,N_11950,N_12823);
or U17251 (N_17251,N_13220,N_11305);
nor U17252 (N_17252,N_10353,N_11401);
nor U17253 (N_17253,N_14902,N_11424);
or U17254 (N_17254,N_11975,N_14533);
nor U17255 (N_17255,N_13310,N_14736);
and U17256 (N_17256,N_13224,N_12976);
nand U17257 (N_17257,N_12692,N_13709);
nand U17258 (N_17258,N_10676,N_11715);
nand U17259 (N_17259,N_13982,N_10293);
xor U17260 (N_17260,N_12715,N_13765);
nor U17261 (N_17261,N_10606,N_11301);
or U17262 (N_17262,N_14640,N_11820);
nor U17263 (N_17263,N_12154,N_14238);
and U17264 (N_17264,N_13916,N_13069);
nor U17265 (N_17265,N_14956,N_11803);
xor U17266 (N_17266,N_10207,N_13244);
nor U17267 (N_17267,N_12217,N_12705);
nor U17268 (N_17268,N_14278,N_13751);
or U17269 (N_17269,N_10310,N_11811);
nand U17270 (N_17270,N_13028,N_10732);
nand U17271 (N_17271,N_11303,N_13648);
nor U17272 (N_17272,N_10122,N_11117);
nand U17273 (N_17273,N_10658,N_14059);
xor U17274 (N_17274,N_14760,N_13366);
nand U17275 (N_17275,N_12592,N_14889);
xor U17276 (N_17276,N_14417,N_13124);
and U17277 (N_17277,N_12130,N_14098);
or U17278 (N_17278,N_10563,N_12131);
and U17279 (N_17279,N_11569,N_13031);
and U17280 (N_17280,N_14963,N_14938);
xor U17281 (N_17281,N_12472,N_10699);
nor U17282 (N_17282,N_14342,N_12573);
and U17283 (N_17283,N_13067,N_13998);
and U17284 (N_17284,N_13888,N_12965);
nand U17285 (N_17285,N_13838,N_12812);
and U17286 (N_17286,N_11286,N_12398);
nor U17287 (N_17287,N_13940,N_11015);
xor U17288 (N_17288,N_11098,N_10305);
xnor U17289 (N_17289,N_14096,N_10964);
xnor U17290 (N_17290,N_14356,N_13335);
xor U17291 (N_17291,N_13102,N_14549);
xor U17292 (N_17292,N_13559,N_14303);
or U17293 (N_17293,N_14368,N_10429);
or U17294 (N_17294,N_10394,N_11183);
and U17295 (N_17295,N_10326,N_11011);
or U17296 (N_17296,N_14072,N_10937);
xnor U17297 (N_17297,N_12978,N_14325);
nor U17298 (N_17298,N_14291,N_10020);
nand U17299 (N_17299,N_12196,N_12612);
xnor U17300 (N_17300,N_13146,N_11697);
and U17301 (N_17301,N_12464,N_11666);
nand U17302 (N_17302,N_14036,N_14398);
xor U17303 (N_17303,N_12681,N_12137);
nor U17304 (N_17304,N_13014,N_12353);
nor U17305 (N_17305,N_11226,N_12394);
nor U17306 (N_17306,N_13877,N_12186);
nand U17307 (N_17307,N_13398,N_12111);
xor U17308 (N_17308,N_12689,N_12552);
xnor U17309 (N_17309,N_12056,N_12076);
nor U17310 (N_17310,N_14997,N_10400);
nor U17311 (N_17311,N_12067,N_11282);
nor U17312 (N_17312,N_14622,N_13140);
and U17313 (N_17313,N_12279,N_14191);
and U17314 (N_17314,N_12841,N_12029);
nor U17315 (N_17315,N_13421,N_11560);
nor U17316 (N_17316,N_13810,N_12204);
or U17317 (N_17317,N_10276,N_12191);
nor U17318 (N_17318,N_14055,N_10753);
nor U17319 (N_17319,N_11378,N_13452);
and U17320 (N_17320,N_10443,N_11952);
and U17321 (N_17321,N_14287,N_10017);
or U17322 (N_17322,N_11326,N_12007);
nor U17323 (N_17323,N_13375,N_12686);
nor U17324 (N_17324,N_12913,N_12733);
nor U17325 (N_17325,N_14957,N_10684);
and U17326 (N_17326,N_14886,N_12755);
nor U17327 (N_17327,N_14713,N_12088);
xor U17328 (N_17328,N_13489,N_10836);
or U17329 (N_17329,N_11167,N_11122);
xnor U17330 (N_17330,N_11392,N_14908);
xnor U17331 (N_17331,N_10428,N_11570);
nor U17332 (N_17332,N_13642,N_12995);
nor U17333 (N_17333,N_11490,N_13458);
xnor U17334 (N_17334,N_14668,N_11214);
xnor U17335 (N_17335,N_11841,N_11219);
or U17336 (N_17336,N_13956,N_10987);
or U17337 (N_17337,N_13586,N_14725);
nand U17338 (N_17338,N_11331,N_10817);
and U17339 (N_17339,N_14319,N_11656);
nand U17340 (N_17340,N_14695,N_14795);
and U17341 (N_17341,N_14024,N_12760);
and U17342 (N_17342,N_10391,N_12919);
xnor U17343 (N_17343,N_14058,N_14670);
nand U17344 (N_17344,N_13144,N_11903);
xnor U17345 (N_17345,N_13300,N_14116);
and U17346 (N_17346,N_12735,N_12477);
nand U17347 (N_17347,N_12957,N_10951);
and U17348 (N_17348,N_14293,N_10232);
nor U17349 (N_17349,N_10721,N_10306);
or U17350 (N_17350,N_14609,N_11588);
and U17351 (N_17351,N_10374,N_14516);
xnor U17352 (N_17352,N_13850,N_13083);
nor U17353 (N_17353,N_10587,N_14971);
xnor U17354 (N_17354,N_14923,N_14374);
and U17355 (N_17355,N_11148,N_10036);
or U17356 (N_17356,N_10788,N_10159);
xnor U17357 (N_17357,N_10687,N_11420);
or U17358 (N_17358,N_12445,N_11801);
nand U17359 (N_17359,N_10933,N_13658);
nor U17360 (N_17360,N_12781,N_14952);
nand U17361 (N_17361,N_13309,N_14007);
or U17362 (N_17362,N_11825,N_14946);
xnor U17363 (N_17363,N_14909,N_11395);
nor U17364 (N_17364,N_14994,N_10844);
xnor U17365 (N_17365,N_10121,N_11900);
nor U17366 (N_17366,N_12551,N_13627);
or U17367 (N_17367,N_11093,N_10155);
nor U17368 (N_17368,N_12199,N_11022);
xnor U17369 (N_17369,N_14605,N_12023);
xnor U17370 (N_17370,N_14264,N_11733);
nor U17371 (N_17371,N_11111,N_12075);
nor U17372 (N_17372,N_10779,N_12773);
or U17373 (N_17373,N_13815,N_10153);
nand U17374 (N_17374,N_14371,N_12939);
or U17375 (N_17375,N_10445,N_10997);
nor U17376 (N_17376,N_14115,N_11033);
and U17377 (N_17377,N_11278,N_13076);
nor U17378 (N_17378,N_12455,N_10505);
nand U17379 (N_17379,N_14220,N_10057);
xnor U17380 (N_17380,N_14379,N_13404);
and U17381 (N_17381,N_14628,N_13159);
xnor U17382 (N_17382,N_12282,N_13976);
or U17383 (N_17383,N_12415,N_10342);
and U17384 (N_17384,N_11746,N_14464);
nor U17385 (N_17385,N_13625,N_10651);
xnor U17386 (N_17386,N_11191,N_14906);
or U17387 (N_17387,N_10451,N_14088);
or U17388 (N_17388,N_12184,N_10918);
nor U17389 (N_17389,N_13505,N_12185);
or U17390 (N_17390,N_11837,N_13897);
nand U17391 (N_17391,N_13188,N_10373);
xnor U17392 (N_17392,N_10440,N_10961);
nand U17393 (N_17393,N_14972,N_10705);
or U17394 (N_17394,N_14989,N_14380);
or U17395 (N_17395,N_10079,N_14219);
nor U17396 (N_17396,N_14084,N_10325);
nor U17397 (N_17397,N_14806,N_10499);
or U17398 (N_17398,N_13308,N_12718);
nand U17399 (N_17399,N_14127,N_10673);
nand U17400 (N_17400,N_11207,N_12360);
xor U17401 (N_17401,N_12054,N_14532);
nand U17402 (N_17402,N_12195,N_13171);
and U17403 (N_17403,N_12949,N_13333);
and U17404 (N_17404,N_14580,N_12133);
or U17405 (N_17405,N_11762,N_14427);
xor U17406 (N_17406,N_10504,N_10092);
and U17407 (N_17407,N_11584,N_12400);
nor U17408 (N_17408,N_11419,N_10389);
nor U17409 (N_17409,N_12975,N_12043);
or U17410 (N_17410,N_10280,N_10413);
and U17411 (N_17411,N_11650,N_12816);
or U17412 (N_17412,N_10808,N_10359);
xnor U17413 (N_17413,N_13816,N_13646);
nand U17414 (N_17414,N_14749,N_12844);
and U17415 (N_17415,N_12821,N_14008);
nor U17416 (N_17416,N_11228,N_11509);
or U17417 (N_17417,N_11972,N_10127);
xnor U17418 (N_17418,N_10126,N_12176);
or U17419 (N_17419,N_12292,N_12038);
nor U17420 (N_17420,N_13984,N_10547);
xor U17421 (N_17421,N_11965,N_12316);
or U17422 (N_17422,N_13510,N_13323);
nor U17423 (N_17423,N_14095,N_11155);
nand U17424 (N_17424,N_12321,N_14104);
or U17425 (N_17425,N_11731,N_10245);
nand U17426 (N_17426,N_13043,N_10766);
nor U17427 (N_17427,N_14075,N_11089);
nand U17428 (N_17428,N_11079,N_14140);
and U17429 (N_17429,N_12041,N_12695);
nand U17430 (N_17430,N_13106,N_10761);
and U17431 (N_17431,N_12277,N_10799);
nand U17432 (N_17432,N_12175,N_12637);
xnor U17433 (N_17433,N_13501,N_10666);
or U17434 (N_17434,N_10187,N_10065);
or U17435 (N_17435,N_14613,N_14097);
nor U17436 (N_17436,N_14553,N_11414);
and U17437 (N_17437,N_14335,N_12391);
xnor U17438 (N_17438,N_13359,N_12459);
nand U17439 (N_17439,N_13992,N_13771);
or U17440 (N_17440,N_10387,N_13832);
or U17441 (N_17441,N_13468,N_13514);
nor U17442 (N_17442,N_14155,N_11316);
nor U17443 (N_17443,N_11150,N_13979);
and U17444 (N_17444,N_12288,N_12648);
nor U17445 (N_17445,N_12334,N_13580);
and U17446 (N_17446,N_10882,N_14326);
nand U17447 (N_17447,N_10192,N_13735);
xnor U17448 (N_17448,N_10349,N_11388);
nand U17449 (N_17449,N_14658,N_11261);
or U17450 (N_17450,N_11321,N_13651);
or U17451 (N_17451,N_12402,N_11894);
nor U17452 (N_17452,N_11673,N_10790);
xor U17453 (N_17453,N_13077,N_12824);
xnor U17454 (N_17454,N_12529,N_11131);
nor U17455 (N_17455,N_12916,N_10053);
and U17456 (N_17456,N_12940,N_12520);
nor U17457 (N_17457,N_10794,N_10220);
nor U17458 (N_17458,N_13536,N_12417);
nor U17459 (N_17459,N_11295,N_11546);
or U17460 (N_17460,N_14915,N_14692);
xnor U17461 (N_17461,N_12717,N_14239);
nand U17462 (N_17462,N_14422,N_11405);
or U17463 (N_17463,N_12327,N_11097);
nor U17464 (N_17464,N_14210,N_11725);
and U17465 (N_17465,N_12774,N_12635);
or U17466 (N_17466,N_10441,N_13784);
or U17467 (N_17467,N_11154,N_11706);
nand U17468 (N_17468,N_11456,N_10821);
xnor U17469 (N_17469,N_11852,N_14212);
nand U17470 (N_17470,N_11514,N_10777);
or U17471 (N_17471,N_13764,N_12274);
nand U17472 (N_17472,N_14596,N_10998);
nor U17473 (N_17473,N_13537,N_14403);
nor U17474 (N_17474,N_12252,N_12095);
nand U17475 (N_17475,N_14732,N_13002);
and U17476 (N_17476,N_14472,N_12497);
xnor U17477 (N_17477,N_10626,N_14525);
and U17478 (N_17478,N_13781,N_12851);
or U17479 (N_17479,N_14870,N_12515);
or U17480 (N_17480,N_12590,N_13223);
nor U17481 (N_17481,N_10528,N_12541);
nand U17482 (N_17482,N_10988,N_10439);
xnor U17483 (N_17483,N_12435,N_12887);
xor U17484 (N_17484,N_13008,N_13190);
xor U17485 (N_17485,N_10281,N_10251);
nor U17486 (N_17486,N_11193,N_14967);
xor U17487 (N_17487,N_14217,N_10177);
xnor U17488 (N_17488,N_12937,N_12941);
nand U17489 (N_17489,N_10521,N_11664);
or U17490 (N_17490,N_10650,N_10592);
xnor U17491 (N_17491,N_13184,N_13552);
xor U17492 (N_17492,N_12428,N_10807);
or U17493 (N_17493,N_10458,N_12628);
xnor U17494 (N_17494,N_11919,N_11838);
nor U17495 (N_17495,N_11272,N_14146);
xor U17496 (N_17496,N_14382,N_10075);
nand U17497 (N_17497,N_14015,N_13934);
xor U17498 (N_17498,N_12739,N_12214);
or U17499 (N_17499,N_11141,N_12496);
xor U17500 (N_17500,N_10113,N_14698);
or U17501 (N_17501,N_11325,N_14482);
nand U17502 (N_17502,N_13723,N_12199);
nand U17503 (N_17503,N_13471,N_12165);
or U17504 (N_17504,N_13349,N_10502);
and U17505 (N_17505,N_12880,N_14884);
nand U17506 (N_17506,N_12598,N_10072);
and U17507 (N_17507,N_10797,N_13938);
and U17508 (N_17508,N_11636,N_11949);
nand U17509 (N_17509,N_14407,N_12491);
nor U17510 (N_17510,N_14083,N_12130);
nand U17511 (N_17511,N_11970,N_10941);
or U17512 (N_17512,N_11893,N_10767);
xor U17513 (N_17513,N_10023,N_14655);
nor U17514 (N_17514,N_12570,N_12309);
nand U17515 (N_17515,N_12805,N_13766);
and U17516 (N_17516,N_13058,N_10945);
or U17517 (N_17517,N_14862,N_13713);
nor U17518 (N_17518,N_11750,N_11670);
nor U17519 (N_17519,N_10683,N_10178);
and U17520 (N_17520,N_11490,N_12584);
nand U17521 (N_17521,N_13224,N_12898);
and U17522 (N_17522,N_12750,N_10456);
xor U17523 (N_17523,N_12443,N_10455);
and U17524 (N_17524,N_11610,N_10000);
xnor U17525 (N_17525,N_14145,N_12352);
or U17526 (N_17526,N_14434,N_12455);
nand U17527 (N_17527,N_12759,N_10935);
or U17528 (N_17528,N_11175,N_10314);
nand U17529 (N_17529,N_13143,N_10770);
xnor U17530 (N_17530,N_12110,N_13848);
nor U17531 (N_17531,N_12942,N_14572);
nor U17532 (N_17532,N_13719,N_11861);
nor U17533 (N_17533,N_11914,N_12105);
or U17534 (N_17534,N_14170,N_10715);
nand U17535 (N_17535,N_13898,N_13870);
nand U17536 (N_17536,N_14905,N_14150);
nor U17537 (N_17537,N_14203,N_14194);
or U17538 (N_17538,N_11794,N_12148);
or U17539 (N_17539,N_11194,N_10964);
nand U17540 (N_17540,N_11919,N_13708);
or U17541 (N_17541,N_13526,N_12488);
xnor U17542 (N_17542,N_12393,N_11321);
or U17543 (N_17543,N_13118,N_11634);
nor U17544 (N_17544,N_12718,N_14844);
or U17545 (N_17545,N_10385,N_11087);
xor U17546 (N_17546,N_10811,N_14936);
or U17547 (N_17547,N_14136,N_12173);
xnor U17548 (N_17548,N_12842,N_14379);
nor U17549 (N_17549,N_10755,N_13811);
nor U17550 (N_17550,N_11837,N_11734);
nand U17551 (N_17551,N_14601,N_12926);
nor U17552 (N_17552,N_10672,N_11227);
and U17553 (N_17553,N_10463,N_10211);
nand U17554 (N_17554,N_12178,N_12664);
and U17555 (N_17555,N_14965,N_10663);
nor U17556 (N_17556,N_13245,N_12459);
and U17557 (N_17557,N_13525,N_13305);
xor U17558 (N_17558,N_11562,N_11482);
nor U17559 (N_17559,N_14315,N_14229);
or U17560 (N_17560,N_10745,N_12580);
xor U17561 (N_17561,N_11325,N_11038);
or U17562 (N_17562,N_11935,N_11152);
and U17563 (N_17563,N_12249,N_10067);
and U17564 (N_17564,N_11196,N_13669);
nand U17565 (N_17565,N_13519,N_11875);
and U17566 (N_17566,N_11348,N_11263);
xnor U17567 (N_17567,N_11792,N_11972);
nor U17568 (N_17568,N_10433,N_14103);
xor U17569 (N_17569,N_11511,N_14243);
or U17570 (N_17570,N_12756,N_10377);
or U17571 (N_17571,N_12144,N_13894);
and U17572 (N_17572,N_14276,N_13834);
nor U17573 (N_17573,N_12198,N_12359);
nor U17574 (N_17574,N_10007,N_14676);
nand U17575 (N_17575,N_10667,N_11271);
nand U17576 (N_17576,N_14041,N_10331);
nor U17577 (N_17577,N_10484,N_12217);
or U17578 (N_17578,N_11845,N_12206);
or U17579 (N_17579,N_12992,N_10184);
xor U17580 (N_17580,N_11453,N_10365);
nand U17581 (N_17581,N_11843,N_14654);
nand U17582 (N_17582,N_13810,N_13680);
nor U17583 (N_17583,N_13529,N_11666);
nand U17584 (N_17584,N_12040,N_12010);
or U17585 (N_17585,N_14756,N_13102);
nor U17586 (N_17586,N_12309,N_13736);
or U17587 (N_17587,N_13234,N_10562);
or U17588 (N_17588,N_12788,N_12442);
xor U17589 (N_17589,N_12970,N_12074);
and U17590 (N_17590,N_12233,N_13411);
and U17591 (N_17591,N_10173,N_13829);
xnor U17592 (N_17592,N_11513,N_10447);
nand U17593 (N_17593,N_11856,N_11260);
nor U17594 (N_17594,N_10282,N_14973);
nand U17595 (N_17595,N_12431,N_11761);
nor U17596 (N_17596,N_10397,N_14172);
nand U17597 (N_17597,N_13461,N_13704);
nand U17598 (N_17598,N_12045,N_12153);
nand U17599 (N_17599,N_10443,N_10101);
nor U17600 (N_17600,N_10323,N_12173);
or U17601 (N_17601,N_13556,N_11810);
and U17602 (N_17602,N_10342,N_14101);
or U17603 (N_17603,N_13086,N_12775);
or U17604 (N_17604,N_12619,N_12483);
or U17605 (N_17605,N_14095,N_10340);
or U17606 (N_17606,N_11225,N_13894);
and U17607 (N_17607,N_10486,N_10086);
nor U17608 (N_17608,N_10835,N_12421);
xnor U17609 (N_17609,N_10058,N_10253);
and U17610 (N_17610,N_13871,N_13015);
nor U17611 (N_17611,N_11733,N_14300);
nand U17612 (N_17612,N_10443,N_11323);
xnor U17613 (N_17613,N_13391,N_12419);
and U17614 (N_17614,N_12848,N_10210);
xnor U17615 (N_17615,N_14934,N_13547);
or U17616 (N_17616,N_13803,N_11438);
xor U17617 (N_17617,N_12251,N_12226);
nor U17618 (N_17618,N_14765,N_12974);
nand U17619 (N_17619,N_14455,N_11972);
or U17620 (N_17620,N_10851,N_13606);
and U17621 (N_17621,N_13363,N_11456);
nor U17622 (N_17622,N_13363,N_11866);
nor U17623 (N_17623,N_12175,N_10629);
and U17624 (N_17624,N_11682,N_13236);
nand U17625 (N_17625,N_12462,N_14069);
or U17626 (N_17626,N_14825,N_11000);
or U17627 (N_17627,N_13447,N_11259);
nand U17628 (N_17628,N_10202,N_12998);
nand U17629 (N_17629,N_12464,N_12539);
or U17630 (N_17630,N_11242,N_14368);
and U17631 (N_17631,N_13980,N_12548);
or U17632 (N_17632,N_13631,N_14511);
nand U17633 (N_17633,N_14270,N_11438);
nand U17634 (N_17634,N_11522,N_11688);
nand U17635 (N_17635,N_13732,N_10739);
or U17636 (N_17636,N_10811,N_14439);
and U17637 (N_17637,N_12745,N_14607);
and U17638 (N_17638,N_14448,N_14136);
nand U17639 (N_17639,N_10553,N_13340);
and U17640 (N_17640,N_11903,N_13469);
nand U17641 (N_17641,N_11385,N_11649);
or U17642 (N_17642,N_14622,N_13962);
and U17643 (N_17643,N_12653,N_14715);
and U17644 (N_17644,N_11460,N_12471);
xnor U17645 (N_17645,N_10149,N_14288);
or U17646 (N_17646,N_10497,N_14775);
xnor U17647 (N_17647,N_10771,N_10612);
nand U17648 (N_17648,N_14315,N_10741);
nand U17649 (N_17649,N_10880,N_14104);
nor U17650 (N_17650,N_13532,N_13097);
or U17651 (N_17651,N_11360,N_11489);
nand U17652 (N_17652,N_12353,N_11093);
xor U17653 (N_17653,N_11161,N_12220);
and U17654 (N_17654,N_12353,N_13291);
nand U17655 (N_17655,N_10324,N_12586);
or U17656 (N_17656,N_13305,N_10670);
xnor U17657 (N_17657,N_12541,N_10661);
nand U17658 (N_17658,N_11271,N_14673);
nor U17659 (N_17659,N_13603,N_14679);
xor U17660 (N_17660,N_12285,N_14387);
or U17661 (N_17661,N_11368,N_13171);
nand U17662 (N_17662,N_10577,N_12290);
or U17663 (N_17663,N_13362,N_10495);
or U17664 (N_17664,N_14681,N_11400);
xor U17665 (N_17665,N_14838,N_13892);
or U17666 (N_17666,N_14100,N_11105);
xor U17667 (N_17667,N_11204,N_11000);
nor U17668 (N_17668,N_11420,N_11556);
and U17669 (N_17669,N_12552,N_11480);
nor U17670 (N_17670,N_10673,N_12320);
nand U17671 (N_17671,N_13722,N_11672);
nor U17672 (N_17672,N_10082,N_14158);
and U17673 (N_17673,N_11990,N_10228);
nor U17674 (N_17674,N_14962,N_12144);
nor U17675 (N_17675,N_12602,N_12283);
xnor U17676 (N_17676,N_10154,N_13591);
nand U17677 (N_17677,N_14447,N_13025);
nor U17678 (N_17678,N_14023,N_14536);
and U17679 (N_17679,N_11601,N_14008);
nor U17680 (N_17680,N_12680,N_14203);
or U17681 (N_17681,N_12193,N_13172);
nor U17682 (N_17682,N_14216,N_10244);
nor U17683 (N_17683,N_11298,N_11450);
nor U17684 (N_17684,N_10539,N_10426);
xnor U17685 (N_17685,N_12247,N_14221);
or U17686 (N_17686,N_12975,N_11569);
and U17687 (N_17687,N_10715,N_13830);
nor U17688 (N_17688,N_10674,N_14723);
nor U17689 (N_17689,N_10271,N_10320);
nand U17690 (N_17690,N_10335,N_10735);
xnor U17691 (N_17691,N_14598,N_14824);
xor U17692 (N_17692,N_12724,N_14584);
nor U17693 (N_17693,N_14288,N_12349);
nand U17694 (N_17694,N_11907,N_14838);
or U17695 (N_17695,N_14799,N_10591);
and U17696 (N_17696,N_10469,N_14216);
nor U17697 (N_17697,N_11496,N_14926);
nor U17698 (N_17698,N_14892,N_12702);
nand U17699 (N_17699,N_10622,N_12784);
nor U17700 (N_17700,N_11463,N_12168);
xor U17701 (N_17701,N_11765,N_12627);
xor U17702 (N_17702,N_11474,N_11793);
and U17703 (N_17703,N_14428,N_11844);
and U17704 (N_17704,N_12412,N_11054);
nand U17705 (N_17705,N_10677,N_10922);
or U17706 (N_17706,N_10222,N_11233);
and U17707 (N_17707,N_11455,N_14691);
nand U17708 (N_17708,N_13110,N_12816);
or U17709 (N_17709,N_12510,N_14556);
or U17710 (N_17710,N_13251,N_12703);
or U17711 (N_17711,N_13440,N_14562);
nor U17712 (N_17712,N_12415,N_11236);
nand U17713 (N_17713,N_12601,N_12294);
or U17714 (N_17714,N_13825,N_11576);
xor U17715 (N_17715,N_14508,N_14365);
xor U17716 (N_17716,N_10981,N_13129);
nor U17717 (N_17717,N_12097,N_13005);
nor U17718 (N_17718,N_11538,N_12812);
or U17719 (N_17719,N_11847,N_14446);
or U17720 (N_17720,N_13825,N_10451);
nand U17721 (N_17721,N_10562,N_13476);
and U17722 (N_17722,N_12372,N_12483);
or U17723 (N_17723,N_14227,N_14071);
nor U17724 (N_17724,N_13421,N_11179);
nand U17725 (N_17725,N_12684,N_10939);
xnor U17726 (N_17726,N_12578,N_12476);
xor U17727 (N_17727,N_12209,N_11823);
or U17728 (N_17728,N_10228,N_10239);
and U17729 (N_17729,N_11086,N_13828);
and U17730 (N_17730,N_14633,N_11807);
and U17731 (N_17731,N_10450,N_13538);
nor U17732 (N_17732,N_10837,N_11909);
nor U17733 (N_17733,N_11253,N_13782);
nor U17734 (N_17734,N_10466,N_14046);
nand U17735 (N_17735,N_12438,N_14642);
and U17736 (N_17736,N_14397,N_12634);
xnor U17737 (N_17737,N_12263,N_14322);
or U17738 (N_17738,N_13865,N_13948);
or U17739 (N_17739,N_12922,N_13549);
xor U17740 (N_17740,N_14561,N_11254);
nand U17741 (N_17741,N_10142,N_14402);
nor U17742 (N_17742,N_10963,N_13591);
nand U17743 (N_17743,N_10961,N_14554);
xor U17744 (N_17744,N_10146,N_10091);
xnor U17745 (N_17745,N_10053,N_11177);
xnor U17746 (N_17746,N_12249,N_13559);
nor U17747 (N_17747,N_14666,N_14712);
xnor U17748 (N_17748,N_14238,N_12086);
xor U17749 (N_17749,N_12149,N_13391);
and U17750 (N_17750,N_11036,N_12653);
nand U17751 (N_17751,N_14734,N_12746);
nor U17752 (N_17752,N_13622,N_13499);
nor U17753 (N_17753,N_13041,N_13184);
nand U17754 (N_17754,N_14899,N_12053);
or U17755 (N_17755,N_11976,N_14821);
xor U17756 (N_17756,N_11762,N_10629);
or U17757 (N_17757,N_12020,N_11096);
xnor U17758 (N_17758,N_11044,N_14617);
and U17759 (N_17759,N_13880,N_14453);
xnor U17760 (N_17760,N_14597,N_10324);
or U17761 (N_17761,N_13054,N_14097);
nand U17762 (N_17762,N_14290,N_13772);
or U17763 (N_17763,N_11464,N_13345);
and U17764 (N_17764,N_13150,N_12311);
and U17765 (N_17765,N_11812,N_12280);
nand U17766 (N_17766,N_11182,N_13426);
and U17767 (N_17767,N_14118,N_10151);
or U17768 (N_17768,N_12981,N_14100);
or U17769 (N_17769,N_13475,N_11633);
xnor U17770 (N_17770,N_14177,N_10913);
nand U17771 (N_17771,N_12553,N_10484);
nand U17772 (N_17772,N_12177,N_13737);
xor U17773 (N_17773,N_14543,N_12967);
and U17774 (N_17774,N_11869,N_12621);
nor U17775 (N_17775,N_12997,N_12187);
xnor U17776 (N_17776,N_11515,N_12503);
nand U17777 (N_17777,N_14790,N_14878);
and U17778 (N_17778,N_14523,N_10859);
and U17779 (N_17779,N_11387,N_10257);
and U17780 (N_17780,N_12197,N_10284);
xnor U17781 (N_17781,N_14233,N_13762);
or U17782 (N_17782,N_12723,N_14527);
xor U17783 (N_17783,N_11863,N_10830);
nand U17784 (N_17784,N_14264,N_13168);
xor U17785 (N_17785,N_10147,N_14317);
nor U17786 (N_17786,N_10317,N_14965);
xor U17787 (N_17787,N_13743,N_14532);
or U17788 (N_17788,N_12147,N_10857);
nor U17789 (N_17789,N_11213,N_12292);
xnor U17790 (N_17790,N_13282,N_10572);
nor U17791 (N_17791,N_10999,N_10798);
nor U17792 (N_17792,N_10791,N_14427);
xor U17793 (N_17793,N_13428,N_14832);
nand U17794 (N_17794,N_14170,N_12971);
and U17795 (N_17795,N_13921,N_13361);
and U17796 (N_17796,N_11882,N_10430);
xor U17797 (N_17797,N_14302,N_12098);
nand U17798 (N_17798,N_12704,N_12822);
nor U17799 (N_17799,N_12309,N_14185);
nor U17800 (N_17800,N_13427,N_11489);
or U17801 (N_17801,N_14942,N_14536);
nand U17802 (N_17802,N_10525,N_14890);
xor U17803 (N_17803,N_14944,N_10848);
or U17804 (N_17804,N_11804,N_13301);
and U17805 (N_17805,N_11039,N_13062);
xnor U17806 (N_17806,N_12679,N_14601);
or U17807 (N_17807,N_13214,N_12398);
nand U17808 (N_17808,N_12683,N_13557);
nor U17809 (N_17809,N_13037,N_13640);
and U17810 (N_17810,N_11791,N_10637);
or U17811 (N_17811,N_14850,N_10935);
nor U17812 (N_17812,N_13025,N_12134);
xor U17813 (N_17813,N_13836,N_12254);
and U17814 (N_17814,N_11845,N_13452);
or U17815 (N_17815,N_12638,N_14992);
and U17816 (N_17816,N_11997,N_14255);
xnor U17817 (N_17817,N_11518,N_10990);
nand U17818 (N_17818,N_11027,N_11823);
nand U17819 (N_17819,N_12602,N_11185);
nor U17820 (N_17820,N_10500,N_12890);
xor U17821 (N_17821,N_10879,N_14002);
and U17822 (N_17822,N_12360,N_11228);
nor U17823 (N_17823,N_14394,N_14056);
or U17824 (N_17824,N_10501,N_12761);
and U17825 (N_17825,N_10709,N_11746);
xnor U17826 (N_17826,N_14819,N_14241);
and U17827 (N_17827,N_12420,N_13604);
nand U17828 (N_17828,N_10018,N_13092);
or U17829 (N_17829,N_14634,N_10963);
and U17830 (N_17830,N_13544,N_13327);
nor U17831 (N_17831,N_13716,N_10114);
nor U17832 (N_17832,N_10243,N_12311);
xnor U17833 (N_17833,N_14177,N_13815);
xor U17834 (N_17834,N_12041,N_12101);
and U17835 (N_17835,N_13313,N_12462);
xnor U17836 (N_17836,N_11155,N_13857);
nand U17837 (N_17837,N_10745,N_12102);
nand U17838 (N_17838,N_10187,N_10790);
xor U17839 (N_17839,N_14070,N_13100);
xnor U17840 (N_17840,N_11300,N_10426);
xor U17841 (N_17841,N_10520,N_12160);
or U17842 (N_17842,N_11883,N_11954);
xnor U17843 (N_17843,N_13975,N_11700);
nand U17844 (N_17844,N_10633,N_10511);
or U17845 (N_17845,N_11006,N_11307);
or U17846 (N_17846,N_10571,N_10205);
nor U17847 (N_17847,N_12913,N_11915);
nor U17848 (N_17848,N_12352,N_11333);
and U17849 (N_17849,N_11282,N_13109);
nor U17850 (N_17850,N_12153,N_11881);
xor U17851 (N_17851,N_14791,N_10838);
and U17852 (N_17852,N_10279,N_10004);
or U17853 (N_17853,N_14688,N_10066);
nand U17854 (N_17854,N_13156,N_13255);
and U17855 (N_17855,N_10464,N_14597);
xnor U17856 (N_17856,N_14661,N_13817);
or U17857 (N_17857,N_10900,N_13805);
or U17858 (N_17858,N_11770,N_10961);
xnor U17859 (N_17859,N_14752,N_11324);
nor U17860 (N_17860,N_10779,N_12914);
xor U17861 (N_17861,N_14533,N_12266);
and U17862 (N_17862,N_10412,N_13302);
nor U17863 (N_17863,N_10745,N_14717);
and U17864 (N_17864,N_11046,N_13683);
or U17865 (N_17865,N_12245,N_11077);
xnor U17866 (N_17866,N_10025,N_10982);
xnor U17867 (N_17867,N_12979,N_10346);
nand U17868 (N_17868,N_11999,N_12541);
xor U17869 (N_17869,N_14855,N_11084);
and U17870 (N_17870,N_12201,N_13233);
and U17871 (N_17871,N_13611,N_11796);
nor U17872 (N_17872,N_12764,N_12439);
and U17873 (N_17873,N_11269,N_11515);
nand U17874 (N_17874,N_12655,N_12659);
xor U17875 (N_17875,N_12355,N_10585);
and U17876 (N_17876,N_14814,N_13896);
nand U17877 (N_17877,N_14703,N_12374);
nand U17878 (N_17878,N_13271,N_12475);
nand U17879 (N_17879,N_13374,N_12116);
nor U17880 (N_17880,N_11997,N_10828);
and U17881 (N_17881,N_12358,N_12361);
nor U17882 (N_17882,N_10110,N_11300);
and U17883 (N_17883,N_11236,N_12980);
nor U17884 (N_17884,N_14939,N_14017);
nor U17885 (N_17885,N_13014,N_12061);
and U17886 (N_17886,N_12708,N_11738);
xnor U17887 (N_17887,N_12637,N_11939);
or U17888 (N_17888,N_11739,N_10622);
xnor U17889 (N_17889,N_13723,N_14141);
nand U17890 (N_17890,N_11878,N_13410);
or U17891 (N_17891,N_13018,N_11300);
and U17892 (N_17892,N_14565,N_12145);
nand U17893 (N_17893,N_12710,N_11635);
and U17894 (N_17894,N_11619,N_14940);
nand U17895 (N_17895,N_11878,N_11799);
or U17896 (N_17896,N_12238,N_11622);
or U17897 (N_17897,N_10633,N_14566);
and U17898 (N_17898,N_10386,N_11245);
nand U17899 (N_17899,N_10099,N_14080);
or U17900 (N_17900,N_11104,N_14190);
xor U17901 (N_17901,N_13542,N_12135);
or U17902 (N_17902,N_14591,N_10387);
nor U17903 (N_17903,N_10751,N_14018);
nor U17904 (N_17904,N_13329,N_10957);
or U17905 (N_17905,N_12880,N_14166);
xnor U17906 (N_17906,N_14593,N_12179);
nor U17907 (N_17907,N_14588,N_10972);
nand U17908 (N_17908,N_11783,N_11190);
and U17909 (N_17909,N_12448,N_12284);
nor U17910 (N_17910,N_13138,N_14869);
and U17911 (N_17911,N_14818,N_10090);
nand U17912 (N_17912,N_11787,N_11062);
or U17913 (N_17913,N_14821,N_14219);
or U17914 (N_17914,N_14253,N_11298);
xnor U17915 (N_17915,N_12921,N_13906);
nand U17916 (N_17916,N_12873,N_11652);
nor U17917 (N_17917,N_14900,N_12907);
or U17918 (N_17918,N_13791,N_11861);
or U17919 (N_17919,N_12918,N_10449);
nand U17920 (N_17920,N_14198,N_12628);
nand U17921 (N_17921,N_12300,N_13047);
or U17922 (N_17922,N_10386,N_11671);
nor U17923 (N_17923,N_10626,N_13009);
and U17924 (N_17924,N_12455,N_13660);
nor U17925 (N_17925,N_12790,N_10836);
and U17926 (N_17926,N_13854,N_12023);
nor U17927 (N_17927,N_11165,N_13365);
nand U17928 (N_17928,N_14507,N_14547);
nor U17929 (N_17929,N_13889,N_10380);
or U17930 (N_17930,N_11373,N_14326);
and U17931 (N_17931,N_13823,N_13450);
or U17932 (N_17932,N_12560,N_14143);
nor U17933 (N_17933,N_12006,N_13176);
and U17934 (N_17934,N_12475,N_13373);
and U17935 (N_17935,N_14971,N_12583);
xnor U17936 (N_17936,N_11432,N_11993);
and U17937 (N_17937,N_10945,N_12040);
nand U17938 (N_17938,N_10738,N_14490);
nand U17939 (N_17939,N_10080,N_12382);
and U17940 (N_17940,N_12022,N_10118);
and U17941 (N_17941,N_12178,N_11414);
nor U17942 (N_17942,N_14441,N_14311);
and U17943 (N_17943,N_13451,N_11250);
nor U17944 (N_17944,N_12678,N_12788);
xnor U17945 (N_17945,N_13616,N_14795);
and U17946 (N_17946,N_13259,N_10601);
nor U17947 (N_17947,N_12672,N_14688);
and U17948 (N_17948,N_13401,N_11612);
xor U17949 (N_17949,N_12013,N_11102);
nand U17950 (N_17950,N_12271,N_11617);
xnor U17951 (N_17951,N_14153,N_13977);
xor U17952 (N_17952,N_12304,N_11325);
xor U17953 (N_17953,N_11136,N_13181);
xor U17954 (N_17954,N_11540,N_14907);
and U17955 (N_17955,N_10381,N_13146);
and U17956 (N_17956,N_13993,N_14508);
nor U17957 (N_17957,N_10876,N_12030);
xor U17958 (N_17958,N_11166,N_13029);
xnor U17959 (N_17959,N_12867,N_14274);
nand U17960 (N_17960,N_14751,N_12255);
or U17961 (N_17961,N_10850,N_10063);
nor U17962 (N_17962,N_13114,N_12854);
nor U17963 (N_17963,N_13127,N_12964);
nand U17964 (N_17964,N_14015,N_12155);
nor U17965 (N_17965,N_10243,N_12356);
nand U17966 (N_17966,N_13631,N_11786);
xnor U17967 (N_17967,N_12177,N_12106);
nor U17968 (N_17968,N_12725,N_10924);
or U17969 (N_17969,N_13412,N_14392);
and U17970 (N_17970,N_10289,N_11996);
nand U17971 (N_17971,N_11711,N_13405);
and U17972 (N_17972,N_12047,N_14222);
nand U17973 (N_17973,N_13376,N_10927);
or U17974 (N_17974,N_12176,N_12988);
nor U17975 (N_17975,N_12584,N_12331);
and U17976 (N_17976,N_10764,N_10282);
nor U17977 (N_17977,N_14109,N_11209);
nor U17978 (N_17978,N_13846,N_11501);
nand U17979 (N_17979,N_11774,N_12322);
and U17980 (N_17980,N_14391,N_12464);
and U17981 (N_17981,N_11551,N_12939);
nor U17982 (N_17982,N_11597,N_14196);
and U17983 (N_17983,N_14805,N_14368);
nor U17984 (N_17984,N_12481,N_14483);
and U17985 (N_17985,N_10677,N_11613);
nand U17986 (N_17986,N_13644,N_13618);
xnor U17987 (N_17987,N_11088,N_12616);
nor U17988 (N_17988,N_14321,N_12981);
xor U17989 (N_17989,N_10189,N_10146);
nor U17990 (N_17990,N_11250,N_12513);
or U17991 (N_17991,N_10686,N_10109);
xor U17992 (N_17992,N_12953,N_11360);
nand U17993 (N_17993,N_10885,N_11927);
or U17994 (N_17994,N_11521,N_14340);
or U17995 (N_17995,N_11741,N_10521);
nor U17996 (N_17996,N_11109,N_14310);
nor U17997 (N_17997,N_13130,N_11504);
and U17998 (N_17998,N_12900,N_11809);
nor U17999 (N_17999,N_10480,N_12560);
or U18000 (N_18000,N_13218,N_10969);
or U18001 (N_18001,N_10207,N_10859);
nand U18002 (N_18002,N_10055,N_13518);
and U18003 (N_18003,N_11111,N_12294);
nor U18004 (N_18004,N_14710,N_13810);
or U18005 (N_18005,N_10890,N_12021);
nor U18006 (N_18006,N_14142,N_10594);
nor U18007 (N_18007,N_12354,N_13207);
xor U18008 (N_18008,N_13591,N_11367);
xnor U18009 (N_18009,N_11820,N_10738);
nor U18010 (N_18010,N_10196,N_13619);
or U18011 (N_18011,N_13126,N_11649);
nand U18012 (N_18012,N_10378,N_10372);
nand U18013 (N_18013,N_12033,N_11434);
and U18014 (N_18014,N_10633,N_11093);
or U18015 (N_18015,N_12789,N_10586);
nor U18016 (N_18016,N_14417,N_12209);
nor U18017 (N_18017,N_14393,N_14795);
and U18018 (N_18018,N_12451,N_13938);
and U18019 (N_18019,N_10875,N_13453);
nand U18020 (N_18020,N_14511,N_13794);
nand U18021 (N_18021,N_11063,N_14247);
nor U18022 (N_18022,N_10696,N_10013);
and U18023 (N_18023,N_12479,N_10590);
and U18024 (N_18024,N_10397,N_10870);
and U18025 (N_18025,N_10958,N_12284);
nand U18026 (N_18026,N_11567,N_13474);
nand U18027 (N_18027,N_13936,N_14805);
nor U18028 (N_18028,N_13809,N_14232);
xnor U18029 (N_18029,N_14130,N_11505);
nor U18030 (N_18030,N_12163,N_12671);
or U18031 (N_18031,N_14769,N_11780);
xnor U18032 (N_18032,N_14762,N_11049);
nand U18033 (N_18033,N_11878,N_13631);
nand U18034 (N_18034,N_12962,N_12307);
xor U18035 (N_18035,N_11233,N_13522);
nor U18036 (N_18036,N_14838,N_12016);
or U18037 (N_18037,N_13165,N_11436);
and U18038 (N_18038,N_13597,N_14638);
and U18039 (N_18039,N_14912,N_14720);
and U18040 (N_18040,N_13721,N_13135);
nor U18041 (N_18041,N_10915,N_13192);
and U18042 (N_18042,N_13940,N_10044);
xor U18043 (N_18043,N_13073,N_11355);
nor U18044 (N_18044,N_10876,N_12334);
and U18045 (N_18045,N_11815,N_12346);
nand U18046 (N_18046,N_14746,N_11591);
nor U18047 (N_18047,N_10189,N_10550);
and U18048 (N_18048,N_14879,N_12047);
xnor U18049 (N_18049,N_13678,N_11629);
xor U18050 (N_18050,N_10547,N_12385);
xor U18051 (N_18051,N_14987,N_10174);
or U18052 (N_18052,N_14608,N_14636);
or U18053 (N_18053,N_11184,N_14451);
and U18054 (N_18054,N_11971,N_10008);
and U18055 (N_18055,N_10745,N_13653);
xor U18056 (N_18056,N_11816,N_13362);
and U18057 (N_18057,N_11811,N_13397);
nor U18058 (N_18058,N_11350,N_13051);
and U18059 (N_18059,N_10465,N_12875);
nand U18060 (N_18060,N_14925,N_14406);
nand U18061 (N_18061,N_10257,N_13147);
and U18062 (N_18062,N_11002,N_12868);
and U18063 (N_18063,N_14102,N_14267);
nand U18064 (N_18064,N_11419,N_14376);
or U18065 (N_18065,N_14845,N_10890);
xnor U18066 (N_18066,N_14060,N_12751);
xor U18067 (N_18067,N_12993,N_10939);
nand U18068 (N_18068,N_11871,N_12572);
xnor U18069 (N_18069,N_13598,N_11142);
or U18070 (N_18070,N_10224,N_13062);
nor U18071 (N_18071,N_10655,N_11784);
xnor U18072 (N_18072,N_13689,N_13100);
nand U18073 (N_18073,N_13349,N_11102);
and U18074 (N_18074,N_14145,N_10579);
or U18075 (N_18075,N_12869,N_10756);
xnor U18076 (N_18076,N_13013,N_10391);
xor U18077 (N_18077,N_12856,N_11622);
xnor U18078 (N_18078,N_11590,N_10728);
or U18079 (N_18079,N_12313,N_14702);
and U18080 (N_18080,N_13688,N_12030);
or U18081 (N_18081,N_13442,N_10653);
or U18082 (N_18082,N_10946,N_10373);
xor U18083 (N_18083,N_12941,N_12567);
and U18084 (N_18084,N_12336,N_14956);
nand U18085 (N_18085,N_13312,N_13597);
or U18086 (N_18086,N_14262,N_13045);
nand U18087 (N_18087,N_14440,N_14197);
or U18088 (N_18088,N_10271,N_10998);
xor U18089 (N_18089,N_13809,N_11641);
xor U18090 (N_18090,N_11534,N_12719);
xor U18091 (N_18091,N_14504,N_10577);
nand U18092 (N_18092,N_12007,N_12939);
nand U18093 (N_18093,N_11752,N_11499);
xnor U18094 (N_18094,N_14480,N_10862);
nand U18095 (N_18095,N_14758,N_13452);
nor U18096 (N_18096,N_14852,N_12738);
nor U18097 (N_18097,N_10815,N_12368);
nor U18098 (N_18098,N_12933,N_10267);
or U18099 (N_18099,N_11450,N_10864);
nand U18100 (N_18100,N_14064,N_13243);
or U18101 (N_18101,N_10147,N_10510);
nor U18102 (N_18102,N_13751,N_14295);
and U18103 (N_18103,N_13210,N_11605);
or U18104 (N_18104,N_14779,N_14888);
and U18105 (N_18105,N_11525,N_12093);
nand U18106 (N_18106,N_11476,N_12944);
or U18107 (N_18107,N_13103,N_11429);
nand U18108 (N_18108,N_11318,N_11130);
nor U18109 (N_18109,N_14145,N_14409);
and U18110 (N_18110,N_11060,N_11837);
or U18111 (N_18111,N_12006,N_12284);
xnor U18112 (N_18112,N_11821,N_10938);
and U18113 (N_18113,N_14416,N_12852);
nor U18114 (N_18114,N_13989,N_12664);
nand U18115 (N_18115,N_13927,N_10372);
nor U18116 (N_18116,N_13441,N_11562);
and U18117 (N_18117,N_13091,N_10190);
and U18118 (N_18118,N_11595,N_11662);
nand U18119 (N_18119,N_14336,N_13827);
nor U18120 (N_18120,N_10503,N_14685);
and U18121 (N_18121,N_12158,N_14005);
xor U18122 (N_18122,N_13885,N_13566);
or U18123 (N_18123,N_14504,N_11840);
and U18124 (N_18124,N_14079,N_11758);
xor U18125 (N_18125,N_13610,N_14584);
xnor U18126 (N_18126,N_10851,N_12446);
nor U18127 (N_18127,N_11752,N_14105);
or U18128 (N_18128,N_12271,N_11933);
and U18129 (N_18129,N_10253,N_11236);
xnor U18130 (N_18130,N_13664,N_14804);
nor U18131 (N_18131,N_14924,N_12495);
or U18132 (N_18132,N_12843,N_13227);
xor U18133 (N_18133,N_14895,N_11199);
xnor U18134 (N_18134,N_12683,N_13825);
or U18135 (N_18135,N_11756,N_10187);
and U18136 (N_18136,N_11717,N_10955);
or U18137 (N_18137,N_14957,N_14009);
nand U18138 (N_18138,N_10540,N_13354);
nand U18139 (N_18139,N_10730,N_14417);
xor U18140 (N_18140,N_12662,N_14202);
nand U18141 (N_18141,N_10503,N_13293);
nand U18142 (N_18142,N_13005,N_12086);
and U18143 (N_18143,N_14579,N_13630);
xor U18144 (N_18144,N_12972,N_14201);
xnor U18145 (N_18145,N_12023,N_11479);
nand U18146 (N_18146,N_14014,N_11544);
xnor U18147 (N_18147,N_12493,N_14786);
or U18148 (N_18148,N_10940,N_13361);
xnor U18149 (N_18149,N_11019,N_13914);
nor U18150 (N_18150,N_13952,N_10919);
xor U18151 (N_18151,N_12200,N_13576);
xor U18152 (N_18152,N_10956,N_10283);
nand U18153 (N_18153,N_10039,N_13928);
nor U18154 (N_18154,N_11826,N_12880);
and U18155 (N_18155,N_13514,N_14858);
and U18156 (N_18156,N_14776,N_13903);
nand U18157 (N_18157,N_11473,N_13282);
nand U18158 (N_18158,N_12362,N_13848);
and U18159 (N_18159,N_12413,N_13892);
nor U18160 (N_18160,N_14105,N_14618);
nand U18161 (N_18161,N_13730,N_11196);
nor U18162 (N_18162,N_11189,N_12275);
nand U18163 (N_18163,N_14725,N_13825);
nand U18164 (N_18164,N_11459,N_13321);
xnor U18165 (N_18165,N_13460,N_14218);
nor U18166 (N_18166,N_14220,N_14680);
or U18167 (N_18167,N_14696,N_11414);
nand U18168 (N_18168,N_13242,N_10719);
nor U18169 (N_18169,N_13770,N_13427);
nand U18170 (N_18170,N_11978,N_14994);
xor U18171 (N_18171,N_14877,N_11567);
and U18172 (N_18172,N_11234,N_11987);
nor U18173 (N_18173,N_11171,N_11640);
nor U18174 (N_18174,N_10824,N_13049);
xor U18175 (N_18175,N_11363,N_12288);
xor U18176 (N_18176,N_13896,N_10850);
nor U18177 (N_18177,N_10213,N_13416);
xor U18178 (N_18178,N_13984,N_13692);
xnor U18179 (N_18179,N_10878,N_11250);
or U18180 (N_18180,N_10609,N_14943);
nand U18181 (N_18181,N_11946,N_10980);
xor U18182 (N_18182,N_11077,N_11421);
nor U18183 (N_18183,N_10268,N_12002);
nand U18184 (N_18184,N_14381,N_12748);
nor U18185 (N_18185,N_13185,N_12808);
or U18186 (N_18186,N_12063,N_14772);
or U18187 (N_18187,N_10831,N_10975);
nand U18188 (N_18188,N_14255,N_13036);
nor U18189 (N_18189,N_10669,N_13904);
or U18190 (N_18190,N_12051,N_14749);
nand U18191 (N_18191,N_12264,N_12499);
nor U18192 (N_18192,N_10957,N_14506);
nand U18193 (N_18193,N_14213,N_14975);
nand U18194 (N_18194,N_13194,N_13495);
nor U18195 (N_18195,N_11651,N_10924);
nand U18196 (N_18196,N_10740,N_13011);
xor U18197 (N_18197,N_13196,N_10744);
or U18198 (N_18198,N_12526,N_10566);
or U18199 (N_18199,N_10040,N_13287);
and U18200 (N_18200,N_11981,N_10691);
and U18201 (N_18201,N_11333,N_12799);
and U18202 (N_18202,N_13173,N_10989);
xnor U18203 (N_18203,N_11889,N_10812);
or U18204 (N_18204,N_13068,N_10610);
and U18205 (N_18205,N_13843,N_13915);
xnor U18206 (N_18206,N_14145,N_12606);
nor U18207 (N_18207,N_10689,N_14506);
nor U18208 (N_18208,N_10670,N_13491);
nor U18209 (N_18209,N_12890,N_14741);
xnor U18210 (N_18210,N_12126,N_12306);
and U18211 (N_18211,N_10049,N_11633);
nor U18212 (N_18212,N_10375,N_11929);
and U18213 (N_18213,N_13702,N_14329);
nand U18214 (N_18214,N_13092,N_13679);
nand U18215 (N_18215,N_10118,N_10020);
xor U18216 (N_18216,N_10260,N_10277);
nor U18217 (N_18217,N_10198,N_13557);
nand U18218 (N_18218,N_13528,N_14619);
and U18219 (N_18219,N_10933,N_13299);
and U18220 (N_18220,N_10089,N_14613);
nand U18221 (N_18221,N_14157,N_12315);
nor U18222 (N_18222,N_14140,N_12137);
nor U18223 (N_18223,N_11313,N_10508);
and U18224 (N_18224,N_10630,N_14850);
nand U18225 (N_18225,N_10143,N_11482);
nand U18226 (N_18226,N_14489,N_11428);
xnor U18227 (N_18227,N_14024,N_10931);
nor U18228 (N_18228,N_14858,N_12175);
and U18229 (N_18229,N_11891,N_13148);
xnor U18230 (N_18230,N_12967,N_13177);
and U18231 (N_18231,N_11780,N_12188);
and U18232 (N_18232,N_12447,N_12769);
and U18233 (N_18233,N_14210,N_12833);
and U18234 (N_18234,N_11577,N_13047);
xor U18235 (N_18235,N_12959,N_10325);
nor U18236 (N_18236,N_13671,N_14774);
nor U18237 (N_18237,N_13876,N_12290);
nor U18238 (N_18238,N_10672,N_13380);
xnor U18239 (N_18239,N_12272,N_14993);
nor U18240 (N_18240,N_13900,N_12133);
and U18241 (N_18241,N_12603,N_10584);
nand U18242 (N_18242,N_10654,N_13760);
nor U18243 (N_18243,N_13952,N_10507);
or U18244 (N_18244,N_14134,N_14230);
or U18245 (N_18245,N_11928,N_12237);
or U18246 (N_18246,N_12830,N_11545);
nand U18247 (N_18247,N_11332,N_14639);
xnor U18248 (N_18248,N_11215,N_12041);
nand U18249 (N_18249,N_14820,N_14379);
nor U18250 (N_18250,N_14116,N_10034);
nor U18251 (N_18251,N_10280,N_14230);
and U18252 (N_18252,N_14543,N_14869);
nor U18253 (N_18253,N_10427,N_11886);
or U18254 (N_18254,N_13329,N_10302);
nand U18255 (N_18255,N_13735,N_10699);
or U18256 (N_18256,N_13279,N_12939);
or U18257 (N_18257,N_12096,N_13318);
xor U18258 (N_18258,N_13659,N_12119);
nor U18259 (N_18259,N_14066,N_13121);
or U18260 (N_18260,N_12662,N_10449);
xnor U18261 (N_18261,N_12355,N_14041);
nor U18262 (N_18262,N_11466,N_13954);
or U18263 (N_18263,N_14249,N_14107);
or U18264 (N_18264,N_11460,N_11877);
nand U18265 (N_18265,N_10262,N_13515);
nor U18266 (N_18266,N_13332,N_12324);
and U18267 (N_18267,N_11548,N_13155);
nor U18268 (N_18268,N_13030,N_12314);
xnor U18269 (N_18269,N_11903,N_13263);
xor U18270 (N_18270,N_14937,N_10371);
xnor U18271 (N_18271,N_14658,N_10239);
and U18272 (N_18272,N_11901,N_10530);
and U18273 (N_18273,N_13721,N_10948);
or U18274 (N_18274,N_10371,N_14281);
and U18275 (N_18275,N_13974,N_12728);
or U18276 (N_18276,N_14756,N_14173);
nand U18277 (N_18277,N_12753,N_10099);
nor U18278 (N_18278,N_10013,N_10235);
xnor U18279 (N_18279,N_11756,N_13445);
nand U18280 (N_18280,N_12190,N_14724);
and U18281 (N_18281,N_14733,N_12925);
or U18282 (N_18282,N_10320,N_13632);
or U18283 (N_18283,N_11678,N_14828);
or U18284 (N_18284,N_10122,N_10705);
nor U18285 (N_18285,N_13661,N_14680);
nand U18286 (N_18286,N_10689,N_10716);
and U18287 (N_18287,N_10176,N_11323);
nand U18288 (N_18288,N_10051,N_11576);
xnor U18289 (N_18289,N_11460,N_12250);
nor U18290 (N_18290,N_10801,N_12776);
xor U18291 (N_18291,N_13908,N_12915);
nand U18292 (N_18292,N_11751,N_14298);
and U18293 (N_18293,N_12665,N_13462);
nand U18294 (N_18294,N_10000,N_13469);
and U18295 (N_18295,N_11729,N_12884);
xor U18296 (N_18296,N_12453,N_14397);
nor U18297 (N_18297,N_12350,N_11441);
nand U18298 (N_18298,N_12191,N_14150);
or U18299 (N_18299,N_11656,N_12011);
nand U18300 (N_18300,N_11484,N_11804);
and U18301 (N_18301,N_12425,N_11640);
or U18302 (N_18302,N_12305,N_11448);
and U18303 (N_18303,N_13132,N_13362);
xnor U18304 (N_18304,N_13860,N_14306);
nor U18305 (N_18305,N_14840,N_12257);
and U18306 (N_18306,N_12682,N_10586);
nor U18307 (N_18307,N_13334,N_12905);
xnor U18308 (N_18308,N_10087,N_11076);
nand U18309 (N_18309,N_10112,N_13073);
or U18310 (N_18310,N_12863,N_13385);
and U18311 (N_18311,N_12665,N_11651);
or U18312 (N_18312,N_13728,N_13330);
xnor U18313 (N_18313,N_12868,N_14405);
or U18314 (N_18314,N_10429,N_12392);
nor U18315 (N_18315,N_12371,N_11570);
nand U18316 (N_18316,N_13890,N_14664);
or U18317 (N_18317,N_11346,N_10830);
or U18318 (N_18318,N_14265,N_14642);
nor U18319 (N_18319,N_10603,N_14671);
nor U18320 (N_18320,N_13757,N_10218);
nor U18321 (N_18321,N_10147,N_12454);
nor U18322 (N_18322,N_13693,N_14214);
or U18323 (N_18323,N_12210,N_12048);
nand U18324 (N_18324,N_14728,N_12366);
nor U18325 (N_18325,N_13765,N_11862);
and U18326 (N_18326,N_11553,N_13855);
or U18327 (N_18327,N_10053,N_10983);
xor U18328 (N_18328,N_14011,N_12331);
or U18329 (N_18329,N_14922,N_13867);
nand U18330 (N_18330,N_10764,N_13873);
or U18331 (N_18331,N_10053,N_10271);
and U18332 (N_18332,N_11551,N_12139);
and U18333 (N_18333,N_11522,N_11311);
and U18334 (N_18334,N_10364,N_13842);
xnor U18335 (N_18335,N_11770,N_14385);
or U18336 (N_18336,N_13803,N_14597);
or U18337 (N_18337,N_10912,N_10594);
or U18338 (N_18338,N_10397,N_11381);
nand U18339 (N_18339,N_10054,N_10011);
and U18340 (N_18340,N_13061,N_14022);
and U18341 (N_18341,N_11583,N_11321);
nand U18342 (N_18342,N_13793,N_14669);
or U18343 (N_18343,N_12626,N_12439);
nand U18344 (N_18344,N_14256,N_14540);
nor U18345 (N_18345,N_11977,N_10631);
nor U18346 (N_18346,N_12638,N_13412);
and U18347 (N_18347,N_13302,N_10204);
nor U18348 (N_18348,N_11318,N_11455);
and U18349 (N_18349,N_12900,N_12249);
nand U18350 (N_18350,N_10191,N_12169);
xnor U18351 (N_18351,N_12730,N_14626);
nand U18352 (N_18352,N_13951,N_10609);
or U18353 (N_18353,N_14573,N_14118);
and U18354 (N_18354,N_14375,N_11988);
or U18355 (N_18355,N_14659,N_14990);
nor U18356 (N_18356,N_13539,N_11580);
or U18357 (N_18357,N_12851,N_13324);
and U18358 (N_18358,N_10987,N_14493);
xnor U18359 (N_18359,N_13128,N_14405);
nand U18360 (N_18360,N_10358,N_12302);
xnor U18361 (N_18361,N_11967,N_12313);
and U18362 (N_18362,N_10447,N_13012);
nor U18363 (N_18363,N_11676,N_13879);
and U18364 (N_18364,N_10978,N_10579);
and U18365 (N_18365,N_13691,N_11753);
xor U18366 (N_18366,N_12645,N_10608);
xor U18367 (N_18367,N_12884,N_13821);
xor U18368 (N_18368,N_11065,N_14253);
or U18369 (N_18369,N_13085,N_10929);
xor U18370 (N_18370,N_10688,N_10278);
xor U18371 (N_18371,N_12856,N_13545);
xnor U18372 (N_18372,N_14262,N_12333);
xor U18373 (N_18373,N_10496,N_14553);
nor U18374 (N_18374,N_11316,N_13363);
or U18375 (N_18375,N_10683,N_14625);
xor U18376 (N_18376,N_14444,N_13903);
and U18377 (N_18377,N_11178,N_12031);
or U18378 (N_18378,N_13929,N_10626);
and U18379 (N_18379,N_14207,N_13051);
nand U18380 (N_18380,N_14296,N_14138);
or U18381 (N_18381,N_14996,N_13741);
nor U18382 (N_18382,N_14330,N_13435);
xnor U18383 (N_18383,N_13527,N_13383);
or U18384 (N_18384,N_12992,N_10259);
and U18385 (N_18385,N_11255,N_13598);
and U18386 (N_18386,N_12353,N_12054);
xnor U18387 (N_18387,N_12146,N_10858);
nand U18388 (N_18388,N_14092,N_14619);
nor U18389 (N_18389,N_11959,N_10822);
nor U18390 (N_18390,N_12399,N_10043);
nand U18391 (N_18391,N_10954,N_11768);
nor U18392 (N_18392,N_13140,N_14767);
xor U18393 (N_18393,N_11964,N_13952);
nor U18394 (N_18394,N_11147,N_14680);
or U18395 (N_18395,N_10880,N_13028);
xor U18396 (N_18396,N_14656,N_10417);
or U18397 (N_18397,N_11938,N_11823);
and U18398 (N_18398,N_10692,N_11430);
or U18399 (N_18399,N_11753,N_12047);
and U18400 (N_18400,N_10673,N_14861);
and U18401 (N_18401,N_14260,N_11296);
nor U18402 (N_18402,N_14299,N_14669);
nor U18403 (N_18403,N_12444,N_11267);
nor U18404 (N_18404,N_11583,N_10654);
and U18405 (N_18405,N_12076,N_12575);
xnor U18406 (N_18406,N_11729,N_13594);
and U18407 (N_18407,N_12223,N_13895);
nand U18408 (N_18408,N_11109,N_12799);
nand U18409 (N_18409,N_11336,N_10056);
nor U18410 (N_18410,N_13637,N_10351);
nand U18411 (N_18411,N_12410,N_11276);
nor U18412 (N_18412,N_12643,N_12116);
and U18413 (N_18413,N_12704,N_12388);
xnor U18414 (N_18414,N_13115,N_14261);
or U18415 (N_18415,N_12293,N_14402);
nor U18416 (N_18416,N_12665,N_12637);
nand U18417 (N_18417,N_14888,N_12916);
xor U18418 (N_18418,N_10124,N_10574);
nor U18419 (N_18419,N_12261,N_12157);
nor U18420 (N_18420,N_12382,N_11095);
nor U18421 (N_18421,N_12711,N_13426);
xnor U18422 (N_18422,N_12818,N_12202);
nor U18423 (N_18423,N_11710,N_10690);
or U18424 (N_18424,N_14490,N_12764);
xnor U18425 (N_18425,N_11307,N_12524);
nand U18426 (N_18426,N_10080,N_13308);
nor U18427 (N_18427,N_10171,N_11462);
nand U18428 (N_18428,N_12689,N_10383);
or U18429 (N_18429,N_14425,N_13916);
nor U18430 (N_18430,N_12702,N_13742);
nand U18431 (N_18431,N_11958,N_14665);
xor U18432 (N_18432,N_14642,N_11351);
nor U18433 (N_18433,N_11115,N_14849);
or U18434 (N_18434,N_10775,N_13572);
nor U18435 (N_18435,N_11326,N_11334);
nand U18436 (N_18436,N_11982,N_12943);
xnor U18437 (N_18437,N_14406,N_14515);
xnor U18438 (N_18438,N_10517,N_10616);
or U18439 (N_18439,N_10355,N_12154);
nor U18440 (N_18440,N_10716,N_14983);
nand U18441 (N_18441,N_13130,N_11047);
or U18442 (N_18442,N_11165,N_11323);
nor U18443 (N_18443,N_10753,N_10211);
and U18444 (N_18444,N_14290,N_14696);
nand U18445 (N_18445,N_14677,N_14503);
and U18446 (N_18446,N_12576,N_10024);
xnor U18447 (N_18447,N_10242,N_11682);
xor U18448 (N_18448,N_11113,N_14103);
or U18449 (N_18449,N_13149,N_11179);
and U18450 (N_18450,N_12208,N_13751);
or U18451 (N_18451,N_11322,N_14928);
nand U18452 (N_18452,N_11457,N_12667);
nand U18453 (N_18453,N_10675,N_13060);
nand U18454 (N_18454,N_14626,N_10409);
nand U18455 (N_18455,N_13068,N_13324);
nor U18456 (N_18456,N_14366,N_11166);
and U18457 (N_18457,N_10267,N_14965);
or U18458 (N_18458,N_13489,N_13038);
nor U18459 (N_18459,N_10040,N_10714);
nor U18460 (N_18460,N_11695,N_11943);
and U18461 (N_18461,N_13140,N_10237);
or U18462 (N_18462,N_10700,N_13170);
and U18463 (N_18463,N_14298,N_12968);
nand U18464 (N_18464,N_13522,N_14415);
xnor U18465 (N_18465,N_11069,N_10131);
and U18466 (N_18466,N_12750,N_14014);
or U18467 (N_18467,N_14080,N_13558);
nand U18468 (N_18468,N_11144,N_14075);
and U18469 (N_18469,N_10466,N_10833);
nor U18470 (N_18470,N_13434,N_12835);
or U18471 (N_18471,N_12211,N_12097);
xnor U18472 (N_18472,N_10480,N_12052);
xor U18473 (N_18473,N_14740,N_13865);
nor U18474 (N_18474,N_12258,N_12402);
and U18475 (N_18475,N_13335,N_11290);
and U18476 (N_18476,N_13573,N_10145);
nor U18477 (N_18477,N_10241,N_13276);
nor U18478 (N_18478,N_13628,N_13412);
and U18479 (N_18479,N_14138,N_12536);
and U18480 (N_18480,N_12488,N_14209);
and U18481 (N_18481,N_14970,N_11026);
nand U18482 (N_18482,N_14570,N_13679);
nand U18483 (N_18483,N_12904,N_14052);
nand U18484 (N_18484,N_13762,N_12011);
nand U18485 (N_18485,N_14891,N_11881);
and U18486 (N_18486,N_10082,N_10546);
nand U18487 (N_18487,N_14309,N_10360);
nand U18488 (N_18488,N_13421,N_12624);
nor U18489 (N_18489,N_14119,N_14306);
xnor U18490 (N_18490,N_13857,N_12080);
or U18491 (N_18491,N_12971,N_10906);
xnor U18492 (N_18492,N_11395,N_13881);
xnor U18493 (N_18493,N_11402,N_10546);
nand U18494 (N_18494,N_10870,N_10886);
xor U18495 (N_18495,N_10283,N_10994);
nand U18496 (N_18496,N_12925,N_14546);
nand U18497 (N_18497,N_14037,N_13561);
and U18498 (N_18498,N_14979,N_12013);
or U18499 (N_18499,N_10121,N_10482);
and U18500 (N_18500,N_10848,N_10414);
xnor U18501 (N_18501,N_14077,N_13755);
xnor U18502 (N_18502,N_13362,N_14711);
xnor U18503 (N_18503,N_14555,N_14284);
xnor U18504 (N_18504,N_12624,N_14097);
nand U18505 (N_18505,N_12236,N_11175);
xor U18506 (N_18506,N_12701,N_13502);
xnor U18507 (N_18507,N_10552,N_10928);
or U18508 (N_18508,N_12076,N_11400);
nand U18509 (N_18509,N_13687,N_14433);
xor U18510 (N_18510,N_13952,N_13260);
xor U18511 (N_18511,N_11931,N_14856);
xnor U18512 (N_18512,N_13710,N_12864);
xor U18513 (N_18513,N_11463,N_14197);
nand U18514 (N_18514,N_12866,N_12560);
nand U18515 (N_18515,N_13363,N_12371);
or U18516 (N_18516,N_14192,N_12676);
or U18517 (N_18517,N_11205,N_13047);
and U18518 (N_18518,N_13884,N_13459);
and U18519 (N_18519,N_13125,N_12887);
nor U18520 (N_18520,N_14839,N_11912);
nor U18521 (N_18521,N_12693,N_11741);
nor U18522 (N_18522,N_12480,N_13370);
nor U18523 (N_18523,N_13051,N_14079);
nor U18524 (N_18524,N_11898,N_12030);
and U18525 (N_18525,N_10667,N_13916);
and U18526 (N_18526,N_13134,N_12322);
and U18527 (N_18527,N_12518,N_13995);
or U18528 (N_18528,N_12760,N_13916);
nand U18529 (N_18529,N_14437,N_13384);
or U18530 (N_18530,N_11792,N_12729);
and U18531 (N_18531,N_13911,N_13800);
nor U18532 (N_18532,N_13116,N_12507);
and U18533 (N_18533,N_11584,N_14430);
nand U18534 (N_18534,N_11387,N_10780);
nand U18535 (N_18535,N_11136,N_11416);
and U18536 (N_18536,N_13847,N_11685);
or U18537 (N_18537,N_13871,N_11573);
xor U18538 (N_18538,N_10912,N_10113);
or U18539 (N_18539,N_13407,N_12220);
xnor U18540 (N_18540,N_12862,N_12373);
nor U18541 (N_18541,N_10415,N_14850);
or U18542 (N_18542,N_12262,N_13979);
or U18543 (N_18543,N_12331,N_14379);
or U18544 (N_18544,N_13291,N_14687);
and U18545 (N_18545,N_14876,N_10400);
nor U18546 (N_18546,N_12061,N_11901);
and U18547 (N_18547,N_13132,N_10999);
and U18548 (N_18548,N_10159,N_12691);
and U18549 (N_18549,N_11370,N_14632);
or U18550 (N_18550,N_14472,N_13647);
and U18551 (N_18551,N_13886,N_12505);
and U18552 (N_18552,N_14062,N_12770);
xor U18553 (N_18553,N_13551,N_14387);
or U18554 (N_18554,N_14861,N_11232);
and U18555 (N_18555,N_12588,N_13594);
and U18556 (N_18556,N_12109,N_11293);
or U18557 (N_18557,N_12187,N_12952);
nor U18558 (N_18558,N_11687,N_13570);
nor U18559 (N_18559,N_11716,N_10109);
xor U18560 (N_18560,N_14665,N_11463);
nor U18561 (N_18561,N_13625,N_11682);
and U18562 (N_18562,N_14749,N_10163);
or U18563 (N_18563,N_12477,N_10594);
and U18564 (N_18564,N_12394,N_12392);
nand U18565 (N_18565,N_10740,N_11591);
nor U18566 (N_18566,N_14066,N_10292);
nor U18567 (N_18567,N_14652,N_12608);
nor U18568 (N_18568,N_11424,N_13306);
xor U18569 (N_18569,N_13647,N_12431);
nand U18570 (N_18570,N_11616,N_11894);
nand U18571 (N_18571,N_12597,N_14779);
xor U18572 (N_18572,N_12712,N_10542);
or U18573 (N_18573,N_11593,N_12098);
and U18574 (N_18574,N_11156,N_12562);
nor U18575 (N_18575,N_10567,N_13954);
nand U18576 (N_18576,N_11570,N_11711);
nor U18577 (N_18577,N_11869,N_10842);
xnor U18578 (N_18578,N_14000,N_14451);
xor U18579 (N_18579,N_10394,N_14282);
nor U18580 (N_18580,N_12632,N_12306);
nand U18581 (N_18581,N_10478,N_12296);
or U18582 (N_18582,N_11089,N_10162);
or U18583 (N_18583,N_14188,N_10612);
nor U18584 (N_18584,N_11254,N_12025);
or U18585 (N_18585,N_14852,N_12539);
nor U18586 (N_18586,N_13553,N_11572);
or U18587 (N_18587,N_14690,N_11861);
nor U18588 (N_18588,N_10137,N_12634);
nand U18589 (N_18589,N_11449,N_12361);
nor U18590 (N_18590,N_11146,N_11114);
and U18591 (N_18591,N_12424,N_11420);
nand U18592 (N_18592,N_11084,N_14325);
nand U18593 (N_18593,N_13606,N_14895);
nor U18594 (N_18594,N_13497,N_14003);
nand U18595 (N_18595,N_14827,N_11615);
and U18596 (N_18596,N_13077,N_10189);
nor U18597 (N_18597,N_11824,N_13227);
and U18598 (N_18598,N_13325,N_13531);
nor U18599 (N_18599,N_13852,N_10852);
nor U18600 (N_18600,N_11996,N_11805);
and U18601 (N_18601,N_14573,N_14383);
nor U18602 (N_18602,N_10038,N_13770);
and U18603 (N_18603,N_10796,N_13980);
xor U18604 (N_18604,N_10316,N_13579);
nand U18605 (N_18605,N_12928,N_14501);
or U18606 (N_18606,N_13552,N_12895);
and U18607 (N_18607,N_10130,N_14634);
and U18608 (N_18608,N_13616,N_13307);
and U18609 (N_18609,N_11417,N_13644);
xnor U18610 (N_18610,N_12430,N_13065);
and U18611 (N_18611,N_12643,N_11780);
nor U18612 (N_18612,N_14539,N_12047);
nor U18613 (N_18613,N_14062,N_10503);
and U18614 (N_18614,N_12650,N_11250);
or U18615 (N_18615,N_11953,N_14836);
and U18616 (N_18616,N_10297,N_12796);
nand U18617 (N_18617,N_14768,N_14350);
nand U18618 (N_18618,N_13709,N_14816);
and U18619 (N_18619,N_13467,N_12949);
nand U18620 (N_18620,N_13531,N_12294);
or U18621 (N_18621,N_14759,N_11648);
and U18622 (N_18622,N_10051,N_11982);
or U18623 (N_18623,N_10845,N_13982);
or U18624 (N_18624,N_14566,N_12623);
or U18625 (N_18625,N_10991,N_11198);
nor U18626 (N_18626,N_10151,N_12274);
nand U18627 (N_18627,N_13239,N_12166);
xnor U18628 (N_18628,N_12585,N_13029);
nand U18629 (N_18629,N_10216,N_10309);
or U18630 (N_18630,N_11435,N_10480);
xor U18631 (N_18631,N_14487,N_14356);
xnor U18632 (N_18632,N_13866,N_10150);
nand U18633 (N_18633,N_14854,N_12747);
xor U18634 (N_18634,N_14134,N_14096);
and U18635 (N_18635,N_10009,N_12210);
nor U18636 (N_18636,N_14586,N_10660);
nor U18637 (N_18637,N_14883,N_14868);
or U18638 (N_18638,N_12675,N_12266);
xnor U18639 (N_18639,N_10878,N_12320);
nor U18640 (N_18640,N_10029,N_10413);
and U18641 (N_18641,N_12358,N_11575);
or U18642 (N_18642,N_14881,N_12103);
and U18643 (N_18643,N_14011,N_12247);
nand U18644 (N_18644,N_13456,N_14146);
and U18645 (N_18645,N_10057,N_10835);
nand U18646 (N_18646,N_11218,N_11723);
xnor U18647 (N_18647,N_13632,N_12683);
nor U18648 (N_18648,N_12277,N_14345);
or U18649 (N_18649,N_12298,N_13938);
nand U18650 (N_18650,N_12895,N_13190);
and U18651 (N_18651,N_10841,N_10207);
nor U18652 (N_18652,N_13215,N_10393);
or U18653 (N_18653,N_14081,N_13696);
and U18654 (N_18654,N_11175,N_11650);
xnor U18655 (N_18655,N_12173,N_13545);
nor U18656 (N_18656,N_14432,N_13261);
xnor U18657 (N_18657,N_10546,N_13700);
nor U18658 (N_18658,N_11828,N_12912);
nand U18659 (N_18659,N_11109,N_12563);
or U18660 (N_18660,N_12296,N_12532);
nand U18661 (N_18661,N_10817,N_10077);
or U18662 (N_18662,N_13774,N_12906);
xnor U18663 (N_18663,N_10057,N_13516);
nand U18664 (N_18664,N_12619,N_14575);
xnor U18665 (N_18665,N_13759,N_10065);
and U18666 (N_18666,N_14760,N_12026);
nor U18667 (N_18667,N_14640,N_14939);
and U18668 (N_18668,N_14549,N_13631);
nand U18669 (N_18669,N_11936,N_13100);
nand U18670 (N_18670,N_14732,N_11688);
nor U18671 (N_18671,N_12257,N_11669);
or U18672 (N_18672,N_10072,N_10155);
and U18673 (N_18673,N_13859,N_13606);
nor U18674 (N_18674,N_12336,N_13930);
nand U18675 (N_18675,N_13494,N_12221);
nand U18676 (N_18676,N_13869,N_12642);
xor U18677 (N_18677,N_12857,N_13102);
and U18678 (N_18678,N_12302,N_13805);
nor U18679 (N_18679,N_13823,N_13852);
and U18680 (N_18680,N_11790,N_12346);
xnor U18681 (N_18681,N_14613,N_13605);
nand U18682 (N_18682,N_10408,N_12459);
nor U18683 (N_18683,N_14712,N_10466);
nor U18684 (N_18684,N_12833,N_10929);
xnor U18685 (N_18685,N_11985,N_10080);
and U18686 (N_18686,N_12489,N_11936);
and U18687 (N_18687,N_13058,N_13613);
and U18688 (N_18688,N_13608,N_12842);
nor U18689 (N_18689,N_12039,N_13780);
or U18690 (N_18690,N_12277,N_13607);
nor U18691 (N_18691,N_14968,N_11940);
and U18692 (N_18692,N_10840,N_11662);
and U18693 (N_18693,N_14309,N_11536);
and U18694 (N_18694,N_10922,N_13576);
and U18695 (N_18695,N_12131,N_13899);
and U18696 (N_18696,N_12625,N_12397);
nor U18697 (N_18697,N_11757,N_13565);
or U18698 (N_18698,N_12825,N_12402);
nor U18699 (N_18699,N_14610,N_14772);
xor U18700 (N_18700,N_10561,N_12130);
xor U18701 (N_18701,N_14892,N_11650);
or U18702 (N_18702,N_10031,N_12577);
nor U18703 (N_18703,N_12443,N_14410);
or U18704 (N_18704,N_11000,N_11294);
nand U18705 (N_18705,N_13439,N_10288);
and U18706 (N_18706,N_12571,N_12772);
nor U18707 (N_18707,N_14270,N_11084);
or U18708 (N_18708,N_12549,N_14828);
nor U18709 (N_18709,N_14353,N_14897);
or U18710 (N_18710,N_10722,N_11084);
nor U18711 (N_18711,N_12805,N_14863);
xor U18712 (N_18712,N_10695,N_11426);
and U18713 (N_18713,N_10718,N_14160);
and U18714 (N_18714,N_11255,N_12175);
xnor U18715 (N_18715,N_12186,N_13200);
nand U18716 (N_18716,N_12482,N_12718);
nor U18717 (N_18717,N_13319,N_14944);
nor U18718 (N_18718,N_14545,N_11573);
nand U18719 (N_18719,N_11888,N_14271);
and U18720 (N_18720,N_14747,N_10745);
or U18721 (N_18721,N_13242,N_13895);
and U18722 (N_18722,N_11168,N_12314);
or U18723 (N_18723,N_10066,N_13455);
nor U18724 (N_18724,N_13707,N_11676);
xor U18725 (N_18725,N_13227,N_13801);
nor U18726 (N_18726,N_14487,N_11778);
and U18727 (N_18727,N_11741,N_10725);
or U18728 (N_18728,N_11902,N_13120);
or U18729 (N_18729,N_13550,N_12060);
nor U18730 (N_18730,N_11618,N_14363);
nor U18731 (N_18731,N_12113,N_10376);
xor U18732 (N_18732,N_14287,N_13557);
or U18733 (N_18733,N_13805,N_10087);
or U18734 (N_18734,N_14480,N_14703);
nand U18735 (N_18735,N_14531,N_13351);
nand U18736 (N_18736,N_12215,N_13301);
or U18737 (N_18737,N_12444,N_11881);
xor U18738 (N_18738,N_11071,N_13079);
or U18739 (N_18739,N_13583,N_13615);
xnor U18740 (N_18740,N_12551,N_10172);
nand U18741 (N_18741,N_10729,N_10538);
xnor U18742 (N_18742,N_12388,N_13394);
or U18743 (N_18743,N_14147,N_14349);
nor U18744 (N_18744,N_12654,N_11614);
nor U18745 (N_18745,N_11502,N_12612);
or U18746 (N_18746,N_13116,N_14477);
xnor U18747 (N_18747,N_14686,N_11042);
xor U18748 (N_18748,N_14519,N_11069);
xnor U18749 (N_18749,N_10756,N_11091);
xor U18750 (N_18750,N_10278,N_11911);
nor U18751 (N_18751,N_12282,N_10090);
and U18752 (N_18752,N_13272,N_13948);
or U18753 (N_18753,N_14132,N_11568);
xnor U18754 (N_18754,N_14574,N_12813);
and U18755 (N_18755,N_13990,N_12921);
or U18756 (N_18756,N_10994,N_11960);
and U18757 (N_18757,N_11751,N_11103);
nand U18758 (N_18758,N_11701,N_10589);
xnor U18759 (N_18759,N_14641,N_14527);
xnor U18760 (N_18760,N_13047,N_10368);
or U18761 (N_18761,N_14235,N_12617);
nor U18762 (N_18762,N_13218,N_14978);
or U18763 (N_18763,N_14950,N_12187);
nor U18764 (N_18764,N_13825,N_10121);
xnor U18765 (N_18765,N_12362,N_13495);
or U18766 (N_18766,N_10762,N_14253);
nand U18767 (N_18767,N_13332,N_12590);
and U18768 (N_18768,N_13891,N_14386);
nand U18769 (N_18769,N_13791,N_11015);
nor U18770 (N_18770,N_10840,N_12362);
xnor U18771 (N_18771,N_10336,N_12401);
xor U18772 (N_18772,N_11341,N_10594);
nand U18773 (N_18773,N_11889,N_14708);
and U18774 (N_18774,N_13549,N_11973);
xor U18775 (N_18775,N_13873,N_10581);
xor U18776 (N_18776,N_12805,N_14679);
or U18777 (N_18777,N_10267,N_12448);
or U18778 (N_18778,N_13903,N_14033);
xor U18779 (N_18779,N_13718,N_13949);
nand U18780 (N_18780,N_10219,N_12854);
and U18781 (N_18781,N_11449,N_10330);
and U18782 (N_18782,N_11981,N_12996);
nor U18783 (N_18783,N_14060,N_10713);
nand U18784 (N_18784,N_14256,N_11567);
xnor U18785 (N_18785,N_14326,N_11183);
nor U18786 (N_18786,N_10245,N_12022);
nor U18787 (N_18787,N_14346,N_13887);
nor U18788 (N_18788,N_13844,N_14945);
and U18789 (N_18789,N_11416,N_14229);
xor U18790 (N_18790,N_12272,N_10767);
xor U18791 (N_18791,N_11791,N_11553);
and U18792 (N_18792,N_12249,N_11348);
xor U18793 (N_18793,N_11374,N_14163);
and U18794 (N_18794,N_13683,N_10516);
nand U18795 (N_18795,N_14912,N_12837);
and U18796 (N_18796,N_10068,N_14321);
and U18797 (N_18797,N_10780,N_14607);
xor U18798 (N_18798,N_11040,N_12952);
and U18799 (N_18799,N_10845,N_11635);
xor U18800 (N_18800,N_13552,N_12159);
nand U18801 (N_18801,N_14455,N_14096);
nand U18802 (N_18802,N_13431,N_11390);
nor U18803 (N_18803,N_12328,N_10513);
nor U18804 (N_18804,N_12795,N_13546);
or U18805 (N_18805,N_14316,N_12694);
nor U18806 (N_18806,N_13792,N_12172);
xnor U18807 (N_18807,N_14537,N_12321);
and U18808 (N_18808,N_12195,N_13812);
nand U18809 (N_18809,N_12867,N_14976);
nor U18810 (N_18810,N_14239,N_10211);
nand U18811 (N_18811,N_10361,N_12550);
nand U18812 (N_18812,N_10665,N_10857);
nand U18813 (N_18813,N_11780,N_12329);
and U18814 (N_18814,N_14178,N_11431);
and U18815 (N_18815,N_11600,N_10893);
xor U18816 (N_18816,N_12400,N_10361);
xnor U18817 (N_18817,N_13494,N_14372);
and U18818 (N_18818,N_10986,N_10240);
or U18819 (N_18819,N_13339,N_11640);
nor U18820 (N_18820,N_10573,N_10686);
or U18821 (N_18821,N_13581,N_10959);
and U18822 (N_18822,N_11687,N_14082);
or U18823 (N_18823,N_11850,N_13839);
nor U18824 (N_18824,N_12042,N_10158);
nor U18825 (N_18825,N_12110,N_10298);
nor U18826 (N_18826,N_13131,N_12134);
xnor U18827 (N_18827,N_11773,N_12685);
nand U18828 (N_18828,N_12010,N_11383);
xnor U18829 (N_18829,N_12138,N_10466);
nor U18830 (N_18830,N_13372,N_10983);
nand U18831 (N_18831,N_11848,N_10650);
xnor U18832 (N_18832,N_14916,N_12054);
or U18833 (N_18833,N_12464,N_14676);
nor U18834 (N_18834,N_12897,N_13039);
xor U18835 (N_18835,N_11789,N_14442);
nor U18836 (N_18836,N_12792,N_10847);
or U18837 (N_18837,N_14800,N_10243);
and U18838 (N_18838,N_14746,N_10561);
nor U18839 (N_18839,N_11548,N_12148);
or U18840 (N_18840,N_10827,N_13693);
nand U18841 (N_18841,N_12095,N_14679);
xnor U18842 (N_18842,N_14440,N_13149);
and U18843 (N_18843,N_11351,N_14473);
and U18844 (N_18844,N_14830,N_13445);
xnor U18845 (N_18845,N_12486,N_13238);
nand U18846 (N_18846,N_11111,N_10236);
or U18847 (N_18847,N_12744,N_12769);
nor U18848 (N_18848,N_12335,N_11804);
nor U18849 (N_18849,N_10524,N_14118);
nor U18850 (N_18850,N_12965,N_14036);
or U18851 (N_18851,N_11291,N_13342);
nor U18852 (N_18852,N_14023,N_13478);
nor U18853 (N_18853,N_11739,N_14135);
xnor U18854 (N_18854,N_10235,N_10605);
nand U18855 (N_18855,N_11711,N_11994);
and U18856 (N_18856,N_11249,N_13348);
or U18857 (N_18857,N_13547,N_14966);
and U18858 (N_18858,N_11843,N_14270);
and U18859 (N_18859,N_14784,N_12792);
or U18860 (N_18860,N_14973,N_10186);
xnor U18861 (N_18861,N_12245,N_13013);
nand U18862 (N_18862,N_11942,N_11042);
nor U18863 (N_18863,N_12217,N_13785);
nand U18864 (N_18864,N_13745,N_13645);
nand U18865 (N_18865,N_11518,N_14230);
xor U18866 (N_18866,N_13378,N_10232);
or U18867 (N_18867,N_13653,N_12495);
and U18868 (N_18868,N_11333,N_10629);
nor U18869 (N_18869,N_11846,N_11750);
xnor U18870 (N_18870,N_11684,N_14390);
or U18871 (N_18871,N_12875,N_10766);
xor U18872 (N_18872,N_14260,N_13002);
or U18873 (N_18873,N_10819,N_13013);
nand U18874 (N_18874,N_12214,N_10156);
nor U18875 (N_18875,N_14715,N_11738);
and U18876 (N_18876,N_14434,N_13111);
or U18877 (N_18877,N_11617,N_11247);
or U18878 (N_18878,N_10436,N_13401);
xor U18879 (N_18879,N_10961,N_14482);
nand U18880 (N_18880,N_14324,N_14752);
nor U18881 (N_18881,N_12814,N_12245);
xnor U18882 (N_18882,N_10875,N_13100);
xor U18883 (N_18883,N_13777,N_12871);
nand U18884 (N_18884,N_10800,N_12683);
xor U18885 (N_18885,N_13774,N_11833);
nand U18886 (N_18886,N_12953,N_13416);
and U18887 (N_18887,N_13067,N_13138);
nor U18888 (N_18888,N_10851,N_10537);
and U18889 (N_18889,N_12926,N_13088);
and U18890 (N_18890,N_11129,N_11653);
or U18891 (N_18891,N_13494,N_13884);
and U18892 (N_18892,N_14557,N_11289);
or U18893 (N_18893,N_13881,N_10832);
nand U18894 (N_18894,N_10007,N_12148);
or U18895 (N_18895,N_12130,N_12442);
nand U18896 (N_18896,N_12499,N_13855);
nor U18897 (N_18897,N_13276,N_11136);
nand U18898 (N_18898,N_10703,N_11682);
and U18899 (N_18899,N_11432,N_14794);
xnor U18900 (N_18900,N_10009,N_12936);
nor U18901 (N_18901,N_14883,N_14099);
xor U18902 (N_18902,N_12933,N_12514);
xor U18903 (N_18903,N_10480,N_10420);
and U18904 (N_18904,N_10638,N_13370);
and U18905 (N_18905,N_14884,N_10612);
xnor U18906 (N_18906,N_11973,N_14740);
nor U18907 (N_18907,N_13562,N_10152);
nand U18908 (N_18908,N_14056,N_10812);
xnor U18909 (N_18909,N_11302,N_14612);
or U18910 (N_18910,N_13577,N_11987);
nand U18911 (N_18911,N_10931,N_11879);
xnor U18912 (N_18912,N_10274,N_12780);
nand U18913 (N_18913,N_12839,N_13730);
or U18914 (N_18914,N_14722,N_13765);
and U18915 (N_18915,N_12250,N_10412);
nand U18916 (N_18916,N_11336,N_12623);
nor U18917 (N_18917,N_10449,N_10104);
xor U18918 (N_18918,N_13529,N_11932);
nand U18919 (N_18919,N_10684,N_12014);
or U18920 (N_18920,N_12655,N_11527);
nand U18921 (N_18921,N_11111,N_13900);
xnor U18922 (N_18922,N_10805,N_12354);
nor U18923 (N_18923,N_11126,N_10564);
nor U18924 (N_18924,N_11563,N_12022);
nand U18925 (N_18925,N_13662,N_12965);
xor U18926 (N_18926,N_13691,N_14020);
nand U18927 (N_18927,N_11441,N_14152);
or U18928 (N_18928,N_13569,N_12905);
or U18929 (N_18929,N_11197,N_12585);
nand U18930 (N_18930,N_14957,N_11797);
or U18931 (N_18931,N_13018,N_13675);
nand U18932 (N_18932,N_12817,N_11863);
or U18933 (N_18933,N_11569,N_12283);
nor U18934 (N_18934,N_11908,N_14325);
or U18935 (N_18935,N_10282,N_10368);
nand U18936 (N_18936,N_13558,N_13803);
nand U18937 (N_18937,N_12395,N_10809);
and U18938 (N_18938,N_13132,N_14999);
xor U18939 (N_18939,N_14409,N_12274);
or U18940 (N_18940,N_10812,N_14998);
and U18941 (N_18941,N_11510,N_13524);
nor U18942 (N_18942,N_11765,N_14743);
and U18943 (N_18943,N_14443,N_11380);
nand U18944 (N_18944,N_12737,N_14921);
nand U18945 (N_18945,N_14794,N_10354);
and U18946 (N_18946,N_14981,N_14881);
xnor U18947 (N_18947,N_13873,N_14116);
or U18948 (N_18948,N_11177,N_13263);
nand U18949 (N_18949,N_13988,N_11188);
xnor U18950 (N_18950,N_14865,N_11910);
nor U18951 (N_18951,N_13592,N_14324);
and U18952 (N_18952,N_11439,N_12667);
xnor U18953 (N_18953,N_11077,N_12033);
or U18954 (N_18954,N_11678,N_12604);
nor U18955 (N_18955,N_11686,N_13176);
or U18956 (N_18956,N_13979,N_10056);
nand U18957 (N_18957,N_13286,N_13373);
or U18958 (N_18958,N_12495,N_10679);
nand U18959 (N_18959,N_14295,N_10197);
and U18960 (N_18960,N_12191,N_12302);
xor U18961 (N_18961,N_12264,N_14734);
nand U18962 (N_18962,N_12736,N_12155);
xnor U18963 (N_18963,N_13945,N_10575);
and U18964 (N_18964,N_12973,N_11205);
and U18965 (N_18965,N_13705,N_12086);
xor U18966 (N_18966,N_11724,N_10703);
nor U18967 (N_18967,N_12125,N_11788);
nand U18968 (N_18968,N_12437,N_10874);
and U18969 (N_18969,N_14699,N_12598);
nand U18970 (N_18970,N_14433,N_12069);
xnor U18971 (N_18971,N_13008,N_14773);
nand U18972 (N_18972,N_10886,N_12375);
or U18973 (N_18973,N_12673,N_11698);
or U18974 (N_18974,N_14438,N_13898);
nand U18975 (N_18975,N_11294,N_10538);
xnor U18976 (N_18976,N_13947,N_14205);
and U18977 (N_18977,N_12209,N_13732);
xor U18978 (N_18978,N_11065,N_12552);
and U18979 (N_18979,N_12584,N_13030);
or U18980 (N_18980,N_10790,N_10276);
or U18981 (N_18981,N_14462,N_14411);
and U18982 (N_18982,N_10291,N_14744);
nand U18983 (N_18983,N_13252,N_12717);
and U18984 (N_18984,N_14792,N_11330);
and U18985 (N_18985,N_12525,N_11585);
or U18986 (N_18986,N_11923,N_10973);
nor U18987 (N_18987,N_11610,N_14146);
or U18988 (N_18988,N_11359,N_14005);
and U18989 (N_18989,N_12683,N_11142);
and U18990 (N_18990,N_10263,N_13983);
nand U18991 (N_18991,N_12493,N_11337);
and U18992 (N_18992,N_14804,N_13288);
or U18993 (N_18993,N_12897,N_13072);
nand U18994 (N_18994,N_13770,N_12481);
nor U18995 (N_18995,N_10591,N_12360);
nand U18996 (N_18996,N_11045,N_12757);
nand U18997 (N_18997,N_12986,N_13049);
and U18998 (N_18998,N_12827,N_10319);
or U18999 (N_18999,N_14019,N_14022);
nor U19000 (N_19000,N_11853,N_12654);
xnor U19001 (N_19001,N_10150,N_13675);
and U19002 (N_19002,N_11956,N_14595);
and U19003 (N_19003,N_14017,N_14535);
nand U19004 (N_19004,N_11921,N_14007);
and U19005 (N_19005,N_14415,N_14272);
or U19006 (N_19006,N_12976,N_11515);
nand U19007 (N_19007,N_11405,N_10472);
and U19008 (N_19008,N_10525,N_11972);
nor U19009 (N_19009,N_13683,N_10270);
xnor U19010 (N_19010,N_13955,N_10087);
and U19011 (N_19011,N_12426,N_11776);
nor U19012 (N_19012,N_14152,N_11646);
or U19013 (N_19013,N_10068,N_10279);
nor U19014 (N_19014,N_14809,N_12563);
nor U19015 (N_19015,N_10297,N_11585);
nor U19016 (N_19016,N_11776,N_10527);
nand U19017 (N_19017,N_13215,N_13163);
or U19018 (N_19018,N_11778,N_12513);
xnor U19019 (N_19019,N_10021,N_14446);
nand U19020 (N_19020,N_13016,N_13334);
nand U19021 (N_19021,N_12798,N_11831);
and U19022 (N_19022,N_14297,N_14405);
xnor U19023 (N_19023,N_10437,N_11248);
and U19024 (N_19024,N_10530,N_10857);
xor U19025 (N_19025,N_10668,N_10720);
nor U19026 (N_19026,N_10680,N_11949);
or U19027 (N_19027,N_14951,N_12766);
nor U19028 (N_19028,N_11562,N_11750);
nand U19029 (N_19029,N_11164,N_10261);
and U19030 (N_19030,N_10293,N_14350);
nor U19031 (N_19031,N_14654,N_14628);
nor U19032 (N_19032,N_12011,N_12837);
nand U19033 (N_19033,N_13775,N_11658);
and U19034 (N_19034,N_11340,N_14011);
nor U19035 (N_19035,N_11163,N_14851);
nor U19036 (N_19036,N_12078,N_13685);
xnor U19037 (N_19037,N_13052,N_11689);
or U19038 (N_19038,N_11321,N_13338);
nor U19039 (N_19039,N_11832,N_12552);
or U19040 (N_19040,N_12470,N_13501);
nor U19041 (N_19041,N_10169,N_12423);
and U19042 (N_19042,N_11043,N_11022);
nor U19043 (N_19043,N_11689,N_14594);
nand U19044 (N_19044,N_12459,N_14363);
and U19045 (N_19045,N_10413,N_10498);
xor U19046 (N_19046,N_12787,N_10355);
or U19047 (N_19047,N_13396,N_12605);
and U19048 (N_19048,N_14934,N_12486);
and U19049 (N_19049,N_13499,N_13296);
or U19050 (N_19050,N_13330,N_12797);
or U19051 (N_19051,N_11128,N_14691);
or U19052 (N_19052,N_11682,N_14140);
xor U19053 (N_19053,N_12498,N_11897);
nor U19054 (N_19054,N_14062,N_10159);
nor U19055 (N_19055,N_11903,N_14040);
or U19056 (N_19056,N_11369,N_11919);
and U19057 (N_19057,N_13975,N_14115);
xor U19058 (N_19058,N_14838,N_12096);
nor U19059 (N_19059,N_12595,N_13027);
nand U19060 (N_19060,N_12207,N_12507);
nor U19061 (N_19061,N_10404,N_10835);
nor U19062 (N_19062,N_11117,N_14035);
nand U19063 (N_19063,N_13257,N_13193);
nor U19064 (N_19064,N_14415,N_13724);
xnor U19065 (N_19065,N_13779,N_10921);
or U19066 (N_19066,N_11156,N_14994);
xnor U19067 (N_19067,N_10475,N_10133);
or U19068 (N_19068,N_12935,N_11828);
nand U19069 (N_19069,N_11024,N_10699);
and U19070 (N_19070,N_10278,N_12197);
xor U19071 (N_19071,N_13495,N_11992);
nor U19072 (N_19072,N_11577,N_13423);
nor U19073 (N_19073,N_10640,N_13330);
and U19074 (N_19074,N_11703,N_12351);
or U19075 (N_19075,N_10833,N_14621);
nand U19076 (N_19076,N_10276,N_13730);
nor U19077 (N_19077,N_13786,N_14311);
or U19078 (N_19078,N_14197,N_14541);
or U19079 (N_19079,N_11021,N_12310);
xnor U19080 (N_19080,N_13149,N_11594);
nor U19081 (N_19081,N_11286,N_11200);
or U19082 (N_19082,N_10698,N_10547);
and U19083 (N_19083,N_14689,N_13475);
nor U19084 (N_19084,N_12784,N_11811);
or U19085 (N_19085,N_12215,N_13719);
nor U19086 (N_19086,N_13948,N_14596);
and U19087 (N_19087,N_10835,N_14120);
xor U19088 (N_19088,N_10950,N_14042);
and U19089 (N_19089,N_14111,N_12406);
or U19090 (N_19090,N_12435,N_12278);
and U19091 (N_19091,N_13437,N_12649);
nor U19092 (N_19092,N_10685,N_14622);
and U19093 (N_19093,N_13529,N_12458);
nand U19094 (N_19094,N_12331,N_10094);
and U19095 (N_19095,N_13959,N_11337);
nor U19096 (N_19096,N_11493,N_14727);
nor U19097 (N_19097,N_12932,N_10124);
or U19098 (N_19098,N_11791,N_11089);
nand U19099 (N_19099,N_10095,N_11672);
nand U19100 (N_19100,N_12617,N_12934);
xor U19101 (N_19101,N_11656,N_13004);
xnor U19102 (N_19102,N_12323,N_12789);
and U19103 (N_19103,N_14840,N_10228);
or U19104 (N_19104,N_10354,N_14287);
and U19105 (N_19105,N_14167,N_11310);
nor U19106 (N_19106,N_11413,N_12684);
nor U19107 (N_19107,N_14119,N_13954);
and U19108 (N_19108,N_10997,N_12443);
xor U19109 (N_19109,N_13933,N_12894);
nor U19110 (N_19110,N_12476,N_10594);
nor U19111 (N_19111,N_12228,N_12801);
and U19112 (N_19112,N_11050,N_12428);
nand U19113 (N_19113,N_13247,N_14131);
and U19114 (N_19114,N_12409,N_11217);
nor U19115 (N_19115,N_13519,N_10003);
or U19116 (N_19116,N_11524,N_13847);
or U19117 (N_19117,N_13555,N_13015);
xor U19118 (N_19118,N_13686,N_14757);
and U19119 (N_19119,N_11234,N_14554);
nand U19120 (N_19120,N_13130,N_12963);
xnor U19121 (N_19121,N_11684,N_14592);
or U19122 (N_19122,N_12608,N_13690);
and U19123 (N_19123,N_10934,N_14991);
nor U19124 (N_19124,N_12822,N_13654);
or U19125 (N_19125,N_11000,N_11113);
or U19126 (N_19126,N_13881,N_10422);
xor U19127 (N_19127,N_13758,N_14175);
nor U19128 (N_19128,N_10134,N_12549);
nor U19129 (N_19129,N_10194,N_10298);
and U19130 (N_19130,N_11710,N_12690);
nand U19131 (N_19131,N_13807,N_13357);
nor U19132 (N_19132,N_13742,N_11372);
and U19133 (N_19133,N_14706,N_11929);
and U19134 (N_19134,N_13161,N_12986);
and U19135 (N_19135,N_10791,N_13231);
and U19136 (N_19136,N_14863,N_13209);
nand U19137 (N_19137,N_12252,N_12815);
nor U19138 (N_19138,N_10899,N_12693);
xnor U19139 (N_19139,N_12410,N_11647);
nor U19140 (N_19140,N_12501,N_10844);
xnor U19141 (N_19141,N_14270,N_11341);
nand U19142 (N_19142,N_12097,N_14655);
nor U19143 (N_19143,N_12372,N_13889);
xnor U19144 (N_19144,N_14369,N_11617);
xor U19145 (N_19145,N_10249,N_13132);
xor U19146 (N_19146,N_11869,N_11210);
nor U19147 (N_19147,N_10729,N_13471);
nor U19148 (N_19148,N_14504,N_14561);
and U19149 (N_19149,N_12689,N_13065);
or U19150 (N_19150,N_12670,N_14078);
nand U19151 (N_19151,N_13216,N_12673);
or U19152 (N_19152,N_11680,N_12801);
nor U19153 (N_19153,N_12587,N_11012);
or U19154 (N_19154,N_11351,N_11301);
nand U19155 (N_19155,N_13909,N_13176);
and U19156 (N_19156,N_12240,N_10603);
nor U19157 (N_19157,N_10680,N_14064);
or U19158 (N_19158,N_11521,N_11282);
nand U19159 (N_19159,N_12021,N_10362);
nand U19160 (N_19160,N_10637,N_10453);
xor U19161 (N_19161,N_10399,N_12560);
nor U19162 (N_19162,N_13931,N_11755);
or U19163 (N_19163,N_13804,N_12038);
or U19164 (N_19164,N_12115,N_12340);
or U19165 (N_19165,N_13341,N_11585);
or U19166 (N_19166,N_12298,N_13454);
and U19167 (N_19167,N_10976,N_13382);
xnor U19168 (N_19168,N_14344,N_11262);
nor U19169 (N_19169,N_10585,N_14738);
or U19170 (N_19170,N_10212,N_11373);
and U19171 (N_19171,N_13134,N_10672);
and U19172 (N_19172,N_13986,N_11761);
or U19173 (N_19173,N_10221,N_11194);
xnor U19174 (N_19174,N_14217,N_12734);
xnor U19175 (N_19175,N_13094,N_12772);
nand U19176 (N_19176,N_14981,N_11561);
nand U19177 (N_19177,N_11494,N_12644);
xor U19178 (N_19178,N_14571,N_11991);
nand U19179 (N_19179,N_14003,N_13983);
xor U19180 (N_19180,N_10949,N_13235);
or U19181 (N_19181,N_12066,N_13644);
xor U19182 (N_19182,N_13356,N_11083);
or U19183 (N_19183,N_13601,N_13719);
xor U19184 (N_19184,N_10582,N_10100);
nand U19185 (N_19185,N_13808,N_14732);
nor U19186 (N_19186,N_14179,N_12928);
or U19187 (N_19187,N_12737,N_14962);
xnor U19188 (N_19188,N_12752,N_14649);
and U19189 (N_19189,N_10390,N_11906);
nor U19190 (N_19190,N_12060,N_10737);
nor U19191 (N_19191,N_12649,N_10053);
nor U19192 (N_19192,N_10878,N_11230);
xnor U19193 (N_19193,N_11394,N_11377);
xor U19194 (N_19194,N_13775,N_10621);
nand U19195 (N_19195,N_11528,N_10237);
or U19196 (N_19196,N_11531,N_12919);
xnor U19197 (N_19197,N_13365,N_10342);
nand U19198 (N_19198,N_10256,N_11133);
nand U19199 (N_19199,N_11475,N_14109);
or U19200 (N_19200,N_12425,N_11625);
nor U19201 (N_19201,N_11274,N_14838);
xnor U19202 (N_19202,N_14822,N_11600);
nand U19203 (N_19203,N_10312,N_12623);
or U19204 (N_19204,N_10936,N_13489);
or U19205 (N_19205,N_14203,N_10060);
or U19206 (N_19206,N_14247,N_14480);
and U19207 (N_19207,N_10400,N_11185);
nand U19208 (N_19208,N_13320,N_14912);
nand U19209 (N_19209,N_13498,N_11511);
nor U19210 (N_19210,N_10320,N_10889);
or U19211 (N_19211,N_10848,N_10868);
or U19212 (N_19212,N_11595,N_10082);
nand U19213 (N_19213,N_13044,N_10592);
nor U19214 (N_19214,N_11605,N_14461);
and U19215 (N_19215,N_13493,N_13097);
or U19216 (N_19216,N_11025,N_13078);
nor U19217 (N_19217,N_13558,N_11242);
or U19218 (N_19218,N_10090,N_11314);
nor U19219 (N_19219,N_14691,N_10386);
nand U19220 (N_19220,N_14743,N_11520);
xor U19221 (N_19221,N_10161,N_12486);
and U19222 (N_19222,N_13611,N_11047);
or U19223 (N_19223,N_13533,N_13127);
or U19224 (N_19224,N_13604,N_13428);
nor U19225 (N_19225,N_14294,N_12146);
or U19226 (N_19226,N_11764,N_10208);
or U19227 (N_19227,N_11227,N_14686);
or U19228 (N_19228,N_12259,N_12836);
nand U19229 (N_19229,N_12317,N_11531);
nor U19230 (N_19230,N_11043,N_11094);
nor U19231 (N_19231,N_10254,N_11453);
xor U19232 (N_19232,N_10379,N_10316);
or U19233 (N_19233,N_14601,N_11533);
and U19234 (N_19234,N_11461,N_12379);
xnor U19235 (N_19235,N_12640,N_14521);
or U19236 (N_19236,N_13564,N_10276);
nand U19237 (N_19237,N_12779,N_10033);
and U19238 (N_19238,N_12354,N_10003);
and U19239 (N_19239,N_12208,N_10386);
nor U19240 (N_19240,N_14547,N_10810);
xor U19241 (N_19241,N_13092,N_10111);
and U19242 (N_19242,N_11872,N_14411);
xor U19243 (N_19243,N_14511,N_10283);
xor U19244 (N_19244,N_12022,N_10590);
or U19245 (N_19245,N_10320,N_11744);
or U19246 (N_19246,N_14288,N_14990);
and U19247 (N_19247,N_10522,N_13846);
or U19248 (N_19248,N_13751,N_12835);
nor U19249 (N_19249,N_10830,N_12509);
and U19250 (N_19250,N_13781,N_12358);
or U19251 (N_19251,N_10705,N_13212);
xnor U19252 (N_19252,N_14421,N_11239);
nor U19253 (N_19253,N_10480,N_14925);
xnor U19254 (N_19254,N_13146,N_10451);
xnor U19255 (N_19255,N_12116,N_10631);
nand U19256 (N_19256,N_14083,N_12836);
or U19257 (N_19257,N_14247,N_10341);
nand U19258 (N_19258,N_10235,N_11974);
nor U19259 (N_19259,N_13621,N_11218);
or U19260 (N_19260,N_14260,N_10605);
nor U19261 (N_19261,N_10622,N_13810);
xnor U19262 (N_19262,N_14631,N_11935);
xnor U19263 (N_19263,N_12920,N_12746);
nor U19264 (N_19264,N_11344,N_11141);
nor U19265 (N_19265,N_11513,N_12157);
or U19266 (N_19266,N_13965,N_12664);
and U19267 (N_19267,N_13150,N_11337);
and U19268 (N_19268,N_13391,N_12513);
and U19269 (N_19269,N_13419,N_12995);
xnor U19270 (N_19270,N_10192,N_13771);
nor U19271 (N_19271,N_12764,N_10420);
xnor U19272 (N_19272,N_14130,N_14089);
and U19273 (N_19273,N_14994,N_12426);
nor U19274 (N_19274,N_11914,N_13939);
and U19275 (N_19275,N_12326,N_13131);
or U19276 (N_19276,N_10651,N_11955);
nand U19277 (N_19277,N_13942,N_10158);
nor U19278 (N_19278,N_11992,N_11930);
nand U19279 (N_19279,N_12190,N_14892);
nor U19280 (N_19280,N_13130,N_13787);
nor U19281 (N_19281,N_10766,N_10861);
or U19282 (N_19282,N_14195,N_12241);
xnor U19283 (N_19283,N_11661,N_13076);
or U19284 (N_19284,N_10540,N_10413);
xnor U19285 (N_19285,N_10093,N_11724);
nand U19286 (N_19286,N_10044,N_10576);
or U19287 (N_19287,N_13268,N_10709);
or U19288 (N_19288,N_12147,N_11348);
or U19289 (N_19289,N_12222,N_14425);
xnor U19290 (N_19290,N_12620,N_14599);
or U19291 (N_19291,N_10258,N_13432);
xor U19292 (N_19292,N_14208,N_12328);
nor U19293 (N_19293,N_13317,N_14970);
nand U19294 (N_19294,N_10213,N_10154);
and U19295 (N_19295,N_13150,N_11911);
and U19296 (N_19296,N_10424,N_11053);
nand U19297 (N_19297,N_13725,N_12912);
or U19298 (N_19298,N_14803,N_12933);
nor U19299 (N_19299,N_10966,N_10872);
nor U19300 (N_19300,N_12562,N_10161);
nor U19301 (N_19301,N_10321,N_11927);
nand U19302 (N_19302,N_11126,N_12360);
nand U19303 (N_19303,N_11991,N_14655);
xor U19304 (N_19304,N_11201,N_11323);
nand U19305 (N_19305,N_10262,N_14368);
xnor U19306 (N_19306,N_13207,N_10611);
or U19307 (N_19307,N_11870,N_10951);
or U19308 (N_19308,N_10511,N_13145);
nand U19309 (N_19309,N_12139,N_13047);
and U19310 (N_19310,N_14715,N_10455);
or U19311 (N_19311,N_10969,N_14381);
nor U19312 (N_19312,N_14442,N_14641);
nand U19313 (N_19313,N_10234,N_11429);
and U19314 (N_19314,N_14422,N_14162);
or U19315 (N_19315,N_13626,N_14494);
nand U19316 (N_19316,N_11342,N_12776);
xor U19317 (N_19317,N_14288,N_10662);
nor U19318 (N_19318,N_14982,N_12526);
nor U19319 (N_19319,N_14536,N_11544);
nand U19320 (N_19320,N_13837,N_13284);
or U19321 (N_19321,N_11847,N_14168);
or U19322 (N_19322,N_13507,N_13754);
nand U19323 (N_19323,N_14418,N_13986);
nand U19324 (N_19324,N_12490,N_11603);
and U19325 (N_19325,N_13514,N_10763);
xor U19326 (N_19326,N_14900,N_10998);
xor U19327 (N_19327,N_10684,N_11101);
nor U19328 (N_19328,N_10478,N_14846);
and U19329 (N_19329,N_14779,N_14199);
nand U19330 (N_19330,N_13443,N_14652);
nand U19331 (N_19331,N_14057,N_14112);
nand U19332 (N_19332,N_13810,N_11639);
xnor U19333 (N_19333,N_14870,N_12498);
nand U19334 (N_19334,N_11927,N_13431);
and U19335 (N_19335,N_10236,N_13559);
and U19336 (N_19336,N_12178,N_13418);
nor U19337 (N_19337,N_10482,N_13427);
or U19338 (N_19338,N_11481,N_13340);
nand U19339 (N_19339,N_14344,N_12121);
and U19340 (N_19340,N_12386,N_14287);
xor U19341 (N_19341,N_11788,N_12733);
or U19342 (N_19342,N_13640,N_11564);
and U19343 (N_19343,N_14327,N_10029);
nor U19344 (N_19344,N_12968,N_13764);
xnor U19345 (N_19345,N_10201,N_11647);
or U19346 (N_19346,N_13829,N_12717);
nand U19347 (N_19347,N_12359,N_10043);
nand U19348 (N_19348,N_10267,N_13340);
nand U19349 (N_19349,N_10255,N_13928);
nor U19350 (N_19350,N_14986,N_10572);
nand U19351 (N_19351,N_10462,N_12907);
or U19352 (N_19352,N_14068,N_10874);
and U19353 (N_19353,N_14871,N_10455);
and U19354 (N_19354,N_12412,N_12535);
xor U19355 (N_19355,N_11597,N_10029);
xnor U19356 (N_19356,N_13346,N_10374);
nand U19357 (N_19357,N_13136,N_11094);
xor U19358 (N_19358,N_11685,N_10234);
nor U19359 (N_19359,N_11379,N_12636);
nor U19360 (N_19360,N_14325,N_11475);
and U19361 (N_19361,N_12164,N_13247);
and U19362 (N_19362,N_12779,N_10981);
nor U19363 (N_19363,N_10094,N_14964);
nand U19364 (N_19364,N_10032,N_13634);
xor U19365 (N_19365,N_12942,N_13051);
nand U19366 (N_19366,N_13961,N_13237);
or U19367 (N_19367,N_11349,N_12342);
nor U19368 (N_19368,N_11441,N_11254);
nand U19369 (N_19369,N_10771,N_10103);
nand U19370 (N_19370,N_14906,N_13804);
nand U19371 (N_19371,N_14271,N_11291);
or U19372 (N_19372,N_11388,N_12285);
or U19373 (N_19373,N_11572,N_10384);
nand U19374 (N_19374,N_14796,N_14149);
or U19375 (N_19375,N_14072,N_13780);
xor U19376 (N_19376,N_12120,N_11747);
nand U19377 (N_19377,N_10695,N_10122);
xor U19378 (N_19378,N_10923,N_14170);
xnor U19379 (N_19379,N_11690,N_13953);
nand U19380 (N_19380,N_10058,N_14969);
and U19381 (N_19381,N_10912,N_10163);
xnor U19382 (N_19382,N_11418,N_10990);
and U19383 (N_19383,N_14258,N_10384);
and U19384 (N_19384,N_10282,N_11742);
or U19385 (N_19385,N_12155,N_12225);
xnor U19386 (N_19386,N_14355,N_10997);
nor U19387 (N_19387,N_11346,N_13986);
xnor U19388 (N_19388,N_12984,N_12604);
and U19389 (N_19389,N_13753,N_11254);
nand U19390 (N_19390,N_13813,N_14676);
nand U19391 (N_19391,N_14650,N_10382);
and U19392 (N_19392,N_14043,N_10846);
or U19393 (N_19393,N_12495,N_11035);
nor U19394 (N_19394,N_12358,N_10354);
xor U19395 (N_19395,N_13590,N_13885);
nor U19396 (N_19396,N_10304,N_14085);
or U19397 (N_19397,N_14594,N_11052);
and U19398 (N_19398,N_13305,N_13066);
nor U19399 (N_19399,N_14278,N_10775);
xor U19400 (N_19400,N_10936,N_10968);
and U19401 (N_19401,N_10659,N_11694);
nor U19402 (N_19402,N_13394,N_13702);
or U19403 (N_19403,N_10581,N_14786);
xnor U19404 (N_19404,N_12147,N_10791);
nand U19405 (N_19405,N_10092,N_13142);
and U19406 (N_19406,N_11251,N_11376);
nand U19407 (N_19407,N_12678,N_10966);
nor U19408 (N_19408,N_14959,N_14025);
nand U19409 (N_19409,N_12488,N_11078);
or U19410 (N_19410,N_14766,N_13193);
or U19411 (N_19411,N_12194,N_13248);
and U19412 (N_19412,N_12944,N_14750);
nand U19413 (N_19413,N_14713,N_10981);
nor U19414 (N_19414,N_13583,N_12707);
nand U19415 (N_19415,N_11652,N_11821);
and U19416 (N_19416,N_11284,N_14224);
and U19417 (N_19417,N_10205,N_10152);
xor U19418 (N_19418,N_12200,N_13392);
and U19419 (N_19419,N_12233,N_13686);
and U19420 (N_19420,N_10472,N_10546);
and U19421 (N_19421,N_14641,N_14346);
nand U19422 (N_19422,N_11289,N_14349);
or U19423 (N_19423,N_12562,N_13216);
nand U19424 (N_19424,N_12730,N_13921);
nor U19425 (N_19425,N_13893,N_10814);
xor U19426 (N_19426,N_10142,N_10086);
xor U19427 (N_19427,N_14186,N_11585);
xnor U19428 (N_19428,N_14809,N_12376);
and U19429 (N_19429,N_12144,N_10451);
nand U19430 (N_19430,N_13157,N_12263);
nand U19431 (N_19431,N_11048,N_13246);
nor U19432 (N_19432,N_12596,N_10723);
and U19433 (N_19433,N_14523,N_10494);
xnor U19434 (N_19434,N_14194,N_13947);
xor U19435 (N_19435,N_11995,N_13544);
xnor U19436 (N_19436,N_14269,N_12879);
nor U19437 (N_19437,N_14556,N_12223);
xor U19438 (N_19438,N_14039,N_12564);
nand U19439 (N_19439,N_13408,N_12873);
and U19440 (N_19440,N_12319,N_13787);
or U19441 (N_19441,N_11391,N_11541);
nor U19442 (N_19442,N_13471,N_12905);
or U19443 (N_19443,N_13251,N_13391);
xnor U19444 (N_19444,N_12950,N_11337);
or U19445 (N_19445,N_12238,N_11955);
or U19446 (N_19446,N_12504,N_11810);
nor U19447 (N_19447,N_11234,N_14148);
xor U19448 (N_19448,N_12780,N_11453);
nor U19449 (N_19449,N_13463,N_11557);
xnor U19450 (N_19450,N_12090,N_13884);
or U19451 (N_19451,N_10591,N_14940);
or U19452 (N_19452,N_12824,N_13586);
nor U19453 (N_19453,N_12775,N_10752);
xor U19454 (N_19454,N_14281,N_14944);
or U19455 (N_19455,N_10504,N_11070);
or U19456 (N_19456,N_14898,N_14957);
nor U19457 (N_19457,N_14964,N_13263);
or U19458 (N_19458,N_10888,N_11467);
or U19459 (N_19459,N_11595,N_11518);
or U19460 (N_19460,N_14977,N_13450);
nand U19461 (N_19461,N_11419,N_14747);
and U19462 (N_19462,N_12400,N_12129);
nor U19463 (N_19463,N_14294,N_14281);
xnor U19464 (N_19464,N_13902,N_11750);
nand U19465 (N_19465,N_14964,N_10253);
nor U19466 (N_19466,N_14715,N_14764);
xor U19467 (N_19467,N_10112,N_10467);
nand U19468 (N_19468,N_10364,N_13890);
xor U19469 (N_19469,N_12606,N_12133);
nor U19470 (N_19470,N_11673,N_10605);
nand U19471 (N_19471,N_13888,N_11396);
nor U19472 (N_19472,N_14883,N_12551);
nor U19473 (N_19473,N_14236,N_11067);
nand U19474 (N_19474,N_11111,N_10885);
nor U19475 (N_19475,N_10899,N_10855);
nand U19476 (N_19476,N_12946,N_13757);
or U19477 (N_19477,N_14389,N_13905);
nor U19478 (N_19478,N_13788,N_12083);
xor U19479 (N_19479,N_12979,N_13072);
nor U19480 (N_19480,N_10233,N_13273);
xor U19481 (N_19481,N_12113,N_13140);
and U19482 (N_19482,N_10960,N_10485);
and U19483 (N_19483,N_11029,N_11067);
nor U19484 (N_19484,N_13949,N_10572);
nor U19485 (N_19485,N_14725,N_12773);
nor U19486 (N_19486,N_13041,N_11685);
nand U19487 (N_19487,N_14468,N_13465);
xor U19488 (N_19488,N_12208,N_11316);
and U19489 (N_19489,N_11509,N_10958);
nor U19490 (N_19490,N_12841,N_13251);
and U19491 (N_19491,N_13278,N_12571);
xor U19492 (N_19492,N_11548,N_11569);
or U19493 (N_19493,N_11098,N_11242);
or U19494 (N_19494,N_14975,N_10194);
xor U19495 (N_19495,N_12748,N_14186);
nand U19496 (N_19496,N_12153,N_11952);
or U19497 (N_19497,N_12998,N_14085);
xor U19498 (N_19498,N_12123,N_11669);
xnor U19499 (N_19499,N_12358,N_14469);
or U19500 (N_19500,N_14619,N_14900);
or U19501 (N_19501,N_14068,N_13649);
nand U19502 (N_19502,N_11361,N_12904);
nor U19503 (N_19503,N_10445,N_10941);
and U19504 (N_19504,N_11343,N_14357);
or U19505 (N_19505,N_12220,N_10162);
or U19506 (N_19506,N_13474,N_12201);
xnor U19507 (N_19507,N_14990,N_12634);
or U19508 (N_19508,N_13354,N_11477);
nand U19509 (N_19509,N_13500,N_12482);
nor U19510 (N_19510,N_12954,N_13564);
or U19511 (N_19511,N_13016,N_12051);
and U19512 (N_19512,N_14750,N_11706);
nand U19513 (N_19513,N_10929,N_10626);
or U19514 (N_19514,N_11044,N_10581);
and U19515 (N_19515,N_10229,N_12988);
nor U19516 (N_19516,N_12241,N_14085);
nand U19517 (N_19517,N_10949,N_14652);
nand U19518 (N_19518,N_13087,N_10761);
nor U19519 (N_19519,N_10576,N_11043);
nor U19520 (N_19520,N_11512,N_11905);
or U19521 (N_19521,N_13221,N_13263);
nand U19522 (N_19522,N_13564,N_12551);
and U19523 (N_19523,N_12542,N_14950);
nor U19524 (N_19524,N_14485,N_14912);
or U19525 (N_19525,N_11883,N_12571);
xnor U19526 (N_19526,N_13306,N_12512);
nand U19527 (N_19527,N_14566,N_12928);
nor U19528 (N_19528,N_14272,N_13777);
or U19529 (N_19529,N_13983,N_14303);
and U19530 (N_19530,N_14164,N_13360);
and U19531 (N_19531,N_13628,N_12419);
and U19532 (N_19532,N_13343,N_10882);
and U19533 (N_19533,N_14205,N_11149);
or U19534 (N_19534,N_13646,N_14820);
xnor U19535 (N_19535,N_13504,N_10830);
nor U19536 (N_19536,N_14100,N_13544);
xor U19537 (N_19537,N_14098,N_10431);
xnor U19538 (N_19538,N_13832,N_10394);
nand U19539 (N_19539,N_13153,N_13613);
xor U19540 (N_19540,N_10316,N_10643);
or U19541 (N_19541,N_13597,N_12375);
xnor U19542 (N_19542,N_14860,N_12043);
and U19543 (N_19543,N_13011,N_10162);
and U19544 (N_19544,N_13530,N_11399);
or U19545 (N_19545,N_14703,N_11494);
nand U19546 (N_19546,N_12924,N_11533);
xnor U19547 (N_19547,N_14497,N_13534);
nand U19548 (N_19548,N_11729,N_13762);
and U19549 (N_19549,N_13366,N_10613);
and U19550 (N_19550,N_12762,N_10628);
or U19551 (N_19551,N_10936,N_12852);
xnor U19552 (N_19552,N_14513,N_13020);
or U19553 (N_19553,N_11859,N_13029);
nand U19554 (N_19554,N_13276,N_11742);
xnor U19555 (N_19555,N_14993,N_12652);
nand U19556 (N_19556,N_11252,N_10513);
nand U19557 (N_19557,N_14415,N_13314);
xnor U19558 (N_19558,N_13872,N_12574);
and U19559 (N_19559,N_13848,N_11628);
nand U19560 (N_19560,N_14835,N_14691);
and U19561 (N_19561,N_10008,N_11985);
nor U19562 (N_19562,N_11282,N_12630);
nor U19563 (N_19563,N_10344,N_13930);
xnor U19564 (N_19564,N_10093,N_11765);
and U19565 (N_19565,N_12351,N_10259);
and U19566 (N_19566,N_11502,N_10835);
nor U19567 (N_19567,N_10239,N_12047);
nand U19568 (N_19568,N_12971,N_10051);
nand U19569 (N_19569,N_14006,N_11957);
nor U19570 (N_19570,N_13798,N_10068);
nor U19571 (N_19571,N_11820,N_14529);
nor U19572 (N_19572,N_11459,N_12120);
and U19573 (N_19573,N_10541,N_11927);
xor U19574 (N_19574,N_12436,N_10225);
nor U19575 (N_19575,N_12531,N_11109);
nand U19576 (N_19576,N_12566,N_14531);
nand U19577 (N_19577,N_10676,N_14109);
nor U19578 (N_19578,N_10930,N_14999);
xor U19579 (N_19579,N_10853,N_14896);
or U19580 (N_19580,N_11710,N_14128);
or U19581 (N_19581,N_10814,N_10022);
and U19582 (N_19582,N_10142,N_12531);
and U19583 (N_19583,N_13264,N_12357);
nor U19584 (N_19584,N_10158,N_13491);
and U19585 (N_19585,N_11317,N_14526);
xor U19586 (N_19586,N_10642,N_12498);
nor U19587 (N_19587,N_11721,N_11981);
nor U19588 (N_19588,N_14415,N_10352);
and U19589 (N_19589,N_13054,N_10475);
nor U19590 (N_19590,N_14818,N_10471);
nand U19591 (N_19591,N_14444,N_11240);
xor U19592 (N_19592,N_13593,N_11190);
and U19593 (N_19593,N_13052,N_11330);
nor U19594 (N_19594,N_13676,N_10909);
nor U19595 (N_19595,N_13265,N_13701);
nor U19596 (N_19596,N_13257,N_12388);
or U19597 (N_19597,N_12714,N_11132);
nand U19598 (N_19598,N_14885,N_14550);
nor U19599 (N_19599,N_12053,N_10217);
xor U19600 (N_19600,N_12687,N_13161);
nand U19601 (N_19601,N_12821,N_12696);
xnor U19602 (N_19602,N_11462,N_10365);
nand U19603 (N_19603,N_14264,N_13148);
nor U19604 (N_19604,N_11394,N_11199);
nand U19605 (N_19605,N_14632,N_10050);
nand U19606 (N_19606,N_14314,N_10760);
and U19607 (N_19607,N_12112,N_11339);
xor U19608 (N_19608,N_11086,N_12373);
and U19609 (N_19609,N_10687,N_12900);
nand U19610 (N_19610,N_11342,N_12332);
nor U19611 (N_19611,N_11155,N_13904);
or U19612 (N_19612,N_12380,N_13140);
or U19613 (N_19613,N_14416,N_14304);
or U19614 (N_19614,N_10054,N_14529);
xnor U19615 (N_19615,N_11271,N_14275);
nand U19616 (N_19616,N_12023,N_14045);
or U19617 (N_19617,N_11533,N_12713);
nor U19618 (N_19618,N_10749,N_14680);
nor U19619 (N_19619,N_11103,N_14979);
nand U19620 (N_19620,N_12610,N_10560);
xnor U19621 (N_19621,N_10364,N_12291);
or U19622 (N_19622,N_14962,N_14829);
xnor U19623 (N_19623,N_10079,N_14740);
or U19624 (N_19624,N_11169,N_11656);
nand U19625 (N_19625,N_10930,N_14899);
xor U19626 (N_19626,N_12718,N_10348);
xor U19627 (N_19627,N_10184,N_10956);
xnor U19628 (N_19628,N_10615,N_11319);
xor U19629 (N_19629,N_13297,N_11013);
nor U19630 (N_19630,N_13633,N_13671);
or U19631 (N_19631,N_10194,N_14399);
xor U19632 (N_19632,N_13899,N_14388);
and U19633 (N_19633,N_14832,N_14592);
xor U19634 (N_19634,N_12069,N_11894);
nor U19635 (N_19635,N_13987,N_13949);
or U19636 (N_19636,N_12644,N_13210);
xnor U19637 (N_19637,N_10589,N_13861);
and U19638 (N_19638,N_12607,N_10723);
and U19639 (N_19639,N_13970,N_12575);
and U19640 (N_19640,N_10763,N_14718);
or U19641 (N_19641,N_14855,N_14560);
xnor U19642 (N_19642,N_12734,N_14548);
and U19643 (N_19643,N_11549,N_10840);
and U19644 (N_19644,N_12921,N_13753);
and U19645 (N_19645,N_10610,N_10305);
nor U19646 (N_19646,N_13081,N_10024);
and U19647 (N_19647,N_14435,N_14050);
nor U19648 (N_19648,N_12402,N_13702);
and U19649 (N_19649,N_11624,N_13165);
xnor U19650 (N_19650,N_12471,N_13055);
or U19651 (N_19651,N_10500,N_10570);
nor U19652 (N_19652,N_10304,N_12536);
nor U19653 (N_19653,N_10627,N_12548);
and U19654 (N_19654,N_12539,N_12076);
or U19655 (N_19655,N_12687,N_12957);
xnor U19656 (N_19656,N_13136,N_10492);
nor U19657 (N_19657,N_13348,N_10031);
and U19658 (N_19658,N_14422,N_11830);
nand U19659 (N_19659,N_10402,N_10878);
and U19660 (N_19660,N_10943,N_13048);
nor U19661 (N_19661,N_14459,N_11730);
xor U19662 (N_19662,N_10782,N_11716);
and U19663 (N_19663,N_11061,N_12514);
nand U19664 (N_19664,N_13556,N_11097);
xnor U19665 (N_19665,N_11147,N_10470);
nor U19666 (N_19666,N_12225,N_13522);
and U19667 (N_19667,N_13346,N_11934);
or U19668 (N_19668,N_12770,N_14915);
nor U19669 (N_19669,N_13284,N_11947);
xor U19670 (N_19670,N_13140,N_14785);
nand U19671 (N_19671,N_12130,N_10420);
xor U19672 (N_19672,N_12065,N_12257);
xnor U19673 (N_19673,N_10334,N_13030);
nor U19674 (N_19674,N_12004,N_14015);
xor U19675 (N_19675,N_13476,N_14256);
nor U19676 (N_19676,N_13526,N_10695);
nand U19677 (N_19677,N_10337,N_13290);
xor U19678 (N_19678,N_14441,N_10171);
or U19679 (N_19679,N_13572,N_13532);
or U19680 (N_19680,N_12719,N_12809);
or U19681 (N_19681,N_14209,N_13998);
nor U19682 (N_19682,N_12423,N_11986);
nand U19683 (N_19683,N_14051,N_14515);
nand U19684 (N_19684,N_10379,N_13582);
or U19685 (N_19685,N_13403,N_12478);
or U19686 (N_19686,N_14957,N_10790);
and U19687 (N_19687,N_13359,N_14533);
xor U19688 (N_19688,N_10574,N_14308);
or U19689 (N_19689,N_13066,N_13527);
nor U19690 (N_19690,N_10756,N_14573);
nor U19691 (N_19691,N_12443,N_13524);
nand U19692 (N_19692,N_14701,N_12735);
nor U19693 (N_19693,N_10846,N_12218);
xor U19694 (N_19694,N_13469,N_13408);
nand U19695 (N_19695,N_14653,N_12013);
nor U19696 (N_19696,N_12338,N_10409);
nand U19697 (N_19697,N_14018,N_14957);
nand U19698 (N_19698,N_11426,N_12868);
or U19699 (N_19699,N_10526,N_10532);
nor U19700 (N_19700,N_10924,N_10784);
xnor U19701 (N_19701,N_12009,N_13033);
or U19702 (N_19702,N_13363,N_11580);
nand U19703 (N_19703,N_14477,N_11162);
nand U19704 (N_19704,N_14773,N_13185);
nand U19705 (N_19705,N_11020,N_10287);
and U19706 (N_19706,N_11173,N_11483);
nor U19707 (N_19707,N_12022,N_10797);
nand U19708 (N_19708,N_10147,N_11643);
nand U19709 (N_19709,N_10697,N_13293);
or U19710 (N_19710,N_13032,N_12060);
xor U19711 (N_19711,N_13030,N_13587);
nor U19712 (N_19712,N_14762,N_10271);
nand U19713 (N_19713,N_13810,N_14454);
and U19714 (N_19714,N_12298,N_12599);
and U19715 (N_19715,N_13198,N_10515);
xor U19716 (N_19716,N_11776,N_14679);
nor U19717 (N_19717,N_14739,N_13781);
and U19718 (N_19718,N_11098,N_10390);
nand U19719 (N_19719,N_11771,N_13996);
or U19720 (N_19720,N_11445,N_11912);
or U19721 (N_19721,N_12478,N_10222);
xnor U19722 (N_19722,N_10330,N_12639);
or U19723 (N_19723,N_12834,N_13989);
nor U19724 (N_19724,N_12604,N_11263);
and U19725 (N_19725,N_12202,N_13823);
xnor U19726 (N_19726,N_13986,N_10865);
and U19727 (N_19727,N_10626,N_13373);
nand U19728 (N_19728,N_12519,N_12424);
and U19729 (N_19729,N_14973,N_14437);
nand U19730 (N_19730,N_12464,N_11599);
nand U19731 (N_19731,N_12995,N_11596);
or U19732 (N_19732,N_10722,N_13549);
nand U19733 (N_19733,N_11561,N_13647);
nor U19734 (N_19734,N_10452,N_11880);
and U19735 (N_19735,N_12043,N_10459);
or U19736 (N_19736,N_14564,N_13774);
and U19737 (N_19737,N_13508,N_11097);
and U19738 (N_19738,N_12670,N_10229);
nand U19739 (N_19739,N_11697,N_14754);
xnor U19740 (N_19740,N_14488,N_11288);
and U19741 (N_19741,N_14083,N_11644);
and U19742 (N_19742,N_11055,N_14453);
xor U19743 (N_19743,N_14037,N_12818);
and U19744 (N_19744,N_12189,N_12343);
nor U19745 (N_19745,N_10519,N_11577);
or U19746 (N_19746,N_10186,N_11147);
nor U19747 (N_19747,N_12955,N_14119);
nand U19748 (N_19748,N_10742,N_12682);
nand U19749 (N_19749,N_10267,N_10369);
nand U19750 (N_19750,N_14520,N_10430);
or U19751 (N_19751,N_14510,N_12978);
nand U19752 (N_19752,N_12743,N_12793);
xor U19753 (N_19753,N_10635,N_13818);
or U19754 (N_19754,N_14279,N_14546);
or U19755 (N_19755,N_13515,N_10343);
or U19756 (N_19756,N_10998,N_10775);
and U19757 (N_19757,N_10364,N_14311);
xnor U19758 (N_19758,N_13889,N_14307);
nand U19759 (N_19759,N_14730,N_12008);
nor U19760 (N_19760,N_14764,N_12249);
nor U19761 (N_19761,N_14891,N_13622);
xor U19762 (N_19762,N_11616,N_14027);
nand U19763 (N_19763,N_11862,N_12016);
and U19764 (N_19764,N_14962,N_10893);
and U19765 (N_19765,N_13785,N_10354);
nor U19766 (N_19766,N_14323,N_12072);
nand U19767 (N_19767,N_11173,N_11928);
and U19768 (N_19768,N_11025,N_13704);
and U19769 (N_19769,N_10810,N_13843);
and U19770 (N_19770,N_14429,N_14943);
nor U19771 (N_19771,N_12049,N_13731);
and U19772 (N_19772,N_10305,N_10474);
nor U19773 (N_19773,N_14721,N_14277);
nand U19774 (N_19774,N_10141,N_14621);
nor U19775 (N_19775,N_11063,N_11449);
xnor U19776 (N_19776,N_14902,N_10912);
xnor U19777 (N_19777,N_10994,N_12145);
nand U19778 (N_19778,N_12582,N_13828);
xnor U19779 (N_19779,N_14731,N_11126);
or U19780 (N_19780,N_10805,N_11343);
xnor U19781 (N_19781,N_11802,N_12735);
or U19782 (N_19782,N_12225,N_14289);
or U19783 (N_19783,N_10506,N_11486);
or U19784 (N_19784,N_14295,N_12312);
nor U19785 (N_19785,N_10976,N_12562);
xor U19786 (N_19786,N_14507,N_13820);
xor U19787 (N_19787,N_12906,N_13880);
xnor U19788 (N_19788,N_10774,N_10287);
nand U19789 (N_19789,N_13004,N_11148);
nor U19790 (N_19790,N_13077,N_11260);
or U19791 (N_19791,N_13696,N_14554);
nand U19792 (N_19792,N_10253,N_13352);
nor U19793 (N_19793,N_12157,N_12394);
or U19794 (N_19794,N_13378,N_12761);
or U19795 (N_19795,N_13874,N_14761);
nor U19796 (N_19796,N_11972,N_14478);
xor U19797 (N_19797,N_13517,N_13633);
nor U19798 (N_19798,N_12239,N_10777);
and U19799 (N_19799,N_14972,N_13150);
or U19800 (N_19800,N_14003,N_14880);
and U19801 (N_19801,N_11174,N_14260);
xnor U19802 (N_19802,N_14341,N_13102);
nor U19803 (N_19803,N_11189,N_12740);
or U19804 (N_19804,N_12134,N_13499);
nor U19805 (N_19805,N_12314,N_13099);
nor U19806 (N_19806,N_12174,N_11781);
or U19807 (N_19807,N_12817,N_14348);
xor U19808 (N_19808,N_11290,N_14598);
nand U19809 (N_19809,N_13349,N_11744);
or U19810 (N_19810,N_14317,N_14035);
or U19811 (N_19811,N_11971,N_11340);
xnor U19812 (N_19812,N_13192,N_13654);
and U19813 (N_19813,N_14523,N_11144);
and U19814 (N_19814,N_14806,N_13533);
xnor U19815 (N_19815,N_14891,N_11308);
or U19816 (N_19816,N_14277,N_14593);
or U19817 (N_19817,N_11800,N_13522);
or U19818 (N_19818,N_12339,N_10391);
nand U19819 (N_19819,N_11832,N_13113);
nand U19820 (N_19820,N_11489,N_12732);
or U19821 (N_19821,N_12385,N_14357);
nor U19822 (N_19822,N_10545,N_10602);
and U19823 (N_19823,N_11796,N_11435);
xor U19824 (N_19824,N_11956,N_14972);
or U19825 (N_19825,N_12397,N_12919);
or U19826 (N_19826,N_12284,N_11198);
nor U19827 (N_19827,N_11558,N_12555);
nor U19828 (N_19828,N_12368,N_11435);
and U19829 (N_19829,N_12297,N_12280);
nand U19830 (N_19830,N_13239,N_12209);
nand U19831 (N_19831,N_11436,N_13416);
and U19832 (N_19832,N_14677,N_11745);
nor U19833 (N_19833,N_11048,N_14875);
or U19834 (N_19834,N_13400,N_13649);
xor U19835 (N_19835,N_10325,N_11048);
or U19836 (N_19836,N_11313,N_12993);
xnor U19837 (N_19837,N_14784,N_11932);
or U19838 (N_19838,N_14598,N_13155);
xor U19839 (N_19839,N_13195,N_12172);
xor U19840 (N_19840,N_11359,N_13913);
nor U19841 (N_19841,N_10418,N_10182);
xnor U19842 (N_19842,N_14974,N_11009);
nor U19843 (N_19843,N_12921,N_14694);
and U19844 (N_19844,N_11313,N_11132);
nand U19845 (N_19845,N_10768,N_10776);
or U19846 (N_19846,N_10268,N_12811);
nor U19847 (N_19847,N_14813,N_10989);
nor U19848 (N_19848,N_11824,N_14364);
nor U19849 (N_19849,N_10657,N_10494);
nor U19850 (N_19850,N_13652,N_10816);
nand U19851 (N_19851,N_11739,N_12740);
xor U19852 (N_19852,N_12273,N_11970);
nand U19853 (N_19853,N_14415,N_12313);
nor U19854 (N_19854,N_10614,N_10658);
xnor U19855 (N_19855,N_11132,N_14880);
and U19856 (N_19856,N_11466,N_11977);
nand U19857 (N_19857,N_13703,N_10749);
nand U19858 (N_19858,N_12213,N_12458);
or U19859 (N_19859,N_12663,N_12436);
nor U19860 (N_19860,N_14041,N_10416);
nor U19861 (N_19861,N_10735,N_14733);
or U19862 (N_19862,N_13268,N_10480);
nand U19863 (N_19863,N_12285,N_13000);
nor U19864 (N_19864,N_14200,N_11729);
nor U19865 (N_19865,N_10472,N_13488);
xnor U19866 (N_19866,N_11195,N_14363);
or U19867 (N_19867,N_12251,N_12569);
xor U19868 (N_19868,N_12073,N_12553);
and U19869 (N_19869,N_11672,N_12557);
nor U19870 (N_19870,N_12281,N_11425);
or U19871 (N_19871,N_14279,N_10734);
xor U19872 (N_19872,N_11410,N_10916);
or U19873 (N_19873,N_11247,N_12795);
nand U19874 (N_19874,N_11282,N_10198);
and U19875 (N_19875,N_11784,N_12132);
xor U19876 (N_19876,N_11109,N_10114);
nor U19877 (N_19877,N_12600,N_12605);
nand U19878 (N_19878,N_12538,N_11809);
nand U19879 (N_19879,N_14060,N_10222);
xor U19880 (N_19880,N_14944,N_10831);
or U19881 (N_19881,N_11260,N_13542);
nand U19882 (N_19882,N_13554,N_12553);
or U19883 (N_19883,N_12330,N_10312);
nor U19884 (N_19884,N_11292,N_12290);
and U19885 (N_19885,N_11882,N_13112);
or U19886 (N_19886,N_13067,N_12213);
nor U19887 (N_19887,N_10250,N_14283);
nor U19888 (N_19888,N_10907,N_14763);
and U19889 (N_19889,N_10759,N_13569);
xor U19890 (N_19890,N_13558,N_10208);
xnor U19891 (N_19891,N_13931,N_14808);
xor U19892 (N_19892,N_13193,N_13071);
and U19893 (N_19893,N_14048,N_10214);
nor U19894 (N_19894,N_14862,N_11699);
or U19895 (N_19895,N_14809,N_11895);
or U19896 (N_19896,N_10725,N_10955);
nand U19897 (N_19897,N_12349,N_13813);
and U19898 (N_19898,N_12742,N_12655);
and U19899 (N_19899,N_10155,N_11945);
nor U19900 (N_19900,N_14493,N_14875);
xnor U19901 (N_19901,N_12098,N_12562);
xor U19902 (N_19902,N_14330,N_13714);
nand U19903 (N_19903,N_10679,N_11458);
nor U19904 (N_19904,N_11969,N_14006);
xor U19905 (N_19905,N_12856,N_14886);
and U19906 (N_19906,N_10213,N_10041);
and U19907 (N_19907,N_14501,N_11315);
and U19908 (N_19908,N_10243,N_12656);
or U19909 (N_19909,N_12589,N_14225);
and U19910 (N_19910,N_14878,N_12251);
nand U19911 (N_19911,N_10893,N_11320);
or U19912 (N_19912,N_12162,N_11195);
xnor U19913 (N_19913,N_14060,N_13661);
or U19914 (N_19914,N_12718,N_14017);
and U19915 (N_19915,N_12809,N_11063);
nor U19916 (N_19916,N_11788,N_11638);
nand U19917 (N_19917,N_10291,N_11530);
nor U19918 (N_19918,N_12869,N_11322);
or U19919 (N_19919,N_12514,N_12219);
nor U19920 (N_19920,N_14021,N_12375);
and U19921 (N_19921,N_11812,N_13199);
xnor U19922 (N_19922,N_12946,N_10163);
or U19923 (N_19923,N_12421,N_13816);
or U19924 (N_19924,N_14531,N_10521);
xnor U19925 (N_19925,N_11914,N_12441);
nand U19926 (N_19926,N_12092,N_14689);
and U19927 (N_19927,N_10868,N_11725);
xor U19928 (N_19928,N_12438,N_11524);
nor U19929 (N_19929,N_11737,N_11101);
and U19930 (N_19930,N_11100,N_12993);
or U19931 (N_19931,N_10684,N_13567);
xor U19932 (N_19932,N_14700,N_13582);
nand U19933 (N_19933,N_10376,N_11600);
or U19934 (N_19934,N_14522,N_10004);
and U19935 (N_19935,N_14721,N_10635);
nor U19936 (N_19936,N_13004,N_14585);
or U19937 (N_19937,N_14804,N_10932);
nand U19938 (N_19938,N_14352,N_12018);
or U19939 (N_19939,N_10104,N_12514);
or U19940 (N_19940,N_11982,N_12935);
xor U19941 (N_19941,N_12377,N_13444);
or U19942 (N_19942,N_10032,N_11792);
nand U19943 (N_19943,N_14863,N_13357);
and U19944 (N_19944,N_12695,N_10538);
nand U19945 (N_19945,N_14478,N_11180);
nor U19946 (N_19946,N_14455,N_13756);
or U19947 (N_19947,N_13395,N_14946);
or U19948 (N_19948,N_12128,N_13826);
or U19949 (N_19949,N_11627,N_12567);
and U19950 (N_19950,N_11753,N_14243);
xnor U19951 (N_19951,N_13181,N_13212);
nand U19952 (N_19952,N_12606,N_11331);
or U19953 (N_19953,N_10285,N_11277);
xor U19954 (N_19954,N_10824,N_10357);
and U19955 (N_19955,N_12191,N_14746);
or U19956 (N_19956,N_10061,N_11900);
and U19957 (N_19957,N_11494,N_12606);
xnor U19958 (N_19958,N_13339,N_14199);
nor U19959 (N_19959,N_13484,N_13131);
nor U19960 (N_19960,N_12220,N_12560);
xnor U19961 (N_19961,N_10308,N_11089);
and U19962 (N_19962,N_14121,N_10838);
nor U19963 (N_19963,N_13913,N_13643);
nor U19964 (N_19964,N_14847,N_12110);
or U19965 (N_19965,N_10424,N_13508);
and U19966 (N_19966,N_10875,N_13306);
or U19967 (N_19967,N_11236,N_13066);
nand U19968 (N_19968,N_11672,N_10335);
or U19969 (N_19969,N_11925,N_13957);
or U19970 (N_19970,N_12931,N_14312);
nor U19971 (N_19971,N_13111,N_10620);
xor U19972 (N_19972,N_12281,N_13403);
nor U19973 (N_19973,N_12257,N_12145);
and U19974 (N_19974,N_14887,N_11414);
nor U19975 (N_19975,N_14392,N_12738);
or U19976 (N_19976,N_14668,N_11288);
or U19977 (N_19977,N_13244,N_13428);
xor U19978 (N_19978,N_13683,N_10369);
nor U19979 (N_19979,N_11256,N_10808);
or U19980 (N_19980,N_12259,N_13253);
and U19981 (N_19981,N_10253,N_13058);
nand U19982 (N_19982,N_13577,N_13980);
or U19983 (N_19983,N_14877,N_14514);
nand U19984 (N_19984,N_14694,N_11008);
or U19985 (N_19985,N_12255,N_12175);
nor U19986 (N_19986,N_14434,N_11977);
xnor U19987 (N_19987,N_14531,N_13023);
and U19988 (N_19988,N_13952,N_12734);
or U19989 (N_19989,N_10331,N_10762);
nand U19990 (N_19990,N_14937,N_10598);
and U19991 (N_19991,N_12294,N_10451);
or U19992 (N_19992,N_12480,N_12548);
nand U19993 (N_19993,N_12339,N_14815);
nand U19994 (N_19994,N_13251,N_11105);
and U19995 (N_19995,N_10779,N_14466);
nor U19996 (N_19996,N_11277,N_10122);
xor U19997 (N_19997,N_14007,N_11842);
or U19998 (N_19998,N_11108,N_11905);
and U19999 (N_19999,N_13913,N_11814);
xor U20000 (N_20000,N_18966,N_19935);
nand U20001 (N_20001,N_18705,N_18531);
or U20002 (N_20002,N_18970,N_16738);
xnor U20003 (N_20003,N_18322,N_19154);
nand U20004 (N_20004,N_19027,N_18530);
xor U20005 (N_20005,N_16389,N_19714);
xor U20006 (N_20006,N_17040,N_15418);
nand U20007 (N_20007,N_16461,N_16057);
or U20008 (N_20008,N_17581,N_17488);
nor U20009 (N_20009,N_18428,N_19582);
or U20010 (N_20010,N_19188,N_19800);
or U20011 (N_20011,N_17139,N_18391);
xor U20012 (N_20012,N_17455,N_18919);
nor U20013 (N_20013,N_19259,N_16876);
and U20014 (N_20014,N_18210,N_17265);
xnor U20015 (N_20015,N_17955,N_19491);
xnor U20016 (N_20016,N_16855,N_17737);
and U20017 (N_20017,N_16789,N_16513);
or U20018 (N_20018,N_17428,N_17402);
or U20019 (N_20019,N_16486,N_17697);
nor U20020 (N_20020,N_17365,N_17819);
nor U20021 (N_20021,N_18466,N_15899);
nand U20022 (N_20022,N_15289,N_16028);
nor U20023 (N_20023,N_15006,N_18289);
and U20024 (N_20024,N_15047,N_16573);
nand U20025 (N_20025,N_19065,N_15551);
xor U20026 (N_20026,N_18288,N_16776);
and U20027 (N_20027,N_17325,N_18098);
and U20028 (N_20028,N_16010,N_15986);
or U20029 (N_20029,N_15647,N_19787);
or U20030 (N_20030,N_19945,N_15482);
nor U20031 (N_20031,N_17881,N_17191);
nand U20032 (N_20032,N_17603,N_16372);
and U20033 (N_20033,N_15913,N_16792);
or U20034 (N_20034,N_16033,N_17640);
xor U20035 (N_20035,N_19980,N_16494);
nand U20036 (N_20036,N_18397,N_16426);
or U20037 (N_20037,N_16233,N_17582);
or U20038 (N_20038,N_19432,N_19576);
xnor U20039 (N_20039,N_17649,N_16140);
and U20040 (N_20040,N_17008,N_19323);
or U20041 (N_20041,N_17965,N_18548);
nor U20042 (N_20042,N_18763,N_15275);
nor U20043 (N_20043,N_17193,N_18868);
or U20044 (N_20044,N_15716,N_15245);
nor U20045 (N_20045,N_19485,N_15579);
and U20046 (N_20046,N_16748,N_16048);
or U20047 (N_20047,N_16169,N_16009);
or U20048 (N_20048,N_19626,N_19856);
xor U20049 (N_20049,N_16602,N_17805);
or U20050 (N_20050,N_19351,N_17216);
nand U20051 (N_20051,N_15445,N_18674);
nor U20052 (N_20052,N_15717,N_17849);
or U20053 (N_20053,N_15121,N_19391);
xnor U20054 (N_20054,N_18483,N_17344);
and U20055 (N_20055,N_17412,N_15204);
nor U20056 (N_20056,N_16291,N_18650);
xor U20057 (N_20057,N_15230,N_17751);
and U20058 (N_20058,N_17151,N_18597);
or U20059 (N_20059,N_17645,N_16710);
or U20060 (N_20060,N_17239,N_17076);
nor U20061 (N_20061,N_15709,N_18279);
or U20062 (N_20062,N_17817,N_19831);
xnor U20063 (N_20063,N_15499,N_19046);
nor U20064 (N_20064,N_18685,N_17197);
and U20065 (N_20065,N_18023,N_19052);
xor U20066 (N_20066,N_15998,N_19581);
and U20067 (N_20067,N_19243,N_16990);
and U20068 (N_20068,N_16022,N_18493);
xor U20069 (N_20069,N_19897,N_16301);
xnor U20070 (N_20070,N_15800,N_18091);
xnor U20071 (N_20071,N_16388,N_15648);
or U20072 (N_20072,N_16078,N_18162);
and U20073 (N_20073,N_15955,N_17561);
and U20074 (N_20074,N_15826,N_19462);
nor U20075 (N_20075,N_15026,N_19803);
or U20076 (N_20076,N_17527,N_15992);
nor U20077 (N_20077,N_17142,N_16126);
and U20078 (N_20078,N_18944,N_17163);
xnor U20079 (N_20079,N_17517,N_15078);
nand U20080 (N_20080,N_18753,N_17534);
or U20081 (N_20081,N_16771,N_17258);
nor U20082 (N_20082,N_15233,N_16263);
nand U20083 (N_20083,N_17600,N_17288);
or U20084 (N_20084,N_19449,N_17834);
and U20085 (N_20085,N_18906,N_17631);
xor U20086 (N_20086,N_16836,N_17933);
nor U20087 (N_20087,N_18673,N_15207);
or U20088 (N_20088,N_16911,N_18861);
nand U20089 (N_20089,N_18815,N_19822);
nand U20090 (N_20090,N_18872,N_15691);
and U20091 (N_20091,N_18386,N_17808);
or U20092 (N_20092,N_17146,N_17028);
or U20093 (N_20093,N_17721,N_18143);
or U20094 (N_20094,N_19907,N_16002);
xor U20095 (N_20095,N_18505,N_18224);
and U20096 (N_20096,N_15801,N_15951);
xnor U20097 (N_20097,N_19678,N_15023);
xor U20098 (N_20098,N_19130,N_16042);
nand U20099 (N_20099,N_19878,N_19567);
or U20100 (N_20100,N_18901,N_16407);
and U20101 (N_20101,N_15880,N_15786);
and U20102 (N_20102,N_16757,N_19645);
or U20103 (N_20103,N_19189,N_17642);
and U20104 (N_20104,N_17058,N_15708);
or U20105 (N_20105,N_16989,N_17828);
and U20106 (N_20106,N_18088,N_19434);
nand U20107 (N_20107,N_18636,N_15031);
or U20108 (N_20108,N_15725,N_16487);
or U20109 (N_20109,N_17311,N_17351);
nand U20110 (N_20110,N_16052,N_18940);
nor U20111 (N_20111,N_17702,N_15701);
xnor U20112 (N_20112,N_18606,N_15122);
and U20113 (N_20113,N_19515,N_18672);
xor U20114 (N_20114,N_16974,N_18514);
xor U20115 (N_20115,N_15001,N_18999);
and U20116 (N_20116,N_19041,N_15273);
xnor U20117 (N_20117,N_15156,N_16274);
and U20118 (N_20118,N_17575,N_18507);
nor U20119 (N_20119,N_18778,N_15112);
nand U20120 (N_20120,N_19841,N_16997);
and U20121 (N_20121,N_16802,N_16801);
xnor U20122 (N_20122,N_15768,N_18890);
and U20123 (N_20123,N_15588,N_19635);
nor U20124 (N_20124,N_17323,N_15432);
xor U20125 (N_20125,N_16806,N_19445);
and U20126 (N_20126,N_17067,N_18599);
nand U20127 (N_20127,N_18435,N_16870);
or U20128 (N_20128,N_15858,N_17857);
and U20129 (N_20129,N_15911,N_17446);
nand U20130 (N_20130,N_15485,N_16725);
nor U20131 (N_20131,N_18326,N_19810);
nor U20132 (N_20132,N_17655,N_15796);
nand U20133 (N_20133,N_18173,N_15162);
or U20134 (N_20134,N_16333,N_15412);
and U20135 (N_20135,N_15444,N_15748);
and U20136 (N_20136,N_18692,N_16913);
nor U20137 (N_20137,N_19798,N_19138);
xnor U20138 (N_20138,N_19767,N_18133);
and U20139 (N_20139,N_16168,N_15043);
nand U20140 (N_20140,N_19681,N_15446);
nor U20141 (N_20141,N_18176,N_17803);
and U20142 (N_20142,N_17509,N_19647);
nor U20143 (N_20143,N_19528,N_16276);
or U20144 (N_20144,N_18429,N_19108);
nand U20145 (N_20145,N_15866,N_16373);
nand U20146 (N_20146,N_15956,N_15168);
or U20147 (N_20147,N_18932,N_18184);
xor U20148 (N_20148,N_17059,N_19586);
or U20149 (N_20149,N_15048,N_15931);
nor U20150 (N_20150,N_19532,N_19152);
xnor U20151 (N_20151,N_17261,N_15227);
nand U20152 (N_20152,N_18484,N_16984);
or U20153 (N_20153,N_17962,N_16371);
and U20154 (N_20154,N_16250,N_16516);
nor U20155 (N_20155,N_16442,N_19320);
nor U20156 (N_20156,N_17930,N_16313);
xor U20157 (N_20157,N_15622,N_16204);
and U20158 (N_20158,N_15301,N_18731);
and U20159 (N_20159,N_16081,N_17785);
xor U20160 (N_20160,N_17319,N_18977);
nand U20161 (N_20161,N_15217,N_17681);
or U20162 (N_20162,N_19178,N_18871);
nor U20163 (N_20163,N_18701,N_16348);
nor U20164 (N_20164,N_19461,N_15804);
xnor U20165 (N_20165,N_18961,N_17406);
xor U20166 (N_20166,N_16628,N_15343);
or U20167 (N_20167,N_18528,N_17557);
or U20168 (N_20168,N_17072,N_17868);
and U20169 (N_20169,N_17490,N_15114);
nand U20170 (N_20170,N_18748,N_19623);
xnor U20171 (N_20171,N_17887,N_19964);
and U20172 (N_20172,N_17423,N_16430);
xnor U20173 (N_20173,N_18555,N_17597);
or U20174 (N_20174,N_18051,N_18516);
and U20175 (N_20175,N_17783,N_15824);
nor U20176 (N_20176,N_15010,N_17203);
and U20177 (N_20177,N_16962,N_17861);
or U20178 (N_20178,N_17532,N_19958);
or U20179 (N_20179,N_15274,N_19395);
xnor U20180 (N_20180,N_19683,N_15739);
nor U20181 (N_20181,N_19842,N_15041);
nand U20182 (N_20182,N_19823,N_19079);
xor U20183 (N_20183,N_17284,N_19616);
nand U20184 (N_20184,N_15308,N_17223);
nand U20185 (N_20185,N_19218,N_16330);
or U20186 (N_20186,N_16485,N_17710);
and U20187 (N_20187,N_15562,N_19469);
nand U20188 (N_20188,N_18069,N_15252);
nand U20189 (N_20189,N_17489,N_17668);
nor U20190 (N_20190,N_15350,N_19442);
xnor U20191 (N_20191,N_16857,N_17945);
nor U20192 (N_20192,N_15727,N_15393);
and U20193 (N_20193,N_18120,N_18262);
nor U20194 (N_20194,N_15077,N_16765);
xor U20195 (N_20195,N_15729,N_19246);
nand U20196 (N_20196,N_18877,N_16179);
and U20197 (N_20197,N_15231,N_16594);
or U20198 (N_20198,N_18801,N_17518);
nor U20199 (N_20199,N_18356,N_18405);
nand U20200 (N_20200,N_16899,N_16008);
and U20201 (N_20201,N_17371,N_17741);
nor U20202 (N_20202,N_15565,N_15816);
nor U20203 (N_20203,N_17009,N_16620);
and U20204 (N_20204,N_16116,N_19298);
or U20205 (N_20205,N_19411,N_18300);
nor U20206 (N_20206,N_18792,N_15058);
nor U20207 (N_20207,N_18233,N_19316);
xor U20208 (N_20208,N_19021,N_17304);
or U20209 (N_20209,N_18302,N_16709);
and U20210 (N_20210,N_15247,N_19295);
and U20211 (N_20211,N_15552,N_19436);
nor U20212 (N_20212,N_19342,N_17352);
xor U20213 (N_20213,N_18371,N_15668);
and U20214 (N_20214,N_15554,N_18205);
xor U20215 (N_20215,N_15116,N_17064);
xor U20216 (N_20216,N_16952,N_16150);
nand U20217 (N_20217,N_15578,N_15991);
xnor U20218 (N_20218,N_19742,N_19499);
nor U20219 (N_20219,N_16760,N_17078);
nor U20220 (N_20220,N_15489,N_18547);
xor U20221 (N_20221,N_18255,N_18100);
nand U20222 (N_20222,N_19571,N_15530);
nor U20223 (N_20223,N_15270,N_19450);
and U20224 (N_20224,N_16827,N_15893);
xor U20225 (N_20225,N_18260,N_19826);
nand U20226 (N_20226,N_16540,N_17407);
xor U20227 (N_20227,N_15973,N_19939);
nand U20228 (N_20228,N_15430,N_18177);
nor U20229 (N_20229,N_19900,N_15277);
nor U20230 (N_20230,N_15392,N_16791);
or U20231 (N_20231,N_15345,N_18773);
nor U20232 (N_20232,N_18167,N_17255);
nand U20233 (N_20233,N_19142,N_15170);
nand U20234 (N_20234,N_19049,N_19556);
nor U20235 (N_20235,N_17224,N_17179);
nand U20236 (N_20236,N_18546,N_18592);
and U20237 (N_20237,N_18577,N_18447);
xnor U20238 (N_20238,N_17210,N_19564);
or U20239 (N_20239,N_19853,N_17144);
nor U20240 (N_20240,N_16766,N_15843);
nand U20241 (N_20241,N_18301,N_16156);
nand U20242 (N_20242,N_19083,N_17650);
or U20243 (N_20243,N_16777,N_19638);
and U20244 (N_20244,N_16125,N_17057);
or U20245 (N_20245,N_18159,N_16515);
nor U20246 (N_20246,N_16110,N_17654);
nor U20247 (N_20247,N_15771,N_19572);
xor U20248 (N_20248,N_17373,N_15420);
nor U20249 (N_20249,N_15529,N_17133);
xor U20250 (N_20250,N_16565,N_18989);
nor U20251 (N_20251,N_19477,N_16003);
and U20252 (N_20252,N_18011,N_19655);
nor U20253 (N_20253,N_19700,N_15637);
nor U20254 (N_20254,N_18040,N_17504);
and U20255 (N_20255,N_17718,N_16365);
nand U20256 (N_20256,N_18508,N_15846);
nor U20257 (N_20257,N_17114,N_16079);
xnor U20258 (N_20258,N_15030,N_19080);
and U20259 (N_20259,N_15436,N_16360);
and U20260 (N_20260,N_18353,N_19084);
and U20261 (N_20261,N_18827,N_18061);
xor U20262 (N_20262,N_17062,N_18380);
and U20263 (N_20263,N_16692,N_17674);
and U20264 (N_20264,N_19552,N_18690);
or U20265 (N_20265,N_17979,N_15073);
xnor U20266 (N_20266,N_19871,N_16036);
xnor U20267 (N_20267,N_17036,N_16174);
and U20268 (N_20268,N_15749,N_16070);
xor U20269 (N_20269,N_18244,N_16640);
or U20270 (N_20270,N_16901,N_19796);
or U20271 (N_20271,N_15580,N_18556);
or U20272 (N_20272,N_18525,N_18367);
and U20273 (N_20273,N_17275,N_15198);
xnor U20274 (N_20274,N_15989,N_16794);
xor U20275 (N_20275,N_16999,N_18216);
nand U20276 (N_20276,N_16477,N_18251);
nor U20277 (N_20277,N_19139,N_19962);
and U20278 (N_20278,N_16681,N_19502);
and U20279 (N_20279,N_17259,N_17119);
nor U20280 (N_20280,N_19183,N_17732);
or U20281 (N_20281,N_17380,N_17844);
or U20282 (N_20282,N_16847,N_19899);
xor U20283 (N_20283,N_15616,N_16818);
nand U20284 (N_20284,N_16719,N_15200);
nand U20285 (N_20285,N_17463,N_18523);
or U20286 (N_20286,N_17154,N_15790);
xnor U20287 (N_20287,N_15649,N_18891);
xnor U20288 (N_20288,N_18022,N_17521);
xor U20289 (N_20289,N_19575,N_18575);
or U20290 (N_20290,N_16254,N_19820);
and U20291 (N_20291,N_16304,N_15433);
and U20292 (N_20292,N_17628,N_19210);
and U20293 (N_20293,N_15071,N_18193);
and U20294 (N_20294,N_18443,N_16082);
or U20295 (N_20295,N_16684,N_17770);
nand U20296 (N_20296,N_17010,N_15318);
and U20297 (N_20297,N_17786,N_18954);
or U20298 (N_20298,N_19845,N_17384);
or U20299 (N_20299,N_18654,N_17332);
xnor U20300 (N_20300,N_15226,N_15471);
nand U20301 (N_20301,N_15752,N_18603);
nand U20302 (N_20302,N_16188,N_17956);
xnor U20303 (N_20303,N_17923,N_18348);
nor U20304 (N_20304,N_16068,N_17104);
or U20305 (N_20305,N_16192,N_18459);
and U20306 (N_20306,N_19176,N_18026);
and U20307 (N_20307,N_19309,N_19925);
xor U20308 (N_20308,N_18726,N_15068);
xor U20309 (N_20309,N_19000,N_16665);
xnor U20310 (N_20310,N_16441,N_17924);
nand U20311 (N_20311,N_16144,N_18407);
and U20312 (N_20312,N_18948,N_16664);
nor U20313 (N_20313,N_16538,N_18319);
and U20314 (N_20314,N_19283,N_18121);
and U20315 (N_20315,N_15653,N_15036);
nor U20316 (N_20316,N_17208,N_15635);
nor U20317 (N_20317,N_19091,N_18841);
and U20318 (N_20318,N_15269,N_19979);
nand U20319 (N_20319,N_19550,N_15062);
xnor U20320 (N_20320,N_19337,N_17473);
or U20321 (N_20321,N_18090,N_18250);
and U20322 (N_20322,N_19966,N_16758);
nand U20323 (N_20323,N_18370,N_15435);
nor U20324 (N_20324,N_15428,N_18219);
and U20325 (N_20325,N_19882,N_15259);
xnor U20326 (N_20326,N_18843,N_19943);
nor U20327 (N_20327,N_18141,N_16155);
xnor U20328 (N_20328,N_15621,N_15857);
nand U20329 (N_20329,N_19860,N_15373);
xor U20330 (N_20330,N_16550,N_17321);
or U20331 (N_20331,N_15862,N_18744);
or U20332 (N_20332,N_19716,N_19728);
or U20333 (N_20333,N_16940,N_19663);
nand U20334 (N_20334,N_17699,N_17516);
and U20335 (N_20335,N_17766,N_16811);
or U20336 (N_20336,N_15864,N_18449);
nand U20337 (N_20337,N_15912,N_15572);
and U20338 (N_20338,N_16588,N_19691);
nand U20339 (N_20339,N_16720,N_15777);
nor U20340 (N_20340,N_19611,N_15574);
nand U20341 (N_20341,N_17734,N_17869);
nor U20342 (N_20342,N_15557,N_19741);
or U20343 (N_20343,N_16100,N_19247);
nor U20344 (N_20344,N_19749,N_17775);
xor U20345 (N_20345,N_18057,N_19131);
or U20346 (N_20346,N_17416,N_16105);
xnor U20347 (N_20347,N_16320,N_17269);
and U20348 (N_20348,N_15987,N_19913);
or U20349 (N_20349,N_18777,N_19513);
or U20350 (N_20350,N_16931,N_18333);
nand U20351 (N_20351,N_18089,N_18683);
and U20352 (N_20352,N_16041,N_18315);
nor U20353 (N_20353,N_17888,N_19559);
nor U20354 (N_20354,N_19870,N_18661);
nand U20355 (N_20355,N_18323,N_18096);
nor U20356 (N_20356,N_15287,N_17499);
xor U20357 (N_20357,N_16656,N_19498);
nand U20358 (N_20358,N_18756,N_16231);
or U20359 (N_20359,N_17898,N_15642);
nand U20360 (N_20360,N_18616,N_16267);
xnor U20361 (N_20361,N_17617,N_17462);
and U20362 (N_20362,N_16088,N_15454);
and U20363 (N_20363,N_16701,N_16410);
or U20364 (N_20364,N_15074,N_15549);
or U20365 (N_20365,N_18077,N_18824);
nand U20366 (N_20366,N_18237,N_19356);
nand U20367 (N_20367,N_18381,N_15472);
nand U20368 (N_20368,N_16775,N_19151);
nand U20369 (N_20369,N_17295,N_18852);
xnor U20370 (N_20370,N_19310,N_15497);
nor U20371 (N_20371,N_15886,N_19598);
and U20372 (N_20372,N_15888,N_15920);
or U20373 (N_20373,N_15266,N_16137);
nand U20374 (N_20374,N_18478,N_16842);
or U20375 (N_20375,N_19506,N_18678);
or U20376 (N_20376,N_19030,N_16386);
nand U20377 (N_20377,N_16904,N_16249);
xor U20378 (N_20378,N_19257,N_15850);
xnor U20379 (N_20379,N_17984,N_15205);
nand U20380 (N_20380,N_15902,N_18007);
nand U20381 (N_20381,N_19954,N_19147);
nand U20382 (N_20382,N_17102,N_19880);
nor U20383 (N_20383,N_19426,N_16569);
or U20384 (N_20384,N_16954,N_19270);
xor U20385 (N_20385,N_17878,N_17876);
nand U20386 (N_20386,N_18000,N_19024);
xor U20387 (N_20387,N_19121,N_18625);
nor U20388 (N_20388,N_18737,N_18408);
or U20389 (N_20389,N_18992,N_16727);
xnor U20390 (N_20390,N_17306,N_18836);
and U20391 (N_20391,N_18109,N_17263);
and U20392 (N_20392,N_15610,N_15526);
or U20393 (N_20393,N_19285,N_15743);
nand U20394 (N_20394,N_19170,N_19816);
nand U20395 (N_20395,N_16624,N_18197);
or U20396 (N_20396,N_19441,N_16316);
and U20397 (N_20397,N_19430,N_15615);
and U20398 (N_20398,N_17214,N_16996);
nor U20399 (N_20399,N_16194,N_17985);
nor U20400 (N_20400,N_15629,N_18713);
nor U20401 (N_20401,N_17141,N_15461);
or U20402 (N_20402,N_17272,N_17950);
nand U20403 (N_20403,N_16167,N_16201);
and U20404 (N_20404,N_16359,N_16542);
nand U20405 (N_20405,N_16966,N_18779);
xor U20406 (N_20406,N_16893,N_17156);
nand U20407 (N_20407,N_16302,N_19983);
and U20408 (N_20408,N_16872,N_15921);
and U20409 (N_20409,N_17394,N_16006);
and U20410 (N_20410,N_15720,N_17594);
xor U20411 (N_20411,N_15940,N_16546);
nor U20412 (N_20412,N_16093,N_16211);
or U20413 (N_20413,N_17995,N_16723);
nor U20414 (N_20414,N_17148,N_19135);
xnor U20415 (N_20415,N_16972,N_18915);
xor U20416 (N_20416,N_15819,N_15403);
or U20417 (N_20417,N_18653,N_17914);
and U20418 (N_20418,N_16280,N_18055);
and U20419 (N_20419,N_16180,N_18545);
and U20420 (N_20420,N_15218,N_15066);
nor U20421 (N_20421,N_19199,N_16804);
and U20422 (N_20422,N_19089,N_16136);
or U20423 (N_20423,N_16805,N_17845);
or U20424 (N_20424,N_19007,N_17020);
and U20425 (N_20425,N_15546,N_18814);
or U20426 (N_20426,N_18171,N_18106);
nor U20427 (N_20427,N_18240,N_16733);
and U20428 (N_20428,N_16662,N_15347);
and U20429 (N_20429,N_19833,N_19971);
or U20430 (N_20430,N_19141,N_15685);
nor U20431 (N_20431,N_19403,N_18311);
xnor U20432 (N_20432,N_15969,N_15892);
or U20433 (N_20433,N_19997,N_16654);
nor U20434 (N_20434,N_19225,N_16815);
or U20435 (N_20435,N_16957,N_18107);
and U20436 (N_20436,N_16527,N_17294);
or U20437 (N_20437,N_17940,N_17068);
xnor U20438 (N_20438,N_18870,N_19358);
or U20439 (N_20439,N_15212,N_15038);
xnor U20440 (N_20440,N_19752,N_17978);
or U20441 (N_20441,N_16482,N_15977);
xnor U20442 (N_20442,N_17368,N_17213);
and U20443 (N_20443,N_15400,N_19965);
xor U20444 (N_20444,N_18957,N_18137);
xor U20445 (N_20445,N_18565,N_16338);
nand U20446 (N_20446,N_16571,N_19264);
nor U20447 (N_20447,N_15561,N_15840);
nand U20448 (N_20448,N_17291,N_19305);
nor U20449 (N_20449,N_15271,N_19808);
nor U20450 (N_20450,N_18033,N_16986);
nand U20451 (N_20451,N_15191,N_15640);
nand U20452 (N_20452,N_19720,N_16391);
nor U20453 (N_20453,N_18025,N_19585);
xor U20454 (N_20454,N_18734,N_19789);
nand U20455 (N_20455,N_15522,N_16751);
nor U20456 (N_20456,N_18579,N_18382);
nand U20457 (N_20457,N_16970,N_15811);
nor U20458 (N_20458,N_15478,N_18629);
and U20459 (N_20459,N_18680,N_18303);
nand U20460 (N_20460,N_16369,N_19908);
xor U20461 (N_20461,N_19843,N_18281);
and U20462 (N_20462,N_16920,N_19297);
xnor U20463 (N_20463,N_16086,N_19832);
xnor U20464 (N_20464,N_15481,N_16919);
nor U20465 (N_20465,N_19360,N_15607);
nor U20466 (N_20466,N_18211,N_18959);
nor U20467 (N_20467,N_16623,N_19016);
xnor U20468 (N_20468,N_19874,N_19633);
and U20469 (N_20469,N_18490,N_17338);
or U20470 (N_20470,N_18456,N_17398);
nor U20471 (N_20471,N_19153,N_15448);
and U20472 (N_20472,N_17405,N_19227);
nor U20473 (N_20473,N_18887,N_16305);
or U20474 (N_20474,N_19412,N_17519);
nand U20475 (N_20475,N_15600,N_18770);
xnor U20476 (N_20476,N_15091,N_15002);
xnor U20477 (N_20477,N_18187,N_16816);
and U20478 (N_20478,N_16699,N_17347);
xor U20479 (N_20479,N_16642,N_18807);
xnor U20480 (N_20480,N_17333,N_16525);
nor U20481 (N_20481,N_16015,N_19215);
xnor U20482 (N_20482,N_16852,N_18875);
or U20483 (N_20483,N_17858,N_15841);
nor U20484 (N_20484,N_17494,N_16458);
or U20485 (N_20485,N_16639,N_15715);
xnor U20486 (N_20486,N_19088,N_16722);
xnor U20487 (N_20487,N_15087,N_15390);
nand U20488 (N_20488,N_19666,N_16029);
nand U20489 (N_20489,N_19724,N_18648);
and U20490 (N_20490,N_19888,N_18103);
or U20491 (N_20491,N_15564,N_19828);
and U20492 (N_20492,N_18444,N_15869);
xnor U20493 (N_20493,N_19641,N_18593);
nand U20494 (N_20494,N_18419,N_18434);
nand U20495 (N_20495,N_18046,N_15431);
and U20496 (N_20496,N_15407,N_15721);
xor U20497 (N_20497,N_17081,N_19415);
and U20498 (N_20498,N_17542,N_17041);
nor U20499 (N_20499,N_15742,N_19595);
and U20500 (N_20500,N_18776,N_19797);
and U20501 (N_20501,N_18923,N_15897);
nand U20502 (N_20502,N_15014,N_15963);
xnor U20503 (N_20503,N_15605,N_18709);
or U20504 (N_20504,N_17121,N_18017);
xnor U20505 (N_20505,N_15050,N_15460);
and U20506 (N_20506,N_19982,N_16428);
or U20507 (N_20507,N_16592,N_18842);
or U20508 (N_20508,N_16772,N_17251);
nand U20509 (N_20509,N_17015,N_15238);
xor U20510 (N_20510,N_15086,N_17472);
nor U20511 (N_20511,N_16764,N_18608);
nor U20512 (N_20512,N_19852,N_18212);
or U20513 (N_20513,N_16653,N_18686);
and U20514 (N_20514,N_16942,N_16945);
nor U20515 (N_20515,N_15958,N_17374);
xnor U20516 (N_20516,N_17007,N_16380);
xnor U20517 (N_20517,N_17906,N_17454);
xnor U20518 (N_20518,N_17289,N_19037);
nand U20519 (N_20519,N_17547,N_18415);
or U20520 (N_20520,N_15820,N_19098);
xnor U20521 (N_20521,N_16505,N_16973);
and U20522 (N_20522,N_16495,N_15630);
nor U20523 (N_20523,N_19127,N_17453);
nor U20524 (N_20524,N_19619,N_17591);
nor U20525 (N_20525,N_15596,N_18830);
and U20526 (N_20526,N_15183,N_16387);
or U20527 (N_20527,N_18882,N_15678);
xnor U20528 (N_20528,N_17424,N_18373);
xnor U20529 (N_20529,N_16488,N_18598);
xor U20530 (N_20530,N_18659,N_15335);
xnor U20531 (N_20531,N_19628,N_17774);
xnor U20532 (N_20532,N_17830,N_16552);
nand U20533 (N_20533,N_18232,N_17705);
nor U20534 (N_20534,N_16099,N_15375);
nand U20535 (N_20535,N_15868,N_17128);
nor U20536 (N_20536,N_19369,N_15612);
nor U20537 (N_20537,N_17236,N_19466);
xnor U20538 (N_20538,N_16435,N_17286);
nand U20539 (N_20539,N_17308,N_16399);
or U20540 (N_20540,N_17643,N_18029);
nor U20541 (N_20541,N_15243,N_19695);
or U20542 (N_20542,N_16523,N_16226);
or U20543 (N_20543,N_16512,N_15126);
xnor U20544 (N_20544,N_18905,N_19919);
nand U20545 (N_20545,N_16413,N_17853);
xor U20546 (N_20546,N_17324,N_19409);
or U20547 (N_20547,N_16191,N_17459);
nand U20548 (N_20548,N_18014,N_19396);
nand U20549 (N_20549,N_16454,N_16671);
and U20550 (N_20550,N_16203,N_16547);
xor U20551 (N_20551,N_19128,N_18857);
nand U20552 (N_20552,N_18412,N_19725);
or U20553 (N_20553,N_19140,N_15063);
or U20554 (N_20554,N_19345,N_16184);
nor U20555 (N_20555,N_18041,N_18471);
xnor U20556 (N_20556,N_19187,N_15474);
xor U20557 (N_20557,N_18457,N_15459);
nor U20558 (N_20558,N_17200,N_15541);
xor U20559 (N_20559,N_18195,N_17647);
nor U20560 (N_20560,N_17696,N_15022);
nand U20561 (N_20561,N_18733,N_19493);
and U20562 (N_20562,N_16287,N_18900);
nand U20563 (N_20563,N_16703,N_15759);
nor U20564 (N_20564,N_17465,N_18273);
nand U20565 (N_20565,N_16027,N_15059);
and U20566 (N_20566,N_19267,N_15125);
and U20567 (N_20567,N_18620,N_19458);
nor U20568 (N_20568,N_18742,N_19460);
and U20569 (N_20569,N_19428,N_18045);
nand U20570 (N_20570,N_17172,N_18699);
xnor U20571 (N_20571,N_18066,N_15492);
and U20572 (N_20572,N_17567,N_16189);
xor U20573 (N_20573,N_17619,N_18132);
nor U20574 (N_20574,N_19117,N_16787);
or U20575 (N_20575,N_16511,N_17354);
and U20576 (N_20576,N_15303,N_19544);
or U20577 (N_20577,N_18151,N_15832);
or U20578 (N_20578,N_18499,N_17963);
and U20579 (N_20579,N_16089,N_19650);
or U20580 (N_20580,N_18420,N_15282);
xor U20581 (N_20581,N_17080,N_15543);
nor U20582 (N_20582,N_19811,N_16878);
or U20583 (N_20583,N_15894,N_16694);
and U20584 (N_20584,N_18020,N_17054);
or U20585 (N_20585,N_18446,N_15106);
xor U20586 (N_20586,N_15201,N_19634);
nor U20587 (N_20587,N_17648,N_15763);
xnor U20588 (N_20588,N_15952,N_16746);
xor U20589 (N_20589,N_18622,N_15349);
and U20590 (N_20590,N_17656,N_18986);
or U20591 (N_20591,N_15654,N_19349);
and U20592 (N_20592,N_15092,N_18067);
and U20593 (N_20593,N_15593,N_17486);
xor U20594 (N_20594,N_18280,N_17113);
or U20595 (N_20595,N_18506,N_15939);
xor U20596 (N_20596,N_19100,N_17181);
nor U20597 (N_20597,N_18052,N_15249);
or U20598 (N_20598,N_18395,N_17124);
nand U20599 (N_20599,N_18413,N_19547);
nor U20600 (N_20600,N_17753,N_15555);
nor U20601 (N_20601,N_18313,N_18527);
and U20602 (N_20602,N_17037,N_19468);
xnor U20603 (N_20603,N_17658,N_16652);
and U20604 (N_20604,N_19781,N_16270);
or U20605 (N_20605,N_18349,N_17262);
nand U20606 (N_20606,N_15663,N_18533);
or U20607 (N_20607,N_17411,N_18762);
and U20608 (N_20608,N_19865,N_16798);
or U20609 (N_20609,N_16142,N_19085);
nand U20610 (N_20610,N_17934,N_19448);
nor U20611 (N_20611,N_16172,N_16631);
and U20612 (N_20612,N_16881,N_15406);
nor U20613 (N_20613,N_16161,N_18520);
or U20614 (N_20614,N_16659,N_17350);
nand U20615 (N_20615,N_17118,N_17168);
nand U20616 (N_20616,N_17801,N_19368);
nor U20617 (N_20617,N_16411,N_16856);
and U20618 (N_20618,N_18488,N_15419);
or U20619 (N_20619,N_17856,N_19622);
or U20620 (N_20620,N_19289,N_17233);
and U20621 (N_20621,N_16232,N_17093);
or U20622 (N_20622,N_19330,N_16377);
and U20623 (N_20623,N_15000,N_17138);
nor U20624 (N_20624,N_15040,N_16091);
nand U20625 (N_20625,N_19413,N_18760);
or U20626 (N_20626,N_19698,N_18626);
or U20627 (N_20627,N_17568,N_17867);
and U20628 (N_20628,N_17616,N_17725);
and U20629 (N_20629,N_19408,N_17541);
or U20630 (N_20630,N_15380,N_16017);
nand U20631 (N_20631,N_16560,N_15339);
xor U20632 (N_20632,N_16129,N_15571);
nor U20633 (N_20633,N_16539,N_16831);
and U20634 (N_20634,N_17740,N_18788);
and U20635 (N_20635,N_17387,N_17162);
and U20636 (N_20636,N_17006,N_16480);
nand U20637 (N_20637,N_16734,N_16311);
or U20638 (N_20638,N_17578,N_18750);
xnor U20639 (N_20639,N_15450,N_17971);
nand U20640 (N_20640,N_17480,N_18147);
xnor U20641 (N_20641,N_15757,N_16382);
or U20642 (N_20642,N_17637,N_19381);
nand U20643 (N_20643,N_18751,N_15936);
nor U20644 (N_20644,N_17614,N_19023);
xor U20645 (N_20645,N_18127,N_18059);
or U20646 (N_20646,N_16223,N_19745);
nor U20647 (N_20647,N_16324,N_18271);
and U20648 (N_20648,N_15664,N_18365);
nand U20649 (N_20649,N_19347,N_18249);
or U20650 (N_20650,N_15325,N_17027);
nor U20651 (N_20651,N_19209,N_16219);
xnor U20652 (N_20652,N_17862,N_17508);
and U20653 (N_20653,N_19244,N_16401);
or U20654 (N_20654,N_16063,N_18738);
nand U20655 (N_20655,N_18951,N_17196);
nor U20656 (N_20656,N_17131,N_16222);
nor U20657 (N_20657,N_15705,N_16510);
nand U20658 (N_20658,N_18696,N_15918);
or U20659 (N_20659,N_19542,N_15128);
nand U20660 (N_20660,N_18234,N_17624);
or U20661 (N_20661,N_19315,N_16178);
xnor U20662 (N_20662,N_19159,N_19352);
and U20663 (N_20663,N_18491,N_18933);
and U20664 (N_20664,N_18352,N_15814);
nor U20665 (N_20665,N_15883,N_19001);
and U20666 (N_20666,N_16529,N_15139);
nand U20667 (N_20667,N_16625,N_16793);
and U20668 (N_20668,N_16567,N_19988);
and U20669 (N_20669,N_17890,N_15263);
and U20670 (N_20670,N_18053,N_19521);
nor U20671 (N_20671,N_19050,N_16185);
nand U20672 (N_20672,N_17874,N_15098);
xnor U20673 (N_20673,N_15427,N_19198);
xor U20674 (N_20674,N_19706,N_15724);
and U20675 (N_20675,N_15861,N_15525);
and U20676 (N_20676,N_15927,N_16995);
or U20677 (N_20677,N_15660,N_17417);
nor U20678 (N_20678,N_15833,N_16367);
nor U20679 (N_20679,N_18013,N_16374);
or U20680 (N_20680,N_16630,N_19812);
nand U20681 (N_20681,N_16603,N_15358);
xnor U20682 (N_20682,N_16312,N_18337);
nor U20683 (N_20683,N_18377,N_19019);
xnor U20684 (N_20684,N_16200,N_16306);
nand U20685 (N_20685,N_17401,N_19656);
nand U20686 (N_20686,N_18498,N_19605);
xor U20687 (N_20687,N_18904,N_18924);
xor U20688 (N_20688,N_16648,N_16612);
nor U20689 (N_20689,N_19119,N_17377);
or U20690 (N_20690,N_16916,N_19268);
nand U20691 (N_20691,N_15094,N_17241);
nand U20692 (N_20692,N_17797,N_17349);
and U20693 (N_20693,N_17155,N_15542);
xor U20694 (N_20694,N_19554,N_19032);
and U20695 (N_20695,N_16107,N_17866);
and U20696 (N_20696,N_17717,N_18359);
and U20697 (N_20697,N_15703,N_15634);
and U20698 (N_20698,N_18142,N_19094);
or U20699 (N_20699,N_17821,N_16884);
nor U20700 (N_20700,N_17065,N_16729);
or U20701 (N_20701,N_19902,N_18470);
nor U20702 (N_20702,N_18829,N_19416);
and U20703 (N_20703,N_19012,N_15049);
xnor U20704 (N_20704,N_18797,N_17225);
nand U20705 (N_20705,N_15783,N_16240);
nor U20706 (N_20706,N_17073,N_17884);
and U20707 (N_20707,N_19516,N_16607);
nor U20708 (N_20708,N_16046,N_16507);
nor U20709 (N_20709,N_16742,N_17314);
and U20710 (N_20710,N_15794,N_19389);
nor U20711 (N_20711,N_15192,N_15328);
and U20712 (N_20712,N_18287,N_17249);
or U20713 (N_20713,N_18393,N_16902);
nand U20714 (N_20714,N_19558,N_18336);
nand U20715 (N_20715,N_16000,N_17436);
nand U20716 (N_20716,N_19770,N_15377);
or U20717 (N_20717,N_16393,N_15680);
nand U20718 (N_20718,N_17590,N_17999);
nand U20719 (N_20719,N_16948,N_17184);
nand U20720 (N_20720,N_16544,N_17871);
nor U20721 (N_20721,N_18647,N_15401);
nand U20722 (N_20722,N_18152,N_16903);
nor U20723 (N_20723,N_17461,N_18328);
xor U20724 (N_20724,N_15521,N_19562);
or U20725 (N_20725,N_19115,N_17936);
nor U20726 (N_20726,N_16698,N_18724);
or U20727 (N_20727,N_16964,N_17784);
and U20728 (N_20728,N_17554,N_18085);
xnor U20729 (N_20729,N_17571,N_19960);
xor U20730 (N_20730,N_19492,N_17611);
nand U20731 (N_20731,N_18087,N_19518);
or U20732 (N_20732,N_19082,N_16745);
and U20733 (N_20733,N_17832,N_18317);
nand U20734 (N_20734,N_16492,N_18740);
and U20735 (N_20735,N_15776,N_19150);
nor U20736 (N_20736,N_15699,N_15239);
xor U20737 (N_20737,N_16460,N_18099);
or U20738 (N_20738,N_19040,N_17620);
and U20739 (N_20739,N_18855,N_19167);
nor U20740 (N_20740,N_18097,N_18795);
or U20741 (N_20741,N_18809,N_17110);
nor U20742 (N_20742,N_15834,N_16897);
or U20743 (N_20743,N_17629,N_18895);
nand U20744 (N_20744,N_15173,N_18312);
nor U20745 (N_20745,N_17904,N_16784);
xnor U20746 (N_20746,N_16930,N_19419);
or U20747 (N_20747,N_18819,N_16173);
and U20748 (N_20748,N_19214,N_15337);
nand U20749 (N_20749,N_18144,N_17279);
nor U20750 (N_20750,N_18853,N_18004);
and U20751 (N_20751,N_17892,N_18082);
nand U20752 (N_20752,N_17548,N_15261);
or U20753 (N_20753,N_17572,N_16900);
xnor U20754 (N_20754,N_16982,N_19095);
nor U20755 (N_20755,N_16596,N_18166);
nor U20756 (N_20756,N_19517,N_15639);
nand U20757 (N_20757,N_16743,N_15550);
and U20758 (N_20758,N_15935,N_17724);
or U20759 (N_20759,N_19677,N_18884);
nor U20760 (N_20760,N_16715,N_16697);
or U20761 (N_20761,N_18453,N_15851);
nand U20762 (N_20762,N_15842,N_18802);
xor U20763 (N_20763,N_19290,N_17589);
or U20764 (N_20764,N_18492,N_18942);
or U20765 (N_20765,N_17176,N_15576);
nand U20766 (N_20766,N_16520,N_19280);
or U20767 (N_20767,N_15661,N_16266);
or U20768 (N_20768,N_17451,N_19066);
and U20769 (N_20769,N_15193,N_16824);
nand U20770 (N_20770,N_17790,N_16318);
xnor U20771 (N_20771,N_19744,N_19956);
nand U20772 (N_20772,N_16785,N_17939);
and U20773 (N_20773,N_19560,N_17713);
or U20774 (N_20774,N_17209,N_15132);
and U20775 (N_20775,N_17467,N_15734);
nor U20776 (N_20776,N_19463,N_16670);
xnor U20777 (N_20777,N_15467,N_18582);
and U20778 (N_20778,N_18800,N_19792);
or U20779 (N_20779,N_18411,N_16094);
nor U20780 (N_20780,N_18921,N_19715);
or U20781 (N_20781,N_19437,N_16627);
nand U20782 (N_20782,N_19439,N_17493);
nand U20783 (N_20783,N_17055,N_16679);
nor U20784 (N_20784,N_15961,N_19388);
or U20785 (N_20785,N_15147,N_17949);
nor U20786 (N_20786,N_16217,N_18345);
xor U20787 (N_20787,N_15582,N_16605);
and U20788 (N_20788,N_18104,N_17458);
and U20789 (N_20789,N_15683,N_17528);
or U20790 (N_20790,N_19407,N_19004);
and U20791 (N_20791,N_18110,N_19579);
or U20792 (N_20792,N_15255,N_15625);
or U20793 (N_20793,N_18965,N_16535);
and U20794 (N_20794,N_16644,N_17254);
nand U20795 (N_20795,N_17372,N_15606);
xor U20796 (N_20796,N_18140,N_18558);
nand U20797 (N_20797,N_16319,N_15302);
or U20798 (N_20798,N_18161,N_19487);
xor U20799 (N_20799,N_18148,N_16066);
nor U20800 (N_20800,N_16894,N_16873);
nand U20801 (N_20801,N_17188,N_19531);
nand U20802 (N_20802,N_19926,N_19456);
nor U20803 (N_20803,N_19950,N_18644);
or U20804 (N_20804,N_19423,N_18422);
and U20805 (N_20805,N_18560,N_15415);
or U20806 (N_20806,N_17382,N_17413);
or U20807 (N_20807,N_18213,N_15476);
and U20808 (N_20808,N_18850,N_18223);
and U20809 (N_20809,N_19508,N_19659);
xor U20810 (N_20810,N_18771,N_15926);
or U20811 (N_20811,N_17870,N_15370);
nand U20812 (N_20812,N_16361,N_16221);
and U20813 (N_20813,N_15410,N_19671);
xnor U20814 (N_20814,N_15229,N_15315);
and U20815 (N_20815,N_16418,N_15441);
and U20816 (N_20816,N_19105,N_15587);
and U20817 (N_20817,N_17608,N_18346);
nor U20818 (N_20818,N_15632,N_19022);
or U20819 (N_20819,N_17891,N_16165);
and U20820 (N_20820,N_17271,N_19390);
or U20821 (N_20821,N_16337,N_18509);
nor U20822 (N_20822,N_17738,N_19318);
or U20823 (N_20823,N_18390,N_15740);
xnor U20824 (N_20824,N_19705,N_19510);
or U20825 (N_20825,N_19203,N_19251);
nand U20826 (N_20826,N_17315,N_17752);
nor U20827 (N_20827,N_17185,N_19081);
or U20828 (N_20828,N_18455,N_18826);
nor U20829 (N_20829,N_15965,N_19265);
xnor U20830 (N_20830,N_16728,N_15037);
or U20831 (N_20831,N_19589,N_16634);
nor U20832 (N_20832,N_15506,N_17492);
xor U20833 (N_20833,N_17404,N_17160);
nand U20834 (N_20834,N_17511,N_17127);
xnor U20835 (N_20835,N_16518,N_17538);
nand U20836 (N_20836,N_18278,N_15590);
nor U20837 (N_20837,N_16693,N_19539);
xnor U20838 (N_20838,N_19735,N_15626);
xnor U20839 (N_20839,N_19930,N_18697);
nor U20840 (N_20840,N_18416,N_18112);
and U20841 (N_20841,N_15344,N_15399);
xnor U20842 (N_20842,N_16153,N_18621);
and U20843 (N_20843,N_17049,N_15187);
nand U20844 (N_20844,N_19104,N_15528);
or U20845 (N_20845,N_19867,N_15075);
nor U20846 (N_20846,N_19630,N_16121);
xor U20847 (N_20847,N_18886,N_17231);
nor U20848 (N_20848,N_16868,N_17242);
xnor U20849 (N_20849,N_17750,N_15437);
nor U20850 (N_20850,N_19162,N_19754);
xnor U20851 (N_20851,N_15028,N_17840);
nor U20852 (N_20852,N_18463,N_15095);
xor U20853 (N_20853,N_18818,N_19624);
or U20854 (N_20854,N_18703,N_17348);
nor U20855 (N_20855,N_19292,N_15129);
or U20856 (N_20856,N_16673,N_15638);
nor U20857 (N_20857,N_17107,N_16967);
and U20858 (N_20858,N_17375,N_18248);
and U20859 (N_20859,N_15473,N_17046);
and U20860 (N_20860,N_15744,N_15948);
and U20861 (N_20861,N_15932,N_19794);
and U20862 (N_20862,N_18720,N_16352);
nor U20863 (N_20863,N_15949,N_18409);
and U20864 (N_20864,N_19934,N_16170);
nor U20865 (N_20865,N_16427,N_18305);
nand U20866 (N_20866,N_18048,N_16479);
nor U20867 (N_20867,N_18247,N_18375);
nand U20868 (N_20868,N_17960,N_18786);
nor U20869 (N_20869,N_19399,N_17432);
nand U20870 (N_20870,N_15117,N_17017);
nor U20871 (N_20871,N_16340,N_15177);
or U20872 (N_20872,N_18392,N_18270);
and U20873 (N_20873,N_18072,N_17426);
or U20874 (N_20874,N_18076,N_18030);
xnor U20875 (N_20875,N_17709,N_15158);
nor U20876 (N_20876,N_19604,N_17550);
nor U20877 (N_20877,N_18657,N_15656);
xnor U20878 (N_20878,N_18687,N_19375);
nor U20879 (N_20879,N_17806,N_16356);
and U20880 (N_20880,N_19599,N_18172);
or U20881 (N_20881,N_16574,N_19464);
or U20882 (N_20882,N_17482,N_15508);
and U20883 (N_20883,N_17171,N_17908);
or U20884 (N_20884,N_18716,N_19760);
or U20885 (N_20885,N_16322,N_16832);
nor U20886 (N_20886,N_17665,N_17238);
and U20887 (N_20887,N_19143,N_17747);
nor U20888 (N_20888,N_16841,N_17873);
nor U20889 (N_20889,N_17651,N_19359);
xor U20890 (N_20890,N_19850,N_17563);
or U20891 (N_20891,N_16444,N_19157);
and U20892 (N_20892,N_17688,N_19869);
nor U20893 (N_20893,N_17274,N_16187);
nor U20894 (N_20894,N_15859,N_19113);
or U20895 (N_20895,N_19782,N_15876);
xor U20896 (N_20896,N_18102,N_15686);
and U20897 (N_20897,N_18781,N_17612);
and U20898 (N_20898,N_17503,N_18922);
and U20899 (N_20899,N_18203,N_18298);
nand U20900 (N_20900,N_19228,N_15310);
or U20901 (N_20901,N_18980,N_16016);
or U20902 (N_20902,N_16317,N_17673);
nor U20903 (N_20903,N_19306,N_17749);
xor U20904 (N_20904,N_19042,N_17599);
or U20905 (N_20905,N_18794,N_16877);
nand U20906 (N_20906,N_19174,N_19169);
xor U20907 (N_20907,N_18261,N_17048);
or U20908 (N_20908,N_15887,N_15879);
nor U20909 (N_20909,N_19989,N_17700);
nand U20910 (N_20910,N_16106,N_16943);
nand U20911 (N_20911,N_18438,N_18486);
and U20912 (N_20912,N_15628,N_15097);
or U20913 (N_20913,N_15990,N_19103);
nor U20914 (N_20914,N_18745,N_18854);
or U20915 (N_20915,N_17230,N_16151);
nor U20916 (N_20916,N_15778,N_15465);
or U20917 (N_20917,N_15142,N_18651);
and U20918 (N_20918,N_18441,N_19718);
or U20919 (N_20919,N_18008,N_15799);
nand U20920 (N_20920,N_15051,N_18156);
and U20921 (N_20921,N_15483,N_19204);
or U20922 (N_20922,N_17693,N_17022);
and U20923 (N_20923,N_18618,N_18757);
nor U20924 (N_20924,N_16905,N_15426);
or U20925 (N_20925,N_18879,N_19249);
and U20926 (N_20926,N_17644,N_16095);
nand U20927 (N_20927,N_19474,N_15875);
nand U20928 (N_20928,N_15280,N_15925);
nor U20929 (N_20929,N_19438,N_17434);
and U20930 (N_20930,N_19981,N_17053);
or U20931 (N_20931,N_19522,N_19005);
nor U20932 (N_20932,N_19778,N_19566);
nor U20933 (N_20933,N_17147,N_16845);
or U20934 (N_20934,N_19577,N_17893);
and U20935 (N_20935,N_16023,N_16175);
or U20936 (N_20936,N_18594,N_16750);
or U20937 (N_20937,N_17419,N_18532);
nand U20938 (N_20938,N_19481,N_19786);
or U20939 (N_20939,N_19281,N_18314);
and U20940 (N_20940,N_16782,N_18682);
nand U20941 (N_20941,N_18955,N_19693);
or U20942 (N_20942,N_17952,N_17475);
xor U20943 (N_20943,N_16666,N_15755);
xor U20944 (N_20944,N_17301,N_18268);
nor U20945 (N_20945,N_17514,N_18623);
xor U20946 (N_20946,N_16347,N_15567);
nor U20947 (N_20947,N_15539,N_17549);
xor U20948 (N_20948,N_18136,N_19020);
xnor U20949 (N_20949,N_18206,N_15439);
and U20950 (N_20950,N_15466,N_16837);
xor U20951 (N_20951,N_18892,N_16880);
and U20952 (N_20952,N_18908,N_16257);
xor U20953 (N_20953,N_18368,N_17595);
or U20954 (N_20954,N_15722,N_17260);
nand U20955 (N_20955,N_17659,N_19201);
and U20956 (N_20956,N_16385,N_19961);
nand U20957 (N_20957,N_16553,N_18743);
xnor U20958 (N_20958,N_17677,N_18318);
nor U20959 (N_20959,N_15486,N_18503);
xnor U20960 (N_20960,N_15414,N_18808);
xnor U20961 (N_20961,N_15353,N_18677);
nor U20962 (N_20962,N_18619,N_17621);
xor U20963 (N_20963,N_17735,N_18765);
and U20964 (N_20964,N_17992,N_19340);
or U20965 (N_20965,N_15443,N_17754);
or U20966 (N_20966,N_16524,N_16436);
or U20967 (N_20967,N_19686,N_18675);
xnor U20968 (N_20968,N_19300,N_18982);
and U20969 (N_20969,N_16706,N_16947);
or U20970 (N_20970,N_16282,N_15135);
and U20971 (N_20971,N_16083,N_17303);
or U20972 (N_20972,N_17842,N_16193);
or U20973 (N_20973,N_15311,N_16230);
and U20974 (N_20974,N_19207,N_16020);
and U20975 (N_20975,N_15495,N_19252);
and U20976 (N_20976,N_19615,N_17177);
and U20977 (N_20977,N_15671,N_16463);
nor U20978 (N_20978,N_18153,N_15681);
nor U20979 (N_20979,N_15954,N_19387);
and U20980 (N_20980,N_15171,N_18388);
nor U20981 (N_20981,N_16958,N_18929);
or U20982 (N_20982,N_16190,N_19986);
nor U20983 (N_20983,N_18844,N_16166);
or U20984 (N_20984,N_17399,N_18976);
and U20985 (N_20985,N_17646,N_17477);
nor U20986 (N_20986,N_16481,N_16408);
nand U20987 (N_20987,N_17000,N_19866);
xor U20988 (N_20988,N_17932,N_16344);
nand U20989 (N_20989,N_17760,N_19465);
nand U20990 (N_20990,N_18003,N_19271);
xor U20991 (N_20991,N_18914,N_16355);
nand U20992 (N_20992,N_16724,N_17126);
nand U20993 (N_20993,N_17798,N_17758);
or U20994 (N_20994,N_18722,N_16981);
nor U20995 (N_20995,N_16491,N_19932);
nor U20996 (N_20996,N_17520,N_18174);
nor U20997 (N_20997,N_15257,N_16786);
or U20998 (N_20998,N_16493,N_19534);
xnor U20999 (N_20999,N_16049,N_16879);
nand U21000 (N_21000,N_19905,N_19064);
or U21001 (N_21001,N_16227,N_17327);
and U21002 (N_21002,N_19353,N_15160);
nor U21003 (N_21003,N_18535,N_19895);
or U21004 (N_21004,N_17004,N_18747);
xnor U21005 (N_21005,N_17746,N_16617);
and U21006 (N_21006,N_17256,N_16783);
xor U21007 (N_21007,N_18079,N_15007);
and U21008 (N_21008,N_16278,N_16849);
and U21009 (N_21009,N_15244,N_16103);
or U21010 (N_21010,N_17035,N_16269);
xor U21011 (N_21011,N_17320,N_19854);
and U21012 (N_21012,N_16045,N_19922);
xor U21013 (N_21013,N_15181,N_18376);
nand U21014 (N_21014,N_19111,N_18406);
nand U21015 (N_21015,N_18343,N_16604);
nand U21016 (N_21016,N_19984,N_16127);
xnor U21017 (N_21017,N_15570,N_15294);
nor U21018 (N_21018,N_16047,N_15942);
or U21019 (N_21019,N_17676,N_19957);
or U21020 (N_21020,N_16563,N_19723);
nor U21021 (N_21021,N_15644,N_17358);
nand U21022 (N_21022,N_15930,N_17183);
or U21023 (N_21023,N_17698,N_18202);
and U21024 (N_21024,N_18611,N_19479);
nand U21025 (N_21025,N_19998,N_16713);
nand U21026 (N_21026,N_15613,N_17356);
nor U21027 (N_21027,N_18344,N_19543);
or U21028 (N_21028,N_16414,N_18693);
and U21029 (N_21029,N_16076,N_18073);
xor U21030 (N_21030,N_19171,N_18718);
and U21031 (N_21031,N_19195,N_16885);
nand U21032 (N_21032,N_16753,N_16985);
or U21033 (N_21033,N_17807,N_16978);
nor U21034 (N_21034,N_18974,N_19992);
nand U21035 (N_21035,N_15830,N_16064);
nor U21036 (N_21036,N_18283,N_18054);
nor U21037 (N_21037,N_18646,N_15793);
or U21038 (N_21038,N_19825,N_17880);
and U21039 (N_21039,N_16014,N_16497);
xnor U21040 (N_21040,N_16363,N_19737);
and U21041 (N_21041,N_19653,N_19751);
or U21042 (N_21042,N_19612,N_15268);
and U21043 (N_21043,N_18780,N_18676);
xor U21044 (N_21044,N_19758,N_16925);
nor U21045 (N_21045,N_17533,N_15583);
or U21046 (N_21046,N_17778,N_17085);
nand U21047 (N_21047,N_18927,N_17357);
nor U21048 (N_21048,N_18190,N_16858);
nand U21049 (N_21049,N_18403,N_16433);
xnor U21050 (N_21050,N_17189,N_18930);
or U21051 (N_21051,N_17167,N_17994);
xnor U21052 (N_21052,N_18960,N_19649);
nand U21053 (N_21053,N_18774,N_19851);
or U21054 (N_21054,N_18361,N_16077);
nand U21055 (N_21055,N_15545,N_19837);
xnor U21056 (N_21056,N_19540,N_15712);
and U21057 (N_21057,N_18038,N_15559);
and U21058 (N_21058,N_18481,N_17622);
nand U21059 (N_21059,N_15100,N_16195);
nand U21060 (N_21060,N_16019,N_18201);
or U21061 (N_21061,N_19048,N_18083);
or U21062 (N_21062,N_16440,N_19688);
and U21063 (N_21063,N_15566,N_15844);
or U21064 (N_21064,N_17777,N_15974);
or U21065 (N_21065,N_15127,N_17001);
nor U21066 (N_21066,N_19561,N_16462);
nand U21067 (N_21067,N_16061,N_16130);
nor U21068 (N_21068,N_15396,N_17313);
or U21069 (N_21069,N_16961,N_18274);
nand U21070 (N_21070,N_18064,N_16038);
and U21071 (N_21071,N_17235,N_15042);
and U21072 (N_21072,N_16788,N_18943);
and U21073 (N_21073,N_18383,N_19158);
and U21074 (N_21074,N_17297,N_18320);
nand U21075 (N_21075,N_17701,N_17011);
or U21076 (N_21076,N_19805,N_15995);
nor U21077 (N_21077,N_18741,N_18462);
nor U21078 (N_21078,N_16424,N_19043);
and U21079 (N_21079,N_17283,N_19166);
and U21080 (N_21080,N_17414,N_19321);
nor U21081 (N_21081,N_16358,N_18464);
nand U21082 (N_21082,N_16026,N_15631);
or U21083 (N_21083,N_19422,N_15067);
nor U21084 (N_21084,N_16867,N_16271);
nand U21085 (N_21085,N_18431,N_18034);
nor U21086 (N_21086,N_19636,N_15975);
xor U21087 (N_21087,N_19658,N_19975);
xor U21088 (N_21088,N_17421,N_19132);
or U21089 (N_21089,N_17137,N_17298);
nand U21090 (N_21090,N_15359,N_15457);
and U21091 (N_21091,N_16290,N_17824);
nand U21092 (N_21092,N_15718,N_15024);
or U21093 (N_21093,N_17559,N_18638);
nand U21094 (N_21094,N_16661,N_19524);
or U21095 (N_21095,N_17328,N_17795);
and U21096 (N_21096,N_19060,N_17598);
nand U21097 (N_21097,N_15692,N_16626);
nand U21098 (N_21098,N_18450,N_16183);
or U21099 (N_21099,N_15111,N_17678);
nand U21100 (N_21100,N_18769,N_16097);
xnor U21101 (N_21101,N_18798,N_19314);
nor U21102 (N_21102,N_17812,N_19313);
or U21103 (N_21103,N_15511,N_19294);
xor U21104 (N_21104,N_19944,N_18538);
or U21105 (N_21105,N_19814,N_15597);
or U21106 (N_21106,N_17487,N_19433);
xor U21107 (N_21107,N_18541,N_16737);
nor U21108 (N_21108,N_16844,N_15871);
xor U21109 (N_21109,N_16423,N_19942);
and U21110 (N_21110,N_15120,N_15753);
nand U21111 (N_21111,N_18204,N_16134);
xor U21112 (N_21112,N_15033,N_16308);
xnor U21113 (N_21113,N_19420,N_17460);
nand U21114 (N_21114,N_17921,N_15865);
nand U21115 (N_21115,N_15341,N_17780);
and U21116 (N_21116,N_19311,N_15141);
or U21117 (N_21117,N_15831,N_18502);
nand U21118 (N_21118,N_19361,N_17632);
xor U21119 (N_21119,N_19350,N_15505);
nor U21120 (N_21120,N_16395,N_16718);
nor U21121 (N_21121,N_19476,N_19620);
nor U21122 (N_21122,N_15624,N_15548);
nand U21123 (N_21123,N_17941,N_17318);
xnor U21124 (N_21124,N_16834,N_18179);
and U21125 (N_21125,N_15623,N_19993);
or U21126 (N_21126,N_17149,N_17140);
or U21127 (N_21127,N_18791,N_16255);
or U21128 (N_21128,N_19840,N_18285);
or U21129 (N_21129,N_18360,N_16705);
nand U21130 (N_21130,N_19708,N_16799);
and U21131 (N_21131,N_16277,N_18996);
or U21132 (N_21132,N_15780,N_17033);
or U21133 (N_21133,N_19335,N_15374);
nor U21134 (N_21134,N_16341,N_16202);
xor U21135 (N_21135,N_17566,N_19341);
nand U21136 (N_21136,N_16284,N_16704);
nor U21137 (N_21137,N_17420,N_15389);
xnor U21138 (N_21138,N_19588,N_19713);
and U21139 (N_21139,N_19182,N_19213);
nand U21140 (N_21140,N_15081,N_18497);
xor U21141 (N_21141,N_19260,N_18275);
and U21142 (N_21142,N_16717,N_18129);
nor U21143 (N_21143,N_17340,N_19847);
or U21144 (N_21144,N_16587,N_16732);
or U21145 (N_21145,N_18831,N_16120);
nor U21146 (N_21146,N_19858,N_17877);
or U21147 (N_21147,N_18170,N_19916);
and U21148 (N_21148,N_16854,N_15735);
or U21149 (N_21149,N_17164,N_15527);
nor U21150 (N_21150,N_19471,N_19551);
xnor U21151 (N_21151,N_15336,N_16141);
nand U21152 (N_21152,N_16206,N_16578);
or U21153 (N_21153,N_17403,N_16595);
nor U21154 (N_21154,N_16366,N_17584);
and U21155 (N_21155,N_17756,N_18817);
xor U21156 (N_21156,N_15881,N_15333);
or U21157 (N_21157,N_15773,N_15919);
xor U21158 (N_21158,N_16429,N_19921);
or U21159 (N_21159,N_15657,N_15312);
nor U21160 (N_21160,N_15558,N_19133);
and U21161 (N_21161,N_15386,N_18953);
xnor U21162 (N_21162,N_19273,N_17951);
nand U21163 (N_21163,N_16256,N_19940);
xnor U21164 (N_21164,N_19296,N_16647);
xor U21165 (N_21165,N_15741,N_19631);
xor U21166 (N_21166,N_15784,N_17526);
nand U21167 (N_21167,N_15003,N_15442);
xor U21168 (N_21168,N_18688,N_17625);
nand U21169 (N_21169,N_15447,N_18656);
xnor U21170 (N_21170,N_18366,N_19059);
nand U21171 (N_21171,N_15982,N_18031);
and U21172 (N_21172,N_17202,N_16422);
or U21173 (N_21173,N_16825,N_16823);
and U21174 (N_21174,N_15713,N_16536);
nor U21175 (N_21175,N_17103,N_17927);
or U21176 (N_21176,N_16133,N_19999);
or U21177 (N_21177,N_18590,N_17363);
xnor U21178 (N_21178,N_16696,N_19242);
nand U21179 (N_21179,N_15765,N_17194);
nor U21180 (N_21180,N_16589,N_19804);
and U21181 (N_21181,N_15195,N_19193);
xor U21182 (N_21182,N_18848,N_18060);
or U21183 (N_21183,N_17744,N_17860);
or U21184 (N_21184,N_19901,N_17112);
xor U21185 (N_21185,N_18551,N_16264);
xnor U21186 (N_21186,N_19149,N_16021);
nand U21187 (N_21187,N_18634,N_18941);
and U21188 (N_21188,N_18263,N_16325);
nand U21189 (N_21189,N_15104,N_16123);
nand U21190 (N_21190,N_19302,N_15772);
or U21191 (N_21191,N_18898,N_16378);
or U21192 (N_21192,N_17763,N_15150);
or U21193 (N_21193,N_19478,N_19578);
and U21194 (N_21194,N_18267,N_17739);
or U21195 (N_21195,N_18433,N_17669);
and U21196 (N_21196,N_16452,N_18163);
or U21197 (N_21197,N_19327,N_19033);
and U21198 (N_21198,N_16419,N_19486);
or U21199 (N_21199,N_19346,N_16475);
or U21200 (N_21200,N_19990,N_19951);
nand U21201 (N_21201,N_18610,N_15011);
nand U21202 (N_21202,N_15914,N_19627);
xor U21203 (N_21203,N_15984,N_15645);
and U21204 (N_21204,N_18474,N_15889);
nand U21205 (N_21205,N_16244,N_17094);
and U21206 (N_21206,N_16310,N_17483);
and U21207 (N_21207,N_19175,N_15340);
nand U21208 (N_21208,N_17896,N_18670);
or U21209 (N_21209,N_19709,N_17947);
xnor U21210 (N_21210,N_19557,N_16224);
nand U21211 (N_21211,N_18549,N_15560);
nor U21212 (N_21212,N_15416,N_19453);
or U21213 (N_21213,N_17326,N_16887);
xor U21214 (N_21214,N_19418,N_17106);
nor U21215 (N_21215,N_17376,N_16601);
or U21216 (N_21216,N_19177,N_18869);
or U21217 (N_21217,N_16677,N_15988);
or U21218 (N_21218,N_19379,N_17809);
or U21219 (N_21219,N_16944,N_18987);
nand U21220 (N_21220,N_15675,N_15032);
nor U21221 (N_21221,N_16044,N_19606);
nand U21222 (N_21222,N_19026,N_15604);
nor U21223 (N_21223,N_18335,N_18482);
or U21224 (N_21224,N_15895,N_18012);
nor U21225 (N_21225,N_16949,N_15291);
xor U21226 (N_21226,N_15144,N_17130);
nor U21227 (N_21227,N_16667,N_19694);
xor U21228 (N_21228,N_19815,N_16040);
and U21229 (N_21229,N_17165,N_18307);
xor U21230 (N_21230,N_19555,N_19326);
and U21231 (N_21231,N_17244,N_16390);
xnor U21232 (N_21232,N_18115,N_15993);
nor U21233 (N_21233,N_19256,N_18524);
nor U21234 (N_21234,N_18787,N_15690);
xor U21235 (N_21235,N_18128,N_16934);
or U21236 (N_21236,N_19455,N_17474);
xor U21237 (N_21237,N_19765,N_17123);
nor U21238 (N_21238,N_19859,N_15005);
nor U21239 (N_21239,N_17207,N_16176);
xnor U21240 (N_21240,N_17879,N_17772);
nand U21241 (N_21241,N_17043,N_18236);
nand U21242 (N_21242,N_19116,N_17974);
or U21243 (N_21243,N_16160,N_19429);
or U21244 (N_21244,N_17100,N_15896);
or U21245 (N_21245,N_18578,N_17431);
xor U21246 (N_21246,N_15905,N_18363);
nand U21247 (N_21247,N_16490,N_16898);
or U21248 (N_21248,N_16869,N_16102);
nor U21249 (N_21249,N_18540,N_18084);
nor U21250 (N_21250,N_17448,N_19322);
and U21251 (N_21251,N_17855,N_17013);
and U21252 (N_21252,N_16122,N_16115);
or U21253 (N_21253,N_17577,N_16579);
and U21254 (N_21254,N_18874,N_17496);
and U21255 (N_21255,N_16294,N_15779);
nand U21256 (N_21256,N_19523,N_17512);
nand U21257 (N_21257,N_15137,N_19580);
xor U21258 (N_21258,N_15134,N_17787);
or U21259 (N_21259,N_19613,N_15298);
or U21260 (N_21260,N_18418,N_15362);
or U21261 (N_21261,N_17685,N_19002);
or U21262 (N_21262,N_17522,N_18182);
or U21263 (N_21263,N_15064,N_17875);
nand U21264 (N_21264,N_16327,N_16850);
or U21265 (N_21265,N_19824,N_19740);
and U21266 (N_21266,N_19757,N_19618);
nand U21267 (N_21267,N_18254,N_19533);
xor U21268 (N_21268,N_19668,N_15279);
xor U21269 (N_21269,N_17742,N_17607);
nand U21270 (N_21270,N_15153,N_17159);
or U21271 (N_21271,N_16621,N_15959);
nand U21272 (N_21272,N_18728,N_18191);
or U21273 (N_21273,N_16914,N_15110);
nor U21274 (N_21274,N_19929,N_18293);
xor U21275 (N_21275,N_19949,N_17217);
or U21276 (N_21276,N_19646,N_16959);
or U21277 (N_21277,N_18039,N_16056);
nand U21278 (N_21278,N_16182,N_19601);
xnor U21279 (N_21279,N_17996,N_17942);
or U21280 (N_21280,N_18828,N_16711);
nor U21281 (N_21281,N_17800,N_19643);
or U21282 (N_21282,N_16992,N_15130);
and U21283 (N_21283,N_16243,N_18768);
nand U21284 (N_21284,N_15535,N_19775);
nand U21285 (N_21285,N_16502,N_19574);
nand U21286 (N_21286,N_19275,N_18047);
nand U21287 (N_21287,N_16001,N_18501);
or U21288 (N_21288,N_16522,N_17707);
nand U21289 (N_21289,N_17158,N_16379);
and U21290 (N_21290,N_15054,N_18385);
nor U21291 (N_21291,N_19563,N_17129);
nand U21292 (N_21292,N_19250,N_19372);
xnor U21293 (N_21293,N_17445,N_17829);
nand U21294 (N_21294,N_17206,N_15408);
and U21295 (N_21295,N_18858,N_16400);
and U21296 (N_21296,N_19241,N_17278);
nand U21297 (N_21297,N_17329,N_19873);
nand U21298 (N_21298,N_19291,N_18225);
nand U21299 (N_21299,N_16545,N_17032);
xnor U21300 (N_21300,N_18962,N_18936);
nor U21301 (N_21301,N_15281,N_18384);
nor U21302 (N_21302,N_15547,N_15278);
nand U21303 (N_21303,N_16465,N_18725);
or U21304 (N_21304,N_17330,N_16598);
xor U21305 (N_21305,N_16521,N_19202);
and U21306 (N_21306,N_17253,N_18851);
nor U21307 (N_21307,N_16111,N_17293);
nand U21308 (N_21308,N_15313,N_18846);
nor U21309 (N_21309,N_17706,N_16459);
nor U21310 (N_21310,N_19727,N_18758);
xor U21311 (N_21311,N_18640,N_18378);
nand U21312 (N_21312,N_19519,N_19784);
or U21313 (N_21313,N_19738,N_17042);
nor U21314 (N_21314,N_19753,N_19472);
nand U21315 (N_21315,N_15646,N_19776);
nand U21316 (N_21316,N_15839,N_16608);
nor U21317 (N_21317,N_16406,N_17981);
or U21318 (N_21318,N_17014,N_18500);
xor U21319 (N_21319,N_18658,N_19239);
nand U21320 (N_21320,N_15016,N_17767);
and U21321 (N_21321,N_18175,N_19891);
nor U21322 (N_21322,N_15807,N_17982);
xor U21323 (N_21323,N_19333,N_19648);
nand U21324 (N_21324,N_15933,N_19672);
nand U21325 (N_21325,N_19497,N_17799);
nand U21326 (N_21326,N_19889,N_19003);
xor U21327 (N_21327,N_18398,N_19075);
xnor U21328 (N_21328,N_17843,N_18185);
xor U21329 (N_21329,N_18208,N_17730);
nand U21330 (N_21330,N_17959,N_16906);
nor U21331 (N_21331,N_15873,N_15397);
nor U21332 (N_21332,N_18963,N_18529);
nor U21333 (N_21333,N_19457,N_19829);
nand U21334 (N_21334,N_17846,N_19163);
and U21335 (N_21335,N_19818,N_16085);
or U21336 (N_21336,N_19903,N_16471);
xnor U21337 (N_21337,N_15586,N_17736);
or U21338 (N_21338,N_19362,N_18910);
xnor U21339 (N_21339,N_18215,N_16331);
or U21340 (N_21340,N_17075,N_16979);
nand U21341 (N_21341,N_16549,N_18862);
xor U21342 (N_21342,N_16412,N_16683);
nand U21343 (N_21343,N_16638,N_18559);
or U21344 (N_21344,N_19338,N_16770);
xnor U21345 (N_21345,N_16875,N_16826);
nor U21346 (N_21346,N_18849,N_18078);
xor U21347 (N_21347,N_17248,N_17342);
and U21348 (N_21348,N_19791,N_17212);
and U21349 (N_21349,N_17439,N_16216);
and U21350 (N_21350,N_18894,N_15487);
nand U21351 (N_21351,N_18518,N_19447);
xor U21352 (N_21352,N_16159,N_17975);
xor U21353 (N_21353,N_19652,N_18150);
and U21354 (N_21354,N_17099,N_15034);
and U21355 (N_21355,N_18325,N_18284);
xor U21356 (N_21356,N_16730,N_19637);
nor U21357 (N_21357,N_19160,N_17604);
xor U21358 (N_21358,N_16329,N_17818);
or U21359 (N_21359,N_19058,N_16994);
or U21360 (N_21360,N_15154,N_16975);
xor U21361 (N_21361,N_17731,N_17498);
and U21362 (N_21362,N_15357,N_17762);
and U21363 (N_21363,N_17359,N_19507);
nand U21364 (N_21364,N_15797,N_19780);
and U21365 (N_21365,N_18912,N_16609);
xor U21366 (N_21366,N_17601,N_16819);
and U21367 (N_21367,N_17953,N_15569);
or U21368 (N_21368,N_15157,N_18821);
xnor U21369 (N_21369,N_15802,N_19629);
and U21370 (N_21370,N_19587,N_15770);
xnor U21371 (N_21371,N_18833,N_17150);
and U21372 (N_21372,N_17998,N_19208);
and U21373 (N_21373,N_17222,N_16531);
and U21374 (N_21374,N_19112,N_15835);
nand U21375 (N_21375,N_19148,N_18473);
nor U21376 (N_21376,N_19123,N_18494);
or U21377 (N_21377,N_16037,N_16851);
xor U21378 (N_21378,N_19380,N_18124);
nand U21379 (N_21379,N_19319,N_16289);
or U21380 (N_21380,N_19924,N_19073);
and U21381 (N_21381,N_16874,N_18329);
and U21382 (N_21382,N_16285,N_16891);
or U21383 (N_21383,N_18539,N_16024);
nor U21384 (N_21384,N_19071,N_19809);
xor U21385 (N_21385,N_15240,N_19393);
xnor U21386 (N_21386,N_15674,N_18949);
nor U21387 (N_21387,N_16262,N_18562);
or U21388 (N_21388,N_18789,N_19670);
and U21389 (N_21389,N_17848,N_15479);
xor U21390 (N_21390,N_18451,N_18973);
nand U21391 (N_21391,N_17680,N_16796);
nand U21392 (N_21392,N_19255,N_15265);
nor U21393 (N_21393,N_17968,N_18476);
or U21394 (N_21394,N_19673,N_19739);
and U21395 (N_21395,N_16716,N_18903);
or U21396 (N_21396,N_19331,N_19205);
nand U21397 (N_21397,N_16935,N_17281);
or U21398 (N_21398,N_15378,N_18241);
nor U21399 (N_21399,N_15346,N_17366);
xor U21400 (N_21400,N_16983,N_19378);
nor U21401 (N_21401,N_18799,N_19421);
nor U21402 (N_21402,N_19654,N_18160);
nand U21403 (N_21403,N_18272,N_15688);
nor U21404 (N_21404,N_16774,N_19704);
nor U21405 (N_21405,N_15221,N_19254);
and U21406 (N_21406,N_18238,N_18157);
xor U21407 (N_21407,N_16346,N_16830);
nor U21408 (N_21408,N_15306,N_16067);
xnor U21409 (N_21409,N_18950,N_18667);
nand U21410 (N_21410,N_15972,N_15296);
or U21411 (N_21411,N_17442,N_15105);
or U21412 (N_21412,N_18291,N_17883);
or U21413 (N_21413,N_18338,N_15670);
nand U21414 (N_21414,N_15253,N_18689);
or U21415 (N_21415,N_19221,N_18146);
and U21416 (N_21416,N_15371,N_16209);
nor U21417 (N_21417,N_17429,N_18417);
nand U21418 (N_21418,N_19107,N_18032);
xnor U21419 (N_21419,N_16145,N_18005);
nand U21420 (N_21420,N_17653,N_19801);
xor U21421 (N_21421,N_17634,N_17682);
nand U21422 (N_21422,N_17186,N_16177);
and U21423 (N_21423,N_17157,N_17418);
and U21424 (N_21424,N_17719,N_15669);
nand U21425 (N_21425,N_19608,N_17728);
nor U21426 (N_21426,N_16396,N_16483);
xnor U21427 (N_21427,N_15563,N_16242);
nand U21428 (N_21428,N_19710,N_19233);
xnor U21429 (N_21429,N_16065,N_15523);
xor U21430 (N_21430,N_15256,N_15813);
nor U21431 (N_21431,N_16298,N_15305);
xnor U21432 (N_21432,N_19134,N_19137);
and U21433 (N_21433,N_17540,N_18220);
or U21434 (N_21434,N_19192,N_15997);
xnor U21435 (N_21435,N_18332,N_19168);
nor U21436 (N_21436,N_17383,N_19120);
xor U21437 (N_21437,N_17660,N_15788);
nand U21438 (N_21438,N_17510,N_17305);
and U21439 (N_21439,N_17623,N_18209);
and U21440 (N_21440,N_19834,N_17989);
nand U21441 (N_21441,N_18601,N_19386);
nor U21442 (N_21442,N_18615,N_17663);
or U21443 (N_21443,N_15262,N_18631);
nor U21444 (N_21444,N_18591,N_16050);
nor U21445 (N_21445,N_17470,N_17287);
and U21446 (N_21446,N_16349,N_18002);
nor U21447 (N_21447,N_17135,N_16650);
xor U21448 (N_21448,N_17615,N_19475);
nand U21449 (N_21449,N_15210,N_15352);
nand U21450 (N_21450,N_19910,N_18820);
nor U21451 (N_21451,N_18134,N_19308);
xor U21452 (N_21452,N_17916,N_16496);
or U21453 (N_21453,N_16808,N_19947);
nand U21454 (N_21454,N_18704,N_17865);
nand U21455 (N_21455,N_15599,N_16862);
xnor U21456 (N_21456,N_15076,N_17958);
nor U21457 (N_21457,N_16859,N_16886);
nand U21458 (N_21458,N_17972,N_16098);
nor U21459 (N_21459,N_19830,N_19488);
nor U21460 (N_21460,N_17173,N_19028);
and U21461 (N_21461,N_16922,N_19931);
xnor U21462 (N_21462,N_16051,N_19667);
and U21463 (N_21463,N_15519,N_17580);
nor U21464 (N_21464,N_18169,N_19736);
nand U21465 (N_21465,N_18994,N_19530);
or U21466 (N_21466,N_17267,N_17250);
nor U21467 (N_21467,N_19009,N_17882);
nor U21468 (N_21468,N_17069,N_16058);
nor U21469 (N_21469,N_19640,N_18101);
nor U21470 (N_21470,N_16438,N_15348);
nand U21471 (N_21471,N_18574,N_16273);
nor U21472 (N_21472,N_17310,N_19750);
or U21473 (N_21473,N_18641,N_18297);
or U21474 (N_21474,N_17336,N_18911);
and U21475 (N_21475,N_19494,N_19489);
and U21476 (N_21476,N_19937,N_18049);
nand U21477 (N_21477,N_18617,N_17204);
xnor U21478 (N_21478,N_18119,N_16199);
nand U21479 (N_21479,N_18252,N_18586);
xnor U21480 (N_21480,N_15910,N_16146);
and U21481 (N_21481,N_17052,N_16498);
and U21482 (N_21482,N_16676,N_19336);
nand U21483 (N_21483,N_16813,N_17029);
nand U21484 (N_21484,N_15502,N_15079);
nand U21485 (N_21485,N_16283,N_15425);
xor U21486 (N_21486,N_19890,N_15146);
xnor U21487 (N_21487,N_17726,N_16731);
and U21488 (N_21488,N_18925,N_15364);
or U21489 (N_21489,N_17993,N_16451);
xor U21490 (N_21490,N_18126,N_16272);
and U21491 (N_21491,N_15983,N_18878);
nor U21492 (N_21492,N_16074,N_17299);
nand U21493 (N_21493,N_15903,N_18909);
nand U21494 (N_21494,N_16398,N_19076);
nor U21495 (N_21495,N_15714,N_19405);
nor U21496 (N_21496,N_15924,N_16797);
nand U21497 (N_21497,N_15676,N_19278);
nand U21498 (N_21498,N_15411,N_16288);
nand U21499 (N_21499,N_15515,N_19354);
or U21500 (N_21500,N_16251,N_19235);
and U21501 (N_21501,N_16712,N_15434);
nand U21502 (N_21502,N_15143,N_19014);
or U21503 (N_21503,N_15324,N_16011);
nor U21504 (N_21504,N_16237,N_15728);
xor U21505 (N_21505,N_17523,N_18331);
xor U21506 (N_21506,N_16861,N_19339);
xnor U21507 (N_21507,N_17781,N_18719);
nand U21508 (N_21508,N_18714,N_18637);
and U21509 (N_21509,N_16357,N_18009);
nor U21510 (N_21510,N_16678,N_18767);
and U21511 (N_21511,N_16300,N_16275);
xor U21512 (N_21512,N_18935,N_17252);
nand U21513 (N_21513,N_17899,N_15369);
nor U21514 (N_21514,N_15509,N_15211);
xnor U21515 (N_21515,N_18605,N_16253);
xnor U21516 (N_21516,N_16113,N_18334);
xnor U21517 (N_21517,N_18702,N_18928);
nor U21518 (N_21518,N_18340,N_15404);
nand U21519 (N_21519,N_19303,N_16286);
nand U21520 (N_21520,N_16154,N_16865);
or U21521 (N_21521,N_15803,N_16472);
nor U21522 (N_21522,N_19181,N_18477);
and U21523 (N_21523,N_18458,N_17961);
nand U21524 (N_21524,N_16031,N_18881);
nor U21525 (N_21525,N_16866,N_18362);
and U21526 (N_21526,N_16364,N_18845);
xnor U21527 (N_21527,N_17243,N_18660);
or U21528 (N_21528,N_15161,N_15659);
xor U21529 (N_21529,N_18480,N_17337);
and U21530 (N_21530,N_17218,N_15853);
nor U21531 (N_21531,N_18522,N_19684);
and U21532 (N_21532,N_16055,N_18264);
nand U21533 (N_21533,N_15666,N_16744);
nand U21534 (N_21534,N_16508,N_18782);
and U21535 (N_21535,N_19367,N_18309);
xnor U21536 (N_21536,N_16342,N_16548);
and U21537 (N_21537,N_17794,N_16929);
or U21538 (N_21538,N_16470,N_19051);
and U21539 (N_21539,N_16108,N_17712);
nor U21540 (N_21540,N_15531,N_15314);
nand U21541 (N_21541,N_19806,N_17593);
and U21542 (N_21542,N_17497,N_18572);
nand U21543 (N_21543,N_17574,N_17907);
nand U21544 (N_21544,N_15206,N_15155);
or U21545 (N_21545,N_15254,N_19883);
or U21546 (N_21546,N_16336,N_17911);
nand U21547 (N_21547,N_15501,N_15451);
xnor U21548 (N_21548,N_16409,N_17553);
nor U21549 (N_21549,N_16132,N_17618);
nand U21550 (N_21550,N_15756,N_16118);
and U21551 (N_21551,N_16468,N_16909);
or U21552 (N_21552,N_15962,N_16636);
xor U21553 (N_21553,N_16915,N_18327);
nand U21554 (N_21554,N_18866,N_18452);
or U21555 (N_21555,N_17793,N_15299);
nand U21556 (N_21556,N_19918,N_19490);
xnor U21557 (N_21557,N_18229,N_15332);
nor U21558 (N_21558,N_18864,N_17531);
and U21559 (N_21559,N_17060,N_19584);
and U21560 (N_21560,N_18918,N_16292);
or U21561 (N_21561,N_19343,N_17715);
and U21562 (N_21562,N_16908,N_16889);
nor U21563 (N_21563,N_18316,N_19087);
xnor U21564 (N_21564,N_18712,N_16072);
nand U21565 (N_21565,N_18604,N_19553);
nor U21566 (N_21566,N_17122,N_18984);
nand U21567 (N_21567,N_18290,N_17847);
xnor U21568 (N_21568,N_18600,N_19090);
and U21569 (N_21569,N_19165,N_17885);
nand U21570 (N_21570,N_18691,N_18028);
and U21571 (N_21571,N_17397,N_18235);
and U21572 (N_21572,N_16164,N_17247);
nor U21573 (N_21573,N_15726,N_19184);
nor U21574 (N_21574,N_16721,N_17543);
or U21575 (N_21575,N_18467,N_18736);
xor U21576 (N_21576,N_18517,N_19565);
nand U21577 (N_21577,N_17215,N_19793);
or U21578 (N_21578,N_18761,N_16112);
nor U21579 (N_21579,N_17997,N_16895);
nand U21580 (N_21580,N_15468,N_16769);
nor U21581 (N_21581,N_19505,N_17525);
nand U21582 (N_21582,N_18979,N_15290);
nand U21583 (N_21583,N_16114,N_16682);
xnor U21584 (N_21584,N_19008,N_18956);
xor U21585 (N_21585,N_19969,N_15323);
xor U21586 (N_21586,N_18643,N_19054);
nand U21587 (N_21587,N_17909,N_15045);
nor U21588 (N_21588,N_15609,N_18246);
or U21589 (N_21589,N_19591,N_19344);
nand U21590 (N_21590,N_16071,N_17334);
nand U21591 (N_21591,N_17630,N_17755);
and U21592 (N_21592,N_15854,N_16633);
nor U21593 (N_21593,N_15589,N_19771);
or U21594 (N_21594,N_17440,N_18896);
and U21595 (N_21595,N_19370,N_19948);
and U21596 (N_21596,N_18662,N_16332);
xnor U21597 (N_21597,N_18105,N_18226);
and U21598 (N_21598,N_16568,N_17018);
nor U21599 (N_21599,N_16220,N_19253);
and U21600 (N_21600,N_17229,N_17457);
nor U21601 (N_21601,N_15027,N_18400);
nand U21602 (N_21602,N_17757,N_16755);
and U21603 (N_21603,N_17976,N_16453);
or U21604 (N_21604,N_15652,N_17913);
or U21605 (N_21605,N_19118,N_18436);
or U21606 (N_21606,N_18865,N_16425);
and U21607 (N_21607,N_15013,N_17280);
nand U21608 (N_21608,N_16025,N_19526);
and U21609 (N_21609,N_16800,N_16822);
or U21610 (N_21610,N_15693,N_19609);
nand U21611 (N_21611,N_18221,N_16838);
nand U21612 (N_21612,N_16597,N_18139);
xnor U21613 (N_21613,N_19970,N_16420);
or U21614 (N_21614,N_15438,N_15331);
nor U21615 (N_21615,N_19262,N_16265);
xor U21616 (N_21616,N_16843,N_16131);
and U21617 (N_21617,N_16848,N_19712);
nand U21618 (N_21618,N_18566,N_15356);
xnor U21619 (N_21619,N_15577,N_17447);
and U21620 (N_21620,N_19145,N_19038);
nand U21621 (N_21621,N_18058,N_19603);
and U21622 (N_21622,N_19417,N_18024);
nor U21623 (N_21623,N_17109,N_18116);
or U21624 (N_21624,N_17782,N_18888);
nor U21625 (N_21625,N_16871,N_19402);
and U21626 (N_21626,N_15304,N_16228);
and U21627 (N_21627,N_16528,N_19756);
or U21628 (N_21628,N_16686,N_19057);
and U21629 (N_21629,N_17221,N_17863);
nor U21630 (N_21630,N_19959,N_19846);
and U21631 (N_21631,N_18243,N_19909);
nor U21632 (N_21632,N_16556,N_18971);
nor U21633 (N_21633,N_15276,N_16781);
or U21634 (N_21634,N_17708,N_15746);
and U21635 (N_21635,N_17227,N_19093);
xnor U21636 (N_21636,N_16688,N_15360);
xor U21637 (N_21637,N_16473,N_15761);
nand U21638 (N_21638,N_18401,N_17025);
nor U21639 (N_21639,N_17667,N_18130);
nand U21640 (N_21640,N_16779,N_18253);
and U21641 (N_21641,N_15909,N_18472);
nor U21642 (N_21642,N_19363,N_16918);
nand U21643 (N_21643,N_18168,N_18158);
nand U21644 (N_21644,N_18445,N_15827);
nand U21645 (N_21645,N_17456,N_19401);
nor U21646 (N_21646,N_17987,N_15731);
nand U21647 (N_21647,N_15267,N_19676);
and U21648 (N_21648,N_15190,N_19047);
nand U21649 (N_21649,N_15242,N_18018);
xnor U21650 (N_21650,N_16437,N_18199);
nand U21651 (N_21651,N_16053,N_16651);
and U21652 (N_21652,N_19875,N_16376);
and U21653 (N_21653,N_18510,N_16820);
xor U21654 (N_21654,N_18665,N_19377);
or U21655 (N_21655,N_15463,N_19592);
and U21656 (N_21656,N_17003,N_17771);
and U21657 (N_21657,N_15760,N_19230);
or U21658 (N_21658,N_17915,N_17443);
and U21659 (N_21659,N_19258,N_17925);
and U21660 (N_21660,N_18063,N_15791);
or U21661 (N_21661,N_17317,N_16299);
xor U21662 (N_21662,N_18256,N_16933);
nand U21663 (N_21663,N_15503,N_17066);
nand U21664 (N_21664,N_19546,N_18310);
and U21665 (N_21665,N_16119,N_19657);
and U21666 (N_21666,N_18145,N_18991);
and U21667 (N_21667,N_15149,N_15945);
or U21668 (N_21668,N_19701,N_18164);
nand U21669 (N_21669,N_15295,N_16484);
nor U21670 (N_21670,N_17282,N_17108);
xnor U21671 (N_21671,N_19365,N_19799);
and U21672 (N_21672,N_15272,N_18245);
and U21673 (N_21673,N_19642,N_17346);
xnor U21674 (N_21674,N_17034,N_16381);
nand U21675 (N_21675,N_19680,N_17082);
nor U21676 (N_21676,N_17364,N_19726);
nand U21677 (N_21677,N_16351,N_17664);
and U21678 (N_21678,N_17187,N_16960);
nand U21679 (N_21679,N_19669,N_15937);
nor U21680 (N_21680,N_17872,N_19454);
nor U21681 (N_21681,N_15215,N_16707);
or U21682 (N_21682,N_18793,N_18465);
and U21683 (N_21683,N_16768,N_16238);
or U21684 (N_21684,N_18785,N_17232);
or U21685 (N_21685,N_15719,N_15355);
or U21686 (N_21686,N_18437,N_17792);
or U21687 (N_21687,N_15617,N_19069);
or U21688 (N_21688,N_19366,N_15781);
xnor U21689 (N_21689,N_16687,N_15928);
nor U21690 (N_21690,N_15898,N_16030);
or U21691 (N_21691,N_19034,N_18065);
xnor U21692 (N_21692,N_17044,N_15351);
nand U21693 (N_21693,N_15960,N_19364);
or U21694 (N_21694,N_17748,N_17061);
nor U21695 (N_21695,N_17501,N_18550);
or U21696 (N_21696,N_16503,N_17098);
or U21697 (N_21697,N_16928,N_16248);
nor U21698 (N_21698,N_17670,N_18015);
nor U21699 (N_21699,N_19355,N_15219);
nand U21700 (N_21700,N_17063,N_19067);
or U21701 (N_21701,N_18042,N_15194);
and U21702 (N_21702,N_15455,N_18081);
xnor U21703 (N_21703,N_15611,N_16084);
xor U21704 (N_21704,N_19017,N_19862);
nand U21705 (N_21705,N_16618,N_18784);
nor U21706 (N_21706,N_18934,N_15222);
or U21707 (N_21707,N_18094,N_16635);
nand U21708 (N_21708,N_18016,N_18294);
and U21709 (N_21709,N_17400,N_19122);
nand U21710 (N_21710,N_16469,N_19953);
xnor U21711 (N_21711,N_16384,N_19610);
xnor U21712 (N_21712,N_16892,N_18227);
nand U21713 (N_21713,N_16585,N_17850);
nor U21714 (N_21714,N_15689,N_15297);
and U21715 (N_21715,N_15540,N_17143);
or U21716 (N_21716,N_16599,N_17425);
or U21717 (N_21717,N_15556,N_16109);
nand U21718 (N_21718,N_15285,N_19625);
or U21719 (N_21719,N_19687,N_19512);
or U21720 (N_21720,N_17312,N_16976);
xnor U21721 (N_21721,N_19301,N_19272);
and U21722 (N_21722,N_15388,N_15575);
or U21723 (N_21723,N_15514,N_15856);
xor U21724 (N_21724,N_15704,N_19240);
nor U21725 (N_21725,N_17226,N_17562);
xnor U21726 (N_21726,N_15874,N_18021);
and U21727 (N_21727,N_18885,N_18321);
xnor U21728 (N_21728,N_17257,N_19906);
xor U21729 (N_21729,N_15762,N_15292);
nor U21730 (N_21730,N_15837,N_16239);
nor U21731 (N_21731,N_17716,N_16279);
and U21732 (N_21732,N_15334,N_17071);
xnor U21733 (N_21733,N_15258,N_17246);
or U21734 (N_21734,N_17609,N_19675);
nand U21735 (N_21735,N_15366,N_16581);
xor U21736 (N_21736,N_16572,N_16564);
nor U21737 (N_21737,N_17788,N_18504);
nand U21738 (N_21738,N_19400,N_18460);
nor U21739 (N_21739,N_15636,N_16968);
or U21740 (N_21740,N_19976,N_18222);
or U21741 (N_21741,N_16963,N_17661);
xnor U21742 (N_21742,N_18519,N_15224);
or U21743 (N_21743,N_17277,N_19029);
nand U21744 (N_21744,N_15405,N_16456);
nand U21745 (N_21745,N_15976,N_17827);
xnor U21746 (N_21746,N_16321,N_16610);
xor U21747 (N_21747,N_18707,N_15822);
xor U21748 (N_21748,N_19194,N_19248);
and U21749 (N_21749,N_18542,N_19774);
nor U21750 (N_21750,N_18357,N_19707);
xnor U21751 (N_21751,N_17826,N_18286);
or U21752 (N_21752,N_17672,N_18978);
or U21753 (N_21753,N_18295,N_15662);
and U21754 (N_21754,N_16362,N_18389);
xnor U21755 (N_21755,N_19690,N_17367);
xor U21756 (N_21756,N_18681,N_18838);
or U21757 (N_21757,N_16307,N_19879);
xor U21758 (N_21758,N_15922,N_17704);
nor U21759 (N_21759,N_19568,N_16104);
nor U21760 (N_21760,N_16478,N_15872);
or U21761 (N_21761,N_19068,N_16955);
or U21762 (N_21762,N_19495,N_18266);
nor U21763 (N_21763,N_17662,N_15385);
xor U21764 (N_21764,N_15573,N_15080);
xor U21765 (N_21765,N_17170,N_18214);
or U21766 (N_21766,N_15069,N_15329);
or U21767 (N_21767,N_16455,N_19570);
nand U21768 (N_21768,N_15537,N_19092);
nand U21769 (N_21769,N_17895,N_16554);
nor U21770 (N_21770,N_17409,N_15878);
or U21771 (N_21771,N_18990,N_15490);
nor U21772 (N_21772,N_17733,N_16987);
nor U21773 (N_21773,N_16537,N_18379);
nand U21774 (N_21774,N_17722,N_18154);
nand U21775 (N_21775,N_16247,N_15732);
nand U21776 (N_21776,N_16991,N_18304);
and U21777 (N_21777,N_17657,N_17764);
and U21778 (N_21778,N_17485,N_16415);
and U21779 (N_21779,N_17983,N_16315);
nand U21780 (N_21780,N_19994,N_17415);
or U21781 (N_21781,N_18230,N_18354);
xnor U21782 (N_21782,N_15241,N_18019);
nand U21783 (N_21783,N_18859,N_16821);
nor U21784 (N_21784,N_16229,N_18355);
nor U21785 (N_21785,N_18913,N_19955);
nor U21786 (N_21786,N_18947,N_16575);
xnor U21787 (N_21787,N_17765,N_16735);
and U21788 (N_21788,N_15469,N_18587);
xnor U21789 (N_21789,N_18342,N_18118);
nand U21790 (N_21790,N_15108,N_19348);
or U21791 (N_21791,N_15968,N_19664);
xnor U21792 (N_21792,N_17024,N_17300);
nor U21793 (N_21793,N_16702,N_19679);
nand U21794 (N_21794,N_18902,N_19538);
or U21795 (N_21795,N_15475,N_17546);
nand U21796 (N_21796,N_17535,N_16632);
and U21797 (N_21797,N_17031,N_18813);
nor U21798 (N_21798,N_16927,N_17045);
nand U21799 (N_21799,N_18496,N_16297);
or U21800 (N_21800,N_18583,N_15994);
and U21801 (N_21801,N_15140,N_17389);
or U21802 (N_21802,N_17920,N_16726);
nand U21803 (N_21803,N_19325,N_16810);
nor U21804 (N_21804,N_15745,N_19483);
or U21805 (N_21805,N_18231,N_19231);
or U21806 (N_21806,N_17449,N_16956);
or U21807 (N_21807,N_19186,N_19872);
xnor U21808 (N_21808,N_15309,N_18571);
or U21809 (N_21809,N_16354,N_17948);
or U21810 (N_21810,N_16439,N_16998);
nand U21811 (N_21811,N_15124,N_16162);
nor U21812 (N_21812,N_16526,N_16807);
nand U21813 (N_21813,N_19136,N_15319);
and U21814 (N_21814,N_19607,N_15917);
or U21815 (N_21815,N_17219,N_15413);
or U21816 (N_21816,N_15070,N_15383);
xor U21817 (N_21817,N_16814,N_16700);
xor U21818 (N_21818,N_18589,N_17720);
and U21819 (N_21819,N_19217,N_18186);
and U21820 (N_21820,N_19696,N_19404);
nor U21821 (N_21821,N_17116,N_19245);
nor U21822 (N_21822,N_17626,N_18181);
and U21823 (N_21823,N_17469,N_19692);
nand U21824 (N_21824,N_17026,N_16917);
nand U21825 (N_21825,N_18569,N_17466);
xor U21826 (N_21826,N_15673,N_17727);
or U21827 (N_21827,N_15119,N_17038);
nor U21828 (N_21828,N_16013,N_19651);
or U21829 (N_21829,N_19790,N_16559);
and U21830 (N_21830,N_17484,N_19376);
xnor U21831 (N_21831,N_18239,N_16622);
and U21832 (N_21832,N_16417,N_17390);
xor U21833 (N_21833,N_16809,N_17088);
nand U21834 (N_21834,N_16615,N_15060);
nor U21835 (N_21835,N_16660,N_19541);
xor U21836 (N_21836,N_18832,N_19894);
or U21837 (N_21837,N_15088,N_19191);
or U21838 (N_21838,N_18364,N_17545);
or U21839 (N_21839,N_19424,N_19785);
nor U21840 (N_21840,N_15484,N_19952);
xor U21841 (N_21841,N_17833,N_18805);
nor U21842 (N_21842,N_19443,N_17931);
xnor U21843 (N_21843,N_17779,N_17789);
xnor U21844 (N_21844,N_15750,N_16937);
nor U21845 (N_21845,N_17986,N_15603);
nor U21846 (N_21846,N_16584,N_16551);
nand U21847 (N_21847,N_19719,N_15402);
and U21848 (N_21848,N_16092,N_17814);
or U21849 (N_21849,N_16128,N_16281);
nand U21850 (N_21850,N_18988,N_19838);
nor U21851 (N_21851,N_15863,N_17859);
nor U21852 (N_21852,N_19759,N_16749);
xnor U21853 (N_21853,N_15017,N_15220);
and U21854 (N_21854,N_18074,N_19282);
nor U21855 (N_21855,N_17132,N_19977);
xnor U21856 (N_21856,N_16946,N_16135);
and U21857 (N_21857,N_19529,N_17433);
and U21858 (N_21858,N_16951,N_15677);
nor U21859 (N_21859,N_16152,N_16910);
or U21860 (N_21860,N_16685,N_16517);
and U21861 (N_21861,N_15115,N_19914);
or U21862 (N_21862,N_18983,N_19172);
or U21863 (N_21863,N_15829,N_18764);
and U21864 (N_21864,N_19266,N_17831);
and U21865 (N_21865,N_15182,N_17723);
nor U21866 (N_21866,N_16489,N_17276);
nor U21867 (N_21867,N_15178,N_17560);
xnor U21868 (N_21868,N_18056,N_18632);
nor U21869 (N_21869,N_16035,N_16474);
xor U21870 (N_21870,N_15387,N_16258);
xor U21871 (N_21871,N_15967,N_16370);
and U21872 (N_21872,N_15695,N_16506);
nand U21873 (N_21873,N_17679,N_16668);
nand U21874 (N_21874,N_15185,N_17900);
or U21875 (N_21875,N_19410,N_15950);
or U21876 (N_21876,N_19817,N_19371);
xnor U21877 (N_21877,N_16252,N_19535);
nand U21878 (N_21878,N_16148,N_15138);
nor U21879 (N_21879,N_19197,N_16923);
nand U21880 (N_21880,N_17341,N_15099);
nor U21881 (N_21881,N_15665,N_19857);
nor U21882 (N_21882,N_17537,N_18952);
and U21883 (N_21883,N_18694,N_18194);
nor U21884 (N_21884,N_17392,N_18668);
nor U21885 (N_21885,N_18746,N_19915);
and U21886 (N_21886,N_16629,N_15496);
nor U21887 (N_21887,N_19783,N_17450);
nand U21888 (N_21888,N_17912,N_18218);
or U21889 (N_21889,N_16467,N_15462);
and U21890 (N_21890,N_17513,N_16586);
xor U21891 (N_21891,N_15758,N_15188);
xor U21892 (N_21892,N_18972,N_15524);
and U21893 (N_21893,N_17195,N_15186);
xnor U21894 (N_21894,N_17966,N_15774);
nand U21895 (N_21895,N_17815,N_18276);
nor U21896 (N_21896,N_16018,N_19733);
and U21897 (N_21897,N_17090,N_19721);
and U21898 (N_21898,N_18369,N_16532);
nor U21899 (N_21899,N_15248,N_18664);
xor U21900 (N_21900,N_16245,N_15096);
and U21901 (N_21901,N_19446,N_15825);
or U21902 (N_21902,N_18071,N_15381);
nor U21903 (N_21903,N_16888,N_17935);
and U21904 (N_21904,N_17051,N_17639);
or U21905 (N_21905,N_16431,N_15516);
nand U21906 (N_21906,N_18299,N_17030);
and U21907 (N_21907,N_17515,N_17588);
and U21908 (N_21908,N_16977,N_15072);
xor U21909 (N_21909,N_19470,N_16339);
xnor U21910 (N_21910,N_18645,N_17928);
and U21911 (N_21911,N_18695,N_15957);
nor U21912 (N_21912,N_19099,N_18070);
nand U21913 (N_21913,N_18526,N_15980);
nand U21914 (N_21914,N_16645,N_19509);
nor U21915 (N_21915,N_19061,N_16828);
nand U21916 (N_21916,N_18217,N_16259);
or U21917 (N_21917,N_19480,N_17021);
nand U21918 (N_21918,N_17479,N_15810);
nand U21919 (N_21919,N_18581,N_16641);
nor U21920 (N_21920,N_18717,N_19236);
xor U21921 (N_21921,N_18257,N_19232);
xor U21922 (N_21922,N_16833,N_19536);
and U21923 (N_21923,N_15477,N_19911);
xor U21924 (N_21924,N_17671,N_18711);
nor U21925 (N_21925,N_18183,N_16314);
xor U21926 (N_21926,N_15929,N_19216);
nor U21927 (N_21927,N_18425,N_18630);
xor U21928 (N_21928,N_19665,N_17285);
or U21929 (N_21929,N_19661,N_15179);
xor U21930 (N_21930,N_16143,N_19644);
xnor U21931 (N_21931,N_15053,N_15283);
or U21932 (N_21932,N_15251,N_18766);
nor U21933 (N_21933,N_17579,N_19717);
nand U21934 (N_21934,N_18131,N_17918);
nand U21935 (N_21935,N_19238,N_15694);
and U21936 (N_21936,N_17703,N_18649);
or U21937 (N_21937,N_15619,N_18149);
nand U21938 (N_21938,N_18123,N_17355);
or U21939 (N_21939,N_18958,N_15751);
xor U21940 (N_21940,N_17395,N_16343);
nor U21941 (N_21941,N_18967,N_15618);
xor U21942 (N_21942,N_17926,N_17813);
and U21943 (N_21943,N_16207,N_15320);
xor U21944 (N_21944,N_18596,N_15934);
and U21945 (N_21945,N_16004,N_18259);
nor U21946 (N_21946,N_18806,N_15823);
nand U21947 (N_21947,N_17500,N_17437);
xor U21948 (N_21948,N_17929,N_16969);
xor U21949 (N_21949,N_17791,N_17977);
nand U21950 (N_21950,N_16060,N_15809);
xnor U21951 (N_21951,N_18424,N_15696);
and U21952 (N_21952,N_17973,N_19324);
or U21953 (N_21953,N_15533,N_16763);
nor U21954 (N_21954,N_16218,N_15532);
and U21955 (N_21955,N_18095,N_18907);
nor U21956 (N_21956,N_17091,N_16643);
nor U21957 (N_21957,N_17919,N_17988);
or U21958 (N_21958,N_18189,N_16214);
nor U21959 (N_21959,N_15518,N_16416);
xor U21960 (N_21960,N_18863,N_18122);
nand U21961 (N_21961,N_19855,N_16241);
or U21962 (N_21962,N_18876,N_15133);
nor U21963 (N_21963,N_16350,N_18430);
xnor U21964 (N_21964,N_17084,N_19451);
xnor U21965 (N_21965,N_17438,N_15512);
nand U21966 (N_21966,N_18584,N_17234);
xor U21967 (N_21967,N_16059,N_18410);
and U21968 (N_21968,N_19985,N_19773);
nor U21969 (N_21969,N_19593,N_15702);
or U21970 (N_21970,N_18228,N_18880);
and U21971 (N_21971,N_17687,N_19972);
nand U21972 (N_21972,N_16309,N_17811);
nand U21973 (N_21973,N_15938,N_19269);
nand U21974 (N_21974,N_19827,N_18920);
xnor U21975 (N_21975,N_17524,N_16090);
nand U21976 (N_21976,N_18043,N_17684);
or U21977 (N_21977,N_19674,N_18803);
xor U21978 (N_21978,N_16353,N_17586);
or U21979 (N_21979,N_19839,N_15151);
xnor U21980 (N_21980,N_15602,N_15395);
xnor U21981 (N_21981,N_17838,N_15877);
nor U21982 (N_21982,N_16860,N_19125);
nand U21983 (N_21983,N_16582,N_17430);
nor U21984 (N_21984,N_17714,N_18613);
xnor U21985 (N_21985,N_18374,N_15517);
nand U21986 (N_21986,N_15061,N_16500);
and U21987 (N_21987,N_17166,N_15055);
nor U21988 (N_21988,N_17944,N_16235);
nor U21989 (N_21989,N_16566,N_19876);
and U21990 (N_21990,N_15250,N_19821);
nor U21991 (N_21991,N_18939,N_17152);
and U21992 (N_21992,N_16780,N_17690);
or U21993 (N_21993,N_18108,N_15237);
and U21994 (N_21994,N_18339,N_15163);
nor U21995 (N_21995,N_16149,N_15166);
and U21996 (N_21996,N_19374,N_16936);
or U21997 (N_21997,N_15598,N_17544);
nand U21998 (N_21998,N_17854,N_17471);
nand U21999 (N_21999,N_15480,N_18196);
and U22000 (N_22000,N_15453,N_18469);
xnor U22001 (N_22001,N_17190,N_15730);
or U22002 (N_22002,N_18883,N_15805);
and U22003 (N_22003,N_17946,N_15363);
nor U22004 (N_22004,N_16840,N_19126);
nor U22005 (N_22005,N_15698,N_17369);
xor U22006 (N_22006,N_19397,N_16965);
nor U22007 (N_22007,N_17393,N_18804);
nor U22008 (N_22008,N_18010,N_17105);
nand U22009 (N_22009,N_19772,N_16649);
or U22010 (N_22010,N_19600,N_19096);
and U22011 (N_22011,N_19548,N_18351);
nand U22012 (N_22012,N_15470,N_17759);
nand U22013 (N_22013,N_15817,N_19053);
and U22014 (N_22014,N_15228,N_16921);
xor U22015 (N_22015,N_19382,N_17464);
xnor U22016 (N_22016,N_16445,N_17495);
and U22017 (N_22017,N_17889,N_16198);
xor U22018 (N_22018,N_18580,N_17444);
or U22019 (N_22019,N_18402,N_16434);
or U22020 (N_22020,N_15978,N_18543);
xnor U22021 (N_22021,N_15684,N_17016);
or U22022 (N_22022,N_19287,N_19013);
nor U22023 (N_22023,N_16450,N_18926);
nor U22024 (N_22024,N_18448,N_15907);
nand U22025 (N_22025,N_18178,N_15174);
xor U22026 (N_22026,N_19920,N_19835);
nor U22027 (N_22027,N_17903,N_17012);
nor U22028 (N_22028,N_16464,N_15018);
and U22029 (N_22029,N_15682,N_16803);
and U22030 (N_22030,N_18588,N_19392);
nor U22031 (N_22031,N_15782,N_16163);
or U22032 (N_22032,N_17569,N_17353);
or U22033 (N_22033,N_15687,N_19031);
and U22034 (N_22034,N_18277,N_18068);
xor U22035 (N_22035,N_16466,N_15815);
xor U22036 (N_22036,N_17769,N_16234);
and U22037 (N_22037,N_18554,N_15223);
nor U22038 (N_22038,N_19662,N_19991);
xor U22039 (N_22039,N_16932,N_15046);
and U22040 (N_22040,N_19129,N_15148);
or U22041 (N_22041,N_16896,N_19473);
nor U22042 (N_22042,N_16101,N_19769);
or U22043 (N_22043,N_19234,N_15107);
xnor U22044 (N_22044,N_16736,N_15330);
or U22045 (N_22045,N_19500,N_19573);
nand U22046 (N_22046,N_17666,N_15458);
xnor U22047 (N_22047,N_19597,N_16069);
nor U22048 (N_22048,N_19406,N_16790);
or U22049 (N_22049,N_19569,N_18666);
nand U22050 (N_22050,N_18823,N_17505);
or U22051 (N_22051,N_17610,N_19006);
and U22052 (N_22052,N_15012,N_15828);
and U22053 (N_22053,N_18825,N_18135);
or U22054 (N_22054,N_18671,N_15836);
and U22055 (N_22055,N_15052,N_16829);
nand U22056 (N_22056,N_18350,N_16186);
nand U22057 (N_22057,N_18684,N_17852);
or U22058 (N_22058,N_17264,N_16555);
xnor U22059 (N_22059,N_17576,N_16039);
and U22060 (N_22060,N_19836,N_18536);
and U22061 (N_22061,N_17083,N_15493);
nand U22062 (N_22062,N_18811,N_17408);
nor U22063 (N_22063,N_17802,N_15710);
or U22064 (N_22064,N_17536,N_15440);
and U22065 (N_22065,N_15083,N_15422);
and U22066 (N_22066,N_16864,N_16580);
or U22067 (N_22067,N_17343,N_19881);
nand U22068 (N_22068,N_18404,N_17136);
xor U22069 (N_22069,N_18639,N_17097);
nor U22070 (N_22070,N_19173,N_15711);
and U22071 (N_22071,N_19819,N_18609);
nor U22072 (N_22072,N_16672,N_15019);
or U22073 (N_22073,N_17245,N_19764);
xnor U22074 (N_22074,N_19974,N_15775);
nor U22075 (N_22075,N_18837,N_19226);
nand U22076 (N_22076,N_16939,N_16208);
or U22077 (N_22077,N_15118,N_19077);
or U22078 (N_22078,N_19602,N_17211);
and U22079 (N_22079,N_17901,N_17240);
xor U22080 (N_22080,N_15985,N_17837);
and U22081 (N_22081,N_19722,N_18700);
and U22082 (N_22082,N_15943,N_17585);
or U22083 (N_22083,N_17070,N_15651);
or U22084 (N_22084,N_18679,N_18552);
nor U22085 (N_22085,N_18847,N_19200);
xor U22086 (N_22086,N_19978,N_17810);
and U22087 (N_22087,N_17917,N_15614);
and U22088 (N_22088,N_15216,N_17385);
and U22089 (N_22089,N_17820,N_17825);
nand U22090 (N_22090,N_18387,N_18727);
and U22091 (N_22091,N_17220,N_17266);
xor U22092 (N_22092,N_16457,N_18125);
and U22093 (N_22093,N_16432,N_17558);
or U22094 (N_22094,N_19941,N_17910);
and U22095 (N_22095,N_16397,N_19144);
xor U22096 (N_22096,N_17117,N_17636);
nand U22097 (N_22097,N_17379,N_17316);
or U22098 (N_22098,N_19224,N_19055);
xor U22099 (N_22099,N_17964,N_16695);
nand U22100 (N_22100,N_19904,N_15736);
xnor U22101 (N_22101,N_19431,N_15706);
xnor U22102 (N_22102,N_18816,N_15510);
nor U22103 (N_22103,N_19279,N_19467);
and U22104 (N_22104,N_18308,N_15585);
xnor U22105 (N_22105,N_16534,N_17441);
and U22106 (N_22106,N_15225,N_18628);
and U22107 (N_22107,N_17641,N_16260);
and U22108 (N_22108,N_17711,N_17237);
nor U22109 (N_22109,N_19394,N_18899);
or U22110 (N_22110,N_19734,N_16614);
nor U22111 (N_22111,N_15591,N_15101);
or U22112 (N_22112,N_16096,N_16863);
or U22113 (N_22113,N_16611,N_18306);
xnor U22114 (N_22114,N_16747,N_17391);
nor U22115 (N_22115,N_18840,N_17292);
or U22116 (N_22116,N_18561,N_19062);
or U22117 (N_22117,N_18006,N_15361);
xnor U22118 (N_22118,N_16591,N_18086);
nand U22119 (N_22119,N_18423,N_19699);
nor U22120 (N_22120,N_17335,N_15429);
nand U22121 (N_22121,N_17087,N_16680);
nand U22122 (N_22122,N_16619,N_17835);
nor U22123 (N_22123,N_16938,N_17270);
xor U22124 (N_22124,N_16296,N_15700);
nand U22125 (N_22125,N_18138,N_19110);
nor U22126 (N_22126,N_16326,N_18534);
xor U22127 (N_22127,N_16335,N_19928);
or U22128 (N_22128,N_16590,N_15658);
or U22129 (N_22129,N_18180,N_18652);
nor U22130 (N_22130,N_18487,N_19501);
or U22131 (N_22131,N_15498,N_19511);
or U22132 (N_22132,N_16557,N_15594);
or U22133 (N_22133,N_16261,N_19877);
xnor U22134 (N_22134,N_17592,N_17822);
or U22135 (N_22135,N_18324,N_16196);
nand U22136 (N_22136,N_16941,N_15109);
or U22137 (N_22137,N_19527,N_19703);
and U22138 (N_22138,N_15855,N_15845);
nor U22139 (N_22139,N_18754,N_19156);
nor U22140 (N_22140,N_18969,N_19161);
nand U22141 (N_22141,N_16447,N_19482);
xnor U22142 (N_22142,N_19312,N_16124);
and U22143 (N_22143,N_15089,N_17836);
and U22144 (N_22144,N_15923,N_15504);
and U22145 (N_22145,N_15581,N_19025);
nand U22146 (N_22146,N_18945,N_15592);
xor U22147 (N_22147,N_17555,N_16293);
nand U22148 (N_22148,N_17153,N_15818);
xnor U22149 (N_22149,N_18997,N_15620);
nor U22150 (N_22150,N_17613,N_19795);
nand U22151 (N_22151,N_18258,N_17773);
nand U22152 (N_22152,N_15667,N_15167);
and U22153 (N_22153,N_15946,N_17745);
nand U22154 (N_22154,N_19963,N_19762);
xnor U22155 (N_22155,N_15747,N_17552);
nand U22156 (N_22156,N_18810,N_15906);
nand U22157 (N_22157,N_15601,N_19155);
and U22158 (N_22158,N_19146,N_17967);
or U22159 (N_22159,N_19039,N_18916);
or U22160 (N_22160,N_17175,N_17079);
nand U22161 (N_22161,N_16558,N_16519);
nor U22162 (N_22162,N_16740,N_19711);
or U22163 (N_22163,N_17969,N_15641);
or U22164 (N_22164,N_16213,N_19109);
nor U22165 (N_22165,N_18834,N_17804);
xnor U22166 (N_22166,N_15608,N_18454);
and U22167 (N_22167,N_16658,N_19102);
or U22168 (N_22168,N_19063,N_15733);
xnor U22169 (N_22169,N_19747,N_19639);
or U22170 (N_22170,N_15553,N_18964);
or U22171 (N_22171,N_17507,N_16912);
or U22172 (N_22172,N_16043,N_15398);
and U22173 (N_22173,N_17897,N_16501);
nand U22174 (N_22174,N_16446,N_17502);
nand U22175 (N_22175,N_19732,N_17902);
nand U22176 (N_22176,N_15513,N_17839);
xor U22177 (N_22177,N_19503,N_15536);
or U22178 (N_22178,N_17120,N_16835);
nand U22179 (N_22179,N_19813,N_18708);
xor U22180 (N_22180,N_17851,N_16577);
or U22181 (N_22181,N_15382,N_18642);
xnor U22182 (N_22182,N_17145,N_15236);
nor U22183 (N_22183,N_19070,N_17388);
and U22184 (N_22184,N_18998,N_15795);
xnor U22185 (N_22185,N_17410,N_19212);
and U22186 (N_22186,N_15180,N_18515);
or U22187 (N_22187,N_18111,N_19010);
xor U22188 (N_22188,N_15500,N_18835);
xor U22189 (N_22189,N_18265,N_17345);
nor U22190 (N_22190,N_19617,N_19766);
xnor U22191 (N_22191,N_15284,N_19229);
xnor U22192 (N_22192,N_15792,N_18485);
nor U22193 (N_22193,N_15102,N_16054);
xnor U22194 (N_22194,N_19286,N_15707);
and U22195 (N_22195,N_16883,N_18396);
xnor U22196 (N_22196,N_19101,N_17174);
xor U22197 (N_22197,N_15391,N_16405);
and U22198 (N_22198,N_16246,N_18614);
or U22199 (N_22199,N_18092,N_16993);
and U22200 (N_22200,N_19427,N_15901);
and U22201 (N_22201,N_15544,N_16514);
or U22202 (N_22202,N_15300,N_16616);
xnor U22203 (N_22203,N_18796,N_15035);
and U22204 (N_22204,N_17023,N_16759);
nor U22205 (N_22205,N_19632,N_19537);
nand U22206 (N_22206,N_18035,N_18873);
or U22207 (N_22207,N_16812,N_16689);
or U22208 (N_22208,N_18576,N_18839);
nand U22209 (N_22209,N_18775,N_15234);
xnor U22210 (N_22210,N_16708,N_15697);
nand U22211 (N_22211,N_17539,N_17125);
or U22212 (N_22212,N_16980,N_18968);
or U22213 (N_22213,N_19504,N_18372);
nor U22214 (N_22214,N_15197,N_17273);
and U22215 (N_22215,N_15870,N_16392);
or U22216 (N_22216,N_17302,N_17386);
xor U22217 (N_22217,N_19884,N_17743);
and U22218 (N_22218,N_18421,N_15136);
nor U22219 (N_22219,N_15867,N_18442);
nand U22220 (N_22220,N_18001,N_19440);
or U22221 (N_22221,N_15787,N_15213);
nand U22222 (N_22222,N_18946,N_17182);
and U22223 (N_22223,N_18812,N_18440);
and U22224 (N_22224,N_17476,N_18399);
xnor U22225 (N_22225,N_16303,N_19373);
and U22226 (N_22226,N_15056,N_15449);
and U22227 (N_22227,N_19011,N_17675);
xor U22228 (N_22228,N_15970,N_16448);
nor U22229 (N_22229,N_15643,N_18394);
or U22230 (N_22230,N_15409,N_19697);
xnor U22231 (N_22231,N_18512,N_16890);
or U22232 (N_22232,N_15004,N_17506);
xor U22233 (N_22233,N_19190,N_17002);
nor U22234 (N_22234,N_16205,N_18553);
nand U22235 (N_22235,N_18426,N_16328);
and U22236 (N_22236,N_19730,N_17111);
nor U22237 (N_22237,N_18585,N_18050);
nor U22238 (N_22238,N_17361,N_16663);
xor U22239 (N_22239,N_19973,N_15039);
nand U22240 (N_22240,N_15568,N_18897);
and U22241 (N_22241,N_19729,N_16675);
nand U22242 (N_22242,N_16032,N_17692);
xnor U22243 (N_22243,N_15507,N_17339);
or U22244 (N_22244,N_19748,N_15317);
xor U22245 (N_22245,N_16062,N_15113);
xor U22246 (N_22246,N_18461,N_16080);
nand U22247 (N_22247,N_19334,N_19237);
and U22248 (N_22248,N_17768,N_15020);
xnor U22249 (N_22249,N_15821,N_15021);
nand U22250 (N_22250,N_19496,N_17776);
nor U22251 (N_22251,N_19398,N_18739);
nor U22252 (N_22252,N_16476,N_17635);
or U22253 (N_22253,N_15421,N_19044);
and U22254 (N_22254,N_17362,N_15947);
or U22255 (N_22255,N_17694,N_16756);
and U22256 (N_22256,N_17047,N_19927);
xor U22257 (N_22257,N_16158,N_19114);
nor U22258 (N_22258,N_18729,N_15384);
and U22259 (N_22259,N_17991,N_17478);
xor U22260 (N_22260,N_15082,N_19328);
nand U22261 (N_22261,N_19886,N_16606);
xor U22262 (N_22262,N_16926,N_16778);
nand U22263 (N_22263,N_16139,N_17686);
nand U22264 (N_22264,N_19938,N_16383);
or U22265 (N_22265,N_18475,N_17570);
xnor U22266 (N_22266,N_15767,N_15342);
and U22267 (N_22267,N_17378,N_15103);
or U22268 (N_22268,N_18155,N_19304);
and U22269 (N_22269,N_16674,N_17381);
nand U22270 (N_22270,N_18567,N_18358);
or U22271 (N_22271,N_15488,N_15165);
and U22272 (N_22272,N_15964,N_15008);
xnor U22273 (N_22273,N_17823,N_18721);
nand U22274 (N_22274,N_18981,N_18544);
nand U22275 (N_22275,N_15847,N_15900);
nand U22276 (N_22276,N_16762,N_16012);
or U22277 (N_22277,N_19452,N_15766);
nand U22278 (N_22278,N_19898,N_15798);
nand U22279 (N_22279,N_16375,N_16295);
xnor U22280 (N_22280,N_18511,N_17886);
nor U22281 (N_22281,N_15131,N_18093);
and U22282 (N_22282,N_16181,N_19807);
or U22283 (N_22283,N_18495,N_18113);
nor U22284 (N_22284,N_19755,N_16212);
or U22285 (N_22285,N_18573,N_15260);
and U22286 (N_22286,N_17583,N_18114);
or U22287 (N_22287,N_16739,N_18557);
or U22288 (N_22288,N_18414,N_17529);
nand U22289 (N_22289,N_17192,N_17937);
or U22290 (N_22290,N_18537,N_18790);
nand U22291 (N_22291,N_15908,N_17606);
nor U22292 (N_22292,N_15214,N_15093);
xnor U22293 (N_22293,N_16504,N_18860);
nor U22294 (N_22294,N_16839,N_17864);
nor U22295 (N_22295,N_17086,N_17841);
and U22296 (N_22296,N_18607,N_19893);
xnor U22297 (N_22297,N_16404,N_18080);
xnor U22298 (N_22298,N_17435,N_16657);
and U22299 (N_22299,N_17056,N_15175);
nor U22300 (N_22300,N_17587,N_15264);
and U22301 (N_22301,N_16754,N_16562);
or U22302 (N_22302,N_16950,N_19015);
and U22303 (N_22303,N_19996,N_19761);
or U22304 (N_22304,N_16583,N_17268);
nand U22305 (N_22305,N_15723,N_19276);
nor U22306 (N_22306,N_16741,N_19685);
nor U22307 (N_22307,N_19222,N_15849);
xnor U22308 (N_22308,N_16752,N_17198);
xnor U22309 (N_22309,N_19844,N_15338);
or U22310 (N_22310,N_19106,N_19896);
xor U22311 (N_22311,N_18468,N_15417);
nor U22312 (N_22312,N_19074,N_15235);
nor U22313 (N_22313,N_15152,N_17980);
nor U22314 (N_22314,N_15326,N_17309);
xor U22315 (N_22315,N_19288,N_15999);
and U22316 (N_22316,N_15044,N_16561);
nand U22317 (N_22317,N_15196,N_18062);
nor U22318 (N_22318,N_18612,N_17954);
or U22319 (N_22319,N_18563,N_16402);
xnor U22320 (N_22320,N_19596,N_16971);
nand U22321 (N_22321,N_18330,N_17092);
nor U22322 (N_22322,N_19284,N_15232);
or U22323 (N_22323,N_19968,N_15169);
and U22324 (N_22324,N_16345,N_18993);
nor U22325 (N_22325,N_16268,N_17396);
xnor U22326 (N_22326,N_17296,N_17627);
nor U22327 (N_22327,N_15491,N_19180);
and U22328 (N_22328,N_18715,N_17938);
and U22329 (N_22329,N_15189,N_18192);
xnor U22330 (N_22330,N_16530,N_19746);
and U22331 (N_22331,N_19885,N_19689);
or U22332 (N_22332,N_15633,N_18432);
nor U22333 (N_22333,N_17370,N_19768);
xor U22334 (N_22334,N_19594,N_18188);
nor U22335 (N_22335,N_15852,N_17565);
nor U22336 (N_22336,N_17422,N_17556);
nor U22337 (N_22337,N_19848,N_15176);
or U22338 (N_22338,N_16443,N_18732);
or U22339 (N_22339,N_18635,N_19520);
nand U22340 (N_22340,N_16368,N_18856);
xnor U22341 (N_22341,N_15246,N_19293);
and U22342 (N_22342,N_19164,N_19660);
and U22343 (N_22343,N_19863,N_17596);
xnor U22344 (N_22344,N_18513,N_15754);
xor U22345 (N_22345,N_15307,N_17095);
xor U22346 (N_22346,N_18772,N_17695);
xnor U22347 (N_22347,N_17894,N_19459);
and U22348 (N_22348,N_15979,N_15884);
xnor U22349 (N_22349,N_18975,N_17101);
nand U22350 (N_22350,N_16449,N_15595);
nor U22351 (N_22351,N_17638,N_17905);
nand U22352 (N_22352,N_15123,N_16924);
and U22353 (N_22353,N_16613,N_19549);
nand U22354 (N_22354,N_17551,N_16075);
and U22355 (N_22355,N_18269,N_17605);
and U22356 (N_22356,N_17322,N_16007);
or U22357 (N_22357,N_17178,N_15322);
nor U22358 (N_22358,N_18292,N_19525);
or U22359 (N_22359,N_19329,N_16005);
or U22360 (N_22360,N_19763,N_15164);
or U22361 (N_22361,N_17564,N_16509);
or U22362 (N_22362,N_19179,N_18669);
xor U22363 (N_22363,N_15981,N_18735);
and U22364 (N_22364,N_16953,N_16655);
nor U22365 (N_22365,N_18627,N_15848);
xnor U22366 (N_22366,N_19414,N_15203);
or U22367 (N_22367,N_18036,N_15365);
and U22368 (N_22368,N_15090,N_15354);
or U22369 (N_22369,N_19206,N_16034);
or U22370 (N_22370,N_15534,N_16117);
xor U22371 (N_22371,N_17290,N_19086);
nand U22372 (N_22372,N_19384,N_19892);
xnor U22373 (N_22373,N_16767,N_15321);
nor U22374 (N_22374,N_16087,N_17005);
or U22375 (N_22375,N_15199,N_19731);
or U22376 (N_22376,N_18027,N_19357);
xnor U22377 (N_22377,N_17922,N_17943);
nand U22378 (N_22378,N_17633,N_16394);
nor U22379 (N_22379,N_18341,N_17683);
nand U22380 (N_22380,N_18938,N_15159);
or U22381 (N_22381,N_17180,N_19861);
nor U22382 (N_22382,N_19274,N_18655);
or U22383 (N_22383,N_17816,N_18489);
nor U22384 (N_22384,N_18759,N_15376);
or U22385 (N_22385,N_19277,N_16691);
nor U22386 (N_22386,N_16157,N_16171);
or U22387 (N_22387,N_16403,N_17228);
and U22388 (N_22388,N_18985,N_16421);
and U22389 (N_22389,N_19097,N_19967);
xnor U22390 (N_22390,N_15891,N_19299);
or U22391 (N_22391,N_18755,N_19196);
nand U22392 (N_22392,N_19917,N_19072);
xor U22393 (N_22393,N_15882,N_15785);
xor U22394 (N_22394,N_17691,N_19946);
nor U22395 (N_22395,N_19219,N_19332);
or U22396 (N_22396,N_17427,N_16690);
nor U22397 (N_22397,N_19124,N_17491);
nand U22398 (N_22398,N_15085,N_17199);
xor U22399 (N_22399,N_19317,N_19514);
or U22400 (N_22400,N_19211,N_15904);
nor U22401 (N_22401,N_18893,N_19078);
or U22402 (N_22402,N_18602,N_15172);
and U22403 (N_22403,N_18570,N_18165);
and U22404 (N_22404,N_15494,N_19307);
nand U22405 (N_22405,N_17039,N_19864);
or U22406 (N_22406,N_15057,N_17652);
or U22407 (N_22407,N_16570,N_19933);
nand U22408 (N_22408,N_15672,N_19995);
or U22409 (N_22409,N_18521,N_19223);
nor U22410 (N_22410,N_18200,N_16593);
xnor U22411 (N_22411,N_17360,N_19220);
nand U22412 (N_22412,N_19385,N_18663);
or U22413 (N_22413,N_17201,N_16334);
xor U22414 (N_22414,N_15286,N_17468);
or U22415 (N_22415,N_19702,N_15184);
xor U22416 (N_22416,N_18698,N_15584);
nor U22417 (N_22417,N_17689,N_15737);
or U22418 (N_22418,N_15885,N_16773);
nor U22419 (N_22419,N_15764,N_17602);
and U22420 (N_22420,N_15944,N_16197);
xor U22421 (N_22421,N_15769,N_19484);
nor U22422 (N_22422,N_18995,N_17050);
nor U22423 (N_22423,N_16907,N_16795);
or U22424 (N_22424,N_19614,N_15025);
nand U22425 (N_22425,N_16846,N_18822);
nand U22426 (N_22426,N_18207,N_15464);
nor U22427 (N_22427,N_16215,N_15084);
or U22428 (N_22428,N_15452,N_19849);
xor U22429 (N_22429,N_17161,N_18706);
xnor U22430 (N_22430,N_19912,N_15424);
and U22431 (N_22431,N_15015,N_19036);
nand U22432 (N_22432,N_17573,N_15860);
xnor U22433 (N_22433,N_15890,N_15368);
nor U22434 (N_22434,N_18723,N_17019);
nand U22435 (N_22435,N_18917,N_17307);
xor U22436 (N_22436,N_18730,N_18752);
xnor U22437 (N_22437,N_16533,N_15208);
nor U22438 (N_22438,N_19682,N_15655);
xor U22439 (N_22439,N_17205,N_16210);
nand U22440 (N_22440,N_18783,N_18867);
nand U22441 (N_22441,N_19056,N_19545);
nand U22442 (N_22442,N_16225,N_17796);
nor U22443 (N_22443,N_19185,N_18889);
nor U22444 (N_22444,N_19788,N_19590);
or U22445 (N_22445,N_17729,N_19802);
and U22446 (N_22446,N_19621,N_19868);
xnor U22447 (N_22447,N_19777,N_16236);
nor U22448 (N_22448,N_19936,N_18296);
xor U22449 (N_22449,N_16669,N_16576);
and U22450 (N_22450,N_17331,N_15812);
nor U22451 (N_22451,N_17077,N_15293);
nand U22452 (N_22452,N_15202,N_16543);
xor U22453 (N_22453,N_18037,N_17530);
xnor U22454 (N_22454,N_16600,N_15145);
nand U22455 (N_22455,N_15971,N_15327);
xnor U22456 (N_22456,N_18242,N_15953);
nor U22457 (N_22457,N_19045,N_19887);
nor U22458 (N_22458,N_18117,N_15288);
and U22459 (N_22459,N_15738,N_16323);
and U22460 (N_22460,N_19583,N_17990);
and U22461 (N_22461,N_15367,N_18347);
and U22462 (N_22462,N_16499,N_18044);
nor U22463 (N_22463,N_15996,N_15916);
xnor U22464 (N_22464,N_16147,N_17169);
xor U22465 (N_22465,N_16853,N_18282);
and U22466 (N_22466,N_18075,N_17096);
and U22467 (N_22467,N_15423,N_15379);
nand U22468 (N_22468,N_15966,N_15806);
nor U22469 (N_22469,N_19261,N_18479);
and U22470 (N_22470,N_17970,N_16714);
nand U22471 (N_22471,N_16817,N_18624);
nand U22472 (N_22472,N_18427,N_17115);
nor U22473 (N_22473,N_15538,N_19425);
xor U22474 (N_22474,N_19779,N_19435);
and U22475 (N_22475,N_18439,N_19035);
nor U22476 (N_22476,N_15372,N_15808);
and U22477 (N_22477,N_15065,N_16882);
xor U22478 (N_22478,N_17089,N_16637);
nor U22479 (N_22479,N_15915,N_18931);
and U22480 (N_22480,N_15009,N_16988);
xnor U22481 (N_22481,N_19987,N_19018);
and U22482 (N_22482,N_18595,N_15941);
or U22483 (N_22483,N_19923,N_15394);
nor U22484 (N_22484,N_17481,N_17074);
nand U22485 (N_22485,N_16138,N_18568);
nand U22486 (N_22486,N_15627,N_18198);
xor U22487 (N_22487,N_19444,N_18564);
xor U22488 (N_22488,N_15838,N_17761);
or U22489 (N_22489,N_18749,N_18710);
nand U22490 (N_22490,N_18937,N_19743);
or U22491 (N_22491,N_17957,N_15650);
nand U22492 (N_22492,N_15789,N_15520);
and U22493 (N_22493,N_17134,N_19263);
nand U22494 (N_22494,N_15029,N_16646);
and U22495 (N_22495,N_18633,N_16761);
or U22496 (N_22496,N_16541,N_19383);
or U22497 (N_22497,N_15456,N_15209);
or U22498 (N_22498,N_17452,N_15679);
xnor U22499 (N_22499,N_16073,N_15316);
xnor U22500 (N_22500,N_18739,N_17599);
xnor U22501 (N_22501,N_17076,N_16975);
or U22502 (N_22502,N_19781,N_17828);
nor U22503 (N_22503,N_18225,N_17715);
and U22504 (N_22504,N_15072,N_19429);
and U22505 (N_22505,N_17900,N_19762);
or U22506 (N_22506,N_19600,N_17002);
nor U22507 (N_22507,N_16880,N_17105);
xor U22508 (N_22508,N_18054,N_19766);
or U22509 (N_22509,N_16670,N_19623);
xnor U22510 (N_22510,N_17320,N_15708);
or U22511 (N_22511,N_17523,N_15016);
or U22512 (N_22512,N_18015,N_16662);
nor U22513 (N_22513,N_18274,N_18224);
nand U22514 (N_22514,N_19960,N_16533);
nor U22515 (N_22515,N_16574,N_17488);
or U22516 (N_22516,N_17658,N_19133);
or U22517 (N_22517,N_18839,N_17142);
nand U22518 (N_22518,N_16864,N_15198);
nand U22519 (N_22519,N_16387,N_18843);
or U22520 (N_22520,N_18849,N_18048);
nand U22521 (N_22521,N_16037,N_19727);
nor U22522 (N_22522,N_16227,N_19259);
and U22523 (N_22523,N_18784,N_18927);
nor U22524 (N_22524,N_15361,N_16567);
xnor U22525 (N_22525,N_19280,N_17029);
nor U22526 (N_22526,N_17377,N_17252);
nand U22527 (N_22527,N_16879,N_17769);
nand U22528 (N_22528,N_16516,N_18530);
and U22529 (N_22529,N_18902,N_19605);
and U22530 (N_22530,N_19446,N_16839);
nor U22531 (N_22531,N_18989,N_19773);
or U22532 (N_22532,N_16327,N_17982);
xor U22533 (N_22533,N_18854,N_16538);
and U22534 (N_22534,N_15556,N_19184);
xnor U22535 (N_22535,N_15458,N_16072);
xor U22536 (N_22536,N_16267,N_17815);
xnor U22537 (N_22537,N_15997,N_17097);
and U22538 (N_22538,N_15349,N_17678);
xor U22539 (N_22539,N_19857,N_19145);
and U22540 (N_22540,N_16966,N_19790);
xnor U22541 (N_22541,N_17022,N_18350);
or U22542 (N_22542,N_15649,N_19310);
xor U22543 (N_22543,N_18860,N_17473);
and U22544 (N_22544,N_18245,N_19267);
and U22545 (N_22545,N_18721,N_17316);
and U22546 (N_22546,N_15809,N_16443);
xor U22547 (N_22547,N_18286,N_16513);
or U22548 (N_22548,N_18735,N_18601);
nor U22549 (N_22549,N_15128,N_17207);
nor U22550 (N_22550,N_18742,N_16534);
xor U22551 (N_22551,N_19866,N_15467);
or U22552 (N_22552,N_19323,N_19375);
or U22553 (N_22553,N_19611,N_18836);
nor U22554 (N_22554,N_17410,N_19909);
nor U22555 (N_22555,N_19344,N_19981);
nand U22556 (N_22556,N_16075,N_18163);
and U22557 (N_22557,N_18481,N_19977);
xnor U22558 (N_22558,N_17114,N_18214);
xnor U22559 (N_22559,N_15081,N_19991);
nor U22560 (N_22560,N_18530,N_15589);
nand U22561 (N_22561,N_18523,N_15423);
xnor U22562 (N_22562,N_18820,N_17330);
nand U22563 (N_22563,N_15771,N_16510);
xor U22564 (N_22564,N_18369,N_16841);
and U22565 (N_22565,N_17677,N_19828);
xor U22566 (N_22566,N_17691,N_16465);
xor U22567 (N_22567,N_19135,N_18367);
and U22568 (N_22568,N_16685,N_17261);
nand U22569 (N_22569,N_16195,N_18606);
or U22570 (N_22570,N_15984,N_19667);
or U22571 (N_22571,N_17009,N_16638);
nor U22572 (N_22572,N_17070,N_18004);
or U22573 (N_22573,N_17717,N_16005);
nand U22574 (N_22574,N_17355,N_18694);
nor U22575 (N_22575,N_19552,N_17174);
and U22576 (N_22576,N_18455,N_17964);
and U22577 (N_22577,N_15300,N_17009);
and U22578 (N_22578,N_15585,N_17302);
and U22579 (N_22579,N_18728,N_19035);
xnor U22580 (N_22580,N_15160,N_16230);
or U22581 (N_22581,N_17634,N_16910);
xor U22582 (N_22582,N_18797,N_17833);
or U22583 (N_22583,N_15165,N_18768);
nand U22584 (N_22584,N_16210,N_15415);
and U22585 (N_22585,N_15878,N_15799);
xnor U22586 (N_22586,N_16955,N_16451);
or U22587 (N_22587,N_15533,N_17837);
nand U22588 (N_22588,N_16098,N_16531);
xnor U22589 (N_22589,N_15970,N_18183);
nand U22590 (N_22590,N_16283,N_16080);
xor U22591 (N_22591,N_17029,N_15849);
nand U22592 (N_22592,N_17103,N_16516);
nand U22593 (N_22593,N_17694,N_19323);
xnor U22594 (N_22594,N_15568,N_15870);
and U22595 (N_22595,N_16618,N_19369);
nor U22596 (N_22596,N_18248,N_19026);
and U22597 (N_22597,N_15676,N_18443);
or U22598 (N_22598,N_19987,N_16200);
xor U22599 (N_22599,N_18715,N_17218);
and U22600 (N_22600,N_19310,N_17229);
and U22601 (N_22601,N_15871,N_16786);
xor U22602 (N_22602,N_18635,N_18322);
xnor U22603 (N_22603,N_15003,N_18770);
xor U22604 (N_22604,N_15759,N_16262);
or U22605 (N_22605,N_15948,N_18965);
nor U22606 (N_22606,N_17768,N_19945);
xor U22607 (N_22607,N_19278,N_17267);
or U22608 (N_22608,N_15913,N_19633);
nor U22609 (N_22609,N_17059,N_16674);
nor U22610 (N_22610,N_17568,N_15482);
nand U22611 (N_22611,N_17416,N_19247);
nand U22612 (N_22612,N_17478,N_17280);
xor U22613 (N_22613,N_17889,N_17943);
xnor U22614 (N_22614,N_15648,N_16653);
nor U22615 (N_22615,N_18599,N_17951);
xor U22616 (N_22616,N_16219,N_19060);
and U22617 (N_22617,N_19523,N_19413);
nor U22618 (N_22618,N_17080,N_18008);
nand U22619 (N_22619,N_17671,N_18505);
nand U22620 (N_22620,N_17451,N_15293);
nor U22621 (N_22621,N_18023,N_17471);
nand U22622 (N_22622,N_19716,N_15500);
nand U22623 (N_22623,N_18059,N_19014);
nand U22624 (N_22624,N_19265,N_16741);
nand U22625 (N_22625,N_16209,N_16037);
nor U22626 (N_22626,N_16767,N_17925);
and U22627 (N_22627,N_15987,N_15642);
or U22628 (N_22628,N_16471,N_19265);
or U22629 (N_22629,N_16272,N_17774);
nor U22630 (N_22630,N_19730,N_18221);
or U22631 (N_22631,N_15321,N_17269);
xnor U22632 (N_22632,N_15481,N_15929);
nand U22633 (N_22633,N_16155,N_17363);
nand U22634 (N_22634,N_17181,N_18239);
or U22635 (N_22635,N_19989,N_19076);
and U22636 (N_22636,N_17459,N_15946);
nor U22637 (N_22637,N_16014,N_15974);
or U22638 (N_22638,N_17045,N_18482);
nand U22639 (N_22639,N_18549,N_17833);
or U22640 (N_22640,N_17839,N_16552);
nand U22641 (N_22641,N_19493,N_18469);
nor U22642 (N_22642,N_17721,N_19497);
nor U22643 (N_22643,N_15370,N_18838);
nor U22644 (N_22644,N_17456,N_17467);
nand U22645 (N_22645,N_15552,N_16382);
nor U22646 (N_22646,N_15343,N_16242);
xor U22647 (N_22647,N_17493,N_18594);
nor U22648 (N_22648,N_15954,N_16938);
nor U22649 (N_22649,N_15695,N_15719);
nor U22650 (N_22650,N_16757,N_19450);
nor U22651 (N_22651,N_15300,N_19042);
nand U22652 (N_22652,N_18081,N_16572);
nor U22653 (N_22653,N_16266,N_15817);
and U22654 (N_22654,N_16805,N_19472);
xnor U22655 (N_22655,N_19033,N_15312);
nand U22656 (N_22656,N_19082,N_18106);
xor U22657 (N_22657,N_19489,N_15366);
xor U22658 (N_22658,N_16956,N_19430);
or U22659 (N_22659,N_19793,N_15903);
and U22660 (N_22660,N_17170,N_17529);
and U22661 (N_22661,N_15991,N_16373);
and U22662 (N_22662,N_17961,N_19111);
nor U22663 (N_22663,N_17504,N_15711);
and U22664 (N_22664,N_15242,N_17011);
nor U22665 (N_22665,N_15676,N_17955);
and U22666 (N_22666,N_15320,N_16199);
and U22667 (N_22667,N_15057,N_17107);
nor U22668 (N_22668,N_15803,N_18004);
and U22669 (N_22669,N_17521,N_18912);
xor U22670 (N_22670,N_19225,N_19970);
or U22671 (N_22671,N_15523,N_15415);
nor U22672 (N_22672,N_17475,N_18914);
or U22673 (N_22673,N_16597,N_15983);
or U22674 (N_22674,N_17651,N_17821);
and U22675 (N_22675,N_16966,N_18582);
nor U22676 (N_22676,N_15568,N_15032);
or U22677 (N_22677,N_19827,N_17903);
nor U22678 (N_22678,N_18673,N_15604);
nand U22679 (N_22679,N_16446,N_16462);
xnor U22680 (N_22680,N_17953,N_16496);
or U22681 (N_22681,N_16197,N_17590);
nor U22682 (N_22682,N_15797,N_19533);
nor U22683 (N_22683,N_15182,N_16694);
or U22684 (N_22684,N_18339,N_18884);
or U22685 (N_22685,N_15421,N_15633);
nand U22686 (N_22686,N_16969,N_17874);
nor U22687 (N_22687,N_15444,N_16683);
xnor U22688 (N_22688,N_16181,N_17791);
and U22689 (N_22689,N_16487,N_17328);
or U22690 (N_22690,N_16754,N_16568);
nand U22691 (N_22691,N_15850,N_16209);
and U22692 (N_22692,N_18913,N_17790);
and U22693 (N_22693,N_17045,N_19220);
xnor U22694 (N_22694,N_19885,N_19263);
or U22695 (N_22695,N_15376,N_16807);
nor U22696 (N_22696,N_15670,N_15079);
xor U22697 (N_22697,N_19357,N_19008);
and U22698 (N_22698,N_16513,N_19629);
or U22699 (N_22699,N_16748,N_16345);
and U22700 (N_22700,N_18198,N_19360);
and U22701 (N_22701,N_16025,N_19307);
or U22702 (N_22702,N_15196,N_19773);
nand U22703 (N_22703,N_16001,N_18109);
and U22704 (N_22704,N_16321,N_17526);
nand U22705 (N_22705,N_18885,N_16701);
or U22706 (N_22706,N_15948,N_18155);
xnor U22707 (N_22707,N_17411,N_15952);
xnor U22708 (N_22708,N_15207,N_18064);
nor U22709 (N_22709,N_17963,N_19879);
and U22710 (N_22710,N_15033,N_15500);
or U22711 (N_22711,N_15296,N_18787);
nor U22712 (N_22712,N_19214,N_18578);
nand U22713 (N_22713,N_19385,N_19130);
nand U22714 (N_22714,N_19189,N_18802);
nand U22715 (N_22715,N_17538,N_19275);
nor U22716 (N_22716,N_18825,N_18056);
or U22717 (N_22717,N_17799,N_15231);
xnor U22718 (N_22718,N_18194,N_19830);
nand U22719 (N_22719,N_19544,N_17882);
nand U22720 (N_22720,N_16262,N_15838);
or U22721 (N_22721,N_16305,N_16616);
nor U22722 (N_22722,N_16709,N_16809);
or U22723 (N_22723,N_15172,N_17087);
nor U22724 (N_22724,N_15908,N_16316);
nor U22725 (N_22725,N_19033,N_18033);
nand U22726 (N_22726,N_16716,N_19752);
and U22727 (N_22727,N_18250,N_19170);
xor U22728 (N_22728,N_18360,N_18468);
or U22729 (N_22729,N_19626,N_19789);
or U22730 (N_22730,N_15776,N_19288);
xor U22731 (N_22731,N_16165,N_17587);
nor U22732 (N_22732,N_19895,N_19957);
nor U22733 (N_22733,N_15639,N_16015);
or U22734 (N_22734,N_17137,N_17433);
and U22735 (N_22735,N_17665,N_15929);
nor U22736 (N_22736,N_19280,N_19429);
or U22737 (N_22737,N_19095,N_18553);
nor U22738 (N_22738,N_18419,N_17594);
nand U22739 (N_22739,N_16400,N_19418);
and U22740 (N_22740,N_17020,N_17817);
and U22741 (N_22741,N_17086,N_16464);
nor U22742 (N_22742,N_17599,N_18027);
and U22743 (N_22743,N_16895,N_15230);
xor U22744 (N_22744,N_16057,N_15608);
xor U22745 (N_22745,N_17310,N_19616);
or U22746 (N_22746,N_19280,N_19004);
or U22747 (N_22747,N_18325,N_15478);
or U22748 (N_22748,N_15598,N_16698);
or U22749 (N_22749,N_16837,N_18623);
and U22750 (N_22750,N_15865,N_15212);
and U22751 (N_22751,N_16170,N_19845);
xor U22752 (N_22752,N_19705,N_17564);
and U22753 (N_22753,N_19751,N_16052);
and U22754 (N_22754,N_16463,N_16104);
or U22755 (N_22755,N_18769,N_15541);
xnor U22756 (N_22756,N_18385,N_18485);
nor U22757 (N_22757,N_18585,N_17187);
and U22758 (N_22758,N_18968,N_15777);
nor U22759 (N_22759,N_19631,N_15513);
nand U22760 (N_22760,N_18376,N_15089);
nand U22761 (N_22761,N_15294,N_17924);
and U22762 (N_22762,N_17620,N_15312);
nand U22763 (N_22763,N_19741,N_17100);
or U22764 (N_22764,N_16229,N_17689);
nand U22765 (N_22765,N_15910,N_17718);
xnor U22766 (N_22766,N_16962,N_16207);
xor U22767 (N_22767,N_19792,N_16413);
or U22768 (N_22768,N_18497,N_17956);
xnor U22769 (N_22769,N_16720,N_16230);
nand U22770 (N_22770,N_19808,N_17853);
xnor U22771 (N_22771,N_18220,N_17837);
nor U22772 (N_22772,N_19023,N_17899);
nor U22773 (N_22773,N_15856,N_17938);
or U22774 (N_22774,N_16956,N_16253);
or U22775 (N_22775,N_15515,N_15852);
nor U22776 (N_22776,N_19345,N_18162);
nand U22777 (N_22777,N_18502,N_18298);
and U22778 (N_22778,N_15979,N_18183);
xnor U22779 (N_22779,N_18266,N_19205);
xnor U22780 (N_22780,N_16006,N_19048);
xnor U22781 (N_22781,N_15227,N_16204);
nand U22782 (N_22782,N_17066,N_18472);
nand U22783 (N_22783,N_17002,N_17825);
nor U22784 (N_22784,N_18622,N_18866);
and U22785 (N_22785,N_15864,N_18150);
nor U22786 (N_22786,N_15450,N_18835);
nand U22787 (N_22787,N_15022,N_19216);
nand U22788 (N_22788,N_16656,N_18559);
or U22789 (N_22789,N_15312,N_16460);
nor U22790 (N_22790,N_19470,N_18089);
or U22791 (N_22791,N_16219,N_16995);
xor U22792 (N_22792,N_17063,N_15239);
or U22793 (N_22793,N_16215,N_17621);
nor U22794 (N_22794,N_15497,N_16478);
nand U22795 (N_22795,N_15503,N_16423);
nand U22796 (N_22796,N_16300,N_15554);
or U22797 (N_22797,N_17485,N_17397);
and U22798 (N_22798,N_16829,N_16913);
or U22799 (N_22799,N_17144,N_17866);
and U22800 (N_22800,N_19849,N_17883);
nand U22801 (N_22801,N_15189,N_16512);
xnor U22802 (N_22802,N_15478,N_15750);
and U22803 (N_22803,N_16570,N_17400);
or U22804 (N_22804,N_19840,N_15062);
nand U22805 (N_22805,N_19472,N_17411);
nor U22806 (N_22806,N_16411,N_18784);
nand U22807 (N_22807,N_15988,N_19562);
and U22808 (N_22808,N_15434,N_18553);
nor U22809 (N_22809,N_18890,N_18732);
xnor U22810 (N_22810,N_16526,N_16997);
or U22811 (N_22811,N_16933,N_18478);
nor U22812 (N_22812,N_17313,N_19552);
nor U22813 (N_22813,N_15850,N_17976);
and U22814 (N_22814,N_19099,N_18031);
nor U22815 (N_22815,N_19982,N_19123);
nand U22816 (N_22816,N_15501,N_18993);
or U22817 (N_22817,N_18372,N_18320);
and U22818 (N_22818,N_19173,N_15723);
or U22819 (N_22819,N_16542,N_17903);
or U22820 (N_22820,N_19594,N_18663);
nand U22821 (N_22821,N_16406,N_19922);
or U22822 (N_22822,N_16946,N_15569);
nand U22823 (N_22823,N_17849,N_17156);
xor U22824 (N_22824,N_18159,N_15755);
or U22825 (N_22825,N_19006,N_16691);
and U22826 (N_22826,N_19920,N_15907);
xor U22827 (N_22827,N_19369,N_15217);
xor U22828 (N_22828,N_15282,N_18118);
or U22829 (N_22829,N_19360,N_15777);
and U22830 (N_22830,N_16341,N_16312);
or U22831 (N_22831,N_16980,N_16414);
nand U22832 (N_22832,N_16094,N_15790);
or U22833 (N_22833,N_18299,N_17100);
nor U22834 (N_22834,N_17506,N_19154);
xor U22835 (N_22835,N_18626,N_18705);
and U22836 (N_22836,N_15838,N_19681);
xnor U22837 (N_22837,N_17817,N_17175);
xnor U22838 (N_22838,N_19845,N_18646);
xor U22839 (N_22839,N_18235,N_17029);
and U22840 (N_22840,N_18647,N_16080);
or U22841 (N_22841,N_15750,N_15819);
nor U22842 (N_22842,N_16993,N_15829);
nand U22843 (N_22843,N_15325,N_19049);
or U22844 (N_22844,N_15015,N_19607);
nor U22845 (N_22845,N_15656,N_18903);
xor U22846 (N_22846,N_17323,N_16722);
and U22847 (N_22847,N_15357,N_16477);
nor U22848 (N_22848,N_17216,N_15390);
nor U22849 (N_22849,N_18923,N_18461);
and U22850 (N_22850,N_18150,N_15484);
or U22851 (N_22851,N_18700,N_17588);
xnor U22852 (N_22852,N_16117,N_19208);
and U22853 (N_22853,N_16915,N_18956);
and U22854 (N_22854,N_17470,N_15960);
or U22855 (N_22855,N_15046,N_16484);
and U22856 (N_22856,N_17310,N_18825);
and U22857 (N_22857,N_19483,N_16726);
xor U22858 (N_22858,N_19245,N_18622);
nor U22859 (N_22859,N_15903,N_17609);
xnor U22860 (N_22860,N_17846,N_19862);
and U22861 (N_22861,N_16116,N_17986);
and U22862 (N_22862,N_19748,N_19382);
xnor U22863 (N_22863,N_15912,N_15108);
xnor U22864 (N_22864,N_17763,N_19553);
xnor U22865 (N_22865,N_17325,N_18332);
or U22866 (N_22866,N_15519,N_15607);
xnor U22867 (N_22867,N_17663,N_18227);
or U22868 (N_22868,N_19006,N_18861);
and U22869 (N_22869,N_17531,N_16044);
nor U22870 (N_22870,N_18849,N_15259);
and U22871 (N_22871,N_18023,N_19325);
or U22872 (N_22872,N_19954,N_18301);
or U22873 (N_22873,N_18102,N_19765);
or U22874 (N_22874,N_15946,N_18726);
and U22875 (N_22875,N_17856,N_16430);
nor U22876 (N_22876,N_19169,N_18262);
or U22877 (N_22877,N_19668,N_18620);
nor U22878 (N_22878,N_15617,N_16715);
nor U22879 (N_22879,N_16473,N_19236);
and U22880 (N_22880,N_16210,N_15623);
nand U22881 (N_22881,N_19173,N_17998);
nor U22882 (N_22882,N_19254,N_18698);
nand U22883 (N_22883,N_18301,N_16191);
nor U22884 (N_22884,N_16163,N_15385);
or U22885 (N_22885,N_15548,N_17216);
and U22886 (N_22886,N_19586,N_18848);
nor U22887 (N_22887,N_15927,N_16556);
and U22888 (N_22888,N_15475,N_19640);
nand U22889 (N_22889,N_19590,N_15005);
and U22890 (N_22890,N_19445,N_19999);
and U22891 (N_22891,N_17959,N_15087);
xnor U22892 (N_22892,N_16019,N_19044);
or U22893 (N_22893,N_17053,N_15385);
xor U22894 (N_22894,N_17468,N_16479);
and U22895 (N_22895,N_19700,N_16523);
nand U22896 (N_22896,N_17560,N_17030);
and U22897 (N_22897,N_18547,N_19811);
or U22898 (N_22898,N_17110,N_17502);
nand U22899 (N_22899,N_18520,N_18979);
and U22900 (N_22900,N_16053,N_19510);
nor U22901 (N_22901,N_16589,N_19479);
xor U22902 (N_22902,N_15583,N_17020);
nor U22903 (N_22903,N_17147,N_15696);
xor U22904 (N_22904,N_15344,N_17826);
nand U22905 (N_22905,N_16697,N_17423);
and U22906 (N_22906,N_19292,N_19934);
and U22907 (N_22907,N_17788,N_19898);
or U22908 (N_22908,N_18012,N_17034);
or U22909 (N_22909,N_19945,N_15392);
nor U22910 (N_22910,N_17207,N_16369);
nand U22911 (N_22911,N_15611,N_17947);
nand U22912 (N_22912,N_16030,N_18277);
or U22913 (N_22913,N_16377,N_19594);
nor U22914 (N_22914,N_19889,N_18487);
or U22915 (N_22915,N_18593,N_19088);
nand U22916 (N_22916,N_15939,N_16349);
and U22917 (N_22917,N_19632,N_18301);
and U22918 (N_22918,N_19425,N_18009);
xnor U22919 (N_22919,N_16487,N_15185);
xnor U22920 (N_22920,N_16823,N_19769);
xor U22921 (N_22921,N_19646,N_17826);
xnor U22922 (N_22922,N_18080,N_19233);
nand U22923 (N_22923,N_16538,N_18808);
and U22924 (N_22924,N_17466,N_15722);
nor U22925 (N_22925,N_18641,N_16365);
and U22926 (N_22926,N_17041,N_18677);
nor U22927 (N_22927,N_15676,N_19762);
or U22928 (N_22928,N_17505,N_15264);
xnor U22929 (N_22929,N_15127,N_17625);
or U22930 (N_22930,N_16825,N_16787);
nand U22931 (N_22931,N_16161,N_15982);
nor U22932 (N_22932,N_17523,N_16661);
or U22933 (N_22933,N_19527,N_17951);
or U22934 (N_22934,N_19302,N_17804);
nand U22935 (N_22935,N_16354,N_15504);
nor U22936 (N_22936,N_15942,N_17801);
nor U22937 (N_22937,N_17492,N_17062);
and U22938 (N_22938,N_19220,N_15116);
nor U22939 (N_22939,N_16589,N_17883);
nor U22940 (N_22940,N_16145,N_16484);
or U22941 (N_22941,N_19938,N_19453);
nand U22942 (N_22942,N_19438,N_19566);
nand U22943 (N_22943,N_18812,N_15998);
nand U22944 (N_22944,N_17291,N_16081);
or U22945 (N_22945,N_18209,N_16905);
or U22946 (N_22946,N_15682,N_19036);
nand U22947 (N_22947,N_18922,N_19846);
or U22948 (N_22948,N_19792,N_16786);
nand U22949 (N_22949,N_17874,N_17274);
nand U22950 (N_22950,N_18730,N_16952);
nor U22951 (N_22951,N_17977,N_16380);
nand U22952 (N_22952,N_17974,N_18793);
xnor U22953 (N_22953,N_19629,N_16795);
xnor U22954 (N_22954,N_19897,N_19131);
nand U22955 (N_22955,N_15274,N_19332);
xnor U22956 (N_22956,N_18442,N_15170);
nor U22957 (N_22957,N_15850,N_18957);
or U22958 (N_22958,N_17133,N_17968);
nor U22959 (N_22959,N_19367,N_15110);
nand U22960 (N_22960,N_17859,N_18055);
nand U22961 (N_22961,N_15832,N_17424);
or U22962 (N_22962,N_19408,N_18049);
xnor U22963 (N_22963,N_19093,N_16664);
xor U22964 (N_22964,N_15647,N_18462);
nor U22965 (N_22965,N_19951,N_16353);
and U22966 (N_22966,N_18292,N_19127);
or U22967 (N_22967,N_19288,N_17528);
and U22968 (N_22968,N_19591,N_19079);
xnor U22969 (N_22969,N_15640,N_19956);
or U22970 (N_22970,N_16016,N_18386);
and U22971 (N_22971,N_19840,N_18658);
and U22972 (N_22972,N_15827,N_19281);
xor U22973 (N_22973,N_18871,N_17077);
or U22974 (N_22974,N_17309,N_19318);
xor U22975 (N_22975,N_15521,N_18550);
or U22976 (N_22976,N_16494,N_15502);
nor U22977 (N_22977,N_19582,N_19443);
and U22978 (N_22978,N_18282,N_15274);
nand U22979 (N_22979,N_15811,N_16570);
xnor U22980 (N_22980,N_18688,N_16807);
or U22981 (N_22981,N_17726,N_16703);
nand U22982 (N_22982,N_17868,N_15076);
or U22983 (N_22983,N_18127,N_15414);
and U22984 (N_22984,N_19505,N_19563);
xor U22985 (N_22985,N_19643,N_18348);
or U22986 (N_22986,N_18442,N_16720);
xor U22987 (N_22987,N_17655,N_16641);
nand U22988 (N_22988,N_15758,N_18718);
nand U22989 (N_22989,N_18789,N_19086);
xor U22990 (N_22990,N_17210,N_18444);
xnor U22991 (N_22991,N_19468,N_16792);
and U22992 (N_22992,N_18003,N_17857);
or U22993 (N_22993,N_16544,N_15386);
or U22994 (N_22994,N_15086,N_16085);
xnor U22995 (N_22995,N_17171,N_18317);
nand U22996 (N_22996,N_16347,N_17453);
nor U22997 (N_22997,N_15829,N_15114);
xnor U22998 (N_22998,N_18158,N_16462);
xnor U22999 (N_22999,N_19585,N_16929);
nand U23000 (N_23000,N_19401,N_18755);
nand U23001 (N_23001,N_17083,N_17557);
or U23002 (N_23002,N_17592,N_17958);
xnor U23003 (N_23003,N_15311,N_15043);
or U23004 (N_23004,N_19529,N_18953);
xor U23005 (N_23005,N_19166,N_18753);
nand U23006 (N_23006,N_18429,N_18290);
and U23007 (N_23007,N_17018,N_16253);
or U23008 (N_23008,N_15091,N_16946);
nand U23009 (N_23009,N_15406,N_15237);
xnor U23010 (N_23010,N_17826,N_15900);
nand U23011 (N_23011,N_15468,N_18098);
nor U23012 (N_23012,N_17647,N_16051);
nand U23013 (N_23013,N_18848,N_19302);
and U23014 (N_23014,N_15728,N_17632);
nor U23015 (N_23015,N_18311,N_15601);
and U23016 (N_23016,N_19595,N_19548);
nor U23017 (N_23017,N_19195,N_15707);
xor U23018 (N_23018,N_17499,N_17278);
or U23019 (N_23019,N_19340,N_18239);
nand U23020 (N_23020,N_17918,N_15262);
xor U23021 (N_23021,N_18698,N_19113);
xor U23022 (N_23022,N_16887,N_18516);
or U23023 (N_23023,N_16800,N_17727);
or U23024 (N_23024,N_19938,N_17426);
or U23025 (N_23025,N_18579,N_15650);
and U23026 (N_23026,N_18208,N_17535);
or U23027 (N_23027,N_17334,N_18420);
nor U23028 (N_23028,N_17348,N_15325);
xor U23029 (N_23029,N_17915,N_15354);
nand U23030 (N_23030,N_16263,N_15550);
or U23031 (N_23031,N_17260,N_19376);
nand U23032 (N_23032,N_18007,N_19949);
nand U23033 (N_23033,N_18121,N_17120);
xor U23034 (N_23034,N_17441,N_18719);
or U23035 (N_23035,N_16007,N_17734);
or U23036 (N_23036,N_16436,N_15286);
xnor U23037 (N_23037,N_16170,N_16385);
or U23038 (N_23038,N_18894,N_18604);
or U23039 (N_23039,N_17365,N_16184);
or U23040 (N_23040,N_19686,N_19814);
or U23041 (N_23041,N_19453,N_18815);
xor U23042 (N_23042,N_17433,N_15633);
nand U23043 (N_23043,N_17022,N_19434);
nor U23044 (N_23044,N_19337,N_17255);
or U23045 (N_23045,N_15468,N_15697);
and U23046 (N_23046,N_16320,N_18932);
or U23047 (N_23047,N_15013,N_16866);
xor U23048 (N_23048,N_19644,N_19232);
or U23049 (N_23049,N_17310,N_19409);
and U23050 (N_23050,N_15341,N_19852);
nor U23051 (N_23051,N_16374,N_19370);
nand U23052 (N_23052,N_17049,N_18238);
xnor U23053 (N_23053,N_18842,N_17697);
nor U23054 (N_23054,N_18243,N_16731);
nor U23055 (N_23055,N_15457,N_15464);
and U23056 (N_23056,N_19749,N_18050);
or U23057 (N_23057,N_17318,N_19548);
nand U23058 (N_23058,N_19817,N_16693);
nor U23059 (N_23059,N_17095,N_18569);
nor U23060 (N_23060,N_16384,N_15944);
or U23061 (N_23061,N_15281,N_17544);
or U23062 (N_23062,N_16696,N_15063);
xnor U23063 (N_23063,N_17744,N_17148);
nor U23064 (N_23064,N_18540,N_18811);
nor U23065 (N_23065,N_16105,N_19183);
and U23066 (N_23066,N_15858,N_19377);
and U23067 (N_23067,N_15058,N_19881);
nand U23068 (N_23068,N_15038,N_15758);
and U23069 (N_23069,N_15461,N_16836);
xor U23070 (N_23070,N_16314,N_15192);
or U23071 (N_23071,N_15155,N_16356);
or U23072 (N_23072,N_18646,N_18547);
nor U23073 (N_23073,N_17295,N_19024);
nand U23074 (N_23074,N_17651,N_17841);
nor U23075 (N_23075,N_16784,N_18784);
or U23076 (N_23076,N_19530,N_17876);
and U23077 (N_23077,N_18173,N_18530);
and U23078 (N_23078,N_16519,N_17369);
or U23079 (N_23079,N_15245,N_19748);
nand U23080 (N_23080,N_16998,N_19725);
nor U23081 (N_23081,N_16351,N_15806);
or U23082 (N_23082,N_17873,N_15005);
xnor U23083 (N_23083,N_19433,N_15107);
xnor U23084 (N_23084,N_16351,N_17576);
nand U23085 (N_23085,N_18520,N_19781);
xnor U23086 (N_23086,N_19093,N_16421);
nor U23087 (N_23087,N_17728,N_19705);
xor U23088 (N_23088,N_19228,N_18301);
and U23089 (N_23089,N_15508,N_16116);
xnor U23090 (N_23090,N_15487,N_18674);
and U23091 (N_23091,N_19362,N_17167);
nor U23092 (N_23092,N_17454,N_16689);
nand U23093 (N_23093,N_16480,N_15547);
or U23094 (N_23094,N_18357,N_15377);
or U23095 (N_23095,N_16926,N_15117);
nor U23096 (N_23096,N_18955,N_16114);
and U23097 (N_23097,N_17729,N_19303);
xor U23098 (N_23098,N_19738,N_18383);
xor U23099 (N_23099,N_15744,N_16374);
nor U23100 (N_23100,N_19690,N_17583);
and U23101 (N_23101,N_19574,N_15367);
nor U23102 (N_23102,N_15142,N_17320);
nand U23103 (N_23103,N_15336,N_15094);
xnor U23104 (N_23104,N_17356,N_17677);
nand U23105 (N_23105,N_16172,N_18761);
and U23106 (N_23106,N_18159,N_16469);
or U23107 (N_23107,N_15361,N_19220);
nor U23108 (N_23108,N_16577,N_17545);
or U23109 (N_23109,N_16761,N_19003);
or U23110 (N_23110,N_19991,N_15365);
xnor U23111 (N_23111,N_19203,N_17223);
or U23112 (N_23112,N_15014,N_16191);
or U23113 (N_23113,N_16787,N_17085);
and U23114 (N_23114,N_19954,N_15423);
xor U23115 (N_23115,N_16910,N_15051);
xnor U23116 (N_23116,N_17293,N_16554);
or U23117 (N_23117,N_18730,N_17168);
xnor U23118 (N_23118,N_17152,N_19634);
xnor U23119 (N_23119,N_16564,N_16247);
nor U23120 (N_23120,N_15906,N_16574);
nand U23121 (N_23121,N_18666,N_17388);
and U23122 (N_23122,N_17948,N_17769);
nor U23123 (N_23123,N_18536,N_19855);
nand U23124 (N_23124,N_18670,N_17213);
nand U23125 (N_23125,N_19372,N_17185);
nand U23126 (N_23126,N_15724,N_19444);
or U23127 (N_23127,N_16630,N_19885);
xor U23128 (N_23128,N_18022,N_15326);
xnor U23129 (N_23129,N_17545,N_19425);
nor U23130 (N_23130,N_18895,N_15391);
and U23131 (N_23131,N_16631,N_15631);
xor U23132 (N_23132,N_19442,N_18330);
xor U23133 (N_23133,N_19299,N_15182);
nand U23134 (N_23134,N_15753,N_19609);
nor U23135 (N_23135,N_18961,N_19938);
and U23136 (N_23136,N_16394,N_19917);
nor U23137 (N_23137,N_15740,N_16411);
nor U23138 (N_23138,N_15036,N_18979);
xnor U23139 (N_23139,N_17064,N_18825);
or U23140 (N_23140,N_19376,N_19662);
or U23141 (N_23141,N_16050,N_15393);
or U23142 (N_23142,N_19783,N_17591);
nor U23143 (N_23143,N_17471,N_19240);
nand U23144 (N_23144,N_16953,N_15822);
nand U23145 (N_23145,N_16506,N_19680);
nor U23146 (N_23146,N_16597,N_15615);
xor U23147 (N_23147,N_19826,N_19629);
or U23148 (N_23148,N_18480,N_17330);
or U23149 (N_23149,N_19580,N_18148);
nand U23150 (N_23150,N_18996,N_17385);
nand U23151 (N_23151,N_16349,N_19443);
nand U23152 (N_23152,N_15233,N_15875);
and U23153 (N_23153,N_18320,N_15046);
xnor U23154 (N_23154,N_16153,N_18648);
or U23155 (N_23155,N_15847,N_19722);
and U23156 (N_23156,N_15452,N_16000);
xor U23157 (N_23157,N_17011,N_16913);
and U23158 (N_23158,N_19462,N_16049);
xor U23159 (N_23159,N_15638,N_17021);
nor U23160 (N_23160,N_19235,N_15435);
nor U23161 (N_23161,N_18668,N_16258);
or U23162 (N_23162,N_17292,N_17364);
xnor U23163 (N_23163,N_16577,N_18065);
nand U23164 (N_23164,N_15434,N_15712);
xor U23165 (N_23165,N_19263,N_16671);
xnor U23166 (N_23166,N_18735,N_17256);
nor U23167 (N_23167,N_19660,N_15044);
or U23168 (N_23168,N_16092,N_16499);
nand U23169 (N_23169,N_15506,N_15450);
nor U23170 (N_23170,N_16080,N_18722);
or U23171 (N_23171,N_16793,N_15140);
nand U23172 (N_23172,N_16092,N_16717);
and U23173 (N_23173,N_18201,N_17876);
and U23174 (N_23174,N_16939,N_16655);
nand U23175 (N_23175,N_19703,N_16266);
nand U23176 (N_23176,N_18045,N_17736);
or U23177 (N_23177,N_17552,N_17874);
nor U23178 (N_23178,N_19759,N_15630);
nand U23179 (N_23179,N_18579,N_16934);
nor U23180 (N_23180,N_19426,N_19582);
xor U23181 (N_23181,N_17942,N_18542);
or U23182 (N_23182,N_18099,N_18372);
nand U23183 (N_23183,N_18795,N_18965);
xor U23184 (N_23184,N_15143,N_15665);
nand U23185 (N_23185,N_16507,N_15444);
nand U23186 (N_23186,N_16101,N_19992);
nand U23187 (N_23187,N_15314,N_19309);
xnor U23188 (N_23188,N_17413,N_16220);
and U23189 (N_23189,N_15847,N_18790);
nand U23190 (N_23190,N_15979,N_15434);
and U23191 (N_23191,N_15823,N_16817);
xnor U23192 (N_23192,N_17561,N_19724);
and U23193 (N_23193,N_17340,N_18540);
or U23194 (N_23194,N_16215,N_18498);
xnor U23195 (N_23195,N_18493,N_18445);
nor U23196 (N_23196,N_15098,N_17607);
and U23197 (N_23197,N_15841,N_18810);
xnor U23198 (N_23198,N_15034,N_16116);
nand U23199 (N_23199,N_15312,N_15576);
or U23200 (N_23200,N_19686,N_15472);
nand U23201 (N_23201,N_15490,N_16075);
xor U23202 (N_23202,N_15733,N_18315);
and U23203 (N_23203,N_19721,N_18000);
nand U23204 (N_23204,N_18521,N_17033);
nor U23205 (N_23205,N_19741,N_17066);
or U23206 (N_23206,N_17853,N_16532);
and U23207 (N_23207,N_18832,N_16800);
nor U23208 (N_23208,N_16272,N_17959);
nor U23209 (N_23209,N_17548,N_17002);
and U23210 (N_23210,N_18015,N_18610);
or U23211 (N_23211,N_15475,N_16747);
or U23212 (N_23212,N_15458,N_18444);
or U23213 (N_23213,N_19022,N_15556);
and U23214 (N_23214,N_15695,N_17867);
xnor U23215 (N_23215,N_15256,N_16783);
nor U23216 (N_23216,N_19160,N_17684);
or U23217 (N_23217,N_18128,N_15690);
or U23218 (N_23218,N_16400,N_17911);
nand U23219 (N_23219,N_17224,N_16001);
or U23220 (N_23220,N_18921,N_19120);
xnor U23221 (N_23221,N_16151,N_17010);
and U23222 (N_23222,N_18766,N_17700);
nor U23223 (N_23223,N_16210,N_15978);
nand U23224 (N_23224,N_17357,N_16628);
and U23225 (N_23225,N_19005,N_19371);
and U23226 (N_23226,N_16513,N_16658);
xor U23227 (N_23227,N_16252,N_19572);
and U23228 (N_23228,N_15521,N_18976);
and U23229 (N_23229,N_15891,N_17560);
nand U23230 (N_23230,N_19121,N_16401);
xnor U23231 (N_23231,N_19672,N_15485);
nand U23232 (N_23232,N_15846,N_15969);
xor U23233 (N_23233,N_17128,N_16110);
nor U23234 (N_23234,N_19818,N_18867);
xnor U23235 (N_23235,N_15361,N_19986);
or U23236 (N_23236,N_19829,N_17839);
nand U23237 (N_23237,N_15642,N_15927);
or U23238 (N_23238,N_15759,N_17168);
xnor U23239 (N_23239,N_16258,N_19447);
nor U23240 (N_23240,N_17818,N_19055);
and U23241 (N_23241,N_18536,N_19423);
nand U23242 (N_23242,N_18320,N_16247);
nand U23243 (N_23243,N_19824,N_15903);
or U23244 (N_23244,N_17290,N_18946);
and U23245 (N_23245,N_18094,N_18631);
or U23246 (N_23246,N_19765,N_16650);
or U23247 (N_23247,N_19763,N_18705);
xnor U23248 (N_23248,N_18618,N_18918);
nand U23249 (N_23249,N_15213,N_17322);
xor U23250 (N_23250,N_15604,N_18852);
xor U23251 (N_23251,N_16128,N_17803);
nor U23252 (N_23252,N_16385,N_18105);
nor U23253 (N_23253,N_15537,N_18162);
xor U23254 (N_23254,N_16627,N_18434);
nor U23255 (N_23255,N_19562,N_19202);
xor U23256 (N_23256,N_17889,N_16762);
nor U23257 (N_23257,N_17605,N_17444);
nor U23258 (N_23258,N_18371,N_19161);
and U23259 (N_23259,N_17321,N_18229);
and U23260 (N_23260,N_19742,N_15839);
xor U23261 (N_23261,N_19470,N_15370);
xor U23262 (N_23262,N_16293,N_15739);
nor U23263 (N_23263,N_19578,N_18949);
nor U23264 (N_23264,N_16073,N_17768);
or U23265 (N_23265,N_15715,N_17287);
nand U23266 (N_23266,N_16552,N_17946);
xnor U23267 (N_23267,N_19389,N_15639);
nand U23268 (N_23268,N_17064,N_15421);
or U23269 (N_23269,N_19164,N_16771);
or U23270 (N_23270,N_18154,N_18658);
and U23271 (N_23271,N_15925,N_17704);
and U23272 (N_23272,N_17293,N_16974);
nand U23273 (N_23273,N_17694,N_17295);
nor U23274 (N_23274,N_18838,N_18084);
or U23275 (N_23275,N_19072,N_15928);
nand U23276 (N_23276,N_17092,N_18024);
nor U23277 (N_23277,N_16184,N_16710);
or U23278 (N_23278,N_18758,N_15659);
nor U23279 (N_23279,N_19684,N_16259);
nand U23280 (N_23280,N_19003,N_19798);
or U23281 (N_23281,N_19330,N_16081);
xor U23282 (N_23282,N_19431,N_19560);
nor U23283 (N_23283,N_18260,N_15853);
or U23284 (N_23284,N_16841,N_18357);
nor U23285 (N_23285,N_16739,N_16762);
nor U23286 (N_23286,N_17616,N_17489);
and U23287 (N_23287,N_16067,N_19238);
and U23288 (N_23288,N_18405,N_16161);
or U23289 (N_23289,N_19476,N_15782);
xor U23290 (N_23290,N_17087,N_16428);
and U23291 (N_23291,N_19461,N_16695);
and U23292 (N_23292,N_16520,N_19657);
or U23293 (N_23293,N_19596,N_18086);
or U23294 (N_23294,N_15276,N_19526);
xnor U23295 (N_23295,N_16530,N_15459);
xnor U23296 (N_23296,N_19448,N_16648);
xor U23297 (N_23297,N_15598,N_17204);
nand U23298 (N_23298,N_19547,N_18770);
nor U23299 (N_23299,N_19517,N_15220);
and U23300 (N_23300,N_17567,N_16581);
or U23301 (N_23301,N_16196,N_17452);
or U23302 (N_23302,N_18558,N_17399);
or U23303 (N_23303,N_15514,N_19415);
nand U23304 (N_23304,N_18748,N_18479);
nor U23305 (N_23305,N_16871,N_15652);
xor U23306 (N_23306,N_18945,N_17152);
or U23307 (N_23307,N_16950,N_16731);
and U23308 (N_23308,N_19249,N_15152);
and U23309 (N_23309,N_15033,N_15503);
nand U23310 (N_23310,N_17002,N_15223);
or U23311 (N_23311,N_17850,N_17048);
nand U23312 (N_23312,N_18170,N_19172);
xor U23313 (N_23313,N_17308,N_17699);
xor U23314 (N_23314,N_17457,N_19224);
nor U23315 (N_23315,N_15828,N_18154);
nor U23316 (N_23316,N_19314,N_15973);
nand U23317 (N_23317,N_15112,N_18233);
and U23318 (N_23318,N_19587,N_19314);
or U23319 (N_23319,N_16285,N_15161);
xor U23320 (N_23320,N_15380,N_19911);
nor U23321 (N_23321,N_15670,N_18916);
nor U23322 (N_23322,N_18257,N_19334);
and U23323 (N_23323,N_18542,N_15910);
nor U23324 (N_23324,N_19192,N_17627);
and U23325 (N_23325,N_16581,N_18009);
nand U23326 (N_23326,N_19312,N_19921);
nand U23327 (N_23327,N_18624,N_19128);
or U23328 (N_23328,N_16949,N_15379);
and U23329 (N_23329,N_18609,N_16246);
xnor U23330 (N_23330,N_15623,N_18569);
nand U23331 (N_23331,N_18505,N_15697);
xnor U23332 (N_23332,N_18242,N_16258);
nor U23333 (N_23333,N_16258,N_17731);
and U23334 (N_23334,N_16451,N_17113);
nor U23335 (N_23335,N_16493,N_19619);
xor U23336 (N_23336,N_18880,N_18117);
and U23337 (N_23337,N_16216,N_19922);
and U23338 (N_23338,N_19270,N_18306);
nand U23339 (N_23339,N_19197,N_15920);
or U23340 (N_23340,N_18774,N_15723);
and U23341 (N_23341,N_19070,N_18843);
or U23342 (N_23342,N_15313,N_16028);
nand U23343 (N_23343,N_19711,N_16539);
nand U23344 (N_23344,N_17958,N_18921);
and U23345 (N_23345,N_16179,N_17821);
or U23346 (N_23346,N_17117,N_19580);
nand U23347 (N_23347,N_18732,N_18752);
nand U23348 (N_23348,N_19533,N_18491);
xnor U23349 (N_23349,N_18075,N_18229);
xor U23350 (N_23350,N_18031,N_19833);
and U23351 (N_23351,N_17370,N_16933);
nor U23352 (N_23352,N_19113,N_16044);
nand U23353 (N_23353,N_17627,N_19831);
or U23354 (N_23354,N_16249,N_17310);
nand U23355 (N_23355,N_19409,N_17482);
nor U23356 (N_23356,N_19901,N_17922);
or U23357 (N_23357,N_17756,N_16067);
nor U23358 (N_23358,N_15392,N_17352);
nand U23359 (N_23359,N_18837,N_17514);
nor U23360 (N_23360,N_16893,N_16516);
nand U23361 (N_23361,N_17022,N_18667);
nand U23362 (N_23362,N_16568,N_18084);
and U23363 (N_23363,N_16758,N_17038);
nor U23364 (N_23364,N_16157,N_15987);
xnor U23365 (N_23365,N_18986,N_16888);
and U23366 (N_23366,N_17219,N_17155);
or U23367 (N_23367,N_16955,N_15817);
nor U23368 (N_23368,N_17832,N_18363);
or U23369 (N_23369,N_17975,N_18022);
nand U23370 (N_23370,N_17595,N_16202);
xnor U23371 (N_23371,N_19173,N_16677);
and U23372 (N_23372,N_17540,N_17338);
and U23373 (N_23373,N_16424,N_16984);
or U23374 (N_23374,N_16257,N_16083);
xnor U23375 (N_23375,N_15378,N_19722);
and U23376 (N_23376,N_19853,N_16916);
and U23377 (N_23377,N_19957,N_15664);
nand U23378 (N_23378,N_19606,N_19753);
xnor U23379 (N_23379,N_16070,N_18502);
and U23380 (N_23380,N_19159,N_19838);
nand U23381 (N_23381,N_18110,N_18538);
nand U23382 (N_23382,N_17766,N_19107);
and U23383 (N_23383,N_17583,N_15332);
nand U23384 (N_23384,N_19381,N_16843);
nor U23385 (N_23385,N_15861,N_18306);
and U23386 (N_23386,N_19389,N_16508);
xnor U23387 (N_23387,N_16702,N_18359);
xnor U23388 (N_23388,N_15499,N_17421);
or U23389 (N_23389,N_16330,N_15403);
or U23390 (N_23390,N_18549,N_19729);
and U23391 (N_23391,N_19238,N_15619);
or U23392 (N_23392,N_17569,N_17640);
nand U23393 (N_23393,N_19550,N_18923);
nor U23394 (N_23394,N_16582,N_17482);
and U23395 (N_23395,N_18121,N_18599);
nor U23396 (N_23396,N_18529,N_18359);
xnor U23397 (N_23397,N_15749,N_15208);
or U23398 (N_23398,N_15485,N_16251);
xnor U23399 (N_23399,N_15899,N_16363);
nand U23400 (N_23400,N_18015,N_17160);
nand U23401 (N_23401,N_19882,N_18736);
and U23402 (N_23402,N_17333,N_17439);
and U23403 (N_23403,N_17940,N_18189);
nand U23404 (N_23404,N_15988,N_16480);
nand U23405 (N_23405,N_15844,N_15896);
and U23406 (N_23406,N_16929,N_16139);
and U23407 (N_23407,N_17293,N_18958);
nor U23408 (N_23408,N_17903,N_16337);
nand U23409 (N_23409,N_19168,N_16310);
and U23410 (N_23410,N_15659,N_16444);
xor U23411 (N_23411,N_17226,N_19995);
nand U23412 (N_23412,N_17900,N_18716);
xor U23413 (N_23413,N_16922,N_16740);
nor U23414 (N_23414,N_15111,N_16943);
or U23415 (N_23415,N_15482,N_15374);
nor U23416 (N_23416,N_19281,N_17862);
and U23417 (N_23417,N_18950,N_17451);
nor U23418 (N_23418,N_16934,N_18633);
and U23419 (N_23419,N_17458,N_19218);
and U23420 (N_23420,N_16291,N_19768);
or U23421 (N_23421,N_17834,N_18102);
nor U23422 (N_23422,N_15444,N_18519);
nor U23423 (N_23423,N_19788,N_18324);
nand U23424 (N_23424,N_19921,N_17106);
nand U23425 (N_23425,N_15528,N_18126);
nand U23426 (N_23426,N_18322,N_19886);
xor U23427 (N_23427,N_18066,N_17902);
nand U23428 (N_23428,N_15526,N_16286);
xnor U23429 (N_23429,N_16790,N_17314);
xor U23430 (N_23430,N_15264,N_16283);
nand U23431 (N_23431,N_17707,N_17082);
or U23432 (N_23432,N_19722,N_18468);
or U23433 (N_23433,N_16635,N_15785);
and U23434 (N_23434,N_17887,N_16357);
nand U23435 (N_23435,N_16084,N_18653);
nor U23436 (N_23436,N_18094,N_19964);
nor U23437 (N_23437,N_18769,N_15849);
xor U23438 (N_23438,N_16257,N_19370);
or U23439 (N_23439,N_18274,N_15779);
xnor U23440 (N_23440,N_16509,N_16467);
nor U23441 (N_23441,N_18718,N_18175);
or U23442 (N_23442,N_15857,N_16763);
or U23443 (N_23443,N_16698,N_17651);
or U23444 (N_23444,N_15448,N_15596);
and U23445 (N_23445,N_15289,N_15771);
nand U23446 (N_23446,N_18171,N_17460);
xor U23447 (N_23447,N_15482,N_19397);
xor U23448 (N_23448,N_17697,N_18358);
nor U23449 (N_23449,N_15014,N_17783);
xnor U23450 (N_23450,N_17730,N_18300);
xor U23451 (N_23451,N_17403,N_16772);
and U23452 (N_23452,N_19213,N_18238);
xor U23453 (N_23453,N_18414,N_17781);
nor U23454 (N_23454,N_15485,N_15008);
or U23455 (N_23455,N_19273,N_19855);
nand U23456 (N_23456,N_17736,N_18404);
and U23457 (N_23457,N_15606,N_16980);
xnor U23458 (N_23458,N_16565,N_18865);
xor U23459 (N_23459,N_17608,N_17029);
nor U23460 (N_23460,N_18448,N_17697);
and U23461 (N_23461,N_17395,N_16630);
and U23462 (N_23462,N_18352,N_19397);
or U23463 (N_23463,N_19941,N_15178);
or U23464 (N_23464,N_19527,N_17850);
nor U23465 (N_23465,N_18119,N_17507);
and U23466 (N_23466,N_18830,N_16481);
nor U23467 (N_23467,N_17699,N_15513);
xor U23468 (N_23468,N_18247,N_19032);
xnor U23469 (N_23469,N_18653,N_17459);
nor U23470 (N_23470,N_16381,N_19222);
and U23471 (N_23471,N_15132,N_15861);
or U23472 (N_23472,N_15117,N_16549);
and U23473 (N_23473,N_18230,N_18365);
or U23474 (N_23474,N_15053,N_19817);
and U23475 (N_23475,N_16500,N_19734);
or U23476 (N_23476,N_17460,N_19982);
and U23477 (N_23477,N_18431,N_17665);
or U23478 (N_23478,N_16194,N_17992);
nand U23479 (N_23479,N_18331,N_19472);
and U23480 (N_23480,N_18216,N_19969);
nand U23481 (N_23481,N_17398,N_19214);
and U23482 (N_23482,N_16579,N_18139);
nor U23483 (N_23483,N_18772,N_18103);
or U23484 (N_23484,N_18448,N_15406);
nand U23485 (N_23485,N_15787,N_17691);
xnor U23486 (N_23486,N_19021,N_15016);
and U23487 (N_23487,N_18872,N_18170);
and U23488 (N_23488,N_18585,N_18762);
and U23489 (N_23489,N_17705,N_18588);
nor U23490 (N_23490,N_17686,N_16134);
xnor U23491 (N_23491,N_17613,N_18526);
xor U23492 (N_23492,N_15222,N_17104);
and U23493 (N_23493,N_18336,N_19021);
and U23494 (N_23494,N_15436,N_18922);
nand U23495 (N_23495,N_17075,N_18473);
xnor U23496 (N_23496,N_15356,N_19966);
or U23497 (N_23497,N_17080,N_18730);
nor U23498 (N_23498,N_19141,N_16036);
xnor U23499 (N_23499,N_18918,N_17787);
and U23500 (N_23500,N_17223,N_18047);
nor U23501 (N_23501,N_15622,N_16416);
nand U23502 (N_23502,N_18600,N_15439);
nor U23503 (N_23503,N_15736,N_18161);
xnor U23504 (N_23504,N_17834,N_18960);
nand U23505 (N_23505,N_15208,N_17912);
xnor U23506 (N_23506,N_15169,N_19317);
or U23507 (N_23507,N_19362,N_15862);
nor U23508 (N_23508,N_18973,N_15884);
or U23509 (N_23509,N_15357,N_19493);
nor U23510 (N_23510,N_16132,N_18378);
and U23511 (N_23511,N_18241,N_16173);
nor U23512 (N_23512,N_17746,N_15246);
xor U23513 (N_23513,N_18717,N_15655);
nor U23514 (N_23514,N_18124,N_17129);
nand U23515 (N_23515,N_17848,N_15491);
nor U23516 (N_23516,N_17959,N_17909);
or U23517 (N_23517,N_17038,N_19415);
and U23518 (N_23518,N_17301,N_16621);
xor U23519 (N_23519,N_18970,N_15034);
or U23520 (N_23520,N_18428,N_18152);
or U23521 (N_23521,N_16186,N_15494);
and U23522 (N_23522,N_18987,N_17119);
nand U23523 (N_23523,N_16086,N_15804);
nor U23524 (N_23524,N_15071,N_19057);
xor U23525 (N_23525,N_18313,N_17905);
or U23526 (N_23526,N_16503,N_19644);
xor U23527 (N_23527,N_17822,N_17264);
nand U23528 (N_23528,N_19058,N_19705);
and U23529 (N_23529,N_17016,N_15060);
nor U23530 (N_23530,N_16348,N_17410);
and U23531 (N_23531,N_15662,N_15796);
and U23532 (N_23532,N_16566,N_18809);
or U23533 (N_23533,N_17269,N_15250);
nand U23534 (N_23534,N_15566,N_16764);
nand U23535 (N_23535,N_15184,N_18995);
nor U23536 (N_23536,N_16519,N_15553);
nor U23537 (N_23537,N_19160,N_18400);
and U23538 (N_23538,N_19239,N_18706);
nand U23539 (N_23539,N_19395,N_19541);
nor U23540 (N_23540,N_18550,N_16902);
nor U23541 (N_23541,N_16072,N_16297);
nor U23542 (N_23542,N_19933,N_16443);
xnor U23543 (N_23543,N_19278,N_16948);
nor U23544 (N_23544,N_19065,N_17721);
xnor U23545 (N_23545,N_19407,N_19940);
or U23546 (N_23546,N_16660,N_16768);
nand U23547 (N_23547,N_18130,N_15454);
xnor U23548 (N_23548,N_19238,N_19909);
or U23549 (N_23549,N_16484,N_16535);
and U23550 (N_23550,N_15761,N_18585);
or U23551 (N_23551,N_19660,N_15577);
xor U23552 (N_23552,N_19374,N_18023);
xnor U23553 (N_23553,N_19661,N_16087);
xor U23554 (N_23554,N_17931,N_17566);
nor U23555 (N_23555,N_16753,N_19016);
and U23556 (N_23556,N_16982,N_15747);
and U23557 (N_23557,N_18107,N_19134);
and U23558 (N_23558,N_17292,N_18647);
nor U23559 (N_23559,N_16584,N_17220);
and U23560 (N_23560,N_17919,N_16772);
nor U23561 (N_23561,N_17423,N_19898);
xor U23562 (N_23562,N_15625,N_15859);
nand U23563 (N_23563,N_15648,N_15579);
nor U23564 (N_23564,N_16416,N_17598);
nand U23565 (N_23565,N_15087,N_15151);
or U23566 (N_23566,N_18427,N_18203);
xor U23567 (N_23567,N_19391,N_17512);
xnor U23568 (N_23568,N_17863,N_15544);
or U23569 (N_23569,N_19886,N_19342);
nand U23570 (N_23570,N_18303,N_16709);
or U23571 (N_23571,N_17969,N_18268);
xnor U23572 (N_23572,N_19673,N_17781);
nand U23573 (N_23573,N_19720,N_17629);
xor U23574 (N_23574,N_15360,N_17823);
nand U23575 (N_23575,N_16675,N_16001);
or U23576 (N_23576,N_19306,N_16539);
nor U23577 (N_23577,N_17381,N_19491);
and U23578 (N_23578,N_15300,N_15782);
nor U23579 (N_23579,N_19809,N_16972);
nor U23580 (N_23580,N_16859,N_16329);
nand U23581 (N_23581,N_15338,N_15171);
and U23582 (N_23582,N_19196,N_18676);
nor U23583 (N_23583,N_19952,N_18708);
xnor U23584 (N_23584,N_17767,N_15452);
or U23585 (N_23585,N_17774,N_15000);
nand U23586 (N_23586,N_17079,N_17649);
or U23587 (N_23587,N_16126,N_19795);
or U23588 (N_23588,N_16173,N_17471);
nor U23589 (N_23589,N_18708,N_16692);
nor U23590 (N_23590,N_16203,N_17696);
nand U23591 (N_23591,N_17300,N_16583);
nand U23592 (N_23592,N_15756,N_16465);
nor U23593 (N_23593,N_15109,N_16664);
nand U23594 (N_23594,N_15945,N_16222);
nand U23595 (N_23595,N_15489,N_18263);
nand U23596 (N_23596,N_15297,N_16547);
or U23597 (N_23597,N_17020,N_19402);
and U23598 (N_23598,N_18656,N_17449);
or U23599 (N_23599,N_18739,N_15241);
and U23600 (N_23600,N_18276,N_18459);
or U23601 (N_23601,N_18901,N_18560);
and U23602 (N_23602,N_19242,N_15100);
nand U23603 (N_23603,N_19531,N_19304);
xnor U23604 (N_23604,N_17631,N_17572);
and U23605 (N_23605,N_19454,N_17407);
or U23606 (N_23606,N_16927,N_18723);
xnor U23607 (N_23607,N_15525,N_15980);
xor U23608 (N_23608,N_19608,N_16146);
and U23609 (N_23609,N_16229,N_16215);
nor U23610 (N_23610,N_15394,N_18772);
nand U23611 (N_23611,N_18990,N_15036);
nor U23612 (N_23612,N_15850,N_16538);
or U23613 (N_23613,N_15394,N_19428);
or U23614 (N_23614,N_16161,N_18492);
nand U23615 (N_23615,N_15381,N_15717);
nand U23616 (N_23616,N_18798,N_17464);
nor U23617 (N_23617,N_18086,N_18056);
and U23618 (N_23618,N_17770,N_18351);
nand U23619 (N_23619,N_15223,N_16035);
nor U23620 (N_23620,N_18153,N_16260);
nand U23621 (N_23621,N_18078,N_19835);
and U23622 (N_23622,N_16585,N_16530);
nand U23623 (N_23623,N_16418,N_15079);
nor U23624 (N_23624,N_16435,N_18712);
and U23625 (N_23625,N_16835,N_15127);
and U23626 (N_23626,N_17296,N_18578);
or U23627 (N_23627,N_15783,N_15096);
or U23628 (N_23628,N_17217,N_18311);
nand U23629 (N_23629,N_17783,N_18454);
or U23630 (N_23630,N_19138,N_16575);
or U23631 (N_23631,N_16676,N_19384);
xor U23632 (N_23632,N_19935,N_17355);
or U23633 (N_23633,N_19904,N_16963);
nor U23634 (N_23634,N_16951,N_15116);
nor U23635 (N_23635,N_15731,N_16261);
or U23636 (N_23636,N_19675,N_15619);
nand U23637 (N_23637,N_19991,N_19914);
xor U23638 (N_23638,N_18291,N_19259);
or U23639 (N_23639,N_16851,N_18935);
xor U23640 (N_23640,N_16562,N_18487);
and U23641 (N_23641,N_15203,N_16103);
nand U23642 (N_23642,N_17430,N_16169);
xor U23643 (N_23643,N_19340,N_15586);
nor U23644 (N_23644,N_17357,N_16405);
and U23645 (N_23645,N_19309,N_15710);
nor U23646 (N_23646,N_15131,N_18825);
xnor U23647 (N_23647,N_19542,N_15586);
and U23648 (N_23648,N_16340,N_18590);
xor U23649 (N_23649,N_18444,N_17000);
or U23650 (N_23650,N_16731,N_18927);
and U23651 (N_23651,N_16417,N_17459);
or U23652 (N_23652,N_15288,N_18486);
nand U23653 (N_23653,N_17884,N_15621);
or U23654 (N_23654,N_19297,N_15911);
nor U23655 (N_23655,N_15467,N_17287);
or U23656 (N_23656,N_17247,N_18999);
xor U23657 (N_23657,N_17252,N_15663);
and U23658 (N_23658,N_19005,N_19464);
xnor U23659 (N_23659,N_18536,N_19863);
or U23660 (N_23660,N_16423,N_17777);
and U23661 (N_23661,N_17401,N_17918);
nor U23662 (N_23662,N_19896,N_17751);
xnor U23663 (N_23663,N_15631,N_19465);
nand U23664 (N_23664,N_19875,N_15866);
or U23665 (N_23665,N_15433,N_15849);
nor U23666 (N_23666,N_19650,N_16461);
xor U23667 (N_23667,N_16219,N_15945);
or U23668 (N_23668,N_15316,N_19622);
nand U23669 (N_23669,N_19783,N_16239);
or U23670 (N_23670,N_17379,N_15406);
nor U23671 (N_23671,N_18642,N_17319);
and U23672 (N_23672,N_19079,N_19866);
and U23673 (N_23673,N_17251,N_17154);
nand U23674 (N_23674,N_17528,N_16385);
or U23675 (N_23675,N_15776,N_19619);
or U23676 (N_23676,N_15565,N_18133);
xor U23677 (N_23677,N_15500,N_19423);
or U23678 (N_23678,N_18629,N_16346);
xor U23679 (N_23679,N_18042,N_19800);
nor U23680 (N_23680,N_18141,N_16293);
xnor U23681 (N_23681,N_17221,N_18759);
and U23682 (N_23682,N_18662,N_18844);
or U23683 (N_23683,N_16895,N_15198);
nor U23684 (N_23684,N_19513,N_15214);
xnor U23685 (N_23685,N_17800,N_17711);
or U23686 (N_23686,N_16077,N_17854);
nor U23687 (N_23687,N_19607,N_19870);
or U23688 (N_23688,N_17168,N_18192);
or U23689 (N_23689,N_15483,N_17706);
nand U23690 (N_23690,N_16611,N_19198);
nand U23691 (N_23691,N_19876,N_17004);
and U23692 (N_23692,N_19085,N_16164);
or U23693 (N_23693,N_18494,N_18634);
nand U23694 (N_23694,N_19957,N_17734);
and U23695 (N_23695,N_15498,N_19419);
xor U23696 (N_23696,N_19950,N_18213);
nor U23697 (N_23697,N_18369,N_18991);
xor U23698 (N_23698,N_19785,N_15313);
nor U23699 (N_23699,N_17456,N_17847);
xor U23700 (N_23700,N_16994,N_19003);
or U23701 (N_23701,N_17084,N_17402);
nor U23702 (N_23702,N_17084,N_17665);
and U23703 (N_23703,N_15231,N_19333);
nor U23704 (N_23704,N_15036,N_15128);
xnor U23705 (N_23705,N_15406,N_15348);
nor U23706 (N_23706,N_18533,N_16928);
and U23707 (N_23707,N_16357,N_15476);
nor U23708 (N_23708,N_18355,N_16862);
and U23709 (N_23709,N_15542,N_15732);
or U23710 (N_23710,N_19488,N_18538);
and U23711 (N_23711,N_19637,N_16842);
or U23712 (N_23712,N_17480,N_17473);
nor U23713 (N_23713,N_19671,N_19167);
nand U23714 (N_23714,N_19354,N_17137);
or U23715 (N_23715,N_19253,N_17241);
nor U23716 (N_23716,N_19141,N_18090);
xnor U23717 (N_23717,N_15875,N_19852);
and U23718 (N_23718,N_17949,N_18951);
or U23719 (N_23719,N_19117,N_16550);
xnor U23720 (N_23720,N_18426,N_16064);
xnor U23721 (N_23721,N_16219,N_18611);
nor U23722 (N_23722,N_18059,N_15143);
and U23723 (N_23723,N_16852,N_19203);
nor U23724 (N_23724,N_18200,N_18032);
or U23725 (N_23725,N_15959,N_19476);
and U23726 (N_23726,N_19124,N_17063);
or U23727 (N_23727,N_18353,N_16847);
and U23728 (N_23728,N_19176,N_15529);
and U23729 (N_23729,N_16940,N_17620);
nor U23730 (N_23730,N_16277,N_19369);
nand U23731 (N_23731,N_19713,N_16132);
xnor U23732 (N_23732,N_17260,N_19884);
or U23733 (N_23733,N_19218,N_18898);
nand U23734 (N_23734,N_17710,N_17169);
or U23735 (N_23735,N_16141,N_18132);
xnor U23736 (N_23736,N_19871,N_19851);
and U23737 (N_23737,N_15929,N_16780);
or U23738 (N_23738,N_15963,N_15960);
nor U23739 (N_23739,N_18502,N_15823);
nand U23740 (N_23740,N_18313,N_17926);
or U23741 (N_23741,N_17894,N_16707);
nor U23742 (N_23742,N_17235,N_17936);
xnor U23743 (N_23743,N_19104,N_16539);
or U23744 (N_23744,N_17318,N_17018);
xnor U23745 (N_23745,N_19896,N_19381);
nor U23746 (N_23746,N_15048,N_17855);
and U23747 (N_23747,N_18251,N_15934);
xnor U23748 (N_23748,N_17258,N_16051);
nand U23749 (N_23749,N_17252,N_18163);
nand U23750 (N_23750,N_15974,N_19816);
xnor U23751 (N_23751,N_19566,N_19123);
and U23752 (N_23752,N_18780,N_16846);
nor U23753 (N_23753,N_15739,N_17613);
nand U23754 (N_23754,N_16697,N_16288);
nor U23755 (N_23755,N_17175,N_17931);
nor U23756 (N_23756,N_16693,N_18576);
and U23757 (N_23757,N_18242,N_17743);
or U23758 (N_23758,N_17855,N_16806);
nand U23759 (N_23759,N_19130,N_18829);
and U23760 (N_23760,N_18088,N_17827);
nor U23761 (N_23761,N_17833,N_16847);
xor U23762 (N_23762,N_15871,N_15750);
nand U23763 (N_23763,N_18754,N_16433);
nand U23764 (N_23764,N_18098,N_15747);
nor U23765 (N_23765,N_15166,N_16717);
nor U23766 (N_23766,N_17260,N_16068);
nor U23767 (N_23767,N_19348,N_18907);
nand U23768 (N_23768,N_19495,N_17955);
nand U23769 (N_23769,N_18175,N_18512);
or U23770 (N_23770,N_15825,N_17877);
or U23771 (N_23771,N_19133,N_16914);
nand U23772 (N_23772,N_18691,N_17657);
xnor U23773 (N_23773,N_15288,N_16156);
and U23774 (N_23774,N_16348,N_18598);
nand U23775 (N_23775,N_15111,N_16564);
and U23776 (N_23776,N_18496,N_16477);
and U23777 (N_23777,N_18571,N_17500);
xor U23778 (N_23778,N_15858,N_19883);
nand U23779 (N_23779,N_15094,N_16928);
xnor U23780 (N_23780,N_19151,N_17595);
or U23781 (N_23781,N_15250,N_16140);
and U23782 (N_23782,N_15835,N_15262);
nor U23783 (N_23783,N_18609,N_18077);
nor U23784 (N_23784,N_16384,N_18352);
nor U23785 (N_23785,N_17044,N_18924);
or U23786 (N_23786,N_17634,N_17098);
and U23787 (N_23787,N_18040,N_15108);
nor U23788 (N_23788,N_18692,N_17146);
or U23789 (N_23789,N_19149,N_18680);
xnor U23790 (N_23790,N_17066,N_16804);
xor U23791 (N_23791,N_18243,N_15120);
xnor U23792 (N_23792,N_15533,N_19710);
nor U23793 (N_23793,N_16905,N_18258);
nor U23794 (N_23794,N_15905,N_16679);
and U23795 (N_23795,N_15220,N_17006);
nor U23796 (N_23796,N_15264,N_16923);
nor U23797 (N_23797,N_17415,N_15608);
xnor U23798 (N_23798,N_17800,N_19490);
nor U23799 (N_23799,N_18715,N_17085);
and U23800 (N_23800,N_17832,N_17342);
and U23801 (N_23801,N_17619,N_17163);
or U23802 (N_23802,N_18732,N_16370);
and U23803 (N_23803,N_17224,N_19797);
or U23804 (N_23804,N_17685,N_17159);
or U23805 (N_23805,N_19215,N_19952);
or U23806 (N_23806,N_15469,N_17560);
nor U23807 (N_23807,N_17081,N_19511);
and U23808 (N_23808,N_19303,N_19146);
xor U23809 (N_23809,N_19117,N_18130);
and U23810 (N_23810,N_16511,N_15138);
nor U23811 (N_23811,N_17771,N_17834);
nand U23812 (N_23812,N_16984,N_15190);
and U23813 (N_23813,N_15821,N_17714);
nor U23814 (N_23814,N_18577,N_17042);
nor U23815 (N_23815,N_19165,N_18078);
or U23816 (N_23816,N_15749,N_19385);
nor U23817 (N_23817,N_18093,N_19876);
nor U23818 (N_23818,N_18292,N_18897);
xnor U23819 (N_23819,N_19456,N_16212);
and U23820 (N_23820,N_18621,N_16683);
nor U23821 (N_23821,N_18381,N_18624);
nand U23822 (N_23822,N_18398,N_17032);
or U23823 (N_23823,N_19843,N_17160);
nor U23824 (N_23824,N_16890,N_18995);
xnor U23825 (N_23825,N_19831,N_16289);
and U23826 (N_23826,N_19731,N_17744);
nor U23827 (N_23827,N_19962,N_18525);
nor U23828 (N_23828,N_16350,N_16018);
nand U23829 (N_23829,N_15201,N_17018);
nand U23830 (N_23830,N_18897,N_19279);
xor U23831 (N_23831,N_19643,N_17872);
nor U23832 (N_23832,N_18535,N_15694);
nor U23833 (N_23833,N_17167,N_16213);
and U23834 (N_23834,N_16440,N_16858);
nand U23835 (N_23835,N_16432,N_16659);
nand U23836 (N_23836,N_17282,N_18992);
xnor U23837 (N_23837,N_18273,N_17606);
nor U23838 (N_23838,N_17814,N_16041);
nor U23839 (N_23839,N_15858,N_19596);
xor U23840 (N_23840,N_15052,N_15988);
nor U23841 (N_23841,N_16697,N_17607);
xnor U23842 (N_23842,N_16160,N_15928);
and U23843 (N_23843,N_15085,N_19428);
or U23844 (N_23844,N_16745,N_18768);
nand U23845 (N_23845,N_18752,N_19079);
and U23846 (N_23846,N_16345,N_15919);
or U23847 (N_23847,N_15853,N_18060);
nor U23848 (N_23848,N_15376,N_15108);
nand U23849 (N_23849,N_18527,N_18581);
xor U23850 (N_23850,N_17231,N_16797);
xor U23851 (N_23851,N_18688,N_16461);
nor U23852 (N_23852,N_15255,N_16416);
or U23853 (N_23853,N_16807,N_15110);
nand U23854 (N_23854,N_16189,N_17111);
nand U23855 (N_23855,N_17210,N_15183);
or U23856 (N_23856,N_16276,N_18163);
nor U23857 (N_23857,N_16681,N_19966);
or U23858 (N_23858,N_19081,N_17324);
nand U23859 (N_23859,N_15993,N_15429);
and U23860 (N_23860,N_15844,N_18728);
and U23861 (N_23861,N_15673,N_15303);
or U23862 (N_23862,N_15625,N_16605);
nor U23863 (N_23863,N_16503,N_19793);
or U23864 (N_23864,N_17757,N_18991);
xor U23865 (N_23865,N_16732,N_15672);
xor U23866 (N_23866,N_18017,N_19128);
nor U23867 (N_23867,N_15894,N_16411);
and U23868 (N_23868,N_18051,N_19499);
or U23869 (N_23869,N_16261,N_15245);
nor U23870 (N_23870,N_19978,N_18872);
nand U23871 (N_23871,N_16409,N_19015);
or U23872 (N_23872,N_15360,N_15642);
nor U23873 (N_23873,N_18848,N_19110);
or U23874 (N_23874,N_19233,N_15582);
nor U23875 (N_23875,N_17713,N_19495);
nand U23876 (N_23876,N_19158,N_19582);
or U23877 (N_23877,N_15363,N_17893);
xor U23878 (N_23878,N_15896,N_16031);
nor U23879 (N_23879,N_16036,N_16208);
and U23880 (N_23880,N_18228,N_18831);
xor U23881 (N_23881,N_19386,N_15045);
xnor U23882 (N_23882,N_15375,N_15699);
xnor U23883 (N_23883,N_15206,N_16370);
and U23884 (N_23884,N_17223,N_17533);
or U23885 (N_23885,N_16070,N_19354);
nor U23886 (N_23886,N_17606,N_18960);
nor U23887 (N_23887,N_17277,N_16143);
or U23888 (N_23888,N_15826,N_19953);
nand U23889 (N_23889,N_15386,N_15160);
xnor U23890 (N_23890,N_16784,N_16048);
or U23891 (N_23891,N_17306,N_19122);
nor U23892 (N_23892,N_17424,N_18264);
nand U23893 (N_23893,N_19455,N_16871);
or U23894 (N_23894,N_18072,N_17377);
nand U23895 (N_23895,N_17608,N_19755);
nand U23896 (N_23896,N_15070,N_16381);
and U23897 (N_23897,N_19757,N_15609);
nor U23898 (N_23898,N_17707,N_17922);
or U23899 (N_23899,N_16402,N_15489);
and U23900 (N_23900,N_18505,N_15471);
xor U23901 (N_23901,N_18506,N_17342);
xnor U23902 (N_23902,N_19002,N_19397);
xnor U23903 (N_23903,N_18652,N_19719);
xnor U23904 (N_23904,N_19711,N_15082);
xnor U23905 (N_23905,N_17329,N_19303);
and U23906 (N_23906,N_17206,N_17411);
nand U23907 (N_23907,N_17547,N_18075);
and U23908 (N_23908,N_18449,N_17181);
xnor U23909 (N_23909,N_15670,N_15700);
xnor U23910 (N_23910,N_18576,N_19444);
or U23911 (N_23911,N_15018,N_17416);
and U23912 (N_23912,N_16935,N_15635);
nor U23913 (N_23913,N_19582,N_18031);
or U23914 (N_23914,N_15540,N_19916);
or U23915 (N_23915,N_15143,N_17755);
xnor U23916 (N_23916,N_16378,N_15402);
nand U23917 (N_23917,N_19849,N_19588);
xor U23918 (N_23918,N_18976,N_18276);
nor U23919 (N_23919,N_17279,N_16380);
nand U23920 (N_23920,N_19221,N_18533);
xnor U23921 (N_23921,N_17816,N_17861);
nand U23922 (N_23922,N_18703,N_18355);
nor U23923 (N_23923,N_15819,N_18666);
xor U23924 (N_23924,N_15163,N_16478);
and U23925 (N_23925,N_17760,N_16473);
or U23926 (N_23926,N_19625,N_18984);
and U23927 (N_23927,N_17973,N_19230);
xor U23928 (N_23928,N_15691,N_17827);
and U23929 (N_23929,N_17578,N_16662);
and U23930 (N_23930,N_18529,N_17980);
xor U23931 (N_23931,N_16232,N_17234);
nor U23932 (N_23932,N_17944,N_19460);
xnor U23933 (N_23933,N_18040,N_18998);
or U23934 (N_23934,N_16237,N_18195);
nand U23935 (N_23935,N_17224,N_18551);
or U23936 (N_23936,N_18601,N_18342);
and U23937 (N_23937,N_17507,N_15308);
or U23938 (N_23938,N_19640,N_18146);
or U23939 (N_23939,N_17706,N_19186);
xor U23940 (N_23940,N_16282,N_18527);
xor U23941 (N_23941,N_17267,N_16803);
and U23942 (N_23942,N_16934,N_15403);
or U23943 (N_23943,N_16627,N_19929);
xnor U23944 (N_23944,N_19278,N_19066);
nor U23945 (N_23945,N_17564,N_18522);
nor U23946 (N_23946,N_17784,N_16476);
nor U23947 (N_23947,N_18789,N_16792);
nor U23948 (N_23948,N_17402,N_18148);
nand U23949 (N_23949,N_15912,N_19511);
xor U23950 (N_23950,N_17666,N_17199);
and U23951 (N_23951,N_18711,N_15886);
or U23952 (N_23952,N_18417,N_16953);
or U23953 (N_23953,N_16826,N_18485);
and U23954 (N_23954,N_19146,N_15464);
and U23955 (N_23955,N_19556,N_17484);
xor U23956 (N_23956,N_18805,N_18034);
nand U23957 (N_23957,N_16477,N_16529);
and U23958 (N_23958,N_18126,N_19613);
or U23959 (N_23959,N_19776,N_18183);
or U23960 (N_23960,N_18002,N_16200);
nand U23961 (N_23961,N_18644,N_19718);
or U23962 (N_23962,N_17212,N_18445);
xnor U23963 (N_23963,N_17561,N_18089);
nand U23964 (N_23964,N_18192,N_15811);
nand U23965 (N_23965,N_16866,N_16836);
xnor U23966 (N_23966,N_15528,N_19497);
and U23967 (N_23967,N_17681,N_15187);
xor U23968 (N_23968,N_16339,N_19802);
nand U23969 (N_23969,N_16432,N_17253);
and U23970 (N_23970,N_18302,N_18134);
nand U23971 (N_23971,N_16878,N_18267);
or U23972 (N_23972,N_18613,N_19426);
nor U23973 (N_23973,N_15339,N_18146);
and U23974 (N_23974,N_17186,N_16671);
or U23975 (N_23975,N_16527,N_19961);
or U23976 (N_23976,N_18736,N_18046);
and U23977 (N_23977,N_17217,N_19089);
and U23978 (N_23978,N_18151,N_15043);
nand U23979 (N_23979,N_15907,N_19451);
xor U23980 (N_23980,N_17807,N_15469);
nand U23981 (N_23981,N_16838,N_19407);
nand U23982 (N_23982,N_18554,N_17419);
nor U23983 (N_23983,N_19512,N_15383);
or U23984 (N_23984,N_16610,N_19408);
nand U23985 (N_23985,N_17000,N_16617);
nor U23986 (N_23986,N_15982,N_18357);
nand U23987 (N_23987,N_15882,N_19870);
nor U23988 (N_23988,N_16099,N_17378);
nand U23989 (N_23989,N_17735,N_18011);
or U23990 (N_23990,N_16307,N_16897);
or U23991 (N_23991,N_18572,N_16416);
nor U23992 (N_23992,N_15189,N_16380);
xnor U23993 (N_23993,N_15199,N_15451);
nor U23994 (N_23994,N_17662,N_17951);
xnor U23995 (N_23995,N_16278,N_19042);
xnor U23996 (N_23996,N_19051,N_17689);
and U23997 (N_23997,N_15018,N_18098);
or U23998 (N_23998,N_18329,N_17556);
xor U23999 (N_23999,N_15576,N_16974);
xnor U24000 (N_24000,N_17405,N_16016);
xor U24001 (N_24001,N_16734,N_19553);
nand U24002 (N_24002,N_17771,N_16599);
or U24003 (N_24003,N_17688,N_17824);
or U24004 (N_24004,N_15545,N_17396);
nor U24005 (N_24005,N_17041,N_18526);
nand U24006 (N_24006,N_17577,N_17266);
and U24007 (N_24007,N_15060,N_18434);
nand U24008 (N_24008,N_18161,N_16790);
xor U24009 (N_24009,N_18396,N_17462);
nand U24010 (N_24010,N_15092,N_15788);
xnor U24011 (N_24011,N_15994,N_16142);
or U24012 (N_24012,N_17614,N_15988);
nor U24013 (N_24013,N_17800,N_17431);
or U24014 (N_24014,N_15902,N_17983);
or U24015 (N_24015,N_16173,N_17941);
nand U24016 (N_24016,N_18072,N_18204);
nand U24017 (N_24017,N_17227,N_17186);
and U24018 (N_24018,N_18651,N_16983);
nor U24019 (N_24019,N_18220,N_17849);
nor U24020 (N_24020,N_16211,N_15409);
nor U24021 (N_24021,N_18957,N_16822);
or U24022 (N_24022,N_15912,N_15974);
xnor U24023 (N_24023,N_17090,N_18400);
nand U24024 (N_24024,N_19781,N_19520);
xor U24025 (N_24025,N_15543,N_15152);
nand U24026 (N_24026,N_16740,N_15443);
and U24027 (N_24027,N_18860,N_18993);
or U24028 (N_24028,N_19371,N_17901);
and U24029 (N_24029,N_19888,N_15576);
xnor U24030 (N_24030,N_16652,N_18692);
and U24031 (N_24031,N_16430,N_18422);
xnor U24032 (N_24032,N_18453,N_19635);
and U24033 (N_24033,N_18700,N_18593);
nand U24034 (N_24034,N_18060,N_15317);
or U24035 (N_24035,N_16581,N_19365);
or U24036 (N_24036,N_17090,N_16378);
and U24037 (N_24037,N_19473,N_19658);
nor U24038 (N_24038,N_17742,N_17035);
nor U24039 (N_24039,N_18714,N_17202);
or U24040 (N_24040,N_15253,N_18221);
xnor U24041 (N_24041,N_19967,N_15776);
and U24042 (N_24042,N_19853,N_16783);
or U24043 (N_24043,N_16842,N_15504);
nor U24044 (N_24044,N_15472,N_15153);
nand U24045 (N_24045,N_18594,N_19957);
xor U24046 (N_24046,N_15353,N_17480);
nand U24047 (N_24047,N_19566,N_16828);
and U24048 (N_24048,N_15264,N_18671);
xor U24049 (N_24049,N_15179,N_16541);
nand U24050 (N_24050,N_17642,N_17587);
xnor U24051 (N_24051,N_15025,N_16159);
and U24052 (N_24052,N_19226,N_19995);
or U24053 (N_24053,N_16478,N_17070);
and U24054 (N_24054,N_16680,N_19833);
nor U24055 (N_24055,N_15833,N_17950);
nand U24056 (N_24056,N_15510,N_16371);
or U24057 (N_24057,N_17318,N_16015);
and U24058 (N_24058,N_16062,N_17634);
nand U24059 (N_24059,N_16385,N_15847);
nor U24060 (N_24060,N_18276,N_19938);
nor U24061 (N_24061,N_18092,N_16066);
nor U24062 (N_24062,N_17002,N_17611);
and U24063 (N_24063,N_15675,N_15814);
and U24064 (N_24064,N_18738,N_17406);
and U24065 (N_24065,N_16446,N_16042);
nor U24066 (N_24066,N_16579,N_18979);
xor U24067 (N_24067,N_17464,N_17278);
or U24068 (N_24068,N_16226,N_18258);
nand U24069 (N_24069,N_17548,N_16240);
and U24070 (N_24070,N_19337,N_18967);
nand U24071 (N_24071,N_15794,N_16507);
nand U24072 (N_24072,N_16941,N_16821);
and U24073 (N_24073,N_18069,N_19715);
xnor U24074 (N_24074,N_15057,N_19918);
or U24075 (N_24075,N_18949,N_18945);
nand U24076 (N_24076,N_15233,N_15923);
nand U24077 (N_24077,N_19671,N_17574);
nor U24078 (N_24078,N_15741,N_17352);
or U24079 (N_24079,N_17764,N_19664);
nand U24080 (N_24080,N_15702,N_16769);
nand U24081 (N_24081,N_18176,N_17314);
or U24082 (N_24082,N_18770,N_16027);
xor U24083 (N_24083,N_15019,N_15361);
or U24084 (N_24084,N_18124,N_19256);
and U24085 (N_24085,N_19403,N_19625);
nand U24086 (N_24086,N_19125,N_17753);
or U24087 (N_24087,N_16888,N_19522);
or U24088 (N_24088,N_17897,N_15053);
xor U24089 (N_24089,N_15617,N_17221);
nand U24090 (N_24090,N_15986,N_18572);
nand U24091 (N_24091,N_15252,N_17104);
xnor U24092 (N_24092,N_16786,N_18487);
nor U24093 (N_24093,N_18910,N_18392);
xnor U24094 (N_24094,N_17618,N_19117);
xor U24095 (N_24095,N_19710,N_16250);
and U24096 (N_24096,N_19568,N_18978);
nand U24097 (N_24097,N_16984,N_18735);
nand U24098 (N_24098,N_16780,N_18714);
or U24099 (N_24099,N_16595,N_15673);
nor U24100 (N_24100,N_19369,N_16624);
nand U24101 (N_24101,N_17182,N_17694);
or U24102 (N_24102,N_15939,N_16411);
and U24103 (N_24103,N_19679,N_15936);
nor U24104 (N_24104,N_15737,N_18677);
nand U24105 (N_24105,N_19910,N_16225);
or U24106 (N_24106,N_16276,N_18589);
and U24107 (N_24107,N_19442,N_17959);
or U24108 (N_24108,N_17362,N_15328);
or U24109 (N_24109,N_18911,N_19590);
nand U24110 (N_24110,N_19939,N_15038);
nor U24111 (N_24111,N_16042,N_19635);
and U24112 (N_24112,N_18084,N_17928);
or U24113 (N_24113,N_17359,N_16882);
or U24114 (N_24114,N_19980,N_18259);
nand U24115 (N_24115,N_15018,N_19713);
or U24116 (N_24116,N_19764,N_16802);
and U24117 (N_24117,N_19577,N_16379);
nand U24118 (N_24118,N_15557,N_15008);
or U24119 (N_24119,N_15443,N_15680);
or U24120 (N_24120,N_19193,N_17304);
or U24121 (N_24121,N_18964,N_15775);
and U24122 (N_24122,N_17417,N_18420);
nand U24123 (N_24123,N_19082,N_15455);
nor U24124 (N_24124,N_15389,N_18875);
or U24125 (N_24125,N_18774,N_16181);
nor U24126 (N_24126,N_15122,N_17147);
xnor U24127 (N_24127,N_15906,N_19638);
xnor U24128 (N_24128,N_16839,N_16711);
xor U24129 (N_24129,N_16170,N_15145);
or U24130 (N_24130,N_19246,N_15084);
nor U24131 (N_24131,N_19635,N_18871);
xor U24132 (N_24132,N_16393,N_17841);
and U24133 (N_24133,N_18221,N_15473);
or U24134 (N_24134,N_19717,N_15078);
nand U24135 (N_24135,N_15290,N_17914);
xnor U24136 (N_24136,N_17237,N_15849);
and U24137 (N_24137,N_16542,N_16235);
nor U24138 (N_24138,N_17276,N_15358);
and U24139 (N_24139,N_16361,N_15106);
or U24140 (N_24140,N_19007,N_17507);
or U24141 (N_24141,N_15726,N_18664);
nor U24142 (N_24142,N_17661,N_19662);
nand U24143 (N_24143,N_19581,N_19061);
and U24144 (N_24144,N_19650,N_18826);
nand U24145 (N_24145,N_16321,N_18563);
xor U24146 (N_24146,N_18710,N_16758);
xor U24147 (N_24147,N_17929,N_18672);
xnor U24148 (N_24148,N_16861,N_16441);
and U24149 (N_24149,N_18177,N_17465);
and U24150 (N_24150,N_18278,N_17997);
nor U24151 (N_24151,N_15170,N_15866);
and U24152 (N_24152,N_19809,N_19696);
xnor U24153 (N_24153,N_17914,N_18592);
xnor U24154 (N_24154,N_17841,N_18361);
xnor U24155 (N_24155,N_19708,N_18638);
nor U24156 (N_24156,N_15037,N_18720);
nor U24157 (N_24157,N_16496,N_16273);
or U24158 (N_24158,N_18127,N_19249);
xor U24159 (N_24159,N_15396,N_19926);
and U24160 (N_24160,N_16043,N_15125);
xor U24161 (N_24161,N_16368,N_17564);
and U24162 (N_24162,N_17871,N_18319);
xnor U24163 (N_24163,N_15641,N_18603);
xnor U24164 (N_24164,N_18888,N_17897);
nand U24165 (N_24165,N_15481,N_18729);
xnor U24166 (N_24166,N_16034,N_18286);
or U24167 (N_24167,N_17219,N_19931);
and U24168 (N_24168,N_16747,N_19391);
and U24169 (N_24169,N_16330,N_15505);
nand U24170 (N_24170,N_15371,N_16490);
and U24171 (N_24171,N_17882,N_18993);
nor U24172 (N_24172,N_19277,N_15945);
or U24173 (N_24173,N_16649,N_16243);
nand U24174 (N_24174,N_16435,N_17517);
or U24175 (N_24175,N_15085,N_17466);
nand U24176 (N_24176,N_18855,N_18092);
nand U24177 (N_24177,N_17224,N_18412);
xor U24178 (N_24178,N_18556,N_17098);
xor U24179 (N_24179,N_15165,N_18201);
nand U24180 (N_24180,N_15809,N_19591);
and U24181 (N_24181,N_16344,N_16354);
nor U24182 (N_24182,N_18725,N_19049);
xor U24183 (N_24183,N_15917,N_19440);
or U24184 (N_24184,N_16884,N_16321);
nor U24185 (N_24185,N_16892,N_17107);
xor U24186 (N_24186,N_18268,N_17236);
and U24187 (N_24187,N_19237,N_18485);
xor U24188 (N_24188,N_16585,N_17447);
and U24189 (N_24189,N_19228,N_19029);
nand U24190 (N_24190,N_15745,N_16379);
nor U24191 (N_24191,N_19418,N_16133);
and U24192 (N_24192,N_15343,N_19890);
or U24193 (N_24193,N_18392,N_19534);
xnor U24194 (N_24194,N_18813,N_16682);
nor U24195 (N_24195,N_18730,N_18586);
and U24196 (N_24196,N_17578,N_15308);
nor U24197 (N_24197,N_19869,N_18274);
and U24198 (N_24198,N_16955,N_17533);
xnor U24199 (N_24199,N_16825,N_17729);
nand U24200 (N_24200,N_17179,N_16038);
or U24201 (N_24201,N_17087,N_17463);
and U24202 (N_24202,N_16179,N_16556);
nor U24203 (N_24203,N_16304,N_18945);
and U24204 (N_24204,N_19620,N_18767);
xnor U24205 (N_24205,N_15576,N_19468);
nand U24206 (N_24206,N_19983,N_19841);
and U24207 (N_24207,N_18592,N_19413);
xnor U24208 (N_24208,N_19296,N_17133);
xor U24209 (N_24209,N_16223,N_18614);
nand U24210 (N_24210,N_16440,N_17307);
nand U24211 (N_24211,N_18565,N_18445);
nor U24212 (N_24212,N_16841,N_19292);
xnor U24213 (N_24213,N_16351,N_16543);
xor U24214 (N_24214,N_16738,N_18525);
nand U24215 (N_24215,N_18278,N_16743);
nand U24216 (N_24216,N_16475,N_15918);
and U24217 (N_24217,N_15263,N_17246);
nor U24218 (N_24218,N_19551,N_18639);
nand U24219 (N_24219,N_16630,N_17396);
nand U24220 (N_24220,N_19686,N_15832);
and U24221 (N_24221,N_18484,N_16524);
nand U24222 (N_24222,N_18253,N_19567);
xor U24223 (N_24223,N_16293,N_17332);
or U24224 (N_24224,N_19292,N_18059);
nor U24225 (N_24225,N_19138,N_16145);
nor U24226 (N_24226,N_17393,N_15296);
or U24227 (N_24227,N_16733,N_16851);
xor U24228 (N_24228,N_18067,N_18919);
nor U24229 (N_24229,N_17516,N_19695);
xor U24230 (N_24230,N_19798,N_19701);
xor U24231 (N_24231,N_15016,N_16292);
xnor U24232 (N_24232,N_19882,N_18889);
xnor U24233 (N_24233,N_17465,N_16997);
nand U24234 (N_24234,N_15377,N_16782);
xor U24235 (N_24235,N_17617,N_19456);
xnor U24236 (N_24236,N_18299,N_19027);
or U24237 (N_24237,N_16240,N_15236);
or U24238 (N_24238,N_19795,N_16956);
xnor U24239 (N_24239,N_19356,N_16614);
or U24240 (N_24240,N_15477,N_19228);
and U24241 (N_24241,N_18266,N_17493);
or U24242 (N_24242,N_15477,N_16693);
or U24243 (N_24243,N_18042,N_15951);
and U24244 (N_24244,N_16951,N_15897);
and U24245 (N_24245,N_18777,N_16043);
nor U24246 (N_24246,N_17236,N_19687);
nand U24247 (N_24247,N_16208,N_17295);
and U24248 (N_24248,N_15402,N_19108);
nor U24249 (N_24249,N_17365,N_18642);
nand U24250 (N_24250,N_16032,N_17284);
and U24251 (N_24251,N_19849,N_15064);
or U24252 (N_24252,N_15446,N_16985);
nor U24253 (N_24253,N_16661,N_16169);
xnor U24254 (N_24254,N_17007,N_17213);
nor U24255 (N_24255,N_19995,N_17433);
nor U24256 (N_24256,N_16427,N_15716);
xnor U24257 (N_24257,N_16110,N_16642);
nor U24258 (N_24258,N_18477,N_18895);
and U24259 (N_24259,N_19928,N_19258);
nand U24260 (N_24260,N_19054,N_19352);
xor U24261 (N_24261,N_16956,N_17403);
or U24262 (N_24262,N_17683,N_18282);
xor U24263 (N_24263,N_19688,N_17832);
nand U24264 (N_24264,N_15238,N_19748);
and U24265 (N_24265,N_18872,N_19410);
xor U24266 (N_24266,N_19291,N_15289);
or U24267 (N_24267,N_17537,N_17957);
nor U24268 (N_24268,N_15771,N_16271);
nand U24269 (N_24269,N_16620,N_17923);
or U24270 (N_24270,N_15488,N_19489);
or U24271 (N_24271,N_19852,N_17565);
or U24272 (N_24272,N_16169,N_18435);
nand U24273 (N_24273,N_19304,N_17932);
nand U24274 (N_24274,N_15967,N_16607);
or U24275 (N_24275,N_17021,N_15887);
and U24276 (N_24276,N_18649,N_15589);
and U24277 (N_24277,N_19339,N_17739);
nor U24278 (N_24278,N_18807,N_17364);
or U24279 (N_24279,N_15117,N_19145);
or U24280 (N_24280,N_17860,N_16044);
or U24281 (N_24281,N_18322,N_19388);
xnor U24282 (N_24282,N_18835,N_16089);
nand U24283 (N_24283,N_19226,N_18717);
nand U24284 (N_24284,N_19640,N_17467);
or U24285 (N_24285,N_15674,N_18443);
and U24286 (N_24286,N_17717,N_15195);
nor U24287 (N_24287,N_15467,N_19376);
xor U24288 (N_24288,N_17273,N_16264);
nand U24289 (N_24289,N_15884,N_15710);
nor U24290 (N_24290,N_17102,N_17445);
and U24291 (N_24291,N_18297,N_15001);
or U24292 (N_24292,N_15442,N_19696);
nand U24293 (N_24293,N_18197,N_16759);
or U24294 (N_24294,N_15359,N_19764);
and U24295 (N_24295,N_19601,N_17781);
or U24296 (N_24296,N_15209,N_17739);
and U24297 (N_24297,N_16995,N_18445);
nand U24298 (N_24298,N_16395,N_15316);
or U24299 (N_24299,N_15612,N_17762);
nor U24300 (N_24300,N_15570,N_19134);
and U24301 (N_24301,N_16230,N_17464);
xor U24302 (N_24302,N_19703,N_18383);
xor U24303 (N_24303,N_18029,N_17867);
xor U24304 (N_24304,N_18789,N_15257);
nand U24305 (N_24305,N_18546,N_15407);
nand U24306 (N_24306,N_18681,N_18130);
or U24307 (N_24307,N_15542,N_17217);
xor U24308 (N_24308,N_16750,N_17386);
or U24309 (N_24309,N_17842,N_19034);
xnor U24310 (N_24310,N_18676,N_15576);
nand U24311 (N_24311,N_16959,N_16863);
and U24312 (N_24312,N_17995,N_19461);
and U24313 (N_24313,N_17851,N_18688);
or U24314 (N_24314,N_18698,N_18059);
nor U24315 (N_24315,N_18523,N_17206);
xor U24316 (N_24316,N_16425,N_18857);
xnor U24317 (N_24317,N_16442,N_17120);
and U24318 (N_24318,N_18108,N_18079);
and U24319 (N_24319,N_17350,N_19294);
or U24320 (N_24320,N_19057,N_18148);
or U24321 (N_24321,N_17089,N_17805);
and U24322 (N_24322,N_18642,N_16208);
nand U24323 (N_24323,N_18581,N_16458);
xnor U24324 (N_24324,N_19925,N_19139);
xnor U24325 (N_24325,N_19272,N_15068);
and U24326 (N_24326,N_19327,N_15288);
nand U24327 (N_24327,N_19579,N_17998);
nor U24328 (N_24328,N_17405,N_18311);
or U24329 (N_24329,N_19697,N_19361);
nor U24330 (N_24330,N_18958,N_16529);
and U24331 (N_24331,N_15000,N_16346);
nand U24332 (N_24332,N_16077,N_17997);
nor U24333 (N_24333,N_19813,N_16396);
nor U24334 (N_24334,N_19668,N_19498);
nand U24335 (N_24335,N_18094,N_15019);
and U24336 (N_24336,N_18276,N_17870);
nor U24337 (N_24337,N_15955,N_16612);
nor U24338 (N_24338,N_18677,N_18403);
nand U24339 (N_24339,N_15608,N_17991);
nor U24340 (N_24340,N_16212,N_17363);
nand U24341 (N_24341,N_19445,N_15479);
xor U24342 (N_24342,N_18335,N_17048);
xor U24343 (N_24343,N_17751,N_16871);
nand U24344 (N_24344,N_19722,N_19556);
xnor U24345 (N_24345,N_15312,N_19018);
nor U24346 (N_24346,N_16803,N_19254);
and U24347 (N_24347,N_19301,N_18802);
xnor U24348 (N_24348,N_16936,N_15861);
and U24349 (N_24349,N_18597,N_17623);
or U24350 (N_24350,N_16121,N_18771);
nor U24351 (N_24351,N_15750,N_19799);
and U24352 (N_24352,N_18839,N_16305);
xor U24353 (N_24353,N_19795,N_16287);
xor U24354 (N_24354,N_18399,N_19393);
xor U24355 (N_24355,N_17592,N_18554);
nor U24356 (N_24356,N_17951,N_15653);
and U24357 (N_24357,N_18874,N_15324);
nor U24358 (N_24358,N_16653,N_19463);
or U24359 (N_24359,N_18345,N_17301);
xor U24360 (N_24360,N_18472,N_16156);
or U24361 (N_24361,N_19061,N_16105);
nand U24362 (N_24362,N_19650,N_16350);
xnor U24363 (N_24363,N_19738,N_15120);
nand U24364 (N_24364,N_16003,N_15817);
nor U24365 (N_24365,N_18057,N_17419);
xnor U24366 (N_24366,N_16577,N_16361);
nor U24367 (N_24367,N_15735,N_19936);
xnor U24368 (N_24368,N_17487,N_19357);
nand U24369 (N_24369,N_19957,N_18032);
or U24370 (N_24370,N_17466,N_15327);
or U24371 (N_24371,N_19529,N_17539);
nor U24372 (N_24372,N_17029,N_17742);
nand U24373 (N_24373,N_15428,N_19874);
and U24374 (N_24374,N_16313,N_17451);
xor U24375 (N_24375,N_19979,N_19076);
nor U24376 (N_24376,N_15336,N_17814);
nor U24377 (N_24377,N_16456,N_15660);
xnor U24378 (N_24378,N_16737,N_15256);
or U24379 (N_24379,N_19310,N_19579);
or U24380 (N_24380,N_15007,N_19322);
nor U24381 (N_24381,N_17465,N_15983);
xor U24382 (N_24382,N_16933,N_18649);
and U24383 (N_24383,N_16084,N_15679);
nand U24384 (N_24384,N_18283,N_17752);
xor U24385 (N_24385,N_16166,N_19083);
or U24386 (N_24386,N_16337,N_15915);
nand U24387 (N_24387,N_17062,N_18743);
nand U24388 (N_24388,N_19302,N_16140);
or U24389 (N_24389,N_17964,N_18850);
or U24390 (N_24390,N_18111,N_17410);
nand U24391 (N_24391,N_19767,N_18608);
nand U24392 (N_24392,N_18080,N_18065);
xor U24393 (N_24393,N_19656,N_17648);
or U24394 (N_24394,N_16904,N_19822);
nor U24395 (N_24395,N_19418,N_15791);
and U24396 (N_24396,N_16123,N_17260);
nor U24397 (N_24397,N_15611,N_17441);
xor U24398 (N_24398,N_15128,N_17630);
xor U24399 (N_24399,N_15741,N_18849);
or U24400 (N_24400,N_18209,N_17344);
and U24401 (N_24401,N_18111,N_18552);
xor U24402 (N_24402,N_19134,N_18189);
or U24403 (N_24403,N_18853,N_15695);
nor U24404 (N_24404,N_16076,N_15962);
xor U24405 (N_24405,N_19789,N_19987);
and U24406 (N_24406,N_19864,N_18570);
xor U24407 (N_24407,N_17051,N_16519);
nand U24408 (N_24408,N_18299,N_18154);
nor U24409 (N_24409,N_18523,N_15456);
xor U24410 (N_24410,N_19746,N_18722);
and U24411 (N_24411,N_19763,N_18504);
nor U24412 (N_24412,N_16322,N_18886);
nor U24413 (N_24413,N_18944,N_18726);
nor U24414 (N_24414,N_16586,N_16000);
nand U24415 (N_24415,N_15763,N_16646);
xnor U24416 (N_24416,N_15050,N_17855);
xor U24417 (N_24417,N_18967,N_18113);
or U24418 (N_24418,N_19041,N_16854);
nor U24419 (N_24419,N_15755,N_17683);
nor U24420 (N_24420,N_18091,N_18448);
or U24421 (N_24421,N_15969,N_19431);
or U24422 (N_24422,N_17060,N_18821);
xnor U24423 (N_24423,N_16415,N_16923);
or U24424 (N_24424,N_19640,N_15356);
or U24425 (N_24425,N_16883,N_15214);
nor U24426 (N_24426,N_19995,N_16505);
nand U24427 (N_24427,N_18137,N_15905);
nand U24428 (N_24428,N_17340,N_19710);
nor U24429 (N_24429,N_19139,N_19395);
nor U24430 (N_24430,N_15970,N_16057);
or U24431 (N_24431,N_19721,N_18774);
or U24432 (N_24432,N_19837,N_15773);
nand U24433 (N_24433,N_18495,N_18810);
or U24434 (N_24434,N_17465,N_15584);
and U24435 (N_24435,N_18251,N_17188);
nor U24436 (N_24436,N_19473,N_19370);
nor U24437 (N_24437,N_16321,N_15747);
or U24438 (N_24438,N_19497,N_18194);
and U24439 (N_24439,N_18671,N_16404);
or U24440 (N_24440,N_16216,N_17458);
nor U24441 (N_24441,N_16240,N_18825);
nand U24442 (N_24442,N_16579,N_17696);
and U24443 (N_24443,N_15981,N_15630);
nor U24444 (N_24444,N_18117,N_17732);
or U24445 (N_24445,N_16763,N_19478);
or U24446 (N_24446,N_18159,N_15640);
and U24447 (N_24447,N_18846,N_15368);
or U24448 (N_24448,N_16735,N_18779);
and U24449 (N_24449,N_19894,N_19121);
xnor U24450 (N_24450,N_16568,N_17900);
or U24451 (N_24451,N_15161,N_15849);
nor U24452 (N_24452,N_15984,N_19544);
nor U24453 (N_24453,N_19977,N_17049);
xnor U24454 (N_24454,N_19194,N_18438);
and U24455 (N_24455,N_16951,N_19932);
and U24456 (N_24456,N_18963,N_15994);
and U24457 (N_24457,N_15590,N_16294);
or U24458 (N_24458,N_18302,N_17942);
xnor U24459 (N_24459,N_17188,N_18553);
or U24460 (N_24460,N_16404,N_18199);
nor U24461 (N_24461,N_15945,N_19690);
xnor U24462 (N_24462,N_15016,N_18492);
and U24463 (N_24463,N_18681,N_17461);
nand U24464 (N_24464,N_15137,N_16475);
nor U24465 (N_24465,N_18533,N_15327);
and U24466 (N_24466,N_19483,N_19968);
or U24467 (N_24467,N_15626,N_15803);
or U24468 (N_24468,N_18019,N_15063);
or U24469 (N_24469,N_15626,N_17557);
nand U24470 (N_24470,N_15844,N_17878);
nand U24471 (N_24471,N_17572,N_16854);
xor U24472 (N_24472,N_17748,N_18842);
nor U24473 (N_24473,N_17812,N_19975);
nand U24474 (N_24474,N_16128,N_16469);
xnor U24475 (N_24475,N_18569,N_19003);
nor U24476 (N_24476,N_16684,N_15676);
or U24477 (N_24477,N_19881,N_16827);
and U24478 (N_24478,N_19271,N_16718);
nand U24479 (N_24479,N_15301,N_18017);
nor U24480 (N_24480,N_18136,N_17828);
nand U24481 (N_24481,N_19940,N_16817);
nor U24482 (N_24482,N_19251,N_15075);
and U24483 (N_24483,N_19620,N_17385);
nand U24484 (N_24484,N_16909,N_15969);
or U24485 (N_24485,N_19312,N_16986);
nand U24486 (N_24486,N_19593,N_19505);
nor U24487 (N_24487,N_15369,N_15980);
nor U24488 (N_24488,N_19678,N_16286);
xnor U24489 (N_24489,N_19416,N_15299);
or U24490 (N_24490,N_15178,N_19854);
and U24491 (N_24491,N_16561,N_17749);
nor U24492 (N_24492,N_16850,N_15270);
or U24493 (N_24493,N_19520,N_19561);
xnor U24494 (N_24494,N_18714,N_18569);
and U24495 (N_24495,N_19797,N_19477);
nand U24496 (N_24496,N_15723,N_19956);
nor U24497 (N_24497,N_18989,N_18941);
xor U24498 (N_24498,N_18463,N_18671);
and U24499 (N_24499,N_17203,N_19417);
xor U24500 (N_24500,N_18414,N_19017);
nand U24501 (N_24501,N_19132,N_17352);
nor U24502 (N_24502,N_16097,N_17957);
xnor U24503 (N_24503,N_18128,N_15046);
nor U24504 (N_24504,N_17205,N_19111);
or U24505 (N_24505,N_16258,N_16844);
or U24506 (N_24506,N_18260,N_15442);
or U24507 (N_24507,N_18285,N_18776);
nor U24508 (N_24508,N_16849,N_17804);
and U24509 (N_24509,N_16981,N_19028);
xnor U24510 (N_24510,N_18703,N_16183);
xor U24511 (N_24511,N_19728,N_19896);
nor U24512 (N_24512,N_18284,N_16544);
xnor U24513 (N_24513,N_19936,N_17859);
xor U24514 (N_24514,N_16938,N_16659);
nor U24515 (N_24515,N_18764,N_15864);
or U24516 (N_24516,N_15075,N_16363);
or U24517 (N_24517,N_17386,N_15517);
xor U24518 (N_24518,N_18527,N_19342);
and U24519 (N_24519,N_16087,N_17870);
or U24520 (N_24520,N_16339,N_17167);
or U24521 (N_24521,N_18378,N_18312);
nor U24522 (N_24522,N_19563,N_18510);
or U24523 (N_24523,N_18461,N_19545);
nor U24524 (N_24524,N_16883,N_17738);
nand U24525 (N_24525,N_18099,N_16238);
nand U24526 (N_24526,N_17807,N_17380);
nor U24527 (N_24527,N_17232,N_17575);
nor U24528 (N_24528,N_17320,N_17267);
nor U24529 (N_24529,N_19108,N_18860);
nor U24530 (N_24530,N_18933,N_17400);
and U24531 (N_24531,N_17930,N_18492);
and U24532 (N_24532,N_17397,N_16074);
nor U24533 (N_24533,N_16196,N_17987);
or U24534 (N_24534,N_19076,N_15507);
nor U24535 (N_24535,N_17679,N_19600);
xnor U24536 (N_24536,N_16165,N_15047);
or U24537 (N_24537,N_16318,N_19132);
nand U24538 (N_24538,N_16486,N_17518);
or U24539 (N_24539,N_19097,N_19355);
nand U24540 (N_24540,N_15447,N_18752);
or U24541 (N_24541,N_18026,N_19872);
and U24542 (N_24542,N_15370,N_18049);
and U24543 (N_24543,N_17459,N_19901);
nand U24544 (N_24544,N_17789,N_15429);
nand U24545 (N_24545,N_18736,N_16100);
nor U24546 (N_24546,N_15746,N_18463);
nor U24547 (N_24547,N_15820,N_16874);
nand U24548 (N_24548,N_15260,N_18718);
nand U24549 (N_24549,N_19012,N_18847);
nand U24550 (N_24550,N_17527,N_17195);
xnor U24551 (N_24551,N_19877,N_18257);
nand U24552 (N_24552,N_16725,N_19452);
nor U24553 (N_24553,N_16225,N_17039);
xor U24554 (N_24554,N_16680,N_17117);
and U24555 (N_24555,N_19012,N_16135);
nand U24556 (N_24556,N_15035,N_16055);
nor U24557 (N_24557,N_19174,N_15879);
xnor U24558 (N_24558,N_19694,N_16417);
and U24559 (N_24559,N_17274,N_17707);
nor U24560 (N_24560,N_16316,N_15897);
xor U24561 (N_24561,N_17202,N_19605);
nor U24562 (N_24562,N_15813,N_15687);
and U24563 (N_24563,N_15996,N_17238);
nor U24564 (N_24564,N_18697,N_15146);
nand U24565 (N_24565,N_17958,N_16608);
and U24566 (N_24566,N_19182,N_19831);
xnor U24567 (N_24567,N_19544,N_17601);
nor U24568 (N_24568,N_18132,N_18601);
and U24569 (N_24569,N_19251,N_19707);
nor U24570 (N_24570,N_17423,N_17853);
and U24571 (N_24571,N_19565,N_17109);
nand U24572 (N_24572,N_15706,N_18323);
and U24573 (N_24573,N_19183,N_16415);
xor U24574 (N_24574,N_19842,N_17469);
nand U24575 (N_24575,N_15372,N_17702);
nor U24576 (N_24576,N_18354,N_16236);
nor U24577 (N_24577,N_18656,N_18722);
nor U24578 (N_24578,N_19404,N_19161);
nor U24579 (N_24579,N_18276,N_17747);
nor U24580 (N_24580,N_17065,N_18689);
nor U24581 (N_24581,N_17114,N_17859);
and U24582 (N_24582,N_17911,N_16782);
nor U24583 (N_24583,N_16594,N_17336);
and U24584 (N_24584,N_16059,N_19166);
or U24585 (N_24585,N_19288,N_16025);
or U24586 (N_24586,N_18517,N_19366);
or U24587 (N_24587,N_15637,N_16237);
xnor U24588 (N_24588,N_16978,N_18877);
or U24589 (N_24589,N_18100,N_16106);
nand U24590 (N_24590,N_17073,N_18795);
nand U24591 (N_24591,N_18145,N_15189);
and U24592 (N_24592,N_19011,N_19931);
nor U24593 (N_24593,N_18473,N_18352);
or U24594 (N_24594,N_18503,N_16812);
xor U24595 (N_24595,N_19388,N_15830);
and U24596 (N_24596,N_17274,N_16031);
nand U24597 (N_24597,N_19603,N_18759);
and U24598 (N_24598,N_17140,N_18524);
and U24599 (N_24599,N_18113,N_17184);
nor U24600 (N_24600,N_18306,N_17580);
and U24601 (N_24601,N_19869,N_15917);
nand U24602 (N_24602,N_19042,N_19814);
xnor U24603 (N_24603,N_19674,N_16667);
and U24604 (N_24604,N_17117,N_18888);
nand U24605 (N_24605,N_18581,N_19495);
nand U24606 (N_24606,N_16925,N_16502);
xor U24607 (N_24607,N_18977,N_15327);
and U24608 (N_24608,N_15007,N_15982);
xnor U24609 (N_24609,N_16286,N_16796);
nand U24610 (N_24610,N_19128,N_16888);
or U24611 (N_24611,N_18131,N_17080);
nand U24612 (N_24612,N_18501,N_16086);
nor U24613 (N_24613,N_18295,N_15156);
and U24614 (N_24614,N_19467,N_19678);
nor U24615 (N_24615,N_15317,N_17184);
nor U24616 (N_24616,N_16920,N_18019);
and U24617 (N_24617,N_16747,N_16463);
nor U24618 (N_24618,N_16305,N_17489);
or U24619 (N_24619,N_15606,N_17735);
and U24620 (N_24620,N_15196,N_16278);
nand U24621 (N_24621,N_18891,N_19956);
nand U24622 (N_24622,N_16938,N_18790);
nor U24623 (N_24623,N_19586,N_18628);
xor U24624 (N_24624,N_16366,N_19937);
or U24625 (N_24625,N_15453,N_15389);
or U24626 (N_24626,N_16722,N_19445);
nand U24627 (N_24627,N_16261,N_17946);
or U24628 (N_24628,N_16007,N_18605);
nand U24629 (N_24629,N_16357,N_19379);
nand U24630 (N_24630,N_16887,N_15333);
nor U24631 (N_24631,N_19202,N_15874);
or U24632 (N_24632,N_18096,N_16627);
and U24633 (N_24633,N_16741,N_17081);
or U24634 (N_24634,N_18549,N_18593);
and U24635 (N_24635,N_18919,N_16326);
nor U24636 (N_24636,N_17003,N_18774);
nor U24637 (N_24637,N_17658,N_18312);
xnor U24638 (N_24638,N_17187,N_16845);
nor U24639 (N_24639,N_19910,N_15939);
xor U24640 (N_24640,N_17018,N_18828);
and U24641 (N_24641,N_19298,N_18792);
and U24642 (N_24642,N_18047,N_17710);
xor U24643 (N_24643,N_17675,N_16677);
and U24644 (N_24644,N_16676,N_18394);
xor U24645 (N_24645,N_17920,N_18680);
and U24646 (N_24646,N_19095,N_17119);
and U24647 (N_24647,N_19709,N_19699);
nand U24648 (N_24648,N_18054,N_15969);
and U24649 (N_24649,N_16116,N_16861);
xnor U24650 (N_24650,N_19847,N_15202);
or U24651 (N_24651,N_16047,N_17766);
or U24652 (N_24652,N_18072,N_19510);
nand U24653 (N_24653,N_16489,N_16298);
xor U24654 (N_24654,N_17993,N_17984);
and U24655 (N_24655,N_16153,N_17534);
or U24656 (N_24656,N_18799,N_16668);
or U24657 (N_24657,N_16803,N_16309);
and U24658 (N_24658,N_19952,N_17370);
nand U24659 (N_24659,N_19227,N_18654);
xnor U24660 (N_24660,N_19400,N_15567);
nor U24661 (N_24661,N_18508,N_18465);
or U24662 (N_24662,N_16813,N_18593);
nor U24663 (N_24663,N_15289,N_16897);
or U24664 (N_24664,N_18945,N_17870);
xor U24665 (N_24665,N_18225,N_17853);
or U24666 (N_24666,N_15401,N_17211);
nand U24667 (N_24667,N_17984,N_16959);
nor U24668 (N_24668,N_15332,N_18138);
nor U24669 (N_24669,N_16681,N_16298);
nor U24670 (N_24670,N_16783,N_19567);
nor U24671 (N_24671,N_15315,N_15414);
and U24672 (N_24672,N_15431,N_19370);
and U24673 (N_24673,N_17161,N_17353);
nand U24674 (N_24674,N_17784,N_16822);
and U24675 (N_24675,N_18837,N_18715);
nor U24676 (N_24676,N_18501,N_19979);
xnor U24677 (N_24677,N_18041,N_15171);
nor U24678 (N_24678,N_16238,N_19915);
or U24679 (N_24679,N_18607,N_18265);
xnor U24680 (N_24680,N_15069,N_17666);
nand U24681 (N_24681,N_19383,N_19877);
or U24682 (N_24682,N_16085,N_16077);
and U24683 (N_24683,N_16907,N_18561);
nand U24684 (N_24684,N_19738,N_19522);
xor U24685 (N_24685,N_15434,N_19429);
xor U24686 (N_24686,N_18317,N_16076);
nand U24687 (N_24687,N_15509,N_17420);
xnor U24688 (N_24688,N_15712,N_19458);
or U24689 (N_24689,N_17822,N_17285);
nor U24690 (N_24690,N_17032,N_15132);
nor U24691 (N_24691,N_18083,N_19650);
nor U24692 (N_24692,N_17180,N_18051);
or U24693 (N_24693,N_15106,N_17090);
xor U24694 (N_24694,N_15696,N_17534);
nor U24695 (N_24695,N_17670,N_15817);
or U24696 (N_24696,N_15470,N_18010);
and U24697 (N_24697,N_17211,N_16788);
or U24698 (N_24698,N_18735,N_16130);
or U24699 (N_24699,N_19998,N_15310);
or U24700 (N_24700,N_15394,N_16950);
and U24701 (N_24701,N_17603,N_19099);
xor U24702 (N_24702,N_17661,N_15121);
nor U24703 (N_24703,N_17827,N_18485);
and U24704 (N_24704,N_15618,N_19579);
and U24705 (N_24705,N_15184,N_18972);
nand U24706 (N_24706,N_19142,N_18903);
xnor U24707 (N_24707,N_15701,N_18893);
nor U24708 (N_24708,N_15951,N_15901);
nand U24709 (N_24709,N_17590,N_18370);
or U24710 (N_24710,N_16632,N_16457);
and U24711 (N_24711,N_19357,N_18694);
and U24712 (N_24712,N_18528,N_18963);
or U24713 (N_24713,N_18534,N_15434);
xnor U24714 (N_24714,N_19741,N_15723);
nor U24715 (N_24715,N_17638,N_18349);
nor U24716 (N_24716,N_19560,N_16395);
nand U24717 (N_24717,N_15939,N_16762);
and U24718 (N_24718,N_15437,N_16089);
and U24719 (N_24719,N_18205,N_15207);
and U24720 (N_24720,N_18941,N_18560);
or U24721 (N_24721,N_17687,N_17958);
and U24722 (N_24722,N_17314,N_19027);
xor U24723 (N_24723,N_19961,N_19069);
nor U24724 (N_24724,N_18761,N_17097);
xor U24725 (N_24725,N_18836,N_19330);
xor U24726 (N_24726,N_16660,N_16637);
or U24727 (N_24727,N_16918,N_19105);
nor U24728 (N_24728,N_15688,N_15437);
nand U24729 (N_24729,N_16357,N_18635);
nor U24730 (N_24730,N_16180,N_18318);
nand U24731 (N_24731,N_16856,N_18699);
or U24732 (N_24732,N_17020,N_17525);
nor U24733 (N_24733,N_17686,N_17840);
nand U24734 (N_24734,N_16357,N_16056);
nor U24735 (N_24735,N_16549,N_17263);
xnor U24736 (N_24736,N_15135,N_17586);
and U24737 (N_24737,N_15668,N_17541);
nor U24738 (N_24738,N_16799,N_19608);
and U24739 (N_24739,N_18268,N_18733);
nor U24740 (N_24740,N_19695,N_17225);
nand U24741 (N_24741,N_16842,N_17769);
nor U24742 (N_24742,N_15896,N_15174);
nand U24743 (N_24743,N_17798,N_15263);
and U24744 (N_24744,N_15910,N_18556);
xor U24745 (N_24745,N_15935,N_15788);
nand U24746 (N_24746,N_15385,N_16008);
xnor U24747 (N_24747,N_16838,N_19256);
or U24748 (N_24748,N_17538,N_16694);
and U24749 (N_24749,N_17887,N_18010);
nor U24750 (N_24750,N_18068,N_19425);
or U24751 (N_24751,N_17207,N_16606);
or U24752 (N_24752,N_16134,N_17341);
nand U24753 (N_24753,N_19388,N_17895);
and U24754 (N_24754,N_17786,N_15993);
or U24755 (N_24755,N_19885,N_19898);
nand U24756 (N_24756,N_17916,N_19815);
nor U24757 (N_24757,N_19856,N_18125);
and U24758 (N_24758,N_19557,N_16887);
nor U24759 (N_24759,N_15841,N_15920);
nor U24760 (N_24760,N_17511,N_19779);
nand U24761 (N_24761,N_15366,N_16231);
and U24762 (N_24762,N_19367,N_19504);
nor U24763 (N_24763,N_15199,N_16816);
or U24764 (N_24764,N_17907,N_16200);
xor U24765 (N_24765,N_17103,N_16281);
nor U24766 (N_24766,N_18693,N_19869);
xor U24767 (N_24767,N_19717,N_15334);
xnor U24768 (N_24768,N_18226,N_16404);
or U24769 (N_24769,N_18075,N_17953);
or U24770 (N_24770,N_15198,N_19544);
nand U24771 (N_24771,N_17786,N_16803);
xnor U24772 (N_24772,N_17161,N_15292);
or U24773 (N_24773,N_17166,N_15154);
nand U24774 (N_24774,N_18012,N_15578);
xnor U24775 (N_24775,N_18715,N_16081);
xnor U24776 (N_24776,N_17564,N_15705);
xnor U24777 (N_24777,N_15912,N_15467);
nand U24778 (N_24778,N_16889,N_16688);
and U24779 (N_24779,N_16720,N_17964);
nand U24780 (N_24780,N_19838,N_18873);
nand U24781 (N_24781,N_16069,N_19856);
and U24782 (N_24782,N_16187,N_17354);
or U24783 (N_24783,N_16623,N_17683);
and U24784 (N_24784,N_19984,N_17220);
nand U24785 (N_24785,N_16474,N_18405);
xor U24786 (N_24786,N_19936,N_19964);
or U24787 (N_24787,N_19421,N_15041);
or U24788 (N_24788,N_18314,N_19611);
nand U24789 (N_24789,N_16795,N_19215);
nand U24790 (N_24790,N_19085,N_18217);
nand U24791 (N_24791,N_16642,N_17423);
and U24792 (N_24792,N_15649,N_16453);
or U24793 (N_24793,N_18145,N_16500);
or U24794 (N_24794,N_16228,N_19746);
nor U24795 (N_24795,N_18585,N_16675);
xor U24796 (N_24796,N_16034,N_18380);
or U24797 (N_24797,N_15757,N_15170);
nand U24798 (N_24798,N_18475,N_17680);
and U24799 (N_24799,N_15854,N_15058);
nand U24800 (N_24800,N_15486,N_17740);
nor U24801 (N_24801,N_17109,N_17481);
xnor U24802 (N_24802,N_17221,N_15211);
nand U24803 (N_24803,N_18678,N_18941);
nand U24804 (N_24804,N_18688,N_17672);
and U24805 (N_24805,N_17070,N_15562);
xor U24806 (N_24806,N_17317,N_15700);
nor U24807 (N_24807,N_19591,N_16475);
xnor U24808 (N_24808,N_18238,N_18003);
nor U24809 (N_24809,N_15388,N_17370);
and U24810 (N_24810,N_19301,N_17259);
xnor U24811 (N_24811,N_16881,N_19331);
nand U24812 (N_24812,N_18558,N_17209);
nand U24813 (N_24813,N_16095,N_17800);
xor U24814 (N_24814,N_15340,N_16801);
and U24815 (N_24815,N_16372,N_16541);
nor U24816 (N_24816,N_18117,N_15299);
and U24817 (N_24817,N_16526,N_16653);
xor U24818 (N_24818,N_16070,N_19026);
nand U24819 (N_24819,N_15089,N_17737);
or U24820 (N_24820,N_18050,N_15572);
nor U24821 (N_24821,N_19241,N_16110);
and U24822 (N_24822,N_16422,N_19312);
and U24823 (N_24823,N_15644,N_17723);
and U24824 (N_24824,N_18845,N_18725);
and U24825 (N_24825,N_19680,N_16521);
nor U24826 (N_24826,N_16846,N_18226);
nor U24827 (N_24827,N_18024,N_15964);
nor U24828 (N_24828,N_18944,N_16806);
and U24829 (N_24829,N_17223,N_17727);
nand U24830 (N_24830,N_19691,N_15638);
nor U24831 (N_24831,N_19190,N_17784);
nor U24832 (N_24832,N_16925,N_18581);
and U24833 (N_24833,N_19907,N_19060);
and U24834 (N_24834,N_17114,N_18468);
xor U24835 (N_24835,N_19967,N_15365);
nor U24836 (N_24836,N_17583,N_19178);
nor U24837 (N_24837,N_16120,N_17621);
or U24838 (N_24838,N_16311,N_15305);
nand U24839 (N_24839,N_18329,N_18423);
and U24840 (N_24840,N_16047,N_18438);
nand U24841 (N_24841,N_18674,N_19625);
nor U24842 (N_24842,N_18439,N_16514);
nand U24843 (N_24843,N_16425,N_19391);
xnor U24844 (N_24844,N_17785,N_15078);
nand U24845 (N_24845,N_17562,N_15963);
or U24846 (N_24846,N_19141,N_15306);
and U24847 (N_24847,N_18815,N_17100);
nand U24848 (N_24848,N_16960,N_16110);
and U24849 (N_24849,N_18478,N_17011);
or U24850 (N_24850,N_19443,N_16208);
nor U24851 (N_24851,N_19877,N_15896);
nand U24852 (N_24852,N_16270,N_18669);
and U24853 (N_24853,N_18075,N_18257);
and U24854 (N_24854,N_19026,N_19629);
xnor U24855 (N_24855,N_18923,N_18798);
or U24856 (N_24856,N_17405,N_19729);
xnor U24857 (N_24857,N_15073,N_15915);
and U24858 (N_24858,N_15285,N_18189);
or U24859 (N_24859,N_16304,N_17643);
nor U24860 (N_24860,N_18389,N_15579);
xor U24861 (N_24861,N_15715,N_19173);
xor U24862 (N_24862,N_16082,N_18990);
or U24863 (N_24863,N_18822,N_19623);
nor U24864 (N_24864,N_17404,N_16600);
or U24865 (N_24865,N_17485,N_17530);
or U24866 (N_24866,N_17659,N_19821);
and U24867 (N_24867,N_19047,N_16696);
xnor U24868 (N_24868,N_19563,N_15658);
and U24869 (N_24869,N_19097,N_15311);
or U24870 (N_24870,N_18496,N_15897);
or U24871 (N_24871,N_19392,N_18416);
and U24872 (N_24872,N_15400,N_17953);
nor U24873 (N_24873,N_16600,N_15492);
nand U24874 (N_24874,N_16362,N_18348);
or U24875 (N_24875,N_15744,N_19120);
nand U24876 (N_24876,N_16521,N_18523);
xor U24877 (N_24877,N_17108,N_18923);
and U24878 (N_24878,N_18861,N_15011);
xnor U24879 (N_24879,N_19036,N_16763);
nand U24880 (N_24880,N_18580,N_17661);
and U24881 (N_24881,N_15053,N_17346);
or U24882 (N_24882,N_18976,N_19523);
and U24883 (N_24883,N_16001,N_17970);
and U24884 (N_24884,N_19643,N_18738);
nor U24885 (N_24885,N_17925,N_18482);
and U24886 (N_24886,N_18612,N_16634);
nand U24887 (N_24887,N_15238,N_18548);
and U24888 (N_24888,N_16052,N_16838);
or U24889 (N_24889,N_16723,N_19992);
and U24890 (N_24890,N_17786,N_17762);
nand U24891 (N_24891,N_19159,N_18485);
nand U24892 (N_24892,N_18981,N_15954);
nor U24893 (N_24893,N_17699,N_15330);
nand U24894 (N_24894,N_18387,N_15177);
or U24895 (N_24895,N_18548,N_17841);
nand U24896 (N_24896,N_17404,N_15574);
or U24897 (N_24897,N_17247,N_19951);
xor U24898 (N_24898,N_17868,N_18209);
or U24899 (N_24899,N_17107,N_16854);
or U24900 (N_24900,N_18782,N_16876);
nor U24901 (N_24901,N_16571,N_19469);
xnor U24902 (N_24902,N_18907,N_18879);
nor U24903 (N_24903,N_18523,N_15036);
xnor U24904 (N_24904,N_17629,N_15797);
or U24905 (N_24905,N_18854,N_15540);
nand U24906 (N_24906,N_15561,N_16859);
nand U24907 (N_24907,N_17910,N_15187);
or U24908 (N_24908,N_16192,N_18383);
and U24909 (N_24909,N_17300,N_17202);
and U24910 (N_24910,N_17120,N_19850);
xnor U24911 (N_24911,N_17698,N_19300);
xor U24912 (N_24912,N_15215,N_16823);
nand U24913 (N_24913,N_16617,N_15222);
nand U24914 (N_24914,N_19726,N_19282);
or U24915 (N_24915,N_15948,N_15738);
nor U24916 (N_24916,N_15962,N_19038);
nor U24917 (N_24917,N_18972,N_19844);
or U24918 (N_24918,N_19911,N_18807);
nand U24919 (N_24919,N_19856,N_15061);
xnor U24920 (N_24920,N_19184,N_17625);
and U24921 (N_24921,N_17434,N_19026);
or U24922 (N_24922,N_17101,N_18117);
xnor U24923 (N_24923,N_16791,N_17351);
xor U24924 (N_24924,N_16027,N_17652);
and U24925 (N_24925,N_15267,N_19538);
and U24926 (N_24926,N_19442,N_18915);
or U24927 (N_24927,N_19109,N_15055);
xnor U24928 (N_24928,N_16363,N_16501);
or U24929 (N_24929,N_15427,N_15528);
nor U24930 (N_24930,N_17931,N_15643);
nor U24931 (N_24931,N_18973,N_17254);
or U24932 (N_24932,N_17204,N_18139);
or U24933 (N_24933,N_15024,N_18515);
xnor U24934 (N_24934,N_16905,N_18741);
xor U24935 (N_24935,N_18803,N_19344);
xnor U24936 (N_24936,N_15752,N_17050);
xor U24937 (N_24937,N_16842,N_17756);
nand U24938 (N_24938,N_18649,N_18706);
or U24939 (N_24939,N_15582,N_16481);
nor U24940 (N_24940,N_18060,N_19641);
or U24941 (N_24941,N_16053,N_18732);
nand U24942 (N_24942,N_19384,N_18303);
and U24943 (N_24943,N_18383,N_19208);
nor U24944 (N_24944,N_18665,N_17985);
xor U24945 (N_24945,N_17724,N_19030);
and U24946 (N_24946,N_16587,N_16896);
nor U24947 (N_24947,N_17922,N_15427);
and U24948 (N_24948,N_18903,N_16222);
nor U24949 (N_24949,N_18688,N_17597);
xnor U24950 (N_24950,N_19738,N_18771);
xor U24951 (N_24951,N_15989,N_18251);
xnor U24952 (N_24952,N_18664,N_17372);
xor U24953 (N_24953,N_15813,N_17634);
and U24954 (N_24954,N_19430,N_17562);
xor U24955 (N_24955,N_18173,N_18106);
or U24956 (N_24956,N_16715,N_18538);
xnor U24957 (N_24957,N_19973,N_16507);
or U24958 (N_24958,N_17519,N_15167);
nor U24959 (N_24959,N_15165,N_16454);
xnor U24960 (N_24960,N_15362,N_16277);
nor U24961 (N_24961,N_15303,N_18566);
and U24962 (N_24962,N_19786,N_15440);
nor U24963 (N_24963,N_17587,N_19639);
and U24964 (N_24964,N_17398,N_15204);
nor U24965 (N_24965,N_18812,N_16161);
nand U24966 (N_24966,N_18352,N_18637);
nand U24967 (N_24967,N_17312,N_16203);
or U24968 (N_24968,N_17824,N_15219);
xnor U24969 (N_24969,N_16859,N_16554);
and U24970 (N_24970,N_19319,N_15605);
xnor U24971 (N_24971,N_15438,N_15650);
nand U24972 (N_24972,N_15676,N_15530);
nand U24973 (N_24973,N_19482,N_15072);
nand U24974 (N_24974,N_17092,N_17978);
nor U24975 (N_24975,N_19485,N_18110);
or U24976 (N_24976,N_19637,N_18983);
or U24977 (N_24977,N_15415,N_16329);
or U24978 (N_24978,N_19194,N_15394);
nor U24979 (N_24979,N_18742,N_18684);
xor U24980 (N_24980,N_18712,N_19366);
and U24981 (N_24981,N_16222,N_18522);
nor U24982 (N_24982,N_18494,N_16256);
xnor U24983 (N_24983,N_15572,N_19911);
nand U24984 (N_24984,N_17120,N_18108);
xnor U24985 (N_24985,N_17933,N_16138);
nor U24986 (N_24986,N_16337,N_19082);
or U24987 (N_24987,N_19210,N_19500);
nand U24988 (N_24988,N_16274,N_17652);
xor U24989 (N_24989,N_17533,N_15617);
and U24990 (N_24990,N_16066,N_17378);
and U24991 (N_24991,N_17197,N_19659);
nand U24992 (N_24992,N_18340,N_16528);
and U24993 (N_24993,N_16565,N_16828);
nand U24994 (N_24994,N_18756,N_17819);
xor U24995 (N_24995,N_15217,N_15215);
nor U24996 (N_24996,N_17624,N_17052);
xor U24997 (N_24997,N_17148,N_17814);
xor U24998 (N_24998,N_16956,N_16534);
nand U24999 (N_24999,N_15775,N_17141);
or UO_0 (O_0,N_23445,N_22762);
or UO_1 (O_1,N_24740,N_24496);
nand UO_2 (O_2,N_24206,N_24352);
nand UO_3 (O_3,N_22019,N_22795);
or UO_4 (O_4,N_23980,N_22985);
or UO_5 (O_5,N_23649,N_22630);
and UO_6 (O_6,N_24945,N_20456);
or UO_7 (O_7,N_23269,N_20614);
nand UO_8 (O_8,N_24299,N_24597);
and UO_9 (O_9,N_21168,N_20340);
and UO_10 (O_10,N_21159,N_21278);
nor UO_11 (O_11,N_23036,N_24116);
nor UO_12 (O_12,N_23519,N_22501);
nor UO_13 (O_13,N_23994,N_23418);
xor UO_14 (O_14,N_22754,N_21678);
xnor UO_15 (O_15,N_22141,N_23689);
or UO_16 (O_16,N_23085,N_21976);
xnor UO_17 (O_17,N_22392,N_23338);
nand UO_18 (O_18,N_22743,N_21876);
and UO_19 (O_19,N_22022,N_23640);
xnor UO_20 (O_20,N_23206,N_24713);
and UO_21 (O_21,N_24710,N_20164);
xor UO_22 (O_22,N_22923,N_22265);
or UO_23 (O_23,N_21936,N_24984);
nand UO_24 (O_24,N_21785,N_24526);
nand UO_25 (O_25,N_21747,N_23196);
or UO_26 (O_26,N_24800,N_24195);
nor UO_27 (O_27,N_21540,N_22473);
nand UO_28 (O_28,N_21194,N_20512);
and UO_29 (O_29,N_20566,N_20243);
nor UO_30 (O_30,N_24636,N_20106);
nor UO_31 (O_31,N_24432,N_22662);
nor UO_32 (O_32,N_21469,N_22936);
and UO_33 (O_33,N_22469,N_23956);
nor UO_34 (O_34,N_23149,N_22775);
xnor UO_35 (O_35,N_21077,N_21686);
xnor UO_36 (O_36,N_22316,N_20572);
and UO_37 (O_37,N_22143,N_24276);
nand UO_38 (O_38,N_23897,N_22162);
or UO_39 (O_39,N_22812,N_20709);
nor UO_40 (O_40,N_24825,N_21072);
and UO_41 (O_41,N_20540,N_24971);
nand UO_42 (O_42,N_23024,N_21724);
nand UO_43 (O_43,N_22319,N_22899);
nand UO_44 (O_44,N_22541,N_21738);
nand UO_45 (O_45,N_22941,N_23840);
or UO_46 (O_46,N_20182,N_24780);
or UO_47 (O_47,N_21269,N_21066);
and UO_48 (O_48,N_24463,N_23458);
and UO_49 (O_49,N_20029,N_22303);
nand UO_50 (O_50,N_23314,N_21277);
or UO_51 (O_51,N_20798,N_22921);
nand UO_52 (O_52,N_22651,N_24030);
nand UO_53 (O_53,N_24831,N_24524);
nand UO_54 (O_54,N_22515,N_23611);
xnor UO_55 (O_55,N_20660,N_20414);
nor UO_56 (O_56,N_24674,N_24689);
nor UO_57 (O_57,N_22197,N_24509);
and UO_58 (O_58,N_24684,N_20543);
or UO_59 (O_59,N_20365,N_20191);
nand UO_60 (O_60,N_23921,N_21948);
nand UO_61 (O_61,N_22081,N_22067);
and UO_62 (O_62,N_20311,N_24832);
or UO_63 (O_63,N_21821,N_22677);
and UO_64 (O_64,N_20576,N_23336);
and UO_65 (O_65,N_23126,N_24391);
nand UO_66 (O_66,N_23614,N_21103);
and UO_67 (O_67,N_22522,N_20315);
xor UO_68 (O_68,N_20948,N_22011);
and UO_69 (O_69,N_21842,N_22159);
nor UO_70 (O_70,N_21388,N_20330);
and UO_71 (O_71,N_20523,N_24819);
and UO_72 (O_72,N_24586,N_21007);
nand UO_73 (O_73,N_23597,N_24686);
xnor UO_74 (O_74,N_20482,N_24326);
and UO_75 (O_75,N_23089,N_22183);
nor UO_76 (O_76,N_21728,N_20210);
nand UO_77 (O_77,N_23226,N_21954);
or UO_78 (O_78,N_20908,N_24778);
nor UO_79 (O_79,N_20617,N_24731);
and UO_80 (O_80,N_20720,N_23411);
nor UO_81 (O_81,N_20701,N_22598);
xnor UO_82 (O_82,N_21105,N_24540);
and UO_83 (O_83,N_24409,N_23742);
or UO_84 (O_84,N_20355,N_24988);
nor UO_85 (O_85,N_24098,N_21493);
xor UO_86 (O_86,N_24578,N_20295);
nand UO_87 (O_87,N_22784,N_20789);
nor UO_88 (O_88,N_20273,N_23214);
or UO_89 (O_89,N_23243,N_23617);
nor UO_90 (O_90,N_23057,N_24477);
nor UO_91 (O_91,N_23694,N_24124);
nand UO_92 (O_92,N_24161,N_20139);
nor UO_93 (O_93,N_22916,N_23761);
and UO_94 (O_94,N_22157,N_21380);
nand UO_95 (O_95,N_23008,N_23468);
nor UO_96 (O_96,N_23238,N_20494);
and UO_97 (O_97,N_23317,N_24271);
and UO_98 (O_98,N_20577,N_20929);
nand UO_99 (O_99,N_22909,N_24753);
or UO_100 (O_100,N_22770,N_21143);
and UO_101 (O_101,N_24628,N_22570);
nor UO_102 (O_102,N_20889,N_22792);
or UO_103 (O_103,N_23902,N_23855);
and UO_104 (O_104,N_24986,N_21695);
or UO_105 (O_105,N_20940,N_23670);
nor UO_106 (O_106,N_24305,N_21795);
nor UO_107 (O_107,N_22969,N_21802);
nor UO_108 (O_108,N_23114,N_22602);
and UO_109 (O_109,N_22978,N_21122);
or UO_110 (O_110,N_20187,N_23178);
nand UO_111 (O_111,N_20035,N_23863);
nor UO_112 (O_112,N_21155,N_20080);
or UO_113 (O_113,N_23351,N_23822);
nor UO_114 (O_114,N_23699,N_20214);
and UO_115 (O_115,N_23661,N_24658);
nand UO_116 (O_116,N_23450,N_24732);
or UO_117 (O_117,N_21710,N_22305);
nand UO_118 (O_118,N_24282,N_21457);
nand UO_119 (O_119,N_24908,N_23015);
and UO_120 (O_120,N_21858,N_21767);
nand UO_121 (O_121,N_21083,N_24422);
nand UO_122 (O_122,N_21619,N_21133);
and UO_123 (O_123,N_20163,N_23010);
and UO_124 (O_124,N_23028,N_23281);
nand UO_125 (O_125,N_20670,N_22358);
nor UO_126 (O_126,N_20902,N_23211);
and UO_127 (O_127,N_23213,N_20329);
nor UO_128 (O_128,N_22235,N_21176);
xor UO_129 (O_129,N_20082,N_20400);
nand UO_130 (O_130,N_21222,N_21937);
or UO_131 (O_131,N_21885,N_20338);
nor UO_132 (O_132,N_22706,N_23716);
and UO_133 (O_133,N_22510,N_20955);
or UO_134 (O_134,N_21193,N_24991);
nor UO_135 (O_135,N_23282,N_24528);
or UO_136 (O_136,N_20802,N_23539);
xor UO_137 (O_137,N_22790,N_21209);
nor UO_138 (O_138,N_22359,N_20057);
or UO_139 (O_139,N_20774,N_23273);
or UO_140 (O_140,N_24965,N_20917);
or UO_141 (O_141,N_24789,N_21171);
nor UO_142 (O_142,N_23465,N_23684);
or UO_143 (O_143,N_24469,N_21572);
xor UO_144 (O_144,N_24699,N_22003);
and UO_145 (O_145,N_20168,N_21129);
xor UO_146 (O_146,N_23722,N_23678);
or UO_147 (O_147,N_22029,N_23557);
and UO_148 (O_148,N_23477,N_22326);
or UO_149 (O_149,N_22604,N_24899);
nor UO_150 (O_150,N_20140,N_23601);
nor UO_151 (O_151,N_24748,N_21512);
nand UO_152 (O_152,N_23785,N_24176);
nor UO_153 (O_153,N_21242,N_22001);
nand UO_154 (O_154,N_21662,N_22256);
or UO_155 (O_155,N_22491,N_23866);
or UO_156 (O_156,N_21900,N_23462);
nand UO_157 (O_157,N_20396,N_24203);
nand UO_158 (O_158,N_23886,N_23032);
and UO_159 (O_159,N_24004,N_22713);
nor UO_160 (O_160,N_21480,N_21568);
xor UO_161 (O_161,N_24256,N_22877);
nor UO_162 (O_162,N_23412,N_22467);
xor UO_163 (O_163,N_20599,N_20552);
or UO_164 (O_164,N_22903,N_23603);
or UO_165 (O_165,N_23847,N_23975);
or UO_166 (O_166,N_21106,N_22328);
and UO_167 (O_167,N_20108,N_22454);
nand UO_168 (O_168,N_21509,N_22149);
xor UO_169 (O_169,N_22874,N_23755);
xnor UO_170 (O_170,N_24095,N_24898);
xor UO_171 (O_171,N_22079,N_22481);
nor UO_172 (O_172,N_23311,N_23109);
nand UO_173 (O_173,N_24723,N_24452);
and UO_174 (O_174,N_24428,N_21889);
and UO_175 (O_175,N_20522,N_23147);
nand UO_176 (O_176,N_23294,N_20370);
xor UO_177 (O_177,N_22951,N_23826);
nand UO_178 (O_178,N_23033,N_23359);
and UO_179 (O_179,N_21350,N_22082);
xnor UO_180 (O_180,N_23594,N_22933);
xnor UO_181 (O_181,N_20287,N_22184);
or UO_182 (O_182,N_23307,N_20706);
nor UO_183 (O_183,N_22724,N_20553);
xor UO_184 (O_184,N_23838,N_20356);
or UO_185 (O_185,N_20195,N_21854);
nor UO_186 (O_186,N_22756,N_20764);
and UO_187 (O_187,N_22374,N_22823);
or UO_188 (O_188,N_22172,N_22869);
and UO_189 (O_189,N_22946,N_20631);
and UO_190 (O_190,N_21893,N_22656);
or UO_191 (O_191,N_22593,N_20111);
and UO_192 (O_192,N_20977,N_22649);
or UO_193 (O_193,N_21386,N_23466);
xor UO_194 (O_194,N_22796,N_22659);
and UO_195 (O_195,N_23854,N_20419);
and UO_196 (O_196,N_21487,N_21593);
or UO_197 (O_197,N_20823,N_21605);
and UO_198 (O_198,N_20067,N_20876);
or UO_199 (O_199,N_23786,N_23917);
nand UO_200 (O_200,N_21684,N_24237);
xnor UO_201 (O_201,N_21217,N_21624);
or UO_202 (O_202,N_23616,N_24358);
or UO_203 (O_203,N_22420,N_20162);
or UO_204 (O_204,N_24716,N_24869);
nor UO_205 (O_205,N_21729,N_24601);
or UO_206 (O_206,N_24475,N_20833);
nor UO_207 (O_207,N_20816,N_21573);
or UO_208 (O_208,N_24870,N_21363);
nand UO_209 (O_209,N_21816,N_21049);
and UO_210 (O_210,N_20367,N_23434);
and UO_211 (O_211,N_24360,N_22477);
nand UO_212 (O_212,N_21846,N_23662);
nor UO_213 (O_213,N_23787,N_23582);
nand UO_214 (O_214,N_20705,N_23623);
nand UO_215 (O_215,N_24361,N_22448);
nand UO_216 (O_216,N_24793,N_24479);
nand UO_217 (O_217,N_24472,N_22311);
nand UO_218 (O_218,N_23610,N_21266);
xor UO_219 (O_219,N_20885,N_23518);
nor UO_220 (O_220,N_24097,N_23306);
and UO_221 (O_221,N_24289,N_23808);
xnor UO_222 (O_222,N_20272,N_21836);
or UO_223 (O_223,N_24523,N_23467);
xor UO_224 (O_224,N_23259,N_20933);
and UO_225 (O_225,N_22304,N_23127);
or UO_226 (O_226,N_22548,N_20749);
nand UO_227 (O_227,N_23774,N_21904);
or UO_228 (O_228,N_21272,N_24955);
nor UO_229 (O_229,N_24756,N_23816);
nand UO_230 (O_230,N_20403,N_23235);
or UO_231 (O_231,N_23247,N_24070);
nand UO_232 (O_232,N_22318,N_20151);
xnor UO_233 (O_233,N_21886,N_23288);
nand UO_234 (O_234,N_22410,N_22308);
nor UO_235 (O_235,N_23343,N_20770);
and UO_236 (O_236,N_24721,N_24633);
nor UO_237 (O_237,N_22582,N_24579);
xor UO_238 (O_238,N_22956,N_22924);
nand UO_239 (O_239,N_20381,N_20918);
or UO_240 (O_240,N_24719,N_24212);
xor UO_241 (O_241,N_23421,N_24934);
or UO_242 (O_242,N_23179,N_21742);
xnor UO_243 (O_243,N_23334,N_20406);
or UO_244 (O_244,N_23102,N_21622);
xnor UO_245 (O_245,N_20483,N_22574);
and UO_246 (O_246,N_24649,N_24390);
nand UO_247 (O_247,N_20775,N_24112);
nand UO_248 (O_248,N_21851,N_20817);
xor UO_249 (O_249,N_23970,N_22834);
or UO_250 (O_250,N_23455,N_20430);
xnor UO_251 (O_251,N_23645,N_20286);
xnor UO_252 (O_252,N_20422,N_21008);
and UO_253 (O_253,N_22664,N_22616);
nand UO_254 (O_254,N_23644,N_21183);
xor UO_255 (O_255,N_20107,N_20088);
and UO_256 (O_256,N_21553,N_20294);
nor UO_257 (O_257,N_24291,N_22204);
or UO_258 (O_258,N_21204,N_20761);
nand UO_259 (O_259,N_20208,N_23497);
xor UO_260 (O_260,N_22538,N_23885);
nor UO_261 (O_261,N_23734,N_20193);
or UO_262 (O_262,N_20820,N_24013);
xnor UO_263 (O_263,N_23471,N_21303);
nor UO_264 (O_264,N_21567,N_20507);
xnor UO_265 (O_265,N_20450,N_24916);
nor UO_266 (O_266,N_24425,N_20492);
and UO_267 (O_267,N_23927,N_22729);
nand UO_268 (O_268,N_21670,N_23055);
xnor UO_269 (O_269,N_22803,N_23919);
and UO_270 (O_270,N_20550,N_23398);
nor UO_271 (O_271,N_21446,N_20136);
nand UO_272 (O_272,N_24108,N_22105);
or UO_273 (O_273,N_21470,N_22334);
nor UO_274 (O_274,N_21507,N_20958);
or UO_275 (O_275,N_20763,N_24808);
or UO_276 (O_276,N_21216,N_21454);
or UO_277 (O_277,N_24368,N_24244);
nor UO_278 (O_278,N_21781,N_20649);
or UO_279 (O_279,N_21826,N_21245);
or UO_280 (O_280,N_20443,N_20711);
or UO_281 (O_281,N_24940,N_22161);
and UO_282 (O_282,N_24111,N_22737);
or UO_283 (O_283,N_24198,N_21319);
nand UO_284 (O_284,N_22250,N_20575);
nor UO_285 (O_285,N_20063,N_21474);
nor UO_286 (O_286,N_21806,N_20344);
and UO_287 (O_287,N_23187,N_22036);
nand UO_288 (O_288,N_24053,N_24419);
and UO_289 (O_289,N_24412,N_21974);
nor UO_290 (O_290,N_20801,N_23945);
and UO_291 (O_291,N_20594,N_23168);
nand UO_292 (O_292,N_21950,N_23503);
xor UO_293 (O_293,N_22258,N_24169);
and UO_294 (O_294,N_20228,N_21790);
xor UO_295 (O_295,N_20987,N_24541);
and UO_296 (O_296,N_20846,N_23331);
xor UO_297 (O_297,N_20203,N_20409);
or UO_298 (O_298,N_23170,N_24671);
nand UO_299 (O_299,N_22399,N_21513);
and UO_300 (O_300,N_24734,N_23498);
or UO_301 (O_301,N_24424,N_21448);
nand UO_302 (O_302,N_24277,N_22479);
xnor UO_303 (O_303,N_24459,N_23797);
nor UO_304 (O_304,N_24338,N_24529);
nor UO_305 (O_305,N_20015,N_21005);
nor UO_306 (O_306,N_23749,N_24351);
or UO_307 (O_307,N_21125,N_22727);
xnor UO_308 (O_308,N_20290,N_24417);
xnor UO_309 (O_309,N_21418,N_24829);
nor UO_310 (O_310,N_22460,N_24458);
or UO_311 (O_311,N_21255,N_22094);
nor UO_312 (O_312,N_21855,N_24306);
and UO_313 (O_313,N_24598,N_20873);
nand UO_314 (O_314,N_21014,N_22742);
nand UO_315 (O_315,N_22698,N_20983);
or UO_316 (O_316,N_22802,N_20531);
nand UO_317 (O_317,N_23612,N_23845);
and UO_318 (O_318,N_22181,N_21748);
nand UO_319 (O_319,N_24345,N_22275);
or UO_320 (O_320,N_20473,N_23002);
or UO_321 (O_321,N_21656,N_20138);
nor UO_322 (O_322,N_20903,N_23704);
nor UO_323 (O_323,N_24830,N_24947);
xnor UO_324 (O_324,N_20514,N_23884);
and UO_325 (O_325,N_20255,N_20325);
nor UO_326 (O_326,N_23150,N_24199);
or UO_327 (O_327,N_23874,N_23739);
and UO_328 (O_328,N_21249,N_24373);
nand UO_329 (O_329,N_22786,N_23744);
or UO_330 (O_330,N_23925,N_23373);
xnor UO_331 (O_331,N_21555,N_24784);
xnor UO_332 (O_332,N_23263,N_22794);
or UO_333 (O_333,N_23248,N_24269);
nand UO_334 (O_334,N_23345,N_23789);
nor UO_335 (O_335,N_23758,N_22290);
nor UO_336 (O_336,N_22405,N_21978);
xnor UO_337 (O_337,N_24733,N_23773);
or UO_338 (O_338,N_20538,N_22382);
or UO_339 (O_339,N_21765,N_20056);
xnor UO_340 (O_340,N_21931,N_20232);
or UO_341 (O_341,N_23949,N_24905);
nor UO_342 (O_342,N_21867,N_20094);
nand UO_343 (O_343,N_23839,N_21101);
nor UO_344 (O_344,N_21685,N_22043);
nor UO_345 (O_345,N_23501,N_24284);
nor UO_346 (O_346,N_21707,N_21680);
or UO_347 (O_347,N_23242,N_22063);
or UO_348 (O_348,N_22870,N_23958);
xor UO_349 (O_349,N_21334,N_24331);
and UO_350 (O_350,N_22988,N_23889);
and UO_351 (O_351,N_20744,N_21651);
or UO_352 (O_352,N_23271,N_20839);
nor UO_353 (O_353,N_21726,N_21840);
nor UO_354 (O_354,N_21276,N_22831);
or UO_355 (O_355,N_23953,N_22010);
or UO_356 (O_356,N_24669,N_20612);
and UO_357 (O_357,N_20464,N_21382);
nand UO_358 (O_358,N_21818,N_24514);
xnor UO_359 (O_359,N_22156,N_20375);
or UO_360 (O_360,N_21231,N_22125);
nor UO_361 (O_361,N_21482,N_20662);
nor UO_362 (O_362,N_24103,N_21238);
or UO_363 (O_363,N_20336,N_24446);
nand UO_364 (O_364,N_24127,N_23449);
nand UO_365 (O_365,N_21672,N_21391);
nand UO_366 (O_366,N_23510,N_22196);
and UO_367 (O_367,N_23129,N_23965);
and UO_368 (O_368,N_24895,N_22563);
nor UO_369 (O_369,N_21475,N_22521);
nand UO_370 (O_370,N_23872,N_22338);
nor UO_371 (O_371,N_20461,N_23066);
and UO_372 (O_372,N_23194,N_22363);
nand UO_373 (O_373,N_21705,N_23375);
nor UO_374 (O_374,N_21863,N_22816);
nand UO_375 (O_375,N_20233,N_22723);
xor UO_376 (O_376,N_21723,N_23976);
nor UO_377 (O_377,N_23309,N_22587);
nand UO_378 (O_378,N_21299,N_22132);
nand UO_379 (O_379,N_24182,N_23829);
nor UO_380 (O_380,N_22503,N_21527);
nand UO_381 (O_381,N_21988,N_23298);
or UO_382 (O_382,N_21288,N_22280);
or UO_383 (O_383,N_23183,N_20048);
nand UO_384 (O_384,N_22212,N_21092);
or UO_385 (O_385,N_22401,N_20758);
and UO_386 (O_386,N_20387,N_20361);
and UO_387 (O_387,N_23481,N_22785);
xor UO_388 (O_388,N_24208,N_24516);
nor UO_389 (O_389,N_20410,N_20073);
xnor UO_390 (O_390,N_22842,N_21692);
or UO_391 (O_391,N_21616,N_23365);
xnor UO_392 (O_392,N_22767,N_22342);
xnor UO_393 (O_393,N_20326,N_21901);
xor UO_394 (O_394,N_21773,N_20352);
or UO_395 (O_395,N_23636,N_24925);
nand UO_396 (O_396,N_24755,N_22669);
or UO_397 (O_397,N_22053,N_23723);
xor UO_398 (O_398,N_22252,N_24462);
nor UO_399 (O_399,N_24726,N_22822);
or UO_400 (O_400,N_24063,N_23220);
nor UO_401 (O_401,N_23190,N_23254);
or UO_402 (O_402,N_24551,N_24420);
xor UO_403 (O_403,N_24570,N_21270);
nand UO_404 (O_404,N_23076,N_24938);
xnor UO_405 (O_405,N_24822,N_23223);
xnor UO_406 (O_406,N_20517,N_23668);
nor UO_407 (O_407,N_22507,N_21459);
xor UO_408 (O_408,N_24029,N_24613);
nand UO_409 (O_409,N_23745,N_21268);
xnor UO_410 (O_410,N_24286,N_22322);
nor UO_411 (O_411,N_22594,N_24010);
nand UO_412 (O_412,N_24367,N_22257);
xnor UO_413 (O_413,N_22488,N_21360);
xnor UO_414 (O_414,N_22124,N_20245);
xor UO_415 (O_415,N_20521,N_24268);
xor UO_416 (O_416,N_20862,N_23717);
nand UO_417 (O_417,N_22462,N_24554);
or UO_418 (O_418,N_21939,N_20875);
xnor UO_419 (O_419,N_24618,N_21991);
nand UO_420 (O_420,N_24466,N_23299);
nand UO_421 (O_421,N_22908,N_23101);
or UO_422 (O_422,N_21263,N_23285);
or UO_423 (O_423,N_20795,N_20511);
nand UO_424 (O_424,N_21503,N_23425);
nor UO_425 (O_425,N_23068,N_21903);
nand UO_426 (O_426,N_21696,N_22291);
xor UO_427 (O_427,N_23056,N_21035);
or UO_428 (O_428,N_22601,N_24301);
or UO_429 (O_429,N_22955,N_23584);
xor UO_430 (O_430,N_24839,N_22373);
nand UO_431 (O_431,N_21113,N_23193);
nor UO_432 (O_432,N_21657,N_21743);
and UO_433 (O_433,N_24884,N_20847);
nand UO_434 (O_434,N_22150,N_20992);
nand UO_435 (O_435,N_24384,N_23877);
nor UO_436 (O_436,N_22211,N_23730);
nand UO_437 (O_437,N_21817,N_22317);
and UO_438 (O_438,N_23920,N_20086);
nand UO_439 (O_439,N_21777,N_20300);
or UO_440 (O_440,N_22636,N_24507);
xor UO_441 (O_441,N_23087,N_23393);
and UO_442 (O_442,N_22209,N_23478);
nand UO_443 (O_443,N_21020,N_23470);
nor UO_444 (O_444,N_20640,N_21722);
and UO_445 (O_445,N_20324,N_20974);
and UO_446 (O_446,N_23818,N_20843);
nor UO_447 (O_447,N_20317,N_24921);
xnor UO_448 (O_448,N_22051,N_23012);
nor UO_449 (O_449,N_23111,N_20923);
nor UO_450 (O_450,N_23119,N_22749);
nand UO_451 (O_451,N_23264,N_23224);
and UO_452 (O_452,N_21312,N_23701);
xnor UO_453 (O_453,N_23506,N_20023);
nand UO_454 (O_454,N_23489,N_21630);
and UO_455 (O_455,N_22832,N_22071);
nand UO_456 (O_456,N_20962,N_24060);
nor UO_457 (O_457,N_21443,N_22153);
or UO_458 (O_458,N_24863,N_20069);
xnor UO_459 (O_459,N_22425,N_21094);
xnor UO_460 (O_460,N_21910,N_20684);
xnor UO_461 (O_461,N_24468,N_21377);
nand UO_462 (O_462,N_22140,N_22623);
and UO_463 (O_463,N_24968,N_23916);
nand UO_464 (O_464,N_20471,N_22938);
xor UO_465 (O_465,N_23553,N_21102);
and UO_466 (O_466,N_20768,N_23669);
nor UO_467 (O_467,N_24123,N_21267);
or UO_468 (O_468,N_23339,N_23687);
xnor UO_469 (O_469,N_22129,N_21500);
nor UO_470 (O_470,N_21523,N_22682);
or UO_471 (O_471,N_23290,N_21230);
nand UO_472 (O_472,N_23574,N_24235);
xnor UO_473 (O_473,N_22525,N_23910);
and UO_474 (O_474,N_20248,N_21601);
and UO_475 (O_475,N_21179,N_22757);
and UO_476 (O_476,N_20603,N_24907);
or UO_477 (O_477,N_23978,N_24985);
or UO_478 (O_478,N_21468,N_20779);
or UO_479 (O_479,N_22381,N_22617);
or UO_480 (O_480,N_22813,N_22885);
xor UO_481 (O_481,N_22409,N_24434);
xnor UO_482 (O_482,N_20913,N_20757);
nand UO_483 (O_483,N_21934,N_22465);
nand UO_484 (O_484,N_21543,N_24642);
nand UO_485 (O_485,N_22958,N_21660);
and UO_486 (O_486,N_24175,N_20173);
and UO_487 (O_487,N_21401,N_23793);
and UO_488 (O_488,N_22745,N_22844);
nand UO_489 (O_489,N_24728,N_23538);
nand UO_490 (O_490,N_23633,N_20537);
or UO_491 (O_491,N_22827,N_20792);
and UO_492 (O_492,N_23416,N_23354);
or UO_493 (O_493,N_24283,N_22348);
nor UO_494 (O_494,N_22239,N_22277);
xor UO_495 (O_495,N_21661,N_21421);
xnor UO_496 (O_496,N_23423,N_24587);
nand UO_497 (O_497,N_23652,N_21966);
nor UO_498 (O_498,N_22913,N_22193);
nand UO_499 (O_499,N_23513,N_21514);
xnor UO_500 (O_500,N_21784,N_23180);
nand UO_501 (O_501,N_24324,N_23302);
nor UO_502 (O_502,N_21989,N_21639);
nand UO_503 (O_503,N_24876,N_23155);
nand UO_504 (O_504,N_24019,N_20383);
nor UO_505 (O_505,N_24241,N_21477);
nand UO_506 (O_506,N_21162,N_20971);
nor UO_507 (O_507,N_20504,N_22000);
nor UO_508 (O_508,N_24050,N_20869);
and UO_509 (O_509,N_20098,N_20124);
and UO_510 (O_510,N_20704,N_23646);
nor UO_511 (O_511,N_20667,N_20683);
or UO_512 (O_512,N_21284,N_24105);
xor UO_513 (O_513,N_21038,N_20341);
nor UO_514 (O_514,N_20737,N_22042);
nand UO_515 (O_515,N_23039,N_21154);
or UO_516 (O_516,N_22809,N_21859);
xor UO_517 (O_517,N_21554,N_22741);
and UO_518 (O_518,N_22353,N_20253);
or UO_519 (O_519,N_20252,N_22249);
nand UO_520 (O_520,N_20131,N_20585);
and UO_521 (O_521,N_21866,N_24664);
and UO_522 (O_522,N_24512,N_22910);
nand UO_523 (O_523,N_24632,N_23041);
xnor UO_524 (O_524,N_22940,N_21979);
nor UO_525 (O_525,N_23939,N_23286);
or UO_526 (O_526,N_24976,N_22968);
xor UO_527 (O_527,N_21987,N_20947);
nor UO_528 (O_528,N_20348,N_21317);
xor UO_529 (O_529,N_22128,N_23990);
or UO_530 (O_530,N_22142,N_21353);
and UO_531 (O_531,N_22194,N_21761);
nand UO_532 (O_532,N_23370,N_23692);
or UO_533 (O_533,N_22652,N_24228);
nand UO_534 (O_534,N_22996,N_20677);
and UO_535 (O_535,N_22963,N_20154);
and UO_536 (O_536,N_23508,N_21652);
nor UO_537 (O_537,N_23367,N_21881);
nand UO_538 (O_538,N_22175,N_24142);
or UO_539 (O_539,N_23079,N_21088);
nand UO_540 (O_540,N_24704,N_23305);
nor UO_541 (O_541,N_24209,N_23315);
or UO_542 (O_542,N_22663,N_22686);
and UO_543 (O_543,N_24891,N_20595);
and UO_544 (O_544,N_20633,N_22609);
nand UO_545 (O_545,N_20167,N_24859);
and UO_546 (O_546,N_24498,N_20624);
and UO_547 (O_547,N_20790,N_20197);
or UO_548 (O_548,N_20448,N_22549);
xor UO_549 (O_549,N_20359,N_24961);
xor UO_550 (O_550,N_24924,N_23997);
xnor UO_551 (O_551,N_22751,N_21805);
nor UO_552 (O_552,N_23494,N_21164);
xor UO_553 (O_553,N_20249,N_20436);
and UO_554 (O_554,N_21239,N_21436);
xor UO_555 (O_555,N_22032,N_24821);
nor UO_556 (O_556,N_24505,N_21865);
nor UO_557 (O_557,N_21613,N_21801);
or UO_558 (O_558,N_24970,N_20687);
xnor UO_559 (O_559,N_22606,N_24173);
and UO_560 (O_560,N_24092,N_22394);
and UO_561 (O_561,N_22155,N_21953);
and UO_562 (O_562,N_20698,N_21766);
nor UO_563 (O_563,N_22271,N_21203);
xnor UO_564 (O_564,N_24234,N_23078);
and UO_565 (O_565,N_23892,N_22207);
and UO_566 (O_566,N_22123,N_21456);
nand UO_567 (O_567,N_24879,N_24718);
nand UO_568 (O_568,N_22111,N_21029);
or UO_569 (O_569,N_23869,N_23632);
xor UO_570 (O_570,N_22675,N_22078);
and UO_571 (O_571,N_23665,N_22596);
and UO_572 (O_572,N_21332,N_23879);
nor UO_573 (O_573,N_23683,N_21434);
or UO_574 (O_574,N_22948,N_23794);
or UO_575 (O_575,N_21845,N_24084);
xor UO_576 (O_576,N_22264,N_23492);
or UO_577 (O_577,N_22625,N_21213);
or UO_578 (O_578,N_22746,N_22559);
or UO_579 (O_579,N_20087,N_24320);
or UO_580 (O_580,N_21010,N_21524);
xor UO_581 (O_581,N_21367,N_23977);
and UO_582 (O_582,N_21392,N_23772);
nor UO_583 (O_583,N_23798,N_20668);
or UO_584 (O_584,N_21135,N_21864);
or UO_585 (O_585,N_21342,N_20474);
or UO_586 (O_586,N_24868,N_20549);
nor UO_587 (O_587,N_23969,N_21960);
nor UO_588 (O_588,N_22138,N_24841);
nand UO_589 (O_589,N_23966,N_20156);
xor UO_590 (O_590,N_22918,N_22398);
or UO_591 (O_591,N_24933,N_20567);
nand UO_592 (O_592,N_20005,N_23570);
or UO_593 (O_593,N_21926,N_20291);
and UO_594 (O_594,N_20010,N_22545);
xnor UO_595 (O_595,N_24980,N_24866);
or UO_596 (O_596,N_22120,N_22562);
and UO_597 (O_597,N_21963,N_20438);
and UO_598 (O_598,N_24318,N_22404);
nand UO_599 (O_599,N_22983,N_24179);
or UO_600 (O_600,N_21951,N_22376);
or UO_601 (O_601,N_22299,N_22360);
nand UO_602 (O_602,N_22765,N_24944);
nor UO_603 (O_603,N_22356,N_23171);
nor UO_604 (O_604,N_20849,N_20544);
xnor UO_605 (O_605,N_24066,N_20797);
xnor UO_606 (O_606,N_24890,N_22950);
nand UO_607 (O_607,N_21052,N_24031);
nand UO_608 (O_608,N_24364,N_22546);
nor UO_609 (O_609,N_20600,N_20518);
nor UO_610 (O_610,N_22436,N_20914);
and UO_611 (O_611,N_23353,N_21944);
and UO_612 (O_612,N_22370,N_21912);
and UO_613 (O_613,N_21001,N_22166);
and UO_614 (O_614,N_23599,N_23783);
xor UO_615 (O_615,N_21282,N_22868);
and UO_616 (O_616,N_21604,N_21563);
or UO_617 (O_617,N_21704,N_24380);
and UO_618 (O_618,N_21861,N_22937);
nor UO_619 (O_619,N_22490,N_20278);
or UO_620 (O_620,N_20616,N_22339);
nand UO_621 (O_621,N_22076,N_20818);
nor UO_622 (O_622,N_23568,N_21228);
or UO_623 (O_623,N_21731,N_23098);
and UO_624 (O_624,N_23819,N_20454);
xnor UO_625 (O_625,N_21727,N_20215);
nand UO_626 (O_626,N_24572,N_23113);
or UO_627 (O_627,N_22015,N_24395);
nor UO_628 (O_628,N_23803,N_23814);
or UO_629 (O_629,N_23210,N_23924);
nor UO_630 (O_630,N_24280,N_21588);
or UO_631 (O_631,N_24547,N_23888);
or UO_632 (O_632,N_23320,N_20316);
xor UO_633 (O_633,N_20815,N_24067);
xor UO_634 (O_634,N_23121,N_23204);
nor UO_635 (O_635,N_23762,N_23544);
or UO_636 (O_636,N_22970,N_21648);
nand UO_637 (O_637,N_21533,N_22561);
xor UO_638 (O_638,N_21211,N_22990);
or UO_639 (O_639,N_23417,N_20783);
and UO_640 (O_640,N_21126,N_20964);
xnor UO_641 (O_641,N_20691,N_20479);
or UO_642 (O_642,N_22413,N_24079);
nor UO_643 (O_643,N_22456,N_21089);
or UO_644 (O_644,N_21030,N_22660);
nand UO_645 (O_645,N_22014,N_24981);
and UO_646 (O_646,N_23409,N_20982);
nor UO_647 (O_647,N_22349,N_20570);
nand UO_648 (O_648,N_23639,N_22466);
xnor UO_649 (O_649,N_24966,N_22453);
or UO_650 (O_650,N_24612,N_20880);
nor UO_651 (O_651,N_23583,N_20384);
nor UO_652 (O_652,N_22423,N_20866);
nand UO_653 (O_653,N_23509,N_22106);
or UO_654 (O_654,N_23757,N_21433);
nor UO_655 (O_655,N_23293,N_23003);
or UO_656 (O_656,N_22945,N_23440);
or UO_657 (O_657,N_20998,N_20546);
nand UO_658 (O_658,N_20493,N_22365);
xnor UO_659 (O_659,N_21196,N_22202);
and UO_660 (O_660,N_24694,N_22728);
xor UO_661 (O_661,N_20225,N_23702);
or UO_662 (O_662,N_24651,N_21946);
nor UO_663 (O_663,N_23933,N_20220);
nand UO_664 (O_664,N_23871,N_24799);
nor UO_665 (O_665,N_21075,N_22061);
or UO_666 (O_666,N_21890,N_24781);
xor UO_667 (O_667,N_22009,N_24405);
nor UO_668 (O_668,N_23769,N_21681);
nand UO_669 (O_669,N_24951,N_24408);
or UO_670 (O_670,N_20495,N_21679);
or UO_671 (O_671,N_23659,N_20613);
xor UO_672 (O_672,N_22272,N_20505);
or UO_673 (O_673,N_21916,N_20500);
nand UO_674 (O_674,N_24926,N_22294);
nor UO_675 (O_675,N_24140,N_20413);
and UO_676 (O_676,N_22873,N_21068);
or UO_677 (O_677,N_23981,N_21227);
nor UO_678 (O_678,N_21632,N_20257);
nand UO_679 (O_679,N_24265,N_24670);
and UO_680 (O_680,N_20209,N_24566);
and UO_681 (O_681,N_21993,N_20194);
nand UO_682 (O_682,N_23605,N_22470);
nand UO_683 (O_683,N_20444,N_20740);
or UO_684 (O_684,N_24444,N_24045);
nor UO_685 (O_685,N_22597,N_21629);
and UO_686 (O_686,N_21180,N_23992);
or UO_687 (O_687,N_24245,N_20629);
and UO_688 (O_688,N_24487,N_21915);
and UO_689 (O_689,N_22234,N_21793);
and UO_690 (O_690,N_22502,N_24770);
nor UO_691 (O_691,N_24037,N_20256);
xnor UO_692 (O_692,N_23324,N_21464);
nand UO_693 (O_693,N_24901,N_21358);
nor UO_694 (O_694,N_23520,N_24171);
nand UO_695 (O_695,N_22049,N_23634);
nand UO_696 (O_696,N_22719,N_23382);
or UO_697 (O_697,N_22007,N_24436);
nor UO_698 (O_698,N_20721,N_20620);
and UO_699 (O_699,N_23212,N_24561);
nand UO_700 (O_700,N_20569,N_20077);
nand UO_701 (O_701,N_22389,N_23971);
or UO_702 (O_702,N_23132,N_21252);
nor UO_703 (O_703,N_23278,N_24023);
or UO_704 (O_704,N_24972,N_24149);
nor UO_705 (O_705,N_21370,N_22646);
nand UO_706 (O_706,N_23631,N_23962);
and UO_707 (O_707,N_24109,N_20049);
nor UO_708 (O_708,N_22856,N_22733);
and UO_709 (O_709,N_21947,N_20360);
xnor UO_710 (O_710,N_23936,N_20799);
or UO_711 (O_711,N_20496,N_24250);
nor UO_712 (O_712,N_24223,N_24363);
nand UO_713 (O_713,N_23771,N_21427);
xnor UO_714 (O_714,N_23711,N_21614);
nor UO_715 (O_715,N_22839,N_22085);
xor UO_716 (O_716,N_24645,N_23360);
or UO_717 (O_717,N_22080,N_24785);
nand UO_718 (O_718,N_22432,N_20224);
and UO_719 (O_719,N_21578,N_22186);
or UO_720 (O_720,N_24874,N_21318);
and UO_721 (O_721,N_23531,N_24975);
or UO_722 (O_722,N_22028,N_21232);
nand UO_723 (O_723,N_22222,N_24575);
nand UO_724 (O_724,N_22351,N_24631);
xnor UO_725 (O_725,N_21787,N_21687);
or UO_726 (O_726,N_22223,N_23112);
or UO_727 (O_727,N_24218,N_21256);
nand UO_728 (O_728,N_20394,N_22312);
xnor UO_729 (O_729,N_24550,N_20039);
xor UO_730 (O_730,N_22555,N_23053);
and UO_731 (O_731,N_23064,N_22400);
nand UO_732 (O_732,N_21432,N_24017);
xor UO_733 (O_733,N_22164,N_21750);
nor UO_734 (O_734,N_23995,N_23430);
nor UO_735 (O_735,N_21062,N_23475);
nand UO_736 (O_736,N_20672,N_20308);
xor UO_737 (O_737,N_23082,N_24057);
nor UO_738 (O_738,N_23729,N_22366);
nand UO_739 (O_739,N_20742,N_23691);
nor UO_740 (O_740,N_23724,N_23485);
and UO_741 (O_741,N_23638,N_24886);
and UO_742 (O_742,N_23124,N_21774);
nor UO_743 (O_743,N_22133,N_20845);
nand UO_744 (O_744,N_20636,N_22151);
and UO_745 (O_745,N_24300,N_21346);
and UO_746 (O_746,N_23363,N_24307);
nand UO_747 (O_747,N_22709,N_21422);
xnor UO_748 (O_748,N_24158,N_24931);
nor UO_749 (O_749,N_22911,N_22438);
or UO_750 (O_750,N_20959,N_24708);
and UO_751 (O_751,N_23767,N_22524);
nor UO_752 (O_752,N_20881,N_24478);
and UO_753 (O_753,N_23156,N_24333);
and UO_754 (O_754,N_24707,N_21643);
or UO_755 (O_755,N_20695,N_20475);
and UO_756 (O_756,N_24805,N_22281);
or UO_757 (O_757,N_20455,N_22768);
nor UO_758 (O_758,N_21788,N_24622);
or UO_759 (O_759,N_22482,N_20472);
nor UO_760 (O_760,N_24827,N_24201);
xnor UO_761 (O_761,N_20842,N_20812);
xnor UO_762 (O_762,N_20986,N_23428);
nand UO_763 (O_763,N_23941,N_24696);
and UO_764 (O_764,N_20593,N_20217);
xnor UO_765 (O_765,N_22995,N_23058);
or UO_766 (O_766,N_24847,N_23942);
nor UO_767 (O_767,N_23203,N_20013);
nor UO_768 (O_768,N_21786,N_23395);
nor UO_769 (O_769,N_23529,N_21586);
nand UO_770 (O_770,N_23833,N_22980);
and UO_771 (O_771,N_21557,N_22861);
or UO_772 (O_772,N_22588,N_24720);
and UO_773 (O_773,N_21302,N_20423);
and UO_774 (O_774,N_22516,N_21606);
xnor UO_775 (O_775,N_20829,N_21356);
and UO_776 (O_776,N_24012,N_20661);
nand UO_777 (O_777,N_22897,N_20223);
xor UO_778 (O_778,N_22680,N_22998);
nand UO_779 (O_779,N_20270,N_24340);
nor UO_780 (O_780,N_24022,N_24615);
nand UO_781 (O_781,N_21151,N_21262);
nand UO_782 (O_782,N_22821,N_23947);
xor UO_783 (O_783,N_22605,N_22627);
nor UO_784 (O_784,N_24205,N_21701);
and UO_785 (O_785,N_24935,N_21511);
nor UO_786 (O_786,N_23490,N_23709);
xor UO_787 (O_787,N_24270,N_23105);
nand UO_788 (O_788,N_21852,N_23256);
xor UO_789 (O_789,N_22122,N_23261);
or UO_790 (O_790,N_22774,N_21307);
nand UO_791 (O_791,N_22891,N_22667);
or UO_792 (O_792,N_20646,N_22097);
nand UO_793 (O_793,N_22730,N_22233);
nand UO_794 (O_794,N_20235,N_21402);
xnor UO_795 (O_795,N_24527,N_22531);
nor UO_796 (O_796,N_23332,N_24746);
or UO_797 (O_797,N_23228,N_24883);
nor UO_798 (O_798,N_20157,N_23782);
nand UO_799 (O_799,N_23993,N_20844);
and UO_800 (O_800,N_21831,N_20765);
xnor UO_801 (O_801,N_23257,N_24294);
and UO_802 (O_802,N_21215,N_24137);
xor UO_803 (O_803,N_22884,N_23598);
and UO_804 (O_804,N_22093,N_23827);
nand UO_805 (O_805,N_21471,N_21494);
nor UO_806 (O_806,N_20568,N_21508);
xnor UO_807 (O_807,N_24862,N_24357);
nor UO_808 (O_808,N_21830,N_24602);
nand UO_809 (O_809,N_24758,N_21040);
nand UO_810 (O_810,N_24193,N_20564);
xor UO_811 (O_811,N_20666,N_22854);
and UO_812 (O_812,N_21977,N_22375);
xor UO_813 (O_813,N_23151,N_21069);
xor UO_814 (O_814,N_21019,N_24456);
nand UO_815 (O_815,N_23384,N_23188);
xnor UO_816 (O_816,N_24760,N_22929);
and UO_817 (O_817,N_24134,N_23473);
and UO_818 (O_818,N_24623,N_23987);
and UO_819 (O_819,N_24197,N_23891);
nand UO_820 (O_820,N_22476,N_20915);
or UO_821 (O_821,N_21579,N_23005);
nand UO_822 (O_822,N_24672,N_20714);
and UO_823 (O_823,N_21271,N_20969);
xnor UO_824 (O_824,N_21721,N_22100);
or UO_825 (O_825,N_24503,N_23760);
xnor UO_826 (O_826,N_24312,N_20837);
xor UO_827 (O_827,N_23253,N_22962);
nand UO_828 (O_828,N_24850,N_22685);
nor UO_829 (O_829,N_21911,N_20042);
xnor UO_830 (O_830,N_22232,N_24220);
or UO_831 (O_831,N_22176,N_21921);
or UO_832 (O_832,N_20467,N_23986);
or UO_833 (O_833,N_20851,N_21775);
xor UO_834 (O_834,N_22333,N_24603);
or UO_835 (O_835,N_21812,N_22437);
or UO_836 (O_836,N_20638,N_24150);
or UO_837 (O_837,N_21057,N_22084);
nor UO_838 (O_838,N_20838,N_22750);
xnor UO_839 (O_839,N_23573,N_23388);
nor UO_840 (O_840,N_20462,N_20078);
nand UO_841 (O_841,N_24077,N_22416);
nor UO_842 (O_842,N_24107,N_21084);
nand UO_843 (O_843,N_24888,N_20800);
xor UO_844 (O_844,N_20598,N_22337);
and UO_845 (O_845,N_21566,N_22287);
or UO_846 (O_846,N_23067,N_21197);
nand UO_847 (O_847,N_24379,N_21789);
nand UO_848 (O_848,N_20354,N_21869);
xnor UO_849 (O_849,N_22583,N_24571);
nor UO_850 (O_850,N_24194,N_21502);
nor UO_851 (O_851,N_24577,N_21927);
and UO_852 (O_852,N_23569,N_21254);
xnor UO_853 (O_853,N_20070,N_24656);
xor UO_854 (O_854,N_21028,N_24287);
or UO_855 (O_855,N_23394,N_23714);
nand UO_856 (O_856,N_24904,N_21177);
or UO_857 (O_857,N_23690,N_22865);
nor UO_858 (O_858,N_22201,N_22379);
nand UO_859 (O_859,N_20114,N_24141);
xor UO_860 (O_860,N_22273,N_23427);
nor UO_861 (O_861,N_22961,N_22089);
nand UO_862 (O_862,N_24659,N_20411);
nor UO_863 (O_863,N_23017,N_24591);
nand UO_864 (O_864,N_23899,N_22815);
and UO_865 (O_865,N_21420,N_22701);
nor UO_866 (O_866,N_22681,N_22444);
and UO_867 (O_867,N_20560,N_20238);
nor UO_868 (O_868,N_22221,N_24143);
nand UO_869 (O_869,N_22378,N_21063);
and UO_870 (O_870,N_23013,N_23400);
nand UO_871 (O_871,N_20226,N_21627);
or UO_872 (O_872,N_20076,N_20834);
and UO_873 (O_873,N_20043,N_24450);
nand UO_874 (O_874,N_22881,N_20489);
and UO_875 (O_875,N_23272,N_22552);
xor UO_876 (O_876,N_22710,N_21546);
and UO_877 (O_877,N_22760,N_24680);
nand UO_878 (O_878,N_20685,N_20378);
nor UO_879 (O_879,N_23934,N_24180);
nor UO_880 (O_880,N_23935,N_22110);
and UO_881 (O_881,N_22798,N_22056);
or UO_882 (O_882,N_24041,N_24590);
and UO_883 (O_883,N_24230,N_23880);
nor UO_884 (O_884,N_22571,N_23567);
and UO_885 (O_885,N_20557,N_20920);
nand UO_886 (O_886,N_22618,N_22887);
nand UO_887 (O_887,N_21732,N_22989);
xor UO_888 (O_888,N_24765,N_20934);
and UO_889 (O_889,N_23656,N_24226);
nor UO_890 (O_890,N_22661,N_22219);
or UO_891 (O_891,N_24717,N_21012);
xor UO_892 (O_892,N_20972,N_20189);
and UO_893 (O_893,N_23329,N_22973);
nor UO_894 (O_894,N_23779,N_24824);
or UO_895 (O_895,N_20282,N_24071);
nand UO_896 (O_896,N_24620,N_23964);
or UO_897 (O_897,N_22185,N_20752);
or UO_898 (O_898,N_20416,N_23943);
nor UO_899 (O_899,N_21534,N_20794);
nand UO_900 (O_900,N_23326,N_23883);
nand UO_901 (O_901,N_23383,N_23229);
nor UO_902 (O_902,N_23735,N_24833);
or UO_903 (O_903,N_20707,N_23551);
and UO_904 (O_904,N_24678,N_24043);
nor UO_905 (O_905,N_20127,N_21815);
nor UO_906 (O_906,N_24377,N_23999);
nand UO_907 (O_907,N_21110,N_23580);
xor UO_908 (O_908,N_24440,N_22560);
xnor UO_909 (O_909,N_21412,N_23624);
nor UO_910 (O_910,N_23115,N_23703);
and UO_911 (O_911,N_20989,N_20404);
nor UO_912 (O_912,N_22174,N_22065);
xnor UO_913 (O_913,N_22535,N_23063);
nor UO_914 (O_914,N_21335,N_21584);
and UO_915 (O_915,N_24872,N_24055);
nand UO_916 (O_916,N_23093,N_20895);
and UO_917 (O_917,N_20793,N_21055);
xor UO_918 (O_918,N_24545,N_24568);
nor UO_919 (O_919,N_22158,N_20981);
nor UO_920 (O_920,N_20103,N_22006);
and UO_921 (O_921,N_20619,N_23609);
nand UO_922 (O_922,N_24222,N_22782);
and UO_923 (O_923,N_23419,N_22247);
xor UO_924 (O_924,N_22241,N_20726);
or UO_925 (O_925,N_20700,N_21314);
and UO_926 (O_926,N_22244,N_24941);
nor UO_927 (O_927,N_24767,N_24074);
or UO_928 (O_928,N_21829,N_22591);
nand UO_929 (O_929,N_21051,N_24703);
or UO_930 (O_930,N_21118,N_22298);
xor UO_931 (O_931,N_22332,N_21495);
nor UO_932 (O_932,N_20513,N_20990);
nor UO_933 (O_933,N_24646,N_23022);
xnor UO_934 (O_934,N_21306,N_20681);
and UO_935 (O_935,N_23726,N_24643);
or UO_936 (O_936,N_22414,N_24701);
and UO_937 (O_937,N_20417,N_21160);
or UO_938 (O_938,N_24394,N_24929);
nor UO_939 (O_939,N_22764,N_21877);
and UO_940 (O_940,N_23671,N_22650);
or UO_941 (O_941,N_23303,N_23843);
or UO_942 (O_942,N_24754,N_20525);
or UO_943 (O_943,N_22900,N_24967);
xor UO_944 (O_944,N_22484,N_23795);
nor UO_945 (O_945,N_21549,N_21120);
nor UO_946 (O_946,N_22313,N_22814);
nand UO_947 (O_947,N_21615,N_20026);
or UO_948 (O_948,N_22324,N_20601);
or UO_949 (O_949,N_21127,N_23088);
xnor UO_950 (O_950,N_24963,N_20893);
and UO_951 (O_951,N_23523,N_20811);
or UO_952 (O_952,N_22347,N_21517);
nor UO_953 (O_953,N_23239,N_21770);
nor UO_954 (O_954,N_23898,N_20426);
and UO_955 (O_955,N_22520,N_23081);
nor UO_956 (O_956,N_20271,N_22780);
nand UO_957 (O_957,N_20349,N_23799);
nand UO_958 (O_958,N_21962,N_21080);
or UO_959 (O_959,N_20647,N_21175);
or UO_960 (O_960,N_22645,N_21833);
and UO_961 (O_961,N_20109,N_22518);
nand UO_962 (O_962,N_20524,N_24647);
nand UO_963 (O_963,N_22753,N_24665);
nor UO_964 (O_964,N_20212,N_21608);
and UO_965 (O_965,N_20244,N_22090);
xnor UO_966 (O_966,N_20606,N_23868);
and UO_967 (O_967,N_21981,N_23448);
nand UO_968 (O_968,N_21354,N_23009);
or UO_969 (O_969,N_23141,N_22863);
nor UO_970 (O_970,N_20002,N_24855);
or UO_971 (O_971,N_20536,N_20083);
xnor UO_972 (O_972,N_24851,N_22058);
nand UO_973 (O_973,N_20776,N_24003);
xor UO_974 (O_974,N_24288,N_22848);
or UO_975 (O_975,N_24836,N_24741);
nor UO_976 (O_976,N_21237,N_21857);
and UO_977 (O_977,N_24914,N_21497);
xnor UO_978 (O_978,N_23084,N_23062);
nand UO_979 (O_979,N_20503,N_23103);
nor UO_980 (O_980,N_24893,N_21577);
nor UO_981 (O_981,N_20024,N_23677);
nor UO_982 (O_982,N_22407,N_21286);
or UO_983 (O_983,N_23844,N_22830);
or UO_984 (O_984,N_22101,N_22578);
or UO_985 (O_985,N_22619,N_21913);
xnor UO_986 (O_986,N_22427,N_24609);
xnor UO_987 (O_987,N_20148,N_24675);
nand UO_988 (O_988,N_23853,N_24310);
nand UO_989 (O_989,N_23358,N_20694);
nand UO_990 (O_990,N_24779,N_24557);
nor UO_991 (O_991,N_22766,N_24489);
nand UO_992 (O_992,N_24263,N_23486);
nor UO_993 (O_993,N_24190,N_21357);
and UO_994 (O_994,N_24560,N_20125);
xnor UO_995 (O_995,N_23560,N_22371);
nor UO_996 (O_996,N_24062,N_24558);
or UO_997 (O_997,N_24744,N_22452);
and UO_998 (O_998,N_20771,N_23460);
or UO_999 (O_999,N_21304,N_20555);
nand UO_1000 (O_1000,N_24588,N_21116);
or UO_1001 (O_1001,N_24125,N_22835);
nand UO_1002 (O_1002,N_20118,N_21037);
or UO_1003 (O_1003,N_20690,N_22883);
xor UO_1004 (O_1004,N_21905,N_22586);
xor UO_1005 (O_1005,N_21535,N_24521);
xnor UO_1006 (O_1006,N_23679,N_21709);
or UO_1007 (O_1007,N_24937,N_21756);
or UO_1008 (O_1008,N_23083,N_22492);
nor UO_1009 (O_1009,N_20274,N_20165);
or UO_1010 (O_1010,N_21712,N_24327);
or UO_1011 (O_1011,N_22878,N_24328);
and UO_1012 (O_1012,N_21301,N_23161);
xor UO_1013 (O_1013,N_21530,N_24997);
xnor UO_1014 (O_1014,N_22505,N_21341);
nor UO_1015 (O_1015,N_24903,N_24290);
nor UO_1016 (O_1016,N_23280,N_21757);
nor UO_1017 (O_1017,N_20123,N_22403);
nand UO_1018 (O_1018,N_20786,N_20449);
nor UO_1019 (O_1019,N_23157,N_22696);
or UO_1020 (O_1020,N_22697,N_24135);
nand UO_1021 (O_1021,N_22668,N_21425);
nor UO_1022 (O_1022,N_24662,N_20032);
nor UO_1023 (O_1023,N_21108,N_24485);
nand UO_1024 (O_1024,N_21034,N_23697);
nor UO_1025 (O_1025,N_20102,N_24154);
xnor UO_1026 (O_1026,N_23232,N_20466);
nand UO_1027 (O_1027,N_21717,N_23676);
nor UO_1028 (O_1028,N_23344,N_24139);
nor UO_1029 (O_1029,N_21698,N_20980);
or UO_1030 (O_1030,N_24537,N_20093);
xnor UO_1031 (O_1031,N_22369,N_24418);
xor UO_1032 (O_1032,N_24787,N_24266);
and UO_1033 (O_1033,N_23389,N_20730);
nand UO_1034 (O_1034,N_24042,N_23810);
nor UO_1035 (O_1035,N_24690,N_24202);
xor UO_1036 (O_1036,N_24882,N_22576);
nand UO_1037 (O_1037,N_20791,N_22550);
nor UO_1038 (O_1038,N_22198,N_24196);
xor UO_1039 (O_1039,N_24593,N_21452);
or UO_1040 (O_1040,N_21725,N_21220);
nand UO_1041 (O_1041,N_20222,N_22380);
or UO_1042 (O_1042,N_23589,N_20246);
nor UO_1043 (O_1043,N_22424,N_24936);
nand UO_1044 (O_1044,N_20509,N_24555);
or UO_1045 (O_1045,N_24687,N_22912);
and UO_1046 (O_1046,N_20671,N_22485);
nand UO_1047 (O_1047,N_23615,N_24619);
and UO_1048 (O_1048,N_23740,N_23094);
nand UO_1049 (O_1049,N_24838,N_24517);
and UO_1050 (O_1050,N_22984,N_21011);
nor UO_1051 (O_1051,N_20122,N_23148);
nand UO_1052 (O_1052,N_22992,N_23104);
nor UO_1053 (O_1053,N_22446,N_22368);
and UO_1054 (O_1054,N_24826,N_21131);
nand UO_1055 (O_1055,N_22771,N_21414);
xnor UO_1056 (O_1056,N_23955,N_20898);
and UO_1057 (O_1057,N_23585,N_24626);
and UO_1058 (O_1058,N_23107,N_22108);
nand UO_1059 (O_1059,N_23781,N_22634);
or UO_1060 (O_1060,N_20868,N_22633);
xnor UO_1061 (O_1061,N_22991,N_22341);
nor UO_1062 (O_1062,N_24178,N_21668);
xnor UO_1063 (O_1063,N_22288,N_24815);
nor UO_1064 (O_1064,N_24314,N_20437);
or UO_1065 (O_1065,N_24455,N_22095);
nor UO_1066 (O_1066,N_20723,N_24712);
and UO_1067 (O_1067,N_20337,N_24596);
xor UO_1068 (O_1068,N_24573,N_23192);
and UO_1069 (O_1069,N_24677,N_21167);
nand UO_1070 (O_1070,N_23613,N_23364);
xnor UO_1071 (O_1071,N_21841,N_21074);
nand UO_1072 (O_1072,N_20054,N_21091);
or UO_1073 (O_1073,N_23823,N_24982);
nand UO_1074 (O_1074,N_23784,N_21995);
nand UO_1075 (O_1075,N_23864,N_20916);
and UO_1076 (O_1076,N_23972,N_20347);
or UO_1077 (O_1077,N_24491,N_23950);
nor UO_1078 (O_1078,N_21548,N_23225);
and UO_1079 (O_1079,N_20941,N_22307);
xor UO_1080 (O_1080,N_23713,N_23991);
nand UO_1081 (O_1081,N_21275,N_21223);
xnor UO_1082 (O_1082,N_22977,N_24993);
nand UO_1083 (O_1083,N_20216,N_22117);
or UO_1084 (O_1084,N_22428,N_20738);
or UO_1085 (O_1085,N_22915,N_20089);
xor UO_1086 (O_1086,N_24354,N_21688);
and UO_1087 (O_1087,N_21945,N_21693);
nor UO_1088 (O_1088,N_23237,N_20954);
xnor UO_1089 (O_1089,N_20051,N_21547);
xnor UO_1090 (O_1090,N_23054,N_24889);
nand UO_1091 (O_1091,N_21892,N_20674);
nor UO_1092 (O_1092,N_20905,N_20044);
or UO_1093 (O_1093,N_24809,N_24088);
xor UO_1094 (O_1094,N_22731,N_24954);
nand UO_1095 (O_1095,N_23802,N_23457);
or UO_1096 (O_1096,N_21929,N_22526);
xnor UO_1097 (O_1097,N_21986,N_21907);
and UO_1098 (O_1098,N_20314,N_23424);
xnor UO_1099 (O_1099,N_21532,N_23209);
xor UO_1100 (O_1100,N_23045,N_23092);
nand UO_1101 (O_1101,N_20407,N_21467);
and UO_1102 (O_1102,N_21938,N_21922);
nand UO_1103 (O_1103,N_21199,N_21891);
nand UO_1104 (O_1104,N_21612,N_23922);
nand UO_1105 (O_1105,N_21515,N_22769);
nand UO_1106 (O_1106,N_24606,N_20459);
nor UO_1107 (O_1107,N_21902,N_24569);
nor UO_1108 (O_1108,N_20867,N_23476);
and UO_1109 (O_1109,N_24927,N_22494);
or UO_1110 (O_1110,N_24794,N_21348);
xnor UO_1111 (O_1111,N_22939,N_24281);
xor UO_1112 (O_1112,N_20930,N_20170);
and UO_1113 (O_1113,N_22450,N_24033);
and UO_1114 (O_1114,N_20497,N_21803);
xor UO_1115 (O_1115,N_24705,N_22957);
and UO_1116 (O_1116,N_22017,N_20739);
and UO_1117 (O_1117,N_21872,N_21413);
or UO_1118 (O_1118,N_22486,N_21488);
and UO_1119 (O_1119,N_22744,N_24969);
nand UO_1120 (O_1120,N_24742,N_24438);
or UO_1121 (O_1121,N_23330,N_21236);
nand UO_1122 (O_1122,N_21763,N_24255);
nand UO_1123 (O_1123,N_21611,N_23131);
nand UO_1124 (O_1124,N_20395,N_23805);
or UO_1125 (O_1125,N_23241,N_23090);
or UO_1126 (O_1126,N_24912,N_22952);
and UO_1127 (O_1127,N_20534,N_24035);
or UO_1128 (O_1128,N_23841,N_22027);
nand UO_1129 (O_1129,N_23759,N_24484);
and UO_1130 (O_1130,N_23696,N_20259);
nand UO_1131 (O_1131,N_21809,N_20020);
nand UO_1132 (O_1132,N_21676,N_22355);
and UO_1133 (O_1133,N_24157,N_22119);
nand UO_1134 (O_1134,N_20152,N_23857);
xnor UO_1135 (O_1135,N_20377,N_22642);
nor UO_1136 (O_1136,N_22031,N_24995);
or UO_1137 (O_1137,N_22801,N_21894);
nand UO_1138 (O_1138,N_23026,N_22556);
nor UO_1139 (O_1139,N_24624,N_20046);
xnor UO_1140 (O_1140,N_24415,N_22044);
or UO_1141 (O_1141,N_20526,N_20186);
nand UO_1142 (O_1142,N_22002,N_24402);
or UO_1143 (O_1143,N_20397,N_23325);
nand UO_1144 (O_1144,N_21708,N_24714);
xnor UO_1145 (O_1145,N_24834,N_23199);
or UO_1146 (O_1146,N_24164,N_24239);
nand UO_1147 (O_1147,N_21751,N_20071);
and UO_1148 (O_1148,N_20320,N_24089);
and UO_1149 (O_1149,N_20822,N_24349);
xor UO_1150 (O_1150,N_21047,N_24168);
and UO_1151 (O_1151,N_20732,N_20865);
nand UO_1152 (O_1152,N_21333,N_21124);
nor UO_1153 (O_1153,N_21054,N_24534);
nor UO_1154 (O_1154,N_20379,N_20268);
xnor UO_1155 (O_1155,N_20858,N_24014);
or UO_1156 (O_1156,N_23511,N_23909);
nand UO_1157 (O_1157,N_20510,N_20571);
xor UO_1158 (O_1158,N_21305,N_24054);
or UO_1159 (O_1159,N_21664,N_24413);
or UO_1160 (O_1160,N_24258,N_22901);
and UO_1161 (O_1161,N_21746,N_23878);
xnor UO_1162 (O_1162,N_23721,N_22738);
or UO_1163 (O_1163,N_21486,N_20388);
and UO_1164 (O_1164,N_20558,N_22300);
or UO_1165 (O_1165,N_20693,N_20266);
xnor UO_1166 (O_1166,N_24481,N_23333);
nor UO_1167 (O_1167,N_21832,N_23848);
or UO_1168 (O_1168,N_21737,N_21172);
or UO_1169 (O_1169,N_24437,N_22074);
xnor UO_1170 (O_1170,N_20239,N_22474);
xnor UO_1171 (O_1171,N_23514,N_21598);
and UO_1172 (O_1172,N_20530,N_23901);
or UO_1173 (O_1173,N_23973,N_20665);
nor UO_1174 (O_1174,N_23042,N_21545);
xor UO_1175 (O_1175,N_23715,N_21352);
nor UO_1176 (O_1176,N_20477,N_23255);
and UO_1177 (O_1177,N_21600,N_22121);
nand UO_1178 (O_1178,N_24715,N_20402);
nor UO_1179 (O_1179,N_24389,N_22572);
or UO_1180 (O_1180,N_21496,N_20956);
and UO_1181 (O_1181,N_20334,N_23136);
xnor UO_1182 (O_1182,N_24525,N_23221);
and UO_1183 (O_1183,N_24073,N_23575);
nor UO_1184 (O_1184,N_21032,N_23700);
nor UO_1185 (O_1185,N_24454,N_22433);
or UO_1186 (O_1186,N_22187,N_24983);
nor UO_1187 (O_1187,N_20926,N_22752);
xnor UO_1188 (O_1188,N_22168,N_22364);
xnor UO_1189 (O_1189,N_22824,N_21621);
nand UO_1190 (O_1190,N_21574,N_20896);
nor UO_1191 (O_1191,N_24353,N_24392);
or UO_1192 (O_1192,N_21906,N_23073);
nor UO_1193 (O_1193,N_23705,N_23630);
nand UO_1194 (O_1194,N_23811,N_20588);
and UO_1195 (O_1195,N_24170,N_21526);
and UO_1196 (O_1196,N_21086,N_20697);
nor UO_1197 (O_1197,N_24130,N_23362);
or UO_1198 (O_1198,N_21758,N_24881);
nor UO_1199 (O_1199,N_24818,N_20158);
or UO_1200 (O_1200,N_21848,N_21453);
or UO_1201 (O_1201,N_23138,N_22498);
nor UO_1202 (O_1202,N_24461,N_20408);
nand UO_1203 (O_1203,N_21646,N_20431);
and UO_1204 (O_1204,N_20441,N_21375);
and UO_1205 (O_1205,N_22483,N_24902);
nand UO_1206 (O_1206,N_24978,N_23602);
nand UO_1207 (O_1207,N_20285,N_20312);
or UO_1208 (O_1208,N_20831,N_20728);
nand UO_1209 (O_1209,N_23244,N_20675);
nand UO_1210 (O_1210,N_23405,N_20421);
xnor UO_1211 (O_1211,N_22251,N_22539);
or UO_1212 (O_1212,N_21968,N_21373);
or UO_1213 (O_1213,N_20066,N_24375);
or UO_1214 (O_1214,N_21675,N_20559);
nor UO_1215 (O_1215,N_23401,N_23698);
xor UO_1216 (O_1216,N_21156,N_22190);
nor UO_1217 (O_1217,N_21581,N_20578);
and UO_1218 (O_1218,N_20743,N_24639);
and UO_1219 (O_1219,N_20608,N_21383);
xnor UO_1220 (O_1220,N_22840,N_21887);
nand UO_1221 (O_1221,N_23731,N_20281);
xor UO_1222 (O_1222,N_21839,N_21111);
xor UO_1223 (O_1223,N_23648,N_24764);
or UO_1224 (O_1224,N_20085,N_22500);
nand UO_1225 (O_1225,N_22012,N_21235);
xnor UO_1226 (O_1226,N_24068,N_21404);
or UO_1227 (O_1227,N_21281,N_23528);
xor UO_1228 (O_1228,N_23751,N_24751);
nand UO_1229 (O_1229,N_20075,N_21145);
nor UO_1230 (O_1230,N_23552,N_23038);
xnor UO_1231 (O_1231,N_23561,N_22928);
nand UO_1232 (O_1232,N_24152,N_22930);
or UO_1233 (O_1233,N_23606,N_20767);
or UO_1234 (O_1234,N_24177,N_20237);
and UO_1235 (O_1235,N_22259,N_20731);
nand UO_1236 (O_1236,N_24752,N_21599);
xnor UO_1237 (O_1237,N_23350,N_23410);
and UO_1238 (O_1238,N_22554,N_20886);
nor UO_1239 (O_1239,N_20009,N_22993);
and UO_1240 (O_1240,N_23399,N_22458);
nor UO_1241 (O_1241,N_21458,N_22357);
nor UO_1242 (O_1242,N_21207,N_21594);
nor UO_1243 (O_1243,N_24544,N_21476);
nand UO_1244 (O_1244,N_24129,N_22920);
or UO_1245 (O_1245,N_23390,N_21381);
and UO_1246 (O_1246,N_23164,N_24381);
xor UO_1247 (O_1247,N_23327,N_22853);
or UO_1248 (O_1248,N_23442,N_22188);
nand UO_1249 (O_1249,N_20353,N_24747);
or UO_1250 (O_1250,N_23347,N_20828);
nand UO_1251 (O_1251,N_22828,N_24700);
and UO_1252 (O_1252,N_23737,N_21702);
nor UO_1253 (O_1253,N_23493,N_24453);
nor UO_1254 (O_1254,N_23618,N_21355);
nor UO_1255 (O_1255,N_21415,N_24165);
xnor UO_1256 (O_1256,N_24443,N_21935);
and UO_1257 (O_1257,N_20741,N_21810);
xnor UO_1258 (O_1258,N_24692,N_22069);
and UO_1259 (O_1259,N_20364,N_23219);
nand UO_1260 (O_1260,N_24610,N_22059);
nand UO_1261 (O_1261,N_23499,N_24650);
or UO_1262 (O_1262,N_24949,N_22098);
or UO_1263 (O_1263,N_21435,N_23842);
nor UO_1264 (O_1264,N_23720,N_24072);
nand UO_1265 (O_1265,N_21243,N_21850);
or UO_1266 (O_1266,N_23502,N_24304);
nand UO_1267 (O_1267,N_24216,N_24006);
or UO_1268 (O_1268,N_21522,N_23181);
nand UO_1269 (O_1269,N_22533,N_23200);
nand UO_1270 (O_1270,N_23967,N_21778);
nor UO_1271 (O_1271,N_22344,N_22480);
nand UO_1272 (O_1272,N_23837,N_23139);
xor UO_1273 (O_1273,N_23870,N_21971);
or UO_1274 (O_1274,N_21033,N_21739);
nor UO_1275 (O_1275,N_22715,N_22216);
nand UO_1276 (O_1276,N_21618,N_22504);
nor UO_1277 (O_1277,N_24735,N_22260);
or UO_1278 (O_1278,N_21718,N_20960);
and UO_1279 (O_1279,N_22245,N_23873);
xor UO_1280 (O_1280,N_24404,N_22062);
nand UO_1281 (O_1281,N_20953,N_21559);
and UO_1282 (O_1282,N_20392,N_23590);
nand UO_1283 (O_1283,N_21397,N_23763);
or UO_1284 (O_1284,N_23034,N_24249);
and UO_1285 (O_1285,N_24261,N_22296);
and UO_1286 (O_1286,N_24823,N_21772);
and UO_1287 (O_1287,N_20064,N_20639);
or UO_1288 (O_1288,N_20298,N_23905);
or UO_1289 (O_1289,N_20478,N_20221);
xor UO_1290 (O_1290,N_20872,N_22262);
xor UO_1291 (O_1291,N_20121,N_21189);
or UO_1292 (O_1292,N_20401,N_20656);
nand UO_1293 (O_1293,N_24008,N_21504);
xor UO_1294 (O_1294,N_24917,N_24167);
nor UO_1295 (O_1295,N_24148,N_20574);
and UO_1296 (O_1296,N_20625,N_21654);
or UO_1297 (O_1297,N_24238,N_23836);
nor UO_1298 (O_1298,N_22999,N_21009);
or UO_1299 (O_1299,N_20147,N_20852);
nor UO_1300 (O_1300,N_23323,N_22944);
or UO_1301 (O_1301,N_24000,N_22974);
nor UO_1302 (O_1302,N_22107,N_22852);
nor UO_1303 (O_1303,N_20622,N_24621);
xnor UO_1304 (O_1304,N_24964,N_21141);
nor UO_1305 (O_1305,N_20602,N_23291);
xnor UO_1306 (O_1306,N_24001,N_23216);
or UO_1307 (O_1307,N_20484,N_20760);
or UO_1308 (O_1308,N_22367,N_24725);
nor UO_1309 (O_1309,N_24943,N_20318);
nand UO_1310 (O_1310,N_23860,N_23604);
xor UO_1311 (O_1311,N_23496,N_20748);
nor UO_1312 (O_1312,N_23397,N_21365);
nor UO_1313 (O_1313,N_24616,N_20351);
or UO_1314 (O_1314,N_21394,N_22013);
or UO_1315 (O_1315,N_21132,N_22218);
xor UO_1316 (O_1316,N_24549,N_20719);
or UO_1317 (O_1317,N_23525,N_20615);
nor UO_1318 (O_1318,N_22024,N_20012);
and UO_1319 (O_1319,N_21096,N_21958);
nand UO_1320 (O_1320,N_21093,N_23366);
nor UO_1321 (O_1321,N_21210,N_24184);
and UO_1322 (O_1322,N_23376,N_22629);
or UO_1323 (O_1323,N_20412,N_21591);
nand UO_1324 (O_1324,N_21883,N_24769);
and UO_1325 (O_1325,N_24225,N_20019);
nor UO_1326 (O_1326,N_20368,N_22654);
and UO_1327 (O_1327,N_20680,N_23413);
nor UO_1328 (O_1328,N_23142,N_23792);
or UO_1329 (O_1329,N_23006,N_21042);
nand UO_1330 (O_1330,N_24078,N_21730);
nand UO_1331 (O_1331,N_21994,N_24210);
or UO_1332 (O_1332,N_22584,N_23047);
nor UO_1333 (O_1333,N_24952,N_23831);
xnor UO_1334 (O_1334,N_24317,N_24445);
nand UO_1335 (O_1335,N_23300,N_21771);
or UO_1336 (O_1336,N_24297,N_21134);
and UO_1337 (O_1337,N_22440,N_20703);
or UO_1338 (O_1338,N_20062,N_21969);
nand UO_1339 (O_1339,N_23459,N_24880);
nand UO_1340 (O_1340,N_20128,N_20358);
nor UO_1341 (O_1341,N_22726,N_23222);
nand UO_1342 (O_1342,N_21313,N_21241);
nand UO_1343 (O_1343,N_23312,N_22114);
and UO_1344 (O_1344,N_20533,N_22229);
nand UO_1345 (O_1345,N_23852,N_23688);
xnor UO_1346 (O_1346,N_24853,N_21472);
and UO_1347 (O_1347,N_20580,N_21139);
nand UO_1348 (O_1348,N_24520,N_21783);
or UO_1349 (O_1349,N_20965,N_20716);
nor UO_1350 (O_1350,N_24181,N_24253);
nor UO_1351 (O_1351,N_21408,N_21364);
xor UO_1352 (O_1352,N_21123,N_23728);
and UO_1353 (O_1353,N_22825,N_21880);
nor UO_1354 (O_1354,N_23537,N_20907);
and UO_1355 (O_1355,N_20736,N_20848);
nor UO_1356 (O_1356,N_22203,N_20547);
nor UO_1357 (O_1357,N_24679,N_23546);
or UO_1358 (O_1358,N_21327,N_20857);
and UO_1359 (O_1359,N_23620,N_23007);
and UO_1360 (O_1360,N_21585,N_24052);
and UO_1361 (O_1361,N_22217,N_21531);
nor UO_1362 (O_1362,N_24064,N_24429);
and UO_1363 (O_1363,N_21715,N_20179);
and UO_1364 (O_1364,N_24913,N_21918);
and UO_1365 (O_1365,N_23642,N_21925);
nor UO_1366 (O_1366,N_21424,N_20342);
nand UO_1367 (O_1367,N_23913,N_22626);
nand UO_1368 (O_1368,N_23048,N_22372);
xnor UO_1369 (O_1369,N_20434,N_20499);
and UO_1370 (O_1370,N_22772,N_23765);
xor UO_1371 (O_1371,N_24110,N_20804);
nor UO_1372 (O_1372,N_22890,N_20199);
xnor UO_1373 (O_1373,N_23524,N_23775);
and UO_1374 (O_1374,N_21264,N_21538);
nor UO_1375 (O_1375,N_23369,N_21844);
or UO_1376 (O_1376,N_23657,N_23619);
and UO_1377 (O_1377,N_21240,N_24247);
nor UO_1378 (O_1378,N_21294,N_24248);
nand UO_1379 (O_1379,N_22514,N_20161);
nand UO_1380 (O_1380,N_24138,N_22858);
or UO_1381 (O_1381,N_20648,N_20390);
and UO_1382 (O_1382,N_21860,N_22496);
nand UO_1383 (O_1383,N_20090,N_20280);
nand UO_1384 (O_1384,N_24200,N_24775);
nor UO_1385 (O_1385,N_20393,N_22254);
nand UO_1386 (O_1386,N_20001,N_20520);
nor UO_1387 (O_1387,N_20650,N_23908);
and UO_1388 (O_1388,N_22612,N_24262);
xor UO_1389 (O_1389,N_20853,N_23743);
nor UO_1390 (O_1390,N_21779,N_20777);
or UO_1391 (O_1391,N_23482,N_22986);
xor UO_1392 (O_1392,N_20323,N_21483);
nand UO_1393 (O_1393,N_24385,N_22859);
or UO_1394 (O_1394,N_22213,N_20946);
and UO_1395 (O_1395,N_24303,N_20304);
and UO_1396 (O_1396,N_21631,N_22457);
nor UO_1397 (O_1397,N_20052,N_22037);
or UO_1398 (O_1398,N_20498,N_21322);
or UO_1399 (O_1399,N_20091,N_21716);
or UO_1400 (O_1400,N_23600,N_24877);
or UO_1401 (O_1401,N_22833,N_20183);
nand UO_1402 (O_1402,N_20824,N_20095);
xnor UO_1403 (O_1403,N_20897,N_23252);
and UO_1404 (O_1404,N_23342,N_23377);
or UO_1405 (O_1405,N_21919,N_24295);
or UO_1406 (O_1406,N_23378,N_21295);
xnor UO_1407 (O_1407,N_20814,N_20979);
xnor UO_1408 (O_1408,N_21856,N_23027);
xor UO_1409 (O_1409,N_21492,N_20573);
and UO_1410 (O_1410,N_20132,N_21590);
and UO_1411 (O_1411,N_22551,N_23100);
xnor UO_1412 (O_1412,N_22819,N_22278);
xor UO_1413 (O_1413,N_20028,N_24329);
and UO_1414 (O_1414,N_24634,N_23856);
xnor UO_1415 (O_1415,N_20284,N_21519);
or UO_1416 (O_1416,N_21449,N_21320);
and UO_1417 (O_1417,N_24504,N_21031);
or UO_1418 (O_1418,N_21273,N_21323);
nand UO_1419 (O_1419,N_21202,N_24580);
xnor UO_1420 (O_1420,N_24530,N_23091);
nor UO_1421 (O_1421,N_23250,N_21561);
nor UO_1422 (O_1422,N_22567,N_22721);
and UO_1423 (O_1423,N_24115,N_24630);
nor UO_1424 (O_1424,N_22845,N_20184);
or UO_1425 (O_1425,N_24172,N_22283);
and UO_1426 (O_1426,N_22329,N_20440);
xor UO_1427 (O_1427,N_20874,N_24923);
nand UO_1428 (O_1428,N_24844,N_24427);
nor UO_1429 (O_1429,N_24511,N_21983);
and UO_1430 (O_1430,N_21460,N_21274);
or UO_1431 (O_1431,N_22655,N_23444);
and UO_1432 (O_1432,N_21634,N_21366);
nand UO_1433 (O_1433,N_21021,N_21558);
nand UO_1434 (O_1434,N_23474,N_20501);
nor UO_1435 (O_1435,N_20307,N_22016);
nor UO_1436 (O_1436,N_22390,N_22511);
nand UO_1437 (O_1437,N_21637,N_20117);
nand UO_1438 (O_1438,N_21187,N_23558);
nor UO_1439 (O_1439,N_20978,N_24382);
xnor UO_1440 (O_1440,N_22227,N_23453);
nand UO_1441 (O_1441,N_24028,N_20110);
xor UO_1442 (O_1442,N_21798,N_23135);
or UO_1443 (O_1443,N_24772,N_23318);
nor UO_1444 (O_1444,N_21326,N_21633);
and UO_1445 (O_1445,N_22047,N_22678);
nor UO_1446 (O_1446,N_24768,N_20610);
nand UO_1447 (O_1447,N_21246,N_23960);
xnor UO_1448 (O_1448,N_21700,N_23249);
nand UO_1449 (O_1449,N_21046,N_24942);
nor UO_1450 (O_1450,N_20563,N_21013);
and UO_1451 (O_1451,N_21339,N_20565);
or UO_1452 (O_1452,N_23938,N_20921);
nor UO_1453 (O_1453,N_23954,N_22384);
or UO_1454 (O_1454,N_23018,N_21142);
and UO_1455 (O_1455,N_21909,N_21212);
nor UO_1456 (O_1456,N_23788,N_22406);
xnor UO_1457 (O_1457,N_23681,N_22388);
or UO_1458 (O_1458,N_22064,N_20372);
xor UO_1459 (O_1459,N_21144,N_21582);
nor UO_1460 (O_1460,N_20781,N_23738);
nand UO_1461 (O_1461,N_24252,N_20836);
xnor UO_1462 (O_1462,N_21498,N_24594);
or UO_1463 (O_1463,N_23926,N_22942);
or UO_1464 (O_1464,N_22720,N_23292);
nor UO_1465 (O_1465,N_22025,N_23963);
nand UO_1466 (O_1466,N_20634,N_22180);
nor UO_1467 (O_1467,N_24396,N_20251);
nor UO_1468 (O_1468,N_22238,N_21760);
nor UO_1469 (O_1469,N_23588,N_20092);
and UO_1470 (O_1470,N_22987,N_20171);
nor UO_1471 (O_1471,N_23517,N_22293);
nand UO_1472 (O_1472,N_21291,N_24346);
and UO_1473 (O_1473,N_21862,N_20655);
or UO_1474 (O_1474,N_22632,N_21745);
xnor UO_1475 (O_1475,N_21564,N_20369);
nor UO_1476 (O_1476,N_23446,N_22997);
or UO_1477 (O_1477,N_24599,N_23587);
xor UO_1478 (O_1478,N_20985,N_22137);
nand UO_1479 (O_1479,N_24009,N_20725);
nor UO_1480 (O_1480,N_20181,N_23277);
xnor UO_1481 (O_1481,N_23266,N_20468);
or UO_1482 (O_1482,N_20014,N_23979);
or UO_1483 (O_1483,N_22806,N_22954);
and UO_1484 (O_1484,N_23851,N_23227);
nor UO_1485 (O_1485,N_23435,N_24729);
xnor UO_1486 (O_1486,N_20007,N_22248);
nor UO_1487 (O_1487,N_20787,N_23217);
nand UO_1488 (O_1488,N_22967,N_23627);
nand UO_1489 (O_1489,N_20040,N_21669);
and UO_1490 (O_1490,N_22131,N_23946);
or UO_1491 (O_1491,N_21107,N_24264);
nor UO_1492 (O_1492,N_21682,N_22397);
xor UO_1493 (O_1493,N_22320,N_23095);
nor UO_1494 (O_1494,N_22021,N_20153);
nor UO_1495 (O_1495,N_23562,N_21949);
nor UO_1496 (O_1496,N_24538,N_22674);
or UO_1497 (O_1497,N_22309,N_20190);
xnor UO_1498 (O_1498,N_20485,N_24015);
and UO_1499 (O_1499,N_20708,N_20399);
xor UO_1500 (O_1500,N_22637,N_24894);
nand UO_1501 (O_1501,N_20870,N_20350);
nor UO_1502 (O_1502,N_21920,N_20306);
nor UO_1503 (O_1503,N_21229,N_21349);
nand UO_1504 (O_1504,N_21015,N_20021);
xor UO_1505 (O_1505,N_24697,N_20265);
xor UO_1506 (O_1506,N_22323,N_23145);
xor UO_1507 (O_1507,N_20611,N_23077);
or UO_1508 (O_1508,N_22246,N_22447);
or UO_1509 (O_1509,N_23146,N_22077);
nor UO_1510 (O_1510,N_21589,N_24242);
nand UO_1511 (O_1511,N_20045,N_24920);
nand UO_1512 (O_1512,N_24783,N_23321);
nand UO_1513 (O_1513,N_23075,N_22284);
nand UO_1514 (O_1514,N_22599,N_24293);
nand UO_1515 (O_1515,N_24430,N_21776);
or UO_1516 (O_1516,N_21085,N_20762);
and UO_1517 (O_1517,N_21287,N_24763);
nor UO_1518 (O_1518,N_22286,N_21814);
and UO_1519 (O_1519,N_22580,N_22783);
xnor UO_1520 (O_1520,N_23452,N_23060);
and UO_1521 (O_1521,N_23719,N_21362);
nand UO_1522 (O_1522,N_21112,N_21233);
xnor UO_1523 (O_1523,N_22200,N_21849);
and UO_1524 (O_1524,N_24423,N_22068);
nand UO_1525 (O_1525,N_21628,N_22635);
xnor UO_1526 (O_1526,N_24865,N_21596);
and UO_1527 (O_1527,N_23957,N_23750);
nor UO_1528 (O_1528,N_22849,N_23283);
or UO_1529 (O_1529,N_21794,N_22243);
or UO_1530 (O_1530,N_22154,N_21828);
xnor UO_1531 (O_1531,N_20813,N_22297);
xnor UO_1532 (O_1532,N_22383,N_23265);
or UO_1533 (O_1533,N_24848,N_23371);
nand UO_1534 (O_1534,N_20301,N_22817);
nor UO_1535 (O_1535,N_21609,N_23426);
or UO_1536 (O_1536,N_21098,N_23174);
and UO_1537 (O_1537,N_21796,N_20806);
and UO_1538 (O_1538,N_23832,N_23859);
or UO_1539 (O_1539,N_20305,N_20321);
nand UO_1540 (O_1540,N_23718,N_20141);
nand UO_1541 (O_1541,N_22512,N_22879);
xnor UO_1542 (O_1542,N_21780,N_24900);
nand UO_1543 (O_1543,N_22116,N_22641);
xor UO_1544 (O_1544,N_23117,N_22445);
or UO_1545 (O_1545,N_21952,N_21407);
or UO_1546 (O_1546,N_20508,N_24637);
xnor UO_1547 (O_1547,N_23166,N_23328);
and UO_1548 (O_1548,N_23535,N_21447);
and UO_1549 (O_1549,N_22875,N_24845);
nand UO_1550 (O_1550,N_20105,N_23186);
nand UO_1551 (O_1551,N_20258,N_24939);
nand UO_1552 (O_1552,N_22099,N_22781);
xnor UO_1553 (O_1553,N_20277,N_21485);
nand UO_1554 (O_1554,N_24321,N_21782);
nor UO_1555 (O_1555,N_24654,N_22060);
or UO_1556 (O_1556,N_20968,N_22614);
nand UO_1557 (O_1557,N_21316,N_20699);
nand UO_1558 (O_1558,N_22530,N_20821);
and UO_1559 (O_1559,N_20653,N_21683);
nand UO_1560 (O_1560,N_24113,N_21395);
nand UO_1561 (O_1561,N_24369,N_20658);
or UO_1562 (O_1562,N_22468,N_23673);
nand UO_1563 (O_1563,N_23074,N_22690);
and UO_1564 (O_1564,N_21749,N_20327);
nand UO_1565 (O_1565,N_20835,N_21208);
xor UO_1566 (O_1566,N_24873,N_21376);
and UO_1567 (O_1567,N_24474,N_20952);
xor UO_1568 (O_1568,N_22860,N_24183);
nand UO_1569 (O_1569,N_21583,N_24251);
xnor UO_1570 (O_1570,N_20418,N_23049);
and UO_1571 (O_1571,N_24406,N_24278);
and UO_1572 (O_1572,N_23695,N_23532);
xnor UO_1573 (O_1573,N_24188,N_22902);
xor UO_1574 (O_1574,N_21932,N_21260);
nand UO_1575 (O_1575,N_20104,N_22182);
nand UO_1576 (O_1576,N_22966,N_21310);
nor UO_1577 (O_1577,N_22714,N_21044);
and UO_1578 (O_1578,N_23133,N_21955);
xnor UO_1579 (O_1579,N_24812,N_22793);
nand UO_1580 (O_1580,N_22671,N_23566);
or UO_1581 (O_1581,N_20516,N_23754);
xor UO_1582 (O_1582,N_23021,N_21649);
nand UO_1583 (O_1583,N_21943,N_20587);
nor UO_1584 (O_1584,N_21285,N_24595);
xnor UO_1585 (O_1585,N_22418,N_23198);
nand UO_1586 (O_1586,N_21544,N_23106);
nand UO_1587 (O_1587,N_20343,N_24163);
and UO_1588 (O_1588,N_22892,N_24786);
and UO_1589 (O_1589,N_20581,N_24400);
and UO_1590 (O_1590,N_23260,N_22199);
nand UO_1591 (O_1591,N_22959,N_24745);
nand UO_1592 (O_1592,N_24653,N_23230);
nand UO_1593 (O_1593,N_20596,N_20909);
and UO_1594 (O_1594,N_20754,N_24102);
nor UO_1595 (O_1595,N_22083,N_24027);
nor UO_1596 (O_1596,N_22431,N_23349);
or UO_1597 (O_1597,N_23801,N_23998);
nor UO_1598 (O_1598,N_24155,N_24442);
nor UO_1599 (O_1599,N_24341,N_22023);
nor UO_1600 (O_1600,N_22558,N_24025);
or UO_1601 (O_1601,N_23507,N_22759);
and UO_1602 (O_1602,N_24473,N_21385);
xor UO_1603 (O_1603,N_24069,N_20296);
nand UO_1604 (O_1604,N_20932,N_20832);
nor UO_1605 (O_1605,N_20727,N_24625);
nand UO_1606 (O_1606,N_23134,N_24801);
and UO_1607 (O_1607,N_24038,N_20937);
nor UO_1608 (O_1608,N_22735,N_21293);
nand UO_1609 (O_1609,N_23404,N_23130);
nor UO_1610 (O_1610,N_20053,N_24214);
or UO_1611 (O_1611,N_22699,N_22676);
or UO_1612 (O_1612,N_20309,N_20362);
xor UO_1613 (O_1613,N_21351,N_22493);
nand UO_1614 (O_1614,N_21128,N_23143);
and UO_1615 (O_1615,N_20943,N_21147);
or UO_1616 (O_1616,N_22836,N_23020);
or UO_1617 (O_1617,N_22872,N_24987);
and UO_1618 (O_1618,N_23791,N_23337);
xor UO_1619 (O_1619,N_20231,N_24081);
and UO_1620 (O_1620,N_20169,N_21870);
nand UO_1621 (O_1621,N_24411,N_22829);
or UO_1622 (O_1622,N_21895,N_24668);
nand UO_1623 (O_1623,N_23019,N_21744);
and UO_1624 (O_1624,N_23172,N_24399);
xnor UO_1625 (O_1625,N_22434,N_21359);
xor UO_1626 (O_1626,N_20527,N_22864);
or UO_1627 (O_1627,N_23414,N_21090);
xor UO_1628 (O_1628,N_20673,N_22566);
or UO_1629 (O_1629,N_20967,N_21827);
xnor UO_1630 (O_1630,N_23675,N_21338);
and UO_1631 (O_1631,N_20134,N_21752);
xor UO_1632 (O_1632,N_22055,N_21309);
nand UO_1633 (O_1633,N_24906,N_21311);
nand UO_1634 (O_1634,N_24316,N_24797);
xnor UO_1635 (O_1635,N_23037,N_24562);
or UO_1636 (O_1636,N_24564,N_20562);
and UO_1637 (O_1637,N_22595,N_24791);
nand UO_1638 (O_1638,N_24257,N_21868);
and UO_1639 (O_1639,N_23893,N_20592);
xor UO_1640 (O_1640,N_22147,N_20144);
or UO_1641 (O_1641,N_20457,N_23591);
or UO_1642 (O_1642,N_22711,N_22906);
xnor UO_1643 (O_1643,N_23576,N_23159);
nor UO_1644 (O_1644,N_24362,N_24804);
xor UO_1645 (O_1645,N_21626,N_24267);
nor UO_1646 (O_1646,N_22804,N_21666);
and UO_1647 (O_1647,N_21924,N_21149);
nor UO_1648 (O_1648,N_20627,N_22943);
nor UO_1649 (O_1649,N_22740,N_22268);
xnor UO_1650 (O_1650,N_22855,N_21837);
xor UO_1651 (O_1651,N_20769,N_22841);
nor UO_1652 (O_1652,N_21078,N_24330);
nand UO_1653 (O_1653,N_24790,N_24644);
and UO_1654 (O_1654,N_22419,N_24020);
or UO_1655 (O_1655,N_24093,N_21539);
nand UO_1656 (O_1656,N_22577,N_20586);
xor UO_1657 (O_1657,N_23406,N_24359);
nand UO_1658 (O_1658,N_22665,N_21499);
or UO_1659 (O_1659,N_23123,N_23403);
or UO_1660 (O_1660,N_24298,N_21290);
xnor UO_1661 (O_1661,N_24959,N_21048);
and UO_1662 (O_1662,N_24973,N_20651);
xnor UO_1663 (O_1663,N_24213,N_20198);
nor UO_1664 (O_1664,N_24581,N_20391);
and UO_1665 (O_1665,N_20008,N_21043);
xor UO_1666 (O_1666,N_20458,N_20936);
nor UO_1667 (O_1667,N_24016,N_22949);
and UO_1668 (O_1668,N_20755,N_23846);
or UO_1669 (O_1669,N_23432,N_22008);
nand UO_1670 (O_1670,N_21340,N_21520);
and UO_1671 (O_1671,N_20515,N_20389);
and UO_1672 (O_1672,N_21297,N_20855);
nor UO_1673 (O_1673,N_22761,N_23940);
and UO_1674 (O_1674,N_24144,N_21026);
or UO_1675 (O_1675,N_23023,N_23682);
or UO_1676 (O_1676,N_21169,N_24047);
and UO_1677 (O_1677,N_24343,N_20529);
and UO_1678 (O_1678,N_23407,N_24771);
and UO_1679 (O_1679,N_22415,N_23821);
xor UO_1680 (O_1680,N_21985,N_20539);
xor UO_1681 (O_1681,N_24535,N_22026);
nand UO_1682 (O_1682,N_24875,N_20782);
and UO_1683 (O_1683,N_21321,N_20679);
nand UO_1684 (O_1684,N_21190,N_22330);
nand UO_1685 (O_1685,N_20542,N_23996);
nand UO_1686 (O_1686,N_22103,N_23296);
xnor UO_1687 (O_1687,N_23461,N_22693);
nand UO_1688 (O_1688,N_20055,N_21537);
and UO_1689 (O_1689,N_23381,N_21703);
xor UO_1690 (O_1690,N_24118,N_23110);
and UO_1691 (O_1691,N_20332,N_20628);
nand UO_1692 (O_1692,N_22231,N_22004);
nand UO_1693 (O_1693,N_24339,N_21463);
and UO_1694 (O_1694,N_24119,N_24693);
xor UO_1695 (O_1695,N_23733,N_20827);
nand UO_1696 (O_1696,N_22104,N_21699);
xnor UO_1697 (O_1697,N_22489,N_24439);
nand UO_1698 (O_1698,N_21640,N_22837);
and UO_1699 (O_1699,N_22192,N_23322);
xor UO_1700 (O_1700,N_22748,N_23207);
nand UO_1701 (O_1701,N_20490,N_22611);
nor UO_1702 (O_1702,N_24897,N_20425);
or UO_1703 (O_1703,N_21691,N_20850);
or UO_1704 (O_1704,N_21428,N_23182);
and UO_1705 (O_1705,N_21562,N_24776);
or UO_1706 (O_1706,N_22179,N_23959);
nand UO_1707 (O_1707,N_21607,N_21959);
nor UO_1708 (O_1708,N_23804,N_24061);
nor UO_1709 (O_1709,N_22553,N_22736);
or UO_1710 (O_1710,N_24999,N_23040);
or UO_1711 (O_1711,N_20299,N_21109);
or UO_1712 (O_1712,N_24500,N_20234);
xor UO_1713 (O_1713,N_22722,N_24499);
xor UO_1714 (O_1714,N_20891,N_24574);
nor UO_1715 (O_1715,N_24641,N_20363);
xor UO_1716 (O_1716,N_22310,N_24370);
nand UO_1717 (O_1717,N_22716,N_22070);
nand UO_1718 (O_1718,N_22417,N_20079);
nor UO_1719 (O_1719,N_23096,N_24811);
and UO_1720 (O_1720,N_21221,N_24661);
and UO_1721 (O_1721,N_22976,N_21378);
xnor UO_1722 (O_1722,N_21510,N_24798);
nor UO_1723 (O_1723,N_22276,N_21368);
and UO_1724 (O_1724,N_24348,N_21635);
xnor UO_1725 (O_1725,N_23441,N_24546);
and UO_1726 (O_1726,N_24998,N_22564);
nand UO_1727 (O_1727,N_24607,N_21516);
or UO_1728 (O_1728,N_22914,N_24629);
and UO_1729 (O_1729,N_24036,N_24065);
nand UO_1730 (O_1730,N_22050,N_20910);
xor UO_1731 (O_1731,N_22302,N_23748);
or UO_1732 (O_1732,N_20427,N_24246);
xnor UO_1733 (O_1733,N_21667,N_20545);
xor UO_1734 (O_1734,N_24814,N_20146);
xnor UO_1735 (O_1735,N_23565,N_20302);
and UO_1736 (O_1736,N_20027,N_21580);
nor UO_1737 (O_1737,N_24486,N_21899);
xor UO_1738 (O_1738,N_24796,N_24309);
xnor UO_1739 (O_1739,N_24431,N_20279);
nor UO_1740 (O_1740,N_22758,N_22441);
nor UO_1741 (O_1741,N_20345,N_23867);
or UO_1742 (O_1742,N_23741,N_20380);
or UO_1743 (O_1743,N_20717,N_24565);
and UO_1744 (O_1744,N_24426,N_20172);
or UO_1745 (O_1745,N_23245,N_21941);
nand UO_1746 (O_1746,N_24342,N_23386);
nand UO_1747 (O_1747,N_21964,N_21550);
nand UO_1748 (O_1748,N_21506,N_21536);
nor UO_1749 (O_1749,N_24447,N_22430);
nand UO_1750 (O_1750,N_23825,N_22543);
or UO_1751 (O_1751,N_24145,N_23030);
or UO_1752 (O_1752,N_23515,N_24049);
nor UO_1753 (O_1753,N_24737,N_20120);
xor UO_1754 (O_1754,N_23491,N_20589);
or UO_1755 (O_1755,N_24376,N_24709);
or UO_1756 (O_1756,N_21838,N_20058);
nand UO_1757 (O_1757,N_23835,N_20807);
and UO_1758 (O_1758,N_23686,N_20722);
nand UO_1759 (O_1759,N_20579,N_22886);
and UO_1760 (O_1760,N_21289,N_20750);
and UO_1761 (O_1761,N_23746,N_21016);
or UO_1762 (O_1762,N_20689,N_24887);
nor UO_1763 (O_1763,N_22867,N_20925);
or UO_1764 (O_1764,N_21871,N_23279);
and UO_1765 (O_1765,N_20061,N_23122);
nor UO_1766 (O_1766,N_24151,N_24388);
xnor UO_1767 (O_1767,N_23930,N_22857);
and UO_1768 (O_1768,N_22171,N_24308);
or UO_1769 (O_1769,N_20970,N_24807);
or UO_1770 (O_1770,N_24739,N_23246);
or UO_1771 (O_1771,N_24918,N_22672);
nor UO_1772 (O_1772,N_20241,N_22377);
nand UO_1773 (O_1773,N_23392,N_21400);
or UO_1774 (O_1774,N_21121,N_24048);
nand UO_1775 (O_1775,N_20213,N_20491);
nand UO_1776 (O_1776,N_21768,N_23778);
nand UO_1777 (O_1777,N_23658,N_22666);
nor UO_1778 (O_1778,N_20676,N_20663);
and UO_1779 (O_1779,N_23051,N_22922);
or UO_1780 (O_1780,N_22253,N_24583);
or UO_1781 (O_1781,N_21575,N_21087);
nor UO_1782 (O_1782,N_23906,N_20030);
or UO_1783 (O_1783,N_20664,N_21119);
nand UO_1784 (O_1784,N_23052,N_22336);
or UO_1785 (O_1785,N_24483,N_21158);
xor UO_1786 (O_1786,N_21214,N_21061);
nor UO_1787 (O_1787,N_20405,N_20433);
and UO_1788 (O_1788,N_23596,N_22882);
xnor UO_1789 (O_1789,N_21560,N_23341);
or UO_1790 (O_1790,N_23543,N_22684);
nand UO_1791 (O_1791,N_21625,N_21296);
or UO_1792 (O_1792,N_21331,N_24398);
or UO_1793 (O_1793,N_22982,N_20944);
nand UO_1794 (O_1794,N_22787,N_21807);
and UO_1795 (O_1795,N_20900,N_21711);
nand UO_1796 (O_1796,N_20751,N_20864);
and UO_1797 (O_1797,N_20016,N_21173);
xnor UO_1798 (O_1798,N_22889,N_24592);
nand UO_1799 (O_1799,N_20996,N_21114);
and UO_1800 (O_1800,N_22134,N_20250);
nand UO_1801 (O_1801,N_21823,N_24366);
xor UO_1802 (O_1802,N_21200,N_24336);
and UO_1803 (O_1803,N_20963,N_23806);
and UO_1804 (O_1804,N_22805,N_21065);
or UO_1805 (O_1805,N_22777,N_24556);
or UO_1806 (O_1806,N_20115,N_22628);
or UO_1807 (O_1807,N_24467,N_23914);
nor UO_1808 (O_1808,N_20006,N_24046);
xor UO_1809 (O_1809,N_20854,N_24187);
nor UO_1810 (O_1810,N_23595,N_23882);
and UO_1811 (O_1811,N_23625,N_23512);
nand UO_1812 (O_1812,N_20861,N_24585);
and UO_1813 (O_1813,N_23035,N_20976);
nand UO_1814 (O_1814,N_24759,N_23429);
nand UO_1815 (O_1815,N_21361,N_22464);
nor UO_1816 (O_1816,N_23628,N_20159);
and UO_1817 (O_1817,N_20877,N_24536);
or UO_1818 (O_1818,N_20335,N_23654);
nor UO_1819 (O_1819,N_21484,N_24492);
nand UO_1820 (O_1820,N_22118,N_21024);
nor UO_1821 (O_1821,N_22224,N_20830);
and UO_1822 (O_1822,N_23097,N_20486);
and UO_1823 (O_1823,N_20632,N_23137);
nand UO_1824 (O_1824,N_20119,N_23348);
and UO_1825 (O_1825,N_24518,N_24990);
and UO_1826 (O_1826,N_20386,N_22972);
nor UO_1827 (O_1827,N_20429,N_24356);
or UO_1828 (O_1828,N_24159,N_24657);
xor UO_1829 (O_1829,N_23408,N_21990);
xor UO_1830 (O_1830,N_22396,N_24864);
and UO_1831 (O_1831,N_24344,N_23215);
nor UO_1832 (O_1832,N_23165,N_20293);
nand UO_1833 (O_1833,N_21095,N_24347);
xor UO_1834 (O_1834,N_23177,N_23086);
and UO_1835 (O_1835,N_20904,N_23961);
nand UO_1836 (O_1836,N_23556,N_20860);
nor UO_1837 (O_1837,N_22528,N_23521);
nor UO_1838 (O_1838,N_24979,N_20966);
or UO_1839 (O_1839,N_22350,N_24335);
nand UO_1840 (O_1840,N_20883,N_23191);
xnor UO_1841 (O_1841,N_21570,N_23185);
nor UO_1842 (O_1842,N_21283,N_20669);
nor UO_1843 (O_1843,N_21961,N_23895);
xnor UO_1844 (O_1844,N_21965,N_24488);
and UO_1845 (O_1845,N_22896,N_21650);
and UO_1846 (O_1846,N_21897,N_21205);
or UO_1847 (O_1847,N_21056,N_21390);
and UO_1848 (O_1848,N_23189,N_23167);
and UO_1849 (O_1849,N_24086,N_20506);
nor UO_1850 (O_1850,N_24695,N_22694);
xor UO_1851 (O_1851,N_21982,N_23861);
or UO_1852 (O_1852,N_24724,N_22115);
xor UO_1853 (O_1853,N_23016,N_21150);
nor UO_1854 (O_1854,N_21438,N_21076);
nor UO_1855 (O_1855,N_22506,N_22568);
nor UO_1856 (O_1856,N_20819,N_21928);
and UO_1857 (O_1857,N_20283,N_20185);
nand UO_1858 (O_1858,N_23849,N_20630);
nor UO_1859 (O_1859,N_24743,N_23197);
nand UO_1860 (O_1860,N_24470,N_20303);
nand UO_1861 (O_1861,N_23516,N_22820);
and UO_1862 (O_1862,N_20894,N_24792);
nor UO_1863 (O_1863,N_20686,N_20050);
xnor UO_1864 (O_1864,N_22139,N_22170);
and UO_1865 (O_1865,N_23850,N_22688);
nor UO_1866 (O_1866,N_22092,N_22683);
nor UO_1867 (O_1867,N_21178,N_21541);
xnor UO_1868 (O_1868,N_20200,N_21071);
and UO_1869 (O_1869,N_20145,N_24090);
xor UO_1870 (O_1870,N_22620,N_20924);
nor UO_1871 (O_1871,N_20805,N_21184);
nand UO_1872 (O_1872,N_20201,N_24034);
nor UO_1873 (O_1873,N_23069,N_22045);
xnor UO_1874 (O_1874,N_24322,N_21734);
nand UO_1875 (O_1875,N_21655,N_23436);
nor UO_1876 (O_1876,N_20975,N_21244);
nor UO_1877 (O_1877,N_23355,N_24552);
nand UO_1878 (O_1878,N_24532,N_23900);
nor UO_1879 (O_1879,N_23437,N_22673);
xnor UO_1880 (O_1880,N_20988,N_22191);
xnor UO_1881 (O_1881,N_20037,N_20100);
nand UO_1882 (O_1882,N_21610,N_21248);
and UO_1883 (O_1883,N_22306,N_21645);
and UO_1884 (O_1884,N_20502,N_21529);
xnor UO_1885 (O_1885,N_24217,N_22421);
and UO_1886 (O_1886,N_21191,N_22932);
or UO_1887 (O_1887,N_22799,N_21879);
and UO_1888 (O_1888,N_24989,N_24858);
and UO_1889 (O_1889,N_20481,N_24795);
or UO_1890 (O_1890,N_24243,N_23385);
xnor UO_1891 (O_1891,N_22523,N_20242);
nor UO_1892 (O_1892,N_21330,N_22893);
and UO_1893 (O_1893,N_20652,N_24960);
nand UO_1894 (O_1894,N_23974,N_24254);
xnor UO_1895 (O_1895,N_23777,N_24788);
or UO_1896 (O_1896,N_21970,N_22904);
nor UO_1897 (O_1897,N_22266,N_21623);
xnor UO_1898 (O_1898,N_21419,N_23536);
nor UO_1899 (O_1899,N_23289,N_21528);
or UO_1900 (O_1900,N_23163,N_24414);
and UO_1901 (O_1901,N_22621,N_21733);
nand UO_1902 (O_1902,N_21371,N_22679);
and UO_1903 (O_1903,N_22778,N_22934);
and UO_1904 (O_1904,N_20130,N_24501);
and UO_1905 (O_1905,N_22818,N_24211);
nand UO_1906 (O_1906,N_21822,N_22261);
or UO_1907 (O_1907,N_22391,N_24051);
or UO_1908 (O_1908,N_20840,N_23070);
nor UO_1909 (O_1909,N_22700,N_24994);
or UO_1910 (O_1910,N_21440,N_24075);
xor UO_1911 (O_1911,N_20688,N_21100);
nor UO_1912 (O_1912,N_22034,N_24387);
nor UO_1913 (O_1913,N_20582,N_21825);
nand UO_1914 (O_1914,N_22540,N_24174);
xor UO_1915 (O_1915,N_23572,N_24189);
and UO_1916 (O_1916,N_23043,N_23065);
xnor UO_1917 (O_1917,N_21565,N_21741);
xnor UO_1918 (O_1918,N_20319,N_20756);
or UO_1919 (O_1919,N_21174,N_20371);
and UO_1920 (O_1920,N_20746,N_20888);
nand UO_1921 (O_1921,N_21152,N_20129);
nor UO_1922 (O_1922,N_22547,N_23968);
or UO_1923 (O_1923,N_21653,N_22113);
nand UO_1924 (O_1924,N_20166,N_22285);
or UO_1925 (O_1925,N_24648,N_20476);
nor UO_1926 (O_1926,N_23464,N_20033);
and UO_1927 (O_1927,N_22402,N_20734);
and UO_1928 (O_1928,N_24374,N_23275);
nand UO_1929 (O_1929,N_23379,N_21218);
nor UO_1930 (O_1930,N_23988,N_21671);
or UO_1931 (O_1931,N_22057,N_24365);
or UO_1932 (O_1932,N_24749,N_21791);
or UO_1933 (O_1933,N_20263,N_21489);
or UO_1934 (O_1934,N_20535,N_24977);
and UO_1935 (O_1935,N_20036,N_20357);
and UO_1936 (O_1936,N_21518,N_22610);
or UO_1937 (O_1937,N_24861,N_21006);
or UO_1938 (O_1938,N_24950,N_20906);
nor UO_1939 (O_1939,N_23554,N_24056);
nand UO_1940 (O_1940,N_24227,N_22289);
nor UO_1941 (O_1941,N_22575,N_22422);
nor UO_1942 (O_1942,N_24867,N_23534);
and UO_1943 (O_1943,N_20192,N_20382);
xor UO_1944 (O_1944,N_20678,N_20261);
nor UO_1945 (O_1945,N_23356,N_22953);
nor UO_1946 (O_1946,N_21138,N_20935);
nand UO_1947 (O_1947,N_23747,N_24100);
or UO_1948 (O_1948,N_24153,N_22385);
and UO_1949 (O_1949,N_21324,N_20659);
nand UO_1950 (O_1950,N_24810,N_20322);
nand UO_1951 (O_1951,N_20927,N_21933);
or UO_1952 (O_1952,N_20826,N_21225);
nor UO_1953 (O_1953,N_21811,N_23014);
nor UO_1954 (O_1954,N_22314,N_24465);
or UO_1955 (O_1955,N_21328,N_23608);
xor UO_1956 (O_1956,N_21769,N_23815);
or UO_1957 (O_1957,N_23915,N_21478);
nand UO_1958 (O_1958,N_24132,N_22717);
xnor UO_1959 (O_1959,N_23912,N_22557);
xor UO_1960 (O_1960,N_24930,N_23483);
nor UO_1961 (O_1961,N_20604,N_21957);
nand UO_1962 (O_1962,N_22791,N_23125);
nand UO_1963 (O_1963,N_23205,N_20446);
or UO_1964 (O_1964,N_20260,N_24698);
xnor UO_1965 (O_1965,N_21181,N_22136);
and UO_1966 (O_1966,N_23479,N_20859);
nor UO_1967 (O_1967,N_21552,N_21234);
or UO_1968 (O_1968,N_21853,N_21417);
xnor UO_1969 (O_1969,N_24761,N_21753);
nand UO_1970 (O_1970,N_22393,N_22981);
or UO_1971 (O_1971,N_22475,N_23422);
xnor UO_1972 (O_1972,N_24946,N_20949);
and UO_1973 (O_1973,N_22130,N_22542);
xnor UO_1974 (O_1974,N_21004,N_20712);
xor UO_1975 (O_1975,N_20882,N_24133);
and UO_1976 (O_1976,N_24513,N_22030);
xnor UO_1977 (O_1977,N_23050,N_22689);
and UO_1978 (O_1978,N_21379,N_21882);
or UO_1979 (O_1979,N_24962,N_23581);
xor UO_1980 (O_1980,N_24279,N_23488);
and UO_1981 (O_1981,N_24660,N_21279);
xnor UO_1982 (O_1982,N_24083,N_24147);
or UO_1983 (O_1983,N_22532,N_20177);
nor UO_1984 (O_1984,N_23234,N_23712);
and UO_1985 (O_1985,N_20452,N_21163);
xor UO_1986 (O_1986,N_20218,N_23154);
nor UO_1987 (O_1987,N_22537,N_24885);
nand UO_1988 (O_1988,N_21878,N_24126);
xor UO_1989 (O_1989,N_24435,N_23128);
nor UO_1990 (O_1990,N_23545,N_20275);
or UO_1991 (O_1991,N_20991,N_21058);
nand UO_1992 (O_1992,N_20328,N_20637);
nand UO_1993 (O_1993,N_21060,N_21442);
nor UO_1994 (O_1994,N_22127,N_21300);
and UO_1995 (O_1995,N_24337,N_20072);
xor UO_1996 (O_1996,N_24433,N_23989);
and UO_1997 (O_1997,N_20892,N_22270);
and UO_1998 (O_1998,N_23268,N_23304);
or UO_1999 (O_1999,N_24204,N_22087);
nor UO_2000 (O_2000,N_23402,N_21325);
xnor UO_2001 (O_2001,N_23918,N_20133);
or UO_2002 (O_2002,N_20942,N_20939);
xor UO_2003 (O_2003,N_22846,N_22850);
or UO_2004 (O_2004,N_22739,N_24911);
xnor UO_2005 (O_2005,N_21345,N_21192);
and UO_2006 (O_2006,N_22734,N_22035);
xnor UO_2007 (O_2007,N_23118,N_23952);
and UO_2008 (O_2008,N_20047,N_20135);
nand UO_2009 (O_2009,N_24910,N_23896);
nand UO_2010 (O_2010,N_24996,N_20796);
and UO_2011 (O_2011,N_22325,N_20692);
nor UO_2012 (O_2012,N_20487,N_21023);
nand UO_2013 (O_2013,N_23876,N_21161);
xnor UO_2014 (O_2014,N_22517,N_22544);
xnor UO_2015 (O_2015,N_22638,N_23495);
or UO_2016 (O_2016,N_20961,N_20825);
and UO_2017 (O_2017,N_24233,N_22495);
xnor UO_2018 (O_2018,N_22590,N_24802);
nand UO_2019 (O_2019,N_24451,N_22895);
nand UO_2020 (O_2020,N_23621,N_24106);
nand UO_2021 (O_2021,N_21641,N_24274);
or UO_2022 (O_2022,N_21130,N_21984);
or UO_2023 (O_2023,N_21073,N_22195);
nor UO_2024 (O_2024,N_24813,N_21067);
and UO_2025 (O_2025,N_24663,N_20729);
nor UO_2026 (O_2026,N_20645,N_24493);
nand UO_2027 (O_2027,N_23708,N_24497);
or UO_2028 (O_2028,N_22687,N_24655);
xor UO_2029 (O_2029,N_23313,N_21967);
nand UO_2030 (O_2030,N_21399,N_21923);
nor UO_2031 (O_2031,N_24773,N_23080);
nor UO_2032 (O_2032,N_23770,N_22648);
and UO_2033 (O_2033,N_23586,N_21002);
or UO_2034 (O_2034,N_21097,N_20288);
nor UO_2035 (O_2035,N_21259,N_24460);
xnor UO_2036 (O_2036,N_22152,N_22925);
or UO_2037 (O_2037,N_21972,N_23809);
nor UO_2038 (O_2038,N_21576,N_22443);
nand UO_2039 (O_2039,N_20584,N_21258);
and UO_2040 (O_2040,N_20901,N_21426);
nand UO_2041 (O_2041,N_24738,N_22705);
or UO_2042 (O_2042,N_24313,N_22236);
nand UO_2043 (O_2043,N_24058,N_22862);
xnor UO_2044 (O_2044,N_24750,N_24652);
nand UO_2045 (O_2045,N_21185,N_21336);
or UO_2046 (O_2046,N_20346,N_21439);
or UO_2047 (O_2047,N_24407,N_20745);
nand UO_2048 (O_2048,N_21595,N_23472);
or UO_2049 (O_2049,N_21137,N_20528);
nor UO_2050 (O_2050,N_21257,N_20605);
nor UO_2051 (O_2051,N_24403,N_20753);
nor UO_2052 (O_2052,N_21571,N_24259);
or UO_2053 (O_2053,N_20994,N_21253);
nand UO_2054 (O_2054,N_24856,N_21759);
and UO_2055 (O_2055,N_23923,N_22228);
or UO_2056 (O_2056,N_22747,N_24490);
nor UO_2057 (O_2057,N_21917,N_21481);
xor UO_2058 (O_2058,N_20995,N_23865);
and UO_2059 (O_2059,N_24548,N_20715);
or UO_2060 (O_2060,N_23001,N_24476);
nor UO_2061 (O_2061,N_22810,N_21473);
or UO_2062 (O_2062,N_22965,N_20205);
nor UO_2063 (O_2063,N_24292,N_24449);
and UO_2064 (O_2064,N_23756,N_21343);
or UO_2065 (O_2065,N_22607,N_23310);
nand UO_2066 (O_2066,N_23813,N_22148);
nand UO_2067 (O_2067,N_21104,N_21719);
or UO_2068 (O_2068,N_21081,N_24378);
and UO_2069 (O_2069,N_21956,N_24457);
or UO_2070 (O_2070,N_22600,N_20175);
or UO_2071 (O_2071,N_21873,N_23693);
and UO_2072 (O_2072,N_21505,N_20038);
nand UO_2073 (O_2073,N_21165,N_24627);
xnor UO_2074 (O_2074,N_23236,N_23655);
xnor UO_2075 (O_2075,N_20641,N_21551);
or UO_2076 (O_2076,N_21479,N_21602);
nand UO_2077 (O_2077,N_21592,N_23820);
xnor UO_2078 (O_2078,N_21079,N_24039);
and UO_2079 (O_2079,N_24393,N_21898);
nor UO_2080 (O_2080,N_22653,N_24567);
nor UO_2081 (O_2081,N_21663,N_23951);
or UO_2082 (O_2082,N_22039,N_23984);
or UO_2083 (O_2083,N_24192,N_22565);
nand UO_2084 (O_2084,N_24495,N_22907);
or UO_2085 (O_2085,N_23707,N_22386);
and UO_2086 (O_2086,N_21017,N_22072);
nand UO_2087 (O_2087,N_22851,N_20180);
nor UO_2088 (O_2088,N_24114,N_20376);
xor UO_2089 (O_2089,N_22497,N_20074);
and UO_2090 (O_2090,N_22919,N_22038);
nand UO_2091 (O_2091,N_21617,N_24302);
or UO_2092 (O_2092,N_20784,N_23577);
nand UO_2093 (O_2093,N_24667,N_22917);
nand UO_2094 (O_2094,N_21673,N_23526);
or UO_2095 (O_2095,N_23116,N_21188);
or UO_2096 (O_2096,N_22173,N_24673);
or UO_2097 (O_2097,N_24722,N_23500);
nand UO_2098 (O_2098,N_21884,N_21713);
nand UO_2099 (O_2099,N_23533,N_22020);
xnor UO_2100 (O_2100,N_24122,N_22215);
or UO_2101 (O_2101,N_23753,N_22345);
xor UO_2102 (O_2102,N_24059,N_24311);
and UO_2103 (O_2103,N_21411,N_20289);
nor UO_2104 (O_2104,N_24011,N_24260);
nand UO_2105 (O_2105,N_22206,N_23433);
nor UO_2106 (O_2106,N_21219,N_21157);
and UO_2107 (O_2107,N_23316,N_23000);
nand UO_2108 (O_2108,N_23352,N_21490);
xnor UO_2109 (O_2109,N_20710,N_20432);
nand UO_2110 (O_2110,N_20084,N_21406);
and UO_2111 (O_2111,N_20143,N_24803);
xor UO_2112 (O_2112,N_21261,N_22210);
or UO_2113 (O_2113,N_22927,N_23176);
nor UO_2114 (O_2114,N_22018,N_23173);
xnor UO_2115 (O_2115,N_22274,N_24018);
nand UO_2116 (O_2116,N_24471,N_21587);
nand UO_2117 (O_2117,N_24676,N_22178);
or UO_2118 (O_2118,N_23828,N_21996);
nor UO_2119 (O_2119,N_24350,N_21053);
nand UO_2120 (O_2120,N_24600,N_22327);
nor UO_2121 (O_2121,N_23169,N_23643);
xor UO_2122 (O_2122,N_22177,N_24448);
and UO_2123 (O_2123,N_21445,N_23540);
xnor UO_2124 (O_2124,N_23548,N_20480);
or UO_2125 (O_2125,N_24816,N_20331);
nor UO_2126 (O_2126,N_24837,N_21542);
xor UO_2127 (O_2127,N_24635,N_24542);
or UO_2128 (O_2128,N_20657,N_24229);
xnor UO_2129 (O_2129,N_24494,N_20788);
or UO_2130 (O_2130,N_20532,N_20463);
and UO_2131 (O_2131,N_23153,N_23308);
and UO_2132 (O_2132,N_20618,N_20276);
and UO_2133 (O_2133,N_20060,N_23641);
and UO_2134 (O_2134,N_20561,N_21099);
nand UO_2135 (O_2135,N_24922,N_23361);
or UO_2136 (O_2136,N_23764,N_20116);
or UO_2137 (O_2137,N_23527,N_21389);
nand UO_2138 (O_2138,N_24871,N_24589);
and UO_2139 (O_2139,N_22033,N_21347);
nor UO_2140 (O_2140,N_20984,N_20204);
nand UO_2141 (O_2141,N_24186,N_23812);
xor UO_2142 (O_2142,N_24857,N_23541);
nor UO_2143 (O_2143,N_20435,N_21755);
nand UO_2144 (O_2144,N_22708,N_20112);
and UO_2145 (O_2145,N_24162,N_22102);
xor UO_2146 (O_2146,N_24032,N_21170);
nor UO_2147 (O_2147,N_24094,N_22926);
xor UO_2148 (O_2148,N_22960,N_23158);
xor UO_2149 (O_2149,N_22622,N_20174);
nor UO_2150 (O_2150,N_20017,N_21706);
xor UO_2151 (O_2151,N_22267,N_24681);
nand UO_2152 (O_2152,N_24974,N_21455);
and UO_2153 (O_2153,N_24285,N_24730);
and UO_2154 (O_2154,N_22066,N_21597);
nor UO_2155 (O_2155,N_21908,N_20607);
nor UO_2156 (O_2156,N_24275,N_21403);
nand UO_2157 (O_2157,N_22838,N_24584);
or UO_2158 (O_2158,N_22387,N_24082);
and UO_2159 (O_2159,N_22354,N_20911);
nand UO_2160 (O_2160,N_21659,N_20928);
or UO_2161 (O_2161,N_24397,N_23504);
nor UO_2162 (O_2162,N_22455,N_24835);
nand UO_2163 (O_2163,N_24666,N_23031);
nand UO_2164 (O_2164,N_22242,N_20428);
and UO_2165 (O_2165,N_23752,N_20445);
nor UO_2166 (O_2166,N_22205,N_23824);
xnor UO_2167 (O_2167,N_20178,N_23894);
and UO_2168 (O_2168,N_23456,N_22165);
and UO_2169 (O_2169,N_23451,N_23160);
or UO_2170 (O_2170,N_23195,N_22459);
nand UO_2171 (O_2171,N_22947,N_20747);
and UO_2172 (O_2172,N_21396,N_20297);
or UO_2173 (O_2173,N_22005,N_21166);
nor UO_2174 (O_2174,N_20541,N_21665);
xor UO_2175 (O_2175,N_20442,N_24711);
nand UO_2176 (O_2176,N_24957,N_23875);
xor UO_2177 (O_2177,N_22691,N_22647);
and UO_2178 (O_2178,N_22880,N_23431);
and UO_2179 (O_2179,N_24240,N_24683);
or UO_2180 (O_2180,N_23152,N_22644);
and UO_2181 (O_2181,N_23162,N_23295);
nor UO_2182 (O_2182,N_24846,N_22163);
or UO_2183 (O_2183,N_21226,N_22657);
or UO_2184 (O_2184,N_23807,N_22779);
xnor UO_2185 (O_2185,N_24221,N_24553);
nand UO_2186 (O_2186,N_21405,N_22169);
nor UO_2187 (O_2187,N_21250,N_22876);
nor UO_2188 (O_2188,N_22898,N_21372);
nor UO_2189 (O_2189,N_20137,N_22321);
xor UO_2190 (O_2190,N_23776,N_20142);
nor UO_2191 (O_2191,N_21556,N_22040);
or UO_2192 (O_2192,N_20374,N_20313);
xnor UO_2193 (O_2193,N_23680,N_20609);
nor UO_2194 (O_2194,N_23706,N_22112);
or UO_2195 (O_2195,N_23374,N_22871);
xor UO_2196 (O_2196,N_22703,N_22519);
xnor UO_2197 (O_2197,N_21888,N_21998);
xor UO_2198 (O_2198,N_23072,N_21808);
and UO_2199 (O_2199,N_21315,N_21423);
nand UO_2200 (O_2200,N_23233,N_23629);
nand UO_2201 (O_2201,N_24506,N_24007);
and UO_2202 (O_2202,N_22755,N_24091);
nand UO_2203 (O_2203,N_22220,N_24319);
xnor UO_2204 (O_2204,N_23297,N_23301);
xnor UO_2205 (O_2205,N_24482,N_22811);
nor UO_2206 (O_2206,N_20912,N_23202);
nor UO_2207 (O_2207,N_23454,N_20635);
nand UO_2208 (O_2208,N_20003,N_23262);
nor UO_2209 (O_2209,N_20590,N_21720);
xor UO_2210 (O_2210,N_24117,N_20879);
or UO_2211 (O_2211,N_21896,N_24325);
xnor UO_2212 (O_2212,N_24576,N_22704);
nand UO_2213 (O_2213,N_22295,N_24762);
nand UO_2214 (O_2214,N_23011,N_20519);
xnor UO_2215 (O_2215,N_24101,N_24121);
or UO_2216 (O_2216,N_21799,N_21186);
and UO_2217 (O_2217,N_24614,N_23563);
nand UO_2218 (O_2218,N_24024,N_24958);
nor UO_2219 (O_2219,N_22592,N_20583);
nand UO_2220 (O_2220,N_22269,N_20059);
or UO_2221 (O_2221,N_22282,N_20554);
or UO_2222 (O_2222,N_23555,N_22451);
and UO_2223 (O_2223,N_22797,N_24605);
nor UO_2224 (O_2224,N_23380,N_24840);
or UO_2225 (O_2225,N_21265,N_22472);
and UO_2226 (O_2226,N_22478,N_22670);
or UO_2227 (O_2227,N_22773,N_20227);
or UO_2228 (O_2228,N_20310,N_21136);
nor UO_2229 (O_2229,N_24099,N_21146);
nor UO_2230 (O_2230,N_21636,N_23505);
nor UO_2231 (O_2231,N_23985,N_24915);
or UO_2232 (O_2232,N_20803,N_23463);
nand UO_2233 (O_2233,N_24355,N_23287);
xor UO_2234 (O_2234,N_22894,N_22145);
and UO_2235 (O_2235,N_22449,N_24909);
nand UO_2236 (O_2236,N_23862,N_23650);
xor UO_2237 (O_2237,N_22346,N_21224);
nand UO_2238 (O_2238,N_22167,N_23387);
or UO_2239 (O_2239,N_22843,N_24774);
nand UO_2240 (O_2240,N_21344,N_21409);
nor UO_2241 (O_2241,N_22579,N_23274);
nand UO_2242 (O_2242,N_24956,N_20097);
and UO_2243 (O_2243,N_22581,N_22411);
or UO_2244 (O_2244,N_22712,N_22237);
and UO_2245 (O_2245,N_22052,N_21374);
nor UO_2246 (O_2246,N_20385,N_22971);
or UO_2247 (O_2247,N_22352,N_23231);
nor UO_2248 (O_2248,N_24156,N_23637);
xor UO_2249 (O_2249,N_22534,N_20211);
and UO_2250 (O_2250,N_21697,N_23415);
xor UO_2251 (O_2251,N_23559,N_22146);
nand UO_2252 (O_2252,N_22343,N_22615);
and UO_2253 (O_2253,N_22695,N_20004);
or UO_2254 (O_2254,N_22126,N_23120);
and UO_2255 (O_2255,N_21148,N_21762);
and UO_2256 (O_2256,N_23469,N_24146);
nand UO_2257 (O_2257,N_24559,N_21647);
nor UO_2258 (O_2258,N_24852,N_23907);
xnor UO_2259 (O_2259,N_22109,N_23439);
xnor UO_2260 (O_2260,N_23357,N_21642);
nor UO_2261 (O_2261,N_23438,N_21430);
nor UO_2262 (O_2262,N_23276,N_22624);
nor UO_2263 (O_2263,N_22603,N_23768);
nand UO_2264 (O_2264,N_20950,N_22487);
nand UO_2265 (O_2265,N_24021,N_20938);
xnor UO_2266 (O_2266,N_20973,N_22471);
and UO_2267 (O_2267,N_21410,N_22725);
or UO_2268 (O_2268,N_20420,N_23059);
xnor UO_2269 (O_2269,N_24828,N_24296);
nand UO_2270 (O_2270,N_20000,N_21064);
or UO_2271 (O_2271,N_22429,N_21416);
nand UO_2272 (O_2272,N_23549,N_21198);
or UO_2273 (O_2273,N_22800,N_22508);
or UO_2274 (O_2274,N_21337,N_22529);
nand UO_2275 (O_2275,N_21834,N_24332);
xor UO_2276 (O_2276,N_21569,N_20469);
xor UO_2277 (O_2277,N_20065,N_20339);
xnor UO_2278 (O_2278,N_24582,N_22230);
nand UO_2279 (O_2279,N_21329,N_23790);
nand UO_2280 (O_2280,N_20155,N_23830);
xnor UO_2281 (O_2281,N_24611,N_21797);
or UO_2282 (O_2282,N_24919,N_23890);
nor UO_2283 (O_2283,N_22589,N_23982);
or UO_2284 (O_2284,N_20773,N_21461);
xnor UO_2285 (O_2285,N_20931,N_24531);
nor UO_2286 (O_2286,N_22331,N_22255);
xnor UO_2287 (O_2287,N_20548,N_24860);
and UO_2288 (O_2288,N_22096,N_24480);
and UO_2289 (O_2289,N_22048,N_23725);
or UO_2290 (O_2290,N_20236,N_24096);
or UO_2291 (O_2291,N_23218,N_23319);
nor UO_2292 (O_2292,N_20373,N_22527);
or UO_2293 (O_2293,N_23674,N_22435);
xor UO_2294 (O_2294,N_24948,N_24315);
and UO_2295 (O_2295,N_23578,N_23592);
or UO_2296 (O_2296,N_21153,N_21674);
nor UO_2297 (O_2297,N_22888,N_22292);
or UO_2298 (O_2298,N_21201,N_24563);
and UO_2299 (O_2299,N_20551,N_24323);
and UO_2300 (O_2300,N_23732,N_22608);
xnor UO_2301 (O_2301,N_24085,N_24464);
and UO_2302 (O_2302,N_24878,N_23368);
nand UO_2303 (O_2303,N_23983,N_21441);
nand UO_2304 (O_2304,N_24727,N_21022);
nor UO_2305 (O_2305,N_22088,N_24953);
or UO_2306 (O_2306,N_22301,N_24224);
nand UO_2307 (O_2307,N_22240,N_20176);
xor UO_2308 (O_2308,N_22041,N_21466);
and UO_2309 (O_2309,N_24044,N_22226);
and UO_2310 (O_2310,N_20424,N_24441);
or UO_2311 (O_2311,N_21754,N_24334);
nand UO_2312 (O_2312,N_22964,N_20025);
xor UO_2313 (O_2313,N_20451,N_22536);
nand UO_2314 (O_2314,N_22569,N_21677);
or UO_2315 (O_2315,N_23710,N_23140);
nor UO_2316 (O_2316,N_22776,N_20856);
and UO_2317 (O_2317,N_22395,N_23184);
or UO_2318 (O_2318,N_20081,N_21603);
or UO_2319 (O_2319,N_20899,N_21251);
nand UO_2320 (O_2320,N_24131,N_23653);
or UO_2321 (O_2321,N_20626,N_22075);
and UO_2322 (O_2322,N_23335,N_23903);
or UO_2323 (O_2323,N_23071,N_21462);
and UO_2324 (O_2324,N_20957,N_20702);
xor UO_2325 (O_2325,N_21140,N_22866);
or UO_2326 (O_2326,N_20398,N_20887);
nand UO_2327 (O_2327,N_22826,N_23667);
and UO_2328 (O_2328,N_20202,N_24005);
nor UO_2329 (O_2329,N_23346,N_20863);
xor UO_2330 (O_2330,N_21039,N_21975);
or UO_2331 (O_2331,N_23284,N_24892);
and UO_2332 (O_2332,N_21800,N_23340);
nor UO_2333 (O_2333,N_22160,N_23647);
or UO_2334 (O_2334,N_21431,N_22086);
or UO_2335 (O_2335,N_20160,N_24026);
nor UO_2336 (O_2336,N_20366,N_20759);
nand UO_2337 (O_2337,N_23571,N_20780);
nor UO_2338 (O_2338,N_23937,N_24682);
and UO_2339 (O_2339,N_23550,N_23663);
and UO_2340 (O_2340,N_20206,N_22135);
or UO_2341 (O_2341,N_21247,N_21036);
or UO_2342 (O_2342,N_21997,N_20884);
nor UO_2343 (O_2343,N_21393,N_20871);
nor UO_2344 (O_2344,N_22361,N_20643);
or UO_2345 (O_2345,N_23834,N_24080);
nor UO_2346 (O_2346,N_20415,N_21835);
and UO_2347 (O_2347,N_20018,N_24539);
nor UO_2348 (O_2348,N_24120,N_22975);
xor UO_2349 (O_2349,N_21764,N_21082);
nor UO_2350 (O_2350,N_20809,N_24386);
nand UO_2351 (O_2351,N_23727,N_24702);
or UO_2352 (O_2352,N_21819,N_21843);
nand UO_2353 (O_2353,N_23607,N_20718);
and UO_2354 (O_2354,N_24522,N_22994);
or UO_2355 (O_2355,N_21620,N_23480);
or UO_2356 (O_2356,N_21465,N_22763);
xor UO_2357 (O_2357,N_21714,N_23372);
or UO_2358 (O_2358,N_20229,N_21930);
xor UO_2359 (O_2359,N_23932,N_22463);
nand UO_2360 (O_2360,N_23420,N_22046);
and UO_2361 (O_2361,N_24166,N_20460);
nand UO_2362 (O_2362,N_24932,N_22931);
or UO_2363 (O_2363,N_20878,N_20041);
nor UO_2364 (O_2364,N_21847,N_20240);
nand UO_2365 (O_2365,N_22208,N_24207);
and UO_2366 (O_2366,N_24777,N_20951);
and UO_2367 (O_2367,N_23542,N_22847);
and UO_2368 (O_2368,N_23240,N_20149);
or UO_2369 (O_2369,N_22639,N_24401);
and UO_2370 (O_2370,N_24854,N_21804);
xor UO_2371 (O_2371,N_20269,N_20096);
nand UO_2372 (O_2372,N_21658,N_20099);
nor UO_2373 (O_2373,N_23928,N_22788);
or UO_2374 (O_2374,N_24782,N_21824);
or UO_2375 (O_2375,N_24849,N_21070);
or UO_2376 (O_2376,N_22707,N_23270);
xor UO_2377 (O_2377,N_22640,N_21000);
and UO_2378 (O_2378,N_20644,N_22189);
or UO_2379 (O_2379,N_21451,N_20126);
nand UO_2380 (O_2380,N_24820,N_24215);
nor UO_2381 (O_2381,N_22315,N_24421);
or UO_2382 (O_2382,N_24502,N_22979);
or UO_2383 (O_2383,N_22585,N_23522);
or UO_2384 (O_2384,N_21369,N_21874);
nor UO_2385 (O_2385,N_23651,N_21973);
and UO_2386 (O_2386,N_24510,N_23099);
nor UO_2387 (O_2387,N_22513,N_24928);
or UO_2388 (O_2388,N_23635,N_24273);
xor UO_2389 (O_2389,N_20196,N_23664);
xor UO_2390 (O_2390,N_24617,N_21206);
xnor UO_2391 (O_2391,N_20696,N_24185);
nor UO_2392 (O_2392,N_22789,N_23881);
or UO_2393 (O_2393,N_23108,N_20267);
nor UO_2394 (O_2394,N_23800,N_20735);
or UO_2395 (O_2395,N_20766,N_20623);
or UO_2396 (O_2396,N_21694,N_22412);
nand UO_2397 (O_2397,N_20778,N_24757);
xnor UO_2398 (O_2398,N_23666,N_20113);
nand UO_2399 (O_2399,N_24604,N_23593);
xor UO_2400 (O_2400,N_22509,N_24543);
nand UO_2401 (O_2401,N_23396,N_22054);
nor UO_2402 (O_2402,N_24128,N_20890);
nor UO_2403 (O_2403,N_22807,N_23564);
nor UO_2404 (O_2404,N_23579,N_21999);
nand UO_2405 (O_2405,N_24736,N_24533);
xor UO_2406 (O_2406,N_21735,N_22439);
nor UO_2407 (O_2407,N_21444,N_22613);
nor UO_2408 (O_2408,N_23487,N_21525);
nand UO_2409 (O_2409,N_24371,N_21638);
xnor UO_2410 (O_2410,N_24519,N_24219);
and UO_2411 (O_2411,N_23201,N_20247);
nand UO_2412 (O_2412,N_21059,N_20439);
and UO_2413 (O_2413,N_24843,N_20993);
or UO_2414 (O_2414,N_22279,N_23251);
or UO_2415 (O_2415,N_22658,N_23796);
nand UO_2416 (O_2416,N_22340,N_21644);
and UO_2417 (O_2417,N_24817,N_23685);
nand UO_2418 (O_2418,N_21384,N_23931);
or UO_2419 (O_2419,N_23208,N_21491);
and UO_2420 (O_2420,N_23267,N_22692);
nand UO_2421 (O_2421,N_20254,N_20447);
xor UO_2422 (O_2422,N_23626,N_24236);
nor UO_2423 (O_2423,N_24104,N_24231);
or UO_2424 (O_2424,N_24608,N_21027);
xnor UO_2425 (O_2425,N_24076,N_21689);
or UO_2426 (O_2426,N_23660,N_22631);
or UO_2427 (O_2427,N_22408,N_20919);
or UO_2428 (O_2428,N_21690,N_24706);
xor UO_2429 (O_2429,N_23144,N_21813);
xor UO_2430 (O_2430,N_20597,N_20785);
xnor UO_2431 (O_2431,N_24416,N_20713);
xnor UO_2432 (O_2432,N_21501,N_20945);
or UO_2433 (O_2433,N_22732,N_24806);
nor UO_2434 (O_2434,N_24992,N_24191);
and UO_2435 (O_2435,N_23025,N_23622);
xor UO_2436 (O_2436,N_21820,N_22073);
nand UO_2437 (O_2437,N_23887,N_21050);
and UO_2438 (O_2438,N_20999,N_21025);
xor UO_2439 (O_2439,N_23766,N_20488);
nor UO_2440 (O_2440,N_21792,N_20034);
xor UO_2441 (O_2441,N_20101,N_20470);
xnor UO_2442 (O_2442,N_23547,N_21387);
or UO_2443 (O_2443,N_20333,N_20591);
or UO_2444 (O_2444,N_20022,N_22702);
and UO_2445 (O_2445,N_20642,N_21429);
nand UO_2446 (O_2446,N_23817,N_24691);
nand UO_2447 (O_2447,N_21195,N_21521);
nand UO_2448 (O_2448,N_23948,N_20654);
nor UO_2449 (O_2449,N_21992,N_20150);
xnor UO_2450 (O_2450,N_21914,N_22214);
nand UO_2451 (O_2451,N_21045,N_24638);
nor UO_2452 (O_2452,N_23443,N_23904);
nor UO_2453 (O_2453,N_24896,N_22718);
xnor UO_2454 (O_2454,N_20997,N_24087);
nor UO_2455 (O_2455,N_22442,N_22362);
or UO_2456 (O_2456,N_20556,N_23929);
or UO_2457 (O_2457,N_23911,N_23484);
nand UO_2458 (O_2458,N_21117,N_22335);
nor UO_2459 (O_2459,N_24002,N_23672);
xnor UO_2460 (O_2460,N_24688,N_20621);
and UO_2461 (O_2461,N_21292,N_20011);
nor UO_2462 (O_2462,N_21003,N_24136);
nor UO_2463 (O_2463,N_20841,N_21740);
nor UO_2464 (O_2464,N_23530,N_20465);
nor UO_2465 (O_2465,N_22935,N_21280);
and UO_2466 (O_2466,N_20219,N_22144);
or UO_2467 (O_2467,N_24232,N_20031);
and UO_2468 (O_2468,N_22573,N_21041);
and UO_2469 (O_2469,N_21875,N_23046);
and UO_2470 (O_2470,N_22091,N_23044);
or UO_2471 (O_2471,N_24842,N_23029);
and UO_2472 (O_2472,N_20068,N_22643);
and UO_2473 (O_2473,N_23258,N_23004);
xor UO_2474 (O_2474,N_20264,N_21942);
nand UO_2475 (O_2475,N_21398,N_21940);
and UO_2476 (O_2476,N_23391,N_20772);
nor UO_2477 (O_2477,N_20453,N_20262);
nor UO_2478 (O_2478,N_20922,N_20207);
and UO_2479 (O_2479,N_20808,N_24040);
nand UO_2480 (O_2480,N_22426,N_23447);
and UO_2481 (O_2481,N_20810,N_22905);
or UO_2482 (O_2482,N_23858,N_21308);
and UO_2483 (O_2483,N_21018,N_21182);
xor UO_2484 (O_2484,N_21298,N_24640);
xor UO_2485 (O_2485,N_22499,N_24766);
or UO_2486 (O_2486,N_23175,N_23061);
or UO_2487 (O_2487,N_20682,N_22461);
nor UO_2488 (O_2488,N_24685,N_21437);
xor UO_2489 (O_2489,N_23736,N_24383);
xnor UO_2490 (O_2490,N_23944,N_24160);
and UO_2491 (O_2491,N_21736,N_20230);
nand UO_2492 (O_2492,N_24272,N_22225);
and UO_2493 (O_2493,N_20733,N_22263);
and UO_2494 (O_2494,N_20724,N_24410);
nand UO_2495 (O_2495,N_22808,N_21980);
or UO_2496 (O_2496,N_24515,N_21115);
nor UO_2497 (O_2497,N_23780,N_24372);
xor UO_2498 (O_2498,N_24508,N_20292);
nor UO_2499 (O_2499,N_20188,N_21450);
and UO_2500 (O_2500,N_21125,N_23277);
nor UO_2501 (O_2501,N_24808,N_23900);
or UO_2502 (O_2502,N_24342,N_21408);
xnor UO_2503 (O_2503,N_23048,N_23624);
xnor UO_2504 (O_2504,N_23800,N_22028);
nor UO_2505 (O_2505,N_20878,N_23758);
and UO_2506 (O_2506,N_23674,N_23441);
nor UO_2507 (O_2507,N_20064,N_22169);
or UO_2508 (O_2508,N_23068,N_20886);
and UO_2509 (O_2509,N_22380,N_23662);
nor UO_2510 (O_2510,N_20688,N_23043);
xnor UO_2511 (O_2511,N_22346,N_24591);
nor UO_2512 (O_2512,N_20129,N_20626);
nor UO_2513 (O_2513,N_24250,N_23422);
nand UO_2514 (O_2514,N_20930,N_20453);
or UO_2515 (O_2515,N_20571,N_23600);
and UO_2516 (O_2516,N_21528,N_20447);
nand UO_2517 (O_2517,N_22352,N_23712);
xor UO_2518 (O_2518,N_24993,N_24572);
xor UO_2519 (O_2519,N_22528,N_22951);
nand UO_2520 (O_2520,N_24059,N_20776);
nand UO_2521 (O_2521,N_23712,N_22973);
nor UO_2522 (O_2522,N_23280,N_24625);
xor UO_2523 (O_2523,N_22066,N_22097);
xnor UO_2524 (O_2524,N_20479,N_20153);
and UO_2525 (O_2525,N_20674,N_20821);
nor UO_2526 (O_2526,N_23551,N_23354);
and UO_2527 (O_2527,N_21961,N_23992);
nor UO_2528 (O_2528,N_20514,N_23285);
xnor UO_2529 (O_2529,N_20379,N_23988);
or UO_2530 (O_2530,N_24991,N_20945);
or UO_2531 (O_2531,N_22612,N_20540);
xnor UO_2532 (O_2532,N_20959,N_22812);
and UO_2533 (O_2533,N_24473,N_21841);
nand UO_2534 (O_2534,N_20164,N_23851);
nor UO_2535 (O_2535,N_23682,N_22121);
and UO_2536 (O_2536,N_21581,N_23899);
and UO_2537 (O_2537,N_23453,N_22747);
nand UO_2538 (O_2538,N_23775,N_22993);
nand UO_2539 (O_2539,N_20803,N_23401);
nand UO_2540 (O_2540,N_24553,N_20979);
and UO_2541 (O_2541,N_23961,N_23561);
xnor UO_2542 (O_2542,N_24537,N_22951);
nor UO_2543 (O_2543,N_22314,N_20173);
nor UO_2544 (O_2544,N_24117,N_24069);
or UO_2545 (O_2545,N_24846,N_21585);
and UO_2546 (O_2546,N_21572,N_23828);
nor UO_2547 (O_2547,N_20432,N_23856);
nor UO_2548 (O_2548,N_22668,N_21648);
or UO_2549 (O_2549,N_21850,N_23975);
or UO_2550 (O_2550,N_22795,N_23147);
nor UO_2551 (O_2551,N_21733,N_21641);
nor UO_2552 (O_2552,N_21892,N_24685);
nor UO_2553 (O_2553,N_20773,N_20784);
nand UO_2554 (O_2554,N_24122,N_20741);
xnor UO_2555 (O_2555,N_23978,N_20966);
xnor UO_2556 (O_2556,N_24232,N_21242);
nand UO_2557 (O_2557,N_23455,N_21965);
xor UO_2558 (O_2558,N_23488,N_22708);
and UO_2559 (O_2559,N_24221,N_23145);
nand UO_2560 (O_2560,N_23653,N_20019);
nand UO_2561 (O_2561,N_21927,N_22949);
nand UO_2562 (O_2562,N_21103,N_21330);
nand UO_2563 (O_2563,N_23635,N_20181);
nand UO_2564 (O_2564,N_22438,N_23754);
nand UO_2565 (O_2565,N_22781,N_21311);
nor UO_2566 (O_2566,N_22884,N_22035);
xor UO_2567 (O_2567,N_20370,N_22883);
or UO_2568 (O_2568,N_20526,N_24968);
nor UO_2569 (O_2569,N_24444,N_20748);
nor UO_2570 (O_2570,N_24861,N_20788);
and UO_2571 (O_2571,N_21002,N_21094);
nor UO_2572 (O_2572,N_24860,N_22793);
or UO_2573 (O_2573,N_23413,N_20196);
nand UO_2574 (O_2574,N_23644,N_21441);
nand UO_2575 (O_2575,N_24910,N_21038);
nor UO_2576 (O_2576,N_22757,N_22481);
xor UO_2577 (O_2577,N_23406,N_21027);
and UO_2578 (O_2578,N_20923,N_23920);
xnor UO_2579 (O_2579,N_20075,N_24753);
or UO_2580 (O_2580,N_20690,N_20272);
nand UO_2581 (O_2581,N_21182,N_23871);
xnor UO_2582 (O_2582,N_22905,N_21204);
or UO_2583 (O_2583,N_23637,N_21528);
and UO_2584 (O_2584,N_21913,N_23741);
nand UO_2585 (O_2585,N_20469,N_21615);
or UO_2586 (O_2586,N_22882,N_24509);
nand UO_2587 (O_2587,N_24018,N_24876);
xor UO_2588 (O_2588,N_22208,N_24390);
xor UO_2589 (O_2589,N_21005,N_23949);
nor UO_2590 (O_2590,N_21073,N_23541);
xor UO_2591 (O_2591,N_24533,N_22943);
xor UO_2592 (O_2592,N_22717,N_23253);
xnor UO_2593 (O_2593,N_20624,N_21862);
nand UO_2594 (O_2594,N_21082,N_20649);
or UO_2595 (O_2595,N_24237,N_20424);
nand UO_2596 (O_2596,N_20215,N_22863);
or UO_2597 (O_2597,N_21523,N_21740);
nand UO_2598 (O_2598,N_21333,N_22294);
xnor UO_2599 (O_2599,N_23056,N_21430);
xnor UO_2600 (O_2600,N_20299,N_22117);
nor UO_2601 (O_2601,N_21040,N_24102);
or UO_2602 (O_2602,N_21816,N_20392);
nor UO_2603 (O_2603,N_22701,N_23045);
xnor UO_2604 (O_2604,N_20673,N_22498);
nor UO_2605 (O_2605,N_20124,N_20638);
and UO_2606 (O_2606,N_24632,N_20860);
and UO_2607 (O_2607,N_21462,N_20928);
and UO_2608 (O_2608,N_24580,N_21748);
nand UO_2609 (O_2609,N_22406,N_24886);
xor UO_2610 (O_2610,N_24631,N_21950);
nor UO_2611 (O_2611,N_22118,N_22079);
nand UO_2612 (O_2612,N_21452,N_24177);
and UO_2613 (O_2613,N_20704,N_23688);
or UO_2614 (O_2614,N_22376,N_24917);
or UO_2615 (O_2615,N_22297,N_20186);
nor UO_2616 (O_2616,N_22048,N_23890);
nor UO_2617 (O_2617,N_23628,N_23803);
nand UO_2618 (O_2618,N_20142,N_24931);
or UO_2619 (O_2619,N_21452,N_21442);
and UO_2620 (O_2620,N_21244,N_21509);
xor UO_2621 (O_2621,N_23694,N_21392);
xor UO_2622 (O_2622,N_23740,N_20312);
or UO_2623 (O_2623,N_23658,N_20008);
nand UO_2624 (O_2624,N_21404,N_20926);
nand UO_2625 (O_2625,N_22571,N_20086);
nor UO_2626 (O_2626,N_24200,N_24418);
or UO_2627 (O_2627,N_21109,N_21438);
xnor UO_2628 (O_2628,N_20732,N_22161);
or UO_2629 (O_2629,N_23721,N_20694);
and UO_2630 (O_2630,N_24812,N_23846);
or UO_2631 (O_2631,N_21744,N_24541);
xnor UO_2632 (O_2632,N_24965,N_21638);
and UO_2633 (O_2633,N_21233,N_23702);
nand UO_2634 (O_2634,N_21484,N_24661);
nand UO_2635 (O_2635,N_24929,N_22299);
and UO_2636 (O_2636,N_21868,N_20632);
xor UO_2637 (O_2637,N_23041,N_22233);
or UO_2638 (O_2638,N_20462,N_20132);
and UO_2639 (O_2639,N_20621,N_20754);
or UO_2640 (O_2640,N_22535,N_22349);
xnor UO_2641 (O_2641,N_22961,N_24246);
nor UO_2642 (O_2642,N_21475,N_21304);
and UO_2643 (O_2643,N_23427,N_20940);
and UO_2644 (O_2644,N_24651,N_20637);
and UO_2645 (O_2645,N_23758,N_20429);
or UO_2646 (O_2646,N_24486,N_21751);
and UO_2647 (O_2647,N_24526,N_24267);
nand UO_2648 (O_2648,N_21215,N_23463);
or UO_2649 (O_2649,N_20180,N_24498);
and UO_2650 (O_2650,N_20603,N_20901);
nor UO_2651 (O_2651,N_20933,N_20988);
xor UO_2652 (O_2652,N_24018,N_23444);
and UO_2653 (O_2653,N_22962,N_21582);
xnor UO_2654 (O_2654,N_23851,N_23982);
nand UO_2655 (O_2655,N_22246,N_24871);
nor UO_2656 (O_2656,N_22704,N_22874);
or UO_2657 (O_2657,N_24079,N_23055);
and UO_2658 (O_2658,N_20525,N_21824);
or UO_2659 (O_2659,N_23882,N_23159);
xnor UO_2660 (O_2660,N_21942,N_24264);
and UO_2661 (O_2661,N_22619,N_22840);
or UO_2662 (O_2662,N_24891,N_24016);
nor UO_2663 (O_2663,N_22091,N_21685);
xor UO_2664 (O_2664,N_23052,N_22749);
nand UO_2665 (O_2665,N_22470,N_22941);
xor UO_2666 (O_2666,N_24016,N_20603);
nand UO_2667 (O_2667,N_20167,N_22617);
and UO_2668 (O_2668,N_22526,N_22337);
nand UO_2669 (O_2669,N_23407,N_23384);
nand UO_2670 (O_2670,N_21476,N_22010);
nand UO_2671 (O_2671,N_21419,N_23284);
or UO_2672 (O_2672,N_24742,N_21271);
xor UO_2673 (O_2673,N_21563,N_23550);
nor UO_2674 (O_2674,N_23069,N_20636);
and UO_2675 (O_2675,N_22465,N_22954);
nor UO_2676 (O_2676,N_22481,N_24936);
and UO_2677 (O_2677,N_22535,N_21942);
nand UO_2678 (O_2678,N_22803,N_24349);
xor UO_2679 (O_2679,N_20893,N_24928);
xor UO_2680 (O_2680,N_24302,N_23162);
xor UO_2681 (O_2681,N_22789,N_22842);
or UO_2682 (O_2682,N_24675,N_24631);
nand UO_2683 (O_2683,N_20999,N_20172);
and UO_2684 (O_2684,N_21374,N_20165);
or UO_2685 (O_2685,N_24430,N_23722);
nand UO_2686 (O_2686,N_23809,N_24055);
nand UO_2687 (O_2687,N_21723,N_21965);
nor UO_2688 (O_2688,N_21027,N_24892);
xnor UO_2689 (O_2689,N_23873,N_23225);
xor UO_2690 (O_2690,N_22934,N_24630);
nor UO_2691 (O_2691,N_20868,N_22521);
nor UO_2692 (O_2692,N_20477,N_24600);
nand UO_2693 (O_2693,N_20990,N_23695);
nor UO_2694 (O_2694,N_23974,N_24829);
or UO_2695 (O_2695,N_24260,N_20177);
and UO_2696 (O_2696,N_23674,N_20225);
xor UO_2697 (O_2697,N_21237,N_20287);
nand UO_2698 (O_2698,N_21856,N_21567);
and UO_2699 (O_2699,N_20425,N_21715);
nor UO_2700 (O_2700,N_23765,N_22673);
or UO_2701 (O_2701,N_22794,N_23837);
and UO_2702 (O_2702,N_22703,N_23903);
and UO_2703 (O_2703,N_24038,N_22166);
and UO_2704 (O_2704,N_20522,N_22154);
and UO_2705 (O_2705,N_21400,N_20835);
nand UO_2706 (O_2706,N_24159,N_21629);
or UO_2707 (O_2707,N_23093,N_22077);
xor UO_2708 (O_2708,N_20382,N_23530);
and UO_2709 (O_2709,N_23064,N_24744);
and UO_2710 (O_2710,N_20681,N_24010);
nand UO_2711 (O_2711,N_20330,N_21735);
and UO_2712 (O_2712,N_20484,N_20893);
nor UO_2713 (O_2713,N_22381,N_20523);
or UO_2714 (O_2714,N_21634,N_20193);
or UO_2715 (O_2715,N_20271,N_22654);
xnor UO_2716 (O_2716,N_21995,N_21002);
nand UO_2717 (O_2717,N_23508,N_21484);
nor UO_2718 (O_2718,N_21089,N_24989);
nand UO_2719 (O_2719,N_24314,N_20336);
and UO_2720 (O_2720,N_20183,N_24395);
and UO_2721 (O_2721,N_23909,N_21746);
or UO_2722 (O_2722,N_21439,N_20131);
and UO_2723 (O_2723,N_24049,N_22865);
and UO_2724 (O_2724,N_22105,N_24714);
or UO_2725 (O_2725,N_24615,N_22974);
nor UO_2726 (O_2726,N_24344,N_22709);
nand UO_2727 (O_2727,N_20967,N_20440);
or UO_2728 (O_2728,N_24423,N_21716);
nand UO_2729 (O_2729,N_21852,N_20646);
xnor UO_2730 (O_2730,N_20704,N_22112);
or UO_2731 (O_2731,N_23306,N_24083);
nor UO_2732 (O_2732,N_21878,N_20031);
nor UO_2733 (O_2733,N_20588,N_23556);
nor UO_2734 (O_2734,N_21840,N_21219);
or UO_2735 (O_2735,N_22325,N_22754);
nor UO_2736 (O_2736,N_22155,N_23435);
and UO_2737 (O_2737,N_21217,N_21159);
nand UO_2738 (O_2738,N_20221,N_23405);
nand UO_2739 (O_2739,N_23703,N_20333);
nor UO_2740 (O_2740,N_23588,N_21524);
and UO_2741 (O_2741,N_24355,N_24329);
and UO_2742 (O_2742,N_21953,N_20716);
nand UO_2743 (O_2743,N_23680,N_24582);
xor UO_2744 (O_2744,N_20655,N_21743);
nor UO_2745 (O_2745,N_20548,N_23857);
or UO_2746 (O_2746,N_23410,N_22957);
and UO_2747 (O_2747,N_21152,N_23753);
nand UO_2748 (O_2748,N_21407,N_24679);
and UO_2749 (O_2749,N_24351,N_22995);
or UO_2750 (O_2750,N_20439,N_23172);
xor UO_2751 (O_2751,N_24932,N_21884);
nand UO_2752 (O_2752,N_24316,N_20680);
xor UO_2753 (O_2753,N_24948,N_22002);
or UO_2754 (O_2754,N_22547,N_22378);
nor UO_2755 (O_2755,N_22307,N_20066);
nor UO_2756 (O_2756,N_24371,N_24219);
nand UO_2757 (O_2757,N_20559,N_21097);
and UO_2758 (O_2758,N_22006,N_21193);
nand UO_2759 (O_2759,N_22485,N_22939);
and UO_2760 (O_2760,N_22681,N_22304);
nand UO_2761 (O_2761,N_24696,N_22922);
nand UO_2762 (O_2762,N_20575,N_23939);
nand UO_2763 (O_2763,N_21180,N_23642);
xnor UO_2764 (O_2764,N_20984,N_20830);
or UO_2765 (O_2765,N_24281,N_24557);
nand UO_2766 (O_2766,N_22202,N_23000);
nor UO_2767 (O_2767,N_20755,N_20381);
and UO_2768 (O_2768,N_22030,N_23347);
or UO_2769 (O_2769,N_24111,N_20053);
xnor UO_2770 (O_2770,N_20752,N_23412);
nor UO_2771 (O_2771,N_24572,N_21438);
and UO_2772 (O_2772,N_21577,N_23308);
and UO_2773 (O_2773,N_21421,N_23911);
nand UO_2774 (O_2774,N_24709,N_22265);
and UO_2775 (O_2775,N_23318,N_24857);
or UO_2776 (O_2776,N_22639,N_21143);
nor UO_2777 (O_2777,N_20150,N_21530);
nand UO_2778 (O_2778,N_21609,N_22649);
nor UO_2779 (O_2779,N_21938,N_21115);
nand UO_2780 (O_2780,N_20454,N_22653);
and UO_2781 (O_2781,N_21986,N_20539);
xor UO_2782 (O_2782,N_24810,N_24874);
nor UO_2783 (O_2783,N_23879,N_20003);
nor UO_2784 (O_2784,N_21824,N_23367);
nand UO_2785 (O_2785,N_22385,N_23373);
and UO_2786 (O_2786,N_22474,N_21029);
xor UO_2787 (O_2787,N_23757,N_20932);
xor UO_2788 (O_2788,N_21198,N_24772);
and UO_2789 (O_2789,N_20641,N_22989);
and UO_2790 (O_2790,N_20313,N_20195);
and UO_2791 (O_2791,N_22749,N_22515);
nor UO_2792 (O_2792,N_24284,N_23993);
xnor UO_2793 (O_2793,N_21991,N_24543);
nor UO_2794 (O_2794,N_21598,N_20800);
nand UO_2795 (O_2795,N_24614,N_20846);
or UO_2796 (O_2796,N_20583,N_23854);
and UO_2797 (O_2797,N_21228,N_21117);
nand UO_2798 (O_2798,N_24616,N_21882);
nand UO_2799 (O_2799,N_22182,N_24754);
and UO_2800 (O_2800,N_24954,N_23561);
nand UO_2801 (O_2801,N_24625,N_23667);
and UO_2802 (O_2802,N_23592,N_21532);
nor UO_2803 (O_2803,N_22343,N_22732);
xnor UO_2804 (O_2804,N_23017,N_21064);
nor UO_2805 (O_2805,N_20278,N_20151);
or UO_2806 (O_2806,N_22655,N_24859);
or UO_2807 (O_2807,N_24801,N_22744);
and UO_2808 (O_2808,N_22738,N_21310);
nand UO_2809 (O_2809,N_23888,N_22942);
or UO_2810 (O_2810,N_20217,N_24468);
nand UO_2811 (O_2811,N_20834,N_22922);
and UO_2812 (O_2812,N_23340,N_20387);
xnor UO_2813 (O_2813,N_22778,N_23361);
nand UO_2814 (O_2814,N_22471,N_23580);
xor UO_2815 (O_2815,N_20640,N_24656);
nand UO_2816 (O_2816,N_21255,N_22700);
nor UO_2817 (O_2817,N_22493,N_23984);
and UO_2818 (O_2818,N_22782,N_21960);
and UO_2819 (O_2819,N_22458,N_22707);
nor UO_2820 (O_2820,N_23906,N_21239);
or UO_2821 (O_2821,N_24321,N_21772);
or UO_2822 (O_2822,N_20878,N_20074);
or UO_2823 (O_2823,N_22422,N_22382);
nor UO_2824 (O_2824,N_23159,N_22029);
and UO_2825 (O_2825,N_20496,N_21393);
nor UO_2826 (O_2826,N_20968,N_23507);
nor UO_2827 (O_2827,N_20891,N_22722);
xnor UO_2828 (O_2828,N_20305,N_23809);
nand UO_2829 (O_2829,N_22589,N_20745);
nor UO_2830 (O_2830,N_20634,N_21843);
and UO_2831 (O_2831,N_23585,N_21181);
or UO_2832 (O_2832,N_23571,N_21323);
and UO_2833 (O_2833,N_20706,N_22654);
or UO_2834 (O_2834,N_22086,N_23252);
xor UO_2835 (O_2835,N_22182,N_24982);
or UO_2836 (O_2836,N_21163,N_24772);
and UO_2837 (O_2837,N_21661,N_24120);
xnor UO_2838 (O_2838,N_23246,N_21009);
or UO_2839 (O_2839,N_20397,N_21958);
xor UO_2840 (O_2840,N_21133,N_24404);
nor UO_2841 (O_2841,N_21999,N_21015);
or UO_2842 (O_2842,N_23000,N_23082);
nor UO_2843 (O_2843,N_23546,N_22272);
xor UO_2844 (O_2844,N_23985,N_21326);
nor UO_2845 (O_2845,N_20725,N_22111);
and UO_2846 (O_2846,N_21555,N_22375);
xor UO_2847 (O_2847,N_24151,N_20887);
and UO_2848 (O_2848,N_20237,N_23343);
and UO_2849 (O_2849,N_22180,N_22289);
and UO_2850 (O_2850,N_20547,N_24947);
xor UO_2851 (O_2851,N_24752,N_21068);
nor UO_2852 (O_2852,N_21285,N_21900);
nand UO_2853 (O_2853,N_20451,N_21495);
xnor UO_2854 (O_2854,N_23317,N_22099);
xor UO_2855 (O_2855,N_20573,N_23106);
or UO_2856 (O_2856,N_22066,N_20402);
xnor UO_2857 (O_2857,N_21505,N_22117);
and UO_2858 (O_2858,N_24091,N_22721);
xor UO_2859 (O_2859,N_24778,N_21868);
or UO_2860 (O_2860,N_23498,N_23403);
nor UO_2861 (O_2861,N_23099,N_24817);
xnor UO_2862 (O_2862,N_22252,N_23463);
nor UO_2863 (O_2863,N_23591,N_23677);
nand UO_2864 (O_2864,N_23687,N_22651);
nor UO_2865 (O_2865,N_23078,N_23823);
xor UO_2866 (O_2866,N_20706,N_21860);
and UO_2867 (O_2867,N_24278,N_22792);
nor UO_2868 (O_2868,N_23127,N_22804);
and UO_2869 (O_2869,N_24699,N_20188);
and UO_2870 (O_2870,N_21453,N_22742);
nand UO_2871 (O_2871,N_24800,N_24250);
nor UO_2872 (O_2872,N_24704,N_22452);
and UO_2873 (O_2873,N_20475,N_23678);
xor UO_2874 (O_2874,N_21233,N_24669);
and UO_2875 (O_2875,N_21466,N_22056);
and UO_2876 (O_2876,N_20459,N_23510);
nand UO_2877 (O_2877,N_20293,N_23736);
nand UO_2878 (O_2878,N_24101,N_24042);
and UO_2879 (O_2879,N_21978,N_20539);
and UO_2880 (O_2880,N_22930,N_21991);
xnor UO_2881 (O_2881,N_23391,N_20628);
xor UO_2882 (O_2882,N_23859,N_20512);
xor UO_2883 (O_2883,N_21556,N_24846);
nand UO_2884 (O_2884,N_23085,N_23120);
or UO_2885 (O_2885,N_21201,N_22021);
and UO_2886 (O_2886,N_22538,N_21563);
xnor UO_2887 (O_2887,N_22200,N_23507);
nor UO_2888 (O_2888,N_20688,N_20722);
and UO_2889 (O_2889,N_23712,N_21373);
and UO_2890 (O_2890,N_21264,N_21849);
nand UO_2891 (O_2891,N_21325,N_20554);
nor UO_2892 (O_2892,N_20723,N_20489);
nand UO_2893 (O_2893,N_21044,N_20440);
nor UO_2894 (O_2894,N_23336,N_24470);
xnor UO_2895 (O_2895,N_23556,N_22552);
nor UO_2896 (O_2896,N_20799,N_23868);
or UO_2897 (O_2897,N_21968,N_20195);
or UO_2898 (O_2898,N_20757,N_24735);
nand UO_2899 (O_2899,N_20756,N_23624);
nor UO_2900 (O_2900,N_22946,N_20939);
or UO_2901 (O_2901,N_21525,N_21800);
nor UO_2902 (O_2902,N_24107,N_20994);
xor UO_2903 (O_2903,N_23755,N_23587);
or UO_2904 (O_2904,N_21661,N_20353);
or UO_2905 (O_2905,N_23719,N_23399);
or UO_2906 (O_2906,N_20650,N_22491);
nand UO_2907 (O_2907,N_21955,N_24774);
or UO_2908 (O_2908,N_24545,N_24433);
nor UO_2909 (O_2909,N_24822,N_24362);
or UO_2910 (O_2910,N_23581,N_24125);
or UO_2911 (O_2911,N_23164,N_20253);
xnor UO_2912 (O_2912,N_22454,N_20074);
nand UO_2913 (O_2913,N_20696,N_21620);
and UO_2914 (O_2914,N_20249,N_22685);
or UO_2915 (O_2915,N_23266,N_23837);
and UO_2916 (O_2916,N_22606,N_22148);
nand UO_2917 (O_2917,N_22099,N_22518);
xnor UO_2918 (O_2918,N_24816,N_20658);
and UO_2919 (O_2919,N_21416,N_20841);
xnor UO_2920 (O_2920,N_24778,N_21400);
xor UO_2921 (O_2921,N_20883,N_22298);
and UO_2922 (O_2922,N_20718,N_24911);
and UO_2923 (O_2923,N_24447,N_22558);
nor UO_2924 (O_2924,N_23634,N_23480);
nor UO_2925 (O_2925,N_20546,N_23118);
nand UO_2926 (O_2926,N_21462,N_21607);
and UO_2927 (O_2927,N_20032,N_20570);
or UO_2928 (O_2928,N_23036,N_21409);
nand UO_2929 (O_2929,N_24646,N_22554);
xnor UO_2930 (O_2930,N_22330,N_23027);
or UO_2931 (O_2931,N_22261,N_22425);
and UO_2932 (O_2932,N_20103,N_21848);
or UO_2933 (O_2933,N_20205,N_24584);
nand UO_2934 (O_2934,N_24468,N_23021);
xnor UO_2935 (O_2935,N_23996,N_21202);
or UO_2936 (O_2936,N_23219,N_20092);
nand UO_2937 (O_2937,N_22137,N_20768);
or UO_2938 (O_2938,N_23463,N_20718);
nand UO_2939 (O_2939,N_20002,N_20931);
and UO_2940 (O_2940,N_24406,N_20793);
and UO_2941 (O_2941,N_20324,N_20381);
xnor UO_2942 (O_2942,N_20282,N_22912);
xor UO_2943 (O_2943,N_21884,N_23259);
nand UO_2944 (O_2944,N_22831,N_24080);
nor UO_2945 (O_2945,N_23791,N_24366);
nand UO_2946 (O_2946,N_24368,N_23801);
and UO_2947 (O_2947,N_23470,N_23875);
xor UO_2948 (O_2948,N_20599,N_23985);
or UO_2949 (O_2949,N_23483,N_23837);
nand UO_2950 (O_2950,N_22860,N_23811);
nor UO_2951 (O_2951,N_23388,N_24229);
or UO_2952 (O_2952,N_20665,N_22547);
and UO_2953 (O_2953,N_24842,N_21496);
xor UO_2954 (O_2954,N_24404,N_22890);
xor UO_2955 (O_2955,N_23575,N_20563);
and UO_2956 (O_2956,N_20768,N_24799);
or UO_2957 (O_2957,N_24452,N_22847);
nand UO_2958 (O_2958,N_20036,N_23665);
xnor UO_2959 (O_2959,N_20925,N_23011);
nor UO_2960 (O_2960,N_21745,N_23285);
nor UO_2961 (O_2961,N_22316,N_22166);
and UO_2962 (O_2962,N_24368,N_24536);
nand UO_2963 (O_2963,N_21554,N_23752);
or UO_2964 (O_2964,N_23848,N_20658);
nor UO_2965 (O_2965,N_22346,N_22164);
xnor UO_2966 (O_2966,N_21185,N_21206);
nand UO_2967 (O_2967,N_24961,N_22164);
nand UO_2968 (O_2968,N_20291,N_23153);
and UO_2969 (O_2969,N_20676,N_20493);
nand UO_2970 (O_2970,N_21959,N_21946);
xor UO_2971 (O_2971,N_23942,N_24177);
nand UO_2972 (O_2972,N_21609,N_20548);
xnor UO_2973 (O_2973,N_23311,N_22519);
and UO_2974 (O_2974,N_23492,N_23609);
nand UO_2975 (O_2975,N_20617,N_23148);
nand UO_2976 (O_2976,N_24130,N_22751);
or UO_2977 (O_2977,N_22328,N_20795);
or UO_2978 (O_2978,N_23404,N_20260);
xnor UO_2979 (O_2979,N_22568,N_21355);
or UO_2980 (O_2980,N_20547,N_23107);
xnor UO_2981 (O_2981,N_22143,N_23305);
nand UO_2982 (O_2982,N_22848,N_23350);
nand UO_2983 (O_2983,N_21141,N_23070);
or UO_2984 (O_2984,N_21085,N_24293);
nand UO_2985 (O_2985,N_20242,N_24834);
and UO_2986 (O_2986,N_22410,N_20581);
nand UO_2987 (O_2987,N_22484,N_20177);
or UO_2988 (O_2988,N_22437,N_24642);
nand UO_2989 (O_2989,N_24144,N_20315);
nand UO_2990 (O_2990,N_20825,N_24576);
xnor UO_2991 (O_2991,N_24103,N_23627);
or UO_2992 (O_2992,N_21860,N_22930);
and UO_2993 (O_2993,N_21924,N_23414);
xnor UO_2994 (O_2994,N_24638,N_22336);
and UO_2995 (O_2995,N_21670,N_21648);
and UO_2996 (O_2996,N_21635,N_24688);
nand UO_2997 (O_2997,N_23216,N_22910);
nor UO_2998 (O_2998,N_20559,N_20419);
and UO_2999 (O_2999,N_24868,N_24133);
endmodule