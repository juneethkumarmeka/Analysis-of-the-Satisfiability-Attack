module basic_1000_10000_1500_50_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_317,In_334);
nand U1 (N_1,In_46,In_790);
and U2 (N_2,In_596,In_810);
xnor U3 (N_3,In_595,In_30);
nor U4 (N_4,In_775,In_246);
nand U5 (N_5,In_678,In_410);
xnor U6 (N_6,In_831,In_181);
nand U7 (N_7,In_239,In_251);
and U8 (N_8,In_74,In_456);
and U9 (N_9,In_808,In_465);
and U10 (N_10,In_539,In_395);
or U11 (N_11,In_579,In_802);
and U12 (N_12,In_608,In_438);
nand U13 (N_13,In_302,In_245);
and U14 (N_14,In_267,In_500);
nor U15 (N_15,In_325,In_144);
xnor U16 (N_16,In_628,In_799);
nor U17 (N_17,In_420,In_795);
or U18 (N_18,In_146,In_152);
or U19 (N_19,In_762,In_649);
or U20 (N_20,In_450,In_263);
nor U21 (N_21,In_25,In_336);
or U22 (N_22,In_236,In_558);
nor U23 (N_23,In_654,In_478);
and U24 (N_24,In_688,In_783);
or U25 (N_25,In_117,In_972);
nor U26 (N_26,In_602,In_407);
nor U27 (N_27,In_924,In_540);
nand U28 (N_28,In_153,In_839);
and U29 (N_29,In_621,In_520);
nor U30 (N_30,In_987,In_753);
nand U31 (N_31,In_91,In_634);
xor U32 (N_32,In_201,In_755);
nand U33 (N_33,In_161,In_817);
nor U34 (N_34,In_448,In_507);
or U35 (N_35,In_912,In_526);
and U36 (N_36,In_778,In_292);
or U37 (N_37,In_531,In_744);
or U38 (N_38,In_761,In_913);
or U39 (N_39,In_707,In_167);
or U40 (N_40,In_561,In_574);
nand U41 (N_41,In_875,In_51);
and U42 (N_42,In_582,In_547);
and U43 (N_43,In_37,In_889);
or U44 (N_44,In_173,In_16);
nor U45 (N_45,In_985,In_211);
and U46 (N_46,In_10,In_66);
nand U47 (N_47,In_850,In_868);
nand U48 (N_48,In_793,In_741);
xor U49 (N_49,In_403,In_459);
or U50 (N_50,In_269,In_720);
nor U51 (N_51,In_320,In_160);
or U52 (N_52,In_339,In_54);
nor U53 (N_53,In_349,In_232);
nand U54 (N_54,In_187,In_952);
nand U55 (N_55,In_936,In_733);
nor U56 (N_56,In_693,In_931);
nand U57 (N_57,In_133,In_928);
or U58 (N_58,In_414,In_244);
and U59 (N_59,In_464,In_75);
nor U60 (N_60,In_248,In_57);
nand U61 (N_61,In_285,In_278);
nor U62 (N_62,In_98,In_169);
and U63 (N_63,In_976,In_726);
or U64 (N_64,In_929,In_600);
and U65 (N_65,In_217,In_105);
nor U66 (N_66,In_184,In_174);
xor U67 (N_67,In_908,In_881);
nand U68 (N_68,In_695,In_882);
or U69 (N_69,In_280,In_282);
nor U70 (N_70,In_318,In_801);
or U71 (N_71,In_65,In_617);
nor U72 (N_72,In_252,In_104);
and U73 (N_73,In_172,In_609);
or U74 (N_74,In_670,In_93);
and U75 (N_75,In_498,In_369);
nor U76 (N_76,In_920,In_299);
and U77 (N_77,In_235,In_304);
or U78 (N_78,In_87,In_67);
xnor U79 (N_79,In_922,In_333);
and U80 (N_80,In_647,In_723);
nand U81 (N_81,In_378,In_439);
or U82 (N_82,In_696,In_107);
or U83 (N_83,In_264,In_657);
or U84 (N_84,In_650,In_309);
nor U85 (N_85,In_163,In_546);
or U86 (N_86,In_15,In_827);
xor U87 (N_87,In_895,In_727);
nor U88 (N_88,In_525,In_396);
nor U89 (N_89,In_798,In_805);
nand U90 (N_90,In_662,In_991);
nand U91 (N_91,In_978,In_892);
and U92 (N_92,In_517,In_295);
or U93 (N_93,In_522,In_88);
xor U94 (N_94,In_939,In_548);
nor U95 (N_95,In_505,In_145);
and U96 (N_96,In_770,In_797);
or U97 (N_97,In_988,In_864);
and U98 (N_98,In_616,In_914);
or U99 (N_99,In_499,In_642);
or U100 (N_100,In_192,In_998);
nand U101 (N_101,In_253,In_425);
nand U102 (N_102,In_923,In_962);
and U103 (N_103,In_434,In_537);
nand U104 (N_104,In_973,In_619);
or U105 (N_105,In_455,In_220);
nor U106 (N_106,In_825,In_210);
nor U107 (N_107,In_360,In_627);
xor U108 (N_108,In_389,In_472);
and U109 (N_109,In_977,In_614);
or U110 (N_110,In_567,In_300);
nor U111 (N_111,In_297,In_159);
and U112 (N_112,In_535,In_927);
xnor U113 (N_113,In_636,In_969);
nor U114 (N_114,In_261,In_832);
xnor U115 (N_115,In_506,In_428);
nor U116 (N_116,In_194,In_288);
nand U117 (N_117,In_326,In_944);
or U118 (N_118,In_963,In_206);
and U119 (N_119,In_125,In_729);
nand U120 (N_120,In_534,In_379);
nor U121 (N_121,In_45,In_121);
or U122 (N_122,In_114,In_854);
and U123 (N_123,In_335,In_675);
nor U124 (N_124,In_466,In_449);
nor U125 (N_125,In_955,In_485);
or U126 (N_126,In_19,In_958);
xnor U127 (N_127,In_277,In_484);
nor U128 (N_128,In_694,In_4);
and U129 (N_129,In_228,In_256);
nor U130 (N_130,In_471,In_178);
or U131 (N_131,In_112,In_492);
nor U132 (N_132,In_667,In_871);
nor U133 (N_133,In_740,In_780);
or U134 (N_134,In_590,In_750);
nand U135 (N_135,In_214,In_932);
or U136 (N_136,In_833,In_73);
and U137 (N_137,In_565,In_873);
xnor U138 (N_138,In_399,In_990);
xor U139 (N_139,In_258,In_965);
or U140 (N_140,In_400,In_847);
xnor U141 (N_141,In_242,In_938);
nor U142 (N_142,In_370,In_397);
nor U143 (N_143,In_686,In_62);
nor U144 (N_144,In_50,In_983);
nor U145 (N_145,In_286,In_732);
and U146 (N_146,In_718,In_734);
nand U147 (N_147,In_524,In_82);
xor U148 (N_148,In_604,In_821);
xor U149 (N_149,In_852,In_247);
and U150 (N_150,In_593,In_878);
xor U151 (N_151,In_714,In_129);
or U152 (N_152,In_836,In_84);
xnor U153 (N_153,In_327,In_512);
or U154 (N_154,In_766,In_354);
or U155 (N_155,In_735,In_441);
nor U156 (N_156,In_196,In_61);
nand U157 (N_157,In_933,In_555);
nor U158 (N_158,In_108,In_863);
nor U159 (N_159,In_33,In_691);
nor U160 (N_160,In_937,In_652);
nor U161 (N_161,In_717,In_861);
xor U162 (N_162,In_655,In_13);
and U163 (N_163,In_890,In_690);
and U164 (N_164,In_32,In_683);
or U165 (N_165,In_166,In_351);
or U166 (N_166,In_527,In_7);
nand U167 (N_167,In_967,In_997);
nand U168 (N_168,In_28,In_305);
nor U169 (N_169,In_571,In_844);
and U170 (N_170,In_993,In_97);
and U171 (N_171,In_496,In_412);
or U172 (N_172,In_941,In_553);
and U173 (N_173,In_791,In_919);
xnor U174 (N_174,In_989,In_860);
and U175 (N_175,In_897,In_509);
and U176 (N_176,In_934,In_366);
nand U177 (N_177,In_664,In_215);
nor U178 (N_178,In_69,In_568);
or U179 (N_179,In_588,In_221);
nor U180 (N_180,In_230,In_130);
nor U181 (N_181,In_809,In_382);
and U182 (N_182,In_728,In_341);
and U183 (N_183,In_829,In_907);
nand U184 (N_184,In_497,In_594);
xor U185 (N_185,In_3,In_24);
nor U186 (N_186,In_869,In_375);
nand U187 (N_187,In_426,In_671);
nand U188 (N_188,In_901,In_515);
or U189 (N_189,In_612,In_234);
or U190 (N_190,In_754,In_90);
nand U191 (N_191,In_979,In_364);
and U192 (N_192,In_227,In_58);
nand U193 (N_193,In_789,In_648);
and U194 (N_194,In_578,In_205);
or U195 (N_195,In_110,In_651);
and U196 (N_196,In_76,In_822);
or U197 (N_197,In_284,In_307);
or U198 (N_198,In_911,In_190);
nand U199 (N_199,In_180,In_229);
nor U200 (N_200,N_175,In_461);
nand U201 (N_201,In_355,N_111);
or U202 (N_202,In_38,In_193);
nor U203 (N_203,N_12,In_346);
nor U204 (N_204,In_606,In_672);
and U205 (N_205,In_641,In_444);
nor U206 (N_206,In_692,In_0);
or U207 (N_207,N_133,In_820);
and U208 (N_208,In_709,In_281);
nor U209 (N_209,N_109,In_536);
nand U210 (N_210,In_758,In_544);
and U211 (N_211,In_489,N_19);
and U212 (N_212,N_106,N_155);
or U213 (N_213,In_131,In_848);
and U214 (N_214,N_7,N_32);
or U215 (N_215,In_446,In_476);
nand U216 (N_216,In_134,In_12);
nand U217 (N_217,N_128,In_814);
and U218 (N_218,In_632,In_519);
or U219 (N_219,N_92,In_964);
or U220 (N_220,N_33,In_898);
or U221 (N_221,In_142,N_20);
nor U222 (N_222,N_187,N_90);
nor U223 (N_223,In_792,N_60);
xnor U224 (N_224,N_182,In_417);
xor U225 (N_225,In_724,In_462);
and U226 (N_226,In_818,In_685);
or U227 (N_227,N_176,In_684);
nand U228 (N_228,In_807,In_583);
and U229 (N_229,In_473,N_174);
nand U230 (N_230,In_823,In_289);
nand U231 (N_231,In_663,In_529);
nor U232 (N_232,In_946,In_404);
or U233 (N_233,In_273,In_80);
nand U234 (N_234,In_501,In_584);
nor U235 (N_235,N_158,In_203);
nand U236 (N_236,In_502,N_57);
or U237 (N_237,In_530,In_330);
and U238 (N_238,N_197,N_67);
nand U239 (N_239,N_64,In_572);
nand U240 (N_240,In_680,In_622);
nand U241 (N_241,In_372,In_219);
nor U242 (N_242,N_84,N_140);
or U243 (N_243,In_625,N_87);
xnor U244 (N_244,N_102,In_705);
nand U245 (N_245,In_840,In_721);
nand U246 (N_246,In_736,In_352);
nor U247 (N_247,In_126,In_971);
xnor U248 (N_248,In_331,In_408);
xor U249 (N_249,N_31,In_513);
nor U250 (N_250,In_569,In_516);
nor U251 (N_251,In_804,In_708);
xor U252 (N_252,In_368,In_787);
nand U253 (N_253,In_402,N_38);
nor U254 (N_254,N_56,In_812);
nor U255 (N_255,N_93,In_383);
nand U256 (N_256,In_452,In_942);
nor U257 (N_257,N_48,N_0);
and U258 (N_258,In_948,In_371);
nand U259 (N_259,In_586,N_3);
and U260 (N_260,In_44,N_72);
nand U261 (N_261,In_262,N_29);
nand U262 (N_262,In_533,In_623);
nand U263 (N_263,N_184,N_74);
or U264 (N_264,In_276,In_150);
nand U265 (N_265,In_342,In_237);
or U266 (N_266,In_601,N_129);
nor U267 (N_267,In_11,N_2);
nand U268 (N_268,In_949,In_638);
nand U269 (N_269,In_240,In_767);
or U270 (N_270,In_154,N_154);
and U271 (N_271,In_697,N_146);
and U272 (N_272,In_510,In_27);
xnor U273 (N_273,In_811,In_776);
xnor U274 (N_274,In_143,In_162);
and U275 (N_275,In_118,In_469);
or U276 (N_276,In_703,In_554);
nor U277 (N_277,N_97,In_470);
nand U278 (N_278,In_746,In_363);
or U279 (N_279,N_61,In_102);
nand U280 (N_280,In_156,In_293);
and U281 (N_281,N_24,In_384);
or U282 (N_282,In_132,In_781);
or U283 (N_283,In_698,N_141);
nand U284 (N_284,In_893,N_37);
or U285 (N_285,In_319,In_306);
or U286 (N_286,In_828,In_806);
and U287 (N_287,In_917,In_443);
nor U288 (N_288,N_54,In_140);
nor U289 (N_289,In_738,N_94);
and U290 (N_290,In_155,In_658);
nor U291 (N_291,N_165,In_870);
and U292 (N_292,N_166,In_199);
nor U293 (N_293,N_120,In_405);
or U294 (N_294,In_918,In_954);
and U295 (N_295,In_824,In_551);
nor U296 (N_296,In_550,In_592);
nand U297 (N_297,In_845,In_643);
nor U298 (N_298,In_52,In_891);
and U299 (N_299,N_139,N_137);
or U300 (N_300,In_197,In_270);
or U301 (N_301,N_99,In_874);
nand U302 (N_302,N_189,In_858);
nor U303 (N_303,In_92,N_142);
and U304 (N_304,In_290,In_296);
or U305 (N_305,In_225,In_390);
or U306 (N_306,In_857,In_745);
or U307 (N_307,N_47,In_376);
or U308 (N_308,In_629,In_423);
xnor U309 (N_309,N_70,In_49);
nor U310 (N_310,N_4,In_86);
or U311 (N_311,In_921,In_774);
or U312 (N_312,In_182,In_999);
nor U313 (N_313,In_148,N_82);
nand U314 (N_314,In_940,N_65);
and U315 (N_315,In_759,In_440);
xnor U316 (N_316,In_315,In_699);
or U317 (N_317,N_118,In_915);
nor U318 (N_318,N_131,In_254);
and U319 (N_319,In_436,In_59);
or U320 (N_320,In_338,In_367);
nand U321 (N_321,N_77,In_14);
nand U322 (N_322,In_661,N_170);
and U323 (N_323,N_163,N_50);
and U324 (N_324,In_216,N_18);
and U325 (N_325,In_170,In_849);
xnor U326 (N_326,In_120,In_504);
xnor U327 (N_327,In_681,In_23);
or U328 (N_328,N_191,In_803);
nor U329 (N_329,In_322,In_916);
nand U330 (N_330,In_816,In_308);
nand U331 (N_331,In_453,In_982);
nor U332 (N_332,In_872,N_110);
and U333 (N_333,N_196,N_15);
and U334 (N_334,In_386,In_984);
or U335 (N_335,In_311,In_265);
and U336 (N_336,N_186,In_859);
nor U337 (N_337,N_161,In_713);
or U338 (N_338,In_344,In_968);
nor U339 (N_339,In_564,In_365);
or U340 (N_340,In_362,N_8);
and U341 (N_341,In_618,In_549);
nor U342 (N_342,In_737,In_250);
nand U343 (N_343,In_60,In_846);
and U344 (N_344,In_381,In_56);
and U345 (N_345,In_149,N_104);
nor U346 (N_346,In_158,In_768);
or U347 (N_347,In_8,In_855);
or U348 (N_348,In_779,In_431);
or U349 (N_349,In_343,In_994);
or U350 (N_350,In_39,In_943);
and U351 (N_351,N_178,N_10);
nor U352 (N_352,N_66,In_218);
and U353 (N_353,In_127,N_152);
and U354 (N_354,N_167,In_992);
or U355 (N_355,N_62,N_40);
nor U356 (N_356,N_122,In_630);
nor U357 (N_357,In_243,In_659);
or U358 (N_358,In_40,In_885);
or U359 (N_359,In_70,N_143);
or U360 (N_360,In_332,In_925);
nor U361 (N_361,In_391,In_486);
xnor U362 (N_362,In_756,In_961);
nand U363 (N_363,In_48,In_1);
or U364 (N_364,In_523,In_359);
nor U365 (N_365,In_960,In_137);
xor U366 (N_366,In_171,In_613);
and U367 (N_367,In_956,In_538);
or U368 (N_368,In_747,N_30);
and U369 (N_369,In_53,N_39);
or U370 (N_370,In_26,In_841);
xnor U371 (N_371,In_427,In_394);
and U372 (N_372,In_393,N_168);
and U373 (N_373,In_626,In_773);
nor U374 (N_374,N_119,N_105);
or U375 (N_375,In_324,In_557);
nand U376 (N_376,In_89,In_175);
xor U377 (N_377,In_36,In_195);
or U378 (N_378,In_581,In_100);
nand U379 (N_379,In_644,In_771);
nand U380 (N_380,In_702,In_796);
and U381 (N_381,In_435,In_9);
and U382 (N_382,In_862,In_541);
or U383 (N_383,In_323,N_160);
nor U384 (N_384,In_570,In_358);
nand U385 (N_385,N_150,In_866);
nor U386 (N_386,In_202,In_457);
or U387 (N_387,In_268,In_411);
nand U388 (N_388,In_79,In_511);
and U389 (N_389,In_508,In_357);
or U390 (N_390,In_442,In_653);
and U391 (N_391,In_639,In_926);
and U392 (N_392,N_181,In_764);
or U393 (N_393,In_906,In_905);
and U394 (N_394,In_677,In_287);
and U395 (N_395,N_151,N_117);
and U396 (N_396,In_765,N_1);
xnor U397 (N_397,N_25,In_55);
nand U398 (N_398,In_731,N_144);
nor U399 (N_399,N_26,In_495);
nor U400 (N_400,N_204,In_348);
or U401 (N_401,N_232,N_53);
nor U402 (N_402,N_313,N_35);
or U403 (N_403,N_330,In_947);
nor U404 (N_404,In_986,N_347);
xnor U405 (N_405,N_100,N_213);
xor U406 (N_406,In_830,In_730);
and U407 (N_407,N_372,N_355);
and U408 (N_408,In_468,In_398);
or U409 (N_409,In_819,In_521);
nand U410 (N_410,N_81,In_573);
nand U411 (N_411,N_185,N_203);
or U412 (N_412,In_867,N_390);
nor U413 (N_413,In_429,N_28);
nor U414 (N_414,N_356,In_479);
or U415 (N_415,N_98,In_266);
and U416 (N_416,N_36,In_722);
nand U417 (N_417,N_162,In_704);
and U418 (N_418,In_904,In_445);
or U419 (N_419,N_121,In_340);
nor U420 (N_420,N_235,N_242);
nor U421 (N_421,N_254,In_970);
or U422 (N_422,N_58,In_208);
or U423 (N_423,In_490,N_243);
nand U424 (N_424,N_135,In_865);
or U425 (N_425,N_252,N_359);
nand U426 (N_426,In_853,In_880);
nor U427 (N_427,N_341,In_314);
nand U428 (N_428,N_262,In_189);
and U429 (N_429,N_136,N_385);
or U430 (N_430,In_635,N_5);
nand U431 (N_431,In_385,In_603);
nor U432 (N_432,N_169,In_94);
and U433 (N_433,N_246,In_168);
xnor U434 (N_434,In_577,N_283);
or U435 (N_435,N_222,In_31);
and U436 (N_436,In_474,In_597);
nor U437 (N_437,N_157,In_209);
nand U438 (N_438,In_380,N_52);
nor U439 (N_439,In_406,In_409);
xor U440 (N_440,N_75,N_207);
and U441 (N_441,N_376,N_343);
xor U442 (N_442,In_179,In_96);
nor U443 (N_443,In_200,In_995);
or U444 (N_444,N_225,N_339);
and U445 (N_445,In_463,In_101);
nand U446 (N_446,In_930,N_362);
nand U447 (N_447,In_815,N_138);
nor U448 (N_448,In_47,N_304);
and U449 (N_449,N_231,N_299);
and U450 (N_450,N_224,In_183);
nor U451 (N_451,N_300,N_229);
or U452 (N_452,In_974,N_171);
nand U453 (N_453,N_321,N_379);
and U454 (N_454,In_122,In_116);
nor U455 (N_455,N_337,N_260);
nor U456 (N_456,In_725,N_269);
nor U457 (N_457,In_598,N_327);
and U458 (N_458,In_701,N_51);
xnor U459 (N_459,N_394,N_380);
or U460 (N_460,N_114,In_834);
or U461 (N_461,In_95,N_272);
nor U462 (N_462,N_149,N_209);
xor U463 (N_463,N_294,N_360);
or U464 (N_464,N_76,In_786);
nor U465 (N_465,In_373,In_945);
and U466 (N_466,N_200,N_253);
or U467 (N_467,N_46,N_126);
xor U468 (N_468,N_258,In_562);
nor U469 (N_469,N_363,N_340);
and U470 (N_470,In_763,N_292);
or U471 (N_471,N_112,In_454);
or U472 (N_472,In_482,N_80);
and U473 (N_473,In_879,N_251);
and U474 (N_474,N_108,In_41);
and U475 (N_475,In_353,In_605);
and U476 (N_476,In_666,N_383);
nand U477 (N_477,N_249,N_153);
nand U478 (N_478,N_384,In_139);
or U479 (N_479,N_16,N_215);
nor U480 (N_480,N_287,In_996);
and U481 (N_481,N_69,N_210);
nand U482 (N_482,In_518,N_298);
nor U483 (N_483,N_49,N_218);
nand U484 (N_484,In_313,In_71);
nor U485 (N_485,N_183,In_585);
nor U486 (N_486,In_413,In_712);
or U487 (N_487,In_416,In_272);
nand U488 (N_488,In_560,N_289);
and U489 (N_489,In_856,N_282);
or U490 (N_490,N_329,N_371);
nor U491 (N_491,N_83,N_198);
nor U492 (N_492,N_22,In_123);
nor U493 (N_493,N_9,N_217);
nor U494 (N_494,In_477,In_903);
nand U495 (N_495,N_309,In_563);
nor U496 (N_496,N_43,In_34);
or U497 (N_497,N_116,In_85);
xor U498 (N_498,N_255,N_214);
and U499 (N_499,In_656,N_370);
or U500 (N_500,N_281,N_202);
xor U501 (N_501,In_430,In_611);
xnor U502 (N_502,In_966,N_395);
and U503 (N_503,In_888,N_6);
nand U504 (N_504,In_599,N_291);
nand U505 (N_505,In_700,In_837);
nand U506 (N_506,In_310,In_682);
xnor U507 (N_507,N_348,In_543);
nor U508 (N_508,N_11,N_320);
nor U509 (N_509,N_228,In_233);
nor U510 (N_510,In_222,N_59);
nor U511 (N_511,In_475,N_244);
or U512 (N_512,In_716,In_345);
or U513 (N_513,In_676,N_350);
nor U514 (N_514,In_164,In_813);
and U515 (N_515,In_886,In_361);
and U516 (N_516,In_576,In_481);
and U517 (N_517,In_843,In_238);
nor U518 (N_518,In_198,In_631);
nand U519 (N_519,In_294,In_552);
nand U520 (N_520,In_17,N_86);
or U521 (N_521,N_132,N_301);
nor U522 (N_522,In_668,N_303);
nor U523 (N_523,In_29,N_219);
nor U524 (N_524,N_288,N_238);
nor U525 (N_525,N_208,N_55);
nor U526 (N_526,N_365,In_566);
and U527 (N_527,N_159,N_257);
nand U528 (N_528,N_353,In_316);
and U529 (N_529,N_393,In_620);
xor U530 (N_530,N_190,In_959);
nor U531 (N_531,In_800,In_78);
xor U532 (N_532,N_336,N_352);
nor U533 (N_533,N_127,In_899);
nand U534 (N_534,In_719,In_260);
nor U535 (N_535,In_589,In_782);
and U536 (N_536,In_910,N_316);
nand U537 (N_537,N_125,In_610);
or U538 (N_538,In_487,N_267);
and U539 (N_539,N_307,N_188);
or U540 (N_540,In_935,In_769);
or U541 (N_541,N_280,N_349);
nand U542 (N_542,N_369,N_233);
or U543 (N_543,In_147,In_424);
or U544 (N_544,In_301,N_164);
or U545 (N_545,In_119,In_392);
nand U546 (N_546,In_711,N_201);
or U547 (N_547,In_226,N_323);
nor U548 (N_548,In_22,In_165);
and U549 (N_549,In_249,N_172);
or U550 (N_550,In_151,In_757);
nand U551 (N_551,N_248,N_279);
and U552 (N_552,N_308,In_5);
nor U553 (N_553,In_419,In_43);
or U554 (N_554,In_637,N_268);
xnor U555 (N_555,N_302,In_415);
nor U556 (N_556,N_354,In_303);
xnor U557 (N_557,In_135,N_241);
nor U558 (N_558,N_239,N_13);
and U559 (N_559,In_274,N_335);
nor U560 (N_560,In_491,In_660);
nor U561 (N_561,In_421,N_324);
or U562 (N_562,N_361,In_951);
and U563 (N_563,In_224,N_389);
nand U564 (N_564,N_314,N_351);
nor U565 (N_565,In_953,N_367);
and U566 (N_566,N_130,In_128);
or U567 (N_567,In_255,N_14);
nor U568 (N_568,In_665,In_749);
and U569 (N_569,N_364,N_377);
nand U570 (N_570,N_230,N_387);
nor U571 (N_571,N_45,N_88);
and U572 (N_572,N_392,In_545);
or U573 (N_573,N_205,In_42);
nor U574 (N_574,In_109,N_295);
or U575 (N_575,In_503,In_99);
nand U576 (N_576,In_231,N_334);
and U577 (N_577,N_177,In_103);
nor U578 (N_578,In_742,N_312);
or U579 (N_579,In_575,In_884);
nand U580 (N_580,N_264,In_138);
and U581 (N_581,N_346,In_640);
or U582 (N_582,In_794,N_236);
nor U583 (N_583,N_325,N_274);
nor U584 (N_584,N_85,In_20);
and U585 (N_585,N_378,N_286);
or U586 (N_586,In_488,In_981);
or U587 (N_587,N_338,In_432);
xnor U588 (N_588,N_68,In_887);
xor U589 (N_589,N_322,N_192);
nand U590 (N_590,In_777,In_883);
nand U591 (N_591,N_344,In_433);
or U592 (N_592,N_227,N_332);
or U593 (N_593,N_226,In_900);
or U594 (N_594,N_234,N_173);
nand U595 (N_595,In_851,N_285);
nor U596 (N_596,N_326,In_788);
nor U597 (N_597,In_213,N_115);
and U598 (N_598,N_21,In_494);
or U599 (N_599,In_673,In_377);
nor U600 (N_600,N_559,N_505);
nand U601 (N_601,N_503,In_18);
nor U602 (N_602,N_555,In_191);
nor U603 (N_603,N_477,In_115);
or U604 (N_604,N_582,N_240);
nor U605 (N_605,N_465,N_468);
or U606 (N_606,In_291,N_578);
and U607 (N_607,N_567,In_356);
or U608 (N_608,N_305,In_957);
xor U609 (N_609,N_550,N_96);
nand U610 (N_610,N_265,N_507);
or U611 (N_611,N_41,In_909);
or U612 (N_612,In_21,N_475);
nand U613 (N_613,N_467,N_402);
and U614 (N_614,N_527,In_6);
or U615 (N_615,N_488,N_560);
xnor U616 (N_616,N_482,N_206);
or U617 (N_617,N_414,N_596);
and U618 (N_618,N_440,N_476);
nand U619 (N_619,N_223,N_409);
or U620 (N_620,In_223,N_566);
nor U621 (N_621,In_633,N_569);
or U622 (N_622,In_674,N_436);
or U623 (N_623,In_607,N_516);
or U624 (N_624,In_279,N_469);
or U625 (N_625,N_595,N_435);
nand U626 (N_626,N_584,N_495);
nand U627 (N_627,N_407,N_266);
nor U628 (N_628,In_388,N_480);
and U629 (N_629,N_408,N_95);
nor U630 (N_630,N_345,N_557);
or U631 (N_631,In_772,In_212);
nor U632 (N_632,N_17,N_506);
nand U633 (N_633,N_89,N_532);
nand U634 (N_634,N_579,N_421);
and U635 (N_635,N_589,N_442);
nand U636 (N_636,N_474,N_461);
nand U637 (N_637,In_559,N_342);
nor U638 (N_638,In_447,N_521);
and U639 (N_639,N_454,N_261);
nand U640 (N_640,N_439,N_382);
or U641 (N_641,N_554,In_186);
xor U642 (N_642,N_552,In_748);
and U643 (N_643,N_573,N_574);
nand U644 (N_644,N_366,N_373);
and U645 (N_645,N_563,N_245);
nor U646 (N_646,In_689,N_511);
or U647 (N_647,In_257,N_145);
or U648 (N_648,N_564,In_706);
nor U649 (N_649,N_401,N_462);
nand U650 (N_650,In_587,N_497);
nor U651 (N_651,In_347,In_624);
or U652 (N_652,N_418,N_478);
and U653 (N_653,N_259,N_451);
or U654 (N_654,In_826,In_532);
or U655 (N_655,N_572,N_277);
and U656 (N_656,In_877,In_752);
or U657 (N_657,N_545,In_374);
or U658 (N_658,In_418,N_508);
and U659 (N_659,N_597,N_276);
or U660 (N_660,N_358,N_78);
nor U661 (N_661,N_107,In_458);
or U662 (N_662,In_157,N_583);
nor U663 (N_663,N_549,N_510);
and U664 (N_664,N_180,N_113);
nor U665 (N_665,N_391,N_428);
xnor U666 (N_666,In_743,In_842);
or U667 (N_667,In_321,In_483);
nor U668 (N_668,In_387,N_296);
and U669 (N_669,N_124,N_463);
nor U670 (N_670,In_687,N_381);
or U671 (N_671,N_523,N_522);
or U672 (N_672,N_73,N_293);
and U673 (N_673,In_63,N_447);
nand U674 (N_674,N_452,In_83);
or U675 (N_675,In_328,N_538);
and U676 (N_676,In_177,N_388);
and U677 (N_677,N_250,In_480);
nor U678 (N_678,N_400,N_221);
nand U679 (N_679,N_63,In_113);
nand U680 (N_680,N_542,N_529);
nor U681 (N_681,N_491,N_431);
and U682 (N_682,N_27,N_466);
and U683 (N_683,N_416,N_518);
or U684 (N_684,In_422,In_894);
xor U685 (N_685,N_101,In_514);
nand U686 (N_686,N_278,N_485);
and U687 (N_687,N_357,N_457);
and U688 (N_688,N_195,In_312);
or U689 (N_689,N_399,N_571);
xor U690 (N_690,N_588,N_450);
nor U691 (N_691,N_501,N_537);
or U692 (N_692,N_446,N_422);
nand U693 (N_693,N_500,In_337);
nand U694 (N_694,N_271,In_980);
and U695 (N_695,In_72,N_484);
nand U696 (N_696,In_710,N_455);
nor U697 (N_697,N_594,N_430);
and U698 (N_698,N_492,N_487);
or U699 (N_699,N_319,N_486);
and U700 (N_700,In_615,N_496);
xnor U701 (N_701,N_576,In_283);
nor U702 (N_702,N_432,N_513);
xor U703 (N_703,In_176,N_275);
nand U704 (N_704,In_271,N_290);
or U705 (N_705,N_548,N_565);
and U706 (N_706,N_591,N_449);
nand U707 (N_707,N_273,N_134);
nand U708 (N_708,N_483,N_396);
xnor U709 (N_709,In_64,N_71);
or U710 (N_710,N_592,N_331);
and U711 (N_711,In_401,In_460);
nor U712 (N_712,N_512,In_669);
nand U713 (N_713,In_838,In_437);
or U714 (N_714,N_443,N_562);
nand U715 (N_715,In_760,N_237);
or U716 (N_716,N_156,In_136);
nor U717 (N_717,N_541,In_493);
nor U718 (N_718,N_490,N_551);
and U719 (N_719,In_591,In_646);
nand U720 (N_720,N_425,N_403);
and U721 (N_721,N_147,N_411);
or U722 (N_722,N_520,N_437);
and U723 (N_723,N_581,N_464);
nand U724 (N_724,N_405,N_216);
or U725 (N_725,N_317,N_593);
or U726 (N_726,N_193,In_950);
or U727 (N_727,N_456,N_458);
and U728 (N_728,In_739,In_715);
xor U729 (N_729,N_445,N_297);
or U730 (N_730,N_412,N_547);
or U731 (N_731,N_535,N_599);
or U732 (N_732,In_2,N_247);
or U733 (N_733,N_553,N_211);
and U734 (N_734,In_645,N_585);
and U735 (N_735,N_498,N_453);
nor U736 (N_736,N_398,N_509);
and U737 (N_737,In_77,N_528);
nor U738 (N_738,In_81,N_459);
xor U739 (N_739,N_410,In_207);
or U740 (N_740,N_423,N_79);
nor U741 (N_741,In_785,N_514);
xor U742 (N_742,N_519,N_499);
nor U743 (N_743,In_111,In_185);
nor U744 (N_744,N_570,N_546);
nand U745 (N_745,In_106,N_438);
and U746 (N_746,N_515,In_975);
nor U747 (N_747,N_284,In_896);
or U748 (N_748,N_91,In_528);
nor U749 (N_749,In_902,In_580);
and U750 (N_750,N_270,In_451);
xnor U751 (N_751,N_460,N_179);
and U752 (N_752,N_420,N_575);
nand U753 (N_753,N_540,N_413);
and U754 (N_754,In_35,N_256);
nor U755 (N_755,N_530,In_679);
nor U756 (N_756,In_329,In_751);
nor U757 (N_757,N_586,N_429);
nand U758 (N_758,In_204,N_199);
or U759 (N_759,N_433,N_34);
or U760 (N_760,N_374,N_424);
nand U761 (N_761,N_23,N_417);
and U762 (N_762,N_368,N_479);
nand U763 (N_763,N_148,N_533);
nand U764 (N_764,N_524,N_311);
and U765 (N_765,N_315,N_489);
or U766 (N_766,N_123,N_472);
nor U767 (N_767,N_481,N_493);
xor U768 (N_768,N_42,N_328);
xor U769 (N_769,In_141,N_539);
xor U770 (N_770,N_526,N_598);
or U771 (N_771,N_502,N_473);
nor U772 (N_772,N_504,N_415);
or U773 (N_773,In_542,In_556);
and U774 (N_774,N_525,In_275);
or U775 (N_775,N_558,N_590);
xnor U776 (N_776,In_298,N_318);
and U777 (N_777,In_350,In_784);
nor U778 (N_778,N_44,N_568);
nor U779 (N_779,N_531,In_124);
nor U780 (N_780,In_241,N_577);
nor U781 (N_781,N_194,In_467);
or U782 (N_782,N_494,N_441);
nand U783 (N_783,N_212,N_444);
nand U784 (N_784,N_333,In_835);
nor U785 (N_785,N_448,N_404);
nand U786 (N_786,N_544,In_188);
nor U787 (N_787,N_534,N_434);
xor U788 (N_788,N_543,In_259);
xnor U789 (N_789,In_68,In_876);
nor U790 (N_790,N_580,N_427);
xnor U791 (N_791,N_587,N_397);
or U792 (N_792,N_375,N_517);
and U793 (N_793,N_561,N_406);
nand U794 (N_794,N_220,N_310);
and U795 (N_795,N_419,N_426);
or U796 (N_796,N_103,N_470);
or U797 (N_797,N_471,N_556);
xnor U798 (N_798,N_306,N_536);
or U799 (N_799,N_386,N_263);
nor U800 (N_800,N_775,N_668);
nand U801 (N_801,N_601,N_796);
or U802 (N_802,N_754,N_744);
and U803 (N_803,N_799,N_696);
nor U804 (N_804,N_629,N_615);
or U805 (N_805,N_706,N_782);
nand U806 (N_806,N_644,N_751);
or U807 (N_807,N_697,N_616);
nand U808 (N_808,N_752,N_678);
nor U809 (N_809,N_654,N_661);
or U810 (N_810,N_603,N_762);
nand U811 (N_811,N_734,N_710);
nor U812 (N_812,N_764,N_620);
nor U813 (N_813,N_667,N_631);
and U814 (N_814,N_643,N_735);
and U815 (N_815,N_784,N_665);
or U816 (N_816,N_666,N_619);
or U817 (N_817,N_771,N_779);
nand U818 (N_818,N_709,N_756);
nor U819 (N_819,N_640,N_691);
or U820 (N_820,N_625,N_653);
or U821 (N_821,N_600,N_611);
nor U822 (N_822,N_770,N_690);
or U823 (N_823,N_730,N_617);
and U824 (N_824,N_648,N_731);
xor U825 (N_825,N_726,N_693);
nor U826 (N_826,N_733,N_685);
nand U827 (N_827,N_659,N_742);
xor U828 (N_828,N_669,N_642);
and U829 (N_829,N_753,N_651);
nor U830 (N_830,N_634,N_767);
or U831 (N_831,N_628,N_676);
or U832 (N_832,N_766,N_757);
and U833 (N_833,N_679,N_739);
or U834 (N_834,N_602,N_633);
nor U835 (N_835,N_637,N_684);
nor U836 (N_836,N_723,N_680);
nor U837 (N_837,N_790,N_740);
or U838 (N_838,N_686,N_785);
nor U839 (N_839,N_621,N_724);
nand U840 (N_840,N_689,N_722);
or U841 (N_841,N_660,N_606);
nor U842 (N_842,N_798,N_647);
or U843 (N_843,N_688,N_604);
nand U844 (N_844,N_708,N_687);
and U845 (N_845,N_732,N_759);
nor U846 (N_846,N_761,N_681);
nor U847 (N_847,N_783,N_698);
and U848 (N_848,N_675,N_704);
or U849 (N_849,N_672,N_774);
nor U850 (N_850,N_677,N_694);
and U851 (N_851,N_765,N_662);
nand U852 (N_852,N_683,N_674);
xor U853 (N_853,N_632,N_618);
nor U854 (N_854,N_746,N_636);
or U855 (N_855,N_773,N_670);
or U856 (N_856,N_786,N_699);
nand U857 (N_857,N_657,N_758);
nand U858 (N_858,N_789,N_741);
or U859 (N_859,N_777,N_695);
or U860 (N_860,N_622,N_788);
xnor U861 (N_861,N_728,N_614);
nand U862 (N_862,N_792,N_692);
xor U863 (N_863,N_797,N_645);
nor U864 (N_864,N_729,N_727);
and U865 (N_865,N_763,N_655);
or U866 (N_866,N_610,N_793);
or U867 (N_867,N_652,N_738);
or U868 (N_868,N_715,N_719);
nand U869 (N_869,N_747,N_748);
nor U870 (N_870,N_635,N_673);
or U871 (N_871,N_701,N_682);
nand U872 (N_872,N_613,N_671);
and U873 (N_873,N_609,N_641);
nand U874 (N_874,N_702,N_781);
or U875 (N_875,N_658,N_720);
xor U876 (N_876,N_718,N_605);
and U877 (N_877,N_760,N_717);
xnor U878 (N_878,N_745,N_649);
nor U879 (N_879,N_711,N_794);
nor U880 (N_880,N_626,N_650);
nand U881 (N_881,N_612,N_627);
nor U882 (N_882,N_736,N_712);
and U883 (N_883,N_716,N_791);
or U884 (N_884,N_721,N_743);
and U885 (N_885,N_663,N_703);
or U886 (N_886,N_769,N_780);
and U887 (N_887,N_749,N_656);
nand U888 (N_888,N_646,N_776);
nand U889 (N_889,N_638,N_700);
nand U890 (N_890,N_755,N_705);
and U891 (N_891,N_737,N_607);
and U892 (N_892,N_787,N_623);
nor U893 (N_893,N_768,N_713);
nand U894 (N_894,N_795,N_778);
nand U895 (N_895,N_725,N_664);
nor U896 (N_896,N_707,N_772);
and U897 (N_897,N_750,N_630);
nor U898 (N_898,N_714,N_624);
and U899 (N_899,N_608,N_639);
nand U900 (N_900,N_769,N_626);
or U901 (N_901,N_789,N_751);
and U902 (N_902,N_705,N_710);
and U903 (N_903,N_730,N_773);
nand U904 (N_904,N_789,N_610);
xnor U905 (N_905,N_731,N_608);
or U906 (N_906,N_671,N_735);
nor U907 (N_907,N_667,N_734);
xor U908 (N_908,N_653,N_610);
and U909 (N_909,N_756,N_710);
and U910 (N_910,N_776,N_691);
nand U911 (N_911,N_697,N_759);
xnor U912 (N_912,N_726,N_788);
nor U913 (N_913,N_776,N_703);
or U914 (N_914,N_653,N_607);
or U915 (N_915,N_751,N_683);
and U916 (N_916,N_695,N_790);
nand U917 (N_917,N_628,N_751);
nand U918 (N_918,N_707,N_659);
and U919 (N_919,N_659,N_679);
and U920 (N_920,N_754,N_632);
and U921 (N_921,N_652,N_680);
nor U922 (N_922,N_763,N_687);
and U923 (N_923,N_706,N_710);
or U924 (N_924,N_793,N_748);
nor U925 (N_925,N_613,N_601);
and U926 (N_926,N_783,N_738);
or U927 (N_927,N_743,N_611);
nor U928 (N_928,N_757,N_684);
or U929 (N_929,N_674,N_688);
and U930 (N_930,N_691,N_703);
nor U931 (N_931,N_710,N_666);
and U932 (N_932,N_728,N_608);
and U933 (N_933,N_714,N_795);
and U934 (N_934,N_757,N_700);
and U935 (N_935,N_613,N_637);
or U936 (N_936,N_753,N_769);
and U937 (N_937,N_653,N_756);
nor U938 (N_938,N_652,N_666);
nor U939 (N_939,N_611,N_701);
or U940 (N_940,N_797,N_736);
and U941 (N_941,N_680,N_778);
and U942 (N_942,N_601,N_741);
or U943 (N_943,N_769,N_609);
nor U944 (N_944,N_668,N_638);
nor U945 (N_945,N_740,N_745);
nor U946 (N_946,N_730,N_779);
nor U947 (N_947,N_793,N_634);
nor U948 (N_948,N_777,N_643);
and U949 (N_949,N_752,N_725);
xor U950 (N_950,N_644,N_768);
and U951 (N_951,N_659,N_648);
or U952 (N_952,N_783,N_658);
xnor U953 (N_953,N_640,N_791);
nand U954 (N_954,N_712,N_668);
or U955 (N_955,N_605,N_763);
nand U956 (N_956,N_641,N_774);
or U957 (N_957,N_790,N_742);
nand U958 (N_958,N_793,N_759);
nand U959 (N_959,N_759,N_721);
xor U960 (N_960,N_643,N_753);
nand U961 (N_961,N_663,N_760);
and U962 (N_962,N_655,N_679);
or U963 (N_963,N_702,N_745);
nand U964 (N_964,N_679,N_626);
xor U965 (N_965,N_798,N_682);
and U966 (N_966,N_608,N_707);
and U967 (N_967,N_644,N_775);
and U968 (N_968,N_694,N_671);
or U969 (N_969,N_645,N_721);
nor U970 (N_970,N_601,N_682);
or U971 (N_971,N_701,N_767);
nor U972 (N_972,N_664,N_738);
or U973 (N_973,N_648,N_711);
nand U974 (N_974,N_655,N_641);
nand U975 (N_975,N_689,N_627);
or U976 (N_976,N_613,N_685);
nor U977 (N_977,N_743,N_787);
xnor U978 (N_978,N_727,N_759);
and U979 (N_979,N_642,N_620);
nand U980 (N_980,N_689,N_751);
xnor U981 (N_981,N_626,N_638);
or U982 (N_982,N_743,N_784);
or U983 (N_983,N_613,N_765);
nor U984 (N_984,N_616,N_618);
or U985 (N_985,N_718,N_799);
nor U986 (N_986,N_770,N_709);
and U987 (N_987,N_771,N_688);
nand U988 (N_988,N_750,N_795);
or U989 (N_989,N_749,N_601);
and U990 (N_990,N_642,N_634);
or U991 (N_991,N_688,N_725);
or U992 (N_992,N_613,N_670);
and U993 (N_993,N_604,N_630);
or U994 (N_994,N_787,N_746);
or U995 (N_995,N_756,N_652);
nand U996 (N_996,N_786,N_640);
xnor U997 (N_997,N_649,N_670);
or U998 (N_998,N_762,N_735);
or U999 (N_999,N_618,N_749);
xnor U1000 (N_1000,N_951,N_814);
or U1001 (N_1001,N_917,N_910);
nand U1002 (N_1002,N_820,N_944);
or U1003 (N_1003,N_872,N_989);
and U1004 (N_1004,N_986,N_976);
nand U1005 (N_1005,N_822,N_840);
nand U1006 (N_1006,N_988,N_992);
xnor U1007 (N_1007,N_816,N_853);
and U1008 (N_1008,N_957,N_905);
nand U1009 (N_1009,N_893,N_963);
and U1010 (N_1010,N_929,N_943);
and U1011 (N_1011,N_983,N_810);
nor U1012 (N_1012,N_881,N_940);
and U1013 (N_1013,N_859,N_911);
and U1014 (N_1014,N_995,N_869);
and U1015 (N_1015,N_952,N_874);
or U1016 (N_1016,N_873,N_980);
nor U1017 (N_1017,N_819,N_839);
xor U1018 (N_1018,N_835,N_804);
or U1019 (N_1019,N_999,N_987);
xor U1020 (N_1020,N_897,N_948);
nor U1021 (N_1021,N_954,N_933);
and U1022 (N_1022,N_808,N_857);
and U1023 (N_1023,N_867,N_908);
nand U1024 (N_1024,N_877,N_896);
nor U1025 (N_1025,N_931,N_899);
nor U1026 (N_1026,N_824,N_817);
nor U1027 (N_1027,N_961,N_997);
nor U1028 (N_1028,N_971,N_856);
or U1029 (N_1029,N_886,N_942);
nand U1030 (N_1030,N_941,N_852);
or U1031 (N_1031,N_918,N_862);
nand U1032 (N_1032,N_876,N_845);
and U1033 (N_1033,N_879,N_902);
xnor U1034 (N_1034,N_937,N_815);
xnor U1035 (N_1035,N_985,N_849);
nor U1036 (N_1036,N_826,N_960);
nand U1037 (N_1037,N_900,N_811);
nor U1038 (N_1038,N_892,N_861);
nor U1039 (N_1039,N_904,N_866);
nor U1040 (N_1040,N_975,N_990);
xor U1041 (N_1041,N_970,N_837);
or U1042 (N_1042,N_928,N_934);
or U1043 (N_1043,N_973,N_972);
nand U1044 (N_1044,N_935,N_907);
nor U1045 (N_1045,N_967,N_883);
and U1046 (N_1046,N_801,N_813);
nand U1047 (N_1047,N_939,N_834);
nand U1048 (N_1048,N_865,N_982);
or U1049 (N_1049,N_821,N_885);
and U1050 (N_1050,N_895,N_964);
nand U1051 (N_1051,N_828,N_851);
xnor U1052 (N_1052,N_906,N_812);
and U1053 (N_1053,N_932,N_833);
or U1054 (N_1054,N_950,N_860);
nor U1055 (N_1055,N_884,N_887);
or U1056 (N_1056,N_930,N_938);
nor U1057 (N_1057,N_946,N_949);
nor U1058 (N_1058,N_844,N_831);
or U1059 (N_1059,N_846,N_855);
or U1060 (N_1060,N_854,N_974);
xnor U1061 (N_1061,N_920,N_875);
or U1062 (N_1062,N_955,N_850);
and U1063 (N_1063,N_889,N_945);
xor U1064 (N_1064,N_864,N_912);
nand U1065 (N_1065,N_962,N_924);
nand U1066 (N_1066,N_806,N_977);
and U1067 (N_1067,N_800,N_991);
nand U1068 (N_1068,N_981,N_996);
nor U1069 (N_1069,N_803,N_979);
and U1070 (N_1070,N_805,N_965);
or U1071 (N_1071,N_830,N_903);
xor U1072 (N_1072,N_802,N_968);
or U1073 (N_1073,N_871,N_858);
nand U1074 (N_1074,N_993,N_901);
and U1075 (N_1075,N_868,N_922);
nand U1076 (N_1076,N_919,N_894);
xnor U1077 (N_1077,N_888,N_916);
and U1078 (N_1078,N_994,N_947);
nor U1079 (N_1079,N_880,N_836);
nand U1080 (N_1080,N_843,N_925);
and U1081 (N_1081,N_923,N_914);
or U1082 (N_1082,N_936,N_847);
nand U1083 (N_1083,N_913,N_915);
nand U1084 (N_1084,N_927,N_823);
xor U1085 (N_1085,N_882,N_838);
and U1086 (N_1086,N_926,N_959);
nand U1087 (N_1087,N_842,N_984);
nor U1088 (N_1088,N_998,N_825);
nand U1089 (N_1089,N_978,N_956);
nor U1090 (N_1090,N_827,N_841);
nor U1091 (N_1091,N_966,N_958);
or U1092 (N_1092,N_809,N_921);
nor U1093 (N_1093,N_969,N_953);
and U1094 (N_1094,N_832,N_848);
or U1095 (N_1095,N_898,N_818);
nor U1096 (N_1096,N_878,N_909);
or U1097 (N_1097,N_807,N_863);
or U1098 (N_1098,N_870,N_829);
and U1099 (N_1099,N_891,N_890);
nor U1100 (N_1100,N_947,N_902);
nor U1101 (N_1101,N_805,N_945);
nand U1102 (N_1102,N_835,N_832);
xnor U1103 (N_1103,N_838,N_973);
nor U1104 (N_1104,N_864,N_834);
or U1105 (N_1105,N_888,N_966);
nor U1106 (N_1106,N_831,N_816);
and U1107 (N_1107,N_923,N_986);
or U1108 (N_1108,N_976,N_949);
and U1109 (N_1109,N_803,N_963);
and U1110 (N_1110,N_837,N_962);
xnor U1111 (N_1111,N_837,N_959);
nor U1112 (N_1112,N_808,N_957);
or U1113 (N_1113,N_908,N_844);
nor U1114 (N_1114,N_911,N_914);
and U1115 (N_1115,N_898,N_835);
or U1116 (N_1116,N_932,N_882);
and U1117 (N_1117,N_983,N_923);
nand U1118 (N_1118,N_990,N_940);
xor U1119 (N_1119,N_992,N_818);
nand U1120 (N_1120,N_939,N_900);
nand U1121 (N_1121,N_865,N_945);
and U1122 (N_1122,N_806,N_901);
nand U1123 (N_1123,N_805,N_894);
or U1124 (N_1124,N_910,N_918);
nor U1125 (N_1125,N_962,N_902);
or U1126 (N_1126,N_898,N_844);
nand U1127 (N_1127,N_810,N_827);
nand U1128 (N_1128,N_935,N_840);
or U1129 (N_1129,N_829,N_835);
xnor U1130 (N_1130,N_835,N_924);
xor U1131 (N_1131,N_925,N_915);
nand U1132 (N_1132,N_880,N_933);
and U1133 (N_1133,N_876,N_813);
and U1134 (N_1134,N_901,N_891);
nor U1135 (N_1135,N_804,N_870);
nor U1136 (N_1136,N_832,N_992);
nor U1137 (N_1137,N_895,N_975);
xor U1138 (N_1138,N_870,N_923);
nand U1139 (N_1139,N_803,N_933);
or U1140 (N_1140,N_926,N_964);
nand U1141 (N_1141,N_916,N_881);
or U1142 (N_1142,N_820,N_977);
xor U1143 (N_1143,N_873,N_878);
nand U1144 (N_1144,N_888,N_926);
and U1145 (N_1145,N_944,N_959);
xor U1146 (N_1146,N_809,N_969);
or U1147 (N_1147,N_911,N_935);
or U1148 (N_1148,N_944,N_867);
nor U1149 (N_1149,N_987,N_895);
nor U1150 (N_1150,N_954,N_958);
xor U1151 (N_1151,N_943,N_864);
nand U1152 (N_1152,N_970,N_807);
nor U1153 (N_1153,N_842,N_949);
or U1154 (N_1154,N_805,N_881);
and U1155 (N_1155,N_831,N_906);
nand U1156 (N_1156,N_836,N_890);
nand U1157 (N_1157,N_905,N_894);
and U1158 (N_1158,N_917,N_873);
nand U1159 (N_1159,N_922,N_923);
xor U1160 (N_1160,N_962,N_921);
nand U1161 (N_1161,N_913,N_956);
xor U1162 (N_1162,N_951,N_894);
or U1163 (N_1163,N_865,N_815);
and U1164 (N_1164,N_914,N_955);
or U1165 (N_1165,N_901,N_964);
or U1166 (N_1166,N_805,N_826);
or U1167 (N_1167,N_980,N_893);
and U1168 (N_1168,N_871,N_984);
nor U1169 (N_1169,N_894,N_910);
nand U1170 (N_1170,N_946,N_929);
nand U1171 (N_1171,N_952,N_986);
or U1172 (N_1172,N_977,N_826);
and U1173 (N_1173,N_986,N_826);
and U1174 (N_1174,N_858,N_922);
or U1175 (N_1175,N_872,N_832);
nand U1176 (N_1176,N_896,N_892);
or U1177 (N_1177,N_852,N_867);
nor U1178 (N_1178,N_942,N_811);
nor U1179 (N_1179,N_801,N_858);
and U1180 (N_1180,N_818,N_944);
nor U1181 (N_1181,N_972,N_857);
nor U1182 (N_1182,N_955,N_848);
xor U1183 (N_1183,N_924,N_883);
nor U1184 (N_1184,N_939,N_821);
or U1185 (N_1185,N_837,N_847);
and U1186 (N_1186,N_852,N_876);
nand U1187 (N_1187,N_985,N_947);
nor U1188 (N_1188,N_879,N_958);
xor U1189 (N_1189,N_807,N_844);
and U1190 (N_1190,N_831,N_936);
nor U1191 (N_1191,N_800,N_898);
xor U1192 (N_1192,N_948,N_887);
nand U1193 (N_1193,N_829,N_937);
nand U1194 (N_1194,N_957,N_920);
and U1195 (N_1195,N_863,N_823);
or U1196 (N_1196,N_977,N_953);
nand U1197 (N_1197,N_851,N_886);
xor U1198 (N_1198,N_978,N_845);
nor U1199 (N_1199,N_930,N_865);
nand U1200 (N_1200,N_1149,N_1182);
or U1201 (N_1201,N_1028,N_1067);
nand U1202 (N_1202,N_1011,N_1018);
or U1203 (N_1203,N_1173,N_1136);
and U1204 (N_1204,N_1021,N_1064);
xnor U1205 (N_1205,N_1057,N_1068);
or U1206 (N_1206,N_1165,N_1087);
and U1207 (N_1207,N_1060,N_1138);
nor U1208 (N_1208,N_1144,N_1192);
nand U1209 (N_1209,N_1184,N_1003);
xnor U1210 (N_1210,N_1131,N_1053);
and U1211 (N_1211,N_1155,N_1098);
xor U1212 (N_1212,N_1110,N_1059);
and U1213 (N_1213,N_1146,N_1049);
and U1214 (N_1214,N_1196,N_1140);
nand U1215 (N_1215,N_1169,N_1020);
or U1216 (N_1216,N_1107,N_1004);
nand U1217 (N_1217,N_1037,N_1164);
nor U1218 (N_1218,N_1034,N_1023);
nand U1219 (N_1219,N_1139,N_1152);
and U1220 (N_1220,N_1074,N_1130);
and U1221 (N_1221,N_1094,N_1002);
or U1222 (N_1222,N_1016,N_1198);
or U1223 (N_1223,N_1190,N_1071);
and U1224 (N_1224,N_1185,N_1084);
and U1225 (N_1225,N_1158,N_1162);
nor U1226 (N_1226,N_1178,N_1006);
xor U1227 (N_1227,N_1135,N_1000);
and U1228 (N_1228,N_1147,N_1113);
nor U1229 (N_1229,N_1056,N_1072);
and U1230 (N_1230,N_1124,N_1096);
or U1231 (N_1231,N_1180,N_1061);
nor U1232 (N_1232,N_1197,N_1177);
nand U1233 (N_1233,N_1103,N_1133);
nor U1234 (N_1234,N_1168,N_1063);
or U1235 (N_1235,N_1013,N_1055);
or U1236 (N_1236,N_1159,N_1121);
or U1237 (N_1237,N_1119,N_1166);
or U1238 (N_1238,N_1123,N_1089);
nand U1239 (N_1239,N_1038,N_1194);
nor U1240 (N_1240,N_1175,N_1154);
nand U1241 (N_1241,N_1191,N_1075);
and U1242 (N_1242,N_1050,N_1052);
nor U1243 (N_1243,N_1007,N_1161);
and U1244 (N_1244,N_1093,N_1025);
nand U1245 (N_1245,N_1145,N_1088);
nand U1246 (N_1246,N_1106,N_1142);
xnor U1247 (N_1247,N_1070,N_1043);
nand U1248 (N_1248,N_1099,N_1044);
or U1249 (N_1249,N_1079,N_1172);
nand U1250 (N_1250,N_1189,N_1112);
or U1251 (N_1251,N_1095,N_1015);
xnor U1252 (N_1252,N_1073,N_1029);
and U1253 (N_1253,N_1195,N_1176);
xnor U1254 (N_1254,N_1125,N_1065);
and U1255 (N_1255,N_1141,N_1010);
nand U1256 (N_1256,N_1024,N_1122);
nand U1257 (N_1257,N_1109,N_1076);
xnor U1258 (N_1258,N_1199,N_1117);
nand U1259 (N_1259,N_1114,N_1081);
and U1260 (N_1260,N_1170,N_1193);
nand U1261 (N_1261,N_1092,N_1128);
nor U1262 (N_1262,N_1156,N_1097);
and U1263 (N_1263,N_1085,N_1188);
nand U1264 (N_1264,N_1080,N_1048);
nand U1265 (N_1265,N_1017,N_1101);
or U1266 (N_1266,N_1134,N_1157);
nor U1267 (N_1267,N_1045,N_1137);
nor U1268 (N_1268,N_1009,N_1127);
nand U1269 (N_1269,N_1160,N_1082);
nand U1270 (N_1270,N_1163,N_1019);
or U1271 (N_1271,N_1181,N_1054);
nand U1272 (N_1272,N_1040,N_1143);
nor U1273 (N_1273,N_1026,N_1041);
nor U1274 (N_1274,N_1078,N_1115);
nor U1275 (N_1275,N_1102,N_1174);
nand U1276 (N_1276,N_1062,N_1046);
xor U1277 (N_1277,N_1083,N_1091);
nand U1278 (N_1278,N_1105,N_1058);
xnor U1279 (N_1279,N_1014,N_1090);
nor U1280 (N_1280,N_1030,N_1118);
nor U1281 (N_1281,N_1012,N_1005);
or U1282 (N_1282,N_1151,N_1153);
or U1283 (N_1283,N_1150,N_1039);
nand U1284 (N_1284,N_1027,N_1051);
and U1285 (N_1285,N_1033,N_1104);
nor U1286 (N_1286,N_1086,N_1171);
or U1287 (N_1287,N_1148,N_1167);
xnor U1288 (N_1288,N_1001,N_1022);
nand U1289 (N_1289,N_1069,N_1187);
nand U1290 (N_1290,N_1179,N_1066);
nand U1291 (N_1291,N_1036,N_1186);
or U1292 (N_1292,N_1047,N_1120);
nor U1293 (N_1293,N_1008,N_1032);
and U1294 (N_1294,N_1111,N_1077);
or U1295 (N_1295,N_1042,N_1100);
nand U1296 (N_1296,N_1132,N_1126);
or U1297 (N_1297,N_1035,N_1108);
xor U1298 (N_1298,N_1116,N_1031);
and U1299 (N_1299,N_1129,N_1183);
nor U1300 (N_1300,N_1161,N_1139);
nor U1301 (N_1301,N_1139,N_1055);
nor U1302 (N_1302,N_1022,N_1170);
nor U1303 (N_1303,N_1002,N_1177);
nor U1304 (N_1304,N_1075,N_1032);
nor U1305 (N_1305,N_1122,N_1084);
and U1306 (N_1306,N_1076,N_1020);
and U1307 (N_1307,N_1165,N_1169);
and U1308 (N_1308,N_1160,N_1093);
nand U1309 (N_1309,N_1121,N_1012);
and U1310 (N_1310,N_1021,N_1166);
nand U1311 (N_1311,N_1120,N_1185);
nand U1312 (N_1312,N_1029,N_1154);
and U1313 (N_1313,N_1156,N_1061);
and U1314 (N_1314,N_1145,N_1044);
and U1315 (N_1315,N_1069,N_1084);
nor U1316 (N_1316,N_1142,N_1090);
and U1317 (N_1317,N_1183,N_1169);
and U1318 (N_1318,N_1141,N_1036);
nand U1319 (N_1319,N_1086,N_1013);
or U1320 (N_1320,N_1178,N_1030);
nor U1321 (N_1321,N_1112,N_1089);
nor U1322 (N_1322,N_1113,N_1177);
or U1323 (N_1323,N_1087,N_1069);
and U1324 (N_1324,N_1178,N_1161);
nand U1325 (N_1325,N_1063,N_1012);
xor U1326 (N_1326,N_1091,N_1159);
nand U1327 (N_1327,N_1101,N_1029);
or U1328 (N_1328,N_1198,N_1028);
or U1329 (N_1329,N_1155,N_1096);
nor U1330 (N_1330,N_1113,N_1050);
xnor U1331 (N_1331,N_1179,N_1115);
nand U1332 (N_1332,N_1005,N_1171);
and U1333 (N_1333,N_1015,N_1166);
and U1334 (N_1334,N_1098,N_1112);
or U1335 (N_1335,N_1054,N_1065);
and U1336 (N_1336,N_1183,N_1038);
or U1337 (N_1337,N_1177,N_1119);
nand U1338 (N_1338,N_1004,N_1018);
xnor U1339 (N_1339,N_1098,N_1080);
nand U1340 (N_1340,N_1074,N_1091);
or U1341 (N_1341,N_1076,N_1166);
xor U1342 (N_1342,N_1045,N_1126);
nor U1343 (N_1343,N_1111,N_1010);
or U1344 (N_1344,N_1194,N_1024);
nand U1345 (N_1345,N_1030,N_1095);
nor U1346 (N_1346,N_1163,N_1143);
nor U1347 (N_1347,N_1040,N_1072);
or U1348 (N_1348,N_1080,N_1197);
and U1349 (N_1349,N_1077,N_1070);
xor U1350 (N_1350,N_1181,N_1108);
nor U1351 (N_1351,N_1164,N_1006);
or U1352 (N_1352,N_1164,N_1016);
or U1353 (N_1353,N_1155,N_1157);
or U1354 (N_1354,N_1106,N_1074);
or U1355 (N_1355,N_1071,N_1083);
nor U1356 (N_1356,N_1125,N_1168);
nand U1357 (N_1357,N_1166,N_1118);
nand U1358 (N_1358,N_1086,N_1000);
nand U1359 (N_1359,N_1185,N_1050);
or U1360 (N_1360,N_1187,N_1140);
xor U1361 (N_1361,N_1145,N_1006);
and U1362 (N_1362,N_1076,N_1139);
xnor U1363 (N_1363,N_1054,N_1157);
or U1364 (N_1364,N_1088,N_1127);
nand U1365 (N_1365,N_1053,N_1103);
nand U1366 (N_1366,N_1146,N_1102);
nand U1367 (N_1367,N_1152,N_1134);
and U1368 (N_1368,N_1031,N_1091);
and U1369 (N_1369,N_1150,N_1107);
and U1370 (N_1370,N_1043,N_1010);
and U1371 (N_1371,N_1091,N_1059);
nor U1372 (N_1372,N_1105,N_1118);
nand U1373 (N_1373,N_1013,N_1083);
nand U1374 (N_1374,N_1169,N_1171);
or U1375 (N_1375,N_1116,N_1012);
nand U1376 (N_1376,N_1077,N_1113);
xnor U1377 (N_1377,N_1191,N_1133);
nor U1378 (N_1378,N_1012,N_1177);
and U1379 (N_1379,N_1196,N_1031);
nor U1380 (N_1380,N_1074,N_1075);
nand U1381 (N_1381,N_1164,N_1059);
and U1382 (N_1382,N_1136,N_1191);
nor U1383 (N_1383,N_1022,N_1008);
xnor U1384 (N_1384,N_1143,N_1017);
xor U1385 (N_1385,N_1046,N_1041);
or U1386 (N_1386,N_1071,N_1088);
nand U1387 (N_1387,N_1168,N_1059);
nor U1388 (N_1388,N_1134,N_1008);
nor U1389 (N_1389,N_1015,N_1115);
nor U1390 (N_1390,N_1064,N_1067);
or U1391 (N_1391,N_1176,N_1090);
nor U1392 (N_1392,N_1153,N_1102);
or U1393 (N_1393,N_1019,N_1161);
nor U1394 (N_1394,N_1181,N_1143);
nand U1395 (N_1395,N_1056,N_1089);
or U1396 (N_1396,N_1157,N_1069);
and U1397 (N_1397,N_1133,N_1150);
nand U1398 (N_1398,N_1097,N_1143);
and U1399 (N_1399,N_1136,N_1074);
nand U1400 (N_1400,N_1261,N_1255);
nand U1401 (N_1401,N_1364,N_1387);
nand U1402 (N_1402,N_1292,N_1313);
and U1403 (N_1403,N_1333,N_1293);
xor U1404 (N_1404,N_1286,N_1268);
or U1405 (N_1405,N_1350,N_1340);
or U1406 (N_1406,N_1221,N_1385);
nand U1407 (N_1407,N_1234,N_1212);
and U1408 (N_1408,N_1321,N_1303);
nor U1409 (N_1409,N_1258,N_1297);
nor U1410 (N_1410,N_1307,N_1248);
xnor U1411 (N_1411,N_1371,N_1305);
nor U1412 (N_1412,N_1356,N_1281);
and U1413 (N_1413,N_1344,N_1322);
nand U1414 (N_1414,N_1289,N_1260);
nor U1415 (N_1415,N_1275,N_1361);
or U1416 (N_1416,N_1218,N_1397);
nor U1417 (N_1417,N_1208,N_1232);
nor U1418 (N_1418,N_1314,N_1379);
or U1419 (N_1419,N_1369,N_1388);
and U1420 (N_1420,N_1376,N_1374);
and U1421 (N_1421,N_1246,N_1296);
nand U1422 (N_1422,N_1318,N_1342);
nand U1423 (N_1423,N_1392,N_1247);
or U1424 (N_1424,N_1316,N_1213);
nand U1425 (N_1425,N_1299,N_1337);
nor U1426 (N_1426,N_1216,N_1271);
xnor U1427 (N_1427,N_1223,N_1290);
and U1428 (N_1428,N_1256,N_1396);
or U1429 (N_1429,N_1257,N_1346);
nor U1430 (N_1430,N_1205,N_1252);
nor U1431 (N_1431,N_1390,N_1381);
nor U1432 (N_1432,N_1354,N_1304);
and U1433 (N_1433,N_1224,N_1311);
nand U1434 (N_1434,N_1283,N_1238);
and U1435 (N_1435,N_1329,N_1382);
or U1436 (N_1436,N_1211,N_1291);
nor U1437 (N_1437,N_1222,N_1267);
nand U1438 (N_1438,N_1345,N_1215);
nand U1439 (N_1439,N_1207,N_1393);
nor U1440 (N_1440,N_1373,N_1270);
nand U1441 (N_1441,N_1230,N_1209);
nand U1442 (N_1442,N_1349,N_1236);
nor U1443 (N_1443,N_1328,N_1279);
nor U1444 (N_1444,N_1284,N_1242);
nor U1445 (N_1445,N_1310,N_1324);
nor U1446 (N_1446,N_1365,N_1214);
or U1447 (N_1447,N_1368,N_1278);
nand U1448 (N_1448,N_1227,N_1272);
and U1449 (N_1449,N_1332,N_1228);
or U1450 (N_1450,N_1210,N_1308);
and U1451 (N_1451,N_1338,N_1217);
nand U1452 (N_1452,N_1363,N_1399);
nor U1453 (N_1453,N_1398,N_1306);
nor U1454 (N_1454,N_1352,N_1288);
or U1455 (N_1455,N_1203,N_1249);
nor U1456 (N_1456,N_1335,N_1285);
xor U1457 (N_1457,N_1300,N_1395);
nor U1458 (N_1458,N_1383,N_1367);
or U1459 (N_1459,N_1315,N_1355);
nor U1460 (N_1460,N_1341,N_1384);
nand U1461 (N_1461,N_1378,N_1343);
and U1462 (N_1462,N_1231,N_1309);
nand U1463 (N_1463,N_1351,N_1263);
or U1464 (N_1464,N_1240,N_1294);
and U1465 (N_1465,N_1370,N_1282);
nand U1466 (N_1466,N_1394,N_1253);
nor U1467 (N_1467,N_1233,N_1273);
or U1468 (N_1468,N_1301,N_1220);
or U1469 (N_1469,N_1204,N_1317);
nand U1470 (N_1470,N_1280,N_1359);
or U1471 (N_1471,N_1225,N_1386);
or U1472 (N_1472,N_1375,N_1243);
or U1473 (N_1473,N_1254,N_1295);
or U1474 (N_1474,N_1330,N_1325);
nand U1475 (N_1475,N_1250,N_1353);
and U1476 (N_1476,N_1274,N_1235);
xnor U1477 (N_1477,N_1262,N_1219);
nor U1478 (N_1478,N_1200,N_1360);
or U1479 (N_1479,N_1287,N_1362);
and U1480 (N_1480,N_1347,N_1276);
nor U1481 (N_1481,N_1251,N_1323);
and U1482 (N_1482,N_1244,N_1201);
nor U1483 (N_1483,N_1265,N_1326);
nand U1484 (N_1484,N_1339,N_1320);
nor U1485 (N_1485,N_1259,N_1380);
and U1486 (N_1486,N_1372,N_1269);
nand U1487 (N_1487,N_1245,N_1319);
xnor U1488 (N_1488,N_1266,N_1298);
nand U1489 (N_1489,N_1366,N_1237);
and U1490 (N_1490,N_1312,N_1336);
nand U1491 (N_1491,N_1327,N_1239);
nor U1492 (N_1492,N_1357,N_1334);
nand U1493 (N_1493,N_1391,N_1302);
nand U1494 (N_1494,N_1202,N_1277);
nand U1495 (N_1495,N_1206,N_1241);
or U1496 (N_1496,N_1348,N_1264);
nand U1497 (N_1497,N_1389,N_1377);
and U1498 (N_1498,N_1331,N_1358);
nand U1499 (N_1499,N_1229,N_1226);
and U1500 (N_1500,N_1251,N_1364);
or U1501 (N_1501,N_1217,N_1229);
nor U1502 (N_1502,N_1252,N_1272);
nand U1503 (N_1503,N_1363,N_1240);
xnor U1504 (N_1504,N_1309,N_1292);
nor U1505 (N_1505,N_1292,N_1257);
or U1506 (N_1506,N_1391,N_1332);
and U1507 (N_1507,N_1322,N_1219);
and U1508 (N_1508,N_1251,N_1305);
nand U1509 (N_1509,N_1283,N_1310);
nor U1510 (N_1510,N_1277,N_1251);
or U1511 (N_1511,N_1290,N_1349);
xor U1512 (N_1512,N_1285,N_1266);
and U1513 (N_1513,N_1377,N_1372);
nor U1514 (N_1514,N_1381,N_1217);
nand U1515 (N_1515,N_1225,N_1206);
and U1516 (N_1516,N_1334,N_1208);
xnor U1517 (N_1517,N_1261,N_1221);
nor U1518 (N_1518,N_1292,N_1265);
xor U1519 (N_1519,N_1324,N_1290);
or U1520 (N_1520,N_1390,N_1324);
and U1521 (N_1521,N_1216,N_1215);
nor U1522 (N_1522,N_1288,N_1327);
nand U1523 (N_1523,N_1327,N_1393);
nor U1524 (N_1524,N_1373,N_1252);
and U1525 (N_1525,N_1280,N_1312);
nor U1526 (N_1526,N_1247,N_1244);
xnor U1527 (N_1527,N_1270,N_1204);
xor U1528 (N_1528,N_1268,N_1322);
and U1529 (N_1529,N_1297,N_1271);
nand U1530 (N_1530,N_1363,N_1246);
or U1531 (N_1531,N_1330,N_1336);
or U1532 (N_1532,N_1360,N_1324);
or U1533 (N_1533,N_1295,N_1314);
nor U1534 (N_1534,N_1357,N_1245);
and U1535 (N_1535,N_1349,N_1263);
nor U1536 (N_1536,N_1316,N_1216);
nand U1537 (N_1537,N_1217,N_1357);
or U1538 (N_1538,N_1391,N_1290);
or U1539 (N_1539,N_1247,N_1313);
nor U1540 (N_1540,N_1259,N_1324);
nor U1541 (N_1541,N_1270,N_1223);
and U1542 (N_1542,N_1256,N_1296);
nand U1543 (N_1543,N_1301,N_1364);
or U1544 (N_1544,N_1341,N_1216);
nand U1545 (N_1545,N_1324,N_1399);
or U1546 (N_1546,N_1373,N_1382);
nand U1547 (N_1547,N_1253,N_1295);
xor U1548 (N_1548,N_1370,N_1327);
or U1549 (N_1549,N_1378,N_1286);
nand U1550 (N_1550,N_1282,N_1362);
nand U1551 (N_1551,N_1310,N_1378);
nand U1552 (N_1552,N_1275,N_1201);
nor U1553 (N_1553,N_1258,N_1226);
nor U1554 (N_1554,N_1382,N_1300);
or U1555 (N_1555,N_1308,N_1203);
or U1556 (N_1556,N_1312,N_1206);
or U1557 (N_1557,N_1314,N_1240);
nand U1558 (N_1558,N_1209,N_1274);
and U1559 (N_1559,N_1220,N_1252);
xnor U1560 (N_1560,N_1263,N_1269);
xor U1561 (N_1561,N_1362,N_1213);
or U1562 (N_1562,N_1333,N_1393);
xnor U1563 (N_1563,N_1339,N_1374);
or U1564 (N_1564,N_1252,N_1256);
nand U1565 (N_1565,N_1332,N_1239);
nor U1566 (N_1566,N_1382,N_1244);
xnor U1567 (N_1567,N_1254,N_1387);
nor U1568 (N_1568,N_1368,N_1234);
nand U1569 (N_1569,N_1206,N_1242);
nor U1570 (N_1570,N_1203,N_1355);
and U1571 (N_1571,N_1383,N_1363);
and U1572 (N_1572,N_1398,N_1279);
xnor U1573 (N_1573,N_1302,N_1260);
nand U1574 (N_1574,N_1332,N_1388);
nor U1575 (N_1575,N_1333,N_1244);
and U1576 (N_1576,N_1234,N_1356);
and U1577 (N_1577,N_1366,N_1277);
nand U1578 (N_1578,N_1284,N_1329);
nor U1579 (N_1579,N_1270,N_1210);
and U1580 (N_1580,N_1314,N_1311);
xnor U1581 (N_1581,N_1357,N_1361);
or U1582 (N_1582,N_1282,N_1391);
and U1583 (N_1583,N_1297,N_1265);
nor U1584 (N_1584,N_1305,N_1341);
nand U1585 (N_1585,N_1376,N_1292);
or U1586 (N_1586,N_1281,N_1213);
nor U1587 (N_1587,N_1301,N_1385);
or U1588 (N_1588,N_1294,N_1277);
xnor U1589 (N_1589,N_1342,N_1301);
nand U1590 (N_1590,N_1325,N_1276);
or U1591 (N_1591,N_1201,N_1339);
or U1592 (N_1592,N_1279,N_1309);
xnor U1593 (N_1593,N_1352,N_1255);
or U1594 (N_1594,N_1322,N_1220);
nor U1595 (N_1595,N_1377,N_1276);
and U1596 (N_1596,N_1263,N_1353);
nor U1597 (N_1597,N_1291,N_1252);
or U1598 (N_1598,N_1203,N_1302);
and U1599 (N_1599,N_1301,N_1288);
nand U1600 (N_1600,N_1565,N_1406);
and U1601 (N_1601,N_1518,N_1481);
nor U1602 (N_1602,N_1497,N_1460);
or U1603 (N_1603,N_1472,N_1485);
nor U1604 (N_1604,N_1514,N_1520);
and U1605 (N_1605,N_1525,N_1567);
or U1606 (N_1606,N_1405,N_1552);
or U1607 (N_1607,N_1457,N_1486);
and U1608 (N_1608,N_1444,N_1451);
and U1609 (N_1609,N_1473,N_1404);
or U1610 (N_1610,N_1575,N_1478);
nor U1611 (N_1611,N_1534,N_1449);
and U1612 (N_1612,N_1423,N_1415);
nor U1613 (N_1613,N_1438,N_1401);
nor U1614 (N_1614,N_1560,N_1566);
nand U1615 (N_1615,N_1557,N_1586);
or U1616 (N_1616,N_1471,N_1576);
and U1617 (N_1617,N_1524,N_1435);
and U1618 (N_1618,N_1446,N_1452);
nor U1619 (N_1619,N_1490,N_1458);
or U1620 (N_1620,N_1550,N_1419);
or U1621 (N_1621,N_1407,N_1500);
nor U1622 (N_1622,N_1496,N_1441);
and U1623 (N_1623,N_1558,N_1453);
nor U1624 (N_1624,N_1426,N_1541);
and U1625 (N_1625,N_1439,N_1516);
nand U1626 (N_1626,N_1455,N_1521);
nand U1627 (N_1627,N_1440,N_1469);
or U1628 (N_1628,N_1542,N_1544);
nor U1629 (N_1629,N_1425,N_1561);
nand U1630 (N_1630,N_1433,N_1450);
nor U1631 (N_1631,N_1447,N_1579);
or U1632 (N_1632,N_1463,N_1408);
nor U1633 (N_1633,N_1417,N_1492);
nor U1634 (N_1634,N_1437,N_1411);
and U1635 (N_1635,N_1597,N_1555);
nand U1636 (N_1636,N_1410,N_1584);
xor U1637 (N_1637,N_1547,N_1533);
xor U1638 (N_1638,N_1468,N_1580);
nor U1639 (N_1639,N_1470,N_1505);
and U1640 (N_1640,N_1531,N_1454);
nand U1641 (N_1641,N_1545,N_1409);
nor U1642 (N_1642,N_1413,N_1416);
and U1643 (N_1643,N_1599,N_1480);
nor U1644 (N_1644,N_1491,N_1475);
or U1645 (N_1645,N_1598,N_1503);
nor U1646 (N_1646,N_1403,N_1515);
nand U1647 (N_1647,N_1588,N_1402);
nor U1648 (N_1648,N_1569,N_1556);
and U1649 (N_1649,N_1522,N_1495);
and U1650 (N_1650,N_1592,N_1498);
nand U1651 (N_1651,N_1467,N_1517);
or U1652 (N_1652,N_1590,N_1532);
or U1653 (N_1653,N_1448,N_1511);
and U1654 (N_1654,N_1523,N_1519);
or U1655 (N_1655,N_1459,N_1583);
and U1656 (N_1656,N_1512,N_1593);
nor U1657 (N_1657,N_1477,N_1504);
and U1658 (N_1658,N_1553,N_1424);
xnor U1659 (N_1659,N_1581,N_1429);
nor U1660 (N_1660,N_1479,N_1539);
or U1661 (N_1661,N_1594,N_1587);
nand U1662 (N_1662,N_1529,N_1549);
xnor U1663 (N_1663,N_1526,N_1510);
nor U1664 (N_1664,N_1559,N_1595);
and U1665 (N_1665,N_1442,N_1564);
nor U1666 (N_1666,N_1571,N_1421);
or U1667 (N_1667,N_1573,N_1422);
nor U1668 (N_1668,N_1456,N_1585);
or U1669 (N_1669,N_1483,N_1513);
nand U1670 (N_1670,N_1551,N_1431);
nor U1671 (N_1671,N_1543,N_1436);
and U1672 (N_1672,N_1418,N_1484);
nor U1673 (N_1673,N_1506,N_1420);
or U1674 (N_1674,N_1465,N_1482);
nor U1675 (N_1675,N_1537,N_1570);
nor U1676 (N_1676,N_1502,N_1412);
and U1677 (N_1677,N_1428,N_1489);
or U1678 (N_1678,N_1493,N_1462);
and U1679 (N_1679,N_1499,N_1572);
and U1680 (N_1680,N_1574,N_1427);
xor U1681 (N_1681,N_1414,N_1535);
nor U1682 (N_1682,N_1554,N_1563);
and U1683 (N_1683,N_1536,N_1548);
nor U1684 (N_1684,N_1445,N_1434);
or U1685 (N_1685,N_1400,N_1430);
or U1686 (N_1686,N_1527,N_1568);
nor U1687 (N_1687,N_1466,N_1507);
and U1688 (N_1688,N_1596,N_1509);
and U1689 (N_1689,N_1432,N_1464);
nor U1690 (N_1690,N_1487,N_1474);
nand U1691 (N_1691,N_1530,N_1461);
nand U1692 (N_1692,N_1501,N_1578);
nand U1693 (N_1693,N_1528,N_1443);
nand U1694 (N_1694,N_1591,N_1577);
and U1695 (N_1695,N_1589,N_1582);
and U1696 (N_1696,N_1476,N_1538);
nor U1697 (N_1697,N_1540,N_1494);
xnor U1698 (N_1698,N_1562,N_1488);
nand U1699 (N_1699,N_1508,N_1546);
nand U1700 (N_1700,N_1422,N_1421);
nor U1701 (N_1701,N_1518,N_1598);
or U1702 (N_1702,N_1505,N_1458);
nand U1703 (N_1703,N_1525,N_1591);
nor U1704 (N_1704,N_1550,N_1569);
nor U1705 (N_1705,N_1566,N_1451);
or U1706 (N_1706,N_1597,N_1514);
or U1707 (N_1707,N_1525,N_1502);
nor U1708 (N_1708,N_1466,N_1412);
nand U1709 (N_1709,N_1460,N_1510);
nor U1710 (N_1710,N_1446,N_1541);
nand U1711 (N_1711,N_1539,N_1410);
or U1712 (N_1712,N_1441,N_1480);
nor U1713 (N_1713,N_1499,N_1598);
and U1714 (N_1714,N_1512,N_1544);
nor U1715 (N_1715,N_1552,N_1454);
or U1716 (N_1716,N_1575,N_1492);
nor U1717 (N_1717,N_1400,N_1448);
and U1718 (N_1718,N_1549,N_1562);
nand U1719 (N_1719,N_1573,N_1435);
nor U1720 (N_1720,N_1451,N_1484);
and U1721 (N_1721,N_1494,N_1476);
xor U1722 (N_1722,N_1498,N_1417);
and U1723 (N_1723,N_1526,N_1482);
xor U1724 (N_1724,N_1406,N_1589);
nand U1725 (N_1725,N_1430,N_1570);
or U1726 (N_1726,N_1412,N_1569);
nand U1727 (N_1727,N_1487,N_1593);
xor U1728 (N_1728,N_1570,N_1567);
nor U1729 (N_1729,N_1439,N_1465);
or U1730 (N_1730,N_1408,N_1592);
or U1731 (N_1731,N_1565,N_1589);
nand U1732 (N_1732,N_1555,N_1504);
nand U1733 (N_1733,N_1400,N_1471);
xnor U1734 (N_1734,N_1599,N_1434);
and U1735 (N_1735,N_1578,N_1590);
or U1736 (N_1736,N_1404,N_1538);
xnor U1737 (N_1737,N_1530,N_1432);
and U1738 (N_1738,N_1533,N_1565);
nor U1739 (N_1739,N_1474,N_1496);
nor U1740 (N_1740,N_1564,N_1401);
and U1741 (N_1741,N_1495,N_1488);
nand U1742 (N_1742,N_1558,N_1500);
or U1743 (N_1743,N_1456,N_1508);
nand U1744 (N_1744,N_1475,N_1409);
or U1745 (N_1745,N_1496,N_1492);
or U1746 (N_1746,N_1552,N_1449);
and U1747 (N_1747,N_1448,N_1532);
xnor U1748 (N_1748,N_1572,N_1566);
nor U1749 (N_1749,N_1519,N_1597);
nand U1750 (N_1750,N_1504,N_1503);
or U1751 (N_1751,N_1576,N_1479);
nand U1752 (N_1752,N_1497,N_1440);
nor U1753 (N_1753,N_1404,N_1483);
nor U1754 (N_1754,N_1523,N_1481);
and U1755 (N_1755,N_1520,N_1526);
nor U1756 (N_1756,N_1411,N_1577);
and U1757 (N_1757,N_1438,N_1521);
nand U1758 (N_1758,N_1479,N_1536);
nand U1759 (N_1759,N_1535,N_1498);
or U1760 (N_1760,N_1573,N_1412);
or U1761 (N_1761,N_1599,N_1447);
nor U1762 (N_1762,N_1473,N_1489);
nand U1763 (N_1763,N_1414,N_1402);
and U1764 (N_1764,N_1528,N_1447);
or U1765 (N_1765,N_1413,N_1526);
nor U1766 (N_1766,N_1544,N_1458);
or U1767 (N_1767,N_1546,N_1543);
nand U1768 (N_1768,N_1422,N_1597);
nor U1769 (N_1769,N_1589,N_1407);
or U1770 (N_1770,N_1528,N_1503);
nand U1771 (N_1771,N_1576,N_1469);
and U1772 (N_1772,N_1452,N_1413);
or U1773 (N_1773,N_1454,N_1562);
nand U1774 (N_1774,N_1528,N_1544);
or U1775 (N_1775,N_1455,N_1475);
or U1776 (N_1776,N_1403,N_1462);
or U1777 (N_1777,N_1516,N_1406);
and U1778 (N_1778,N_1441,N_1439);
nand U1779 (N_1779,N_1480,N_1592);
and U1780 (N_1780,N_1408,N_1596);
nor U1781 (N_1781,N_1577,N_1401);
or U1782 (N_1782,N_1485,N_1591);
nand U1783 (N_1783,N_1479,N_1480);
and U1784 (N_1784,N_1528,N_1498);
xnor U1785 (N_1785,N_1501,N_1573);
nand U1786 (N_1786,N_1491,N_1568);
nand U1787 (N_1787,N_1558,N_1530);
xor U1788 (N_1788,N_1444,N_1421);
nand U1789 (N_1789,N_1423,N_1566);
nand U1790 (N_1790,N_1420,N_1427);
or U1791 (N_1791,N_1434,N_1556);
xnor U1792 (N_1792,N_1427,N_1493);
nand U1793 (N_1793,N_1497,N_1539);
and U1794 (N_1794,N_1446,N_1561);
nand U1795 (N_1795,N_1464,N_1487);
and U1796 (N_1796,N_1597,N_1490);
or U1797 (N_1797,N_1575,N_1570);
nor U1798 (N_1798,N_1473,N_1537);
or U1799 (N_1799,N_1533,N_1575);
nor U1800 (N_1800,N_1745,N_1788);
or U1801 (N_1801,N_1692,N_1611);
or U1802 (N_1802,N_1701,N_1703);
nor U1803 (N_1803,N_1707,N_1766);
and U1804 (N_1804,N_1624,N_1674);
and U1805 (N_1805,N_1776,N_1778);
and U1806 (N_1806,N_1730,N_1774);
nor U1807 (N_1807,N_1762,N_1601);
or U1808 (N_1808,N_1648,N_1608);
or U1809 (N_1809,N_1772,N_1631);
nand U1810 (N_1810,N_1653,N_1609);
xnor U1811 (N_1811,N_1708,N_1717);
and U1812 (N_1812,N_1647,N_1635);
nand U1813 (N_1813,N_1736,N_1729);
nor U1814 (N_1814,N_1628,N_1740);
and U1815 (N_1815,N_1682,N_1790);
nand U1816 (N_1816,N_1769,N_1709);
nand U1817 (N_1817,N_1605,N_1799);
and U1818 (N_1818,N_1721,N_1699);
and U1819 (N_1819,N_1765,N_1786);
nand U1820 (N_1820,N_1650,N_1691);
nand U1821 (N_1821,N_1673,N_1646);
or U1822 (N_1822,N_1723,N_1632);
xor U1823 (N_1823,N_1775,N_1695);
or U1824 (N_1824,N_1770,N_1606);
nand U1825 (N_1825,N_1602,N_1696);
xnor U1826 (N_1826,N_1731,N_1755);
nand U1827 (N_1827,N_1649,N_1704);
and U1828 (N_1828,N_1621,N_1686);
nor U1829 (N_1829,N_1796,N_1616);
nand U1830 (N_1830,N_1771,N_1715);
nand U1831 (N_1831,N_1760,N_1728);
and U1832 (N_1832,N_1764,N_1603);
xor U1833 (N_1833,N_1694,N_1720);
and U1834 (N_1834,N_1678,N_1787);
nor U1835 (N_1835,N_1685,N_1664);
nand U1836 (N_1836,N_1761,N_1743);
and U1837 (N_1837,N_1798,N_1744);
nand U1838 (N_1838,N_1725,N_1718);
nor U1839 (N_1839,N_1711,N_1697);
nand U1840 (N_1840,N_1722,N_1633);
nor U1841 (N_1841,N_1733,N_1756);
xor U1842 (N_1842,N_1794,N_1612);
or U1843 (N_1843,N_1660,N_1658);
or U1844 (N_1844,N_1767,N_1714);
xor U1845 (N_1845,N_1746,N_1702);
nand U1846 (N_1846,N_1637,N_1629);
and U1847 (N_1847,N_1615,N_1610);
or U1848 (N_1848,N_1689,N_1656);
nand U1849 (N_1849,N_1747,N_1669);
and U1850 (N_1850,N_1706,N_1681);
nor U1851 (N_1851,N_1789,N_1644);
nor U1852 (N_1852,N_1661,N_1734);
xnor U1853 (N_1853,N_1600,N_1748);
xnor U1854 (N_1854,N_1690,N_1780);
and U1855 (N_1855,N_1652,N_1665);
nand U1856 (N_1856,N_1655,N_1750);
or U1857 (N_1857,N_1677,N_1642);
and U1858 (N_1858,N_1751,N_1659);
or U1859 (N_1859,N_1687,N_1670);
nand U1860 (N_1860,N_1630,N_1618);
and U1861 (N_1861,N_1698,N_1613);
nand U1862 (N_1862,N_1742,N_1738);
and U1863 (N_1863,N_1741,N_1791);
xor U1864 (N_1864,N_1634,N_1724);
and U1865 (N_1865,N_1727,N_1607);
or U1866 (N_1866,N_1758,N_1754);
nand U1867 (N_1867,N_1620,N_1795);
and U1868 (N_1868,N_1749,N_1623);
nand U1869 (N_1869,N_1777,N_1732);
and U1870 (N_1870,N_1739,N_1638);
nand U1871 (N_1871,N_1683,N_1693);
or U1872 (N_1872,N_1710,N_1713);
nand U1873 (N_1873,N_1640,N_1622);
or U1874 (N_1874,N_1700,N_1625);
nand U1875 (N_1875,N_1792,N_1712);
and U1876 (N_1876,N_1757,N_1737);
and U1877 (N_1877,N_1735,N_1654);
or U1878 (N_1878,N_1705,N_1641);
nand U1879 (N_1879,N_1657,N_1667);
nor U1880 (N_1880,N_1784,N_1783);
or U1881 (N_1881,N_1753,N_1679);
nand U1882 (N_1882,N_1604,N_1626);
and U1883 (N_1883,N_1636,N_1651);
nor U1884 (N_1884,N_1773,N_1719);
and U1885 (N_1885,N_1763,N_1688);
xnor U1886 (N_1886,N_1619,N_1617);
nand U1887 (N_1887,N_1662,N_1779);
and U1888 (N_1888,N_1645,N_1793);
and U1889 (N_1889,N_1666,N_1759);
and U1890 (N_1890,N_1627,N_1614);
and U1891 (N_1891,N_1781,N_1663);
nor U1892 (N_1892,N_1672,N_1675);
nand U1893 (N_1893,N_1726,N_1684);
or U1894 (N_1894,N_1671,N_1785);
nor U1895 (N_1895,N_1643,N_1752);
and U1896 (N_1896,N_1676,N_1680);
or U1897 (N_1897,N_1639,N_1797);
nor U1898 (N_1898,N_1716,N_1782);
or U1899 (N_1899,N_1768,N_1668);
nand U1900 (N_1900,N_1669,N_1703);
or U1901 (N_1901,N_1643,N_1637);
nand U1902 (N_1902,N_1777,N_1680);
nor U1903 (N_1903,N_1686,N_1663);
nand U1904 (N_1904,N_1614,N_1721);
nand U1905 (N_1905,N_1649,N_1770);
and U1906 (N_1906,N_1792,N_1785);
or U1907 (N_1907,N_1755,N_1796);
nor U1908 (N_1908,N_1766,N_1726);
nand U1909 (N_1909,N_1644,N_1799);
or U1910 (N_1910,N_1704,N_1719);
nand U1911 (N_1911,N_1601,N_1644);
nand U1912 (N_1912,N_1750,N_1638);
and U1913 (N_1913,N_1739,N_1662);
and U1914 (N_1914,N_1711,N_1779);
or U1915 (N_1915,N_1769,N_1648);
and U1916 (N_1916,N_1705,N_1627);
and U1917 (N_1917,N_1799,N_1658);
or U1918 (N_1918,N_1795,N_1745);
and U1919 (N_1919,N_1793,N_1740);
or U1920 (N_1920,N_1723,N_1627);
nor U1921 (N_1921,N_1714,N_1695);
or U1922 (N_1922,N_1744,N_1737);
and U1923 (N_1923,N_1685,N_1765);
nor U1924 (N_1924,N_1733,N_1766);
xor U1925 (N_1925,N_1754,N_1639);
nand U1926 (N_1926,N_1686,N_1797);
and U1927 (N_1927,N_1702,N_1798);
xnor U1928 (N_1928,N_1718,N_1772);
or U1929 (N_1929,N_1713,N_1695);
xor U1930 (N_1930,N_1770,N_1600);
nor U1931 (N_1931,N_1771,N_1665);
and U1932 (N_1932,N_1762,N_1659);
nand U1933 (N_1933,N_1749,N_1744);
or U1934 (N_1934,N_1793,N_1630);
nand U1935 (N_1935,N_1765,N_1770);
and U1936 (N_1936,N_1711,N_1647);
nand U1937 (N_1937,N_1773,N_1635);
or U1938 (N_1938,N_1627,N_1601);
nand U1939 (N_1939,N_1794,N_1628);
nor U1940 (N_1940,N_1715,N_1761);
nand U1941 (N_1941,N_1750,N_1789);
nor U1942 (N_1942,N_1663,N_1713);
and U1943 (N_1943,N_1712,N_1708);
nand U1944 (N_1944,N_1739,N_1763);
or U1945 (N_1945,N_1610,N_1776);
or U1946 (N_1946,N_1678,N_1704);
and U1947 (N_1947,N_1708,N_1791);
nand U1948 (N_1948,N_1631,N_1683);
and U1949 (N_1949,N_1629,N_1739);
and U1950 (N_1950,N_1633,N_1649);
nor U1951 (N_1951,N_1720,N_1659);
xor U1952 (N_1952,N_1619,N_1701);
or U1953 (N_1953,N_1702,N_1683);
nor U1954 (N_1954,N_1699,N_1621);
nor U1955 (N_1955,N_1725,N_1717);
nand U1956 (N_1956,N_1695,N_1783);
or U1957 (N_1957,N_1766,N_1611);
and U1958 (N_1958,N_1781,N_1782);
or U1959 (N_1959,N_1619,N_1789);
xnor U1960 (N_1960,N_1628,N_1609);
xnor U1961 (N_1961,N_1713,N_1765);
nor U1962 (N_1962,N_1769,N_1757);
nand U1963 (N_1963,N_1692,N_1641);
nor U1964 (N_1964,N_1699,N_1665);
or U1965 (N_1965,N_1745,N_1612);
nor U1966 (N_1966,N_1789,N_1689);
xnor U1967 (N_1967,N_1729,N_1767);
and U1968 (N_1968,N_1740,N_1703);
or U1969 (N_1969,N_1633,N_1715);
nor U1970 (N_1970,N_1616,N_1726);
nand U1971 (N_1971,N_1704,N_1632);
xnor U1972 (N_1972,N_1768,N_1605);
and U1973 (N_1973,N_1617,N_1643);
or U1974 (N_1974,N_1680,N_1668);
nand U1975 (N_1975,N_1781,N_1699);
and U1976 (N_1976,N_1723,N_1733);
and U1977 (N_1977,N_1786,N_1683);
and U1978 (N_1978,N_1653,N_1720);
and U1979 (N_1979,N_1654,N_1625);
or U1980 (N_1980,N_1760,N_1655);
nor U1981 (N_1981,N_1767,N_1755);
nand U1982 (N_1982,N_1602,N_1720);
nand U1983 (N_1983,N_1777,N_1617);
and U1984 (N_1984,N_1798,N_1780);
nor U1985 (N_1985,N_1795,N_1727);
and U1986 (N_1986,N_1798,N_1669);
and U1987 (N_1987,N_1770,N_1720);
and U1988 (N_1988,N_1681,N_1766);
or U1989 (N_1989,N_1662,N_1603);
nor U1990 (N_1990,N_1720,N_1700);
nor U1991 (N_1991,N_1779,N_1699);
and U1992 (N_1992,N_1640,N_1682);
xor U1993 (N_1993,N_1702,N_1614);
xor U1994 (N_1994,N_1691,N_1752);
nand U1995 (N_1995,N_1632,N_1680);
xnor U1996 (N_1996,N_1773,N_1672);
nor U1997 (N_1997,N_1622,N_1647);
xnor U1998 (N_1998,N_1693,N_1731);
nand U1999 (N_1999,N_1688,N_1727);
and U2000 (N_2000,N_1949,N_1817);
nand U2001 (N_2001,N_1819,N_1960);
nand U2002 (N_2002,N_1859,N_1948);
and U2003 (N_2003,N_1847,N_1954);
or U2004 (N_2004,N_1898,N_1882);
nor U2005 (N_2005,N_1923,N_1982);
xnor U2006 (N_2006,N_1976,N_1853);
or U2007 (N_2007,N_1893,N_1897);
nor U2008 (N_2008,N_1955,N_1851);
nand U2009 (N_2009,N_1956,N_1947);
nand U2010 (N_2010,N_1945,N_1998);
xnor U2011 (N_2011,N_1916,N_1848);
and U2012 (N_2012,N_1974,N_1888);
nor U2013 (N_2013,N_1828,N_1852);
nor U2014 (N_2014,N_1878,N_1992);
nor U2015 (N_2015,N_1972,N_1966);
or U2016 (N_2016,N_1810,N_1830);
or U2017 (N_2017,N_1845,N_1806);
nor U2018 (N_2018,N_1889,N_1823);
nor U2019 (N_2019,N_1912,N_1927);
nand U2020 (N_2020,N_1844,N_1909);
nor U2021 (N_2021,N_1862,N_1940);
nor U2022 (N_2022,N_1991,N_1850);
or U2023 (N_2023,N_1822,N_1987);
and U2024 (N_2024,N_1855,N_1812);
nor U2025 (N_2025,N_1809,N_1800);
nand U2026 (N_2026,N_1841,N_1924);
and U2027 (N_2027,N_1928,N_1986);
nand U2028 (N_2028,N_1997,N_1867);
nor U2029 (N_2029,N_1995,N_1894);
or U2030 (N_2030,N_1838,N_1807);
and U2031 (N_2031,N_1890,N_1869);
xor U2032 (N_2032,N_1858,N_1903);
nor U2033 (N_2033,N_1864,N_1939);
nand U2034 (N_2034,N_1994,N_1929);
and U2035 (N_2035,N_1963,N_1876);
and U2036 (N_2036,N_1921,N_1895);
nand U2037 (N_2037,N_1905,N_1971);
nor U2038 (N_2038,N_1846,N_1907);
and U2039 (N_2039,N_1919,N_1832);
xor U2040 (N_2040,N_1826,N_1910);
nor U2041 (N_2041,N_1970,N_1820);
or U2042 (N_2042,N_1829,N_1942);
and U2043 (N_2043,N_1941,N_1854);
and U2044 (N_2044,N_1977,N_1964);
nor U2045 (N_2045,N_1899,N_1989);
nor U2046 (N_2046,N_1926,N_1975);
nor U2047 (N_2047,N_1833,N_1896);
nor U2048 (N_2048,N_1871,N_1886);
and U2049 (N_2049,N_1849,N_1801);
and U2050 (N_2050,N_1865,N_1816);
nand U2051 (N_2051,N_1920,N_1874);
and U2052 (N_2052,N_1868,N_1915);
and U2053 (N_2053,N_1925,N_1873);
nand U2054 (N_2054,N_1825,N_1944);
nand U2055 (N_2055,N_1999,N_1811);
xor U2056 (N_2056,N_1877,N_1946);
and U2057 (N_2057,N_1861,N_1891);
and U2058 (N_2058,N_1880,N_1979);
nor U2059 (N_2059,N_1887,N_1857);
and U2060 (N_2060,N_1802,N_1908);
or U2061 (N_2061,N_1834,N_1978);
xnor U2062 (N_2062,N_1881,N_1917);
and U2063 (N_2063,N_1803,N_1953);
xor U2064 (N_2064,N_1856,N_1937);
nor U2065 (N_2065,N_1892,N_1837);
and U2066 (N_2066,N_1983,N_1879);
nor U2067 (N_2067,N_1981,N_1935);
and U2068 (N_2068,N_1936,N_1813);
and U2069 (N_2069,N_1965,N_1958);
and U2070 (N_2070,N_1918,N_1969);
and U2071 (N_2071,N_1900,N_1815);
and U2072 (N_2072,N_1870,N_1993);
nor U2073 (N_2073,N_1957,N_1885);
nand U2074 (N_2074,N_1950,N_1831);
and U2075 (N_2075,N_1985,N_1914);
and U2076 (N_2076,N_1968,N_1808);
nor U2077 (N_2077,N_1996,N_1906);
nor U2078 (N_2078,N_1824,N_1902);
or U2079 (N_2079,N_1931,N_1943);
or U2080 (N_2080,N_1863,N_1821);
nor U2081 (N_2081,N_1930,N_1990);
nor U2082 (N_2082,N_1952,N_1843);
or U2083 (N_2083,N_1884,N_1840);
nand U2084 (N_2084,N_1805,N_1959);
nor U2085 (N_2085,N_1938,N_1961);
nor U2086 (N_2086,N_1836,N_1866);
nand U2087 (N_2087,N_1973,N_1934);
and U2088 (N_2088,N_1860,N_1883);
and U2089 (N_2089,N_1933,N_1835);
nor U2090 (N_2090,N_1988,N_1842);
and U2091 (N_2091,N_1911,N_1922);
or U2092 (N_2092,N_1932,N_1872);
nor U2093 (N_2093,N_1913,N_1818);
and U2094 (N_2094,N_1804,N_1962);
nor U2095 (N_2095,N_1951,N_1814);
nor U2096 (N_2096,N_1839,N_1980);
and U2097 (N_2097,N_1967,N_1827);
xor U2098 (N_2098,N_1904,N_1984);
and U2099 (N_2099,N_1901,N_1875);
and U2100 (N_2100,N_1901,N_1873);
nand U2101 (N_2101,N_1996,N_1800);
or U2102 (N_2102,N_1923,N_1905);
nand U2103 (N_2103,N_1978,N_1960);
xor U2104 (N_2104,N_1912,N_1869);
nand U2105 (N_2105,N_1861,N_1968);
nand U2106 (N_2106,N_1861,N_1898);
nor U2107 (N_2107,N_1840,N_1819);
or U2108 (N_2108,N_1897,N_1966);
or U2109 (N_2109,N_1992,N_1909);
nor U2110 (N_2110,N_1894,N_1901);
or U2111 (N_2111,N_1922,N_1946);
nor U2112 (N_2112,N_1907,N_1940);
nand U2113 (N_2113,N_1942,N_1879);
nand U2114 (N_2114,N_1997,N_1953);
and U2115 (N_2115,N_1909,N_1954);
or U2116 (N_2116,N_1968,N_1964);
xor U2117 (N_2117,N_1876,N_1823);
nand U2118 (N_2118,N_1907,N_1815);
nor U2119 (N_2119,N_1984,N_1865);
nor U2120 (N_2120,N_1877,N_1904);
and U2121 (N_2121,N_1909,N_1938);
or U2122 (N_2122,N_1821,N_1808);
and U2123 (N_2123,N_1934,N_1878);
and U2124 (N_2124,N_1877,N_1924);
nand U2125 (N_2125,N_1968,N_1887);
nand U2126 (N_2126,N_1949,N_1955);
nand U2127 (N_2127,N_1919,N_1826);
and U2128 (N_2128,N_1992,N_1974);
xor U2129 (N_2129,N_1949,N_1822);
nor U2130 (N_2130,N_1980,N_1921);
and U2131 (N_2131,N_1833,N_1959);
nor U2132 (N_2132,N_1837,N_1804);
and U2133 (N_2133,N_1868,N_1996);
or U2134 (N_2134,N_1902,N_1891);
and U2135 (N_2135,N_1935,N_1862);
nor U2136 (N_2136,N_1815,N_1873);
nor U2137 (N_2137,N_1854,N_1889);
nor U2138 (N_2138,N_1981,N_1930);
and U2139 (N_2139,N_1825,N_1975);
and U2140 (N_2140,N_1871,N_1863);
or U2141 (N_2141,N_1970,N_1936);
nand U2142 (N_2142,N_1820,N_1909);
nor U2143 (N_2143,N_1846,N_1863);
and U2144 (N_2144,N_1851,N_1854);
nand U2145 (N_2145,N_1953,N_1979);
xor U2146 (N_2146,N_1965,N_1995);
nand U2147 (N_2147,N_1829,N_1966);
nor U2148 (N_2148,N_1913,N_1962);
nor U2149 (N_2149,N_1952,N_1829);
xnor U2150 (N_2150,N_1800,N_1965);
or U2151 (N_2151,N_1957,N_1851);
xor U2152 (N_2152,N_1999,N_1959);
or U2153 (N_2153,N_1807,N_1803);
and U2154 (N_2154,N_1858,N_1884);
or U2155 (N_2155,N_1935,N_1814);
and U2156 (N_2156,N_1958,N_1809);
nand U2157 (N_2157,N_1939,N_1818);
nand U2158 (N_2158,N_1919,N_1963);
and U2159 (N_2159,N_1823,N_1828);
nor U2160 (N_2160,N_1858,N_1939);
nand U2161 (N_2161,N_1802,N_1900);
and U2162 (N_2162,N_1945,N_1891);
or U2163 (N_2163,N_1961,N_1874);
xnor U2164 (N_2164,N_1966,N_1930);
and U2165 (N_2165,N_1964,N_1984);
xor U2166 (N_2166,N_1967,N_1999);
and U2167 (N_2167,N_1950,N_1986);
or U2168 (N_2168,N_1900,N_1887);
and U2169 (N_2169,N_1814,N_1883);
or U2170 (N_2170,N_1971,N_1872);
xnor U2171 (N_2171,N_1948,N_1928);
or U2172 (N_2172,N_1855,N_1912);
and U2173 (N_2173,N_1881,N_1975);
or U2174 (N_2174,N_1925,N_1851);
and U2175 (N_2175,N_1869,N_1943);
and U2176 (N_2176,N_1933,N_1880);
or U2177 (N_2177,N_1992,N_1965);
nor U2178 (N_2178,N_1840,N_1895);
or U2179 (N_2179,N_1811,N_1897);
or U2180 (N_2180,N_1853,N_1855);
nand U2181 (N_2181,N_1834,N_1963);
or U2182 (N_2182,N_1871,N_1887);
or U2183 (N_2183,N_1901,N_1976);
or U2184 (N_2184,N_1903,N_1968);
xor U2185 (N_2185,N_1968,N_1860);
nand U2186 (N_2186,N_1878,N_1912);
nor U2187 (N_2187,N_1849,N_1966);
and U2188 (N_2188,N_1879,N_1897);
and U2189 (N_2189,N_1811,N_1926);
nor U2190 (N_2190,N_1931,N_1889);
nand U2191 (N_2191,N_1879,N_1903);
nor U2192 (N_2192,N_1948,N_1809);
nor U2193 (N_2193,N_1976,N_1967);
nor U2194 (N_2194,N_1801,N_1921);
and U2195 (N_2195,N_1983,N_1892);
or U2196 (N_2196,N_1918,N_1968);
xor U2197 (N_2197,N_1891,N_1880);
nor U2198 (N_2198,N_1896,N_1867);
nand U2199 (N_2199,N_1805,N_1936);
nand U2200 (N_2200,N_2018,N_2055);
nand U2201 (N_2201,N_2157,N_2088);
and U2202 (N_2202,N_2148,N_2044);
nor U2203 (N_2203,N_2076,N_2134);
nand U2204 (N_2204,N_2027,N_2115);
or U2205 (N_2205,N_2104,N_2140);
or U2206 (N_2206,N_2120,N_2121);
nor U2207 (N_2207,N_2067,N_2078);
xor U2208 (N_2208,N_2166,N_2059);
nand U2209 (N_2209,N_2072,N_2045);
or U2210 (N_2210,N_2191,N_2178);
nor U2211 (N_2211,N_2080,N_2012);
or U2212 (N_2212,N_2083,N_2029);
or U2213 (N_2213,N_2186,N_2193);
nor U2214 (N_2214,N_2093,N_2108);
or U2215 (N_2215,N_2123,N_2173);
nor U2216 (N_2216,N_2165,N_2152);
and U2217 (N_2217,N_2139,N_2103);
nand U2218 (N_2218,N_2130,N_2180);
xnor U2219 (N_2219,N_2006,N_2061);
and U2220 (N_2220,N_2023,N_2026);
nand U2221 (N_2221,N_2011,N_2133);
nor U2222 (N_2222,N_2100,N_2020);
or U2223 (N_2223,N_2184,N_2009);
nand U2224 (N_2224,N_2089,N_2110);
nand U2225 (N_2225,N_2058,N_2098);
and U2226 (N_2226,N_2113,N_2051);
nor U2227 (N_2227,N_2075,N_2032);
nor U2228 (N_2228,N_2106,N_2146);
and U2229 (N_2229,N_2159,N_2174);
or U2230 (N_2230,N_2050,N_2099);
and U2231 (N_2231,N_2064,N_2001);
and U2232 (N_2232,N_2069,N_2153);
or U2233 (N_2233,N_2046,N_2107);
nand U2234 (N_2234,N_2094,N_2131);
or U2235 (N_2235,N_2028,N_2129);
nor U2236 (N_2236,N_2016,N_2062);
or U2237 (N_2237,N_2169,N_2084);
nor U2238 (N_2238,N_2082,N_2022);
or U2239 (N_2239,N_2161,N_2112);
nand U2240 (N_2240,N_2063,N_2198);
and U2241 (N_2241,N_2122,N_2005);
and U2242 (N_2242,N_2014,N_2003);
and U2243 (N_2243,N_2085,N_2071);
nor U2244 (N_2244,N_2164,N_2156);
nand U2245 (N_2245,N_2150,N_2070);
nor U2246 (N_2246,N_2136,N_2041);
nor U2247 (N_2247,N_2127,N_2049);
nor U2248 (N_2248,N_2160,N_2025);
and U2249 (N_2249,N_2034,N_2137);
or U2250 (N_2250,N_2101,N_2079);
nor U2251 (N_2251,N_2176,N_2181);
and U2252 (N_2252,N_2149,N_2043);
or U2253 (N_2253,N_2144,N_2086);
nand U2254 (N_2254,N_2010,N_2054);
or U2255 (N_2255,N_2102,N_2158);
nor U2256 (N_2256,N_2002,N_2039);
or U2257 (N_2257,N_2163,N_2143);
xor U2258 (N_2258,N_2013,N_2081);
nand U2259 (N_2259,N_2036,N_2197);
and U2260 (N_2260,N_2030,N_2188);
and U2261 (N_2261,N_2135,N_2042);
or U2262 (N_2262,N_2092,N_2168);
or U2263 (N_2263,N_2141,N_2096);
nor U2264 (N_2264,N_2024,N_2015);
or U2265 (N_2265,N_2048,N_2128);
nand U2266 (N_2266,N_2124,N_2119);
nand U2267 (N_2267,N_2057,N_2118);
or U2268 (N_2268,N_2179,N_2147);
xnor U2269 (N_2269,N_2170,N_2167);
nand U2270 (N_2270,N_2155,N_2056);
and U2271 (N_2271,N_2047,N_2114);
and U2272 (N_2272,N_2035,N_2019);
nor U2273 (N_2273,N_2073,N_2196);
nor U2274 (N_2274,N_2154,N_2068);
or U2275 (N_2275,N_2008,N_2109);
nand U2276 (N_2276,N_2138,N_2185);
or U2277 (N_2277,N_2172,N_2031);
and U2278 (N_2278,N_2090,N_2195);
nor U2279 (N_2279,N_2132,N_2192);
xnor U2280 (N_2280,N_2066,N_2007);
nand U2281 (N_2281,N_2116,N_2097);
nand U2282 (N_2282,N_2182,N_2171);
or U2283 (N_2283,N_2190,N_2151);
nand U2284 (N_2284,N_2145,N_2033);
xor U2285 (N_2285,N_2199,N_2162);
or U2286 (N_2286,N_2000,N_2194);
or U2287 (N_2287,N_2189,N_2053);
nor U2288 (N_2288,N_2074,N_2105);
and U2289 (N_2289,N_2117,N_2187);
or U2290 (N_2290,N_2175,N_2111);
xor U2291 (N_2291,N_2126,N_2052);
nor U2292 (N_2292,N_2065,N_2183);
nand U2293 (N_2293,N_2060,N_2038);
nor U2294 (N_2294,N_2077,N_2040);
and U2295 (N_2295,N_2021,N_2177);
nand U2296 (N_2296,N_2087,N_2095);
nand U2297 (N_2297,N_2091,N_2004);
and U2298 (N_2298,N_2017,N_2142);
nand U2299 (N_2299,N_2037,N_2125);
and U2300 (N_2300,N_2114,N_2095);
and U2301 (N_2301,N_2188,N_2184);
and U2302 (N_2302,N_2120,N_2041);
xor U2303 (N_2303,N_2007,N_2099);
nor U2304 (N_2304,N_2107,N_2089);
and U2305 (N_2305,N_2106,N_2066);
nand U2306 (N_2306,N_2156,N_2109);
nor U2307 (N_2307,N_2057,N_2139);
and U2308 (N_2308,N_2104,N_2105);
and U2309 (N_2309,N_2156,N_2167);
or U2310 (N_2310,N_2064,N_2075);
nand U2311 (N_2311,N_2152,N_2081);
nand U2312 (N_2312,N_2156,N_2071);
or U2313 (N_2313,N_2132,N_2181);
or U2314 (N_2314,N_2056,N_2077);
and U2315 (N_2315,N_2189,N_2191);
nor U2316 (N_2316,N_2119,N_2078);
and U2317 (N_2317,N_2052,N_2108);
or U2318 (N_2318,N_2110,N_2093);
or U2319 (N_2319,N_2199,N_2133);
nand U2320 (N_2320,N_2139,N_2101);
and U2321 (N_2321,N_2163,N_2115);
nand U2322 (N_2322,N_2105,N_2053);
and U2323 (N_2323,N_2192,N_2188);
and U2324 (N_2324,N_2020,N_2062);
or U2325 (N_2325,N_2057,N_2059);
or U2326 (N_2326,N_2112,N_2190);
or U2327 (N_2327,N_2145,N_2173);
nand U2328 (N_2328,N_2038,N_2056);
nand U2329 (N_2329,N_2135,N_2070);
and U2330 (N_2330,N_2106,N_2168);
nor U2331 (N_2331,N_2061,N_2182);
xnor U2332 (N_2332,N_2014,N_2102);
nor U2333 (N_2333,N_2011,N_2063);
nand U2334 (N_2334,N_2111,N_2040);
or U2335 (N_2335,N_2000,N_2190);
nand U2336 (N_2336,N_2027,N_2169);
or U2337 (N_2337,N_2031,N_2060);
nor U2338 (N_2338,N_2128,N_2174);
and U2339 (N_2339,N_2067,N_2141);
or U2340 (N_2340,N_2152,N_2130);
and U2341 (N_2341,N_2162,N_2049);
nor U2342 (N_2342,N_2103,N_2057);
or U2343 (N_2343,N_2000,N_2157);
or U2344 (N_2344,N_2125,N_2150);
and U2345 (N_2345,N_2157,N_2023);
and U2346 (N_2346,N_2011,N_2161);
nor U2347 (N_2347,N_2013,N_2068);
or U2348 (N_2348,N_2146,N_2199);
and U2349 (N_2349,N_2096,N_2043);
or U2350 (N_2350,N_2085,N_2096);
and U2351 (N_2351,N_2159,N_2018);
nor U2352 (N_2352,N_2094,N_2058);
or U2353 (N_2353,N_2158,N_2000);
nand U2354 (N_2354,N_2037,N_2042);
nor U2355 (N_2355,N_2186,N_2152);
nand U2356 (N_2356,N_2019,N_2015);
or U2357 (N_2357,N_2100,N_2152);
or U2358 (N_2358,N_2036,N_2169);
or U2359 (N_2359,N_2042,N_2046);
nand U2360 (N_2360,N_2077,N_2087);
or U2361 (N_2361,N_2150,N_2087);
nor U2362 (N_2362,N_2191,N_2126);
nand U2363 (N_2363,N_2142,N_2012);
and U2364 (N_2364,N_2086,N_2189);
nand U2365 (N_2365,N_2073,N_2000);
nor U2366 (N_2366,N_2019,N_2111);
xor U2367 (N_2367,N_2143,N_2003);
nand U2368 (N_2368,N_2152,N_2174);
nor U2369 (N_2369,N_2048,N_2077);
or U2370 (N_2370,N_2088,N_2065);
nor U2371 (N_2371,N_2182,N_2107);
or U2372 (N_2372,N_2101,N_2032);
nand U2373 (N_2373,N_2145,N_2175);
nand U2374 (N_2374,N_2091,N_2054);
and U2375 (N_2375,N_2068,N_2155);
or U2376 (N_2376,N_2150,N_2094);
and U2377 (N_2377,N_2062,N_2131);
nand U2378 (N_2378,N_2098,N_2198);
xor U2379 (N_2379,N_2043,N_2101);
or U2380 (N_2380,N_2111,N_2115);
nor U2381 (N_2381,N_2192,N_2134);
nor U2382 (N_2382,N_2141,N_2048);
or U2383 (N_2383,N_2011,N_2023);
nand U2384 (N_2384,N_2028,N_2094);
nor U2385 (N_2385,N_2004,N_2146);
and U2386 (N_2386,N_2050,N_2056);
or U2387 (N_2387,N_2110,N_2039);
xor U2388 (N_2388,N_2138,N_2002);
and U2389 (N_2389,N_2185,N_2021);
or U2390 (N_2390,N_2089,N_2087);
nor U2391 (N_2391,N_2100,N_2033);
xor U2392 (N_2392,N_2087,N_2002);
and U2393 (N_2393,N_2044,N_2115);
xor U2394 (N_2394,N_2166,N_2124);
nand U2395 (N_2395,N_2139,N_2144);
xor U2396 (N_2396,N_2161,N_2141);
or U2397 (N_2397,N_2167,N_2036);
xnor U2398 (N_2398,N_2198,N_2090);
and U2399 (N_2399,N_2088,N_2109);
and U2400 (N_2400,N_2271,N_2300);
or U2401 (N_2401,N_2307,N_2256);
nor U2402 (N_2402,N_2309,N_2247);
xor U2403 (N_2403,N_2306,N_2357);
nor U2404 (N_2404,N_2296,N_2318);
nor U2405 (N_2405,N_2250,N_2333);
and U2406 (N_2406,N_2223,N_2397);
or U2407 (N_2407,N_2208,N_2351);
nor U2408 (N_2408,N_2217,N_2316);
nor U2409 (N_2409,N_2272,N_2252);
xor U2410 (N_2410,N_2265,N_2280);
and U2411 (N_2411,N_2381,N_2387);
or U2412 (N_2412,N_2311,N_2260);
and U2413 (N_2413,N_2382,N_2205);
and U2414 (N_2414,N_2365,N_2320);
and U2415 (N_2415,N_2339,N_2201);
or U2416 (N_2416,N_2375,N_2364);
or U2417 (N_2417,N_2249,N_2344);
and U2418 (N_2418,N_2359,N_2373);
nand U2419 (N_2419,N_2213,N_2353);
nor U2420 (N_2420,N_2334,N_2259);
nor U2421 (N_2421,N_2376,N_2354);
or U2422 (N_2422,N_2386,N_2228);
nor U2423 (N_2423,N_2352,N_2241);
or U2424 (N_2424,N_2370,N_2244);
and U2425 (N_2425,N_2284,N_2206);
nand U2426 (N_2426,N_2248,N_2358);
xor U2427 (N_2427,N_2356,N_2200);
nor U2428 (N_2428,N_2362,N_2343);
and U2429 (N_2429,N_2276,N_2288);
nand U2430 (N_2430,N_2313,N_2299);
nand U2431 (N_2431,N_2328,N_2347);
nand U2432 (N_2432,N_2211,N_2337);
and U2433 (N_2433,N_2292,N_2360);
or U2434 (N_2434,N_2261,N_2240);
or U2435 (N_2435,N_2219,N_2254);
nor U2436 (N_2436,N_2218,N_2236);
nor U2437 (N_2437,N_2349,N_2202);
and U2438 (N_2438,N_2380,N_2281);
nor U2439 (N_2439,N_2212,N_2327);
nor U2440 (N_2440,N_2295,N_2204);
or U2441 (N_2441,N_2310,N_2342);
and U2442 (N_2442,N_2341,N_2222);
xnor U2443 (N_2443,N_2394,N_2203);
or U2444 (N_2444,N_2209,N_2279);
and U2445 (N_2445,N_2245,N_2298);
or U2446 (N_2446,N_2392,N_2361);
and U2447 (N_2447,N_2258,N_2378);
and U2448 (N_2448,N_2274,N_2338);
nor U2449 (N_2449,N_2267,N_2233);
or U2450 (N_2450,N_2291,N_2231);
nor U2451 (N_2451,N_2257,N_2348);
or U2452 (N_2452,N_2326,N_2270);
or U2453 (N_2453,N_2297,N_2224);
nand U2454 (N_2454,N_2329,N_2210);
nand U2455 (N_2455,N_2369,N_2383);
nand U2456 (N_2456,N_2264,N_2301);
and U2457 (N_2457,N_2278,N_2346);
nor U2458 (N_2458,N_2216,N_2230);
and U2459 (N_2459,N_2234,N_2385);
nand U2460 (N_2460,N_2304,N_2302);
or U2461 (N_2461,N_2229,N_2350);
nand U2462 (N_2462,N_2377,N_2289);
and U2463 (N_2463,N_2253,N_2239);
nand U2464 (N_2464,N_2321,N_2235);
nor U2465 (N_2465,N_2323,N_2287);
and U2466 (N_2466,N_2315,N_2393);
or U2467 (N_2467,N_2367,N_2324);
nor U2468 (N_2468,N_2332,N_2322);
and U2469 (N_2469,N_2389,N_2384);
or U2470 (N_2470,N_2374,N_2336);
or U2471 (N_2471,N_2345,N_2319);
and U2472 (N_2472,N_2331,N_2340);
and U2473 (N_2473,N_2221,N_2398);
nand U2474 (N_2474,N_2363,N_2390);
and U2475 (N_2475,N_2325,N_2372);
and U2476 (N_2476,N_2395,N_2399);
nand U2477 (N_2477,N_2282,N_2396);
nand U2478 (N_2478,N_2246,N_2227);
nand U2479 (N_2479,N_2242,N_2285);
nor U2480 (N_2480,N_2290,N_2314);
nand U2481 (N_2481,N_2251,N_2293);
nor U2482 (N_2482,N_2317,N_2286);
xnor U2483 (N_2483,N_2238,N_2215);
nor U2484 (N_2484,N_2273,N_2237);
and U2485 (N_2485,N_2330,N_2391);
xnor U2486 (N_2486,N_2312,N_2232);
or U2487 (N_2487,N_2214,N_2262);
or U2488 (N_2488,N_2207,N_2268);
or U2489 (N_2489,N_2266,N_2355);
or U2490 (N_2490,N_2379,N_2243);
and U2491 (N_2491,N_2368,N_2388);
or U2492 (N_2492,N_2226,N_2275);
nand U2493 (N_2493,N_2283,N_2366);
nand U2494 (N_2494,N_2220,N_2335);
nor U2495 (N_2495,N_2255,N_2294);
or U2496 (N_2496,N_2269,N_2277);
or U2497 (N_2497,N_2303,N_2225);
xnor U2498 (N_2498,N_2308,N_2263);
xnor U2499 (N_2499,N_2305,N_2371);
or U2500 (N_2500,N_2259,N_2294);
or U2501 (N_2501,N_2246,N_2333);
nor U2502 (N_2502,N_2393,N_2334);
and U2503 (N_2503,N_2271,N_2237);
xor U2504 (N_2504,N_2307,N_2388);
xnor U2505 (N_2505,N_2249,N_2241);
or U2506 (N_2506,N_2269,N_2234);
and U2507 (N_2507,N_2284,N_2289);
and U2508 (N_2508,N_2230,N_2247);
and U2509 (N_2509,N_2397,N_2391);
and U2510 (N_2510,N_2302,N_2324);
and U2511 (N_2511,N_2398,N_2342);
and U2512 (N_2512,N_2252,N_2344);
and U2513 (N_2513,N_2276,N_2226);
or U2514 (N_2514,N_2283,N_2270);
or U2515 (N_2515,N_2371,N_2368);
nor U2516 (N_2516,N_2388,N_2347);
and U2517 (N_2517,N_2232,N_2390);
nor U2518 (N_2518,N_2397,N_2232);
or U2519 (N_2519,N_2320,N_2213);
nor U2520 (N_2520,N_2200,N_2207);
nand U2521 (N_2521,N_2317,N_2303);
nor U2522 (N_2522,N_2317,N_2380);
nand U2523 (N_2523,N_2263,N_2335);
nand U2524 (N_2524,N_2315,N_2209);
and U2525 (N_2525,N_2397,N_2372);
and U2526 (N_2526,N_2216,N_2387);
and U2527 (N_2527,N_2329,N_2319);
nand U2528 (N_2528,N_2331,N_2228);
nand U2529 (N_2529,N_2200,N_2309);
nor U2530 (N_2530,N_2216,N_2325);
nand U2531 (N_2531,N_2338,N_2223);
and U2532 (N_2532,N_2353,N_2212);
nand U2533 (N_2533,N_2374,N_2259);
xor U2534 (N_2534,N_2301,N_2298);
nand U2535 (N_2535,N_2382,N_2329);
and U2536 (N_2536,N_2315,N_2261);
nand U2537 (N_2537,N_2223,N_2345);
and U2538 (N_2538,N_2333,N_2311);
and U2539 (N_2539,N_2310,N_2206);
nand U2540 (N_2540,N_2337,N_2236);
and U2541 (N_2541,N_2267,N_2202);
nand U2542 (N_2542,N_2346,N_2356);
nor U2543 (N_2543,N_2205,N_2296);
xnor U2544 (N_2544,N_2292,N_2254);
nand U2545 (N_2545,N_2312,N_2287);
nand U2546 (N_2546,N_2222,N_2330);
nor U2547 (N_2547,N_2361,N_2213);
nor U2548 (N_2548,N_2285,N_2202);
nor U2549 (N_2549,N_2281,N_2302);
or U2550 (N_2550,N_2359,N_2257);
nor U2551 (N_2551,N_2221,N_2350);
xnor U2552 (N_2552,N_2205,N_2311);
or U2553 (N_2553,N_2353,N_2362);
xor U2554 (N_2554,N_2318,N_2268);
nor U2555 (N_2555,N_2298,N_2250);
or U2556 (N_2556,N_2390,N_2366);
or U2557 (N_2557,N_2308,N_2213);
xnor U2558 (N_2558,N_2256,N_2266);
and U2559 (N_2559,N_2276,N_2355);
and U2560 (N_2560,N_2327,N_2241);
nor U2561 (N_2561,N_2327,N_2332);
and U2562 (N_2562,N_2379,N_2254);
or U2563 (N_2563,N_2294,N_2251);
or U2564 (N_2564,N_2365,N_2311);
nand U2565 (N_2565,N_2325,N_2306);
nand U2566 (N_2566,N_2375,N_2288);
or U2567 (N_2567,N_2345,N_2255);
nand U2568 (N_2568,N_2369,N_2262);
nand U2569 (N_2569,N_2239,N_2385);
nor U2570 (N_2570,N_2328,N_2204);
nor U2571 (N_2571,N_2261,N_2212);
nand U2572 (N_2572,N_2338,N_2252);
or U2573 (N_2573,N_2289,N_2212);
nand U2574 (N_2574,N_2288,N_2226);
xnor U2575 (N_2575,N_2266,N_2337);
nor U2576 (N_2576,N_2203,N_2379);
nand U2577 (N_2577,N_2378,N_2278);
or U2578 (N_2578,N_2317,N_2382);
nor U2579 (N_2579,N_2262,N_2201);
or U2580 (N_2580,N_2242,N_2317);
or U2581 (N_2581,N_2250,N_2275);
nor U2582 (N_2582,N_2283,N_2384);
or U2583 (N_2583,N_2272,N_2247);
or U2584 (N_2584,N_2334,N_2251);
nand U2585 (N_2585,N_2250,N_2324);
nor U2586 (N_2586,N_2350,N_2202);
nand U2587 (N_2587,N_2228,N_2205);
xnor U2588 (N_2588,N_2332,N_2339);
and U2589 (N_2589,N_2306,N_2267);
nand U2590 (N_2590,N_2299,N_2306);
nor U2591 (N_2591,N_2322,N_2358);
xnor U2592 (N_2592,N_2306,N_2327);
nor U2593 (N_2593,N_2271,N_2354);
and U2594 (N_2594,N_2276,N_2358);
or U2595 (N_2595,N_2360,N_2254);
nand U2596 (N_2596,N_2340,N_2278);
nand U2597 (N_2597,N_2352,N_2361);
nand U2598 (N_2598,N_2237,N_2391);
and U2599 (N_2599,N_2243,N_2310);
or U2600 (N_2600,N_2537,N_2400);
xnor U2601 (N_2601,N_2436,N_2482);
xnor U2602 (N_2602,N_2512,N_2473);
nor U2603 (N_2603,N_2552,N_2491);
nor U2604 (N_2604,N_2487,N_2430);
and U2605 (N_2605,N_2456,N_2495);
and U2606 (N_2606,N_2501,N_2465);
or U2607 (N_2607,N_2493,N_2422);
or U2608 (N_2608,N_2407,N_2450);
nand U2609 (N_2609,N_2571,N_2448);
or U2610 (N_2610,N_2574,N_2590);
nor U2611 (N_2611,N_2471,N_2500);
xor U2612 (N_2612,N_2541,N_2599);
or U2613 (N_2613,N_2470,N_2401);
or U2614 (N_2614,N_2536,N_2412);
or U2615 (N_2615,N_2404,N_2429);
nor U2616 (N_2616,N_2521,N_2484);
and U2617 (N_2617,N_2560,N_2524);
nand U2618 (N_2618,N_2591,N_2423);
nor U2619 (N_2619,N_2587,N_2554);
and U2620 (N_2620,N_2504,N_2455);
nor U2621 (N_2621,N_2592,N_2567);
nor U2622 (N_2622,N_2489,N_2457);
and U2623 (N_2623,N_2435,N_2546);
xnor U2624 (N_2624,N_2462,N_2507);
nand U2625 (N_2625,N_2481,N_2566);
and U2626 (N_2626,N_2589,N_2438);
nor U2627 (N_2627,N_2562,N_2476);
nor U2628 (N_2628,N_2413,N_2515);
nor U2629 (N_2629,N_2472,N_2461);
or U2630 (N_2630,N_2446,N_2403);
or U2631 (N_2631,N_2505,N_2540);
nand U2632 (N_2632,N_2568,N_2522);
and U2633 (N_2633,N_2518,N_2497);
nand U2634 (N_2634,N_2533,N_2449);
or U2635 (N_2635,N_2596,N_2502);
or U2636 (N_2636,N_2486,N_2576);
or U2637 (N_2637,N_2535,N_2459);
nor U2638 (N_2638,N_2563,N_2514);
nand U2639 (N_2639,N_2556,N_2555);
xnor U2640 (N_2640,N_2437,N_2424);
xnor U2641 (N_2641,N_2573,N_2490);
xnor U2642 (N_2642,N_2539,N_2506);
nor U2643 (N_2643,N_2509,N_2542);
and U2644 (N_2644,N_2468,N_2585);
or U2645 (N_2645,N_2519,N_2498);
and U2646 (N_2646,N_2543,N_2477);
xor U2647 (N_2647,N_2452,N_2494);
nand U2648 (N_2648,N_2416,N_2408);
xor U2649 (N_2649,N_2582,N_2588);
or U2650 (N_2650,N_2525,N_2474);
or U2651 (N_2651,N_2434,N_2410);
and U2652 (N_2652,N_2425,N_2578);
nor U2653 (N_2653,N_2523,N_2460);
nor U2654 (N_2654,N_2564,N_2420);
or U2655 (N_2655,N_2415,N_2508);
and U2656 (N_2656,N_2458,N_2510);
and U2657 (N_2657,N_2469,N_2426);
or U2658 (N_2658,N_2526,N_2547);
and U2659 (N_2659,N_2475,N_2534);
xor U2660 (N_2660,N_2516,N_2527);
nand U2661 (N_2661,N_2451,N_2447);
nor U2662 (N_2662,N_2586,N_2569);
nand U2663 (N_2663,N_2584,N_2443);
or U2664 (N_2664,N_2577,N_2545);
xnor U2665 (N_2665,N_2432,N_2549);
or U2666 (N_2666,N_2419,N_2551);
nand U2667 (N_2667,N_2480,N_2597);
or U2668 (N_2668,N_2439,N_2467);
nor U2669 (N_2669,N_2414,N_2544);
nand U2670 (N_2670,N_2503,N_2579);
or U2671 (N_2671,N_2417,N_2479);
xnor U2672 (N_2672,N_2427,N_2593);
nand U2673 (N_2673,N_2406,N_2421);
nand U2674 (N_2674,N_2442,N_2409);
nor U2675 (N_2675,N_2531,N_2538);
and U2676 (N_2676,N_2492,N_2553);
nor U2677 (N_2677,N_2453,N_2583);
xor U2678 (N_2678,N_2511,N_2598);
or U2679 (N_2679,N_2464,N_2444);
nand U2680 (N_2680,N_2513,N_2463);
nand U2681 (N_2681,N_2496,N_2581);
nor U2682 (N_2682,N_2405,N_2532);
or U2683 (N_2683,N_2485,N_2433);
nand U2684 (N_2684,N_2528,N_2557);
nand U2685 (N_2685,N_2488,N_2411);
nand U2686 (N_2686,N_2428,N_2440);
and U2687 (N_2687,N_2580,N_2454);
nand U2688 (N_2688,N_2565,N_2517);
and U2689 (N_2689,N_2561,N_2402);
nor U2690 (N_2690,N_2595,N_2483);
or U2691 (N_2691,N_2572,N_2530);
nand U2692 (N_2692,N_2441,N_2466);
or U2693 (N_2693,N_2445,N_2529);
nand U2694 (N_2694,N_2548,N_2575);
and U2695 (N_2695,N_2558,N_2418);
or U2696 (N_2696,N_2520,N_2431);
nor U2697 (N_2697,N_2559,N_2550);
and U2698 (N_2698,N_2594,N_2570);
or U2699 (N_2699,N_2499,N_2478);
nand U2700 (N_2700,N_2404,N_2591);
nand U2701 (N_2701,N_2438,N_2516);
or U2702 (N_2702,N_2593,N_2503);
nor U2703 (N_2703,N_2520,N_2435);
nor U2704 (N_2704,N_2461,N_2519);
or U2705 (N_2705,N_2539,N_2528);
or U2706 (N_2706,N_2578,N_2555);
nor U2707 (N_2707,N_2488,N_2583);
nor U2708 (N_2708,N_2451,N_2563);
or U2709 (N_2709,N_2549,N_2455);
and U2710 (N_2710,N_2506,N_2474);
and U2711 (N_2711,N_2585,N_2484);
nor U2712 (N_2712,N_2489,N_2454);
nor U2713 (N_2713,N_2533,N_2535);
and U2714 (N_2714,N_2565,N_2595);
and U2715 (N_2715,N_2537,N_2409);
nor U2716 (N_2716,N_2462,N_2553);
nand U2717 (N_2717,N_2502,N_2594);
and U2718 (N_2718,N_2415,N_2584);
and U2719 (N_2719,N_2567,N_2453);
nor U2720 (N_2720,N_2597,N_2599);
xor U2721 (N_2721,N_2597,N_2524);
or U2722 (N_2722,N_2466,N_2436);
and U2723 (N_2723,N_2456,N_2501);
or U2724 (N_2724,N_2474,N_2554);
and U2725 (N_2725,N_2528,N_2495);
nand U2726 (N_2726,N_2519,N_2471);
nor U2727 (N_2727,N_2482,N_2419);
nand U2728 (N_2728,N_2470,N_2516);
nand U2729 (N_2729,N_2573,N_2407);
or U2730 (N_2730,N_2534,N_2448);
and U2731 (N_2731,N_2468,N_2523);
and U2732 (N_2732,N_2407,N_2535);
nand U2733 (N_2733,N_2551,N_2517);
nor U2734 (N_2734,N_2422,N_2561);
or U2735 (N_2735,N_2510,N_2592);
nand U2736 (N_2736,N_2491,N_2591);
nor U2737 (N_2737,N_2406,N_2558);
or U2738 (N_2738,N_2460,N_2579);
xnor U2739 (N_2739,N_2459,N_2581);
xnor U2740 (N_2740,N_2468,N_2474);
nor U2741 (N_2741,N_2555,N_2481);
xnor U2742 (N_2742,N_2462,N_2481);
nor U2743 (N_2743,N_2523,N_2581);
or U2744 (N_2744,N_2428,N_2483);
nand U2745 (N_2745,N_2545,N_2497);
nand U2746 (N_2746,N_2518,N_2567);
nand U2747 (N_2747,N_2572,N_2500);
nand U2748 (N_2748,N_2599,N_2402);
nand U2749 (N_2749,N_2574,N_2522);
or U2750 (N_2750,N_2475,N_2419);
and U2751 (N_2751,N_2400,N_2515);
nor U2752 (N_2752,N_2591,N_2579);
and U2753 (N_2753,N_2465,N_2547);
nand U2754 (N_2754,N_2530,N_2558);
nand U2755 (N_2755,N_2557,N_2545);
nand U2756 (N_2756,N_2509,N_2425);
or U2757 (N_2757,N_2411,N_2438);
and U2758 (N_2758,N_2506,N_2599);
nor U2759 (N_2759,N_2545,N_2408);
or U2760 (N_2760,N_2409,N_2592);
xor U2761 (N_2761,N_2571,N_2457);
nor U2762 (N_2762,N_2597,N_2572);
and U2763 (N_2763,N_2593,N_2414);
nand U2764 (N_2764,N_2528,N_2526);
nand U2765 (N_2765,N_2522,N_2525);
and U2766 (N_2766,N_2541,N_2597);
nand U2767 (N_2767,N_2456,N_2428);
or U2768 (N_2768,N_2590,N_2533);
nand U2769 (N_2769,N_2459,N_2482);
or U2770 (N_2770,N_2567,N_2487);
nor U2771 (N_2771,N_2437,N_2412);
or U2772 (N_2772,N_2555,N_2434);
nor U2773 (N_2773,N_2487,N_2598);
or U2774 (N_2774,N_2511,N_2591);
or U2775 (N_2775,N_2423,N_2532);
xnor U2776 (N_2776,N_2507,N_2426);
xnor U2777 (N_2777,N_2448,N_2539);
xnor U2778 (N_2778,N_2557,N_2457);
nand U2779 (N_2779,N_2575,N_2437);
nand U2780 (N_2780,N_2524,N_2526);
nand U2781 (N_2781,N_2546,N_2538);
or U2782 (N_2782,N_2558,N_2515);
and U2783 (N_2783,N_2451,N_2406);
or U2784 (N_2784,N_2582,N_2494);
nor U2785 (N_2785,N_2495,N_2443);
nor U2786 (N_2786,N_2518,N_2542);
or U2787 (N_2787,N_2513,N_2444);
nand U2788 (N_2788,N_2595,N_2504);
or U2789 (N_2789,N_2528,N_2472);
xor U2790 (N_2790,N_2492,N_2574);
and U2791 (N_2791,N_2417,N_2598);
or U2792 (N_2792,N_2580,N_2543);
or U2793 (N_2793,N_2527,N_2486);
nor U2794 (N_2794,N_2460,N_2592);
or U2795 (N_2795,N_2587,N_2515);
nor U2796 (N_2796,N_2563,N_2518);
or U2797 (N_2797,N_2474,N_2589);
xnor U2798 (N_2798,N_2467,N_2562);
nor U2799 (N_2799,N_2533,N_2526);
nor U2800 (N_2800,N_2784,N_2600);
and U2801 (N_2801,N_2733,N_2788);
nand U2802 (N_2802,N_2698,N_2686);
xor U2803 (N_2803,N_2735,N_2718);
or U2804 (N_2804,N_2662,N_2756);
xnor U2805 (N_2805,N_2769,N_2675);
nand U2806 (N_2806,N_2665,N_2615);
nor U2807 (N_2807,N_2731,N_2645);
nor U2808 (N_2808,N_2751,N_2630);
or U2809 (N_2809,N_2725,N_2714);
nor U2810 (N_2810,N_2746,N_2642);
nand U2811 (N_2811,N_2652,N_2684);
and U2812 (N_2812,N_2604,N_2711);
nand U2813 (N_2813,N_2708,N_2669);
or U2814 (N_2814,N_2749,N_2750);
xnor U2815 (N_2815,N_2752,N_2779);
and U2816 (N_2816,N_2639,N_2795);
nor U2817 (N_2817,N_2623,N_2780);
and U2818 (N_2818,N_2719,N_2762);
and U2819 (N_2819,N_2608,N_2712);
or U2820 (N_2820,N_2744,N_2758);
nor U2821 (N_2821,N_2619,N_2793);
xor U2822 (N_2822,N_2760,N_2678);
nand U2823 (N_2823,N_2730,N_2786);
or U2824 (N_2824,N_2606,N_2612);
or U2825 (N_2825,N_2660,N_2628);
nand U2826 (N_2826,N_2626,N_2768);
and U2827 (N_2827,N_2705,N_2759);
nand U2828 (N_2828,N_2763,N_2697);
or U2829 (N_2829,N_2681,N_2723);
xnor U2830 (N_2830,N_2778,N_2636);
and U2831 (N_2831,N_2741,N_2605);
or U2832 (N_2832,N_2611,N_2656);
and U2833 (N_2833,N_2745,N_2776);
and U2834 (N_2834,N_2674,N_2740);
or U2835 (N_2835,N_2620,N_2783);
nor U2836 (N_2836,N_2610,N_2794);
nand U2837 (N_2837,N_2755,N_2624);
xnor U2838 (N_2838,N_2707,N_2618);
nor U2839 (N_2839,N_2693,N_2706);
nand U2840 (N_2840,N_2797,N_2632);
nand U2841 (N_2841,N_2650,N_2704);
nor U2842 (N_2842,N_2754,N_2690);
xor U2843 (N_2843,N_2774,N_2689);
nand U2844 (N_2844,N_2777,N_2692);
nor U2845 (N_2845,N_2677,N_2709);
or U2846 (N_2846,N_2748,N_2694);
and U2847 (N_2847,N_2631,N_2622);
and U2848 (N_2848,N_2721,N_2775);
and U2849 (N_2849,N_2664,N_2696);
nand U2850 (N_2850,N_2781,N_2753);
nor U2851 (N_2851,N_2661,N_2720);
and U2852 (N_2852,N_2603,N_2643);
xor U2853 (N_2853,N_2787,N_2700);
nand U2854 (N_2854,N_2770,N_2742);
nand U2855 (N_2855,N_2743,N_2773);
nand U2856 (N_2856,N_2683,N_2771);
and U2857 (N_2857,N_2738,N_2616);
nand U2858 (N_2858,N_2695,N_2621);
nand U2859 (N_2859,N_2799,N_2614);
or U2860 (N_2860,N_2676,N_2727);
nor U2861 (N_2861,N_2654,N_2666);
and U2862 (N_2862,N_2757,N_2798);
nand U2863 (N_2863,N_2617,N_2633);
nor U2864 (N_2864,N_2792,N_2634);
or U2865 (N_2865,N_2637,N_2737);
or U2866 (N_2866,N_2739,N_2641);
and U2867 (N_2867,N_2644,N_2673);
nor U2868 (N_2868,N_2668,N_2717);
or U2869 (N_2869,N_2657,N_2638);
and U2870 (N_2870,N_2682,N_2734);
nor U2871 (N_2871,N_2635,N_2796);
nor U2872 (N_2872,N_2767,N_2648);
xor U2873 (N_2873,N_2715,N_2761);
nor U2874 (N_2874,N_2728,N_2703);
and U2875 (N_2875,N_2640,N_2766);
nor U2876 (N_2876,N_2724,N_2627);
or U2877 (N_2877,N_2670,N_2649);
nor U2878 (N_2878,N_2672,N_2671);
nor U2879 (N_2879,N_2651,N_2782);
and U2880 (N_2880,N_2685,N_2765);
nand U2881 (N_2881,N_2732,N_2691);
or U2882 (N_2882,N_2716,N_2790);
and U2883 (N_2883,N_2713,N_2601);
nand U2884 (N_2884,N_2679,N_2785);
or U2885 (N_2885,N_2722,N_2613);
or U2886 (N_2886,N_2747,N_2602);
and U2887 (N_2887,N_2791,N_2653);
xnor U2888 (N_2888,N_2607,N_2646);
or U2889 (N_2889,N_2687,N_2729);
or U2890 (N_2890,N_2629,N_2764);
and U2891 (N_2891,N_2688,N_2647);
nor U2892 (N_2892,N_2655,N_2667);
xnor U2893 (N_2893,N_2789,N_2658);
nand U2894 (N_2894,N_2609,N_2710);
nor U2895 (N_2895,N_2680,N_2772);
nor U2896 (N_2896,N_2625,N_2726);
xor U2897 (N_2897,N_2699,N_2663);
nor U2898 (N_2898,N_2736,N_2659);
nand U2899 (N_2899,N_2702,N_2701);
and U2900 (N_2900,N_2734,N_2732);
nand U2901 (N_2901,N_2748,N_2640);
or U2902 (N_2902,N_2789,N_2631);
and U2903 (N_2903,N_2786,N_2610);
nand U2904 (N_2904,N_2701,N_2663);
xnor U2905 (N_2905,N_2674,N_2647);
or U2906 (N_2906,N_2631,N_2777);
or U2907 (N_2907,N_2794,N_2682);
nor U2908 (N_2908,N_2659,N_2781);
nor U2909 (N_2909,N_2745,N_2699);
or U2910 (N_2910,N_2680,N_2701);
or U2911 (N_2911,N_2613,N_2687);
or U2912 (N_2912,N_2772,N_2694);
nand U2913 (N_2913,N_2740,N_2605);
and U2914 (N_2914,N_2689,N_2766);
and U2915 (N_2915,N_2602,N_2615);
or U2916 (N_2916,N_2767,N_2666);
xnor U2917 (N_2917,N_2780,N_2714);
nand U2918 (N_2918,N_2614,N_2717);
or U2919 (N_2919,N_2714,N_2641);
or U2920 (N_2920,N_2617,N_2606);
xor U2921 (N_2921,N_2767,N_2743);
and U2922 (N_2922,N_2604,N_2799);
nor U2923 (N_2923,N_2609,N_2681);
and U2924 (N_2924,N_2678,N_2623);
nor U2925 (N_2925,N_2612,N_2763);
nor U2926 (N_2926,N_2741,N_2737);
nand U2927 (N_2927,N_2657,N_2645);
nor U2928 (N_2928,N_2643,N_2701);
and U2929 (N_2929,N_2716,N_2616);
nor U2930 (N_2930,N_2677,N_2650);
and U2931 (N_2931,N_2797,N_2688);
nand U2932 (N_2932,N_2744,N_2780);
and U2933 (N_2933,N_2676,N_2755);
nand U2934 (N_2934,N_2646,N_2709);
or U2935 (N_2935,N_2784,N_2643);
or U2936 (N_2936,N_2731,N_2732);
nand U2937 (N_2937,N_2729,N_2761);
nand U2938 (N_2938,N_2762,N_2738);
nor U2939 (N_2939,N_2703,N_2777);
and U2940 (N_2940,N_2763,N_2667);
or U2941 (N_2941,N_2663,N_2698);
nor U2942 (N_2942,N_2730,N_2635);
nand U2943 (N_2943,N_2772,N_2692);
or U2944 (N_2944,N_2668,N_2769);
and U2945 (N_2945,N_2615,N_2649);
or U2946 (N_2946,N_2740,N_2691);
or U2947 (N_2947,N_2664,N_2628);
and U2948 (N_2948,N_2620,N_2662);
and U2949 (N_2949,N_2668,N_2734);
nand U2950 (N_2950,N_2613,N_2661);
xnor U2951 (N_2951,N_2764,N_2761);
nor U2952 (N_2952,N_2777,N_2743);
and U2953 (N_2953,N_2722,N_2690);
or U2954 (N_2954,N_2741,N_2683);
and U2955 (N_2955,N_2648,N_2674);
nand U2956 (N_2956,N_2688,N_2705);
and U2957 (N_2957,N_2687,N_2611);
nand U2958 (N_2958,N_2790,N_2683);
nor U2959 (N_2959,N_2688,N_2640);
xor U2960 (N_2960,N_2600,N_2663);
nand U2961 (N_2961,N_2743,N_2703);
or U2962 (N_2962,N_2753,N_2752);
or U2963 (N_2963,N_2752,N_2654);
or U2964 (N_2964,N_2774,N_2688);
and U2965 (N_2965,N_2726,N_2715);
and U2966 (N_2966,N_2701,N_2705);
nand U2967 (N_2967,N_2744,N_2656);
nor U2968 (N_2968,N_2633,N_2665);
and U2969 (N_2969,N_2693,N_2697);
nand U2970 (N_2970,N_2626,N_2764);
or U2971 (N_2971,N_2667,N_2639);
and U2972 (N_2972,N_2667,N_2735);
or U2973 (N_2973,N_2628,N_2686);
nor U2974 (N_2974,N_2771,N_2741);
nor U2975 (N_2975,N_2731,N_2693);
or U2976 (N_2976,N_2660,N_2732);
nor U2977 (N_2977,N_2602,N_2666);
and U2978 (N_2978,N_2756,N_2795);
nand U2979 (N_2979,N_2641,N_2614);
nand U2980 (N_2980,N_2603,N_2661);
nand U2981 (N_2981,N_2663,N_2743);
nor U2982 (N_2982,N_2749,N_2658);
nor U2983 (N_2983,N_2746,N_2787);
nand U2984 (N_2984,N_2666,N_2638);
or U2985 (N_2985,N_2663,N_2707);
and U2986 (N_2986,N_2623,N_2744);
or U2987 (N_2987,N_2617,N_2719);
and U2988 (N_2988,N_2627,N_2709);
or U2989 (N_2989,N_2722,N_2673);
nand U2990 (N_2990,N_2766,N_2792);
nand U2991 (N_2991,N_2769,N_2756);
nand U2992 (N_2992,N_2757,N_2659);
nor U2993 (N_2993,N_2624,N_2685);
nand U2994 (N_2994,N_2763,N_2620);
nand U2995 (N_2995,N_2689,N_2718);
xnor U2996 (N_2996,N_2688,N_2719);
nor U2997 (N_2997,N_2674,N_2750);
xor U2998 (N_2998,N_2734,N_2669);
or U2999 (N_2999,N_2669,N_2664);
and U3000 (N_3000,N_2816,N_2886);
or U3001 (N_3001,N_2853,N_2960);
or U3002 (N_3002,N_2876,N_2963);
nor U3003 (N_3003,N_2897,N_2926);
xnor U3004 (N_3004,N_2843,N_2943);
or U3005 (N_3005,N_2978,N_2942);
nor U3006 (N_3006,N_2845,N_2988);
nor U3007 (N_3007,N_2894,N_2927);
nor U3008 (N_3008,N_2891,N_2850);
and U3009 (N_3009,N_2923,N_2907);
or U3010 (N_3010,N_2858,N_2861);
nand U3011 (N_3011,N_2870,N_2854);
nand U3012 (N_3012,N_2893,N_2903);
nor U3013 (N_3013,N_2892,N_2972);
nor U3014 (N_3014,N_2838,N_2970);
or U3015 (N_3015,N_2940,N_2920);
nor U3016 (N_3016,N_2958,N_2971);
or U3017 (N_3017,N_2931,N_2924);
xor U3018 (N_3018,N_2864,N_2915);
and U3019 (N_3019,N_2840,N_2828);
nand U3020 (N_3020,N_2977,N_2994);
nand U3021 (N_3021,N_2914,N_2967);
nand U3022 (N_3022,N_2944,N_2883);
nand U3023 (N_3023,N_2992,N_2947);
or U3024 (N_3024,N_2936,N_2820);
and U3025 (N_3025,N_2811,N_2812);
and U3026 (N_3026,N_2884,N_2996);
or U3027 (N_3027,N_2941,N_2909);
or U3028 (N_3028,N_2986,N_2800);
and U3029 (N_3029,N_2991,N_2844);
nor U3030 (N_3030,N_2881,N_2921);
nand U3031 (N_3031,N_2846,N_2832);
nand U3032 (N_3032,N_2849,N_2929);
or U3033 (N_3033,N_2852,N_2842);
nand U3034 (N_3034,N_2899,N_2887);
and U3035 (N_3035,N_2813,N_2865);
nand U3036 (N_3036,N_2801,N_2857);
and U3037 (N_3037,N_2949,N_2868);
nor U3038 (N_3038,N_2895,N_2910);
nor U3039 (N_3039,N_2980,N_2961);
or U3040 (N_3040,N_2912,N_2911);
nor U3041 (N_3041,N_2898,N_2888);
xor U3042 (N_3042,N_2872,N_2904);
nor U3043 (N_3043,N_2965,N_2847);
and U3044 (N_3044,N_2950,N_2873);
and U3045 (N_3045,N_2976,N_2815);
nor U3046 (N_3046,N_2835,N_2954);
nand U3047 (N_3047,N_2998,N_2863);
nor U3048 (N_3048,N_2932,N_2827);
nor U3049 (N_3049,N_2959,N_2885);
nand U3050 (N_3050,N_2928,N_2839);
or U3051 (N_3051,N_2948,N_2836);
and U3052 (N_3052,N_2818,N_2829);
nor U3053 (N_3053,N_2803,N_2952);
xor U3054 (N_3054,N_2995,N_2878);
and U3055 (N_3055,N_2862,N_2964);
and U3056 (N_3056,N_2946,N_2937);
and U3057 (N_3057,N_2997,N_2826);
xnor U3058 (N_3058,N_2807,N_2804);
nor U3059 (N_3059,N_2908,N_2848);
nand U3060 (N_3060,N_2825,N_2900);
and U3061 (N_3061,N_2830,N_2981);
nand U3062 (N_3062,N_2985,N_2817);
nand U3063 (N_3063,N_2860,N_2837);
nand U3064 (N_3064,N_2880,N_2957);
and U3065 (N_3065,N_2906,N_2821);
or U3066 (N_3066,N_2993,N_2953);
nor U3067 (N_3067,N_2859,N_2851);
or U3068 (N_3068,N_2919,N_2866);
nand U3069 (N_3069,N_2938,N_2999);
or U3070 (N_3070,N_2984,N_2974);
nor U3071 (N_3071,N_2975,N_2833);
and U3072 (N_3072,N_2905,N_2918);
nor U3073 (N_3073,N_2982,N_2831);
nor U3074 (N_3074,N_2869,N_2916);
or U3075 (N_3075,N_2955,N_2902);
or U3076 (N_3076,N_2896,N_2979);
and U3077 (N_3077,N_2934,N_2969);
nand U3078 (N_3078,N_2856,N_2824);
or U3079 (N_3079,N_2871,N_2874);
and U3080 (N_3080,N_2990,N_2930);
xnor U3081 (N_3081,N_2823,N_2841);
and U3082 (N_3082,N_2962,N_2933);
nand U3083 (N_3083,N_2935,N_2882);
nor U3084 (N_3084,N_2890,N_2819);
or U3085 (N_3085,N_2917,N_2968);
nor U3086 (N_3086,N_2901,N_2939);
nor U3087 (N_3087,N_2855,N_2802);
nand U3088 (N_3088,N_2951,N_2913);
and U3089 (N_3089,N_2925,N_2814);
and U3090 (N_3090,N_2922,N_2809);
and U3091 (N_3091,N_2966,N_2945);
nand U3092 (N_3092,N_2875,N_2805);
or U3093 (N_3093,N_2983,N_2956);
nor U3094 (N_3094,N_2889,N_2806);
nand U3095 (N_3095,N_2973,N_2822);
xor U3096 (N_3096,N_2987,N_2989);
and U3097 (N_3097,N_2808,N_2810);
and U3098 (N_3098,N_2879,N_2877);
nand U3099 (N_3099,N_2834,N_2867);
and U3100 (N_3100,N_2967,N_2827);
and U3101 (N_3101,N_2899,N_2894);
or U3102 (N_3102,N_2976,N_2907);
or U3103 (N_3103,N_2821,N_2940);
xor U3104 (N_3104,N_2893,N_2829);
or U3105 (N_3105,N_2803,N_2960);
or U3106 (N_3106,N_2822,N_2843);
nand U3107 (N_3107,N_2896,N_2906);
and U3108 (N_3108,N_2990,N_2964);
nor U3109 (N_3109,N_2985,N_2875);
or U3110 (N_3110,N_2908,N_2931);
and U3111 (N_3111,N_2809,N_2972);
nor U3112 (N_3112,N_2847,N_2925);
nand U3113 (N_3113,N_2911,N_2922);
or U3114 (N_3114,N_2908,N_2899);
nor U3115 (N_3115,N_2877,N_2801);
or U3116 (N_3116,N_2994,N_2874);
or U3117 (N_3117,N_2836,N_2870);
and U3118 (N_3118,N_2936,N_2843);
and U3119 (N_3119,N_2993,N_2982);
nand U3120 (N_3120,N_2845,N_2946);
xnor U3121 (N_3121,N_2913,N_2991);
or U3122 (N_3122,N_2815,N_2986);
nor U3123 (N_3123,N_2949,N_2935);
or U3124 (N_3124,N_2873,N_2803);
nand U3125 (N_3125,N_2891,N_2852);
or U3126 (N_3126,N_2897,N_2915);
or U3127 (N_3127,N_2874,N_2899);
xnor U3128 (N_3128,N_2988,N_2867);
nand U3129 (N_3129,N_2956,N_2965);
nand U3130 (N_3130,N_2932,N_2891);
and U3131 (N_3131,N_2999,N_2836);
or U3132 (N_3132,N_2850,N_2948);
and U3133 (N_3133,N_2861,N_2852);
nand U3134 (N_3134,N_2892,N_2911);
or U3135 (N_3135,N_2859,N_2967);
and U3136 (N_3136,N_2989,N_2801);
nor U3137 (N_3137,N_2955,N_2834);
nor U3138 (N_3138,N_2871,N_2860);
or U3139 (N_3139,N_2988,N_2837);
or U3140 (N_3140,N_2830,N_2839);
or U3141 (N_3141,N_2937,N_2811);
xnor U3142 (N_3142,N_2851,N_2852);
nand U3143 (N_3143,N_2936,N_2892);
or U3144 (N_3144,N_2867,N_2920);
nand U3145 (N_3145,N_2864,N_2859);
and U3146 (N_3146,N_2908,N_2865);
or U3147 (N_3147,N_2825,N_2820);
xor U3148 (N_3148,N_2911,N_2935);
or U3149 (N_3149,N_2976,N_2861);
and U3150 (N_3150,N_2860,N_2864);
nor U3151 (N_3151,N_2916,N_2952);
nor U3152 (N_3152,N_2866,N_2841);
xnor U3153 (N_3153,N_2846,N_2923);
nor U3154 (N_3154,N_2811,N_2983);
or U3155 (N_3155,N_2852,N_2967);
nor U3156 (N_3156,N_2981,N_2955);
or U3157 (N_3157,N_2830,N_2904);
or U3158 (N_3158,N_2845,N_2902);
nand U3159 (N_3159,N_2880,N_2833);
xor U3160 (N_3160,N_2864,N_2900);
nor U3161 (N_3161,N_2827,N_2961);
nor U3162 (N_3162,N_2894,N_2829);
xnor U3163 (N_3163,N_2827,N_2940);
xor U3164 (N_3164,N_2835,N_2813);
nor U3165 (N_3165,N_2871,N_2961);
nand U3166 (N_3166,N_2882,N_2970);
nand U3167 (N_3167,N_2804,N_2924);
or U3168 (N_3168,N_2888,N_2865);
or U3169 (N_3169,N_2898,N_2939);
and U3170 (N_3170,N_2903,N_2917);
nor U3171 (N_3171,N_2849,N_2867);
nor U3172 (N_3172,N_2888,N_2928);
and U3173 (N_3173,N_2870,N_2861);
or U3174 (N_3174,N_2815,N_2861);
and U3175 (N_3175,N_2933,N_2826);
nor U3176 (N_3176,N_2966,N_2866);
xor U3177 (N_3177,N_2999,N_2820);
nand U3178 (N_3178,N_2975,N_2874);
or U3179 (N_3179,N_2877,N_2826);
xnor U3180 (N_3180,N_2825,N_2933);
and U3181 (N_3181,N_2835,N_2960);
and U3182 (N_3182,N_2875,N_2871);
nand U3183 (N_3183,N_2898,N_2822);
nand U3184 (N_3184,N_2878,N_2829);
nand U3185 (N_3185,N_2985,N_2863);
and U3186 (N_3186,N_2831,N_2947);
nor U3187 (N_3187,N_2924,N_2906);
or U3188 (N_3188,N_2869,N_2910);
or U3189 (N_3189,N_2987,N_2948);
nor U3190 (N_3190,N_2917,N_2858);
xor U3191 (N_3191,N_2888,N_2877);
xor U3192 (N_3192,N_2806,N_2973);
or U3193 (N_3193,N_2849,N_2831);
and U3194 (N_3194,N_2802,N_2828);
nand U3195 (N_3195,N_2804,N_2900);
nand U3196 (N_3196,N_2818,N_2915);
or U3197 (N_3197,N_2863,N_2834);
and U3198 (N_3198,N_2864,N_2985);
nor U3199 (N_3199,N_2983,N_2972);
and U3200 (N_3200,N_3023,N_3126);
or U3201 (N_3201,N_3027,N_3085);
or U3202 (N_3202,N_3135,N_3131);
nor U3203 (N_3203,N_3180,N_3002);
nor U3204 (N_3204,N_3094,N_3179);
or U3205 (N_3205,N_3021,N_3127);
and U3206 (N_3206,N_3093,N_3003);
and U3207 (N_3207,N_3182,N_3087);
nand U3208 (N_3208,N_3080,N_3071);
nand U3209 (N_3209,N_3194,N_3000);
nand U3210 (N_3210,N_3175,N_3177);
xnor U3211 (N_3211,N_3061,N_3103);
xor U3212 (N_3212,N_3189,N_3178);
nor U3213 (N_3213,N_3114,N_3163);
nand U3214 (N_3214,N_3084,N_3174);
or U3215 (N_3215,N_3157,N_3143);
or U3216 (N_3216,N_3048,N_3079);
nand U3217 (N_3217,N_3173,N_3113);
nor U3218 (N_3218,N_3054,N_3035);
nand U3219 (N_3219,N_3133,N_3187);
and U3220 (N_3220,N_3044,N_3160);
and U3221 (N_3221,N_3089,N_3146);
xnor U3222 (N_3222,N_3176,N_3001);
and U3223 (N_3223,N_3156,N_3168);
xor U3224 (N_3224,N_3170,N_3104);
nor U3225 (N_3225,N_3040,N_3106);
nand U3226 (N_3226,N_3012,N_3062);
nand U3227 (N_3227,N_3077,N_3092);
or U3228 (N_3228,N_3016,N_3041);
or U3229 (N_3229,N_3145,N_3043);
and U3230 (N_3230,N_3196,N_3121);
nor U3231 (N_3231,N_3192,N_3183);
or U3232 (N_3232,N_3117,N_3090);
nor U3233 (N_3233,N_3075,N_3019);
nand U3234 (N_3234,N_3086,N_3051);
or U3235 (N_3235,N_3172,N_3128);
nand U3236 (N_3236,N_3130,N_3036);
and U3237 (N_3237,N_3142,N_3099);
nand U3238 (N_3238,N_3153,N_3185);
and U3239 (N_3239,N_3070,N_3052);
or U3240 (N_3240,N_3129,N_3055);
nor U3241 (N_3241,N_3109,N_3042);
or U3242 (N_3242,N_3038,N_3060);
and U3243 (N_3243,N_3100,N_3101);
xnor U3244 (N_3244,N_3063,N_3088);
or U3245 (N_3245,N_3065,N_3020);
nor U3246 (N_3246,N_3032,N_3154);
and U3247 (N_3247,N_3081,N_3110);
xor U3248 (N_3248,N_3164,N_3056);
or U3249 (N_3249,N_3057,N_3144);
xor U3250 (N_3250,N_3150,N_3125);
or U3251 (N_3251,N_3190,N_3017);
and U3252 (N_3252,N_3188,N_3031);
or U3253 (N_3253,N_3096,N_3013);
or U3254 (N_3254,N_3167,N_3181);
nand U3255 (N_3255,N_3053,N_3024);
nor U3256 (N_3256,N_3004,N_3137);
and U3257 (N_3257,N_3158,N_3030);
nand U3258 (N_3258,N_3059,N_3049);
nor U3259 (N_3259,N_3132,N_3037);
nand U3260 (N_3260,N_3166,N_3171);
nor U3261 (N_3261,N_3026,N_3006);
nor U3262 (N_3262,N_3091,N_3107);
or U3263 (N_3263,N_3082,N_3047);
nand U3264 (N_3264,N_3139,N_3152);
or U3265 (N_3265,N_3014,N_3193);
nand U3266 (N_3266,N_3076,N_3169);
and U3267 (N_3267,N_3074,N_3010);
and U3268 (N_3268,N_3149,N_3159);
nand U3269 (N_3269,N_3115,N_3095);
or U3270 (N_3270,N_3008,N_3102);
or U3271 (N_3271,N_3067,N_3033);
nand U3272 (N_3272,N_3184,N_3072);
nand U3273 (N_3273,N_3025,N_3122);
nor U3274 (N_3274,N_3140,N_3165);
or U3275 (N_3275,N_3138,N_3098);
nand U3276 (N_3276,N_3136,N_3045);
nand U3277 (N_3277,N_3083,N_3015);
xnor U3278 (N_3278,N_3018,N_3034);
nand U3279 (N_3279,N_3148,N_3123);
nor U3280 (N_3280,N_3011,N_3124);
nand U3281 (N_3281,N_3151,N_3078);
nor U3282 (N_3282,N_3108,N_3112);
nor U3283 (N_3283,N_3147,N_3111);
nand U3284 (N_3284,N_3066,N_3073);
nand U3285 (N_3285,N_3191,N_3161);
nor U3286 (N_3286,N_3186,N_3022);
nor U3287 (N_3287,N_3097,N_3039);
nor U3288 (N_3288,N_3162,N_3118);
or U3289 (N_3289,N_3050,N_3119);
and U3290 (N_3290,N_3199,N_3198);
or U3291 (N_3291,N_3134,N_3068);
and U3292 (N_3292,N_3195,N_3007);
nand U3293 (N_3293,N_3028,N_3155);
nor U3294 (N_3294,N_3009,N_3046);
nor U3295 (N_3295,N_3105,N_3120);
nor U3296 (N_3296,N_3058,N_3064);
or U3297 (N_3297,N_3069,N_3116);
or U3298 (N_3298,N_3005,N_3197);
and U3299 (N_3299,N_3141,N_3029);
nand U3300 (N_3300,N_3078,N_3005);
and U3301 (N_3301,N_3162,N_3144);
and U3302 (N_3302,N_3013,N_3146);
nand U3303 (N_3303,N_3129,N_3127);
nand U3304 (N_3304,N_3191,N_3157);
nand U3305 (N_3305,N_3132,N_3026);
nor U3306 (N_3306,N_3171,N_3057);
nor U3307 (N_3307,N_3056,N_3001);
and U3308 (N_3308,N_3193,N_3131);
nand U3309 (N_3309,N_3028,N_3052);
nand U3310 (N_3310,N_3166,N_3027);
nor U3311 (N_3311,N_3129,N_3143);
nand U3312 (N_3312,N_3026,N_3095);
nor U3313 (N_3313,N_3007,N_3059);
xnor U3314 (N_3314,N_3081,N_3171);
or U3315 (N_3315,N_3116,N_3035);
and U3316 (N_3316,N_3180,N_3014);
nor U3317 (N_3317,N_3118,N_3012);
or U3318 (N_3318,N_3116,N_3174);
xor U3319 (N_3319,N_3156,N_3050);
or U3320 (N_3320,N_3172,N_3050);
xnor U3321 (N_3321,N_3046,N_3135);
or U3322 (N_3322,N_3009,N_3193);
or U3323 (N_3323,N_3022,N_3119);
and U3324 (N_3324,N_3029,N_3018);
or U3325 (N_3325,N_3057,N_3111);
or U3326 (N_3326,N_3007,N_3091);
nor U3327 (N_3327,N_3155,N_3066);
nor U3328 (N_3328,N_3174,N_3183);
nand U3329 (N_3329,N_3094,N_3140);
nand U3330 (N_3330,N_3021,N_3164);
nor U3331 (N_3331,N_3065,N_3148);
and U3332 (N_3332,N_3187,N_3045);
nand U3333 (N_3333,N_3143,N_3172);
and U3334 (N_3334,N_3143,N_3164);
and U3335 (N_3335,N_3123,N_3049);
and U3336 (N_3336,N_3084,N_3089);
nor U3337 (N_3337,N_3161,N_3013);
or U3338 (N_3338,N_3090,N_3146);
and U3339 (N_3339,N_3082,N_3195);
xnor U3340 (N_3340,N_3000,N_3102);
nor U3341 (N_3341,N_3021,N_3097);
and U3342 (N_3342,N_3114,N_3164);
and U3343 (N_3343,N_3123,N_3166);
and U3344 (N_3344,N_3088,N_3097);
nand U3345 (N_3345,N_3006,N_3113);
or U3346 (N_3346,N_3039,N_3171);
nor U3347 (N_3347,N_3120,N_3013);
or U3348 (N_3348,N_3122,N_3138);
or U3349 (N_3349,N_3022,N_3089);
nand U3350 (N_3350,N_3000,N_3114);
nand U3351 (N_3351,N_3028,N_3013);
or U3352 (N_3352,N_3121,N_3056);
nor U3353 (N_3353,N_3051,N_3024);
or U3354 (N_3354,N_3072,N_3155);
and U3355 (N_3355,N_3027,N_3078);
and U3356 (N_3356,N_3124,N_3140);
nand U3357 (N_3357,N_3141,N_3169);
xor U3358 (N_3358,N_3017,N_3013);
xor U3359 (N_3359,N_3000,N_3116);
nand U3360 (N_3360,N_3156,N_3007);
or U3361 (N_3361,N_3120,N_3017);
xnor U3362 (N_3362,N_3160,N_3108);
nand U3363 (N_3363,N_3029,N_3102);
xnor U3364 (N_3364,N_3053,N_3163);
nor U3365 (N_3365,N_3150,N_3035);
or U3366 (N_3366,N_3065,N_3030);
nor U3367 (N_3367,N_3053,N_3196);
nand U3368 (N_3368,N_3166,N_3174);
and U3369 (N_3369,N_3196,N_3009);
nand U3370 (N_3370,N_3072,N_3104);
nor U3371 (N_3371,N_3166,N_3137);
nor U3372 (N_3372,N_3158,N_3067);
or U3373 (N_3373,N_3136,N_3146);
and U3374 (N_3374,N_3195,N_3164);
and U3375 (N_3375,N_3149,N_3050);
nand U3376 (N_3376,N_3005,N_3109);
or U3377 (N_3377,N_3139,N_3146);
nand U3378 (N_3378,N_3034,N_3121);
nand U3379 (N_3379,N_3149,N_3085);
nand U3380 (N_3380,N_3175,N_3031);
and U3381 (N_3381,N_3182,N_3074);
nand U3382 (N_3382,N_3191,N_3125);
nor U3383 (N_3383,N_3019,N_3178);
nand U3384 (N_3384,N_3189,N_3165);
nand U3385 (N_3385,N_3074,N_3174);
xnor U3386 (N_3386,N_3047,N_3006);
or U3387 (N_3387,N_3034,N_3178);
xnor U3388 (N_3388,N_3140,N_3126);
nor U3389 (N_3389,N_3181,N_3063);
nand U3390 (N_3390,N_3171,N_3122);
nor U3391 (N_3391,N_3026,N_3044);
nand U3392 (N_3392,N_3116,N_3196);
and U3393 (N_3393,N_3155,N_3091);
nand U3394 (N_3394,N_3156,N_3140);
or U3395 (N_3395,N_3190,N_3113);
nand U3396 (N_3396,N_3001,N_3142);
and U3397 (N_3397,N_3055,N_3062);
xor U3398 (N_3398,N_3007,N_3121);
or U3399 (N_3399,N_3135,N_3198);
nor U3400 (N_3400,N_3330,N_3322);
xor U3401 (N_3401,N_3256,N_3271);
nor U3402 (N_3402,N_3277,N_3320);
or U3403 (N_3403,N_3270,N_3205);
nand U3404 (N_3404,N_3201,N_3382);
nand U3405 (N_3405,N_3223,N_3312);
xnor U3406 (N_3406,N_3289,N_3244);
nand U3407 (N_3407,N_3286,N_3341);
or U3408 (N_3408,N_3337,N_3309);
nand U3409 (N_3409,N_3370,N_3297);
nor U3410 (N_3410,N_3266,N_3376);
xnor U3411 (N_3411,N_3378,N_3300);
or U3412 (N_3412,N_3272,N_3317);
nand U3413 (N_3413,N_3319,N_3398);
nand U3414 (N_3414,N_3357,N_3298);
or U3415 (N_3415,N_3374,N_3233);
and U3416 (N_3416,N_3208,N_3220);
or U3417 (N_3417,N_3218,N_3287);
nor U3418 (N_3418,N_3221,N_3384);
xor U3419 (N_3419,N_3396,N_3225);
and U3420 (N_3420,N_3213,N_3294);
or U3421 (N_3421,N_3202,N_3227);
and U3422 (N_3422,N_3333,N_3359);
or U3423 (N_3423,N_3386,N_3217);
nor U3424 (N_3424,N_3399,N_3389);
nand U3425 (N_3425,N_3234,N_3347);
nor U3426 (N_3426,N_3246,N_3274);
nor U3427 (N_3427,N_3315,N_3257);
or U3428 (N_3428,N_3303,N_3241);
or U3429 (N_3429,N_3200,N_3393);
and U3430 (N_3430,N_3348,N_3212);
and U3431 (N_3431,N_3306,N_3259);
nand U3432 (N_3432,N_3362,N_3388);
nand U3433 (N_3433,N_3314,N_3344);
nor U3434 (N_3434,N_3283,N_3245);
or U3435 (N_3435,N_3260,N_3381);
nor U3436 (N_3436,N_3302,N_3224);
and U3437 (N_3437,N_3351,N_3358);
and U3438 (N_3438,N_3332,N_3237);
nand U3439 (N_3439,N_3325,N_3295);
nor U3440 (N_3440,N_3232,N_3216);
nor U3441 (N_3441,N_3292,N_3343);
nand U3442 (N_3442,N_3250,N_3375);
nor U3443 (N_3443,N_3211,N_3385);
or U3444 (N_3444,N_3355,N_3236);
nor U3445 (N_3445,N_3318,N_3268);
nor U3446 (N_3446,N_3361,N_3339);
xor U3447 (N_3447,N_3251,N_3331);
and U3448 (N_3448,N_3327,N_3258);
and U3449 (N_3449,N_3369,N_3379);
and U3450 (N_3450,N_3282,N_3383);
xor U3451 (N_3451,N_3360,N_3279);
xor U3452 (N_3452,N_3335,N_3254);
nor U3453 (N_3453,N_3299,N_3372);
and U3454 (N_3454,N_3278,N_3334);
nor U3455 (N_3455,N_3313,N_3323);
or U3456 (N_3456,N_3242,N_3356);
or U3457 (N_3457,N_3229,N_3366);
and U3458 (N_3458,N_3349,N_3345);
or U3459 (N_3459,N_3252,N_3228);
and U3460 (N_3460,N_3392,N_3316);
and U3461 (N_3461,N_3394,N_3276);
and U3462 (N_3462,N_3215,N_3263);
or U3463 (N_3463,N_3203,N_3353);
or U3464 (N_3464,N_3346,N_3284);
nor U3465 (N_3465,N_3321,N_3243);
xor U3466 (N_3466,N_3281,N_3340);
or U3467 (N_3467,N_3364,N_3373);
nor U3468 (N_3468,N_3280,N_3238);
nor U3469 (N_3469,N_3328,N_3267);
or U3470 (N_3470,N_3307,N_3288);
nand U3471 (N_3471,N_3336,N_3311);
nand U3472 (N_3472,N_3249,N_3371);
or U3473 (N_3473,N_3308,N_3255);
nand U3474 (N_3474,N_3273,N_3324);
nor U3475 (N_3475,N_3247,N_3350);
nand U3476 (N_3476,N_3235,N_3231);
nand U3477 (N_3477,N_3264,N_3352);
xor U3478 (N_3478,N_3326,N_3261);
nand U3479 (N_3479,N_3305,N_3391);
nor U3480 (N_3480,N_3304,N_3275);
nor U3481 (N_3481,N_3397,N_3363);
nand U3482 (N_3482,N_3206,N_3338);
and U3483 (N_3483,N_3354,N_3207);
nand U3484 (N_3484,N_3291,N_3293);
nor U3485 (N_3485,N_3285,N_3380);
and U3486 (N_3486,N_3395,N_3262);
nor U3487 (N_3487,N_3222,N_3230);
nor U3488 (N_3488,N_3290,N_3387);
nor U3489 (N_3489,N_3210,N_3253);
nand U3490 (N_3490,N_3240,N_3265);
xor U3491 (N_3491,N_3296,N_3204);
nand U3492 (N_3492,N_3239,N_3368);
nor U3493 (N_3493,N_3329,N_3214);
and U3494 (N_3494,N_3367,N_3390);
and U3495 (N_3495,N_3209,N_3310);
and U3496 (N_3496,N_3226,N_3342);
nor U3497 (N_3497,N_3301,N_3365);
and U3498 (N_3498,N_3377,N_3248);
and U3499 (N_3499,N_3269,N_3219);
nor U3500 (N_3500,N_3309,N_3389);
and U3501 (N_3501,N_3216,N_3335);
and U3502 (N_3502,N_3347,N_3267);
nand U3503 (N_3503,N_3225,N_3214);
and U3504 (N_3504,N_3370,N_3306);
nor U3505 (N_3505,N_3257,N_3360);
nand U3506 (N_3506,N_3399,N_3318);
or U3507 (N_3507,N_3306,N_3326);
or U3508 (N_3508,N_3361,N_3358);
xor U3509 (N_3509,N_3343,N_3380);
nor U3510 (N_3510,N_3333,N_3240);
nand U3511 (N_3511,N_3357,N_3211);
nand U3512 (N_3512,N_3321,N_3239);
or U3513 (N_3513,N_3250,N_3228);
or U3514 (N_3514,N_3311,N_3233);
or U3515 (N_3515,N_3324,N_3346);
nand U3516 (N_3516,N_3280,N_3240);
nor U3517 (N_3517,N_3346,N_3358);
and U3518 (N_3518,N_3201,N_3333);
or U3519 (N_3519,N_3377,N_3235);
nor U3520 (N_3520,N_3292,N_3315);
nand U3521 (N_3521,N_3248,N_3249);
xnor U3522 (N_3522,N_3368,N_3302);
or U3523 (N_3523,N_3367,N_3292);
and U3524 (N_3524,N_3254,N_3287);
nor U3525 (N_3525,N_3290,N_3306);
and U3526 (N_3526,N_3224,N_3246);
nor U3527 (N_3527,N_3264,N_3391);
and U3528 (N_3528,N_3319,N_3276);
or U3529 (N_3529,N_3356,N_3206);
or U3530 (N_3530,N_3244,N_3274);
or U3531 (N_3531,N_3291,N_3366);
xor U3532 (N_3532,N_3352,N_3224);
nor U3533 (N_3533,N_3238,N_3233);
and U3534 (N_3534,N_3231,N_3302);
nand U3535 (N_3535,N_3240,N_3259);
nand U3536 (N_3536,N_3295,N_3303);
nand U3537 (N_3537,N_3390,N_3253);
nand U3538 (N_3538,N_3300,N_3276);
nand U3539 (N_3539,N_3312,N_3307);
nand U3540 (N_3540,N_3293,N_3236);
nand U3541 (N_3541,N_3309,N_3326);
or U3542 (N_3542,N_3326,N_3292);
and U3543 (N_3543,N_3357,N_3387);
nand U3544 (N_3544,N_3384,N_3291);
nand U3545 (N_3545,N_3230,N_3291);
and U3546 (N_3546,N_3200,N_3211);
xor U3547 (N_3547,N_3296,N_3388);
nand U3548 (N_3548,N_3371,N_3350);
and U3549 (N_3549,N_3330,N_3209);
nor U3550 (N_3550,N_3301,N_3351);
or U3551 (N_3551,N_3216,N_3321);
nand U3552 (N_3552,N_3202,N_3259);
and U3553 (N_3553,N_3306,N_3334);
and U3554 (N_3554,N_3367,N_3351);
nand U3555 (N_3555,N_3282,N_3201);
nor U3556 (N_3556,N_3212,N_3241);
nand U3557 (N_3557,N_3399,N_3237);
and U3558 (N_3558,N_3260,N_3294);
nor U3559 (N_3559,N_3380,N_3395);
nor U3560 (N_3560,N_3399,N_3255);
nor U3561 (N_3561,N_3249,N_3261);
or U3562 (N_3562,N_3317,N_3201);
nor U3563 (N_3563,N_3290,N_3225);
nor U3564 (N_3564,N_3295,N_3221);
or U3565 (N_3565,N_3349,N_3222);
or U3566 (N_3566,N_3388,N_3232);
nand U3567 (N_3567,N_3269,N_3221);
nor U3568 (N_3568,N_3287,N_3238);
xor U3569 (N_3569,N_3235,N_3283);
or U3570 (N_3570,N_3303,N_3378);
or U3571 (N_3571,N_3305,N_3228);
xnor U3572 (N_3572,N_3375,N_3223);
and U3573 (N_3573,N_3274,N_3222);
nor U3574 (N_3574,N_3342,N_3293);
and U3575 (N_3575,N_3273,N_3384);
and U3576 (N_3576,N_3367,N_3383);
nor U3577 (N_3577,N_3296,N_3277);
nand U3578 (N_3578,N_3380,N_3206);
nor U3579 (N_3579,N_3308,N_3296);
or U3580 (N_3580,N_3268,N_3276);
and U3581 (N_3581,N_3375,N_3297);
or U3582 (N_3582,N_3328,N_3258);
and U3583 (N_3583,N_3361,N_3321);
or U3584 (N_3584,N_3279,N_3374);
and U3585 (N_3585,N_3361,N_3382);
and U3586 (N_3586,N_3370,N_3330);
and U3587 (N_3587,N_3279,N_3397);
nand U3588 (N_3588,N_3201,N_3352);
nor U3589 (N_3589,N_3276,N_3233);
nand U3590 (N_3590,N_3288,N_3217);
nand U3591 (N_3591,N_3266,N_3381);
or U3592 (N_3592,N_3339,N_3366);
nand U3593 (N_3593,N_3380,N_3398);
nor U3594 (N_3594,N_3262,N_3232);
nor U3595 (N_3595,N_3260,N_3210);
nand U3596 (N_3596,N_3371,N_3320);
or U3597 (N_3597,N_3368,N_3261);
or U3598 (N_3598,N_3222,N_3373);
nand U3599 (N_3599,N_3398,N_3251);
nor U3600 (N_3600,N_3452,N_3510);
and U3601 (N_3601,N_3523,N_3552);
or U3602 (N_3602,N_3546,N_3592);
or U3603 (N_3603,N_3488,N_3457);
xnor U3604 (N_3604,N_3545,N_3470);
or U3605 (N_3605,N_3521,N_3493);
or U3606 (N_3606,N_3496,N_3487);
and U3607 (N_3607,N_3400,N_3535);
nand U3608 (N_3608,N_3514,N_3464);
nor U3609 (N_3609,N_3438,N_3558);
nor U3610 (N_3610,N_3499,N_3486);
and U3611 (N_3611,N_3557,N_3524);
nor U3612 (N_3612,N_3477,N_3412);
xnor U3613 (N_3613,N_3599,N_3575);
and U3614 (N_3614,N_3563,N_3576);
nor U3615 (N_3615,N_3583,N_3430);
nand U3616 (N_3616,N_3489,N_3436);
nand U3617 (N_3617,N_3474,N_3542);
and U3618 (N_3618,N_3589,N_3429);
xnor U3619 (N_3619,N_3459,N_3569);
or U3620 (N_3620,N_3403,N_3409);
and U3621 (N_3621,N_3570,N_3568);
nand U3622 (N_3622,N_3500,N_3597);
nor U3623 (N_3623,N_3567,N_3402);
nor U3624 (N_3624,N_3505,N_3519);
or U3625 (N_3625,N_3468,N_3465);
and U3626 (N_3626,N_3455,N_3553);
nand U3627 (N_3627,N_3417,N_3461);
nor U3628 (N_3628,N_3561,N_3579);
xnor U3629 (N_3629,N_3444,N_3442);
nand U3630 (N_3630,N_3588,N_3462);
or U3631 (N_3631,N_3598,N_3541);
nand U3632 (N_3632,N_3432,N_3591);
nor U3633 (N_3633,N_3481,N_3504);
and U3634 (N_3634,N_3536,N_3596);
and U3635 (N_3635,N_3437,N_3447);
nand U3636 (N_3636,N_3419,N_3483);
xnor U3637 (N_3637,N_3418,N_3564);
nand U3638 (N_3638,N_3456,N_3485);
nor U3639 (N_3639,N_3414,N_3428);
nand U3640 (N_3640,N_3533,N_3406);
and U3641 (N_3641,N_3478,N_3475);
xnor U3642 (N_3642,N_3467,N_3508);
or U3643 (N_3643,N_3476,N_3503);
and U3644 (N_3644,N_3404,N_3450);
nor U3645 (N_3645,N_3534,N_3540);
nand U3646 (N_3646,N_3526,N_3482);
and U3647 (N_3647,N_3416,N_3415);
nand U3648 (N_3648,N_3427,N_3492);
nor U3649 (N_3649,N_3449,N_3543);
xor U3650 (N_3650,N_3559,N_3562);
or U3651 (N_3651,N_3539,N_3527);
or U3652 (N_3652,N_3547,N_3466);
nand U3653 (N_3653,N_3423,N_3420);
xnor U3654 (N_3654,N_3440,N_3448);
nor U3655 (N_3655,N_3435,N_3560);
and U3656 (N_3656,N_3401,N_3425);
xnor U3657 (N_3657,N_3408,N_3593);
or U3658 (N_3658,N_3550,N_3515);
or U3659 (N_3659,N_3507,N_3445);
or U3660 (N_3660,N_3439,N_3453);
nand U3661 (N_3661,N_3573,N_3517);
and U3662 (N_3662,N_3580,N_3458);
and U3663 (N_3663,N_3511,N_3585);
or U3664 (N_3664,N_3512,N_3454);
nand U3665 (N_3665,N_3538,N_3469);
nand U3666 (N_3666,N_3446,N_3497);
or U3667 (N_3667,N_3594,N_3590);
and U3668 (N_3668,N_3525,N_3581);
nor U3669 (N_3669,N_3577,N_3460);
xor U3670 (N_3670,N_3407,N_3516);
nand U3671 (N_3671,N_3551,N_3413);
or U3672 (N_3672,N_3480,N_3502);
or U3673 (N_3673,N_3441,N_3528);
and U3674 (N_3674,N_3565,N_3513);
or U3675 (N_3675,N_3491,N_3431);
and U3676 (N_3676,N_3548,N_3582);
or U3677 (N_3677,N_3584,N_3451);
or U3678 (N_3678,N_3555,N_3586);
or U3679 (N_3679,N_3537,N_3556);
or U3680 (N_3680,N_3422,N_3554);
nand U3681 (N_3681,N_3424,N_3495);
nand U3682 (N_3682,N_3484,N_3421);
or U3683 (N_3683,N_3411,N_3574);
nand U3684 (N_3684,N_3518,N_3494);
nor U3685 (N_3685,N_3571,N_3509);
or U3686 (N_3686,N_3498,N_3544);
and U3687 (N_3687,N_3471,N_3433);
xnor U3688 (N_3688,N_3473,N_3532);
nor U3689 (N_3689,N_3463,N_3530);
nor U3690 (N_3690,N_3479,N_3472);
or U3691 (N_3691,N_3566,N_3587);
or U3692 (N_3692,N_3529,N_3410);
or U3693 (N_3693,N_3426,N_3531);
nor U3694 (N_3694,N_3572,N_3549);
and U3695 (N_3695,N_3443,N_3522);
and U3696 (N_3696,N_3501,N_3405);
xor U3697 (N_3697,N_3506,N_3434);
nand U3698 (N_3698,N_3578,N_3595);
and U3699 (N_3699,N_3520,N_3490);
and U3700 (N_3700,N_3403,N_3416);
or U3701 (N_3701,N_3594,N_3542);
nand U3702 (N_3702,N_3518,N_3467);
or U3703 (N_3703,N_3425,N_3518);
nand U3704 (N_3704,N_3416,N_3559);
nand U3705 (N_3705,N_3522,N_3492);
nor U3706 (N_3706,N_3566,N_3441);
and U3707 (N_3707,N_3532,N_3475);
or U3708 (N_3708,N_3411,N_3526);
or U3709 (N_3709,N_3413,N_3425);
nand U3710 (N_3710,N_3548,N_3546);
or U3711 (N_3711,N_3586,N_3515);
and U3712 (N_3712,N_3503,N_3441);
nor U3713 (N_3713,N_3576,N_3401);
and U3714 (N_3714,N_3587,N_3568);
nor U3715 (N_3715,N_3477,N_3423);
xnor U3716 (N_3716,N_3459,N_3556);
nand U3717 (N_3717,N_3476,N_3558);
nor U3718 (N_3718,N_3441,N_3469);
nor U3719 (N_3719,N_3430,N_3593);
or U3720 (N_3720,N_3513,N_3537);
and U3721 (N_3721,N_3476,N_3516);
nor U3722 (N_3722,N_3436,N_3503);
and U3723 (N_3723,N_3438,N_3567);
xor U3724 (N_3724,N_3533,N_3577);
and U3725 (N_3725,N_3547,N_3462);
nor U3726 (N_3726,N_3540,N_3459);
nor U3727 (N_3727,N_3406,N_3425);
nand U3728 (N_3728,N_3509,N_3406);
nand U3729 (N_3729,N_3534,N_3576);
nor U3730 (N_3730,N_3452,N_3415);
nor U3731 (N_3731,N_3496,N_3539);
xor U3732 (N_3732,N_3514,N_3433);
nand U3733 (N_3733,N_3546,N_3532);
nor U3734 (N_3734,N_3447,N_3582);
and U3735 (N_3735,N_3556,N_3573);
nand U3736 (N_3736,N_3403,N_3475);
xor U3737 (N_3737,N_3564,N_3429);
or U3738 (N_3738,N_3508,N_3439);
nand U3739 (N_3739,N_3566,N_3438);
and U3740 (N_3740,N_3455,N_3469);
nor U3741 (N_3741,N_3475,N_3446);
or U3742 (N_3742,N_3448,N_3513);
and U3743 (N_3743,N_3423,N_3455);
nand U3744 (N_3744,N_3419,N_3586);
and U3745 (N_3745,N_3430,N_3463);
xnor U3746 (N_3746,N_3476,N_3575);
nand U3747 (N_3747,N_3494,N_3567);
or U3748 (N_3748,N_3415,N_3519);
or U3749 (N_3749,N_3539,N_3584);
nand U3750 (N_3750,N_3501,N_3442);
nor U3751 (N_3751,N_3410,N_3516);
and U3752 (N_3752,N_3544,N_3458);
nor U3753 (N_3753,N_3566,N_3468);
and U3754 (N_3754,N_3559,N_3557);
and U3755 (N_3755,N_3419,N_3472);
and U3756 (N_3756,N_3486,N_3458);
or U3757 (N_3757,N_3431,N_3573);
and U3758 (N_3758,N_3438,N_3445);
nand U3759 (N_3759,N_3561,N_3530);
or U3760 (N_3760,N_3487,N_3497);
xor U3761 (N_3761,N_3446,N_3541);
and U3762 (N_3762,N_3418,N_3501);
or U3763 (N_3763,N_3562,N_3451);
and U3764 (N_3764,N_3482,N_3581);
nor U3765 (N_3765,N_3420,N_3502);
xor U3766 (N_3766,N_3440,N_3438);
or U3767 (N_3767,N_3411,N_3463);
nor U3768 (N_3768,N_3576,N_3554);
nor U3769 (N_3769,N_3506,N_3500);
and U3770 (N_3770,N_3495,N_3510);
nand U3771 (N_3771,N_3449,N_3558);
xor U3772 (N_3772,N_3493,N_3467);
xor U3773 (N_3773,N_3595,N_3553);
nor U3774 (N_3774,N_3436,N_3523);
xor U3775 (N_3775,N_3470,N_3414);
nor U3776 (N_3776,N_3419,N_3522);
nor U3777 (N_3777,N_3496,N_3413);
or U3778 (N_3778,N_3501,N_3519);
or U3779 (N_3779,N_3592,N_3468);
nand U3780 (N_3780,N_3429,N_3483);
nand U3781 (N_3781,N_3552,N_3509);
nor U3782 (N_3782,N_3410,N_3460);
nor U3783 (N_3783,N_3485,N_3597);
nor U3784 (N_3784,N_3564,N_3595);
or U3785 (N_3785,N_3478,N_3531);
nand U3786 (N_3786,N_3478,N_3462);
and U3787 (N_3787,N_3404,N_3534);
and U3788 (N_3788,N_3507,N_3451);
xor U3789 (N_3789,N_3586,N_3594);
nor U3790 (N_3790,N_3536,N_3418);
and U3791 (N_3791,N_3467,N_3403);
and U3792 (N_3792,N_3552,N_3412);
and U3793 (N_3793,N_3518,N_3424);
nor U3794 (N_3794,N_3435,N_3581);
nor U3795 (N_3795,N_3403,N_3491);
xnor U3796 (N_3796,N_3509,N_3597);
or U3797 (N_3797,N_3402,N_3505);
nor U3798 (N_3798,N_3532,N_3504);
and U3799 (N_3799,N_3511,N_3458);
nor U3800 (N_3800,N_3679,N_3707);
nor U3801 (N_3801,N_3641,N_3669);
nand U3802 (N_3802,N_3628,N_3785);
nand U3803 (N_3803,N_3681,N_3631);
xor U3804 (N_3804,N_3731,N_3717);
nor U3805 (N_3805,N_3721,N_3757);
nor U3806 (N_3806,N_3771,N_3786);
nor U3807 (N_3807,N_3759,N_3646);
nand U3808 (N_3808,N_3649,N_3633);
nand U3809 (N_3809,N_3670,N_3756);
nor U3810 (N_3810,N_3782,N_3763);
nand U3811 (N_3811,N_3619,N_3788);
nand U3812 (N_3812,N_3699,N_3792);
nand U3813 (N_3813,N_3607,N_3748);
xor U3814 (N_3814,N_3660,N_3709);
nor U3815 (N_3815,N_3621,N_3667);
nand U3816 (N_3816,N_3609,N_3722);
nand U3817 (N_3817,N_3711,N_3603);
nor U3818 (N_3818,N_3701,N_3634);
or U3819 (N_3819,N_3650,N_3752);
nor U3820 (N_3820,N_3687,N_3776);
and U3821 (N_3821,N_3613,N_3662);
nor U3822 (N_3822,N_3637,N_3651);
xnor U3823 (N_3823,N_3738,N_3610);
and U3824 (N_3824,N_3682,N_3769);
or U3825 (N_3825,N_3636,N_3724);
or U3826 (N_3826,N_3758,N_3790);
nand U3827 (N_3827,N_3606,N_3766);
nand U3828 (N_3828,N_3787,N_3652);
nor U3829 (N_3829,N_3668,N_3625);
and U3830 (N_3830,N_3653,N_3632);
and U3831 (N_3831,N_3629,N_3744);
or U3832 (N_3832,N_3730,N_3614);
or U3833 (N_3833,N_3640,N_3616);
and U3834 (N_3834,N_3658,N_3762);
nand U3835 (N_3835,N_3693,N_3765);
nand U3836 (N_3836,N_3689,N_3737);
or U3837 (N_3837,N_3797,N_3725);
nor U3838 (N_3838,N_3615,N_3674);
and U3839 (N_3839,N_3655,N_3661);
or U3840 (N_3840,N_3691,N_3645);
and U3841 (N_3841,N_3751,N_3611);
or U3842 (N_3842,N_3779,N_3695);
xor U3843 (N_3843,N_3755,N_3665);
nand U3844 (N_3844,N_3784,N_3686);
or U3845 (N_3845,N_3704,N_3753);
nor U3846 (N_3846,N_3747,N_3783);
and U3847 (N_3847,N_3671,N_3600);
nand U3848 (N_3848,N_3732,N_3749);
xor U3849 (N_3849,N_3768,N_3643);
and U3850 (N_3850,N_3639,N_3627);
or U3851 (N_3851,N_3690,N_3648);
and U3852 (N_3852,N_3781,N_3718);
xnor U3853 (N_3853,N_3723,N_3720);
or U3854 (N_3854,N_3692,N_3688);
nand U3855 (N_3855,N_3663,N_3623);
nand U3856 (N_3856,N_3703,N_3608);
and U3857 (N_3857,N_3789,N_3685);
nand U3858 (N_3858,N_3713,N_3777);
or U3859 (N_3859,N_3684,N_3742);
nand U3860 (N_3860,N_3739,N_3715);
and U3861 (N_3861,N_3624,N_3657);
or U3862 (N_3862,N_3735,N_3673);
nand U3863 (N_3863,N_3694,N_3745);
xor U3864 (N_3864,N_3635,N_3672);
nand U3865 (N_3865,N_3605,N_3676);
or U3866 (N_3866,N_3677,N_3678);
xor U3867 (N_3867,N_3659,N_3794);
and U3868 (N_3868,N_3602,N_3799);
nor U3869 (N_3869,N_3760,N_3626);
nor U3870 (N_3870,N_3736,N_3706);
nor U3871 (N_3871,N_3716,N_3683);
and U3872 (N_3872,N_3750,N_3618);
nor U3873 (N_3873,N_3710,N_3740);
xor U3874 (N_3874,N_3795,N_3743);
or U3875 (N_3875,N_3767,N_3729);
nor U3876 (N_3876,N_3680,N_3727);
nand U3877 (N_3877,N_3664,N_3714);
nand U3878 (N_3878,N_3746,N_3697);
nand U3879 (N_3879,N_3772,N_3741);
or U3880 (N_3880,N_3675,N_3764);
or U3881 (N_3881,N_3601,N_3644);
xor U3882 (N_3882,N_3793,N_3761);
xnor U3883 (N_3883,N_3617,N_3698);
xnor U3884 (N_3884,N_3630,N_3798);
or U3885 (N_3885,N_3791,N_3734);
nor U3886 (N_3886,N_3780,N_3770);
or U3887 (N_3887,N_3622,N_3696);
nor U3888 (N_3888,N_3604,N_3700);
nand U3889 (N_3889,N_3666,N_3647);
xor U3890 (N_3890,N_3796,N_3612);
and U3891 (N_3891,N_3773,N_3620);
nor U3892 (N_3892,N_3728,N_3638);
and U3893 (N_3893,N_3775,N_3654);
nor U3894 (N_3894,N_3702,N_3754);
xnor U3895 (N_3895,N_3778,N_3719);
nand U3896 (N_3896,N_3708,N_3774);
nand U3897 (N_3897,N_3712,N_3642);
xor U3898 (N_3898,N_3726,N_3656);
and U3899 (N_3899,N_3733,N_3705);
nor U3900 (N_3900,N_3722,N_3765);
xor U3901 (N_3901,N_3768,N_3616);
and U3902 (N_3902,N_3764,N_3758);
nand U3903 (N_3903,N_3776,N_3723);
nand U3904 (N_3904,N_3792,N_3673);
nand U3905 (N_3905,N_3764,N_3629);
xnor U3906 (N_3906,N_3731,N_3653);
and U3907 (N_3907,N_3775,N_3736);
and U3908 (N_3908,N_3656,N_3635);
and U3909 (N_3909,N_3654,N_3721);
and U3910 (N_3910,N_3610,N_3707);
nor U3911 (N_3911,N_3790,N_3739);
xnor U3912 (N_3912,N_3751,N_3738);
xor U3913 (N_3913,N_3656,N_3649);
nand U3914 (N_3914,N_3689,N_3797);
nand U3915 (N_3915,N_3665,N_3718);
xor U3916 (N_3916,N_3790,N_3763);
or U3917 (N_3917,N_3743,N_3780);
xor U3918 (N_3918,N_3688,N_3637);
and U3919 (N_3919,N_3738,N_3620);
nand U3920 (N_3920,N_3656,N_3798);
or U3921 (N_3921,N_3748,N_3758);
xnor U3922 (N_3922,N_3778,N_3782);
nor U3923 (N_3923,N_3710,N_3607);
and U3924 (N_3924,N_3665,N_3679);
nand U3925 (N_3925,N_3665,N_3744);
or U3926 (N_3926,N_3640,N_3766);
and U3927 (N_3927,N_3792,N_3723);
and U3928 (N_3928,N_3636,N_3628);
and U3929 (N_3929,N_3605,N_3769);
nand U3930 (N_3930,N_3731,N_3655);
xnor U3931 (N_3931,N_3788,N_3779);
nand U3932 (N_3932,N_3780,N_3726);
or U3933 (N_3933,N_3710,N_3606);
nor U3934 (N_3934,N_3709,N_3615);
nor U3935 (N_3935,N_3778,N_3752);
and U3936 (N_3936,N_3666,N_3613);
and U3937 (N_3937,N_3673,N_3632);
and U3938 (N_3938,N_3654,N_3703);
xor U3939 (N_3939,N_3775,N_3708);
nor U3940 (N_3940,N_3652,N_3691);
and U3941 (N_3941,N_3633,N_3750);
nand U3942 (N_3942,N_3658,N_3783);
xor U3943 (N_3943,N_3745,N_3645);
or U3944 (N_3944,N_3782,N_3642);
xnor U3945 (N_3945,N_3752,N_3708);
or U3946 (N_3946,N_3722,N_3710);
or U3947 (N_3947,N_3746,N_3786);
xnor U3948 (N_3948,N_3770,N_3617);
or U3949 (N_3949,N_3696,N_3636);
or U3950 (N_3950,N_3719,N_3625);
nor U3951 (N_3951,N_3609,N_3780);
nor U3952 (N_3952,N_3699,N_3798);
and U3953 (N_3953,N_3680,N_3670);
and U3954 (N_3954,N_3737,N_3736);
nor U3955 (N_3955,N_3712,N_3766);
and U3956 (N_3956,N_3786,N_3662);
or U3957 (N_3957,N_3600,N_3721);
nor U3958 (N_3958,N_3640,N_3799);
nand U3959 (N_3959,N_3635,N_3667);
nand U3960 (N_3960,N_3686,N_3775);
and U3961 (N_3961,N_3774,N_3796);
or U3962 (N_3962,N_3784,N_3714);
nand U3963 (N_3963,N_3694,N_3602);
or U3964 (N_3964,N_3714,N_3647);
or U3965 (N_3965,N_3730,N_3788);
nand U3966 (N_3966,N_3786,N_3680);
xor U3967 (N_3967,N_3645,N_3629);
or U3968 (N_3968,N_3798,N_3682);
nor U3969 (N_3969,N_3725,N_3747);
and U3970 (N_3970,N_3729,N_3618);
nand U3971 (N_3971,N_3686,N_3672);
or U3972 (N_3972,N_3734,N_3659);
nor U3973 (N_3973,N_3708,N_3639);
xnor U3974 (N_3974,N_3774,N_3637);
nor U3975 (N_3975,N_3650,N_3673);
nand U3976 (N_3976,N_3778,N_3762);
or U3977 (N_3977,N_3777,N_3606);
and U3978 (N_3978,N_3722,N_3694);
or U3979 (N_3979,N_3733,N_3688);
xor U3980 (N_3980,N_3645,N_3747);
nand U3981 (N_3981,N_3639,N_3602);
and U3982 (N_3982,N_3603,N_3654);
nor U3983 (N_3983,N_3695,N_3748);
or U3984 (N_3984,N_3638,N_3771);
nand U3985 (N_3985,N_3794,N_3770);
or U3986 (N_3986,N_3759,N_3720);
and U3987 (N_3987,N_3733,N_3601);
nor U3988 (N_3988,N_3666,N_3728);
or U3989 (N_3989,N_3748,N_3778);
or U3990 (N_3990,N_3714,N_3674);
nor U3991 (N_3991,N_3758,N_3780);
xor U3992 (N_3992,N_3708,N_3777);
nor U3993 (N_3993,N_3632,N_3772);
xor U3994 (N_3994,N_3793,N_3785);
nor U3995 (N_3995,N_3690,N_3673);
nand U3996 (N_3996,N_3749,N_3783);
or U3997 (N_3997,N_3767,N_3636);
or U3998 (N_3998,N_3694,N_3795);
or U3999 (N_3999,N_3618,N_3604);
nand U4000 (N_4000,N_3846,N_3973);
and U4001 (N_4001,N_3953,N_3954);
xor U4002 (N_4002,N_3955,N_3950);
nand U4003 (N_4003,N_3891,N_3952);
nor U4004 (N_4004,N_3989,N_3958);
or U4005 (N_4005,N_3892,N_3998);
nand U4006 (N_4006,N_3923,N_3865);
and U4007 (N_4007,N_3978,N_3844);
nor U4008 (N_4008,N_3984,N_3916);
nor U4009 (N_4009,N_3801,N_3999);
nand U4010 (N_4010,N_3841,N_3895);
nand U4011 (N_4011,N_3887,N_3960);
nor U4012 (N_4012,N_3969,N_3888);
nor U4013 (N_4013,N_3949,N_3871);
nand U4014 (N_4014,N_3864,N_3824);
or U4015 (N_4015,N_3970,N_3980);
nand U4016 (N_4016,N_3933,N_3802);
or U4017 (N_4017,N_3830,N_3991);
and U4018 (N_4018,N_3807,N_3927);
or U4019 (N_4019,N_3829,N_3917);
nand U4020 (N_4020,N_3948,N_3833);
xor U4021 (N_4021,N_3956,N_3805);
and U4022 (N_4022,N_3874,N_3913);
xnor U4023 (N_4023,N_3918,N_3907);
and U4024 (N_4024,N_3821,N_3834);
or U4025 (N_4025,N_3966,N_3890);
xor U4026 (N_4026,N_3808,N_3855);
nor U4027 (N_4027,N_3932,N_3873);
nand U4028 (N_4028,N_3868,N_3836);
nand U4029 (N_4029,N_3852,N_3814);
nor U4030 (N_4030,N_3972,N_3920);
nor U4031 (N_4031,N_3894,N_3809);
nor U4032 (N_4032,N_3912,N_3883);
and U4033 (N_4033,N_3854,N_3945);
nor U4034 (N_4034,N_3898,N_3908);
xor U4035 (N_4035,N_3951,N_3910);
and U4036 (N_4036,N_3828,N_3992);
nand U4037 (N_4037,N_3817,N_3982);
xor U4038 (N_4038,N_3939,N_3832);
and U4039 (N_4039,N_3938,N_3901);
nand U4040 (N_4040,N_3937,N_3911);
nand U4041 (N_4041,N_3922,N_3944);
and U4042 (N_4042,N_3831,N_3964);
nand U4043 (N_4043,N_3827,N_3947);
nand U4044 (N_4044,N_3959,N_3860);
nor U4045 (N_4045,N_3957,N_3993);
xor U4046 (N_4046,N_3995,N_3816);
or U4047 (N_4047,N_3915,N_3819);
or U4048 (N_4048,N_3988,N_3943);
nor U4049 (N_4049,N_3936,N_3847);
xnor U4050 (N_4050,N_3977,N_3946);
and U4051 (N_4051,N_3812,N_3983);
nor U4052 (N_4052,N_3879,N_3842);
nor U4053 (N_4053,N_3881,N_3840);
nor U4054 (N_4054,N_3906,N_3893);
or U4055 (N_4055,N_3843,N_3930);
nor U4056 (N_4056,N_3962,N_3997);
nand U4057 (N_4057,N_3961,N_3851);
and U4058 (N_4058,N_3872,N_3905);
or U4059 (N_4059,N_3928,N_3994);
nor U4060 (N_4060,N_3990,N_3974);
and U4061 (N_4061,N_3825,N_3903);
and U4062 (N_4062,N_3965,N_3979);
nand U4063 (N_4063,N_3925,N_3909);
nor U4064 (N_4064,N_3929,N_3835);
or U4065 (N_4065,N_3940,N_3934);
nand U4066 (N_4066,N_3976,N_3985);
nand U4067 (N_4067,N_3869,N_3889);
or U4068 (N_4068,N_3880,N_3803);
and U4069 (N_4069,N_3885,N_3882);
and U4070 (N_4070,N_3810,N_3813);
nand U4071 (N_4071,N_3820,N_3823);
xnor U4072 (N_4072,N_3826,N_3896);
and U4073 (N_4073,N_3987,N_3837);
and U4074 (N_4074,N_3902,N_3857);
or U4075 (N_4075,N_3996,N_3921);
xor U4076 (N_4076,N_3838,N_3876);
nand U4077 (N_4077,N_3877,N_3866);
nand U4078 (N_4078,N_3804,N_3870);
nand U4079 (N_4079,N_3818,N_3861);
xor U4080 (N_4080,N_3941,N_3968);
nand U4081 (N_4081,N_3863,N_3942);
nor U4082 (N_4082,N_3878,N_3867);
or U4083 (N_4083,N_3886,N_3963);
and U4084 (N_4084,N_3900,N_3845);
nor U4085 (N_4085,N_3862,N_3897);
or U4086 (N_4086,N_3884,N_3926);
and U4087 (N_4087,N_3899,N_3975);
and U4088 (N_4088,N_3919,N_3859);
nor U4089 (N_4089,N_3967,N_3815);
xor U4090 (N_4090,N_3931,N_3849);
and U4091 (N_4091,N_3822,N_3875);
nor U4092 (N_4092,N_3904,N_3924);
nand U4093 (N_4093,N_3858,N_3800);
nand U4094 (N_4094,N_3856,N_3981);
or U4095 (N_4095,N_3935,N_3853);
nand U4096 (N_4096,N_3839,N_3848);
nor U4097 (N_4097,N_3806,N_3986);
and U4098 (N_4098,N_3850,N_3811);
or U4099 (N_4099,N_3971,N_3914);
xor U4100 (N_4100,N_3921,N_3830);
nor U4101 (N_4101,N_3806,N_3811);
nand U4102 (N_4102,N_3897,N_3872);
nor U4103 (N_4103,N_3987,N_3831);
nand U4104 (N_4104,N_3804,N_3883);
xnor U4105 (N_4105,N_3966,N_3840);
nor U4106 (N_4106,N_3982,N_3924);
or U4107 (N_4107,N_3912,N_3939);
or U4108 (N_4108,N_3819,N_3832);
and U4109 (N_4109,N_3832,N_3869);
and U4110 (N_4110,N_3879,N_3901);
nand U4111 (N_4111,N_3888,N_3895);
nand U4112 (N_4112,N_3851,N_3947);
nor U4113 (N_4113,N_3851,N_3842);
xor U4114 (N_4114,N_3904,N_3847);
or U4115 (N_4115,N_3842,N_3839);
or U4116 (N_4116,N_3962,N_3955);
nand U4117 (N_4117,N_3863,N_3952);
or U4118 (N_4118,N_3968,N_3910);
or U4119 (N_4119,N_3896,N_3938);
xor U4120 (N_4120,N_3925,N_3842);
nor U4121 (N_4121,N_3820,N_3827);
nor U4122 (N_4122,N_3934,N_3994);
or U4123 (N_4123,N_3965,N_3875);
xor U4124 (N_4124,N_3888,N_3993);
and U4125 (N_4125,N_3817,N_3951);
or U4126 (N_4126,N_3874,N_3826);
and U4127 (N_4127,N_3942,N_3893);
nand U4128 (N_4128,N_3809,N_3976);
and U4129 (N_4129,N_3883,N_3907);
nand U4130 (N_4130,N_3915,N_3802);
nand U4131 (N_4131,N_3884,N_3835);
nand U4132 (N_4132,N_3866,N_3990);
nor U4133 (N_4133,N_3969,N_3881);
and U4134 (N_4134,N_3964,N_3877);
xnor U4135 (N_4135,N_3982,N_3820);
xor U4136 (N_4136,N_3882,N_3802);
xor U4137 (N_4137,N_3823,N_3813);
or U4138 (N_4138,N_3997,N_3931);
nand U4139 (N_4139,N_3869,N_3984);
xor U4140 (N_4140,N_3852,N_3880);
and U4141 (N_4141,N_3898,N_3867);
and U4142 (N_4142,N_3932,N_3813);
nand U4143 (N_4143,N_3837,N_3920);
or U4144 (N_4144,N_3976,N_3869);
nand U4145 (N_4145,N_3866,N_3885);
and U4146 (N_4146,N_3881,N_3880);
nor U4147 (N_4147,N_3830,N_3920);
xnor U4148 (N_4148,N_3944,N_3978);
nor U4149 (N_4149,N_3877,N_3887);
or U4150 (N_4150,N_3848,N_3864);
and U4151 (N_4151,N_3884,N_3979);
nor U4152 (N_4152,N_3866,N_3886);
or U4153 (N_4153,N_3809,N_3859);
or U4154 (N_4154,N_3838,N_3952);
nor U4155 (N_4155,N_3820,N_3975);
nand U4156 (N_4156,N_3944,N_3981);
nor U4157 (N_4157,N_3899,N_3994);
nand U4158 (N_4158,N_3958,N_3910);
nor U4159 (N_4159,N_3987,N_3872);
nand U4160 (N_4160,N_3858,N_3980);
and U4161 (N_4161,N_3901,N_3918);
or U4162 (N_4162,N_3852,N_3900);
nor U4163 (N_4163,N_3810,N_3956);
nor U4164 (N_4164,N_3915,N_3883);
and U4165 (N_4165,N_3879,N_3945);
and U4166 (N_4166,N_3922,N_3847);
nand U4167 (N_4167,N_3801,N_3836);
xnor U4168 (N_4168,N_3946,N_3816);
or U4169 (N_4169,N_3965,N_3822);
nor U4170 (N_4170,N_3810,N_3862);
and U4171 (N_4171,N_3946,N_3912);
xor U4172 (N_4172,N_3842,N_3830);
or U4173 (N_4173,N_3895,N_3900);
nand U4174 (N_4174,N_3871,N_3928);
nand U4175 (N_4175,N_3813,N_3875);
and U4176 (N_4176,N_3960,N_3866);
or U4177 (N_4177,N_3807,N_3925);
nor U4178 (N_4178,N_3845,N_3923);
xnor U4179 (N_4179,N_3956,N_3990);
and U4180 (N_4180,N_3936,N_3817);
or U4181 (N_4181,N_3997,N_3876);
and U4182 (N_4182,N_3836,N_3889);
nand U4183 (N_4183,N_3901,N_3990);
nand U4184 (N_4184,N_3802,N_3867);
and U4185 (N_4185,N_3860,N_3891);
nand U4186 (N_4186,N_3828,N_3958);
and U4187 (N_4187,N_3919,N_3863);
nor U4188 (N_4188,N_3922,N_3833);
nor U4189 (N_4189,N_3994,N_3988);
and U4190 (N_4190,N_3801,N_3883);
nand U4191 (N_4191,N_3843,N_3910);
and U4192 (N_4192,N_3931,N_3830);
nor U4193 (N_4193,N_3968,N_3872);
or U4194 (N_4194,N_3821,N_3818);
or U4195 (N_4195,N_3843,N_3936);
nor U4196 (N_4196,N_3863,N_3902);
nor U4197 (N_4197,N_3931,N_3971);
nor U4198 (N_4198,N_3856,N_3811);
nor U4199 (N_4199,N_3948,N_3944);
or U4200 (N_4200,N_4192,N_4143);
nor U4201 (N_4201,N_4125,N_4156);
nand U4202 (N_4202,N_4172,N_4046);
nor U4203 (N_4203,N_4187,N_4097);
or U4204 (N_4204,N_4113,N_4191);
or U4205 (N_4205,N_4152,N_4020);
or U4206 (N_4206,N_4195,N_4140);
and U4207 (N_4207,N_4110,N_4010);
nor U4208 (N_4208,N_4185,N_4069);
or U4209 (N_4209,N_4027,N_4164);
and U4210 (N_4210,N_4062,N_4009);
and U4211 (N_4211,N_4123,N_4112);
nand U4212 (N_4212,N_4126,N_4053);
and U4213 (N_4213,N_4129,N_4153);
nand U4214 (N_4214,N_4047,N_4144);
and U4215 (N_4215,N_4175,N_4000);
and U4216 (N_4216,N_4089,N_4006);
nand U4217 (N_4217,N_4190,N_4060);
nand U4218 (N_4218,N_4109,N_4163);
nand U4219 (N_4219,N_4077,N_4100);
and U4220 (N_4220,N_4173,N_4142);
and U4221 (N_4221,N_4134,N_4198);
or U4222 (N_4222,N_4167,N_4001);
xnor U4223 (N_4223,N_4122,N_4032);
or U4224 (N_4224,N_4029,N_4072);
xor U4225 (N_4225,N_4038,N_4042);
or U4226 (N_4226,N_4101,N_4007);
or U4227 (N_4227,N_4104,N_4075);
nor U4228 (N_4228,N_4111,N_4138);
nor U4229 (N_4229,N_4088,N_4155);
nand U4230 (N_4230,N_4068,N_4035);
and U4231 (N_4231,N_4085,N_4115);
or U4232 (N_4232,N_4074,N_4044);
xnor U4233 (N_4233,N_4061,N_4130);
nor U4234 (N_4234,N_4120,N_4067);
xor U4235 (N_4235,N_4082,N_4103);
nor U4236 (N_4236,N_4127,N_4018);
nand U4237 (N_4237,N_4124,N_4002);
or U4238 (N_4238,N_4117,N_4141);
nand U4239 (N_4239,N_4013,N_4108);
nand U4240 (N_4240,N_4146,N_4043);
xor U4241 (N_4241,N_4147,N_4178);
and U4242 (N_4242,N_4031,N_4080);
nand U4243 (N_4243,N_4090,N_4099);
and U4244 (N_4244,N_4193,N_4045);
or U4245 (N_4245,N_4168,N_4148);
nor U4246 (N_4246,N_4137,N_4011);
nand U4247 (N_4247,N_4086,N_4128);
or U4248 (N_4248,N_4041,N_4161);
nor U4249 (N_4249,N_4081,N_4183);
nand U4250 (N_4250,N_4024,N_4083);
nor U4251 (N_4251,N_4008,N_4057);
nor U4252 (N_4252,N_4188,N_4078);
xor U4253 (N_4253,N_4048,N_4119);
nor U4254 (N_4254,N_4151,N_4017);
xor U4255 (N_4255,N_4025,N_4165);
nor U4256 (N_4256,N_4073,N_4014);
and U4257 (N_4257,N_4087,N_4093);
and U4258 (N_4258,N_4154,N_4003);
nand U4259 (N_4259,N_4066,N_4037);
nor U4260 (N_4260,N_4034,N_4094);
nand U4261 (N_4261,N_4189,N_4054);
nor U4262 (N_4262,N_4065,N_4171);
and U4263 (N_4263,N_4040,N_4036);
and U4264 (N_4264,N_4004,N_4196);
nor U4265 (N_4265,N_4114,N_4170);
xor U4266 (N_4266,N_4118,N_4028);
nand U4267 (N_4267,N_4022,N_4106);
nand U4268 (N_4268,N_4182,N_4102);
and U4269 (N_4269,N_4012,N_4181);
or U4270 (N_4270,N_4158,N_4166);
nor U4271 (N_4271,N_4030,N_4105);
or U4272 (N_4272,N_4079,N_4092);
nand U4273 (N_4273,N_4063,N_4059);
nand U4274 (N_4274,N_4197,N_4159);
nand U4275 (N_4275,N_4064,N_4076);
and U4276 (N_4276,N_4095,N_4121);
nor U4277 (N_4277,N_4162,N_4132);
or U4278 (N_4278,N_4049,N_4005);
nand U4279 (N_4279,N_4026,N_4174);
xnor U4280 (N_4280,N_4039,N_4021);
nor U4281 (N_4281,N_4019,N_4139);
or U4282 (N_4282,N_4050,N_4194);
and U4283 (N_4283,N_4186,N_4145);
and U4284 (N_4284,N_4070,N_4051);
and U4285 (N_4285,N_4084,N_4058);
nand U4286 (N_4286,N_4016,N_4015);
and U4287 (N_4287,N_4150,N_4023);
nand U4288 (N_4288,N_4169,N_4199);
and U4289 (N_4289,N_4116,N_4033);
nand U4290 (N_4290,N_4098,N_4133);
nor U4291 (N_4291,N_4157,N_4180);
or U4292 (N_4292,N_4177,N_4179);
and U4293 (N_4293,N_4071,N_4091);
nand U4294 (N_4294,N_4131,N_4160);
nor U4295 (N_4295,N_4135,N_4136);
or U4296 (N_4296,N_4055,N_4184);
nand U4297 (N_4297,N_4149,N_4176);
or U4298 (N_4298,N_4056,N_4052);
nor U4299 (N_4299,N_4096,N_4107);
nand U4300 (N_4300,N_4146,N_4099);
and U4301 (N_4301,N_4092,N_4197);
nand U4302 (N_4302,N_4029,N_4171);
nand U4303 (N_4303,N_4061,N_4168);
and U4304 (N_4304,N_4027,N_4007);
or U4305 (N_4305,N_4112,N_4115);
xnor U4306 (N_4306,N_4002,N_4078);
or U4307 (N_4307,N_4055,N_4136);
nor U4308 (N_4308,N_4036,N_4103);
and U4309 (N_4309,N_4166,N_4124);
xor U4310 (N_4310,N_4087,N_4085);
or U4311 (N_4311,N_4146,N_4084);
nand U4312 (N_4312,N_4103,N_4113);
or U4313 (N_4313,N_4081,N_4040);
nand U4314 (N_4314,N_4148,N_4043);
nor U4315 (N_4315,N_4173,N_4148);
or U4316 (N_4316,N_4174,N_4024);
and U4317 (N_4317,N_4146,N_4123);
nand U4318 (N_4318,N_4178,N_4139);
and U4319 (N_4319,N_4192,N_4182);
and U4320 (N_4320,N_4180,N_4189);
or U4321 (N_4321,N_4039,N_4108);
xnor U4322 (N_4322,N_4155,N_4002);
and U4323 (N_4323,N_4161,N_4141);
nor U4324 (N_4324,N_4181,N_4159);
nand U4325 (N_4325,N_4026,N_4119);
nand U4326 (N_4326,N_4157,N_4020);
xnor U4327 (N_4327,N_4041,N_4160);
nand U4328 (N_4328,N_4174,N_4109);
nor U4329 (N_4329,N_4073,N_4043);
or U4330 (N_4330,N_4067,N_4193);
and U4331 (N_4331,N_4012,N_4047);
xor U4332 (N_4332,N_4076,N_4111);
and U4333 (N_4333,N_4186,N_4162);
nand U4334 (N_4334,N_4131,N_4033);
nor U4335 (N_4335,N_4150,N_4102);
and U4336 (N_4336,N_4008,N_4039);
xor U4337 (N_4337,N_4176,N_4161);
or U4338 (N_4338,N_4105,N_4018);
or U4339 (N_4339,N_4097,N_4134);
and U4340 (N_4340,N_4182,N_4152);
or U4341 (N_4341,N_4102,N_4069);
or U4342 (N_4342,N_4196,N_4179);
and U4343 (N_4343,N_4090,N_4044);
and U4344 (N_4344,N_4111,N_4170);
nor U4345 (N_4345,N_4104,N_4011);
nor U4346 (N_4346,N_4074,N_4165);
and U4347 (N_4347,N_4008,N_4014);
nor U4348 (N_4348,N_4023,N_4190);
nand U4349 (N_4349,N_4158,N_4051);
nor U4350 (N_4350,N_4038,N_4175);
or U4351 (N_4351,N_4146,N_4169);
nand U4352 (N_4352,N_4169,N_4194);
nand U4353 (N_4353,N_4136,N_4085);
nor U4354 (N_4354,N_4109,N_4161);
and U4355 (N_4355,N_4013,N_4014);
xnor U4356 (N_4356,N_4068,N_4088);
and U4357 (N_4357,N_4098,N_4190);
nor U4358 (N_4358,N_4089,N_4108);
and U4359 (N_4359,N_4185,N_4092);
xor U4360 (N_4360,N_4147,N_4049);
or U4361 (N_4361,N_4145,N_4116);
or U4362 (N_4362,N_4029,N_4175);
and U4363 (N_4363,N_4139,N_4062);
and U4364 (N_4364,N_4114,N_4089);
nor U4365 (N_4365,N_4069,N_4132);
and U4366 (N_4366,N_4016,N_4123);
nor U4367 (N_4367,N_4171,N_4022);
nand U4368 (N_4368,N_4165,N_4012);
and U4369 (N_4369,N_4081,N_4174);
nor U4370 (N_4370,N_4035,N_4078);
nor U4371 (N_4371,N_4009,N_4088);
xor U4372 (N_4372,N_4021,N_4042);
or U4373 (N_4373,N_4055,N_4084);
and U4374 (N_4374,N_4110,N_4015);
and U4375 (N_4375,N_4174,N_4029);
xor U4376 (N_4376,N_4028,N_4041);
xor U4377 (N_4377,N_4111,N_4062);
xnor U4378 (N_4378,N_4188,N_4131);
nor U4379 (N_4379,N_4137,N_4043);
xnor U4380 (N_4380,N_4141,N_4175);
xnor U4381 (N_4381,N_4038,N_4107);
or U4382 (N_4382,N_4114,N_4041);
and U4383 (N_4383,N_4117,N_4097);
nor U4384 (N_4384,N_4152,N_4168);
nand U4385 (N_4385,N_4186,N_4068);
nand U4386 (N_4386,N_4025,N_4184);
or U4387 (N_4387,N_4180,N_4181);
and U4388 (N_4388,N_4019,N_4094);
and U4389 (N_4389,N_4040,N_4124);
nor U4390 (N_4390,N_4176,N_4056);
nor U4391 (N_4391,N_4192,N_4152);
nor U4392 (N_4392,N_4022,N_4071);
nor U4393 (N_4393,N_4017,N_4132);
or U4394 (N_4394,N_4069,N_4019);
and U4395 (N_4395,N_4007,N_4023);
nor U4396 (N_4396,N_4081,N_4193);
or U4397 (N_4397,N_4177,N_4036);
nand U4398 (N_4398,N_4140,N_4153);
nand U4399 (N_4399,N_4030,N_4063);
nor U4400 (N_4400,N_4364,N_4213);
and U4401 (N_4401,N_4303,N_4291);
nor U4402 (N_4402,N_4356,N_4389);
or U4403 (N_4403,N_4396,N_4357);
and U4404 (N_4404,N_4289,N_4315);
or U4405 (N_4405,N_4381,N_4298);
xor U4406 (N_4406,N_4328,N_4290);
nand U4407 (N_4407,N_4386,N_4341);
nand U4408 (N_4408,N_4217,N_4243);
and U4409 (N_4409,N_4374,N_4241);
nand U4410 (N_4410,N_4220,N_4270);
nor U4411 (N_4411,N_4203,N_4311);
nor U4412 (N_4412,N_4344,N_4230);
or U4413 (N_4413,N_4295,N_4376);
nand U4414 (N_4414,N_4225,N_4262);
or U4415 (N_4415,N_4227,N_4255);
nor U4416 (N_4416,N_4369,N_4370);
and U4417 (N_4417,N_4308,N_4271);
and U4418 (N_4418,N_4246,N_4383);
or U4419 (N_4419,N_4379,N_4350);
nand U4420 (N_4420,N_4275,N_4274);
or U4421 (N_4421,N_4391,N_4380);
or U4422 (N_4422,N_4251,N_4318);
nor U4423 (N_4423,N_4222,N_4272);
or U4424 (N_4424,N_4362,N_4268);
nor U4425 (N_4425,N_4329,N_4278);
nor U4426 (N_4426,N_4221,N_4252);
or U4427 (N_4427,N_4332,N_4236);
nand U4428 (N_4428,N_4336,N_4306);
nand U4429 (N_4429,N_4353,N_4337);
nor U4430 (N_4430,N_4207,N_4216);
or U4431 (N_4431,N_4322,N_4257);
nand U4432 (N_4432,N_4265,N_4373);
and U4433 (N_4433,N_4202,N_4277);
nor U4434 (N_4434,N_4297,N_4247);
and U4435 (N_4435,N_4253,N_4313);
nor U4436 (N_4436,N_4205,N_4346);
and U4437 (N_4437,N_4288,N_4263);
nand U4438 (N_4438,N_4232,N_4248);
and U4439 (N_4439,N_4299,N_4280);
nand U4440 (N_4440,N_4384,N_4388);
or U4441 (N_4441,N_4365,N_4237);
nand U4442 (N_4442,N_4340,N_4325);
or U4443 (N_4443,N_4398,N_4385);
nand U4444 (N_4444,N_4208,N_4234);
or U4445 (N_4445,N_4375,N_4285);
nor U4446 (N_4446,N_4260,N_4201);
nand U4447 (N_4447,N_4267,N_4331);
nand U4448 (N_4448,N_4343,N_4371);
nor U4449 (N_4449,N_4397,N_4395);
and U4450 (N_4450,N_4347,N_4283);
nand U4451 (N_4451,N_4249,N_4309);
or U4452 (N_4452,N_4212,N_4273);
and U4453 (N_4453,N_4269,N_4352);
and U4454 (N_4454,N_4361,N_4228);
nor U4455 (N_4455,N_4394,N_4206);
or U4456 (N_4456,N_4215,N_4366);
xor U4457 (N_4457,N_4242,N_4360);
and U4458 (N_4458,N_4266,N_4226);
nand U4459 (N_4459,N_4312,N_4305);
nand U4460 (N_4460,N_4214,N_4256);
and U4461 (N_4461,N_4349,N_4233);
nand U4462 (N_4462,N_4279,N_4323);
nand U4463 (N_4463,N_4261,N_4304);
or U4464 (N_4464,N_4363,N_4209);
nand U4465 (N_4465,N_4334,N_4218);
nand U4466 (N_4466,N_4348,N_4200);
nand U4467 (N_4467,N_4382,N_4239);
nor U4468 (N_4468,N_4392,N_4368);
xnor U4469 (N_4469,N_4210,N_4335);
nand U4470 (N_4470,N_4301,N_4317);
nand U4471 (N_4471,N_4293,N_4399);
nor U4472 (N_4472,N_4287,N_4231);
nand U4473 (N_4473,N_4223,N_4393);
nor U4474 (N_4474,N_4286,N_4250);
nand U4475 (N_4475,N_4354,N_4367);
or U4476 (N_4476,N_4292,N_4338);
or U4477 (N_4477,N_4390,N_4320);
and U4478 (N_4478,N_4316,N_4281);
nand U4479 (N_4479,N_4204,N_4229);
and U4480 (N_4480,N_4264,N_4321);
and U4481 (N_4481,N_4211,N_4314);
or U4482 (N_4482,N_4240,N_4302);
and U4483 (N_4483,N_4342,N_4359);
and U4484 (N_4484,N_4235,N_4294);
nor U4485 (N_4485,N_4333,N_4238);
or U4486 (N_4486,N_4358,N_4387);
nand U4487 (N_4487,N_4339,N_4377);
nand U4488 (N_4488,N_4326,N_4245);
or U4489 (N_4489,N_4284,N_4351);
nand U4490 (N_4490,N_4307,N_4330);
nor U4491 (N_4491,N_4282,N_4345);
nor U4492 (N_4492,N_4244,N_4258);
nor U4493 (N_4493,N_4259,N_4319);
or U4494 (N_4494,N_4372,N_4276);
or U4495 (N_4495,N_4224,N_4355);
nor U4496 (N_4496,N_4254,N_4378);
or U4497 (N_4497,N_4296,N_4324);
nand U4498 (N_4498,N_4300,N_4219);
or U4499 (N_4499,N_4327,N_4310);
nand U4500 (N_4500,N_4256,N_4301);
nand U4501 (N_4501,N_4322,N_4360);
nor U4502 (N_4502,N_4223,N_4302);
xnor U4503 (N_4503,N_4350,N_4305);
and U4504 (N_4504,N_4373,N_4383);
and U4505 (N_4505,N_4320,N_4267);
nor U4506 (N_4506,N_4250,N_4379);
nor U4507 (N_4507,N_4395,N_4279);
or U4508 (N_4508,N_4364,N_4206);
or U4509 (N_4509,N_4273,N_4293);
nand U4510 (N_4510,N_4287,N_4353);
or U4511 (N_4511,N_4373,N_4237);
or U4512 (N_4512,N_4291,N_4344);
nand U4513 (N_4513,N_4236,N_4314);
or U4514 (N_4514,N_4261,N_4264);
and U4515 (N_4515,N_4246,N_4214);
and U4516 (N_4516,N_4299,N_4379);
nor U4517 (N_4517,N_4287,N_4398);
or U4518 (N_4518,N_4360,N_4249);
nor U4519 (N_4519,N_4207,N_4278);
nand U4520 (N_4520,N_4394,N_4357);
nand U4521 (N_4521,N_4248,N_4301);
nor U4522 (N_4522,N_4355,N_4329);
nand U4523 (N_4523,N_4387,N_4236);
nand U4524 (N_4524,N_4212,N_4230);
and U4525 (N_4525,N_4385,N_4330);
nand U4526 (N_4526,N_4279,N_4368);
xnor U4527 (N_4527,N_4325,N_4243);
nand U4528 (N_4528,N_4278,N_4244);
nor U4529 (N_4529,N_4269,N_4259);
xor U4530 (N_4530,N_4224,N_4352);
and U4531 (N_4531,N_4373,N_4389);
or U4532 (N_4532,N_4261,N_4381);
xor U4533 (N_4533,N_4371,N_4247);
nand U4534 (N_4534,N_4269,N_4206);
nor U4535 (N_4535,N_4345,N_4362);
nor U4536 (N_4536,N_4356,N_4376);
nor U4537 (N_4537,N_4253,N_4294);
nor U4538 (N_4538,N_4387,N_4356);
nor U4539 (N_4539,N_4320,N_4225);
and U4540 (N_4540,N_4315,N_4238);
and U4541 (N_4541,N_4349,N_4318);
nand U4542 (N_4542,N_4316,N_4306);
or U4543 (N_4543,N_4217,N_4309);
nor U4544 (N_4544,N_4360,N_4237);
xnor U4545 (N_4545,N_4299,N_4237);
and U4546 (N_4546,N_4276,N_4269);
xor U4547 (N_4547,N_4361,N_4243);
or U4548 (N_4548,N_4200,N_4294);
and U4549 (N_4549,N_4236,N_4341);
nor U4550 (N_4550,N_4338,N_4324);
and U4551 (N_4551,N_4216,N_4344);
nor U4552 (N_4552,N_4392,N_4374);
or U4553 (N_4553,N_4286,N_4313);
xnor U4554 (N_4554,N_4370,N_4321);
nor U4555 (N_4555,N_4252,N_4212);
nor U4556 (N_4556,N_4392,N_4268);
and U4557 (N_4557,N_4335,N_4260);
and U4558 (N_4558,N_4235,N_4251);
nand U4559 (N_4559,N_4273,N_4291);
nor U4560 (N_4560,N_4266,N_4282);
and U4561 (N_4561,N_4268,N_4351);
nand U4562 (N_4562,N_4233,N_4273);
nor U4563 (N_4563,N_4290,N_4227);
or U4564 (N_4564,N_4333,N_4285);
nor U4565 (N_4565,N_4290,N_4356);
and U4566 (N_4566,N_4261,N_4223);
nand U4567 (N_4567,N_4390,N_4234);
or U4568 (N_4568,N_4281,N_4326);
and U4569 (N_4569,N_4397,N_4237);
nor U4570 (N_4570,N_4245,N_4297);
and U4571 (N_4571,N_4303,N_4292);
nor U4572 (N_4572,N_4221,N_4265);
and U4573 (N_4573,N_4291,N_4395);
and U4574 (N_4574,N_4242,N_4373);
nor U4575 (N_4575,N_4390,N_4235);
and U4576 (N_4576,N_4384,N_4278);
nor U4577 (N_4577,N_4381,N_4204);
nor U4578 (N_4578,N_4331,N_4349);
and U4579 (N_4579,N_4384,N_4242);
or U4580 (N_4580,N_4226,N_4394);
nor U4581 (N_4581,N_4256,N_4235);
and U4582 (N_4582,N_4378,N_4364);
nand U4583 (N_4583,N_4260,N_4302);
nor U4584 (N_4584,N_4328,N_4269);
nor U4585 (N_4585,N_4369,N_4384);
nand U4586 (N_4586,N_4225,N_4340);
or U4587 (N_4587,N_4328,N_4276);
and U4588 (N_4588,N_4319,N_4364);
nand U4589 (N_4589,N_4313,N_4387);
nand U4590 (N_4590,N_4206,N_4369);
or U4591 (N_4591,N_4288,N_4267);
nor U4592 (N_4592,N_4260,N_4337);
and U4593 (N_4593,N_4374,N_4348);
and U4594 (N_4594,N_4391,N_4284);
and U4595 (N_4595,N_4285,N_4267);
nor U4596 (N_4596,N_4287,N_4308);
nand U4597 (N_4597,N_4277,N_4335);
or U4598 (N_4598,N_4394,N_4364);
nand U4599 (N_4599,N_4335,N_4217);
xor U4600 (N_4600,N_4513,N_4503);
or U4601 (N_4601,N_4588,N_4585);
nand U4602 (N_4602,N_4564,N_4426);
nor U4603 (N_4603,N_4582,N_4515);
nand U4604 (N_4604,N_4523,N_4591);
nor U4605 (N_4605,N_4490,N_4530);
or U4606 (N_4606,N_4406,N_4464);
xnor U4607 (N_4607,N_4492,N_4590);
nor U4608 (N_4608,N_4405,N_4495);
or U4609 (N_4609,N_4497,N_4470);
and U4610 (N_4610,N_4493,N_4430);
or U4611 (N_4611,N_4556,N_4504);
and U4612 (N_4612,N_4598,N_4593);
xor U4613 (N_4613,N_4473,N_4512);
nand U4614 (N_4614,N_4409,N_4579);
and U4615 (N_4615,N_4509,N_4531);
and U4616 (N_4616,N_4476,N_4547);
nand U4617 (N_4617,N_4510,N_4458);
nand U4618 (N_4618,N_4520,N_4465);
nor U4619 (N_4619,N_4437,N_4420);
nor U4620 (N_4620,N_4486,N_4533);
nand U4621 (N_4621,N_4545,N_4522);
and U4622 (N_4622,N_4500,N_4400);
nor U4623 (N_4623,N_4519,N_4407);
nor U4624 (N_4624,N_4537,N_4596);
nor U4625 (N_4625,N_4568,N_4505);
and U4626 (N_4626,N_4555,N_4548);
and U4627 (N_4627,N_4566,N_4471);
nand U4628 (N_4628,N_4488,N_4413);
nor U4629 (N_4629,N_4482,N_4587);
and U4630 (N_4630,N_4551,N_4485);
or U4631 (N_4631,N_4529,N_4434);
nor U4632 (N_4632,N_4542,N_4452);
nand U4633 (N_4633,N_4518,N_4421);
nor U4634 (N_4634,N_4438,N_4448);
xor U4635 (N_4635,N_4549,N_4416);
or U4636 (N_4636,N_4414,N_4472);
nand U4637 (N_4637,N_4573,N_4467);
xnor U4638 (N_4638,N_4535,N_4563);
nor U4639 (N_4639,N_4469,N_4418);
and U4640 (N_4640,N_4599,N_4571);
xnor U4641 (N_4641,N_4480,N_4450);
or U4642 (N_4642,N_4479,N_4457);
or U4643 (N_4643,N_4594,N_4511);
or U4644 (N_4644,N_4433,N_4578);
or U4645 (N_4645,N_4539,N_4461);
or U4646 (N_4646,N_4502,N_4570);
and U4647 (N_4647,N_4487,N_4552);
nor U4648 (N_4648,N_4595,N_4553);
or U4649 (N_4649,N_4419,N_4525);
nor U4650 (N_4650,N_4401,N_4475);
xnor U4651 (N_4651,N_4572,N_4466);
and U4652 (N_4652,N_4443,N_4454);
and U4653 (N_4653,N_4411,N_4481);
nand U4654 (N_4654,N_4489,N_4446);
xnor U4655 (N_4655,N_4415,N_4562);
and U4656 (N_4656,N_4417,N_4575);
or U4657 (N_4657,N_4567,N_4445);
and U4658 (N_4658,N_4569,N_4447);
xor U4659 (N_4659,N_4432,N_4439);
and U4660 (N_4660,N_4577,N_4514);
and U4661 (N_4661,N_4449,N_4423);
nor U4662 (N_4662,N_4554,N_4498);
nand U4663 (N_4663,N_4451,N_4477);
nor U4664 (N_4664,N_4410,N_4559);
nand U4665 (N_4665,N_4583,N_4455);
nand U4666 (N_4666,N_4544,N_4532);
nor U4667 (N_4667,N_4546,N_4483);
or U4668 (N_4668,N_4521,N_4494);
nand U4669 (N_4669,N_4534,N_4431);
nor U4670 (N_4670,N_4527,N_4404);
nor U4671 (N_4671,N_4462,N_4526);
or U4672 (N_4672,N_4536,N_4574);
nor U4673 (N_4673,N_4560,N_4425);
nand U4674 (N_4674,N_4581,N_4580);
or U4675 (N_4675,N_4441,N_4460);
or U4676 (N_4676,N_4584,N_4528);
nor U4677 (N_4677,N_4444,N_4435);
xnor U4678 (N_4678,N_4538,N_4589);
xor U4679 (N_4679,N_4403,N_4474);
nand U4680 (N_4680,N_4408,N_4484);
nand U4681 (N_4681,N_4456,N_4508);
or U4682 (N_4682,N_4436,N_4586);
or U4683 (N_4683,N_4428,N_4557);
and U4684 (N_4684,N_4459,N_4597);
and U4685 (N_4685,N_4499,N_4427);
nand U4686 (N_4686,N_4541,N_4543);
or U4687 (N_4687,N_4524,N_4453);
and U4688 (N_4688,N_4507,N_4429);
or U4689 (N_4689,N_4576,N_4592);
or U4690 (N_4690,N_4468,N_4565);
xor U4691 (N_4691,N_4442,N_4424);
and U4692 (N_4692,N_4506,N_4501);
xnor U4693 (N_4693,N_4550,N_4412);
or U4694 (N_4694,N_4491,N_4463);
nor U4695 (N_4695,N_4440,N_4496);
nor U4696 (N_4696,N_4517,N_4516);
nor U4697 (N_4697,N_4402,N_4558);
and U4698 (N_4698,N_4561,N_4478);
or U4699 (N_4699,N_4422,N_4540);
or U4700 (N_4700,N_4404,N_4576);
or U4701 (N_4701,N_4508,N_4495);
xor U4702 (N_4702,N_4421,N_4578);
nor U4703 (N_4703,N_4500,N_4593);
and U4704 (N_4704,N_4582,N_4530);
nand U4705 (N_4705,N_4523,N_4416);
and U4706 (N_4706,N_4423,N_4518);
or U4707 (N_4707,N_4569,N_4598);
nor U4708 (N_4708,N_4567,N_4472);
and U4709 (N_4709,N_4421,N_4403);
nor U4710 (N_4710,N_4583,N_4520);
nand U4711 (N_4711,N_4413,N_4594);
nand U4712 (N_4712,N_4566,N_4448);
nand U4713 (N_4713,N_4563,N_4544);
nor U4714 (N_4714,N_4422,N_4594);
xnor U4715 (N_4715,N_4473,N_4490);
and U4716 (N_4716,N_4589,N_4507);
nor U4717 (N_4717,N_4459,N_4517);
nor U4718 (N_4718,N_4592,N_4421);
nand U4719 (N_4719,N_4469,N_4455);
nor U4720 (N_4720,N_4410,N_4517);
or U4721 (N_4721,N_4520,N_4486);
nor U4722 (N_4722,N_4402,N_4453);
nand U4723 (N_4723,N_4579,N_4531);
nand U4724 (N_4724,N_4452,N_4413);
and U4725 (N_4725,N_4490,N_4459);
or U4726 (N_4726,N_4438,N_4449);
and U4727 (N_4727,N_4576,N_4584);
xnor U4728 (N_4728,N_4505,N_4403);
or U4729 (N_4729,N_4405,N_4542);
nand U4730 (N_4730,N_4588,N_4466);
nor U4731 (N_4731,N_4406,N_4490);
and U4732 (N_4732,N_4596,N_4495);
nand U4733 (N_4733,N_4581,N_4420);
and U4734 (N_4734,N_4530,N_4532);
nor U4735 (N_4735,N_4532,N_4492);
nor U4736 (N_4736,N_4550,N_4418);
or U4737 (N_4737,N_4490,N_4502);
and U4738 (N_4738,N_4434,N_4460);
or U4739 (N_4739,N_4405,N_4471);
nand U4740 (N_4740,N_4487,N_4500);
nand U4741 (N_4741,N_4461,N_4506);
xnor U4742 (N_4742,N_4438,N_4495);
nand U4743 (N_4743,N_4541,N_4570);
nand U4744 (N_4744,N_4531,N_4576);
and U4745 (N_4745,N_4553,N_4496);
and U4746 (N_4746,N_4483,N_4407);
or U4747 (N_4747,N_4476,N_4467);
or U4748 (N_4748,N_4470,N_4547);
or U4749 (N_4749,N_4535,N_4442);
nand U4750 (N_4750,N_4471,N_4505);
nand U4751 (N_4751,N_4437,N_4477);
xor U4752 (N_4752,N_4421,N_4591);
and U4753 (N_4753,N_4536,N_4493);
nor U4754 (N_4754,N_4544,N_4461);
nand U4755 (N_4755,N_4533,N_4577);
and U4756 (N_4756,N_4588,N_4510);
or U4757 (N_4757,N_4486,N_4494);
nand U4758 (N_4758,N_4477,N_4542);
or U4759 (N_4759,N_4520,N_4493);
and U4760 (N_4760,N_4563,N_4548);
nand U4761 (N_4761,N_4593,N_4477);
and U4762 (N_4762,N_4528,N_4498);
and U4763 (N_4763,N_4592,N_4468);
nand U4764 (N_4764,N_4435,N_4400);
and U4765 (N_4765,N_4541,N_4597);
and U4766 (N_4766,N_4474,N_4545);
nand U4767 (N_4767,N_4467,N_4462);
nand U4768 (N_4768,N_4567,N_4542);
xor U4769 (N_4769,N_4573,N_4462);
xnor U4770 (N_4770,N_4433,N_4571);
nor U4771 (N_4771,N_4489,N_4480);
or U4772 (N_4772,N_4569,N_4440);
nor U4773 (N_4773,N_4594,N_4487);
nor U4774 (N_4774,N_4524,N_4596);
nand U4775 (N_4775,N_4552,N_4538);
or U4776 (N_4776,N_4428,N_4477);
nor U4777 (N_4777,N_4536,N_4412);
and U4778 (N_4778,N_4590,N_4493);
nor U4779 (N_4779,N_4424,N_4402);
and U4780 (N_4780,N_4484,N_4540);
nor U4781 (N_4781,N_4436,N_4408);
or U4782 (N_4782,N_4433,N_4514);
and U4783 (N_4783,N_4484,N_4585);
and U4784 (N_4784,N_4414,N_4476);
or U4785 (N_4785,N_4556,N_4490);
nor U4786 (N_4786,N_4454,N_4497);
nand U4787 (N_4787,N_4537,N_4459);
nand U4788 (N_4788,N_4534,N_4570);
or U4789 (N_4789,N_4500,N_4442);
and U4790 (N_4790,N_4402,N_4477);
nand U4791 (N_4791,N_4430,N_4576);
nor U4792 (N_4792,N_4584,N_4580);
and U4793 (N_4793,N_4491,N_4404);
nand U4794 (N_4794,N_4432,N_4561);
nor U4795 (N_4795,N_4573,N_4583);
nand U4796 (N_4796,N_4535,N_4505);
nor U4797 (N_4797,N_4527,N_4586);
xnor U4798 (N_4798,N_4489,N_4472);
xor U4799 (N_4799,N_4490,N_4572);
nand U4800 (N_4800,N_4779,N_4682);
nand U4801 (N_4801,N_4751,N_4626);
nor U4802 (N_4802,N_4729,N_4747);
nand U4803 (N_4803,N_4683,N_4793);
nand U4804 (N_4804,N_4690,N_4776);
nor U4805 (N_4805,N_4780,N_4686);
nand U4806 (N_4806,N_4726,N_4764);
or U4807 (N_4807,N_4796,N_4749);
nor U4808 (N_4808,N_4705,N_4714);
nor U4809 (N_4809,N_4717,N_4752);
nor U4810 (N_4810,N_4720,N_4716);
xnor U4811 (N_4811,N_4711,N_4679);
and U4812 (N_4812,N_4708,N_4706);
and U4813 (N_4813,N_4658,N_4653);
nand U4814 (N_4814,N_4631,N_4629);
and U4815 (N_4815,N_4633,N_4732);
xnor U4816 (N_4816,N_4667,N_4661);
nand U4817 (N_4817,N_4638,N_4715);
or U4818 (N_4818,N_4784,N_4738);
nor U4819 (N_4819,N_4794,N_4725);
and U4820 (N_4820,N_4713,N_4703);
or U4821 (N_4821,N_4724,N_4628);
xor U4822 (N_4822,N_4759,N_4730);
and U4823 (N_4823,N_4662,N_4758);
nor U4824 (N_4824,N_4659,N_4689);
or U4825 (N_4825,N_4736,N_4742);
xor U4826 (N_4826,N_4616,N_4761);
xor U4827 (N_4827,N_4790,N_4684);
or U4828 (N_4828,N_4668,N_4657);
and U4829 (N_4829,N_4783,N_4606);
nor U4830 (N_4830,N_4673,N_4680);
and U4831 (N_4831,N_4767,N_4763);
or U4832 (N_4832,N_4798,N_4791);
xnor U4833 (N_4833,N_4670,N_4678);
or U4834 (N_4834,N_4632,N_4622);
nor U4835 (N_4835,N_4674,N_4733);
nand U4836 (N_4836,N_4727,N_4754);
xnor U4837 (N_4837,N_4701,N_4692);
xnor U4838 (N_4838,N_4617,N_4781);
nor U4839 (N_4839,N_4672,N_4619);
and U4840 (N_4840,N_4646,N_4637);
nor U4841 (N_4841,N_4797,N_4675);
xor U4842 (N_4842,N_4698,N_4602);
or U4843 (N_4843,N_4772,N_4723);
nand U4844 (N_4844,N_4748,N_4652);
nand U4845 (N_4845,N_4694,N_4750);
nand U4846 (N_4846,N_4787,N_4607);
nand U4847 (N_4847,N_4641,N_4687);
nand U4848 (N_4848,N_4696,N_4789);
or U4849 (N_4849,N_4697,N_4691);
nor U4850 (N_4850,N_4608,N_4665);
nor U4851 (N_4851,N_4688,N_4644);
and U4852 (N_4852,N_4639,N_4604);
nand U4853 (N_4853,N_4611,N_4768);
or U4854 (N_4854,N_4669,N_4785);
and U4855 (N_4855,N_4664,N_4634);
xnor U4856 (N_4856,N_4741,N_4745);
and U4857 (N_4857,N_4625,N_4609);
and U4858 (N_4858,N_4650,N_4719);
nand U4859 (N_4859,N_4766,N_4601);
nor U4860 (N_4860,N_4627,N_4778);
nand U4861 (N_4861,N_4677,N_4610);
and U4862 (N_4862,N_4605,N_4799);
and U4863 (N_4863,N_4621,N_4676);
xor U4864 (N_4864,N_4600,N_4615);
or U4865 (N_4865,N_4707,N_4651);
or U4866 (N_4866,N_4699,N_4795);
xnor U4867 (N_4867,N_4739,N_4718);
nor U4868 (N_4868,N_4695,N_4731);
xor U4869 (N_4869,N_4744,N_4735);
nor U4870 (N_4870,N_4775,N_4756);
nor U4871 (N_4871,N_4782,N_4612);
or U4872 (N_4872,N_4770,N_4649);
nand U4873 (N_4873,N_4613,N_4642);
nand U4874 (N_4874,N_4734,N_4693);
nand U4875 (N_4875,N_4762,N_4663);
or U4876 (N_4876,N_4618,N_4648);
nand U4877 (N_4877,N_4620,N_4722);
nor U4878 (N_4878,N_4666,N_4769);
and U4879 (N_4879,N_4753,N_4765);
or U4880 (N_4880,N_4774,N_4635);
or U4881 (N_4881,N_4623,N_4777);
xnor U4882 (N_4882,N_4728,N_4704);
and U4883 (N_4883,N_4786,N_4681);
nand U4884 (N_4884,N_4743,N_4773);
and U4885 (N_4885,N_4740,N_4700);
nor U4886 (N_4886,N_4645,N_4614);
xor U4887 (N_4887,N_4660,N_4671);
nor U4888 (N_4888,N_4643,N_4656);
and U4889 (N_4889,N_4630,N_4654);
nand U4890 (N_4890,N_4771,N_4603);
and U4891 (N_4891,N_4712,N_4640);
xor U4892 (N_4892,N_4647,N_4737);
xor U4893 (N_4893,N_4702,N_4624);
or U4894 (N_4894,N_4760,N_4636);
nor U4895 (N_4895,N_4755,N_4792);
and U4896 (N_4896,N_4746,N_4685);
nand U4897 (N_4897,N_4721,N_4709);
nand U4898 (N_4898,N_4757,N_4788);
nand U4899 (N_4899,N_4655,N_4710);
and U4900 (N_4900,N_4780,N_4696);
nor U4901 (N_4901,N_4678,N_4699);
nor U4902 (N_4902,N_4610,N_4652);
nand U4903 (N_4903,N_4694,N_4644);
xnor U4904 (N_4904,N_4623,N_4707);
and U4905 (N_4905,N_4720,N_4643);
and U4906 (N_4906,N_4795,N_4673);
and U4907 (N_4907,N_4775,N_4767);
xor U4908 (N_4908,N_4733,N_4625);
nor U4909 (N_4909,N_4766,N_4606);
or U4910 (N_4910,N_4670,N_4721);
or U4911 (N_4911,N_4770,N_4699);
nand U4912 (N_4912,N_4630,N_4726);
nand U4913 (N_4913,N_4737,N_4748);
and U4914 (N_4914,N_4735,N_4644);
and U4915 (N_4915,N_4679,N_4658);
and U4916 (N_4916,N_4692,N_4696);
or U4917 (N_4917,N_4648,N_4606);
xor U4918 (N_4918,N_4672,N_4661);
and U4919 (N_4919,N_4627,N_4798);
nand U4920 (N_4920,N_4725,N_4713);
or U4921 (N_4921,N_4699,N_4766);
nand U4922 (N_4922,N_4604,N_4749);
nand U4923 (N_4923,N_4670,N_4702);
xor U4924 (N_4924,N_4767,N_4667);
nand U4925 (N_4925,N_4717,N_4739);
xnor U4926 (N_4926,N_4703,N_4628);
nand U4927 (N_4927,N_4682,N_4647);
and U4928 (N_4928,N_4622,N_4771);
xor U4929 (N_4929,N_4613,N_4720);
nand U4930 (N_4930,N_4623,N_4666);
nand U4931 (N_4931,N_4728,N_4624);
nand U4932 (N_4932,N_4640,N_4715);
and U4933 (N_4933,N_4664,N_4790);
and U4934 (N_4934,N_4671,N_4796);
nor U4935 (N_4935,N_4659,N_4684);
and U4936 (N_4936,N_4746,N_4788);
nand U4937 (N_4937,N_4713,N_4775);
or U4938 (N_4938,N_4751,N_4711);
xnor U4939 (N_4939,N_4734,N_4786);
or U4940 (N_4940,N_4660,N_4622);
nor U4941 (N_4941,N_4752,N_4623);
nand U4942 (N_4942,N_4602,N_4616);
nor U4943 (N_4943,N_4778,N_4797);
nand U4944 (N_4944,N_4710,N_4794);
or U4945 (N_4945,N_4726,N_4698);
nand U4946 (N_4946,N_4619,N_4786);
and U4947 (N_4947,N_4795,N_4667);
nor U4948 (N_4948,N_4784,N_4668);
and U4949 (N_4949,N_4775,N_4654);
or U4950 (N_4950,N_4790,N_4744);
or U4951 (N_4951,N_4783,N_4760);
xor U4952 (N_4952,N_4661,N_4769);
or U4953 (N_4953,N_4646,N_4751);
xor U4954 (N_4954,N_4751,N_4655);
or U4955 (N_4955,N_4661,N_4765);
or U4956 (N_4956,N_4612,N_4631);
and U4957 (N_4957,N_4634,N_4799);
nor U4958 (N_4958,N_4644,N_4611);
or U4959 (N_4959,N_4678,N_4632);
or U4960 (N_4960,N_4797,N_4612);
nand U4961 (N_4961,N_4622,N_4681);
nand U4962 (N_4962,N_4698,N_4763);
nand U4963 (N_4963,N_4625,N_4645);
nand U4964 (N_4964,N_4610,N_4764);
or U4965 (N_4965,N_4782,N_4741);
or U4966 (N_4966,N_4722,N_4732);
nor U4967 (N_4967,N_4673,N_4683);
xnor U4968 (N_4968,N_4600,N_4748);
nor U4969 (N_4969,N_4640,N_4750);
nand U4970 (N_4970,N_4739,N_4725);
nand U4971 (N_4971,N_4712,N_4738);
nand U4972 (N_4972,N_4793,N_4782);
and U4973 (N_4973,N_4616,N_4788);
nand U4974 (N_4974,N_4634,N_4608);
nor U4975 (N_4975,N_4742,N_4759);
nand U4976 (N_4976,N_4715,N_4662);
xnor U4977 (N_4977,N_4643,N_4623);
and U4978 (N_4978,N_4711,N_4700);
and U4979 (N_4979,N_4692,N_4668);
nor U4980 (N_4980,N_4744,N_4691);
nand U4981 (N_4981,N_4678,N_4799);
and U4982 (N_4982,N_4692,N_4703);
and U4983 (N_4983,N_4687,N_4665);
and U4984 (N_4984,N_4624,N_4712);
xor U4985 (N_4985,N_4664,N_4723);
nand U4986 (N_4986,N_4692,N_4655);
or U4987 (N_4987,N_4664,N_4720);
nand U4988 (N_4988,N_4649,N_4743);
nand U4989 (N_4989,N_4637,N_4695);
or U4990 (N_4990,N_4645,N_4786);
xnor U4991 (N_4991,N_4753,N_4725);
or U4992 (N_4992,N_4611,N_4663);
and U4993 (N_4993,N_4678,N_4768);
xor U4994 (N_4994,N_4738,N_4672);
nor U4995 (N_4995,N_4662,N_4696);
or U4996 (N_4996,N_4742,N_4611);
and U4997 (N_4997,N_4676,N_4650);
xor U4998 (N_4998,N_4658,N_4628);
or U4999 (N_4999,N_4736,N_4642);
and U5000 (N_5000,N_4914,N_4850);
nand U5001 (N_5001,N_4978,N_4863);
nand U5002 (N_5002,N_4999,N_4980);
nand U5003 (N_5003,N_4841,N_4890);
and U5004 (N_5004,N_4936,N_4957);
nand U5005 (N_5005,N_4885,N_4874);
nand U5006 (N_5006,N_4814,N_4943);
and U5007 (N_5007,N_4831,N_4990);
and U5008 (N_5008,N_4838,N_4950);
and U5009 (N_5009,N_4899,N_4830);
or U5010 (N_5010,N_4949,N_4947);
nand U5011 (N_5011,N_4807,N_4816);
or U5012 (N_5012,N_4916,N_4925);
nand U5013 (N_5013,N_4989,N_4877);
or U5014 (N_5014,N_4854,N_4820);
nand U5015 (N_5015,N_4839,N_4963);
and U5016 (N_5016,N_4867,N_4888);
nand U5017 (N_5017,N_4840,N_4806);
nor U5018 (N_5018,N_4915,N_4905);
or U5019 (N_5019,N_4879,N_4804);
and U5020 (N_5020,N_4986,N_4895);
and U5021 (N_5021,N_4985,N_4842);
and U5022 (N_5022,N_4903,N_4945);
or U5023 (N_5023,N_4801,N_4852);
or U5024 (N_5024,N_4817,N_4984);
or U5025 (N_5025,N_4912,N_4901);
xor U5026 (N_5026,N_4876,N_4815);
xor U5027 (N_5027,N_4859,N_4952);
nor U5028 (N_5028,N_4971,N_4832);
nor U5029 (N_5029,N_4875,N_4848);
xnor U5030 (N_5030,N_4858,N_4828);
or U5031 (N_5031,N_4887,N_4956);
and U5032 (N_5032,N_4881,N_4974);
nand U5033 (N_5033,N_4853,N_4940);
nor U5034 (N_5034,N_4845,N_4997);
nor U5035 (N_5035,N_4871,N_4846);
and U5036 (N_5036,N_4923,N_4918);
or U5037 (N_5037,N_4900,N_4946);
or U5038 (N_5038,N_4958,N_4893);
and U5039 (N_5039,N_4995,N_4939);
and U5040 (N_5040,N_4926,N_4920);
nand U5041 (N_5041,N_4965,N_4913);
nor U5042 (N_5042,N_4886,N_4805);
and U5043 (N_5043,N_4860,N_4961);
or U5044 (N_5044,N_4812,N_4894);
nor U5045 (N_5045,N_4932,N_4970);
and U5046 (N_5046,N_4866,N_4937);
or U5047 (N_5047,N_4992,N_4891);
nand U5048 (N_5048,N_4968,N_4809);
nand U5049 (N_5049,N_4878,N_4954);
nand U5050 (N_5050,N_4959,N_4811);
or U5051 (N_5051,N_4967,N_4810);
nor U5052 (N_5052,N_4813,N_4896);
and U5053 (N_5053,N_4991,N_4802);
and U5054 (N_5054,N_4977,N_4909);
or U5055 (N_5055,N_4906,N_4969);
nor U5056 (N_5056,N_4982,N_4933);
nor U5057 (N_5057,N_4825,N_4836);
or U5058 (N_5058,N_4821,N_4919);
nor U5059 (N_5059,N_4833,N_4981);
nor U5060 (N_5060,N_4934,N_4953);
nand U5061 (N_5061,N_4979,N_4847);
or U5062 (N_5062,N_4998,N_4883);
xnor U5063 (N_5063,N_4921,N_4861);
nand U5064 (N_5064,N_4922,N_4824);
nand U5065 (N_5065,N_4819,N_4929);
nor U5066 (N_5066,N_4862,N_4851);
nor U5067 (N_5067,N_4892,N_4837);
or U5068 (N_5068,N_4962,N_4930);
and U5069 (N_5069,N_4955,N_4976);
nand U5070 (N_5070,N_4987,N_4988);
nand U5071 (N_5071,N_4849,N_4941);
nand U5072 (N_5072,N_4857,N_4873);
nor U5073 (N_5073,N_4931,N_4864);
nand U5074 (N_5074,N_4964,N_4823);
or U5075 (N_5075,N_4870,N_4884);
and U5076 (N_5076,N_4935,N_4902);
nor U5077 (N_5077,N_4924,N_4803);
or U5078 (N_5078,N_4898,N_4889);
nor U5079 (N_5079,N_4827,N_4983);
nor U5080 (N_5080,N_4856,N_4993);
or U5081 (N_5081,N_4822,N_4973);
nor U5082 (N_5082,N_4868,N_4869);
nand U5083 (N_5083,N_4917,N_4855);
xor U5084 (N_5084,N_4800,N_4818);
or U5085 (N_5085,N_4938,N_4835);
or U5086 (N_5086,N_4844,N_4910);
and U5087 (N_5087,N_4944,N_4808);
nor U5088 (N_5088,N_4927,N_4972);
nand U5089 (N_5089,N_4904,N_4975);
nand U5090 (N_5090,N_4960,N_4880);
xor U5091 (N_5091,N_4908,N_4829);
xnor U5092 (N_5092,N_4834,N_4911);
nand U5093 (N_5093,N_4907,N_4865);
xnor U5094 (N_5094,N_4996,N_4948);
or U5095 (N_5095,N_4994,N_4928);
nand U5096 (N_5096,N_4951,N_4826);
and U5097 (N_5097,N_4882,N_4897);
xnor U5098 (N_5098,N_4843,N_4872);
and U5099 (N_5099,N_4942,N_4966);
or U5100 (N_5100,N_4955,N_4823);
or U5101 (N_5101,N_4963,N_4808);
or U5102 (N_5102,N_4909,N_4857);
nand U5103 (N_5103,N_4864,N_4911);
and U5104 (N_5104,N_4982,N_4850);
xor U5105 (N_5105,N_4838,N_4998);
nand U5106 (N_5106,N_4838,N_4837);
nand U5107 (N_5107,N_4810,N_4983);
nand U5108 (N_5108,N_4915,N_4909);
or U5109 (N_5109,N_4814,N_4921);
nor U5110 (N_5110,N_4993,N_4808);
xor U5111 (N_5111,N_4936,N_4895);
nand U5112 (N_5112,N_4836,N_4833);
or U5113 (N_5113,N_4839,N_4820);
nor U5114 (N_5114,N_4997,N_4859);
or U5115 (N_5115,N_4847,N_4905);
xor U5116 (N_5116,N_4899,N_4805);
nor U5117 (N_5117,N_4965,N_4909);
or U5118 (N_5118,N_4880,N_4989);
nand U5119 (N_5119,N_4968,N_4845);
or U5120 (N_5120,N_4918,N_4843);
and U5121 (N_5121,N_4932,N_4925);
and U5122 (N_5122,N_4995,N_4933);
and U5123 (N_5123,N_4973,N_4945);
or U5124 (N_5124,N_4940,N_4950);
and U5125 (N_5125,N_4964,N_4947);
nand U5126 (N_5126,N_4964,N_4934);
nor U5127 (N_5127,N_4856,N_4808);
or U5128 (N_5128,N_4965,N_4978);
and U5129 (N_5129,N_4975,N_4886);
nand U5130 (N_5130,N_4877,N_4961);
nor U5131 (N_5131,N_4857,N_4867);
or U5132 (N_5132,N_4880,N_4866);
or U5133 (N_5133,N_4883,N_4877);
nand U5134 (N_5134,N_4843,N_4994);
and U5135 (N_5135,N_4866,N_4832);
nor U5136 (N_5136,N_4912,N_4837);
or U5137 (N_5137,N_4869,N_4954);
nor U5138 (N_5138,N_4845,N_4922);
xor U5139 (N_5139,N_4933,N_4918);
or U5140 (N_5140,N_4923,N_4941);
and U5141 (N_5141,N_4866,N_4924);
and U5142 (N_5142,N_4915,N_4997);
nor U5143 (N_5143,N_4877,N_4956);
nor U5144 (N_5144,N_4959,N_4974);
nor U5145 (N_5145,N_4876,N_4991);
nand U5146 (N_5146,N_4816,N_4947);
and U5147 (N_5147,N_4888,N_4834);
or U5148 (N_5148,N_4902,N_4889);
or U5149 (N_5149,N_4864,N_4808);
nor U5150 (N_5150,N_4897,N_4810);
or U5151 (N_5151,N_4988,N_4884);
nand U5152 (N_5152,N_4905,N_4812);
or U5153 (N_5153,N_4875,N_4945);
nor U5154 (N_5154,N_4939,N_4964);
nand U5155 (N_5155,N_4857,N_4889);
nand U5156 (N_5156,N_4992,N_4870);
nand U5157 (N_5157,N_4843,N_4931);
and U5158 (N_5158,N_4877,N_4910);
and U5159 (N_5159,N_4933,N_4990);
nand U5160 (N_5160,N_4980,N_4970);
xor U5161 (N_5161,N_4988,N_4926);
nand U5162 (N_5162,N_4837,N_4952);
or U5163 (N_5163,N_4914,N_4868);
or U5164 (N_5164,N_4892,N_4975);
nand U5165 (N_5165,N_4838,N_4903);
and U5166 (N_5166,N_4991,N_4949);
nor U5167 (N_5167,N_4912,N_4991);
or U5168 (N_5168,N_4814,N_4829);
or U5169 (N_5169,N_4969,N_4992);
nand U5170 (N_5170,N_4829,N_4885);
nand U5171 (N_5171,N_4924,N_4847);
xnor U5172 (N_5172,N_4917,N_4825);
nor U5173 (N_5173,N_4983,N_4851);
nor U5174 (N_5174,N_4852,N_4980);
nand U5175 (N_5175,N_4872,N_4806);
nand U5176 (N_5176,N_4929,N_4877);
nand U5177 (N_5177,N_4926,N_4973);
nor U5178 (N_5178,N_4827,N_4811);
or U5179 (N_5179,N_4955,N_4876);
and U5180 (N_5180,N_4857,N_4810);
nor U5181 (N_5181,N_4936,N_4852);
nor U5182 (N_5182,N_4949,N_4917);
nor U5183 (N_5183,N_4801,N_4872);
nor U5184 (N_5184,N_4890,N_4850);
and U5185 (N_5185,N_4973,N_4815);
or U5186 (N_5186,N_4999,N_4878);
and U5187 (N_5187,N_4990,N_4813);
and U5188 (N_5188,N_4946,N_4937);
nor U5189 (N_5189,N_4908,N_4825);
or U5190 (N_5190,N_4838,N_4925);
or U5191 (N_5191,N_4862,N_4972);
nand U5192 (N_5192,N_4883,N_4987);
nor U5193 (N_5193,N_4821,N_4842);
and U5194 (N_5194,N_4869,N_4932);
nand U5195 (N_5195,N_4995,N_4919);
and U5196 (N_5196,N_4943,N_4924);
nor U5197 (N_5197,N_4935,N_4993);
or U5198 (N_5198,N_4900,N_4847);
nand U5199 (N_5199,N_4881,N_4891);
or U5200 (N_5200,N_5188,N_5067);
xor U5201 (N_5201,N_5167,N_5115);
and U5202 (N_5202,N_5014,N_5000);
nor U5203 (N_5203,N_5120,N_5173);
and U5204 (N_5204,N_5160,N_5175);
or U5205 (N_5205,N_5084,N_5137);
nor U5206 (N_5206,N_5073,N_5028);
nor U5207 (N_5207,N_5124,N_5196);
nand U5208 (N_5208,N_5070,N_5020);
nand U5209 (N_5209,N_5030,N_5112);
or U5210 (N_5210,N_5139,N_5085);
and U5211 (N_5211,N_5176,N_5130);
and U5212 (N_5212,N_5123,N_5192);
nor U5213 (N_5213,N_5090,N_5093);
or U5214 (N_5214,N_5118,N_5079);
or U5215 (N_5215,N_5069,N_5190);
xnor U5216 (N_5216,N_5038,N_5143);
and U5217 (N_5217,N_5049,N_5193);
xnor U5218 (N_5218,N_5106,N_5055);
or U5219 (N_5219,N_5159,N_5078);
and U5220 (N_5220,N_5027,N_5184);
nand U5221 (N_5221,N_5061,N_5105);
or U5222 (N_5222,N_5097,N_5095);
nand U5223 (N_5223,N_5019,N_5145);
nand U5224 (N_5224,N_5074,N_5114);
nand U5225 (N_5225,N_5102,N_5004);
or U5226 (N_5226,N_5023,N_5082);
nor U5227 (N_5227,N_5109,N_5017);
nand U5228 (N_5228,N_5029,N_5146);
nand U5229 (N_5229,N_5001,N_5087);
nand U5230 (N_5230,N_5016,N_5153);
nand U5231 (N_5231,N_5044,N_5110);
or U5232 (N_5232,N_5009,N_5024);
and U5233 (N_5233,N_5062,N_5158);
or U5234 (N_5234,N_5104,N_5039);
and U5235 (N_5235,N_5101,N_5051);
nand U5236 (N_5236,N_5100,N_5040);
and U5237 (N_5237,N_5163,N_5053);
and U5238 (N_5238,N_5046,N_5125);
or U5239 (N_5239,N_5091,N_5180);
nand U5240 (N_5240,N_5177,N_5172);
and U5241 (N_5241,N_5077,N_5048);
or U5242 (N_5242,N_5005,N_5072);
nand U5243 (N_5243,N_5198,N_5058);
nand U5244 (N_5244,N_5128,N_5041);
nor U5245 (N_5245,N_5012,N_5047);
xor U5246 (N_5246,N_5168,N_5036);
or U5247 (N_5247,N_5018,N_5089);
and U5248 (N_5248,N_5189,N_5068);
or U5249 (N_5249,N_5026,N_5010);
nand U5250 (N_5250,N_5134,N_5197);
nor U5251 (N_5251,N_5013,N_5170);
and U5252 (N_5252,N_5194,N_5126);
nor U5253 (N_5253,N_5133,N_5144);
nor U5254 (N_5254,N_5081,N_5199);
nand U5255 (N_5255,N_5043,N_5065);
nand U5256 (N_5256,N_5156,N_5092);
or U5257 (N_5257,N_5025,N_5161);
nor U5258 (N_5258,N_5076,N_5136);
nand U5259 (N_5259,N_5154,N_5083);
xor U5260 (N_5260,N_5121,N_5096);
and U5261 (N_5261,N_5052,N_5182);
nor U5262 (N_5262,N_5155,N_5147);
nand U5263 (N_5263,N_5122,N_5116);
nand U5264 (N_5264,N_5185,N_5002);
and U5265 (N_5265,N_5056,N_5164);
or U5266 (N_5266,N_5015,N_5150);
and U5267 (N_5267,N_5045,N_5071);
or U5268 (N_5268,N_5127,N_5006);
and U5269 (N_5269,N_5035,N_5191);
and U5270 (N_5270,N_5003,N_5075);
xor U5271 (N_5271,N_5117,N_5108);
nand U5272 (N_5272,N_5099,N_5034);
xnor U5273 (N_5273,N_5008,N_5140);
and U5274 (N_5274,N_5094,N_5179);
or U5275 (N_5275,N_5011,N_5141);
or U5276 (N_5276,N_5022,N_5181);
nor U5277 (N_5277,N_5132,N_5166);
nor U5278 (N_5278,N_5171,N_5098);
or U5279 (N_5279,N_5064,N_5032);
and U5280 (N_5280,N_5059,N_5165);
nor U5281 (N_5281,N_5186,N_5111);
xnor U5282 (N_5282,N_5138,N_5054);
nand U5283 (N_5283,N_5178,N_5187);
or U5284 (N_5284,N_5149,N_5050);
and U5285 (N_5285,N_5021,N_5151);
or U5286 (N_5286,N_5080,N_5007);
or U5287 (N_5287,N_5033,N_5088);
nor U5288 (N_5288,N_5162,N_5057);
nand U5289 (N_5289,N_5148,N_5129);
nor U5290 (N_5290,N_5113,N_5037);
nand U5291 (N_5291,N_5131,N_5152);
xnor U5292 (N_5292,N_5086,N_5183);
nand U5293 (N_5293,N_5142,N_5169);
nor U5294 (N_5294,N_5195,N_5103);
and U5295 (N_5295,N_5042,N_5031);
xnor U5296 (N_5296,N_5157,N_5066);
and U5297 (N_5297,N_5107,N_5060);
nand U5298 (N_5298,N_5174,N_5063);
nor U5299 (N_5299,N_5119,N_5135);
nand U5300 (N_5300,N_5176,N_5109);
nor U5301 (N_5301,N_5039,N_5154);
and U5302 (N_5302,N_5173,N_5026);
nand U5303 (N_5303,N_5105,N_5010);
nand U5304 (N_5304,N_5176,N_5057);
and U5305 (N_5305,N_5029,N_5116);
nand U5306 (N_5306,N_5125,N_5180);
or U5307 (N_5307,N_5136,N_5011);
or U5308 (N_5308,N_5076,N_5087);
nand U5309 (N_5309,N_5015,N_5121);
or U5310 (N_5310,N_5029,N_5121);
and U5311 (N_5311,N_5017,N_5049);
nand U5312 (N_5312,N_5021,N_5006);
nand U5313 (N_5313,N_5034,N_5096);
and U5314 (N_5314,N_5183,N_5127);
or U5315 (N_5315,N_5078,N_5016);
nand U5316 (N_5316,N_5153,N_5035);
or U5317 (N_5317,N_5033,N_5045);
and U5318 (N_5318,N_5008,N_5161);
nor U5319 (N_5319,N_5193,N_5092);
nor U5320 (N_5320,N_5089,N_5145);
and U5321 (N_5321,N_5007,N_5184);
nand U5322 (N_5322,N_5034,N_5170);
xnor U5323 (N_5323,N_5001,N_5127);
nor U5324 (N_5324,N_5153,N_5117);
nor U5325 (N_5325,N_5113,N_5193);
or U5326 (N_5326,N_5128,N_5009);
nor U5327 (N_5327,N_5190,N_5005);
and U5328 (N_5328,N_5064,N_5068);
or U5329 (N_5329,N_5084,N_5136);
or U5330 (N_5330,N_5132,N_5004);
or U5331 (N_5331,N_5139,N_5013);
nor U5332 (N_5332,N_5006,N_5180);
nor U5333 (N_5333,N_5012,N_5063);
or U5334 (N_5334,N_5178,N_5110);
nand U5335 (N_5335,N_5025,N_5141);
nand U5336 (N_5336,N_5027,N_5199);
xnor U5337 (N_5337,N_5067,N_5143);
or U5338 (N_5338,N_5110,N_5015);
or U5339 (N_5339,N_5066,N_5067);
and U5340 (N_5340,N_5026,N_5086);
and U5341 (N_5341,N_5004,N_5070);
nand U5342 (N_5342,N_5122,N_5105);
nor U5343 (N_5343,N_5083,N_5169);
xnor U5344 (N_5344,N_5002,N_5059);
or U5345 (N_5345,N_5043,N_5018);
nor U5346 (N_5346,N_5012,N_5064);
nor U5347 (N_5347,N_5186,N_5100);
nand U5348 (N_5348,N_5067,N_5060);
xor U5349 (N_5349,N_5147,N_5121);
nand U5350 (N_5350,N_5101,N_5165);
nor U5351 (N_5351,N_5093,N_5162);
nor U5352 (N_5352,N_5089,N_5103);
nand U5353 (N_5353,N_5067,N_5152);
nand U5354 (N_5354,N_5135,N_5026);
and U5355 (N_5355,N_5171,N_5030);
nand U5356 (N_5356,N_5071,N_5198);
nand U5357 (N_5357,N_5011,N_5142);
nand U5358 (N_5358,N_5187,N_5181);
or U5359 (N_5359,N_5101,N_5045);
nand U5360 (N_5360,N_5063,N_5037);
and U5361 (N_5361,N_5022,N_5029);
nor U5362 (N_5362,N_5198,N_5088);
and U5363 (N_5363,N_5178,N_5072);
or U5364 (N_5364,N_5045,N_5104);
and U5365 (N_5365,N_5046,N_5081);
nand U5366 (N_5366,N_5156,N_5178);
and U5367 (N_5367,N_5079,N_5089);
or U5368 (N_5368,N_5139,N_5174);
and U5369 (N_5369,N_5017,N_5159);
nor U5370 (N_5370,N_5155,N_5034);
nand U5371 (N_5371,N_5130,N_5022);
nand U5372 (N_5372,N_5108,N_5140);
or U5373 (N_5373,N_5157,N_5003);
nand U5374 (N_5374,N_5071,N_5160);
and U5375 (N_5375,N_5031,N_5013);
and U5376 (N_5376,N_5051,N_5170);
nor U5377 (N_5377,N_5118,N_5049);
nand U5378 (N_5378,N_5156,N_5124);
nand U5379 (N_5379,N_5151,N_5161);
xor U5380 (N_5380,N_5122,N_5160);
or U5381 (N_5381,N_5188,N_5041);
or U5382 (N_5382,N_5065,N_5158);
nand U5383 (N_5383,N_5185,N_5128);
nor U5384 (N_5384,N_5125,N_5105);
nand U5385 (N_5385,N_5106,N_5111);
nor U5386 (N_5386,N_5095,N_5147);
nand U5387 (N_5387,N_5040,N_5120);
or U5388 (N_5388,N_5085,N_5038);
nor U5389 (N_5389,N_5154,N_5010);
and U5390 (N_5390,N_5056,N_5049);
nand U5391 (N_5391,N_5157,N_5176);
xnor U5392 (N_5392,N_5038,N_5111);
nand U5393 (N_5393,N_5147,N_5178);
nor U5394 (N_5394,N_5049,N_5066);
and U5395 (N_5395,N_5138,N_5106);
or U5396 (N_5396,N_5046,N_5179);
xnor U5397 (N_5397,N_5051,N_5124);
or U5398 (N_5398,N_5141,N_5160);
nand U5399 (N_5399,N_5043,N_5104);
and U5400 (N_5400,N_5277,N_5348);
nand U5401 (N_5401,N_5255,N_5359);
nand U5402 (N_5402,N_5232,N_5222);
xnor U5403 (N_5403,N_5272,N_5321);
or U5404 (N_5404,N_5227,N_5394);
and U5405 (N_5405,N_5373,N_5286);
and U5406 (N_5406,N_5289,N_5228);
and U5407 (N_5407,N_5204,N_5318);
nand U5408 (N_5408,N_5279,N_5396);
nor U5409 (N_5409,N_5284,N_5283);
or U5410 (N_5410,N_5266,N_5350);
or U5411 (N_5411,N_5238,N_5358);
and U5412 (N_5412,N_5211,N_5252);
or U5413 (N_5413,N_5292,N_5271);
nor U5414 (N_5414,N_5370,N_5345);
or U5415 (N_5415,N_5297,N_5319);
nor U5416 (N_5416,N_5260,N_5234);
and U5417 (N_5417,N_5285,N_5390);
nand U5418 (N_5418,N_5366,N_5282);
nand U5419 (N_5419,N_5332,N_5356);
nand U5420 (N_5420,N_5317,N_5273);
xnor U5421 (N_5421,N_5342,N_5290);
xor U5422 (N_5422,N_5361,N_5375);
and U5423 (N_5423,N_5258,N_5337);
or U5424 (N_5424,N_5347,N_5339);
or U5425 (N_5425,N_5214,N_5261);
or U5426 (N_5426,N_5300,N_5315);
nand U5427 (N_5427,N_5335,N_5326);
and U5428 (N_5428,N_5240,N_5386);
and U5429 (N_5429,N_5363,N_5309);
nor U5430 (N_5430,N_5262,N_5338);
nand U5431 (N_5431,N_5330,N_5333);
xor U5432 (N_5432,N_5298,N_5243);
nor U5433 (N_5433,N_5368,N_5295);
and U5434 (N_5434,N_5341,N_5387);
and U5435 (N_5435,N_5354,N_5274);
nand U5436 (N_5436,N_5372,N_5210);
and U5437 (N_5437,N_5294,N_5399);
xor U5438 (N_5438,N_5328,N_5220);
xor U5439 (N_5439,N_5205,N_5223);
xor U5440 (N_5440,N_5215,N_5235);
and U5441 (N_5441,N_5365,N_5381);
and U5442 (N_5442,N_5313,N_5382);
nor U5443 (N_5443,N_5376,N_5307);
nand U5444 (N_5444,N_5264,N_5320);
or U5445 (N_5445,N_5389,N_5362);
and U5446 (N_5446,N_5398,N_5249);
and U5447 (N_5447,N_5391,N_5208);
nand U5448 (N_5448,N_5340,N_5267);
nor U5449 (N_5449,N_5265,N_5242);
nand U5450 (N_5450,N_5247,N_5327);
or U5451 (N_5451,N_5275,N_5304);
nand U5452 (N_5452,N_5291,N_5241);
and U5453 (N_5453,N_5216,N_5237);
nor U5454 (N_5454,N_5256,N_5322);
and U5455 (N_5455,N_5226,N_5352);
nor U5456 (N_5456,N_5244,N_5357);
or U5457 (N_5457,N_5351,N_5236);
nor U5458 (N_5458,N_5306,N_5303);
nor U5459 (N_5459,N_5201,N_5325);
nor U5460 (N_5460,N_5224,N_5383);
and U5461 (N_5461,N_5207,N_5250);
and U5462 (N_5462,N_5344,N_5374);
nor U5463 (N_5463,N_5206,N_5203);
nand U5464 (N_5464,N_5378,N_5343);
nand U5465 (N_5465,N_5253,N_5248);
nand U5466 (N_5466,N_5349,N_5314);
nand U5467 (N_5467,N_5397,N_5288);
and U5468 (N_5468,N_5296,N_5225);
and U5469 (N_5469,N_5219,N_5209);
nor U5470 (N_5470,N_5246,N_5364);
nand U5471 (N_5471,N_5200,N_5212);
nand U5472 (N_5472,N_5281,N_5251);
nand U5473 (N_5473,N_5202,N_5287);
nand U5474 (N_5474,N_5346,N_5311);
nor U5475 (N_5475,N_5230,N_5324);
xnor U5476 (N_5476,N_5384,N_5329);
or U5477 (N_5477,N_5336,N_5257);
or U5478 (N_5478,N_5245,N_5395);
and U5479 (N_5479,N_5293,N_5388);
xnor U5480 (N_5480,N_5278,N_5269);
or U5481 (N_5481,N_5316,N_5323);
nand U5482 (N_5482,N_5231,N_5239);
xnor U5483 (N_5483,N_5301,N_5221);
nor U5484 (N_5484,N_5305,N_5392);
and U5485 (N_5485,N_5355,N_5308);
nor U5486 (N_5486,N_5334,N_5393);
or U5487 (N_5487,N_5377,N_5299);
or U5488 (N_5488,N_5259,N_5371);
or U5489 (N_5489,N_5310,N_5217);
nand U5490 (N_5490,N_5276,N_5302);
nor U5491 (N_5491,N_5367,N_5331);
nor U5492 (N_5492,N_5218,N_5280);
and U5493 (N_5493,N_5379,N_5213);
nor U5494 (N_5494,N_5229,N_5254);
xnor U5495 (N_5495,N_5360,N_5369);
nand U5496 (N_5496,N_5263,N_5268);
and U5497 (N_5497,N_5233,N_5353);
or U5498 (N_5498,N_5380,N_5385);
nand U5499 (N_5499,N_5312,N_5270);
nand U5500 (N_5500,N_5323,N_5232);
or U5501 (N_5501,N_5367,N_5303);
nor U5502 (N_5502,N_5209,N_5341);
and U5503 (N_5503,N_5206,N_5252);
xor U5504 (N_5504,N_5275,N_5225);
nand U5505 (N_5505,N_5390,N_5314);
xor U5506 (N_5506,N_5389,N_5396);
and U5507 (N_5507,N_5311,N_5309);
or U5508 (N_5508,N_5253,N_5295);
and U5509 (N_5509,N_5367,N_5376);
or U5510 (N_5510,N_5288,N_5286);
and U5511 (N_5511,N_5375,N_5380);
or U5512 (N_5512,N_5212,N_5369);
nand U5513 (N_5513,N_5200,N_5331);
nor U5514 (N_5514,N_5344,N_5228);
nor U5515 (N_5515,N_5282,N_5222);
nand U5516 (N_5516,N_5212,N_5258);
and U5517 (N_5517,N_5275,N_5338);
nand U5518 (N_5518,N_5359,N_5210);
nor U5519 (N_5519,N_5354,N_5394);
and U5520 (N_5520,N_5218,N_5227);
or U5521 (N_5521,N_5224,N_5389);
nor U5522 (N_5522,N_5241,N_5369);
or U5523 (N_5523,N_5230,N_5231);
xnor U5524 (N_5524,N_5361,N_5219);
nor U5525 (N_5525,N_5297,N_5374);
nand U5526 (N_5526,N_5224,N_5218);
and U5527 (N_5527,N_5314,N_5352);
and U5528 (N_5528,N_5352,N_5279);
nor U5529 (N_5529,N_5291,N_5301);
nor U5530 (N_5530,N_5278,N_5397);
or U5531 (N_5531,N_5341,N_5396);
and U5532 (N_5532,N_5256,N_5214);
or U5533 (N_5533,N_5254,N_5382);
or U5534 (N_5534,N_5262,N_5344);
or U5535 (N_5535,N_5342,N_5212);
or U5536 (N_5536,N_5220,N_5377);
nor U5537 (N_5537,N_5232,N_5290);
nand U5538 (N_5538,N_5377,N_5349);
or U5539 (N_5539,N_5265,N_5313);
nand U5540 (N_5540,N_5347,N_5399);
and U5541 (N_5541,N_5207,N_5386);
and U5542 (N_5542,N_5218,N_5257);
or U5543 (N_5543,N_5345,N_5262);
and U5544 (N_5544,N_5248,N_5362);
nand U5545 (N_5545,N_5259,N_5264);
nor U5546 (N_5546,N_5284,N_5346);
nor U5547 (N_5547,N_5307,N_5257);
xnor U5548 (N_5548,N_5212,N_5390);
or U5549 (N_5549,N_5326,N_5242);
and U5550 (N_5550,N_5281,N_5372);
and U5551 (N_5551,N_5276,N_5317);
nor U5552 (N_5552,N_5288,N_5373);
nor U5553 (N_5553,N_5222,N_5225);
nor U5554 (N_5554,N_5397,N_5370);
or U5555 (N_5555,N_5397,N_5373);
nor U5556 (N_5556,N_5242,N_5394);
nor U5557 (N_5557,N_5304,N_5281);
or U5558 (N_5558,N_5320,N_5254);
nand U5559 (N_5559,N_5316,N_5282);
or U5560 (N_5560,N_5322,N_5223);
or U5561 (N_5561,N_5324,N_5233);
and U5562 (N_5562,N_5287,N_5238);
nand U5563 (N_5563,N_5260,N_5204);
or U5564 (N_5564,N_5397,N_5345);
or U5565 (N_5565,N_5283,N_5306);
nand U5566 (N_5566,N_5338,N_5325);
nor U5567 (N_5567,N_5348,N_5325);
xnor U5568 (N_5568,N_5329,N_5215);
nor U5569 (N_5569,N_5330,N_5319);
and U5570 (N_5570,N_5220,N_5349);
and U5571 (N_5571,N_5250,N_5237);
and U5572 (N_5572,N_5254,N_5214);
and U5573 (N_5573,N_5238,N_5273);
or U5574 (N_5574,N_5310,N_5275);
and U5575 (N_5575,N_5275,N_5246);
nand U5576 (N_5576,N_5241,N_5267);
or U5577 (N_5577,N_5315,N_5229);
nor U5578 (N_5578,N_5317,N_5299);
and U5579 (N_5579,N_5399,N_5374);
and U5580 (N_5580,N_5209,N_5363);
nor U5581 (N_5581,N_5283,N_5218);
nand U5582 (N_5582,N_5319,N_5339);
or U5583 (N_5583,N_5398,N_5229);
or U5584 (N_5584,N_5259,N_5217);
nand U5585 (N_5585,N_5299,N_5206);
nor U5586 (N_5586,N_5224,N_5324);
xor U5587 (N_5587,N_5322,N_5305);
nor U5588 (N_5588,N_5273,N_5398);
or U5589 (N_5589,N_5295,N_5266);
and U5590 (N_5590,N_5276,N_5220);
or U5591 (N_5591,N_5205,N_5297);
nand U5592 (N_5592,N_5234,N_5331);
nand U5593 (N_5593,N_5278,N_5331);
nand U5594 (N_5594,N_5204,N_5233);
and U5595 (N_5595,N_5376,N_5245);
nor U5596 (N_5596,N_5343,N_5310);
or U5597 (N_5597,N_5318,N_5292);
xnor U5598 (N_5598,N_5318,N_5272);
nor U5599 (N_5599,N_5295,N_5312);
nand U5600 (N_5600,N_5434,N_5506);
and U5601 (N_5601,N_5420,N_5519);
nor U5602 (N_5602,N_5522,N_5439);
nor U5603 (N_5603,N_5440,N_5438);
nor U5604 (N_5604,N_5587,N_5413);
nor U5605 (N_5605,N_5436,N_5411);
nand U5606 (N_5606,N_5495,N_5516);
and U5607 (N_5607,N_5541,N_5469);
and U5608 (N_5608,N_5414,N_5509);
and U5609 (N_5609,N_5575,N_5498);
nand U5610 (N_5610,N_5504,N_5507);
nor U5611 (N_5611,N_5421,N_5456);
nor U5612 (N_5612,N_5583,N_5589);
nand U5613 (N_5613,N_5510,N_5481);
nor U5614 (N_5614,N_5511,N_5468);
nand U5615 (N_5615,N_5463,N_5544);
nor U5616 (N_5616,N_5465,N_5572);
nand U5617 (N_5617,N_5400,N_5447);
or U5618 (N_5618,N_5497,N_5462);
xor U5619 (N_5619,N_5599,N_5479);
and U5620 (N_5620,N_5426,N_5559);
nand U5621 (N_5621,N_5445,N_5480);
nor U5622 (N_5622,N_5531,N_5596);
nand U5623 (N_5623,N_5543,N_5492);
and U5624 (N_5624,N_5424,N_5533);
nand U5625 (N_5625,N_5483,N_5571);
and U5626 (N_5626,N_5521,N_5588);
nor U5627 (N_5627,N_5500,N_5488);
nor U5628 (N_5628,N_5432,N_5529);
or U5629 (N_5629,N_5402,N_5403);
or U5630 (N_5630,N_5406,N_5472);
or U5631 (N_5631,N_5470,N_5513);
or U5632 (N_5632,N_5429,N_5597);
nor U5633 (N_5633,N_5553,N_5476);
nor U5634 (N_5634,N_5530,N_5579);
xor U5635 (N_5635,N_5535,N_5525);
and U5636 (N_5636,N_5404,N_5561);
nand U5637 (N_5637,N_5407,N_5524);
nor U5638 (N_5638,N_5410,N_5556);
nand U5639 (N_5639,N_5508,N_5557);
nor U5640 (N_5640,N_5464,N_5582);
and U5641 (N_5641,N_5550,N_5489);
nor U5642 (N_5642,N_5409,N_5555);
and U5643 (N_5643,N_5460,N_5501);
and U5644 (N_5644,N_5592,N_5539);
xor U5645 (N_5645,N_5546,N_5598);
or U5646 (N_5646,N_5520,N_5514);
nor U5647 (N_5647,N_5570,N_5566);
nor U5648 (N_5648,N_5461,N_5534);
and U5649 (N_5649,N_5485,N_5585);
and U5650 (N_5650,N_5482,N_5532);
nand U5651 (N_5651,N_5528,N_5416);
or U5652 (N_5652,N_5450,N_5554);
or U5653 (N_5653,N_5423,N_5428);
and U5654 (N_5654,N_5569,N_5540);
or U5655 (N_5655,N_5549,N_5484);
and U5656 (N_5656,N_5491,N_5496);
nor U5657 (N_5657,N_5580,N_5446);
nand U5658 (N_5658,N_5593,N_5527);
or U5659 (N_5659,N_5515,N_5551);
or U5660 (N_5660,N_5591,N_5475);
nand U5661 (N_5661,N_5412,N_5408);
nand U5662 (N_5662,N_5454,N_5453);
nor U5663 (N_5663,N_5574,N_5590);
nor U5664 (N_5664,N_5562,N_5486);
nand U5665 (N_5665,N_5474,N_5537);
nand U5666 (N_5666,N_5435,N_5526);
nand U5667 (N_5667,N_5448,N_5564);
or U5668 (N_5668,N_5427,N_5422);
nand U5669 (N_5669,N_5443,N_5425);
nand U5670 (N_5670,N_5466,N_5471);
or U5671 (N_5671,N_5487,N_5577);
xnor U5672 (N_5672,N_5493,N_5467);
nor U5673 (N_5673,N_5536,N_5478);
and U5674 (N_5674,N_5584,N_5581);
xor U5675 (N_5675,N_5573,N_5494);
nor U5676 (N_5676,N_5594,N_5538);
and U5677 (N_5677,N_5563,N_5451);
and U5678 (N_5678,N_5512,N_5523);
nor U5679 (N_5679,N_5576,N_5567);
nor U5680 (N_5680,N_5452,N_5547);
nor U5681 (N_5681,N_5586,N_5401);
nand U5682 (N_5682,N_5545,N_5405);
nand U5683 (N_5683,N_5441,N_5442);
or U5684 (N_5684,N_5437,N_5565);
nor U5685 (N_5685,N_5542,N_5419);
xor U5686 (N_5686,N_5517,N_5415);
nand U5687 (N_5687,N_5502,N_5548);
nor U5688 (N_5688,N_5595,N_5455);
nand U5689 (N_5689,N_5578,N_5418);
or U5690 (N_5690,N_5560,N_5568);
or U5691 (N_5691,N_5477,N_5459);
xor U5692 (N_5692,N_5433,N_5558);
nand U5693 (N_5693,N_5473,N_5417);
nand U5694 (N_5694,N_5552,N_5499);
xor U5695 (N_5695,N_5490,N_5458);
xor U5696 (N_5696,N_5505,N_5457);
nor U5697 (N_5697,N_5444,N_5431);
nand U5698 (N_5698,N_5430,N_5503);
xor U5699 (N_5699,N_5518,N_5449);
or U5700 (N_5700,N_5576,N_5414);
xor U5701 (N_5701,N_5456,N_5490);
nor U5702 (N_5702,N_5509,N_5472);
nand U5703 (N_5703,N_5465,N_5412);
nor U5704 (N_5704,N_5568,N_5510);
nor U5705 (N_5705,N_5420,N_5558);
nor U5706 (N_5706,N_5549,N_5560);
or U5707 (N_5707,N_5425,N_5572);
xnor U5708 (N_5708,N_5463,N_5528);
or U5709 (N_5709,N_5509,N_5571);
and U5710 (N_5710,N_5487,N_5507);
nor U5711 (N_5711,N_5523,N_5454);
and U5712 (N_5712,N_5457,N_5436);
nand U5713 (N_5713,N_5443,N_5588);
nor U5714 (N_5714,N_5575,N_5584);
nor U5715 (N_5715,N_5451,N_5522);
or U5716 (N_5716,N_5545,N_5451);
nor U5717 (N_5717,N_5594,N_5442);
and U5718 (N_5718,N_5545,N_5486);
nor U5719 (N_5719,N_5479,N_5516);
nor U5720 (N_5720,N_5529,N_5416);
nand U5721 (N_5721,N_5588,N_5549);
nor U5722 (N_5722,N_5412,N_5496);
nand U5723 (N_5723,N_5559,N_5583);
or U5724 (N_5724,N_5458,N_5531);
and U5725 (N_5725,N_5461,N_5501);
nand U5726 (N_5726,N_5432,N_5479);
or U5727 (N_5727,N_5438,N_5482);
or U5728 (N_5728,N_5400,N_5414);
or U5729 (N_5729,N_5574,N_5511);
nand U5730 (N_5730,N_5447,N_5401);
and U5731 (N_5731,N_5525,N_5539);
nor U5732 (N_5732,N_5490,N_5449);
and U5733 (N_5733,N_5528,N_5422);
nand U5734 (N_5734,N_5464,N_5532);
nor U5735 (N_5735,N_5530,N_5528);
nand U5736 (N_5736,N_5563,N_5479);
or U5737 (N_5737,N_5488,N_5420);
or U5738 (N_5738,N_5519,N_5501);
or U5739 (N_5739,N_5428,N_5585);
nor U5740 (N_5740,N_5432,N_5453);
and U5741 (N_5741,N_5548,N_5415);
nand U5742 (N_5742,N_5531,N_5569);
xor U5743 (N_5743,N_5436,N_5535);
nand U5744 (N_5744,N_5512,N_5489);
nand U5745 (N_5745,N_5585,N_5595);
nand U5746 (N_5746,N_5593,N_5420);
nand U5747 (N_5747,N_5548,N_5511);
and U5748 (N_5748,N_5518,N_5555);
and U5749 (N_5749,N_5512,N_5575);
xor U5750 (N_5750,N_5432,N_5504);
and U5751 (N_5751,N_5512,N_5502);
and U5752 (N_5752,N_5468,N_5577);
and U5753 (N_5753,N_5458,N_5598);
and U5754 (N_5754,N_5410,N_5561);
and U5755 (N_5755,N_5564,N_5483);
and U5756 (N_5756,N_5572,N_5486);
and U5757 (N_5757,N_5436,N_5477);
or U5758 (N_5758,N_5581,N_5555);
or U5759 (N_5759,N_5489,N_5576);
and U5760 (N_5760,N_5536,N_5549);
nand U5761 (N_5761,N_5484,N_5410);
and U5762 (N_5762,N_5474,N_5542);
nand U5763 (N_5763,N_5430,N_5402);
nor U5764 (N_5764,N_5436,N_5434);
or U5765 (N_5765,N_5416,N_5559);
and U5766 (N_5766,N_5429,N_5478);
nand U5767 (N_5767,N_5528,N_5587);
nor U5768 (N_5768,N_5501,N_5416);
nand U5769 (N_5769,N_5545,N_5487);
and U5770 (N_5770,N_5544,N_5492);
and U5771 (N_5771,N_5445,N_5405);
nor U5772 (N_5772,N_5559,N_5526);
or U5773 (N_5773,N_5455,N_5594);
xnor U5774 (N_5774,N_5486,N_5435);
and U5775 (N_5775,N_5462,N_5510);
nand U5776 (N_5776,N_5491,N_5413);
nor U5777 (N_5777,N_5401,N_5427);
and U5778 (N_5778,N_5564,N_5472);
xor U5779 (N_5779,N_5497,N_5465);
or U5780 (N_5780,N_5547,N_5400);
or U5781 (N_5781,N_5425,N_5577);
nor U5782 (N_5782,N_5510,N_5514);
nor U5783 (N_5783,N_5535,N_5596);
xor U5784 (N_5784,N_5479,N_5445);
and U5785 (N_5785,N_5555,N_5418);
or U5786 (N_5786,N_5429,N_5461);
or U5787 (N_5787,N_5544,N_5464);
and U5788 (N_5788,N_5546,N_5497);
nand U5789 (N_5789,N_5439,N_5549);
nand U5790 (N_5790,N_5589,N_5581);
or U5791 (N_5791,N_5510,N_5439);
nand U5792 (N_5792,N_5424,N_5409);
or U5793 (N_5793,N_5592,N_5473);
or U5794 (N_5794,N_5563,N_5598);
and U5795 (N_5795,N_5527,N_5406);
nand U5796 (N_5796,N_5437,N_5448);
and U5797 (N_5797,N_5444,N_5406);
xor U5798 (N_5798,N_5570,N_5554);
nand U5799 (N_5799,N_5531,N_5512);
or U5800 (N_5800,N_5686,N_5754);
and U5801 (N_5801,N_5617,N_5658);
nand U5802 (N_5802,N_5719,N_5660);
nor U5803 (N_5803,N_5751,N_5772);
nand U5804 (N_5804,N_5694,N_5657);
and U5805 (N_5805,N_5625,N_5668);
or U5806 (N_5806,N_5642,N_5655);
nand U5807 (N_5807,N_5608,N_5680);
nand U5808 (N_5808,N_5693,N_5614);
nand U5809 (N_5809,N_5644,N_5741);
or U5810 (N_5810,N_5687,N_5723);
nor U5811 (N_5811,N_5663,N_5676);
xnor U5812 (N_5812,N_5633,N_5629);
or U5813 (N_5813,N_5696,N_5770);
nor U5814 (N_5814,N_5643,N_5649);
or U5815 (N_5815,N_5735,N_5626);
or U5816 (N_5816,N_5769,N_5775);
nor U5817 (N_5817,N_5677,N_5606);
or U5818 (N_5818,N_5797,N_5665);
nor U5819 (N_5819,N_5700,N_5776);
or U5820 (N_5820,N_5782,N_5604);
and U5821 (N_5821,N_5795,N_5793);
nor U5822 (N_5822,N_5777,N_5695);
nand U5823 (N_5823,N_5619,N_5618);
or U5824 (N_5824,N_5683,N_5717);
nand U5825 (N_5825,N_5673,N_5631);
and U5826 (N_5826,N_5790,N_5699);
nand U5827 (N_5827,N_5714,N_5771);
or U5828 (N_5828,N_5767,N_5786);
and U5829 (N_5829,N_5610,N_5798);
and U5830 (N_5830,N_5710,N_5706);
xor U5831 (N_5831,N_5750,N_5623);
nand U5832 (N_5832,N_5671,N_5742);
xnor U5833 (N_5833,N_5725,N_5622);
nand U5834 (N_5834,N_5749,N_5779);
nand U5835 (N_5835,N_5768,N_5731);
and U5836 (N_5836,N_5744,N_5627);
nand U5837 (N_5837,N_5661,N_5603);
xnor U5838 (N_5838,N_5791,N_5692);
nor U5839 (N_5839,N_5799,N_5654);
or U5840 (N_5840,N_5641,N_5716);
and U5841 (N_5841,N_5774,N_5702);
or U5842 (N_5842,N_5620,N_5624);
nor U5843 (N_5843,N_5781,N_5713);
or U5844 (N_5844,N_5728,N_5732);
or U5845 (N_5845,N_5762,N_5639);
and U5846 (N_5846,N_5647,N_5746);
nand U5847 (N_5847,N_5697,N_5794);
nand U5848 (N_5848,N_5729,N_5785);
and U5849 (N_5849,N_5783,N_5734);
or U5850 (N_5850,N_5612,N_5737);
and U5851 (N_5851,N_5602,N_5636);
xnor U5852 (N_5852,N_5712,N_5615);
and U5853 (N_5853,N_5659,N_5650);
or U5854 (N_5854,N_5711,N_5780);
nor U5855 (N_5855,N_5638,N_5730);
nor U5856 (N_5856,N_5652,N_5646);
and U5857 (N_5857,N_5698,N_5688);
and U5858 (N_5858,N_5709,N_5669);
nand U5859 (N_5859,N_5740,N_5681);
or U5860 (N_5860,N_5763,N_5758);
nor U5861 (N_5861,N_5648,N_5667);
nand U5862 (N_5862,N_5760,N_5664);
nand U5863 (N_5863,N_5672,N_5720);
or U5864 (N_5864,N_5611,N_5748);
nor U5865 (N_5865,N_5721,N_5651);
nand U5866 (N_5866,N_5628,N_5653);
nand U5867 (N_5867,N_5645,N_5609);
or U5868 (N_5868,N_5670,N_5705);
xnor U5869 (N_5869,N_5765,N_5784);
nand U5870 (N_5870,N_5759,N_5613);
and U5871 (N_5871,N_5722,N_5766);
xor U5872 (N_5872,N_5691,N_5707);
xnor U5873 (N_5873,N_5616,N_5736);
nor U5874 (N_5874,N_5752,N_5607);
and U5875 (N_5875,N_5685,N_5747);
nor U5876 (N_5876,N_5733,N_5789);
nor U5877 (N_5877,N_5632,N_5764);
and U5878 (N_5878,N_5755,N_5708);
nand U5879 (N_5879,N_5678,N_5684);
or U5880 (N_5880,N_5757,N_5718);
and U5881 (N_5881,N_5689,N_5682);
nor U5882 (N_5882,N_5662,N_5724);
nand U5883 (N_5883,N_5787,N_5656);
and U5884 (N_5884,N_5679,N_5600);
and U5885 (N_5885,N_5792,N_5778);
nor U5886 (N_5886,N_5605,N_5703);
nand U5887 (N_5887,N_5761,N_5726);
or U5888 (N_5888,N_5690,N_5743);
nand U5889 (N_5889,N_5704,N_5701);
or U5890 (N_5890,N_5753,N_5756);
nor U5891 (N_5891,N_5796,N_5634);
or U5892 (N_5892,N_5635,N_5715);
or U5893 (N_5893,N_5630,N_5666);
nand U5894 (N_5894,N_5773,N_5745);
and U5895 (N_5895,N_5601,N_5637);
and U5896 (N_5896,N_5727,N_5621);
nand U5897 (N_5897,N_5675,N_5640);
and U5898 (N_5898,N_5788,N_5674);
and U5899 (N_5899,N_5739,N_5738);
and U5900 (N_5900,N_5721,N_5625);
nand U5901 (N_5901,N_5790,N_5683);
nand U5902 (N_5902,N_5757,N_5735);
nor U5903 (N_5903,N_5602,N_5695);
or U5904 (N_5904,N_5731,N_5781);
nor U5905 (N_5905,N_5723,N_5732);
or U5906 (N_5906,N_5611,N_5603);
nor U5907 (N_5907,N_5796,N_5623);
nand U5908 (N_5908,N_5755,N_5642);
and U5909 (N_5909,N_5633,N_5648);
nor U5910 (N_5910,N_5721,N_5668);
or U5911 (N_5911,N_5672,N_5768);
nor U5912 (N_5912,N_5616,N_5755);
or U5913 (N_5913,N_5704,N_5637);
nor U5914 (N_5914,N_5687,N_5646);
and U5915 (N_5915,N_5692,N_5709);
nor U5916 (N_5916,N_5760,N_5679);
and U5917 (N_5917,N_5671,N_5619);
and U5918 (N_5918,N_5648,N_5745);
nand U5919 (N_5919,N_5613,N_5676);
nor U5920 (N_5920,N_5795,N_5783);
nor U5921 (N_5921,N_5720,N_5789);
or U5922 (N_5922,N_5647,N_5765);
nand U5923 (N_5923,N_5692,N_5610);
xnor U5924 (N_5924,N_5791,N_5785);
or U5925 (N_5925,N_5656,N_5781);
nor U5926 (N_5926,N_5741,N_5634);
xnor U5927 (N_5927,N_5660,N_5784);
nor U5928 (N_5928,N_5787,N_5753);
and U5929 (N_5929,N_5772,N_5736);
or U5930 (N_5930,N_5708,N_5662);
nand U5931 (N_5931,N_5686,N_5662);
and U5932 (N_5932,N_5656,N_5686);
and U5933 (N_5933,N_5664,N_5754);
nand U5934 (N_5934,N_5690,N_5794);
xnor U5935 (N_5935,N_5691,N_5790);
or U5936 (N_5936,N_5749,N_5772);
nand U5937 (N_5937,N_5710,N_5776);
and U5938 (N_5938,N_5706,N_5601);
or U5939 (N_5939,N_5627,N_5786);
and U5940 (N_5940,N_5797,N_5788);
or U5941 (N_5941,N_5775,N_5703);
nand U5942 (N_5942,N_5674,N_5692);
nand U5943 (N_5943,N_5686,N_5767);
and U5944 (N_5944,N_5672,N_5756);
nor U5945 (N_5945,N_5619,N_5710);
or U5946 (N_5946,N_5686,N_5750);
and U5947 (N_5947,N_5619,N_5605);
nor U5948 (N_5948,N_5646,N_5610);
and U5949 (N_5949,N_5635,N_5619);
or U5950 (N_5950,N_5651,N_5754);
nor U5951 (N_5951,N_5774,N_5708);
and U5952 (N_5952,N_5786,N_5728);
nor U5953 (N_5953,N_5742,N_5747);
or U5954 (N_5954,N_5600,N_5699);
nor U5955 (N_5955,N_5772,N_5724);
or U5956 (N_5956,N_5757,N_5647);
or U5957 (N_5957,N_5605,N_5729);
nor U5958 (N_5958,N_5714,N_5617);
nand U5959 (N_5959,N_5686,N_5735);
and U5960 (N_5960,N_5739,N_5786);
or U5961 (N_5961,N_5603,N_5679);
nand U5962 (N_5962,N_5771,N_5631);
nor U5963 (N_5963,N_5715,N_5723);
and U5964 (N_5964,N_5795,N_5717);
or U5965 (N_5965,N_5763,N_5673);
and U5966 (N_5966,N_5695,N_5689);
xnor U5967 (N_5967,N_5761,N_5778);
or U5968 (N_5968,N_5792,N_5767);
nand U5969 (N_5969,N_5705,N_5650);
nor U5970 (N_5970,N_5780,N_5645);
and U5971 (N_5971,N_5609,N_5706);
nand U5972 (N_5972,N_5670,N_5731);
nor U5973 (N_5973,N_5689,N_5728);
nand U5974 (N_5974,N_5689,N_5700);
or U5975 (N_5975,N_5699,N_5784);
and U5976 (N_5976,N_5697,N_5600);
and U5977 (N_5977,N_5775,N_5620);
nor U5978 (N_5978,N_5689,N_5794);
or U5979 (N_5979,N_5723,N_5793);
nor U5980 (N_5980,N_5783,N_5641);
nor U5981 (N_5981,N_5626,N_5791);
nand U5982 (N_5982,N_5633,N_5780);
and U5983 (N_5983,N_5684,N_5799);
nand U5984 (N_5984,N_5666,N_5757);
nand U5985 (N_5985,N_5623,N_5754);
and U5986 (N_5986,N_5606,N_5696);
xor U5987 (N_5987,N_5724,N_5633);
nor U5988 (N_5988,N_5653,N_5639);
nor U5989 (N_5989,N_5681,N_5798);
and U5990 (N_5990,N_5732,N_5674);
and U5991 (N_5991,N_5622,N_5746);
nand U5992 (N_5992,N_5722,N_5619);
and U5993 (N_5993,N_5641,N_5639);
and U5994 (N_5994,N_5605,N_5763);
and U5995 (N_5995,N_5733,N_5659);
and U5996 (N_5996,N_5773,N_5720);
nand U5997 (N_5997,N_5705,N_5674);
xor U5998 (N_5998,N_5723,N_5740);
or U5999 (N_5999,N_5782,N_5623);
and U6000 (N_6000,N_5984,N_5989);
nor U6001 (N_6001,N_5837,N_5969);
or U6002 (N_6002,N_5971,N_5929);
and U6003 (N_6003,N_5890,N_5871);
and U6004 (N_6004,N_5909,N_5950);
nand U6005 (N_6005,N_5846,N_5867);
and U6006 (N_6006,N_5964,N_5901);
xor U6007 (N_6007,N_5982,N_5931);
and U6008 (N_6008,N_5810,N_5852);
nor U6009 (N_6009,N_5943,N_5900);
nor U6010 (N_6010,N_5829,N_5895);
nor U6011 (N_6011,N_5862,N_5975);
nor U6012 (N_6012,N_5991,N_5802);
and U6013 (N_6013,N_5869,N_5819);
nor U6014 (N_6014,N_5844,N_5960);
or U6015 (N_6015,N_5826,N_5833);
nor U6016 (N_6016,N_5908,N_5997);
nor U6017 (N_6017,N_5841,N_5903);
or U6018 (N_6018,N_5805,N_5992);
or U6019 (N_6019,N_5899,N_5861);
nor U6020 (N_6020,N_5917,N_5998);
or U6021 (N_6021,N_5912,N_5881);
xor U6022 (N_6022,N_5876,N_5967);
and U6023 (N_6023,N_5849,N_5985);
nor U6024 (N_6024,N_5886,N_5811);
or U6025 (N_6025,N_5949,N_5814);
or U6026 (N_6026,N_5916,N_5934);
or U6027 (N_6027,N_5994,N_5956);
or U6028 (N_6028,N_5965,N_5959);
and U6029 (N_6029,N_5990,N_5866);
or U6030 (N_6030,N_5968,N_5888);
or U6031 (N_6031,N_5887,N_5944);
and U6032 (N_6032,N_5856,N_5945);
nor U6033 (N_6033,N_5999,N_5882);
nand U6034 (N_6034,N_5865,N_5958);
nand U6035 (N_6035,N_5995,N_5822);
nor U6036 (N_6036,N_5878,N_5806);
nand U6037 (N_6037,N_5891,N_5921);
and U6038 (N_6038,N_5868,N_5920);
nor U6039 (N_6039,N_5962,N_5823);
or U6040 (N_6040,N_5848,N_5840);
or U6041 (N_6041,N_5941,N_5813);
nor U6042 (N_6042,N_5948,N_5818);
nor U6043 (N_6043,N_5863,N_5854);
nand U6044 (N_6044,N_5880,N_5904);
nor U6045 (N_6045,N_5864,N_5923);
or U6046 (N_6046,N_5815,N_5963);
or U6047 (N_6047,N_5850,N_5966);
nor U6048 (N_6048,N_5947,N_5843);
or U6049 (N_6049,N_5970,N_5807);
or U6050 (N_6050,N_5932,N_5927);
and U6051 (N_6051,N_5896,N_5816);
and U6052 (N_6052,N_5834,N_5853);
and U6053 (N_6053,N_5938,N_5922);
nor U6054 (N_6054,N_5800,N_5855);
nand U6055 (N_6055,N_5809,N_5979);
nand U6056 (N_6056,N_5894,N_5919);
nor U6057 (N_6057,N_5851,N_5859);
nand U6058 (N_6058,N_5924,N_5911);
or U6059 (N_6059,N_5925,N_5845);
nand U6060 (N_6060,N_5928,N_5936);
xor U6061 (N_6061,N_5832,N_5996);
or U6062 (N_6062,N_5884,N_5972);
and U6063 (N_6063,N_5801,N_5892);
or U6064 (N_6064,N_5827,N_5951);
and U6065 (N_6065,N_5906,N_5812);
nor U6066 (N_6066,N_5898,N_5980);
or U6067 (N_6067,N_5926,N_5933);
nand U6068 (N_6068,N_5847,N_5993);
or U6069 (N_6069,N_5874,N_5976);
nor U6070 (N_6070,N_5877,N_5803);
nor U6071 (N_6071,N_5952,N_5954);
xnor U6072 (N_6072,N_5937,N_5957);
nor U6073 (N_6073,N_5913,N_5820);
nand U6074 (N_6074,N_5838,N_5873);
nor U6075 (N_6075,N_5981,N_5883);
or U6076 (N_6076,N_5930,N_5987);
nand U6077 (N_6077,N_5824,N_5889);
nor U6078 (N_6078,N_5872,N_5860);
or U6079 (N_6079,N_5918,N_5978);
nor U6080 (N_6080,N_5910,N_5983);
nand U6081 (N_6081,N_5988,N_5817);
and U6082 (N_6082,N_5885,N_5905);
xor U6083 (N_6083,N_5935,N_5828);
xnor U6084 (N_6084,N_5825,N_5942);
or U6085 (N_6085,N_5808,N_5879);
or U6086 (N_6086,N_5839,N_5835);
nor U6087 (N_6087,N_5939,N_5875);
and U6088 (N_6088,N_5955,N_5907);
nand U6089 (N_6089,N_5973,N_5977);
or U6090 (N_6090,N_5836,N_5974);
or U6091 (N_6091,N_5914,N_5940);
nor U6092 (N_6092,N_5821,N_5953);
nor U6093 (N_6093,N_5857,N_5986);
nor U6094 (N_6094,N_5858,N_5915);
and U6095 (N_6095,N_5842,N_5893);
and U6096 (N_6096,N_5831,N_5946);
or U6097 (N_6097,N_5897,N_5870);
nand U6098 (N_6098,N_5804,N_5830);
xnor U6099 (N_6099,N_5961,N_5902);
nor U6100 (N_6100,N_5872,N_5928);
or U6101 (N_6101,N_5861,N_5877);
and U6102 (N_6102,N_5809,N_5910);
xnor U6103 (N_6103,N_5926,N_5974);
xor U6104 (N_6104,N_5919,N_5824);
nor U6105 (N_6105,N_5803,N_5989);
nor U6106 (N_6106,N_5970,N_5814);
and U6107 (N_6107,N_5809,N_5948);
xnor U6108 (N_6108,N_5871,N_5807);
nor U6109 (N_6109,N_5866,N_5872);
nand U6110 (N_6110,N_5800,N_5864);
or U6111 (N_6111,N_5960,N_5870);
and U6112 (N_6112,N_5987,N_5943);
and U6113 (N_6113,N_5913,N_5824);
and U6114 (N_6114,N_5802,N_5932);
nor U6115 (N_6115,N_5944,N_5839);
and U6116 (N_6116,N_5827,N_5938);
or U6117 (N_6117,N_5929,N_5811);
nor U6118 (N_6118,N_5982,N_5897);
nor U6119 (N_6119,N_5829,N_5978);
nor U6120 (N_6120,N_5811,N_5959);
nor U6121 (N_6121,N_5867,N_5891);
nand U6122 (N_6122,N_5889,N_5821);
and U6123 (N_6123,N_5802,N_5801);
nor U6124 (N_6124,N_5985,N_5807);
nand U6125 (N_6125,N_5946,N_5965);
nor U6126 (N_6126,N_5977,N_5995);
nand U6127 (N_6127,N_5938,N_5931);
or U6128 (N_6128,N_5933,N_5874);
xor U6129 (N_6129,N_5848,N_5831);
nor U6130 (N_6130,N_5869,N_5836);
nand U6131 (N_6131,N_5901,N_5936);
and U6132 (N_6132,N_5955,N_5986);
nor U6133 (N_6133,N_5995,N_5921);
nand U6134 (N_6134,N_5817,N_5872);
nor U6135 (N_6135,N_5872,N_5870);
xor U6136 (N_6136,N_5906,N_5996);
and U6137 (N_6137,N_5988,N_5978);
and U6138 (N_6138,N_5821,N_5845);
and U6139 (N_6139,N_5974,N_5896);
nand U6140 (N_6140,N_5879,N_5933);
nor U6141 (N_6141,N_5863,N_5814);
nor U6142 (N_6142,N_5839,N_5989);
and U6143 (N_6143,N_5936,N_5866);
or U6144 (N_6144,N_5806,N_5854);
nor U6145 (N_6145,N_5809,N_5966);
or U6146 (N_6146,N_5832,N_5876);
or U6147 (N_6147,N_5971,N_5999);
xnor U6148 (N_6148,N_5981,N_5857);
xnor U6149 (N_6149,N_5986,N_5938);
and U6150 (N_6150,N_5977,N_5813);
or U6151 (N_6151,N_5849,N_5815);
nor U6152 (N_6152,N_5853,N_5817);
or U6153 (N_6153,N_5988,N_5837);
and U6154 (N_6154,N_5865,N_5964);
nand U6155 (N_6155,N_5842,N_5870);
nand U6156 (N_6156,N_5926,N_5832);
nor U6157 (N_6157,N_5818,N_5823);
xnor U6158 (N_6158,N_5996,N_5955);
or U6159 (N_6159,N_5990,N_5974);
nor U6160 (N_6160,N_5968,N_5856);
nor U6161 (N_6161,N_5968,N_5929);
and U6162 (N_6162,N_5889,N_5812);
xor U6163 (N_6163,N_5968,N_5971);
nand U6164 (N_6164,N_5977,N_5840);
or U6165 (N_6165,N_5987,N_5942);
or U6166 (N_6166,N_5952,N_5953);
nor U6167 (N_6167,N_5917,N_5928);
or U6168 (N_6168,N_5805,N_5917);
nand U6169 (N_6169,N_5840,N_5934);
xnor U6170 (N_6170,N_5974,N_5934);
or U6171 (N_6171,N_5876,N_5854);
or U6172 (N_6172,N_5885,N_5862);
nand U6173 (N_6173,N_5904,N_5946);
nand U6174 (N_6174,N_5978,N_5939);
or U6175 (N_6175,N_5957,N_5929);
nand U6176 (N_6176,N_5966,N_5836);
or U6177 (N_6177,N_5923,N_5825);
nor U6178 (N_6178,N_5830,N_5870);
and U6179 (N_6179,N_5935,N_5938);
nand U6180 (N_6180,N_5836,N_5856);
nor U6181 (N_6181,N_5933,N_5991);
xor U6182 (N_6182,N_5995,N_5842);
or U6183 (N_6183,N_5901,N_5985);
nor U6184 (N_6184,N_5919,N_5884);
nor U6185 (N_6185,N_5842,N_5896);
and U6186 (N_6186,N_5802,N_5917);
xor U6187 (N_6187,N_5975,N_5860);
and U6188 (N_6188,N_5838,N_5875);
and U6189 (N_6189,N_5876,N_5919);
nand U6190 (N_6190,N_5963,N_5927);
xnor U6191 (N_6191,N_5846,N_5912);
nand U6192 (N_6192,N_5851,N_5893);
or U6193 (N_6193,N_5903,N_5943);
and U6194 (N_6194,N_5922,N_5874);
or U6195 (N_6195,N_5858,N_5965);
or U6196 (N_6196,N_5954,N_5911);
or U6197 (N_6197,N_5990,N_5971);
or U6198 (N_6198,N_5977,N_5998);
nand U6199 (N_6199,N_5800,N_5962);
nand U6200 (N_6200,N_6101,N_6022);
nand U6201 (N_6201,N_6154,N_6125);
xor U6202 (N_6202,N_6082,N_6121);
or U6203 (N_6203,N_6053,N_6138);
and U6204 (N_6204,N_6198,N_6040);
nor U6205 (N_6205,N_6073,N_6019);
or U6206 (N_6206,N_6185,N_6192);
and U6207 (N_6207,N_6176,N_6106);
or U6208 (N_6208,N_6095,N_6130);
or U6209 (N_6209,N_6084,N_6134);
xor U6210 (N_6210,N_6144,N_6177);
nand U6211 (N_6211,N_6039,N_6173);
nand U6212 (N_6212,N_6074,N_6030);
nand U6213 (N_6213,N_6048,N_6007);
nand U6214 (N_6214,N_6104,N_6175);
nor U6215 (N_6215,N_6029,N_6140);
or U6216 (N_6216,N_6115,N_6066);
and U6217 (N_6217,N_6117,N_6085);
or U6218 (N_6218,N_6190,N_6124);
nand U6219 (N_6219,N_6118,N_6102);
nor U6220 (N_6220,N_6052,N_6027);
and U6221 (N_6221,N_6145,N_6083);
nor U6222 (N_6222,N_6188,N_6093);
xor U6223 (N_6223,N_6096,N_6132);
nand U6224 (N_6224,N_6010,N_6142);
xor U6225 (N_6225,N_6090,N_6133);
and U6226 (N_6226,N_6072,N_6076);
nand U6227 (N_6227,N_6161,N_6024);
or U6228 (N_6228,N_6005,N_6150);
or U6229 (N_6229,N_6146,N_6080);
nand U6230 (N_6230,N_6127,N_6119);
or U6231 (N_6231,N_6172,N_6179);
nor U6232 (N_6232,N_6041,N_6191);
nand U6233 (N_6233,N_6032,N_6160);
and U6234 (N_6234,N_6178,N_6078);
nor U6235 (N_6235,N_6086,N_6062);
and U6236 (N_6236,N_6038,N_6165);
nand U6237 (N_6237,N_6169,N_6186);
nor U6238 (N_6238,N_6061,N_6114);
nor U6239 (N_6239,N_6045,N_6153);
and U6240 (N_6240,N_6120,N_6049);
nor U6241 (N_6241,N_6158,N_6189);
or U6242 (N_6242,N_6050,N_6099);
xnor U6243 (N_6243,N_6111,N_6094);
or U6244 (N_6244,N_6021,N_6064);
or U6245 (N_6245,N_6129,N_6092);
nor U6246 (N_6246,N_6157,N_6008);
nand U6247 (N_6247,N_6028,N_6059);
or U6248 (N_6248,N_6057,N_6156);
or U6249 (N_6249,N_6167,N_6025);
or U6250 (N_6250,N_6164,N_6143);
nor U6251 (N_6251,N_6199,N_6098);
or U6252 (N_6252,N_6103,N_6141);
nor U6253 (N_6253,N_6004,N_6105);
and U6254 (N_6254,N_6126,N_6071);
nand U6255 (N_6255,N_6148,N_6136);
nor U6256 (N_6256,N_6170,N_6168);
or U6257 (N_6257,N_6108,N_6152);
xor U6258 (N_6258,N_6075,N_6110);
or U6259 (N_6259,N_6012,N_6014);
and U6260 (N_6260,N_6006,N_6036);
or U6261 (N_6261,N_6003,N_6034);
nand U6262 (N_6262,N_6013,N_6079);
nand U6263 (N_6263,N_6107,N_6183);
nand U6264 (N_6264,N_6026,N_6000);
xor U6265 (N_6265,N_6051,N_6044);
nor U6266 (N_6266,N_6155,N_6097);
or U6267 (N_6267,N_6017,N_6151);
xor U6268 (N_6268,N_6055,N_6011);
nand U6269 (N_6269,N_6109,N_6182);
nor U6270 (N_6270,N_6187,N_6058);
or U6271 (N_6271,N_6002,N_6122);
nand U6272 (N_6272,N_6171,N_6087);
xnor U6273 (N_6273,N_6162,N_6068);
xnor U6274 (N_6274,N_6091,N_6077);
and U6275 (N_6275,N_6047,N_6056);
and U6276 (N_6276,N_6197,N_6139);
nor U6277 (N_6277,N_6020,N_6149);
and U6278 (N_6278,N_6174,N_6116);
or U6279 (N_6279,N_6100,N_6015);
and U6280 (N_6280,N_6046,N_6031);
and U6281 (N_6281,N_6131,N_6037);
nand U6282 (N_6282,N_6042,N_6193);
and U6283 (N_6283,N_6196,N_6033);
or U6284 (N_6284,N_6018,N_6060);
or U6285 (N_6285,N_6184,N_6054);
nor U6286 (N_6286,N_6112,N_6016);
xor U6287 (N_6287,N_6043,N_6181);
or U6288 (N_6288,N_6135,N_6195);
or U6289 (N_6289,N_6001,N_6023);
nand U6290 (N_6290,N_6035,N_6137);
and U6291 (N_6291,N_6159,N_6088);
nor U6292 (N_6292,N_6166,N_6113);
and U6293 (N_6293,N_6147,N_6081);
or U6294 (N_6294,N_6180,N_6123);
or U6295 (N_6295,N_6069,N_6194);
nand U6296 (N_6296,N_6128,N_6067);
or U6297 (N_6297,N_6070,N_6065);
or U6298 (N_6298,N_6063,N_6163);
nor U6299 (N_6299,N_6089,N_6009);
or U6300 (N_6300,N_6056,N_6137);
and U6301 (N_6301,N_6112,N_6010);
nand U6302 (N_6302,N_6173,N_6075);
nor U6303 (N_6303,N_6183,N_6074);
nand U6304 (N_6304,N_6059,N_6160);
xor U6305 (N_6305,N_6025,N_6127);
or U6306 (N_6306,N_6034,N_6112);
or U6307 (N_6307,N_6119,N_6186);
and U6308 (N_6308,N_6093,N_6156);
or U6309 (N_6309,N_6157,N_6095);
or U6310 (N_6310,N_6159,N_6144);
or U6311 (N_6311,N_6149,N_6135);
or U6312 (N_6312,N_6155,N_6060);
and U6313 (N_6313,N_6181,N_6148);
or U6314 (N_6314,N_6037,N_6128);
nand U6315 (N_6315,N_6173,N_6143);
or U6316 (N_6316,N_6009,N_6114);
nand U6317 (N_6317,N_6051,N_6095);
and U6318 (N_6318,N_6017,N_6058);
and U6319 (N_6319,N_6087,N_6023);
or U6320 (N_6320,N_6083,N_6177);
nor U6321 (N_6321,N_6004,N_6019);
or U6322 (N_6322,N_6164,N_6026);
nand U6323 (N_6323,N_6136,N_6196);
and U6324 (N_6324,N_6074,N_6099);
and U6325 (N_6325,N_6120,N_6199);
or U6326 (N_6326,N_6075,N_6041);
and U6327 (N_6327,N_6041,N_6180);
or U6328 (N_6328,N_6153,N_6008);
nor U6329 (N_6329,N_6061,N_6094);
or U6330 (N_6330,N_6156,N_6060);
and U6331 (N_6331,N_6100,N_6052);
nor U6332 (N_6332,N_6088,N_6075);
and U6333 (N_6333,N_6185,N_6005);
or U6334 (N_6334,N_6075,N_6103);
nand U6335 (N_6335,N_6091,N_6195);
nand U6336 (N_6336,N_6055,N_6113);
or U6337 (N_6337,N_6198,N_6168);
nand U6338 (N_6338,N_6160,N_6073);
nand U6339 (N_6339,N_6179,N_6123);
and U6340 (N_6340,N_6018,N_6077);
nand U6341 (N_6341,N_6078,N_6073);
and U6342 (N_6342,N_6031,N_6025);
nor U6343 (N_6343,N_6095,N_6109);
nand U6344 (N_6344,N_6147,N_6028);
xnor U6345 (N_6345,N_6051,N_6192);
nor U6346 (N_6346,N_6153,N_6113);
nand U6347 (N_6347,N_6032,N_6102);
nand U6348 (N_6348,N_6191,N_6150);
or U6349 (N_6349,N_6146,N_6145);
and U6350 (N_6350,N_6090,N_6057);
nand U6351 (N_6351,N_6090,N_6168);
and U6352 (N_6352,N_6018,N_6143);
nand U6353 (N_6353,N_6062,N_6045);
nor U6354 (N_6354,N_6006,N_6126);
or U6355 (N_6355,N_6047,N_6140);
nand U6356 (N_6356,N_6097,N_6123);
and U6357 (N_6357,N_6174,N_6040);
or U6358 (N_6358,N_6137,N_6071);
or U6359 (N_6359,N_6167,N_6091);
and U6360 (N_6360,N_6167,N_6163);
or U6361 (N_6361,N_6033,N_6076);
nand U6362 (N_6362,N_6151,N_6069);
or U6363 (N_6363,N_6107,N_6119);
nand U6364 (N_6364,N_6169,N_6175);
or U6365 (N_6365,N_6197,N_6140);
or U6366 (N_6366,N_6006,N_6148);
nand U6367 (N_6367,N_6052,N_6049);
nor U6368 (N_6368,N_6045,N_6056);
xnor U6369 (N_6369,N_6022,N_6017);
xor U6370 (N_6370,N_6012,N_6182);
and U6371 (N_6371,N_6102,N_6124);
and U6372 (N_6372,N_6193,N_6155);
nand U6373 (N_6373,N_6164,N_6094);
and U6374 (N_6374,N_6181,N_6055);
nor U6375 (N_6375,N_6048,N_6102);
nand U6376 (N_6376,N_6138,N_6046);
nor U6377 (N_6377,N_6133,N_6121);
xor U6378 (N_6378,N_6089,N_6127);
or U6379 (N_6379,N_6199,N_6132);
or U6380 (N_6380,N_6157,N_6018);
nor U6381 (N_6381,N_6064,N_6129);
or U6382 (N_6382,N_6031,N_6036);
or U6383 (N_6383,N_6037,N_6099);
or U6384 (N_6384,N_6131,N_6071);
and U6385 (N_6385,N_6119,N_6082);
or U6386 (N_6386,N_6176,N_6166);
xor U6387 (N_6387,N_6091,N_6089);
xor U6388 (N_6388,N_6076,N_6182);
nor U6389 (N_6389,N_6157,N_6042);
or U6390 (N_6390,N_6090,N_6189);
nor U6391 (N_6391,N_6088,N_6082);
and U6392 (N_6392,N_6021,N_6125);
or U6393 (N_6393,N_6093,N_6144);
or U6394 (N_6394,N_6079,N_6115);
and U6395 (N_6395,N_6087,N_6036);
and U6396 (N_6396,N_6097,N_6193);
nand U6397 (N_6397,N_6195,N_6069);
or U6398 (N_6398,N_6013,N_6146);
nand U6399 (N_6399,N_6138,N_6023);
or U6400 (N_6400,N_6398,N_6384);
or U6401 (N_6401,N_6262,N_6229);
and U6402 (N_6402,N_6255,N_6336);
and U6403 (N_6403,N_6359,N_6298);
nor U6404 (N_6404,N_6273,N_6316);
and U6405 (N_6405,N_6259,N_6236);
and U6406 (N_6406,N_6373,N_6244);
or U6407 (N_6407,N_6221,N_6296);
and U6408 (N_6408,N_6237,N_6228);
nor U6409 (N_6409,N_6383,N_6242);
or U6410 (N_6410,N_6202,N_6210);
nand U6411 (N_6411,N_6230,N_6274);
nand U6412 (N_6412,N_6203,N_6223);
xor U6413 (N_6413,N_6265,N_6303);
and U6414 (N_6414,N_6397,N_6270);
nand U6415 (N_6415,N_6266,N_6337);
nand U6416 (N_6416,N_6363,N_6300);
or U6417 (N_6417,N_6287,N_6215);
xnor U6418 (N_6418,N_6299,N_6355);
or U6419 (N_6419,N_6284,N_6286);
and U6420 (N_6420,N_6331,N_6375);
or U6421 (N_6421,N_6365,N_6216);
nand U6422 (N_6422,N_6251,N_6217);
xor U6423 (N_6423,N_6332,N_6370);
and U6424 (N_6424,N_6322,N_6388);
nor U6425 (N_6425,N_6341,N_6311);
nand U6426 (N_6426,N_6234,N_6289);
or U6427 (N_6427,N_6288,N_6366);
nor U6428 (N_6428,N_6238,N_6334);
and U6429 (N_6429,N_6218,N_6256);
and U6430 (N_6430,N_6321,N_6302);
nand U6431 (N_6431,N_6310,N_6374);
and U6432 (N_6432,N_6247,N_6279);
or U6433 (N_6433,N_6282,N_6291);
and U6434 (N_6434,N_6313,N_6330);
nand U6435 (N_6435,N_6209,N_6305);
nor U6436 (N_6436,N_6350,N_6200);
or U6437 (N_6437,N_6390,N_6391);
or U6438 (N_6438,N_6250,N_6263);
or U6439 (N_6439,N_6357,N_6371);
nand U6440 (N_6440,N_6392,N_6278);
or U6441 (N_6441,N_6241,N_6243);
and U6442 (N_6442,N_6354,N_6314);
nor U6443 (N_6443,N_6283,N_6204);
nor U6444 (N_6444,N_6233,N_6208);
nor U6445 (N_6445,N_6301,N_6380);
or U6446 (N_6446,N_6294,N_6297);
or U6447 (N_6447,N_6222,N_6285);
nor U6448 (N_6448,N_6346,N_6214);
or U6449 (N_6449,N_6343,N_6220);
nand U6450 (N_6450,N_6349,N_6324);
and U6451 (N_6451,N_6269,N_6290);
nor U6452 (N_6452,N_6272,N_6264);
nor U6453 (N_6453,N_6377,N_6212);
and U6454 (N_6454,N_6226,N_6277);
nor U6455 (N_6455,N_6395,N_6225);
nand U6456 (N_6456,N_6258,N_6317);
nand U6457 (N_6457,N_6319,N_6352);
and U6458 (N_6458,N_6335,N_6245);
nor U6459 (N_6459,N_6368,N_6348);
xnor U6460 (N_6460,N_6268,N_6275);
nand U6461 (N_6461,N_6351,N_6280);
and U6462 (N_6462,N_6309,N_6304);
or U6463 (N_6463,N_6246,N_6249);
nor U6464 (N_6464,N_6323,N_6260);
nor U6465 (N_6465,N_6342,N_6292);
xor U6466 (N_6466,N_6367,N_6396);
nand U6467 (N_6467,N_6387,N_6338);
or U6468 (N_6468,N_6211,N_6207);
and U6469 (N_6469,N_6293,N_6358);
or U6470 (N_6470,N_6308,N_6276);
nand U6471 (N_6471,N_6267,N_6379);
or U6472 (N_6472,N_6320,N_6386);
nor U6473 (N_6473,N_6307,N_6385);
nor U6474 (N_6474,N_6306,N_6329);
xor U6475 (N_6475,N_6315,N_6382);
nor U6476 (N_6476,N_6253,N_6345);
nor U6477 (N_6477,N_6205,N_6360);
or U6478 (N_6478,N_6328,N_6394);
nand U6479 (N_6479,N_6356,N_6327);
nor U6480 (N_6480,N_6393,N_6364);
nor U6481 (N_6481,N_6206,N_6295);
nor U6482 (N_6482,N_6227,N_6252);
or U6483 (N_6483,N_6361,N_6344);
and U6484 (N_6484,N_6399,N_6239);
nor U6485 (N_6485,N_6254,N_6232);
or U6486 (N_6486,N_6333,N_6353);
xor U6487 (N_6487,N_6271,N_6312);
nor U6488 (N_6488,N_6248,N_6372);
and U6489 (N_6489,N_6213,N_6389);
nand U6490 (N_6490,N_6219,N_6378);
nor U6491 (N_6491,N_6339,N_6318);
nor U6492 (N_6492,N_6240,N_6257);
xnor U6493 (N_6493,N_6381,N_6281);
nor U6494 (N_6494,N_6231,N_6261);
and U6495 (N_6495,N_6369,N_6325);
and U6496 (N_6496,N_6376,N_6362);
or U6497 (N_6497,N_6201,N_6224);
or U6498 (N_6498,N_6347,N_6340);
and U6499 (N_6499,N_6326,N_6235);
xor U6500 (N_6500,N_6262,N_6365);
nand U6501 (N_6501,N_6388,N_6305);
or U6502 (N_6502,N_6226,N_6391);
nand U6503 (N_6503,N_6351,N_6232);
nor U6504 (N_6504,N_6219,N_6228);
and U6505 (N_6505,N_6272,N_6326);
nand U6506 (N_6506,N_6381,N_6220);
or U6507 (N_6507,N_6386,N_6390);
nand U6508 (N_6508,N_6278,N_6311);
and U6509 (N_6509,N_6307,N_6232);
or U6510 (N_6510,N_6335,N_6282);
nand U6511 (N_6511,N_6353,N_6248);
nand U6512 (N_6512,N_6253,N_6224);
or U6513 (N_6513,N_6388,N_6279);
xor U6514 (N_6514,N_6330,N_6232);
or U6515 (N_6515,N_6370,N_6338);
xnor U6516 (N_6516,N_6342,N_6270);
nand U6517 (N_6517,N_6201,N_6285);
nand U6518 (N_6518,N_6330,N_6307);
xor U6519 (N_6519,N_6343,N_6224);
or U6520 (N_6520,N_6259,N_6268);
or U6521 (N_6521,N_6271,N_6334);
xor U6522 (N_6522,N_6360,N_6327);
nor U6523 (N_6523,N_6277,N_6238);
and U6524 (N_6524,N_6380,N_6288);
or U6525 (N_6525,N_6272,N_6315);
nor U6526 (N_6526,N_6303,N_6255);
nand U6527 (N_6527,N_6229,N_6397);
nand U6528 (N_6528,N_6305,N_6244);
and U6529 (N_6529,N_6213,N_6351);
nor U6530 (N_6530,N_6253,N_6276);
nor U6531 (N_6531,N_6334,N_6382);
nor U6532 (N_6532,N_6384,N_6203);
and U6533 (N_6533,N_6278,N_6276);
and U6534 (N_6534,N_6308,N_6215);
nand U6535 (N_6535,N_6385,N_6251);
nor U6536 (N_6536,N_6203,N_6360);
and U6537 (N_6537,N_6344,N_6295);
and U6538 (N_6538,N_6370,N_6266);
xnor U6539 (N_6539,N_6294,N_6274);
xnor U6540 (N_6540,N_6382,N_6373);
and U6541 (N_6541,N_6384,N_6301);
and U6542 (N_6542,N_6373,N_6320);
nor U6543 (N_6543,N_6397,N_6204);
xnor U6544 (N_6544,N_6390,N_6296);
nor U6545 (N_6545,N_6242,N_6396);
and U6546 (N_6546,N_6327,N_6228);
or U6547 (N_6547,N_6280,N_6334);
or U6548 (N_6548,N_6363,N_6225);
nor U6549 (N_6549,N_6325,N_6280);
and U6550 (N_6550,N_6342,N_6334);
or U6551 (N_6551,N_6228,N_6380);
nand U6552 (N_6552,N_6320,N_6360);
or U6553 (N_6553,N_6353,N_6236);
and U6554 (N_6554,N_6290,N_6394);
and U6555 (N_6555,N_6209,N_6380);
xnor U6556 (N_6556,N_6324,N_6269);
xor U6557 (N_6557,N_6268,N_6306);
nor U6558 (N_6558,N_6201,N_6238);
or U6559 (N_6559,N_6212,N_6292);
xnor U6560 (N_6560,N_6236,N_6328);
nor U6561 (N_6561,N_6376,N_6208);
nor U6562 (N_6562,N_6225,N_6293);
nand U6563 (N_6563,N_6226,N_6323);
and U6564 (N_6564,N_6280,N_6392);
nor U6565 (N_6565,N_6316,N_6248);
nand U6566 (N_6566,N_6233,N_6313);
nand U6567 (N_6567,N_6238,N_6329);
xnor U6568 (N_6568,N_6340,N_6364);
or U6569 (N_6569,N_6330,N_6355);
nand U6570 (N_6570,N_6206,N_6300);
nor U6571 (N_6571,N_6330,N_6269);
or U6572 (N_6572,N_6349,N_6255);
nor U6573 (N_6573,N_6348,N_6300);
nor U6574 (N_6574,N_6333,N_6306);
nand U6575 (N_6575,N_6259,N_6272);
or U6576 (N_6576,N_6291,N_6284);
nand U6577 (N_6577,N_6282,N_6343);
nor U6578 (N_6578,N_6261,N_6296);
nor U6579 (N_6579,N_6320,N_6362);
xor U6580 (N_6580,N_6279,N_6241);
nor U6581 (N_6581,N_6279,N_6355);
xnor U6582 (N_6582,N_6396,N_6245);
or U6583 (N_6583,N_6284,N_6335);
and U6584 (N_6584,N_6302,N_6358);
nor U6585 (N_6585,N_6212,N_6227);
nand U6586 (N_6586,N_6271,N_6264);
or U6587 (N_6587,N_6364,N_6323);
or U6588 (N_6588,N_6222,N_6334);
nor U6589 (N_6589,N_6370,N_6368);
and U6590 (N_6590,N_6300,N_6296);
xor U6591 (N_6591,N_6333,N_6301);
xor U6592 (N_6592,N_6390,N_6239);
nor U6593 (N_6593,N_6206,N_6397);
xnor U6594 (N_6594,N_6286,N_6205);
nor U6595 (N_6595,N_6214,N_6222);
and U6596 (N_6596,N_6350,N_6275);
nor U6597 (N_6597,N_6209,N_6342);
nor U6598 (N_6598,N_6331,N_6295);
xor U6599 (N_6599,N_6356,N_6348);
and U6600 (N_6600,N_6573,N_6581);
and U6601 (N_6601,N_6475,N_6484);
or U6602 (N_6602,N_6522,N_6412);
or U6603 (N_6603,N_6564,N_6447);
or U6604 (N_6604,N_6508,N_6593);
nor U6605 (N_6605,N_6458,N_6529);
xnor U6606 (N_6606,N_6521,N_6494);
or U6607 (N_6607,N_6477,N_6424);
nor U6608 (N_6608,N_6551,N_6454);
or U6609 (N_6609,N_6496,N_6414);
nor U6610 (N_6610,N_6487,N_6462);
or U6611 (N_6611,N_6509,N_6434);
nor U6612 (N_6612,N_6489,N_6531);
and U6613 (N_6613,N_6548,N_6544);
or U6614 (N_6614,N_6427,N_6507);
or U6615 (N_6615,N_6570,N_6542);
or U6616 (N_6616,N_6530,N_6480);
and U6617 (N_6617,N_6552,N_6467);
or U6618 (N_6618,N_6580,N_6425);
nand U6619 (N_6619,N_6550,N_6422);
or U6620 (N_6620,N_6589,N_6441);
or U6621 (N_6621,N_6532,N_6557);
or U6622 (N_6622,N_6466,N_6463);
or U6623 (N_6623,N_6519,N_6599);
xor U6624 (N_6624,N_6429,N_6537);
nand U6625 (N_6625,N_6518,N_6418);
or U6626 (N_6626,N_6416,N_6415);
nor U6627 (N_6627,N_6421,N_6590);
or U6628 (N_6628,N_6493,N_6549);
and U6629 (N_6629,N_6520,N_6404);
nor U6630 (N_6630,N_6543,N_6411);
nand U6631 (N_6631,N_6406,N_6515);
and U6632 (N_6632,N_6474,N_6438);
and U6633 (N_6633,N_6553,N_6584);
nand U6634 (N_6634,N_6547,N_6565);
and U6635 (N_6635,N_6491,N_6476);
nand U6636 (N_6636,N_6478,N_6402);
or U6637 (N_6637,N_6569,N_6516);
nor U6638 (N_6638,N_6417,N_6588);
and U6639 (N_6639,N_6436,N_6513);
nor U6640 (N_6640,N_6448,N_6559);
nor U6641 (N_6641,N_6409,N_6413);
or U6642 (N_6642,N_6428,N_6598);
xor U6643 (N_6643,N_6437,N_6511);
nor U6644 (N_6644,N_6452,N_6453);
nor U6645 (N_6645,N_6596,N_6539);
nand U6646 (N_6646,N_6456,N_6533);
nor U6647 (N_6647,N_6574,N_6483);
nor U6648 (N_6648,N_6578,N_6464);
and U6649 (N_6649,N_6469,N_6432);
or U6650 (N_6650,N_6444,N_6535);
or U6651 (N_6651,N_6419,N_6545);
nand U6652 (N_6652,N_6426,N_6457);
nand U6653 (N_6653,N_6440,N_6488);
nand U6654 (N_6654,N_6512,N_6500);
nand U6655 (N_6655,N_6481,N_6492);
or U6656 (N_6656,N_6485,N_6517);
nor U6657 (N_6657,N_6470,N_6443);
nand U6658 (N_6658,N_6541,N_6465);
nor U6659 (N_6659,N_6451,N_6403);
or U6660 (N_6660,N_6439,N_6433);
and U6661 (N_6661,N_6410,N_6576);
nor U6662 (N_6662,N_6526,N_6423);
and U6663 (N_6663,N_6594,N_6446);
xor U6664 (N_6664,N_6435,N_6527);
and U6665 (N_6665,N_6442,N_6461);
and U6666 (N_6666,N_6568,N_6534);
or U6667 (N_6667,N_6571,N_6585);
nor U6668 (N_6668,N_6566,N_6592);
and U6669 (N_6669,N_6591,N_6554);
and U6670 (N_6670,N_6506,N_6504);
nor U6671 (N_6671,N_6471,N_6499);
nand U6672 (N_6672,N_6431,N_6503);
nand U6673 (N_6673,N_6586,N_6430);
and U6674 (N_6674,N_6495,N_6408);
or U6675 (N_6675,N_6567,N_6555);
or U6676 (N_6676,N_6405,N_6528);
or U6677 (N_6677,N_6577,N_6472);
nor U6678 (N_6678,N_6502,N_6460);
or U6679 (N_6679,N_6536,N_6546);
and U6680 (N_6680,N_6579,N_6563);
nand U6681 (N_6681,N_6525,N_6595);
or U6682 (N_6682,N_6514,N_6575);
nand U6683 (N_6683,N_6505,N_6498);
and U6684 (N_6684,N_6538,N_6473);
nand U6685 (N_6685,N_6510,N_6556);
xnor U6686 (N_6686,N_6468,N_6401);
nor U6687 (N_6687,N_6479,N_6482);
or U6688 (N_6688,N_6501,N_6486);
nor U6689 (N_6689,N_6455,N_6490);
nor U6690 (N_6690,N_6407,N_6524);
nor U6691 (N_6691,N_6582,N_6558);
nand U6692 (N_6692,N_6562,N_6572);
and U6693 (N_6693,N_6587,N_6540);
nand U6694 (N_6694,N_6459,N_6583);
xnor U6695 (N_6695,N_6449,N_6560);
nor U6696 (N_6696,N_6450,N_6445);
nand U6697 (N_6697,N_6400,N_6420);
nand U6698 (N_6698,N_6523,N_6597);
nor U6699 (N_6699,N_6561,N_6497);
nor U6700 (N_6700,N_6476,N_6478);
xor U6701 (N_6701,N_6479,N_6472);
xor U6702 (N_6702,N_6581,N_6542);
nor U6703 (N_6703,N_6444,N_6486);
nand U6704 (N_6704,N_6486,N_6579);
or U6705 (N_6705,N_6536,N_6586);
or U6706 (N_6706,N_6521,N_6463);
and U6707 (N_6707,N_6589,N_6529);
nand U6708 (N_6708,N_6548,N_6480);
or U6709 (N_6709,N_6453,N_6574);
nor U6710 (N_6710,N_6583,N_6534);
xnor U6711 (N_6711,N_6598,N_6491);
nand U6712 (N_6712,N_6521,N_6481);
xor U6713 (N_6713,N_6529,N_6582);
nand U6714 (N_6714,N_6513,N_6510);
or U6715 (N_6715,N_6554,N_6574);
or U6716 (N_6716,N_6458,N_6579);
or U6717 (N_6717,N_6545,N_6495);
or U6718 (N_6718,N_6547,N_6591);
nand U6719 (N_6719,N_6597,N_6496);
or U6720 (N_6720,N_6551,N_6593);
xnor U6721 (N_6721,N_6515,N_6442);
nand U6722 (N_6722,N_6518,N_6502);
nor U6723 (N_6723,N_6520,N_6581);
or U6724 (N_6724,N_6420,N_6518);
nor U6725 (N_6725,N_6405,N_6518);
nor U6726 (N_6726,N_6422,N_6545);
nor U6727 (N_6727,N_6567,N_6415);
xnor U6728 (N_6728,N_6531,N_6421);
nand U6729 (N_6729,N_6496,N_6591);
or U6730 (N_6730,N_6579,N_6406);
nand U6731 (N_6731,N_6574,N_6548);
nor U6732 (N_6732,N_6580,N_6598);
nor U6733 (N_6733,N_6516,N_6527);
xor U6734 (N_6734,N_6577,N_6550);
nand U6735 (N_6735,N_6541,N_6502);
and U6736 (N_6736,N_6531,N_6548);
nor U6737 (N_6737,N_6455,N_6452);
nor U6738 (N_6738,N_6423,N_6501);
nor U6739 (N_6739,N_6558,N_6417);
or U6740 (N_6740,N_6504,N_6480);
and U6741 (N_6741,N_6487,N_6463);
nor U6742 (N_6742,N_6496,N_6446);
or U6743 (N_6743,N_6562,N_6570);
nand U6744 (N_6744,N_6433,N_6409);
nor U6745 (N_6745,N_6539,N_6405);
and U6746 (N_6746,N_6549,N_6505);
and U6747 (N_6747,N_6435,N_6408);
nor U6748 (N_6748,N_6475,N_6561);
nand U6749 (N_6749,N_6521,N_6499);
and U6750 (N_6750,N_6453,N_6514);
or U6751 (N_6751,N_6410,N_6418);
nand U6752 (N_6752,N_6571,N_6410);
nand U6753 (N_6753,N_6490,N_6534);
nand U6754 (N_6754,N_6505,N_6575);
nand U6755 (N_6755,N_6563,N_6513);
and U6756 (N_6756,N_6415,N_6563);
or U6757 (N_6757,N_6485,N_6447);
and U6758 (N_6758,N_6540,N_6477);
or U6759 (N_6759,N_6440,N_6594);
and U6760 (N_6760,N_6521,N_6506);
nand U6761 (N_6761,N_6576,N_6540);
nor U6762 (N_6762,N_6587,N_6476);
and U6763 (N_6763,N_6451,N_6435);
and U6764 (N_6764,N_6580,N_6589);
and U6765 (N_6765,N_6486,N_6412);
or U6766 (N_6766,N_6532,N_6517);
nand U6767 (N_6767,N_6568,N_6524);
or U6768 (N_6768,N_6433,N_6451);
nand U6769 (N_6769,N_6507,N_6463);
nor U6770 (N_6770,N_6405,N_6511);
and U6771 (N_6771,N_6447,N_6522);
nor U6772 (N_6772,N_6436,N_6522);
xor U6773 (N_6773,N_6424,N_6439);
nand U6774 (N_6774,N_6494,N_6424);
and U6775 (N_6775,N_6562,N_6585);
or U6776 (N_6776,N_6401,N_6415);
nor U6777 (N_6777,N_6498,N_6530);
nor U6778 (N_6778,N_6459,N_6575);
and U6779 (N_6779,N_6422,N_6466);
or U6780 (N_6780,N_6491,N_6570);
nor U6781 (N_6781,N_6599,N_6557);
nor U6782 (N_6782,N_6512,N_6564);
and U6783 (N_6783,N_6518,N_6479);
or U6784 (N_6784,N_6560,N_6579);
nand U6785 (N_6785,N_6577,N_6449);
nand U6786 (N_6786,N_6560,N_6435);
and U6787 (N_6787,N_6575,N_6469);
nor U6788 (N_6788,N_6447,N_6519);
xor U6789 (N_6789,N_6547,N_6506);
or U6790 (N_6790,N_6440,N_6568);
or U6791 (N_6791,N_6519,N_6424);
and U6792 (N_6792,N_6599,N_6584);
nor U6793 (N_6793,N_6433,N_6580);
and U6794 (N_6794,N_6518,N_6430);
nor U6795 (N_6795,N_6466,N_6578);
or U6796 (N_6796,N_6524,N_6488);
nand U6797 (N_6797,N_6557,N_6562);
nand U6798 (N_6798,N_6490,N_6514);
and U6799 (N_6799,N_6560,N_6499);
nand U6800 (N_6800,N_6618,N_6738);
or U6801 (N_6801,N_6631,N_6679);
nor U6802 (N_6802,N_6633,N_6625);
nand U6803 (N_6803,N_6773,N_6605);
and U6804 (N_6804,N_6636,N_6656);
nor U6805 (N_6805,N_6739,N_6790);
and U6806 (N_6806,N_6639,N_6614);
nand U6807 (N_6807,N_6774,N_6740);
nor U6808 (N_6808,N_6711,N_6662);
and U6809 (N_6809,N_6748,N_6620);
nor U6810 (N_6810,N_6681,N_6690);
or U6811 (N_6811,N_6694,N_6772);
nor U6812 (N_6812,N_6665,N_6643);
xnor U6813 (N_6813,N_6783,N_6791);
nor U6814 (N_6814,N_6635,N_6743);
nand U6815 (N_6815,N_6661,N_6684);
or U6816 (N_6816,N_6727,N_6629);
nor U6817 (N_6817,N_6638,N_6601);
and U6818 (N_6818,N_6677,N_6664);
nand U6819 (N_6819,N_6715,N_6630);
nand U6820 (N_6820,N_6733,N_6615);
or U6821 (N_6821,N_6792,N_6749);
nand U6822 (N_6822,N_6680,N_6756);
and U6823 (N_6823,N_6660,N_6617);
nand U6824 (N_6824,N_6771,N_6759);
nand U6825 (N_6825,N_6746,N_6623);
and U6826 (N_6826,N_6688,N_6701);
xor U6827 (N_6827,N_6619,N_6788);
nand U6828 (N_6828,N_6722,N_6692);
and U6829 (N_6829,N_6725,N_6670);
nand U6830 (N_6830,N_6603,N_6699);
and U6831 (N_6831,N_6775,N_6626);
xnor U6832 (N_6832,N_6768,N_6611);
and U6833 (N_6833,N_6634,N_6781);
or U6834 (N_6834,N_6678,N_6627);
or U6835 (N_6835,N_6644,N_6785);
xnor U6836 (N_6836,N_6673,N_6794);
nand U6837 (N_6837,N_6776,N_6784);
or U6838 (N_6838,N_6793,N_6645);
xor U6839 (N_6839,N_6765,N_6700);
nor U6840 (N_6840,N_6745,N_6607);
and U6841 (N_6841,N_6649,N_6762);
nand U6842 (N_6842,N_6764,N_6609);
nand U6843 (N_6843,N_6786,N_6724);
nand U6844 (N_6844,N_6653,N_6663);
or U6845 (N_6845,N_6602,N_6695);
or U6846 (N_6846,N_6693,N_6697);
nand U6847 (N_6847,N_6742,N_6718);
and U6848 (N_6848,N_6797,N_6689);
or U6849 (N_6849,N_6728,N_6741);
and U6850 (N_6850,N_6709,N_6766);
nand U6851 (N_6851,N_6632,N_6683);
and U6852 (N_6852,N_6787,N_6622);
nor U6853 (N_6853,N_6696,N_6613);
nand U6854 (N_6854,N_6608,N_6606);
nor U6855 (N_6855,N_6778,N_6777);
and U6856 (N_6856,N_6737,N_6650);
or U6857 (N_6857,N_6779,N_6666);
and U6858 (N_6858,N_6652,N_6640);
nand U6859 (N_6859,N_6747,N_6676);
nand U6860 (N_6860,N_6682,N_6687);
nor U6861 (N_6861,N_6642,N_6647);
nor U6862 (N_6862,N_6760,N_6686);
or U6863 (N_6863,N_6717,N_6621);
nor U6864 (N_6864,N_6754,N_6753);
nand U6865 (N_6865,N_6735,N_6710);
nand U6866 (N_6866,N_6731,N_6769);
nand U6867 (N_6867,N_6674,N_6668);
nand U6868 (N_6868,N_6651,N_6761);
nand U6869 (N_6869,N_6705,N_6767);
and U6870 (N_6870,N_6707,N_6755);
nand U6871 (N_6871,N_6763,N_6714);
nor U6872 (N_6872,N_6780,N_6648);
nor U6873 (N_6873,N_6721,N_6655);
or U6874 (N_6874,N_6757,N_6719);
nand U6875 (N_6875,N_6770,N_6782);
and U6876 (N_6876,N_6704,N_6669);
nand U6877 (N_6877,N_6628,N_6600);
or U6878 (N_6878,N_6723,N_6716);
xnor U6879 (N_6879,N_6744,N_6657);
nor U6880 (N_6880,N_6604,N_6726);
nor U6881 (N_6881,N_6646,N_6685);
and U6882 (N_6882,N_6708,N_6616);
nor U6883 (N_6883,N_6667,N_6712);
and U6884 (N_6884,N_6671,N_6799);
and U6885 (N_6885,N_6672,N_6706);
or U6886 (N_6886,N_6654,N_6612);
nand U6887 (N_6887,N_6691,N_6610);
or U6888 (N_6888,N_6659,N_6795);
nand U6889 (N_6889,N_6641,N_6758);
or U6890 (N_6890,N_6736,N_6624);
nor U6891 (N_6891,N_6796,N_6730);
xnor U6892 (N_6892,N_6751,N_6798);
and U6893 (N_6893,N_6703,N_6720);
nand U6894 (N_6894,N_6637,N_6713);
xnor U6895 (N_6895,N_6752,N_6698);
xnor U6896 (N_6896,N_6702,N_6675);
or U6897 (N_6897,N_6789,N_6658);
and U6898 (N_6898,N_6750,N_6734);
nand U6899 (N_6899,N_6732,N_6729);
and U6900 (N_6900,N_6674,N_6704);
and U6901 (N_6901,N_6673,N_6725);
nand U6902 (N_6902,N_6750,N_6704);
or U6903 (N_6903,N_6695,N_6745);
nor U6904 (N_6904,N_6634,N_6707);
or U6905 (N_6905,N_6610,N_6651);
xnor U6906 (N_6906,N_6774,N_6692);
nand U6907 (N_6907,N_6642,N_6785);
or U6908 (N_6908,N_6778,N_6758);
or U6909 (N_6909,N_6784,N_6603);
and U6910 (N_6910,N_6651,N_6601);
nand U6911 (N_6911,N_6663,N_6629);
or U6912 (N_6912,N_6617,N_6756);
or U6913 (N_6913,N_6734,N_6621);
and U6914 (N_6914,N_6748,N_6621);
or U6915 (N_6915,N_6614,N_6708);
and U6916 (N_6916,N_6741,N_6665);
nor U6917 (N_6917,N_6661,N_6724);
or U6918 (N_6918,N_6642,N_6724);
nand U6919 (N_6919,N_6740,N_6656);
nor U6920 (N_6920,N_6611,N_6747);
or U6921 (N_6921,N_6711,N_6788);
or U6922 (N_6922,N_6790,N_6725);
nor U6923 (N_6923,N_6777,N_6799);
nor U6924 (N_6924,N_6723,N_6751);
nand U6925 (N_6925,N_6707,N_6744);
and U6926 (N_6926,N_6617,N_6667);
and U6927 (N_6927,N_6742,N_6746);
nor U6928 (N_6928,N_6679,N_6713);
nand U6929 (N_6929,N_6740,N_6683);
or U6930 (N_6930,N_6626,N_6697);
nand U6931 (N_6931,N_6609,N_6620);
nor U6932 (N_6932,N_6625,N_6724);
nor U6933 (N_6933,N_6783,N_6752);
and U6934 (N_6934,N_6687,N_6665);
or U6935 (N_6935,N_6753,N_6629);
and U6936 (N_6936,N_6699,N_6740);
nor U6937 (N_6937,N_6725,N_6694);
xor U6938 (N_6938,N_6653,N_6734);
nor U6939 (N_6939,N_6676,N_6765);
or U6940 (N_6940,N_6789,N_6691);
nand U6941 (N_6941,N_6783,N_6609);
or U6942 (N_6942,N_6705,N_6796);
or U6943 (N_6943,N_6622,N_6687);
xnor U6944 (N_6944,N_6632,N_6745);
or U6945 (N_6945,N_6750,N_6656);
or U6946 (N_6946,N_6733,N_6653);
nand U6947 (N_6947,N_6630,N_6776);
or U6948 (N_6948,N_6614,N_6684);
xnor U6949 (N_6949,N_6755,N_6788);
or U6950 (N_6950,N_6604,N_6725);
nor U6951 (N_6951,N_6792,N_6783);
nand U6952 (N_6952,N_6603,N_6760);
and U6953 (N_6953,N_6705,N_6682);
xor U6954 (N_6954,N_6779,N_6678);
xor U6955 (N_6955,N_6685,N_6731);
nand U6956 (N_6956,N_6763,N_6794);
xor U6957 (N_6957,N_6727,N_6683);
nand U6958 (N_6958,N_6629,N_6678);
nor U6959 (N_6959,N_6668,N_6614);
nand U6960 (N_6960,N_6667,N_6660);
nor U6961 (N_6961,N_6696,N_6738);
or U6962 (N_6962,N_6796,N_6697);
nor U6963 (N_6963,N_6602,N_6727);
or U6964 (N_6964,N_6669,N_6677);
or U6965 (N_6965,N_6621,N_6718);
nor U6966 (N_6966,N_6782,N_6619);
nor U6967 (N_6967,N_6767,N_6605);
and U6968 (N_6968,N_6648,N_6740);
nand U6969 (N_6969,N_6699,N_6674);
xnor U6970 (N_6970,N_6643,N_6604);
nor U6971 (N_6971,N_6755,N_6734);
nor U6972 (N_6972,N_6678,N_6780);
xnor U6973 (N_6973,N_6776,N_6600);
or U6974 (N_6974,N_6753,N_6718);
xor U6975 (N_6975,N_6733,N_6643);
or U6976 (N_6976,N_6636,N_6679);
nand U6977 (N_6977,N_6673,N_6736);
and U6978 (N_6978,N_6704,N_6717);
nand U6979 (N_6979,N_6652,N_6727);
or U6980 (N_6980,N_6658,N_6732);
xor U6981 (N_6981,N_6634,N_6778);
nand U6982 (N_6982,N_6795,N_6719);
or U6983 (N_6983,N_6737,N_6799);
nand U6984 (N_6984,N_6625,N_6688);
or U6985 (N_6985,N_6796,N_6714);
nor U6986 (N_6986,N_6644,N_6786);
xnor U6987 (N_6987,N_6744,N_6660);
or U6988 (N_6988,N_6753,N_6642);
and U6989 (N_6989,N_6622,N_6747);
nand U6990 (N_6990,N_6603,N_6798);
and U6991 (N_6991,N_6739,N_6664);
or U6992 (N_6992,N_6627,N_6744);
and U6993 (N_6993,N_6647,N_6634);
nand U6994 (N_6994,N_6766,N_6631);
nor U6995 (N_6995,N_6626,N_6663);
nand U6996 (N_6996,N_6792,N_6745);
or U6997 (N_6997,N_6686,N_6677);
or U6998 (N_6998,N_6656,N_6650);
nor U6999 (N_6999,N_6619,N_6757);
and U7000 (N_7000,N_6845,N_6866);
or U7001 (N_7001,N_6871,N_6832);
nor U7002 (N_7002,N_6925,N_6827);
nor U7003 (N_7003,N_6971,N_6933);
or U7004 (N_7004,N_6847,N_6964);
or U7005 (N_7005,N_6915,N_6970);
xor U7006 (N_7006,N_6893,N_6946);
and U7007 (N_7007,N_6816,N_6892);
or U7008 (N_7008,N_6987,N_6834);
nor U7009 (N_7009,N_6843,N_6813);
nand U7010 (N_7010,N_6858,N_6920);
or U7011 (N_7011,N_6846,N_6903);
nor U7012 (N_7012,N_6868,N_6801);
nand U7013 (N_7013,N_6914,N_6808);
and U7014 (N_7014,N_6839,N_6862);
nor U7015 (N_7015,N_6944,N_6902);
or U7016 (N_7016,N_6899,N_6997);
nor U7017 (N_7017,N_6835,N_6947);
nor U7018 (N_7018,N_6949,N_6958);
xor U7019 (N_7019,N_6821,N_6826);
nand U7020 (N_7020,N_6905,N_6950);
or U7021 (N_7021,N_6966,N_6981);
and U7022 (N_7022,N_6926,N_6955);
nand U7023 (N_7023,N_6838,N_6999);
xnor U7024 (N_7024,N_6810,N_6937);
nand U7025 (N_7025,N_6812,N_6895);
nand U7026 (N_7026,N_6954,N_6841);
nor U7027 (N_7027,N_6831,N_6890);
and U7028 (N_7028,N_6864,N_6819);
nor U7029 (N_7029,N_6972,N_6996);
nand U7030 (N_7030,N_6940,N_6900);
xnor U7031 (N_7031,N_6818,N_6945);
or U7032 (N_7032,N_6874,N_6990);
nor U7033 (N_7033,N_6849,N_6885);
xnor U7034 (N_7034,N_6921,N_6860);
nor U7035 (N_7035,N_6837,N_6924);
nor U7036 (N_7036,N_6941,N_6873);
nand U7037 (N_7037,N_6817,N_6928);
and U7038 (N_7038,N_6965,N_6979);
and U7039 (N_7039,N_6836,N_6894);
and U7040 (N_7040,N_6989,N_6901);
nand U7041 (N_7041,N_6891,N_6913);
nand U7042 (N_7042,N_6910,N_6992);
nor U7043 (N_7043,N_6815,N_6982);
or U7044 (N_7044,N_6842,N_6888);
or U7045 (N_7045,N_6939,N_6875);
xor U7046 (N_7046,N_6848,N_6806);
nand U7047 (N_7047,N_6850,N_6865);
or U7048 (N_7048,N_6911,N_6830);
xor U7049 (N_7049,N_6881,N_6896);
and U7050 (N_7050,N_6985,N_6986);
nor U7051 (N_7051,N_6867,N_6994);
nand U7052 (N_7052,N_6889,N_6930);
xnor U7053 (N_7053,N_6886,N_6825);
nand U7054 (N_7054,N_6983,N_6919);
nand U7055 (N_7055,N_6877,N_6828);
nor U7056 (N_7056,N_6880,N_6863);
nor U7057 (N_7057,N_6870,N_6988);
xnor U7058 (N_7058,N_6953,N_6974);
nor U7059 (N_7059,N_6978,N_6820);
nor U7060 (N_7060,N_6936,N_6922);
and U7061 (N_7061,N_6840,N_6887);
nand U7062 (N_7062,N_6991,N_6929);
nand U7063 (N_7063,N_6942,N_6811);
and U7064 (N_7064,N_6803,N_6968);
nor U7065 (N_7065,N_6822,N_6829);
nor U7066 (N_7066,N_6916,N_6918);
nand U7067 (N_7067,N_6973,N_6814);
nor U7068 (N_7068,N_6856,N_6906);
and U7069 (N_7069,N_6952,N_6963);
nor U7070 (N_7070,N_6809,N_6857);
or U7071 (N_7071,N_6927,N_6935);
nand U7072 (N_7072,N_6800,N_6853);
or U7073 (N_7073,N_6912,N_6934);
nor U7074 (N_7074,N_6969,N_6876);
and U7075 (N_7075,N_6908,N_6962);
and U7076 (N_7076,N_6923,N_6869);
and U7077 (N_7077,N_6823,N_6851);
and U7078 (N_7078,N_6956,N_6957);
nor U7079 (N_7079,N_6861,N_6976);
nor U7080 (N_7080,N_6961,N_6855);
or U7081 (N_7081,N_6938,N_6872);
and U7082 (N_7082,N_6993,N_6804);
xnor U7083 (N_7083,N_6833,N_6959);
xor U7084 (N_7084,N_6943,N_6951);
or U7085 (N_7085,N_6859,N_6805);
nand U7086 (N_7086,N_6931,N_6948);
or U7087 (N_7087,N_6967,N_6917);
xnor U7088 (N_7088,N_6909,N_6878);
nand U7089 (N_7089,N_6882,N_6824);
or U7090 (N_7090,N_6854,N_6995);
and U7091 (N_7091,N_6884,N_6998);
or U7092 (N_7092,N_6960,N_6898);
nand U7093 (N_7093,N_6852,N_6932);
nand U7094 (N_7094,N_6802,N_6844);
and U7095 (N_7095,N_6883,N_6897);
xor U7096 (N_7096,N_6907,N_6977);
nand U7097 (N_7097,N_6980,N_6984);
nor U7098 (N_7098,N_6904,N_6975);
and U7099 (N_7099,N_6807,N_6879);
nor U7100 (N_7100,N_6911,N_6901);
and U7101 (N_7101,N_6832,N_6957);
or U7102 (N_7102,N_6801,N_6855);
or U7103 (N_7103,N_6914,N_6900);
nand U7104 (N_7104,N_6867,N_6946);
nand U7105 (N_7105,N_6948,N_6861);
xnor U7106 (N_7106,N_6931,N_6824);
nor U7107 (N_7107,N_6941,N_6955);
nand U7108 (N_7108,N_6950,N_6993);
xnor U7109 (N_7109,N_6871,N_6841);
and U7110 (N_7110,N_6946,N_6858);
nor U7111 (N_7111,N_6953,N_6996);
nor U7112 (N_7112,N_6824,N_6977);
or U7113 (N_7113,N_6991,N_6965);
and U7114 (N_7114,N_6898,N_6938);
nand U7115 (N_7115,N_6990,N_6827);
or U7116 (N_7116,N_6909,N_6916);
and U7117 (N_7117,N_6915,N_6862);
or U7118 (N_7118,N_6939,N_6978);
nor U7119 (N_7119,N_6885,N_6883);
nor U7120 (N_7120,N_6816,N_6811);
or U7121 (N_7121,N_6975,N_6960);
and U7122 (N_7122,N_6908,N_6828);
and U7123 (N_7123,N_6953,N_6837);
or U7124 (N_7124,N_6864,N_6802);
nor U7125 (N_7125,N_6802,N_6843);
nor U7126 (N_7126,N_6822,N_6974);
nand U7127 (N_7127,N_6889,N_6907);
nand U7128 (N_7128,N_6906,N_6839);
nor U7129 (N_7129,N_6908,N_6834);
nor U7130 (N_7130,N_6922,N_6998);
nor U7131 (N_7131,N_6931,N_6894);
nand U7132 (N_7132,N_6876,N_6903);
or U7133 (N_7133,N_6820,N_6996);
nand U7134 (N_7134,N_6900,N_6847);
xnor U7135 (N_7135,N_6858,N_6930);
or U7136 (N_7136,N_6867,N_6940);
nand U7137 (N_7137,N_6819,N_6889);
nor U7138 (N_7138,N_6964,N_6949);
nand U7139 (N_7139,N_6812,N_6857);
xnor U7140 (N_7140,N_6805,N_6878);
nor U7141 (N_7141,N_6983,N_6897);
nand U7142 (N_7142,N_6895,N_6906);
or U7143 (N_7143,N_6816,N_6911);
and U7144 (N_7144,N_6834,N_6924);
nor U7145 (N_7145,N_6918,N_6928);
nand U7146 (N_7146,N_6908,N_6870);
or U7147 (N_7147,N_6819,N_6932);
or U7148 (N_7148,N_6818,N_6957);
nor U7149 (N_7149,N_6965,N_6974);
nand U7150 (N_7150,N_6914,N_6813);
or U7151 (N_7151,N_6862,N_6813);
xnor U7152 (N_7152,N_6940,N_6969);
nand U7153 (N_7153,N_6848,N_6835);
and U7154 (N_7154,N_6881,N_6910);
and U7155 (N_7155,N_6898,N_6888);
or U7156 (N_7156,N_6925,N_6834);
and U7157 (N_7157,N_6960,N_6971);
nand U7158 (N_7158,N_6816,N_6807);
nor U7159 (N_7159,N_6945,N_6927);
xor U7160 (N_7160,N_6914,N_6870);
and U7161 (N_7161,N_6849,N_6878);
or U7162 (N_7162,N_6921,N_6811);
nor U7163 (N_7163,N_6987,N_6986);
nor U7164 (N_7164,N_6867,N_6848);
or U7165 (N_7165,N_6830,N_6947);
nor U7166 (N_7166,N_6979,N_6868);
or U7167 (N_7167,N_6970,N_6842);
nor U7168 (N_7168,N_6941,N_6837);
nand U7169 (N_7169,N_6875,N_6853);
and U7170 (N_7170,N_6826,N_6902);
and U7171 (N_7171,N_6940,N_6873);
xnor U7172 (N_7172,N_6885,N_6827);
and U7173 (N_7173,N_6869,N_6987);
nor U7174 (N_7174,N_6981,N_6889);
nand U7175 (N_7175,N_6953,N_6809);
xor U7176 (N_7176,N_6866,N_6892);
and U7177 (N_7177,N_6860,N_6995);
nand U7178 (N_7178,N_6806,N_6958);
nor U7179 (N_7179,N_6979,N_6821);
nor U7180 (N_7180,N_6821,N_6804);
or U7181 (N_7181,N_6824,N_6829);
nand U7182 (N_7182,N_6857,N_6971);
or U7183 (N_7183,N_6831,N_6805);
nand U7184 (N_7184,N_6872,N_6926);
and U7185 (N_7185,N_6941,N_6894);
nand U7186 (N_7186,N_6844,N_6883);
and U7187 (N_7187,N_6911,N_6991);
nor U7188 (N_7188,N_6839,N_6985);
xnor U7189 (N_7189,N_6947,N_6831);
nor U7190 (N_7190,N_6815,N_6884);
and U7191 (N_7191,N_6804,N_6917);
nor U7192 (N_7192,N_6844,N_6850);
nor U7193 (N_7193,N_6818,N_6904);
nor U7194 (N_7194,N_6943,N_6872);
nor U7195 (N_7195,N_6822,N_6954);
xnor U7196 (N_7196,N_6945,N_6857);
nor U7197 (N_7197,N_6902,N_6908);
or U7198 (N_7198,N_6843,N_6986);
or U7199 (N_7199,N_6906,N_6962);
or U7200 (N_7200,N_7138,N_7102);
or U7201 (N_7201,N_7177,N_7027);
and U7202 (N_7202,N_7068,N_7124);
or U7203 (N_7203,N_7192,N_7196);
nor U7204 (N_7204,N_7149,N_7039);
nor U7205 (N_7205,N_7013,N_7088);
and U7206 (N_7206,N_7048,N_7037);
nand U7207 (N_7207,N_7029,N_7028);
and U7208 (N_7208,N_7105,N_7060);
nor U7209 (N_7209,N_7104,N_7100);
nor U7210 (N_7210,N_7030,N_7054);
nor U7211 (N_7211,N_7103,N_7141);
nor U7212 (N_7212,N_7148,N_7093);
and U7213 (N_7213,N_7059,N_7078);
nor U7214 (N_7214,N_7108,N_7136);
or U7215 (N_7215,N_7010,N_7167);
or U7216 (N_7216,N_7081,N_7131);
nand U7217 (N_7217,N_7058,N_7005);
xnor U7218 (N_7218,N_7125,N_7188);
xor U7219 (N_7219,N_7187,N_7014);
nand U7220 (N_7220,N_7157,N_7166);
nor U7221 (N_7221,N_7020,N_7174);
and U7222 (N_7222,N_7042,N_7052);
nor U7223 (N_7223,N_7116,N_7038);
and U7224 (N_7224,N_7023,N_7006);
and U7225 (N_7225,N_7050,N_7147);
nand U7226 (N_7226,N_7120,N_7034);
nor U7227 (N_7227,N_7067,N_7032);
or U7228 (N_7228,N_7071,N_7075);
nand U7229 (N_7229,N_7079,N_7072);
xor U7230 (N_7230,N_7156,N_7090);
and U7231 (N_7231,N_7087,N_7190);
nand U7232 (N_7232,N_7009,N_7171);
or U7233 (N_7233,N_7169,N_7119);
or U7234 (N_7234,N_7110,N_7094);
or U7235 (N_7235,N_7070,N_7160);
and U7236 (N_7236,N_7140,N_7083);
and U7237 (N_7237,N_7115,N_7063);
or U7238 (N_7238,N_7056,N_7164);
nand U7239 (N_7239,N_7184,N_7001);
nand U7240 (N_7240,N_7130,N_7176);
nor U7241 (N_7241,N_7109,N_7180);
or U7242 (N_7242,N_7175,N_7082);
nor U7243 (N_7243,N_7162,N_7051);
nor U7244 (N_7244,N_7183,N_7073);
and U7245 (N_7245,N_7182,N_7185);
and U7246 (N_7246,N_7133,N_7085);
nand U7247 (N_7247,N_7158,N_7002);
nand U7248 (N_7248,N_7007,N_7099);
nor U7249 (N_7249,N_7053,N_7043);
or U7250 (N_7250,N_7170,N_7172);
or U7251 (N_7251,N_7018,N_7076);
and U7252 (N_7252,N_7161,N_7064);
or U7253 (N_7253,N_7049,N_7061);
nor U7254 (N_7254,N_7163,N_7155);
nand U7255 (N_7255,N_7173,N_7146);
or U7256 (N_7256,N_7139,N_7055);
or U7257 (N_7257,N_7122,N_7040);
and U7258 (N_7258,N_7191,N_7019);
nor U7259 (N_7259,N_7069,N_7041);
and U7260 (N_7260,N_7086,N_7101);
and U7261 (N_7261,N_7021,N_7047);
nor U7262 (N_7262,N_7189,N_7017);
nand U7263 (N_7263,N_7107,N_7011);
nand U7264 (N_7264,N_7181,N_7153);
nor U7265 (N_7265,N_7199,N_7132);
xnor U7266 (N_7266,N_7062,N_7178);
nor U7267 (N_7267,N_7198,N_7126);
and U7268 (N_7268,N_7150,N_7168);
nand U7269 (N_7269,N_7144,N_7118);
or U7270 (N_7270,N_7065,N_7004);
xnor U7271 (N_7271,N_7151,N_7000);
or U7272 (N_7272,N_7096,N_7033);
nor U7273 (N_7273,N_7095,N_7145);
nor U7274 (N_7274,N_7128,N_7127);
and U7275 (N_7275,N_7026,N_7045);
and U7276 (N_7276,N_7117,N_7003);
nor U7277 (N_7277,N_7193,N_7135);
or U7278 (N_7278,N_7031,N_7022);
nand U7279 (N_7279,N_7091,N_7194);
nor U7280 (N_7280,N_7097,N_7092);
nand U7281 (N_7281,N_7121,N_7025);
or U7282 (N_7282,N_7008,N_7016);
and U7283 (N_7283,N_7142,N_7152);
xor U7284 (N_7284,N_7066,N_7012);
nor U7285 (N_7285,N_7112,N_7098);
nand U7286 (N_7286,N_7186,N_7123);
or U7287 (N_7287,N_7036,N_7024);
or U7288 (N_7288,N_7154,N_7080);
nor U7289 (N_7289,N_7084,N_7111);
nor U7290 (N_7290,N_7035,N_7114);
nor U7291 (N_7291,N_7195,N_7057);
nor U7292 (N_7292,N_7106,N_7077);
or U7293 (N_7293,N_7179,N_7015);
and U7294 (N_7294,N_7143,N_7089);
and U7295 (N_7295,N_7134,N_7046);
and U7296 (N_7296,N_7165,N_7197);
or U7297 (N_7297,N_7113,N_7137);
nor U7298 (N_7298,N_7044,N_7074);
and U7299 (N_7299,N_7129,N_7159);
or U7300 (N_7300,N_7161,N_7009);
nand U7301 (N_7301,N_7189,N_7116);
and U7302 (N_7302,N_7076,N_7172);
and U7303 (N_7303,N_7070,N_7034);
nand U7304 (N_7304,N_7131,N_7036);
or U7305 (N_7305,N_7123,N_7053);
nor U7306 (N_7306,N_7034,N_7144);
nor U7307 (N_7307,N_7026,N_7117);
or U7308 (N_7308,N_7039,N_7103);
nand U7309 (N_7309,N_7001,N_7183);
xnor U7310 (N_7310,N_7172,N_7181);
or U7311 (N_7311,N_7003,N_7052);
nor U7312 (N_7312,N_7034,N_7020);
xor U7313 (N_7313,N_7142,N_7020);
nand U7314 (N_7314,N_7155,N_7132);
or U7315 (N_7315,N_7172,N_7021);
or U7316 (N_7316,N_7132,N_7149);
nand U7317 (N_7317,N_7187,N_7058);
nand U7318 (N_7318,N_7084,N_7025);
and U7319 (N_7319,N_7128,N_7103);
nor U7320 (N_7320,N_7062,N_7093);
nand U7321 (N_7321,N_7182,N_7168);
nor U7322 (N_7322,N_7128,N_7156);
nand U7323 (N_7323,N_7054,N_7038);
or U7324 (N_7324,N_7089,N_7148);
nor U7325 (N_7325,N_7051,N_7007);
xnor U7326 (N_7326,N_7120,N_7083);
nor U7327 (N_7327,N_7158,N_7048);
or U7328 (N_7328,N_7122,N_7052);
and U7329 (N_7329,N_7082,N_7129);
xor U7330 (N_7330,N_7014,N_7126);
or U7331 (N_7331,N_7065,N_7178);
and U7332 (N_7332,N_7005,N_7036);
and U7333 (N_7333,N_7095,N_7049);
nor U7334 (N_7334,N_7041,N_7110);
xnor U7335 (N_7335,N_7059,N_7105);
and U7336 (N_7336,N_7189,N_7042);
nor U7337 (N_7337,N_7123,N_7076);
and U7338 (N_7338,N_7036,N_7038);
or U7339 (N_7339,N_7106,N_7027);
and U7340 (N_7340,N_7152,N_7078);
nor U7341 (N_7341,N_7067,N_7117);
and U7342 (N_7342,N_7053,N_7184);
nand U7343 (N_7343,N_7104,N_7132);
or U7344 (N_7344,N_7034,N_7164);
nand U7345 (N_7345,N_7004,N_7030);
and U7346 (N_7346,N_7103,N_7082);
nor U7347 (N_7347,N_7142,N_7139);
nor U7348 (N_7348,N_7050,N_7079);
or U7349 (N_7349,N_7181,N_7050);
nor U7350 (N_7350,N_7026,N_7030);
nand U7351 (N_7351,N_7029,N_7024);
or U7352 (N_7352,N_7093,N_7130);
or U7353 (N_7353,N_7167,N_7099);
nand U7354 (N_7354,N_7118,N_7030);
nor U7355 (N_7355,N_7027,N_7172);
nand U7356 (N_7356,N_7038,N_7195);
nand U7357 (N_7357,N_7084,N_7162);
and U7358 (N_7358,N_7193,N_7108);
nand U7359 (N_7359,N_7097,N_7042);
or U7360 (N_7360,N_7038,N_7132);
or U7361 (N_7361,N_7168,N_7100);
and U7362 (N_7362,N_7094,N_7134);
nor U7363 (N_7363,N_7052,N_7031);
xor U7364 (N_7364,N_7140,N_7067);
and U7365 (N_7365,N_7101,N_7030);
or U7366 (N_7366,N_7177,N_7019);
nand U7367 (N_7367,N_7194,N_7060);
nor U7368 (N_7368,N_7056,N_7199);
and U7369 (N_7369,N_7006,N_7109);
or U7370 (N_7370,N_7082,N_7011);
xnor U7371 (N_7371,N_7054,N_7095);
or U7372 (N_7372,N_7176,N_7013);
nor U7373 (N_7373,N_7187,N_7138);
xnor U7374 (N_7374,N_7174,N_7166);
nand U7375 (N_7375,N_7080,N_7170);
nand U7376 (N_7376,N_7018,N_7014);
or U7377 (N_7377,N_7135,N_7183);
and U7378 (N_7378,N_7178,N_7177);
nor U7379 (N_7379,N_7007,N_7147);
and U7380 (N_7380,N_7102,N_7141);
nor U7381 (N_7381,N_7051,N_7192);
nand U7382 (N_7382,N_7062,N_7120);
nor U7383 (N_7383,N_7056,N_7010);
nor U7384 (N_7384,N_7026,N_7084);
and U7385 (N_7385,N_7087,N_7076);
nand U7386 (N_7386,N_7052,N_7140);
and U7387 (N_7387,N_7057,N_7090);
nor U7388 (N_7388,N_7074,N_7184);
nand U7389 (N_7389,N_7191,N_7108);
or U7390 (N_7390,N_7135,N_7196);
nor U7391 (N_7391,N_7017,N_7176);
nor U7392 (N_7392,N_7170,N_7114);
nand U7393 (N_7393,N_7150,N_7070);
nor U7394 (N_7394,N_7051,N_7084);
nor U7395 (N_7395,N_7084,N_7053);
and U7396 (N_7396,N_7184,N_7157);
nand U7397 (N_7397,N_7062,N_7066);
nand U7398 (N_7398,N_7053,N_7044);
or U7399 (N_7399,N_7100,N_7072);
nor U7400 (N_7400,N_7275,N_7340);
or U7401 (N_7401,N_7355,N_7298);
nor U7402 (N_7402,N_7364,N_7286);
nor U7403 (N_7403,N_7390,N_7331);
and U7404 (N_7404,N_7247,N_7282);
nand U7405 (N_7405,N_7241,N_7376);
nor U7406 (N_7406,N_7329,N_7213);
and U7407 (N_7407,N_7326,N_7293);
and U7408 (N_7408,N_7334,N_7348);
nor U7409 (N_7409,N_7232,N_7264);
or U7410 (N_7410,N_7330,N_7276);
nor U7411 (N_7411,N_7283,N_7371);
nand U7412 (N_7412,N_7302,N_7208);
nand U7413 (N_7413,N_7354,N_7342);
or U7414 (N_7414,N_7352,N_7291);
and U7415 (N_7415,N_7290,N_7363);
or U7416 (N_7416,N_7273,N_7328);
nor U7417 (N_7417,N_7219,N_7216);
xor U7418 (N_7418,N_7357,N_7211);
or U7419 (N_7419,N_7381,N_7396);
nand U7420 (N_7420,N_7385,N_7256);
nand U7421 (N_7421,N_7315,N_7224);
or U7422 (N_7422,N_7307,N_7395);
xor U7423 (N_7423,N_7246,N_7312);
nor U7424 (N_7424,N_7345,N_7372);
or U7425 (N_7425,N_7323,N_7252);
and U7426 (N_7426,N_7305,N_7332);
nand U7427 (N_7427,N_7397,N_7251);
nor U7428 (N_7428,N_7316,N_7274);
and U7429 (N_7429,N_7382,N_7226);
and U7430 (N_7430,N_7341,N_7319);
or U7431 (N_7431,N_7386,N_7253);
nor U7432 (N_7432,N_7394,N_7349);
xnor U7433 (N_7433,N_7221,N_7205);
or U7434 (N_7434,N_7248,N_7212);
nor U7435 (N_7435,N_7258,N_7344);
nor U7436 (N_7436,N_7222,N_7347);
nor U7437 (N_7437,N_7346,N_7321);
nand U7438 (N_7438,N_7288,N_7284);
nand U7439 (N_7439,N_7369,N_7367);
and U7440 (N_7440,N_7242,N_7384);
nand U7441 (N_7441,N_7304,N_7261);
nor U7442 (N_7442,N_7306,N_7398);
nor U7443 (N_7443,N_7351,N_7327);
and U7444 (N_7444,N_7237,N_7230);
nor U7445 (N_7445,N_7285,N_7217);
nand U7446 (N_7446,N_7207,N_7260);
or U7447 (N_7447,N_7227,N_7308);
nand U7448 (N_7448,N_7380,N_7203);
or U7449 (N_7449,N_7214,N_7263);
and U7450 (N_7450,N_7249,N_7268);
and U7451 (N_7451,N_7265,N_7383);
xor U7452 (N_7452,N_7377,N_7210);
nor U7453 (N_7453,N_7292,N_7368);
and U7454 (N_7454,N_7374,N_7389);
or U7455 (N_7455,N_7324,N_7281);
nor U7456 (N_7456,N_7399,N_7365);
and U7457 (N_7457,N_7257,N_7297);
nand U7458 (N_7458,N_7336,N_7300);
nor U7459 (N_7459,N_7322,N_7361);
and U7460 (N_7460,N_7279,N_7343);
or U7461 (N_7461,N_7223,N_7201);
and U7462 (N_7462,N_7392,N_7234);
nand U7463 (N_7463,N_7356,N_7235);
or U7464 (N_7464,N_7303,N_7313);
nor U7465 (N_7465,N_7267,N_7339);
nand U7466 (N_7466,N_7206,N_7280);
or U7467 (N_7467,N_7295,N_7259);
and U7468 (N_7468,N_7337,N_7362);
or U7469 (N_7469,N_7320,N_7220);
and U7470 (N_7470,N_7335,N_7271);
nor U7471 (N_7471,N_7360,N_7350);
nor U7472 (N_7472,N_7272,N_7294);
and U7473 (N_7473,N_7243,N_7236);
nor U7474 (N_7474,N_7228,N_7209);
nor U7475 (N_7475,N_7296,N_7317);
nand U7476 (N_7476,N_7366,N_7388);
nor U7477 (N_7477,N_7318,N_7314);
nor U7478 (N_7478,N_7287,N_7373);
or U7479 (N_7479,N_7289,N_7278);
nor U7480 (N_7480,N_7378,N_7301);
xor U7481 (N_7481,N_7309,N_7393);
nor U7482 (N_7482,N_7333,N_7218);
and U7483 (N_7483,N_7299,N_7277);
nand U7484 (N_7484,N_7266,N_7375);
xnor U7485 (N_7485,N_7204,N_7269);
nor U7486 (N_7486,N_7387,N_7200);
nor U7487 (N_7487,N_7202,N_7338);
or U7488 (N_7488,N_7229,N_7353);
or U7489 (N_7489,N_7391,N_7240);
nand U7490 (N_7490,N_7379,N_7238);
xnor U7491 (N_7491,N_7215,N_7231);
nor U7492 (N_7492,N_7255,N_7370);
and U7493 (N_7493,N_7325,N_7359);
and U7494 (N_7494,N_7244,N_7358);
and U7495 (N_7495,N_7245,N_7233);
nor U7496 (N_7496,N_7311,N_7239);
and U7497 (N_7497,N_7250,N_7225);
or U7498 (N_7498,N_7310,N_7262);
xor U7499 (N_7499,N_7254,N_7270);
xnor U7500 (N_7500,N_7215,N_7375);
nand U7501 (N_7501,N_7203,N_7315);
and U7502 (N_7502,N_7309,N_7367);
xor U7503 (N_7503,N_7366,N_7275);
nand U7504 (N_7504,N_7318,N_7289);
xnor U7505 (N_7505,N_7311,N_7351);
nor U7506 (N_7506,N_7247,N_7270);
and U7507 (N_7507,N_7208,N_7354);
xor U7508 (N_7508,N_7244,N_7256);
nor U7509 (N_7509,N_7307,N_7393);
nor U7510 (N_7510,N_7368,N_7229);
and U7511 (N_7511,N_7343,N_7376);
and U7512 (N_7512,N_7238,N_7218);
or U7513 (N_7513,N_7270,N_7206);
or U7514 (N_7514,N_7355,N_7241);
and U7515 (N_7515,N_7375,N_7307);
or U7516 (N_7516,N_7278,N_7286);
or U7517 (N_7517,N_7394,N_7206);
nor U7518 (N_7518,N_7340,N_7288);
nor U7519 (N_7519,N_7263,N_7381);
and U7520 (N_7520,N_7378,N_7288);
nand U7521 (N_7521,N_7328,N_7387);
nand U7522 (N_7522,N_7335,N_7266);
or U7523 (N_7523,N_7208,N_7372);
and U7524 (N_7524,N_7397,N_7300);
nand U7525 (N_7525,N_7389,N_7264);
nor U7526 (N_7526,N_7319,N_7340);
nand U7527 (N_7527,N_7222,N_7251);
nand U7528 (N_7528,N_7219,N_7248);
nor U7529 (N_7529,N_7226,N_7350);
nor U7530 (N_7530,N_7238,N_7205);
nor U7531 (N_7531,N_7214,N_7239);
nor U7532 (N_7532,N_7313,N_7205);
nand U7533 (N_7533,N_7223,N_7292);
or U7534 (N_7534,N_7338,N_7291);
or U7535 (N_7535,N_7394,N_7376);
or U7536 (N_7536,N_7284,N_7382);
nand U7537 (N_7537,N_7330,N_7228);
and U7538 (N_7538,N_7374,N_7283);
nor U7539 (N_7539,N_7350,N_7323);
and U7540 (N_7540,N_7287,N_7225);
xor U7541 (N_7541,N_7320,N_7392);
xnor U7542 (N_7542,N_7353,N_7366);
xor U7543 (N_7543,N_7301,N_7368);
xor U7544 (N_7544,N_7365,N_7283);
nand U7545 (N_7545,N_7201,N_7316);
nor U7546 (N_7546,N_7322,N_7364);
xnor U7547 (N_7547,N_7231,N_7358);
or U7548 (N_7548,N_7348,N_7382);
nor U7549 (N_7549,N_7264,N_7278);
or U7550 (N_7550,N_7211,N_7255);
or U7551 (N_7551,N_7273,N_7359);
or U7552 (N_7552,N_7238,N_7369);
nand U7553 (N_7553,N_7304,N_7342);
nor U7554 (N_7554,N_7308,N_7393);
and U7555 (N_7555,N_7386,N_7320);
or U7556 (N_7556,N_7290,N_7268);
nand U7557 (N_7557,N_7293,N_7380);
or U7558 (N_7558,N_7323,N_7352);
and U7559 (N_7559,N_7267,N_7212);
nor U7560 (N_7560,N_7348,N_7239);
or U7561 (N_7561,N_7228,N_7202);
xor U7562 (N_7562,N_7217,N_7286);
nor U7563 (N_7563,N_7341,N_7240);
or U7564 (N_7564,N_7256,N_7381);
nor U7565 (N_7565,N_7220,N_7370);
xnor U7566 (N_7566,N_7318,N_7216);
and U7567 (N_7567,N_7231,N_7236);
and U7568 (N_7568,N_7274,N_7219);
nor U7569 (N_7569,N_7222,N_7358);
nand U7570 (N_7570,N_7250,N_7359);
or U7571 (N_7571,N_7264,N_7215);
nor U7572 (N_7572,N_7203,N_7351);
nand U7573 (N_7573,N_7345,N_7257);
and U7574 (N_7574,N_7295,N_7232);
or U7575 (N_7575,N_7241,N_7288);
or U7576 (N_7576,N_7278,N_7239);
nor U7577 (N_7577,N_7336,N_7353);
and U7578 (N_7578,N_7217,N_7203);
and U7579 (N_7579,N_7378,N_7214);
or U7580 (N_7580,N_7295,N_7323);
or U7581 (N_7581,N_7278,N_7367);
and U7582 (N_7582,N_7315,N_7391);
nand U7583 (N_7583,N_7365,N_7379);
or U7584 (N_7584,N_7284,N_7299);
or U7585 (N_7585,N_7285,N_7341);
or U7586 (N_7586,N_7244,N_7210);
nand U7587 (N_7587,N_7235,N_7275);
xor U7588 (N_7588,N_7369,N_7276);
nor U7589 (N_7589,N_7359,N_7339);
and U7590 (N_7590,N_7373,N_7268);
nor U7591 (N_7591,N_7261,N_7315);
nand U7592 (N_7592,N_7393,N_7322);
and U7593 (N_7593,N_7267,N_7391);
nand U7594 (N_7594,N_7330,N_7333);
xnor U7595 (N_7595,N_7266,N_7332);
nand U7596 (N_7596,N_7200,N_7365);
xnor U7597 (N_7597,N_7393,N_7320);
or U7598 (N_7598,N_7297,N_7282);
or U7599 (N_7599,N_7265,N_7357);
nor U7600 (N_7600,N_7597,N_7547);
or U7601 (N_7601,N_7550,N_7429);
or U7602 (N_7602,N_7572,N_7596);
nand U7603 (N_7603,N_7495,N_7434);
xnor U7604 (N_7604,N_7585,N_7408);
or U7605 (N_7605,N_7482,N_7439);
nand U7606 (N_7606,N_7407,N_7502);
or U7607 (N_7607,N_7558,N_7406);
nor U7608 (N_7608,N_7409,N_7538);
nor U7609 (N_7609,N_7404,N_7450);
or U7610 (N_7610,N_7489,N_7445);
and U7611 (N_7611,N_7480,N_7527);
and U7612 (N_7612,N_7470,N_7432);
xnor U7613 (N_7613,N_7496,N_7462);
or U7614 (N_7614,N_7467,N_7461);
nor U7615 (N_7615,N_7566,N_7548);
or U7616 (N_7616,N_7457,N_7587);
xnor U7617 (N_7617,N_7512,N_7567);
or U7618 (N_7618,N_7528,N_7400);
nor U7619 (N_7619,N_7431,N_7544);
and U7620 (N_7620,N_7413,N_7551);
nor U7621 (N_7621,N_7446,N_7412);
or U7622 (N_7622,N_7532,N_7458);
nor U7623 (N_7623,N_7580,N_7594);
and U7624 (N_7624,N_7485,N_7456);
and U7625 (N_7625,N_7592,N_7589);
nor U7626 (N_7626,N_7483,N_7490);
and U7627 (N_7627,N_7443,N_7599);
nor U7628 (N_7628,N_7510,N_7455);
xnor U7629 (N_7629,N_7565,N_7542);
nand U7630 (N_7630,N_7537,N_7442);
or U7631 (N_7631,N_7477,N_7531);
nor U7632 (N_7632,N_7522,N_7486);
nor U7633 (N_7633,N_7546,N_7511);
nor U7634 (N_7634,N_7424,N_7557);
and U7635 (N_7635,N_7509,N_7451);
and U7636 (N_7636,N_7453,N_7523);
nor U7637 (N_7637,N_7574,N_7520);
and U7638 (N_7638,N_7459,N_7568);
nor U7639 (N_7639,N_7578,N_7479);
nand U7640 (N_7640,N_7518,N_7500);
and U7641 (N_7641,N_7469,N_7478);
and U7642 (N_7642,N_7493,N_7414);
and U7643 (N_7643,N_7519,N_7582);
and U7644 (N_7644,N_7463,N_7472);
or U7645 (N_7645,N_7573,N_7583);
and U7646 (N_7646,N_7498,N_7579);
or U7647 (N_7647,N_7436,N_7541);
and U7648 (N_7648,N_7590,N_7586);
nor U7649 (N_7649,N_7452,N_7494);
nand U7650 (N_7650,N_7475,N_7556);
and U7651 (N_7651,N_7517,N_7464);
and U7652 (N_7652,N_7561,N_7421);
and U7653 (N_7653,N_7552,N_7549);
nor U7654 (N_7654,N_7543,N_7491);
and U7655 (N_7655,N_7402,N_7417);
nand U7656 (N_7656,N_7405,N_7437);
nor U7657 (N_7657,N_7427,N_7591);
nor U7658 (N_7658,N_7575,N_7540);
or U7659 (N_7659,N_7473,N_7569);
nand U7660 (N_7660,N_7466,N_7422);
and U7661 (N_7661,N_7492,N_7416);
or U7662 (N_7662,N_7420,N_7499);
or U7663 (N_7663,N_7539,N_7508);
nor U7664 (N_7664,N_7529,N_7468);
nor U7665 (N_7665,N_7449,N_7530);
nor U7666 (N_7666,N_7545,N_7430);
nor U7667 (N_7667,N_7465,N_7415);
nand U7668 (N_7668,N_7438,N_7513);
nor U7669 (N_7669,N_7503,N_7576);
and U7670 (N_7670,N_7411,N_7448);
nor U7671 (N_7671,N_7571,N_7553);
nor U7672 (N_7672,N_7515,N_7555);
and U7673 (N_7673,N_7506,N_7526);
and U7674 (N_7674,N_7559,N_7564);
or U7675 (N_7675,N_7441,N_7504);
nand U7676 (N_7676,N_7460,N_7454);
xnor U7677 (N_7677,N_7584,N_7435);
and U7678 (N_7678,N_7440,N_7554);
and U7679 (N_7679,N_7433,N_7524);
nand U7680 (N_7680,N_7521,N_7501);
nand U7681 (N_7681,N_7581,N_7401);
nand U7682 (N_7682,N_7418,N_7444);
nand U7683 (N_7683,N_7593,N_7533);
nand U7684 (N_7684,N_7598,N_7425);
and U7685 (N_7685,N_7588,N_7423);
nand U7686 (N_7686,N_7505,N_7562);
nor U7687 (N_7687,N_7474,N_7403);
nor U7688 (N_7688,N_7560,N_7426);
nand U7689 (N_7689,N_7536,N_7525);
nor U7690 (N_7690,N_7488,N_7476);
or U7691 (N_7691,N_7481,N_7507);
nand U7692 (N_7692,N_7563,N_7484);
or U7693 (N_7693,N_7516,N_7497);
and U7694 (N_7694,N_7535,N_7428);
nor U7695 (N_7695,N_7487,N_7410);
and U7696 (N_7696,N_7534,N_7570);
or U7697 (N_7697,N_7447,N_7577);
nor U7698 (N_7698,N_7514,N_7419);
nor U7699 (N_7699,N_7595,N_7471);
nor U7700 (N_7700,N_7536,N_7412);
nand U7701 (N_7701,N_7402,N_7507);
nand U7702 (N_7702,N_7466,N_7413);
nand U7703 (N_7703,N_7551,N_7590);
nor U7704 (N_7704,N_7535,N_7475);
xor U7705 (N_7705,N_7579,N_7455);
xnor U7706 (N_7706,N_7570,N_7499);
and U7707 (N_7707,N_7557,N_7540);
nor U7708 (N_7708,N_7555,N_7411);
nor U7709 (N_7709,N_7416,N_7463);
nor U7710 (N_7710,N_7481,N_7490);
nand U7711 (N_7711,N_7546,N_7528);
nand U7712 (N_7712,N_7402,N_7483);
and U7713 (N_7713,N_7421,N_7450);
and U7714 (N_7714,N_7416,N_7474);
nor U7715 (N_7715,N_7498,N_7591);
and U7716 (N_7716,N_7492,N_7423);
or U7717 (N_7717,N_7587,N_7468);
or U7718 (N_7718,N_7415,N_7567);
and U7719 (N_7719,N_7553,N_7513);
nor U7720 (N_7720,N_7479,N_7492);
xor U7721 (N_7721,N_7521,N_7440);
or U7722 (N_7722,N_7531,N_7520);
nand U7723 (N_7723,N_7454,N_7439);
nor U7724 (N_7724,N_7536,N_7492);
or U7725 (N_7725,N_7587,N_7552);
and U7726 (N_7726,N_7475,N_7574);
and U7727 (N_7727,N_7585,N_7477);
nand U7728 (N_7728,N_7507,N_7486);
nor U7729 (N_7729,N_7488,N_7522);
nor U7730 (N_7730,N_7573,N_7465);
nor U7731 (N_7731,N_7472,N_7460);
nand U7732 (N_7732,N_7506,N_7403);
nand U7733 (N_7733,N_7455,N_7533);
or U7734 (N_7734,N_7592,N_7570);
xnor U7735 (N_7735,N_7502,N_7557);
nand U7736 (N_7736,N_7508,N_7483);
or U7737 (N_7737,N_7503,N_7513);
nor U7738 (N_7738,N_7549,N_7474);
nand U7739 (N_7739,N_7515,N_7450);
nor U7740 (N_7740,N_7465,N_7450);
and U7741 (N_7741,N_7556,N_7570);
nor U7742 (N_7742,N_7448,N_7401);
or U7743 (N_7743,N_7583,N_7489);
and U7744 (N_7744,N_7459,N_7555);
and U7745 (N_7745,N_7535,N_7494);
nor U7746 (N_7746,N_7538,N_7485);
nand U7747 (N_7747,N_7537,N_7514);
nor U7748 (N_7748,N_7423,N_7518);
and U7749 (N_7749,N_7473,N_7503);
or U7750 (N_7750,N_7548,N_7483);
and U7751 (N_7751,N_7515,N_7475);
nor U7752 (N_7752,N_7562,N_7523);
or U7753 (N_7753,N_7455,N_7401);
and U7754 (N_7754,N_7506,N_7585);
or U7755 (N_7755,N_7487,N_7536);
nor U7756 (N_7756,N_7509,N_7500);
and U7757 (N_7757,N_7494,N_7428);
and U7758 (N_7758,N_7598,N_7477);
nand U7759 (N_7759,N_7427,N_7423);
or U7760 (N_7760,N_7535,N_7438);
nor U7761 (N_7761,N_7460,N_7440);
nor U7762 (N_7762,N_7447,N_7590);
nor U7763 (N_7763,N_7454,N_7402);
nor U7764 (N_7764,N_7596,N_7442);
nor U7765 (N_7765,N_7560,N_7472);
nand U7766 (N_7766,N_7509,N_7589);
and U7767 (N_7767,N_7453,N_7586);
or U7768 (N_7768,N_7406,N_7559);
nand U7769 (N_7769,N_7431,N_7568);
xor U7770 (N_7770,N_7491,N_7530);
or U7771 (N_7771,N_7475,N_7441);
nor U7772 (N_7772,N_7599,N_7471);
nand U7773 (N_7773,N_7460,N_7480);
nor U7774 (N_7774,N_7415,N_7426);
or U7775 (N_7775,N_7436,N_7475);
nand U7776 (N_7776,N_7464,N_7467);
or U7777 (N_7777,N_7597,N_7457);
or U7778 (N_7778,N_7531,N_7555);
or U7779 (N_7779,N_7473,N_7507);
and U7780 (N_7780,N_7579,N_7488);
nor U7781 (N_7781,N_7555,N_7516);
nor U7782 (N_7782,N_7571,N_7597);
and U7783 (N_7783,N_7458,N_7467);
xnor U7784 (N_7784,N_7513,N_7442);
or U7785 (N_7785,N_7505,N_7417);
and U7786 (N_7786,N_7480,N_7495);
xor U7787 (N_7787,N_7589,N_7586);
xnor U7788 (N_7788,N_7400,N_7515);
nor U7789 (N_7789,N_7495,N_7411);
and U7790 (N_7790,N_7577,N_7496);
nand U7791 (N_7791,N_7403,N_7565);
xnor U7792 (N_7792,N_7449,N_7564);
nor U7793 (N_7793,N_7429,N_7467);
or U7794 (N_7794,N_7540,N_7453);
and U7795 (N_7795,N_7552,N_7472);
and U7796 (N_7796,N_7568,N_7503);
nand U7797 (N_7797,N_7443,N_7548);
or U7798 (N_7798,N_7463,N_7567);
and U7799 (N_7799,N_7540,N_7433);
or U7800 (N_7800,N_7795,N_7742);
nand U7801 (N_7801,N_7613,N_7713);
and U7802 (N_7802,N_7749,N_7685);
and U7803 (N_7803,N_7793,N_7763);
nor U7804 (N_7804,N_7669,N_7661);
nor U7805 (N_7805,N_7721,N_7640);
and U7806 (N_7806,N_7738,N_7643);
nand U7807 (N_7807,N_7706,N_7603);
nand U7808 (N_7808,N_7744,N_7671);
nand U7809 (N_7809,N_7644,N_7797);
and U7810 (N_7810,N_7759,N_7645);
and U7811 (N_7811,N_7715,N_7748);
nor U7812 (N_7812,N_7746,N_7701);
or U7813 (N_7813,N_7660,N_7614);
nor U7814 (N_7814,N_7646,N_7667);
nor U7815 (N_7815,N_7764,N_7704);
and U7816 (N_7816,N_7761,N_7609);
and U7817 (N_7817,N_7691,N_7703);
and U7818 (N_7818,N_7647,N_7769);
and U7819 (N_7819,N_7752,N_7710);
or U7820 (N_7820,N_7794,N_7698);
nand U7821 (N_7821,N_7650,N_7753);
and U7822 (N_7822,N_7773,N_7679);
nand U7823 (N_7823,N_7728,N_7618);
and U7824 (N_7824,N_7781,N_7754);
and U7825 (N_7825,N_7686,N_7736);
xnor U7826 (N_7826,N_7690,N_7700);
or U7827 (N_7827,N_7648,N_7725);
xnor U7828 (N_7828,N_7642,N_7621);
xnor U7829 (N_7829,N_7676,N_7664);
nand U7830 (N_7830,N_7735,N_7737);
nand U7831 (N_7831,N_7626,N_7636);
nand U7832 (N_7832,N_7638,N_7780);
and U7833 (N_7833,N_7757,N_7771);
or U7834 (N_7834,N_7796,N_7601);
nor U7835 (N_7835,N_7668,N_7762);
nor U7836 (N_7836,N_7782,N_7730);
and U7837 (N_7837,N_7677,N_7639);
nor U7838 (N_7838,N_7635,N_7740);
and U7839 (N_7839,N_7770,N_7756);
and U7840 (N_7840,N_7717,N_7637);
nor U7841 (N_7841,N_7727,N_7617);
nand U7842 (N_7842,N_7696,N_7705);
and U7843 (N_7843,N_7624,N_7629);
nor U7844 (N_7844,N_7674,N_7760);
or U7845 (N_7845,N_7692,N_7790);
nand U7846 (N_7846,N_7658,N_7707);
nor U7847 (N_7847,N_7714,N_7608);
nor U7848 (N_7848,N_7689,N_7654);
or U7849 (N_7849,N_7678,N_7693);
or U7850 (N_7850,N_7697,N_7768);
and U7851 (N_7851,N_7610,N_7649);
nor U7852 (N_7852,N_7765,N_7708);
and U7853 (N_7853,N_7767,N_7716);
nand U7854 (N_7854,N_7680,N_7784);
xor U7855 (N_7855,N_7743,N_7619);
or U7856 (N_7856,N_7791,N_7731);
or U7857 (N_7857,N_7627,N_7606);
xor U7858 (N_7858,N_7659,N_7651);
and U7859 (N_7859,N_7750,N_7788);
xor U7860 (N_7860,N_7672,N_7681);
nand U7861 (N_7861,N_7774,N_7652);
or U7862 (N_7862,N_7662,N_7632);
or U7863 (N_7863,N_7630,N_7776);
or U7864 (N_7864,N_7687,N_7653);
nor U7865 (N_7865,N_7663,N_7711);
xor U7866 (N_7866,N_7747,N_7755);
or U7867 (N_7867,N_7656,N_7605);
nand U7868 (N_7868,N_7695,N_7600);
or U7869 (N_7869,N_7675,N_7751);
and U7870 (N_7870,N_7783,N_7620);
nand U7871 (N_7871,N_7655,N_7604);
nand U7872 (N_7872,N_7688,N_7724);
or U7873 (N_7873,N_7745,N_7772);
or U7874 (N_7874,N_7732,N_7670);
nor U7875 (N_7875,N_7628,N_7777);
and U7876 (N_7876,N_7615,N_7673);
and U7877 (N_7877,N_7602,N_7766);
or U7878 (N_7878,N_7792,N_7785);
nor U7879 (N_7879,N_7786,N_7612);
nand U7880 (N_7880,N_7616,N_7789);
or U7881 (N_7881,N_7739,N_7694);
nor U7882 (N_7882,N_7798,N_7778);
or U7883 (N_7883,N_7666,N_7702);
or U7884 (N_7884,N_7684,N_7726);
nor U7885 (N_7885,N_7718,N_7799);
nand U7886 (N_7886,N_7625,N_7741);
nor U7887 (N_7887,N_7723,N_7631);
xnor U7888 (N_7888,N_7611,N_7622);
or U7889 (N_7889,N_7682,N_7720);
nand U7890 (N_7890,N_7719,N_7734);
and U7891 (N_7891,N_7787,N_7699);
xnor U7892 (N_7892,N_7758,N_7733);
or U7893 (N_7893,N_7623,N_7775);
and U7894 (N_7894,N_7633,N_7657);
and U7895 (N_7895,N_7641,N_7779);
nand U7896 (N_7896,N_7712,N_7607);
xnor U7897 (N_7897,N_7634,N_7729);
nand U7898 (N_7898,N_7722,N_7709);
and U7899 (N_7899,N_7665,N_7683);
or U7900 (N_7900,N_7799,N_7620);
nand U7901 (N_7901,N_7640,N_7782);
nor U7902 (N_7902,N_7773,N_7664);
nor U7903 (N_7903,N_7609,N_7759);
and U7904 (N_7904,N_7794,N_7624);
xor U7905 (N_7905,N_7678,N_7763);
xnor U7906 (N_7906,N_7754,N_7744);
nor U7907 (N_7907,N_7609,N_7731);
and U7908 (N_7908,N_7790,N_7604);
or U7909 (N_7909,N_7629,N_7779);
or U7910 (N_7910,N_7752,N_7781);
or U7911 (N_7911,N_7730,N_7758);
or U7912 (N_7912,N_7628,N_7622);
and U7913 (N_7913,N_7671,N_7735);
and U7914 (N_7914,N_7644,N_7789);
and U7915 (N_7915,N_7664,N_7669);
nor U7916 (N_7916,N_7623,N_7783);
and U7917 (N_7917,N_7679,N_7754);
nor U7918 (N_7918,N_7776,N_7603);
nand U7919 (N_7919,N_7629,N_7743);
or U7920 (N_7920,N_7635,N_7785);
nor U7921 (N_7921,N_7612,N_7748);
or U7922 (N_7922,N_7705,N_7774);
and U7923 (N_7923,N_7624,N_7772);
or U7924 (N_7924,N_7676,N_7743);
nor U7925 (N_7925,N_7727,N_7670);
nor U7926 (N_7926,N_7627,N_7709);
and U7927 (N_7927,N_7681,N_7722);
nor U7928 (N_7928,N_7765,N_7797);
nand U7929 (N_7929,N_7760,N_7692);
xnor U7930 (N_7930,N_7738,N_7737);
and U7931 (N_7931,N_7677,N_7661);
or U7932 (N_7932,N_7656,N_7776);
and U7933 (N_7933,N_7748,N_7714);
or U7934 (N_7934,N_7648,N_7740);
nand U7935 (N_7935,N_7739,N_7604);
nand U7936 (N_7936,N_7683,N_7715);
and U7937 (N_7937,N_7645,N_7798);
nor U7938 (N_7938,N_7687,N_7793);
nand U7939 (N_7939,N_7672,N_7674);
xor U7940 (N_7940,N_7702,N_7650);
or U7941 (N_7941,N_7715,N_7731);
nand U7942 (N_7942,N_7760,N_7771);
nand U7943 (N_7943,N_7697,N_7641);
and U7944 (N_7944,N_7637,N_7788);
and U7945 (N_7945,N_7769,N_7740);
or U7946 (N_7946,N_7784,N_7643);
or U7947 (N_7947,N_7713,N_7754);
nand U7948 (N_7948,N_7799,N_7658);
nand U7949 (N_7949,N_7790,N_7644);
nor U7950 (N_7950,N_7676,N_7719);
and U7951 (N_7951,N_7799,N_7628);
or U7952 (N_7952,N_7685,N_7736);
and U7953 (N_7953,N_7648,N_7639);
and U7954 (N_7954,N_7722,N_7764);
nor U7955 (N_7955,N_7748,N_7665);
nand U7956 (N_7956,N_7616,N_7608);
and U7957 (N_7957,N_7757,N_7651);
nand U7958 (N_7958,N_7695,N_7687);
and U7959 (N_7959,N_7722,N_7736);
nand U7960 (N_7960,N_7689,N_7745);
or U7961 (N_7961,N_7755,N_7750);
and U7962 (N_7962,N_7662,N_7755);
and U7963 (N_7963,N_7630,N_7698);
or U7964 (N_7964,N_7601,N_7779);
or U7965 (N_7965,N_7758,N_7645);
and U7966 (N_7966,N_7647,N_7626);
and U7967 (N_7967,N_7710,N_7628);
and U7968 (N_7968,N_7659,N_7767);
nand U7969 (N_7969,N_7648,N_7749);
or U7970 (N_7970,N_7798,N_7622);
xor U7971 (N_7971,N_7658,N_7633);
nor U7972 (N_7972,N_7642,N_7781);
and U7973 (N_7973,N_7737,N_7719);
or U7974 (N_7974,N_7754,N_7655);
and U7975 (N_7975,N_7663,N_7636);
or U7976 (N_7976,N_7651,N_7602);
and U7977 (N_7977,N_7697,N_7761);
nor U7978 (N_7978,N_7717,N_7711);
xnor U7979 (N_7979,N_7665,N_7754);
nand U7980 (N_7980,N_7614,N_7647);
and U7981 (N_7981,N_7605,N_7629);
and U7982 (N_7982,N_7784,N_7711);
nor U7983 (N_7983,N_7608,N_7601);
nor U7984 (N_7984,N_7755,N_7707);
nand U7985 (N_7985,N_7601,N_7633);
or U7986 (N_7986,N_7732,N_7733);
or U7987 (N_7987,N_7782,N_7609);
and U7988 (N_7988,N_7751,N_7653);
and U7989 (N_7989,N_7777,N_7798);
nand U7990 (N_7990,N_7683,N_7611);
and U7991 (N_7991,N_7728,N_7781);
or U7992 (N_7992,N_7711,N_7686);
nand U7993 (N_7993,N_7602,N_7751);
nand U7994 (N_7994,N_7749,N_7785);
nand U7995 (N_7995,N_7687,N_7738);
or U7996 (N_7996,N_7742,N_7678);
and U7997 (N_7997,N_7791,N_7779);
nor U7998 (N_7998,N_7780,N_7772);
nand U7999 (N_7999,N_7728,N_7771);
and U8000 (N_8000,N_7823,N_7839);
and U8001 (N_8001,N_7919,N_7960);
or U8002 (N_8002,N_7860,N_7817);
nor U8003 (N_8003,N_7807,N_7924);
and U8004 (N_8004,N_7851,N_7829);
or U8005 (N_8005,N_7950,N_7991);
nand U8006 (N_8006,N_7930,N_7844);
nor U8007 (N_8007,N_7842,N_7867);
nor U8008 (N_8008,N_7893,N_7902);
nor U8009 (N_8009,N_7800,N_7853);
and U8010 (N_8010,N_7918,N_7885);
nor U8011 (N_8011,N_7959,N_7875);
or U8012 (N_8012,N_7951,N_7891);
or U8013 (N_8013,N_7838,N_7929);
or U8014 (N_8014,N_7808,N_7928);
and U8015 (N_8015,N_7856,N_7909);
or U8016 (N_8016,N_7922,N_7944);
and U8017 (N_8017,N_7819,N_7814);
nor U8018 (N_8018,N_7926,N_7888);
nand U8019 (N_8019,N_7958,N_7970);
nand U8020 (N_8020,N_7858,N_7957);
nand U8021 (N_8021,N_7884,N_7892);
or U8022 (N_8022,N_7947,N_7973);
or U8023 (N_8023,N_7980,N_7832);
nand U8024 (N_8024,N_7913,N_7835);
nand U8025 (N_8025,N_7910,N_7837);
xor U8026 (N_8026,N_7868,N_7932);
xnor U8027 (N_8027,N_7996,N_7914);
or U8028 (N_8028,N_7849,N_7995);
nor U8029 (N_8029,N_7916,N_7900);
nor U8030 (N_8030,N_7816,N_7953);
nand U8031 (N_8031,N_7968,N_7828);
xor U8032 (N_8032,N_7825,N_7869);
or U8033 (N_8033,N_7852,N_7933);
nor U8034 (N_8034,N_7964,N_7982);
xnor U8035 (N_8035,N_7946,N_7896);
nor U8036 (N_8036,N_7861,N_7988);
nand U8037 (N_8037,N_7952,N_7976);
and U8038 (N_8038,N_7941,N_7989);
and U8039 (N_8039,N_7859,N_7863);
and U8040 (N_8040,N_7881,N_7984);
or U8041 (N_8041,N_7834,N_7820);
or U8042 (N_8042,N_7843,N_7812);
or U8043 (N_8043,N_7879,N_7890);
xnor U8044 (N_8044,N_7809,N_7985);
xnor U8045 (N_8045,N_7865,N_7945);
nand U8046 (N_8046,N_7850,N_7971);
nor U8047 (N_8047,N_7855,N_7877);
nand U8048 (N_8048,N_7912,N_7998);
nand U8049 (N_8049,N_7978,N_7811);
and U8050 (N_8050,N_7871,N_7937);
or U8051 (N_8051,N_7904,N_7975);
and U8052 (N_8052,N_7961,N_7899);
or U8053 (N_8053,N_7986,N_7931);
and U8054 (N_8054,N_7894,N_7872);
and U8055 (N_8055,N_7954,N_7873);
nor U8056 (N_8056,N_7848,N_7939);
nor U8057 (N_8057,N_7956,N_7936);
nor U8058 (N_8058,N_7818,N_7925);
or U8059 (N_8059,N_7907,N_7921);
and U8060 (N_8060,N_7955,N_7830);
or U8061 (N_8061,N_7948,N_7847);
or U8062 (N_8062,N_7864,N_7805);
and U8063 (N_8063,N_7898,N_7927);
and U8064 (N_8064,N_7942,N_7870);
nor U8065 (N_8065,N_7857,N_7827);
nor U8066 (N_8066,N_7846,N_7878);
or U8067 (N_8067,N_7963,N_7840);
or U8068 (N_8068,N_7979,N_7962);
nor U8069 (N_8069,N_7802,N_7806);
nand U8070 (N_8070,N_7949,N_7908);
or U8071 (N_8071,N_7997,N_7969);
and U8072 (N_8072,N_7990,N_7915);
nand U8073 (N_8073,N_7874,N_7935);
nand U8074 (N_8074,N_7826,N_7972);
and U8075 (N_8075,N_7999,N_7813);
nand U8076 (N_8076,N_7886,N_7845);
nor U8077 (N_8077,N_7889,N_7895);
or U8078 (N_8078,N_7824,N_7993);
nand U8079 (N_8079,N_7883,N_7822);
nor U8080 (N_8080,N_7882,N_7801);
and U8081 (N_8081,N_7943,N_7803);
nor U8082 (N_8082,N_7876,N_7831);
or U8083 (N_8083,N_7974,N_7836);
and U8084 (N_8084,N_7887,N_7862);
xor U8085 (N_8085,N_7880,N_7992);
nor U8086 (N_8086,N_7901,N_7897);
and U8087 (N_8087,N_7854,N_7967);
nand U8088 (N_8088,N_7994,N_7810);
nor U8089 (N_8089,N_7923,N_7934);
nor U8090 (N_8090,N_7815,N_7917);
nand U8091 (N_8091,N_7841,N_7983);
or U8092 (N_8092,N_7905,N_7866);
and U8093 (N_8093,N_7821,N_7906);
or U8094 (N_8094,N_7987,N_7911);
nor U8095 (N_8095,N_7965,N_7833);
nand U8096 (N_8096,N_7903,N_7940);
or U8097 (N_8097,N_7938,N_7804);
nor U8098 (N_8098,N_7966,N_7981);
xnor U8099 (N_8099,N_7977,N_7920);
nor U8100 (N_8100,N_7802,N_7973);
nand U8101 (N_8101,N_7814,N_7866);
nand U8102 (N_8102,N_7982,N_7899);
nand U8103 (N_8103,N_7966,N_7903);
xor U8104 (N_8104,N_7899,N_7897);
or U8105 (N_8105,N_7840,N_7817);
xor U8106 (N_8106,N_7825,N_7888);
and U8107 (N_8107,N_7839,N_7979);
or U8108 (N_8108,N_7987,N_7957);
xnor U8109 (N_8109,N_7991,N_7912);
and U8110 (N_8110,N_7816,N_7861);
and U8111 (N_8111,N_7813,N_7850);
or U8112 (N_8112,N_7816,N_7833);
nand U8113 (N_8113,N_7817,N_7991);
and U8114 (N_8114,N_7847,N_7869);
nor U8115 (N_8115,N_7847,N_7852);
and U8116 (N_8116,N_7868,N_7971);
nand U8117 (N_8117,N_7976,N_7896);
or U8118 (N_8118,N_7816,N_7842);
and U8119 (N_8119,N_7838,N_7837);
nand U8120 (N_8120,N_7964,N_7949);
nor U8121 (N_8121,N_7956,N_7861);
nor U8122 (N_8122,N_7858,N_7966);
nor U8123 (N_8123,N_7888,N_7953);
nor U8124 (N_8124,N_7949,N_7918);
or U8125 (N_8125,N_7917,N_7940);
nor U8126 (N_8126,N_7832,N_7935);
or U8127 (N_8127,N_7975,N_7848);
nand U8128 (N_8128,N_7821,N_7824);
or U8129 (N_8129,N_7847,N_7918);
and U8130 (N_8130,N_7807,N_7860);
and U8131 (N_8131,N_7863,N_7852);
nor U8132 (N_8132,N_7992,N_7911);
nand U8133 (N_8133,N_7823,N_7846);
nand U8134 (N_8134,N_7925,N_7884);
nand U8135 (N_8135,N_7994,N_7906);
or U8136 (N_8136,N_7966,N_7827);
and U8137 (N_8137,N_7975,N_7968);
nor U8138 (N_8138,N_7898,N_7932);
xnor U8139 (N_8139,N_7884,N_7849);
nor U8140 (N_8140,N_7877,N_7932);
and U8141 (N_8141,N_7980,N_7853);
and U8142 (N_8142,N_7919,N_7987);
nor U8143 (N_8143,N_7982,N_7823);
or U8144 (N_8144,N_7893,N_7884);
xnor U8145 (N_8145,N_7903,N_7812);
nand U8146 (N_8146,N_7887,N_7872);
nand U8147 (N_8147,N_7987,N_7905);
nor U8148 (N_8148,N_7893,N_7989);
and U8149 (N_8149,N_7856,N_7962);
nand U8150 (N_8150,N_7802,N_7949);
or U8151 (N_8151,N_7858,N_7891);
nor U8152 (N_8152,N_7960,N_7953);
xor U8153 (N_8153,N_7897,N_7822);
nand U8154 (N_8154,N_7982,N_7849);
or U8155 (N_8155,N_7844,N_7853);
or U8156 (N_8156,N_7969,N_7957);
or U8157 (N_8157,N_7942,N_7925);
or U8158 (N_8158,N_7991,N_7847);
and U8159 (N_8159,N_7851,N_7983);
nor U8160 (N_8160,N_7871,N_7862);
or U8161 (N_8161,N_7885,N_7967);
or U8162 (N_8162,N_7986,N_7871);
nor U8163 (N_8163,N_7824,N_7978);
nand U8164 (N_8164,N_7895,N_7955);
nor U8165 (N_8165,N_7953,N_7815);
nand U8166 (N_8166,N_7967,N_7844);
xnor U8167 (N_8167,N_7977,N_7864);
xnor U8168 (N_8168,N_7909,N_7905);
or U8169 (N_8169,N_7806,N_7814);
and U8170 (N_8170,N_7935,N_7892);
and U8171 (N_8171,N_7957,N_7880);
nor U8172 (N_8172,N_7847,N_7932);
nor U8173 (N_8173,N_7919,N_7957);
nand U8174 (N_8174,N_7872,N_7993);
or U8175 (N_8175,N_7930,N_7977);
xnor U8176 (N_8176,N_7875,N_7828);
or U8177 (N_8177,N_7866,N_7901);
nor U8178 (N_8178,N_7999,N_7873);
or U8179 (N_8179,N_7879,N_7960);
xor U8180 (N_8180,N_7810,N_7915);
nand U8181 (N_8181,N_7864,N_7832);
nor U8182 (N_8182,N_7851,N_7957);
or U8183 (N_8183,N_7801,N_7970);
and U8184 (N_8184,N_7862,N_7805);
xor U8185 (N_8185,N_7931,N_7937);
nor U8186 (N_8186,N_7899,N_7913);
or U8187 (N_8187,N_7911,N_7954);
nor U8188 (N_8188,N_7869,N_7836);
or U8189 (N_8189,N_7879,N_7911);
nand U8190 (N_8190,N_7978,N_7896);
or U8191 (N_8191,N_7880,N_7847);
nor U8192 (N_8192,N_7814,N_7996);
nand U8193 (N_8193,N_7961,N_7834);
nor U8194 (N_8194,N_7980,N_7929);
nor U8195 (N_8195,N_7869,N_7854);
and U8196 (N_8196,N_7934,N_7945);
nand U8197 (N_8197,N_7841,N_7955);
nand U8198 (N_8198,N_7834,N_7856);
nor U8199 (N_8199,N_7816,N_7826);
and U8200 (N_8200,N_8060,N_8122);
or U8201 (N_8201,N_8033,N_8096);
and U8202 (N_8202,N_8013,N_8084);
and U8203 (N_8203,N_8154,N_8164);
nor U8204 (N_8204,N_8098,N_8146);
or U8205 (N_8205,N_8037,N_8088);
or U8206 (N_8206,N_8021,N_8167);
and U8207 (N_8207,N_8192,N_8162);
xor U8208 (N_8208,N_8017,N_8090);
and U8209 (N_8209,N_8077,N_8151);
nor U8210 (N_8210,N_8115,N_8067);
and U8211 (N_8211,N_8168,N_8030);
nand U8212 (N_8212,N_8047,N_8080);
and U8213 (N_8213,N_8092,N_8005);
nor U8214 (N_8214,N_8051,N_8139);
and U8215 (N_8215,N_8123,N_8172);
nand U8216 (N_8216,N_8052,N_8045);
nand U8217 (N_8217,N_8012,N_8050);
or U8218 (N_8218,N_8023,N_8097);
nand U8219 (N_8219,N_8155,N_8177);
nor U8220 (N_8220,N_8141,N_8100);
nor U8221 (N_8221,N_8016,N_8102);
nor U8222 (N_8222,N_8114,N_8056);
and U8223 (N_8223,N_8101,N_8048);
nor U8224 (N_8224,N_8156,N_8130);
nand U8225 (N_8225,N_8059,N_8027);
or U8226 (N_8226,N_8093,N_8001);
xor U8227 (N_8227,N_8113,N_8182);
nand U8228 (N_8228,N_8178,N_8112);
nor U8229 (N_8229,N_8035,N_8198);
and U8230 (N_8230,N_8064,N_8085);
or U8231 (N_8231,N_8002,N_8186);
or U8232 (N_8232,N_8135,N_8194);
nor U8233 (N_8233,N_8118,N_8127);
or U8234 (N_8234,N_8148,N_8058);
nand U8235 (N_8235,N_8110,N_8036);
or U8236 (N_8236,N_8028,N_8150);
and U8237 (N_8237,N_8137,N_8007);
nand U8238 (N_8238,N_8095,N_8171);
nor U8239 (N_8239,N_8116,N_8176);
and U8240 (N_8240,N_8000,N_8189);
nand U8241 (N_8241,N_8166,N_8183);
and U8242 (N_8242,N_8180,N_8163);
and U8243 (N_8243,N_8055,N_8145);
nor U8244 (N_8244,N_8074,N_8026);
xnor U8245 (N_8245,N_8143,N_8065);
nand U8246 (N_8246,N_8117,N_8108);
nor U8247 (N_8247,N_8069,N_8039);
xnor U8248 (N_8248,N_8041,N_8042);
nor U8249 (N_8249,N_8157,N_8132);
nor U8250 (N_8250,N_8054,N_8008);
or U8251 (N_8251,N_8179,N_8019);
and U8252 (N_8252,N_8111,N_8086);
nand U8253 (N_8253,N_8099,N_8073);
or U8254 (N_8254,N_8004,N_8089);
xor U8255 (N_8255,N_8032,N_8181);
xor U8256 (N_8256,N_8131,N_8107);
nor U8257 (N_8257,N_8044,N_8124);
xor U8258 (N_8258,N_8106,N_8191);
and U8259 (N_8259,N_8072,N_8003);
nor U8260 (N_8260,N_8199,N_8109);
nand U8261 (N_8261,N_8015,N_8062);
nor U8262 (N_8262,N_8120,N_8147);
nor U8263 (N_8263,N_8082,N_8057);
and U8264 (N_8264,N_8066,N_8121);
and U8265 (N_8265,N_8128,N_8197);
or U8266 (N_8266,N_8138,N_8031);
nand U8267 (N_8267,N_8076,N_8175);
and U8268 (N_8268,N_8094,N_8075);
and U8269 (N_8269,N_8185,N_8125);
nor U8270 (N_8270,N_8068,N_8024);
and U8271 (N_8271,N_8020,N_8129);
and U8272 (N_8272,N_8144,N_8025);
nand U8273 (N_8273,N_8104,N_8195);
or U8274 (N_8274,N_8142,N_8152);
and U8275 (N_8275,N_8136,N_8070);
nor U8276 (N_8276,N_8061,N_8196);
or U8277 (N_8277,N_8034,N_8149);
nand U8278 (N_8278,N_8119,N_8193);
or U8279 (N_8279,N_8006,N_8091);
xnor U8280 (N_8280,N_8046,N_8173);
nand U8281 (N_8281,N_8018,N_8029);
and U8282 (N_8282,N_8010,N_8159);
and U8283 (N_8283,N_8083,N_8134);
or U8284 (N_8284,N_8187,N_8011);
xnor U8285 (N_8285,N_8190,N_8014);
nor U8286 (N_8286,N_8103,N_8022);
nor U8287 (N_8287,N_8169,N_8184);
nor U8288 (N_8288,N_8160,N_8165);
xor U8289 (N_8289,N_8038,N_8079);
nand U8290 (N_8290,N_8174,N_8071);
nor U8291 (N_8291,N_8040,N_8078);
nand U8292 (N_8292,N_8009,N_8133);
nand U8293 (N_8293,N_8043,N_8170);
nor U8294 (N_8294,N_8188,N_8105);
nor U8295 (N_8295,N_8081,N_8087);
and U8296 (N_8296,N_8053,N_8063);
nand U8297 (N_8297,N_8126,N_8161);
and U8298 (N_8298,N_8049,N_8140);
nand U8299 (N_8299,N_8158,N_8153);
xnor U8300 (N_8300,N_8037,N_8157);
nand U8301 (N_8301,N_8170,N_8096);
nor U8302 (N_8302,N_8084,N_8045);
and U8303 (N_8303,N_8099,N_8142);
nor U8304 (N_8304,N_8164,N_8112);
or U8305 (N_8305,N_8183,N_8003);
and U8306 (N_8306,N_8020,N_8032);
nand U8307 (N_8307,N_8141,N_8104);
and U8308 (N_8308,N_8063,N_8111);
nand U8309 (N_8309,N_8019,N_8184);
nor U8310 (N_8310,N_8027,N_8058);
or U8311 (N_8311,N_8034,N_8081);
nor U8312 (N_8312,N_8112,N_8131);
and U8313 (N_8313,N_8068,N_8166);
or U8314 (N_8314,N_8058,N_8183);
and U8315 (N_8315,N_8094,N_8144);
or U8316 (N_8316,N_8110,N_8145);
nand U8317 (N_8317,N_8183,N_8168);
nand U8318 (N_8318,N_8198,N_8012);
or U8319 (N_8319,N_8038,N_8072);
or U8320 (N_8320,N_8181,N_8178);
nor U8321 (N_8321,N_8011,N_8046);
and U8322 (N_8322,N_8106,N_8077);
and U8323 (N_8323,N_8186,N_8177);
nand U8324 (N_8324,N_8047,N_8026);
nand U8325 (N_8325,N_8047,N_8020);
or U8326 (N_8326,N_8044,N_8183);
nor U8327 (N_8327,N_8090,N_8098);
and U8328 (N_8328,N_8101,N_8015);
nand U8329 (N_8329,N_8020,N_8068);
or U8330 (N_8330,N_8141,N_8071);
nor U8331 (N_8331,N_8115,N_8125);
nand U8332 (N_8332,N_8015,N_8198);
and U8333 (N_8333,N_8084,N_8126);
nor U8334 (N_8334,N_8053,N_8132);
nor U8335 (N_8335,N_8080,N_8020);
nor U8336 (N_8336,N_8028,N_8059);
nand U8337 (N_8337,N_8182,N_8114);
or U8338 (N_8338,N_8160,N_8177);
xnor U8339 (N_8339,N_8186,N_8089);
nand U8340 (N_8340,N_8192,N_8010);
and U8341 (N_8341,N_8182,N_8142);
or U8342 (N_8342,N_8042,N_8119);
and U8343 (N_8343,N_8083,N_8070);
nor U8344 (N_8344,N_8193,N_8157);
or U8345 (N_8345,N_8049,N_8070);
nor U8346 (N_8346,N_8034,N_8127);
nand U8347 (N_8347,N_8010,N_8174);
nand U8348 (N_8348,N_8151,N_8141);
nor U8349 (N_8349,N_8046,N_8121);
xnor U8350 (N_8350,N_8185,N_8042);
and U8351 (N_8351,N_8175,N_8046);
and U8352 (N_8352,N_8141,N_8069);
or U8353 (N_8353,N_8039,N_8030);
nor U8354 (N_8354,N_8069,N_8191);
nand U8355 (N_8355,N_8108,N_8097);
nor U8356 (N_8356,N_8048,N_8073);
and U8357 (N_8357,N_8055,N_8047);
nand U8358 (N_8358,N_8111,N_8171);
and U8359 (N_8359,N_8087,N_8168);
nand U8360 (N_8360,N_8020,N_8082);
nor U8361 (N_8361,N_8061,N_8098);
nor U8362 (N_8362,N_8097,N_8056);
or U8363 (N_8363,N_8050,N_8061);
nor U8364 (N_8364,N_8159,N_8000);
nand U8365 (N_8365,N_8052,N_8011);
nor U8366 (N_8366,N_8124,N_8057);
nor U8367 (N_8367,N_8029,N_8034);
nor U8368 (N_8368,N_8131,N_8080);
nand U8369 (N_8369,N_8050,N_8188);
nor U8370 (N_8370,N_8042,N_8050);
and U8371 (N_8371,N_8139,N_8095);
nor U8372 (N_8372,N_8188,N_8013);
or U8373 (N_8373,N_8023,N_8076);
nor U8374 (N_8374,N_8065,N_8166);
or U8375 (N_8375,N_8058,N_8113);
nor U8376 (N_8376,N_8194,N_8030);
nor U8377 (N_8377,N_8116,N_8036);
or U8378 (N_8378,N_8198,N_8041);
nand U8379 (N_8379,N_8062,N_8090);
or U8380 (N_8380,N_8191,N_8123);
xnor U8381 (N_8381,N_8058,N_8087);
and U8382 (N_8382,N_8067,N_8000);
or U8383 (N_8383,N_8079,N_8071);
xnor U8384 (N_8384,N_8198,N_8052);
nand U8385 (N_8385,N_8018,N_8187);
xnor U8386 (N_8386,N_8162,N_8177);
nand U8387 (N_8387,N_8030,N_8152);
nand U8388 (N_8388,N_8087,N_8006);
nor U8389 (N_8389,N_8029,N_8064);
nand U8390 (N_8390,N_8026,N_8107);
and U8391 (N_8391,N_8146,N_8014);
or U8392 (N_8392,N_8131,N_8001);
nor U8393 (N_8393,N_8002,N_8067);
nand U8394 (N_8394,N_8147,N_8161);
nand U8395 (N_8395,N_8096,N_8125);
xor U8396 (N_8396,N_8114,N_8092);
nor U8397 (N_8397,N_8181,N_8110);
and U8398 (N_8398,N_8072,N_8151);
or U8399 (N_8399,N_8012,N_8119);
nand U8400 (N_8400,N_8292,N_8288);
nand U8401 (N_8401,N_8228,N_8224);
xnor U8402 (N_8402,N_8332,N_8327);
nand U8403 (N_8403,N_8230,N_8213);
and U8404 (N_8404,N_8218,N_8319);
nor U8405 (N_8405,N_8347,N_8343);
nand U8406 (N_8406,N_8296,N_8291);
and U8407 (N_8407,N_8317,N_8246);
nor U8408 (N_8408,N_8366,N_8265);
and U8409 (N_8409,N_8346,N_8293);
nor U8410 (N_8410,N_8252,N_8242);
xor U8411 (N_8411,N_8380,N_8338);
nor U8412 (N_8412,N_8391,N_8305);
or U8413 (N_8413,N_8370,N_8356);
nand U8414 (N_8414,N_8303,N_8386);
or U8415 (N_8415,N_8276,N_8358);
and U8416 (N_8416,N_8304,N_8244);
nand U8417 (N_8417,N_8340,N_8235);
xor U8418 (N_8418,N_8255,N_8282);
or U8419 (N_8419,N_8378,N_8368);
xnor U8420 (N_8420,N_8257,N_8362);
nor U8421 (N_8421,N_8321,N_8234);
and U8422 (N_8422,N_8207,N_8328);
and U8423 (N_8423,N_8239,N_8220);
or U8424 (N_8424,N_8385,N_8278);
nand U8425 (N_8425,N_8384,N_8333);
nor U8426 (N_8426,N_8295,N_8351);
or U8427 (N_8427,N_8229,N_8302);
or U8428 (N_8428,N_8271,N_8337);
and U8429 (N_8429,N_8249,N_8330);
nor U8430 (N_8430,N_8397,N_8399);
and U8431 (N_8431,N_8254,N_8212);
and U8432 (N_8432,N_8201,N_8313);
nand U8433 (N_8433,N_8318,N_8316);
nand U8434 (N_8434,N_8352,N_8222);
and U8435 (N_8435,N_8208,N_8205);
nand U8436 (N_8436,N_8240,N_8398);
nor U8437 (N_8437,N_8396,N_8261);
or U8438 (N_8438,N_8245,N_8393);
nor U8439 (N_8439,N_8355,N_8206);
or U8440 (N_8440,N_8273,N_8280);
and U8441 (N_8441,N_8367,N_8307);
or U8442 (N_8442,N_8357,N_8379);
xnor U8443 (N_8443,N_8204,N_8348);
nor U8444 (N_8444,N_8217,N_8350);
and U8445 (N_8445,N_8241,N_8359);
nor U8446 (N_8446,N_8232,N_8312);
nand U8447 (N_8447,N_8284,N_8383);
nor U8448 (N_8448,N_8376,N_8388);
or U8449 (N_8449,N_8311,N_8381);
xnor U8450 (N_8450,N_8285,N_8334);
nand U8451 (N_8451,N_8270,N_8286);
nor U8452 (N_8452,N_8315,N_8267);
and U8453 (N_8453,N_8353,N_8266);
nor U8454 (N_8454,N_8223,N_8236);
xor U8455 (N_8455,N_8221,N_8344);
or U8456 (N_8456,N_8210,N_8211);
or U8457 (N_8457,N_8309,N_8268);
nor U8458 (N_8458,N_8365,N_8226);
or U8459 (N_8459,N_8320,N_8325);
nand U8460 (N_8460,N_8203,N_8294);
and U8461 (N_8461,N_8287,N_8256);
nand U8462 (N_8462,N_8237,N_8300);
nor U8463 (N_8463,N_8275,N_8247);
nand U8464 (N_8464,N_8277,N_8243);
nor U8465 (N_8465,N_8377,N_8324);
or U8466 (N_8466,N_8323,N_8336);
and U8467 (N_8467,N_8390,N_8341);
and U8468 (N_8468,N_8250,N_8345);
nand U8469 (N_8469,N_8363,N_8349);
and U8470 (N_8470,N_8361,N_8299);
and U8471 (N_8471,N_8251,N_8301);
and U8472 (N_8472,N_8354,N_8297);
xor U8473 (N_8473,N_8269,N_8253);
nor U8474 (N_8474,N_8342,N_8289);
nor U8475 (N_8475,N_8274,N_8231);
and U8476 (N_8476,N_8372,N_8214);
and U8477 (N_8477,N_8290,N_8279);
nand U8478 (N_8478,N_8248,N_8225);
nand U8479 (N_8479,N_8310,N_8308);
nand U8480 (N_8480,N_8202,N_8314);
nand U8481 (N_8481,N_8306,N_8389);
and U8482 (N_8482,N_8259,N_8298);
nand U8483 (N_8483,N_8373,N_8394);
and U8484 (N_8484,N_8331,N_8264);
or U8485 (N_8485,N_8326,N_8375);
and U8486 (N_8486,N_8216,N_8371);
or U8487 (N_8487,N_8200,N_8322);
and U8488 (N_8488,N_8360,N_8329);
xor U8489 (N_8489,N_8258,N_8215);
and U8490 (N_8490,N_8395,N_8227);
nor U8491 (N_8491,N_8262,N_8219);
or U8492 (N_8492,N_8339,N_8364);
or U8493 (N_8493,N_8283,N_8260);
nand U8494 (N_8494,N_8272,N_8392);
nor U8495 (N_8495,N_8233,N_8374);
nor U8496 (N_8496,N_8238,N_8369);
nand U8497 (N_8497,N_8281,N_8263);
and U8498 (N_8498,N_8335,N_8382);
nor U8499 (N_8499,N_8387,N_8209);
xnor U8500 (N_8500,N_8338,N_8371);
nor U8501 (N_8501,N_8279,N_8376);
and U8502 (N_8502,N_8248,N_8343);
or U8503 (N_8503,N_8237,N_8292);
nand U8504 (N_8504,N_8339,N_8350);
or U8505 (N_8505,N_8241,N_8324);
or U8506 (N_8506,N_8383,N_8237);
nand U8507 (N_8507,N_8359,N_8333);
nor U8508 (N_8508,N_8252,N_8201);
or U8509 (N_8509,N_8270,N_8206);
or U8510 (N_8510,N_8232,N_8240);
nand U8511 (N_8511,N_8200,N_8232);
or U8512 (N_8512,N_8330,N_8337);
nand U8513 (N_8513,N_8297,N_8341);
and U8514 (N_8514,N_8304,N_8318);
or U8515 (N_8515,N_8304,N_8351);
nand U8516 (N_8516,N_8241,N_8320);
and U8517 (N_8517,N_8205,N_8280);
and U8518 (N_8518,N_8389,N_8355);
or U8519 (N_8519,N_8275,N_8307);
and U8520 (N_8520,N_8322,N_8350);
nor U8521 (N_8521,N_8351,N_8267);
xor U8522 (N_8522,N_8399,N_8328);
nor U8523 (N_8523,N_8311,N_8262);
nand U8524 (N_8524,N_8250,N_8263);
and U8525 (N_8525,N_8205,N_8276);
nand U8526 (N_8526,N_8250,N_8374);
and U8527 (N_8527,N_8231,N_8351);
or U8528 (N_8528,N_8244,N_8356);
nor U8529 (N_8529,N_8344,N_8330);
nor U8530 (N_8530,N_8250,N_8236);
or U8531 (N_8531,N_8390,N_8209);
and U8532 (N_8532,N_8252,N_8235);
nor U8533 (N_8533,N_8271,N_8219);
nand U8534 (N_8534,N_8203,N_8306);
or U8535 (N_8535,N_8294,N_8301);
nor U8536 (N_8536,N_8291,N_8239);
xor U8537 (N_8537,N_8250,N_8300);
xor U8538 (N_8538,N_8260,N_8241);
nand U8539 (N_8539,N_8225,N_8397);
nor U8540 (N_8540,N_8394,N_8285);
nand U8541 (N_8541,N_8234,N_8339);
and U8542 (N_8542,N_8302,N_8367);
and U8543 (N_8543,N_8278,N_8292);
nand U8544 (N_8544,N_8233,N_8316);
nand U8545 (N_8545,N_8249,N_8399);
or U8546 (N_8546,N_8372,N_8360);
nor U8547 (N_8547,N_8341,N_8353);
xnor U8548 (N_8548,N_8398,N_8362);
or U8549 (N_8549,N_8214,N_8284);
or U8550 (N_8550,N_8241,N_8347);
xnor U8551 (N_8551,N_8351,N_8299);
nand U8552 (N_8552,N_8251,N_8391);
and U8553 (N_8553,N_8395,N_8285);
and U8554 (N_8554,N_8398,N_8367);
and U8555 (N_8555,N_8311,N_8305);
or U8556 (N_8556,N_8258,N_8297);
xor U8557 (N_8557,N_8293,N_8327);
or U8558 (N_8558,N_8257,N_8309);
nor U8559 (N_8559,N_8354,N_8271);
or U8560 (N_8560,N_8366,N_8271);
or U8561 (N_8561,N_8233,N_8251);
nor U8562 (N_8562,N_8207,N_8307);
nand U8563 (N_8563,N_8328,N_8214);
xor U8564 (N_8564,N_8305,N_8389);
nand U8565 (N_8565,N_8302,N_8233);
and U8566 (N_8566,N_8393,N_8223);
and U8567 (N_8567,N_8271,N_8316);
nand U8568 (N_8568,N_8299,N_8277);
or U8569 (N_8569,N_8330,N_8332);
nand U8570 (N_8570,N_8265,N_8223);
and U8571 (N_8571,N_8313,N_8356);
and U8572 (N_8572,N_8335,N_8305);
nand U8573 (N_8573,N_8346,N_8255);
nand U8574 (N_8574,N_8310,N_8321);
and U8575 (N_8575,N_8256,N_8332);
and U8576 (N_8576,N_8305,N_8212);
nand U8577 (N_8577,N_8231,N_8365);
nand U8578 (N_8578,N_8244,N_8380);
nor U8579 (N_8579,N_8238,N_8203);
or U8580 (N_8580,N_8211,N_8391);
nand U8581 (N_8581,N_8385,N_8310);
and U8582 (N_8582,N_8349,N_8352);
and U8583 (N_8583,N_8323,N_8256);
xor U8584 (N_8584,N_8332,N_8391);
xor U8585 (N_8585,N_8271,N_8222);
nand U8586 (N_8586,N_8225,N_8258);
and U8587 (N_8587,N_8293,N_8254);
or U8588 (N_8588,N_8317,N_8257);
nand U8589 (N_8589,N_8260,N_8337);
and U8590 (N_8590,N_8205,N_8236);
nand U8591 (N_8591,N_8200,N_8221);
and U8592 (N_8592,N_8384,N_8392);
nor U8593 (N_8593,N_8311,N_8265);
xor U8594 (N_8594,N_8394,N_8269);
nor U8595 (N_8595,N_8342,N_8204);
and U8596 (N_8596,N_8219,N_8380);
nand U8597 (N_8597,N_8398,N_8324);
nand U8598 (N_8598,N_8341,N_8357);
or U8599 (N_8599,N_8326,N_8245);
xor U8600 (N_8600,N_8504,N_8452);
or U8601 (N_8601,N_8535,N_8496);
nand U8602 (N_8602,N_8514,N_8587);
nor U8603 (N_8603,N_8444,N_8435);
nor U8604 (N_8604,N_8489,N_8508);
and U8605 (N_8605,N_8499,N_8505);
nor U8606 (N_8606,N_8558,N_8468);
and U8607 (N_8607,N_8471,N_8577);
or U8608 (N_8608,N_8556,N_8475);
nand U8609 (N_8609,N_8594,N_8526);
or U8610 (N_8610,N_8456,N_8509);
xor U8611 (N_8611,N_8498,N_8406);
nor U8612 (N_8612,N_8433,N_8573);
or U8613 (N_8613,N_8545,N_8527);
and U8614 (N_8614,N_8497,N_8408);
nor U8615 (N_8615,N_8400,N_8513);
and U8616 (N_8616,N_8418,N_8450);
and U8617 (N_8617,N_8551,N_8448);
xor U8618 (N_8618,N_8552,N_8531);
or U8619 (N_8619,N_8439,N_8485);
and U8620 (N_8620,N_8455,N_8589);
or U8621 (N_8621,N_8595,N_8580);
or U8622 (N_8622,N_8491,N_8454);
or U8623 (N_8623,N_8451,N_8506);
nor U8624 (N_8624,N_8410,N_8554);
nor U8625 (N_8625,N_8518,N_8528);
nand U8626 (N_8626,N_8466,N_8517);
or U8627 (N_8627,N_8578,N_8405);
xnor U8628 (N_8628,N_8481,N_8598);
nor U8629 (N_8629,N_8476,N_8585);
nor U8630 (N_8630,N_8460,N_8576);
or U8631 (N_8631,N_8520,N_8427);
nand U8632 (N_8632,N_8566,N_8474);
or U8633 (N_8633,N_8425,N_8547);
and U8634 (N_8634,N_8442,N_8546);
or U8635 (N_8635,N_8430,N_8540);
and U8636 (N_8636,N_8592,N_8411);
nand U8637 (N_8637,N_8431,N_8412);
and U8638 (N_8638,N_8541,N_8569);
nor U8639 (N_8639,N_8438,N_8416);
nand U8640 (N_8640,N_8525,N_8544);
and U8641 (N_8641,N_8443,N_8420);
nand U8642 (N_8642,N_8424,N_8515);
nand U8643 (N_8643,N_8512,N_8434);
nor U8644 (N_8644,N_8429,N_8523);
or U8645 (N_8645,N_8560,N_8565);
and U8646 (N_8646,N_8524,N_8593);
xor U8647 (N_8647,N_8422,N_8483);
nand U8648 (N_8648,N_8597,N_8529);
nor U8649 (N_8649,N_8486,N_8519);
and U8650 (N_8650,N_8543,N_8413);
nor U8651 (N_8651,N_8599,N_8462);
or U8652 (N_8652,N_8563,N_8473);
nand U8653 (N_8653,N_8579,N_8446);
nor U8654 (N_8654,N_8419,N_8488);
nor U8655 (N_8655,N_8507,N_8472);
or U8656 (N_8656,N_8449,N_8447);
nand U8657 (N_8657,N_8536,N_8494);
or U8658 (N_8658,N_8409,N_8537);
xnor U8659 (N_8659,N_8533,N_8570);
nor U8660 (N_8660,N_8493,N_8500);
nand U8661 (N_8661,N_8440,N_8542);
nand U8662 (N_8662,N_8557,N_8561);
nand U8663 (N_8663,N_8503,N_8467);
and U8664 (N_8664,N_8403,N_8437);
nand U8665 (N_8665,N_8516,N_8550);
or U8666 (N_8666,N_8596,N_8477);
or U8667 (N_8667,N_8490,N_8465);
or U8668 (N_8668,N_8464,N_8584);
nand U8669 (N_8669,N_8539,N_8501);
nor U8670 (N_8670,N_8495,N_8511);
nor U8671 (N_8671,N_8469,N_8417);
or U8672 (N_8672,N_8479,N_8571);
and U8673 (N_8673,N_8463,N_8478);
xor U8674 (N_8674,N_8415,N_8470);
or U8675 (N_8675,N_8453,N_8549);
and U8676 (N_8676,N_8553,N_8436);
and U8677 (N_8677,N_8441,N_8484);
nand U8678 (N_8678,N_8457,N_8530);
or U8679 (N_8679,N_8590,N_8404);
nand U8680 (N_8680,N_8575,N_8534);
and U8681 (N_8681,N_8459,N_8564);
nor U8682 (N_8682,N_8572,N_8583);
nor U8683 (N_8683,N_8568,N_8586);
nor U8684 (N_8684,N_8426,N_8581);
nor U8685 (N_8685,N_8555,N_8521);
or U8686 (N_8686,N_8522,N_8428);
nand U8687 (N_8687,N_8574,N_8401);
and U8688 (N_8688,N_8510,N_8407);
or U8689 (N_8689,N_8458,N_8461);
or U8690 (N_8690,N_8492,N_8548);
xnor U8691 (N_8691,N_8559,N_8402);
and U8692 (N_8692,N_8588,N_8502);
nor U8693 (N_8693,N_8432,N_8480);
nor U8694 (N_8694,N_8482,N_8567);
nor U8695 (N_8695,N_8421,N_8591);
and U8696 (N_8696,N_8538,N_8423);
or U8697 (N_8697,N_8414,N_8562);
nor U8698 (N_8698,N_8487,N_8445);
nand U8699 (N_8699,N_8532,N_8582);
nor U8700 (N_8700,N_8579,N_8565);
nor U8701 (N_8701,N_8598,N_8456);
or U8702 (N_8702,N_8469,N_8435);
xor U8703 (N_8703,N_8570,N_8468);
and U8704 (N_8704,N_8467,N_8547);
xnor U8705 (N_8705,N_8547,N_8544);
nand U8706 (N_8706,N_8575,N_8480);
or U8707 (N_8707,N_8478,N_8473);
xor U8708 (N_8708,N_8457,N_8473);
and U8709 (N_8709,N_8438,N_8442);
and U8710 (N_8710,N_8474,N_8546);
nor U8711 (N_8711,N_8494,N_8563);
nor U8712 (N_8712,N_8420,N_8526);
nand U8713 (N_8713,N_8501,N_8512);
xnor U8714 (N_8714,N_8513,N_8509);
nand U8715 (N_8715,N_8588,N_8418);
nand U8716 (N_8716,N_8483,N_8544);
and U8717 (N_8717,N_8427,N_8433);
nand U8718 (N_8718,N_8571,N_8574);
and U8719 (N_8719,N_8548,N_8565);
and U8720 (N_8720,N_8420,N_8444);
and U8721 (N_8721,N_8475,N_8516);
or U8722 (N_8722,N_8446,N_8505);
nor U8723 (N_8723,N_8550,N_8530);
and U8724 (N_8724,N_8426,N_8555);
or U8725 (N_8725,N_8538,N_8489);
or U8726 (N_8726,N_8500,N_8538);
nor U8727 (N_8727,N_8517,N_8424);
or U8728 (N_8728,N_8564,N_8502);
nand U8729 (N_8729,N_8562,N_8569);
or U8730 (N_8730,N_8571,N_8518);
xor U8731 (N_8731,N_8492,N_8413);
and U8732 (N_8732,N_8588,N_8445);
and U8733 (N_8733,N_8449,N_8588);
nand U8734 (N_8734,N_8460,N_8490);
and U8735 (N_8735,N_8525,N_8508);
nand U8736 (N_8736,N_8586,N_8405);
nand U8737 (N_8737,N_8444,N_8513);
nor U8738 (N_8738,N_8422,N_8554);
nor U8739 (N_8739,N_8418,N_8426);
or U8740 (N_8740,N_8488,N_8486);
xnor U8741 (N_8741,N_8586,N_8549);
or U8742 (N_8742,N_8593,N_8480);
nand U8743 (N_8743,N_8445,N_8562);
xnor U8744 (N_8744,N_8402,N_8495);
nor U8745 (N_8745,N_8582,N_8415);
nand U8746 (N_8746,N_8406,N_8552);
xor U8747 (N_8747,N_8462,N_8476);
xor U8748 (N_8748,N_8590,N_8490);
nand U8749 (N_8749,N_8486,N_8542);
nand U8750 (N_8750,N_8523,N_8570);
nor U8751 (N_8751,N_8418,N_8403);
nand U8752 (N_8752,N_8466,N_8463);
or U8753 (N_8753,N_8435,N_8413);
and U8754 (N_8754,N_8451,N_8584);
or U8755 (N_8755,N_8401,N_8462);
nand U8756 (N_8756,N_8518,N_8471);
nand U8757 (N_8757,N_8538,N_8449);
nand U8758 (N_8758,N_8452,N_8407);
or U8759 (N_8759,N_8470,N_8516);
nor U8760 (N_8760,N_8486,N_8555);
nor U8761 (N_8761,N_8483,N_8541);
nor U8762 (N_8762,N_8505,N_8475);
nor U8763 (N_8763,N_8597,N_8547);
nand U8764 (N_8764,N_8545,N_8432);
nand U8765 (N_8765,N_8528,N_8455);
nand U8766 (N_8766,N_8539,N_8546);
or U8767 (N_8767,N_8539,N_8585);
and U8768 (N_8768,N_8484,N_8478);
or U8769 (N_8769,N_8412,N_8514);
and U8770 (N_8770,N_8476,N_8539);
or U8771 (N_8771,N_8555,N_8423);
nor U8772 (N_8772,N_8495,N_8590);
nand U8773 (N_8773,N_8488,N_8577);
and U8774 (N_8774,N_8561,N_8524);
xor U8775 (N_8775,N_8479,N_8437);
and U8776 (N_8776,N_8549,N_8512);
xor U8777 (N_8777,N_8575,N_8535);
and U8778 (N_8778,N_8456,N_8534);
nor U8779 (N_8779,N_8497,N_8522);
nor U8780 (N_8780,N_8593,N_8583);
nor U8781 (N_8781,N_8552,N_8508);
nand U8782 (N_8782,N_8574,N_8436);
or U8783 (N_8783,N_8566,N_8437);
nand U8784 (N_8784,N_8426,N_8508);
nand U8785 (N_8785,N_8522,N_8481);
or U8786 (N_8786,N_8575,N_8565);
nand U8787 (N_8787,N_8480,N_8468);
and U8788 (N_8788,N_8423,N_8587);
nand U8789 (N_8789,N_8528,N_8477);
or U8790 (N_8790,N_8434,N_8588);
nor U8791 (N_8791,N_8577,N_8506);
and U8792 (N_8792,N_8411,N_8447);
and U8793 (N_8793,N_8445,N_8584);
or U8794 (N_8794,N_8402,N_8421);
nand U8795 (N_8795,N_8548,N_8427);
nand U8796 (N_8796,N_8427,N_8400);
or U8797 (N_8797,N_8528,N_8461);
and U8798 (N_8798,N_8486,N_8593);
nor U8799 (N_8799,N_8590,N_8492);
nand U8800 (N_8800,N_8783,N_8668);
or U8801 (N_8801,N_8725,N_8672);
nand U8802 (N_8802,N_8767,N_8773);
and U8803 (N_8803,N_8721,N_8791);
and U8804 (N_8804,N_8792,N_8716);
or U8805 (N_8805,N_8740,N_8723);
and U8806 (N_8806,N_8770,N_8772);
xnor U8807 (N_8807,N_8646,N_8678);
and U8808 (N_8808,N_8709,N_8621);
xor U8809 (N_8809,N_8613,N_8797);
xor U8810 (N_8810,N_8690,N_8688);
xor U8811 (N_8811,N_8691,N_8776);
or U8812 (N_8812,N_8648,N_8611);
xor U8813 (N_8813,N_8653,N_8609);
nor U8814 (N_8814,N_8781,N_8670);
nand U8815 (N_8815,N_8727,N_8684);
and U8816 (N_8816,N_8707,N_8622);
xnor U8817 (N_8817,N_8625,N_8726);
or U8818 (N_8818,N_8699,N_8711);
nor U8819 (N_8819,N_8654,N_8718);
or U8820 (N_8820,N_8765,N_8751);
nand U8821 (N_8821,N_8616,N_8766);
or U8822 (N_8822,N_8754,N_8680);
nand U8823 (N_8823,N_8750,N_8729);
and U8824 (N_8824,N_8730,N_8758);
and U8825 (N_8825,N_8656,N_8608);
xor U8826 (N_8826,N_8736,N_8756);
xnor U8827 (N_8827,N_8697,N_8657);
nand U8828 (N_8828,N_8719,N_8640);
nand U8829 (N_8829,N_8655,N_8760);
and U8830 (N_8830,N_8687,N_8745);
nor U8831 (N_8831,N_8626,N_8752);
and U8832 (N_8832,N_8780,N_8698);
or U8833 (N_8833,N_8794,N_8681);
nor U8834 (N_8834,N_8706,N_8602);
nor U8835 (N_8835,N_8620,N_8764);
xor U8836 (N_8836,N_8641,N_8617);
nor U8837 (N_8837,N_8636,N_8662);
nand U8838 (N_8838,N_8722,N_8628);
and U8839 (N_8839,N_8658,N_8642);
or U8840 (N_8840,N_8735,N_8650);
or U8841 (N_8841,N_8600,N_8674);
and U8842 (N_8842,N_8633,N_8753);
nor U8843 (N_8843,N_8612,N_8755);
nand U8844 (N_8844,N_8624,N_8649);
or U8845 (N_8845,N_8747,N_8720);
and U8846 (N_8846,N_8771,N_8786);
and U8847 (N_8847,N_8663,N_8683);
nor U8848 (N_8848,N_8774,N_8733);
and U8849 (N_8849,N_8739,N_8601);
nor U8850 (N_8850,N_8741,N_8788);
or U8851 (N_8851,N_8623,N_8666);
and U8852 (N_8852,N_8717,N_8652);
nand U8853 (N_8853,N_8604,N_8700);
nor U8854 (N_8854,N_8714,N_8695);
and U8855 (N_8855,N_8669,N_8664);
and U8856 (N_8856,N_8661,N_8630);
nor U8857 (N_8857,N_8763,N_8677);
nand U8858 (N_8858,N_8702,N_8694);
nand U8859 (N_8859,N_8692,N_8632);
and U8860 (N_8860,N_8749,N_8769);
or U8861 (N_8861,N_8732,N_8713);
or U8862 (N_8862,N_8686,N_8742);
xnor U8863 (N_8863,N_8782,N_8785);
nor U8864 (N_8864,N_8693,N_8610);
or U8865 (N_8865,N_8790,N_8704);
and U8866 (N_8866,N_8761,N_8660);
nand U8867 (N_8867,N_8679,N_8795);
and U8868 (N_8868,N_8768,N_8724);
nor U8869 (N_8869,N_8614,N_8715);
or U8870 (N_8870,N_8671,N_8746);
or U8871 (N_8871,N_8793,N_8667);
nand U8872 (N_8872,N_8635,N_8665);
or U8873 (N_8873,N_8637,N_8748);
nor U8874 (N_8874,N_8631,N_8743);
xor U8875 (N_8875,N_8651,N_8784);
xor U8876 (N_8876,N_8618,N_8682);
and U8877 (N_8877,N_8710,N_8728);
or U8878 (N_8878,N_8789,N_8619);
nor U8879 (N_8879,N_8615,N_8647);
nand U8880 (N_8880,N_8659,N_8603);
or U8881 (N_8881,N_8762,N_8605);
and U8882 (N_8882,N_8644,N_8734);
xnor U8883 (N_8883,N_8703,N_8738);
and U8884 (N_8884,N_8779,N_8775);
and U8885 (N_8885,N_8757,N_8606);
and U8886 (N_8886,N_8629,N_8701);
nor U8887 (N_8887,N_8689,N_8696);
or U8888 (N_8888,N_8799,N_8627);
nand U8889 (N_8889,N_8639,N_8643);
nand U8890 (N_8890,N_8708,N_8777);
or U8891 (N_8891,N_8737,N_8676);
nor U8892 (N_8892,N_8731,N_8778);
nand U8893 (N_8893,N_8634,N_8638);
or U8894 (N_8894,N_8787,N_8645);
or U8895 (N_8895,N_8744,N_8673);
or U8896 (N_8896,N_8685,N_8712);
nor U8897 (N_8897,N_8796,N_8607);
nand U8898 (N_8898,N_8675,N_8705);
xnor U8899 (N_8899,N_8759,N_8798);
and U8900 (N_8900,N_8630,N_8683);
or U8901 (N_8901,N_8605,N_8778);
or U8902 (N_8902,N_8695,N_8600);
or U8903 (N_8903,N_8702,N_8776);
or U8904 (N_8904,N_8654,N_8613);
xor U8905 (N_8905,N_8797,N_8778);
nor U8906 (N_8906,N_8673,N_8713);
or U8907 (N_8907,N_8614,N_8636);
nor U8908 (N_8908,N_8602,N_8784);
and U8909 (N_8909,N_8678,N_8735);
xnor U8910 (N_8910,N_8754,N_8788);
or U8911 (N_8911,N_8741,N_8627);
nor U8912 (N_8912,N_8657,N_8605);
nor U8913 (N_8913,N_8778,N_8799);
and U8914 (N_8914,N_8632,N_8713);
and U8915 (N_8915,N_8654,N_8647);
and U8916 (N_8916,N_8615,N_8760);
and U8917 (N_8917,N_8739,N_8670);
and U8918 (N_8918,N_8736,N_8724);
nand U8919 (N_8919,N_8622,N_8629);
xor U8920 (N_8920,N_8771,N_8691);
nor U8921 (N_8921,N_8769,N_8734);
nand U8922 (N_8922,N_8760,N_8646);
nand U8923 (N_8923,N_8794,N_8646);
and U8924 (N_8924,N_8708,N_8718);
nor U8925 (N_8925,N_8663,N_8755);
nor U8926 (N_8926,N_8609,N_8660);
nor U8927 (N_8927,N_8722,N_8602);
and U8928 (N_8928,N_8657,N_8770);
nor U8929 (N_8929,N_8678,N_8797);
nand U8930 (N_8930,N_8626,N_8644);
or U8931 (N_8931,N_8697,N_8784);
nor U8932 (N_8932,N_8609,N_8600);
nor U8933 (N_8933,N_8659,N_8621);
or U8934 (N_8934,N_8685,N_8664);
or U8935 (N_8935,N_8664,N_8748);
or U8936 (N_8936,N_8639,N_8731);
and U8937 (N_8937,N_8642,N_8720);
nand U8938 (N_8938,N_8702,N_8614);
nor U8939 (N_8939,N_8750,N_8744);
xor U8940 (N_8940,N_8606,N_8640);
nand U8941 (N_8941,N_8612,N_8678);
nand U8942 (N_8942,N_8651,N_8620);
nor U8943 (N_8943,N_8654,N_8713);
or U8944 (N_8944,N_8661,N_8751);
xor U8945 (N_8945,N_8646,N_8746);
and U8946 (N_8946,N_8762,N_8663);
or U8947 (N_8947,N_8715,N_8711);
xnor U8948 (N_8948,N_8620,N_8649);
xor U8949 (N_8949,N_8695,N_8724);
and U8950 (N_8950,N_8665,N_8707);
nand U8951 (N_8951,N_8642,N_8790);
nor U8952 (N_8952,N_8736,N_8603);
nand U8953 (N_8953,N_8655,N_8679);
or U8954 (N_8954,N_8749,N_8618);
and U8955 (N_8955,N_8627,N_8716);
and U8956 (N_8956,N_8650,N_8763);
xnor U8957 (N_8957,N_8666,N_8730);
nor U8958 (N_8958,N_8684,N_8628);
nor U8959 (N_8959,N_8654,N_8618);
or U8960 (N_8960,N_8646,N_8618);
nor U8961 (N_8961,N_8601,N_8761);
xnor U8962 (N_8962,N_8774,N_8615);
and U8963 (N_8963,N_8720,N_8792);
nor U8964 (N_8964,N_8731,N_8663);
nand U8965 (N_8965,N_8661,N_8660);
xnor U8966 (N_8966,N_8603,N_8772);
or U8967 (N_8967,N_8704,N_8666);
or U8968 (N_8968,N_8790,N_8703);
nand U8969 (N_8969,N_8620,N_8660);
nand U8970 (N_8970,N_8659,N_8638);
nor U8971 (N_8971,N_8686,N_8653);
xor U8972 (N_8972,N_8651,N_8787);
xnor U8973 (N_8973,N_8753,N_8746);
nand U8974 (N_8974,N_8741,N_8662);
nand U8975 (N_8975,N_8739,N_8710);
or U8976 (N_8976,N_8706,N_8612);
nand U8977 (N_8977,N_8748,N_8613);
nor U8978 (N_8978,N_8732,N_8746);
or U8979 (N_8979,N_8688,N_8725);
nor U8980 (N_8980,N_8728,N_8626);
and U8981 (N_8981,N_8759,N_8644);
xor U8982 (N_8982,N_8621,N_8657);
nor U8983 (N_8983,N_8657,N_8636);
nor U8984 (N_8984,N_8615,N_8650);
or U8985 (N_8985,N_8728,N_8662);
nand U8986 (N_8986,N_8616,N_8736);
xnor U8987 (N_8987,N_8662,N_8793);
nand U8988 (N_8988,N_8756,N_8797);
and U8989 (N_8989,N_8796,N_8694);
or U8990 (N_8990,N_8784,N_8679);
nor U8991 (N_8991,N_8604,N_8647);
or U8992 (N_8992,N_8676,N_8732);
or U8993 (N_8993,N_8764,N_8677);
and U8994 (N_8994,N_8664,N_8626);
or U8995 (N_8995,N_8710,N_8607);
nor U8996 (N_8996,N_8799,N_8785);
nand U8997 (N_8997,N_8638,N_8762);
and U8998 (N_8998,N_8792,N_8609);
nand U8999 (N_8999,N_8725,N_8653);
xor U9000 (N_9000,N_8985,N_8897);
nor U9001 (N_9001,N_8824,N_8956);
or U9002 (N_9002,N_8911,N_8944);
or U9003 (N_9003,N_8848,N_8872);
xor U9004 (N_9004,N_8979,N_8929);
xnor U9005 (N_9005,N_8925,N_8957);
nand U9006 (N_9006,N_8913,N_8809);
or U9007 (N_9007,N_8899,N_8839);
and U9008 (N_9008,N_8965,N_8973);
nand U9009 (N_9009,N_8998,N_8800);
and U9010 (N_9010,N_8989,N_8914);
nand U9011 (N_9011,N_8894,N_8813);
nand U9012 (N_9012,N_8954,N_8963);
nor U9013 (N_9013,N_8858,N_8938);
nor U9014 (N_9014,N_8801,N_8964);
or U9015 (N_9015,N_8924,N_8833);
or U9016 (N_9016,N_8870,N_8907);
and U9017 (N_9017,N_8902,N_8818);
and U9018 (N_9018,N_8997,N_8857);
or U9019 (N_9019,N_8949,N_8970);
nand U9020 (N_9020,N_8862,N_8923);
nor U9021 (N_9021,N_8971,N_8974);
nand U9022 (N_9022,N_8856,N_8891);
nor U9023 (N_9023,N_8805,N_8827);
nor U9024 (N_9024,N_8961,N_8920);
xnor U9025 (N_9025,N_8823,N_8978);
and U9026 (N_9026,N_8822,N_8812);
xor U9027 (N_9027,N_8868,N_8828);
or U9028 (N_9028,N_8855,N_8987);
or U9029 (N_9029,N_8884,N_8832);
nand U9030 (N_9030,N_8881,N_8843);
or U9031 (N_9031,N_8864,N_8808);
nor U9032 (N_9032,N_8927,N_8951);
nand U9033 (N_9033,N_8810,N_8893);
or U9034 (N_9034,N_8816,N_8948);
or U9035 (N_9035,N_8955,N_8887);
nand U9036 (N_9036,N_8901,N_8815);
xnor U9037 (N_9037,N_8992,N_8986);
nand U9038 (N_9038,N_8874,N_8922);
nand U9039 (N_9039,N_8869,N_8886);
nand U9040 (N_9040,N_8926,N_8936);
nand U9041 (N_9041,N_8969,N_8994);
nand U9042 (N_9042,N_8983,N_8942);
nor U9043 (N_9043,N_8980,N_8885);
and U9044 (N_9044,N_8918,N_8840);
xnor U9045 (N_9045,N_8947,N_8995);
nor U9046 (N_9046,N_8976,N_8958);
nor U9047 (N_9047,N_8866,N_8904);
nor U9048 (N_9048,N_8898,N_8906);
or U9049 (N_9049,N_8841,N_8962);
or U9050 (N_9050,N_8959,N_8953);
nand U9051 (N_9051,N_8836,N_8854);
nor U9052 (N_9052,N_8867,N_8908);
or U9053 (N_9053,N_8940,N_8819);
xnor U9054 (N_9054,N_8915,N_8878);
or U9055 (N_9055,N_8941,N_8909);
and U9056 (N_9056,N_8831,N_8966);
and U9057 (N_9057,N_8849,N_8993);
nor U9058 (N_9058,N_8834,N_8883);
nand U9059 (N_9059,N_8943,N_8982);
or U9060 (N_9060,N_8890,N_8931);
and U9061 (N_9061,N_8811,N_8967);
nand U9062 (N_9062,N_8996,N_8875);
or U9063 (N_9063,N_8803,N_8928);
and U9064 (N_9064,N_8873,N_8851);
or U9065 (N_9065,N_8945,N_8830);
or U9066 (N_9066,N_8863,N_8903);
nand U9067 (N_9067,N_8999,N_8829);
nor U9068 (N_9068,N_8937,N_8919);
nand U9069 (N_9069,N_8905,N_8814);
or U9070 (N_9070,N_8933,N_8879);
nand U9071 (N_9071,N_8880,N_8934);
nand U9072 (N_9072,N_8932,N_8876);
nor U9073 (N_9073,N_8990,N_8817);
nand U9074 (N_9074,N_8860,N_8842);
nand U9075 (N_9075,N_8835,N_8847);
and U9076 (N_9076,N_8806,N_8888);
nand U9077 (N_9077,N_8802,N_8807);
nor U9078 (N_9078,N_8859,N_8820);
or U9079 (N_9079,N_8988,N_8892);
and U9080 (N_9080,N_8917,N_8900);
nand U9081 (N_9081,N_8972,N_8871);
and U9082 (N_9082,N_8853,N_8844);
nand U9083 (N_9083,N_8946,N_8850);
or U9084 (N_9084,N_8889,N_8977);
nor U9085 (N_9085,N_8895,N_8804);
nor U9086 (N_9086,N_8865,N_8975);
or U9087 (N_9087,N_8882,N_8950);
xnor U9088 (N_9088,N_8984,N_8921);
and U9089 (N_9089,N_8952,N_8930);
and U9090 (N_9090,N_8838,N_8846);
nand U9091 (N_9091,N_8861,N_8910);
nand U9092 (N_9092,N_8825,N_8935);
nor U9093 (N_9093,N_8981,N_8939);
nor U9094 (N_9094,N_8852,N_8837);
and U9095 (N_9095,N_8896,N_8912);
nor U9096 (N_9096,N_8968,N_8877);
nand U9097 (N_9097,N_8960,N_8845);
nor U9098 (N_9098,N_8916,N_8821);
nor U9099 (N_9099,N_8991,N_8826);
nor U9100 (N_9100,N_8873,N_8905);
nand U9101 (N_9101,N_8988,N_8962);
or U9102 (N_9102,N_8862,N_8966);
or U9103 (N_9103,N_8909,N_8871);
or U9104 (N_9104,N_8822,N_8901);
nand U9105 (N_9105,N_8915,N_8966);
nand U9106 (N_9106,N_8870,N_8824);
and U9107 (N_9107,N_8906,N_8804);
or U9108 (N_9108,N_8949,N_8993);
or U9109 (N_9109,N_8903,N_8995);
nand U9110 (N_9110,N_8859,N_8826);
xor U9111 (N_9111,N_8870,N_8977);
and U9112 (N_9112,N_8972,N_8816);
nor U9113 (N_9113,N_8861,N_8814);
nand U9114 (N_9114,N_8976,N_8911);
nor U9115 (N_9115,N_8972,N_8958);
or U9116 (N_9116,N_8826,N_8802);
and U9117 (N_9117,N_8867,N_8880);
xor U9118 (N_9118,N_8875,N_8960);
nor U9119 (N_9119,N_8895,N_8914);
xnor U9120 (N_9120,N_8914,N_8890);
nor U9121 (N_9121,N_8875,N_8833);
nand U9122 (N_9122,N_8852,N_8919);
and U9123 (N_9123,N_8894,N_8942);
and U9124 (N_9124,N_8838,N_8845);
or U9125 (N_9125,N_8963,N_8863);
nor U9126 (N_9126,N_8887,N_8830);
xnor U9127 (N_9127,N_8918,N_8836);
nor U9128 (N_9128,N_8839,N_8917);
nor U9129 (N_9129,N_8872,N_8954);
and U9130 (N_9130,N_8908,N_8970);
and U9131 (N_9131,N_8929,N_8920);
and U9132 (N_9132,N_8812,N_8921);
nor U9133 (N_9133,N_8895,N_8851);
or U9134 (N_9134,N_8984,N_8829);
nand U9135 (N_9135,N_8812,N_8872);
xnor U9136 (N_9136,N_8961,N_8884);
or U9137 (N_9137,N_8896,N_8964);
xor U9138 (N_9138,N_8941,N_8998);
xor U9139 (N_9139,N_8828,N_8922);
nor U9140 (N_9140,N_8934,N_8981);
nor U9141 (N_9141,N_8871,N_8942);
nand U9142 (N_9142,N_8860,N_8806);
or U9143 (N_9143,N_8905,N_8888);
nor U9144 (N_9144,N_8803,N_8984);
and U9145 (N_9145,N_8917,N_8940);
and U9146 (N_9146,N_8950,N_8949);
nand U9147 (N_9147,N_8848,N_8961);
nand U9148 (N_9148,N_8923,N_8979);
nor U9149 (N_9149,N_8854,N_8842);
and U9150 (N_9150,N_8964,N_8959);
nor U9151 (N_9151,N_8867,N_8928);
or U9152 (N_9152,N_8950,N_8959);
or U9153 (N_9153,N_8883,N_8872);
and U9154 (N_9154,N_8828,N_8899);
and U9155 (N_9155,N_8951,N_8855);
and U9156 (N_9156,N_8976,N_8971);
xnor U9157 (N_9157,N_8980,N_8874);
nor U9158 (N_9158,N_8934,N_8936);
or U9159 (N_9159,N_8911,N_8820);
xnor U9160 (N_9160,N_8968,N_8963);
nor U9161 (N_9161,N_8943,N_8968);
nor U9162 (N_9162,N_8932,N_8913);
and U9163 (N_9163,N_8808,N_8995);
or U9164 (N_9164,N_8871,N_8931);
nand U9165 (N_9165,N_8987,N_8983);
nor U9166 (N_9166,N_8972,N_8979);
nand U9167 (N_9167,N_8848,N_8959);
xor U9168 (N_9168,N_8937,N_8832);
nand U9169 (N_9169,N_8955,N_8812);
or U9170 (N_9170,N_8990,N_8865);
nor U9171 (N_9171,N_8921,N_8803);
and U9172 (N_9172,N_8870,N_8862);
nor U9173 (N_9173,N_8937,N_8877);
nand U9174 (N_9174,N_8939,N_8867);
and U9175 (N_9175,N_8881,N_8915);
nor U9176 (N_9176,N_8919,N_8891);
and U9177 (N_9177,N_8802,N_8981);
nand U9178 (N_9178,N_8968,N_8813);
or U9179 (N_9179,N_8904,N_8920);
nor U9180 (N_9180,N_8840,N_8853);
or U9181 (N_9181,N_8901,N_8938);
nor U9182 (N_9182,N_8803,N_8969);
and U9183 (N_9183,N_8835,N_8974);
nor U9184 (N_9184,N_8867,N_8931);
and U9185 (N_9185,N_8936,N_8890);
or U9186 (N_9186,N_8807,N_8811);
nor U9187 (N_9187,N_8900,N_8940);
nor U9188 (N_9188,N_8975,N_8888);
nor U9189 (N_9189,N_8997,N_8949);
or U9190 (N_9190,N_8913,N_8857);
or U9191 (N_9191,N_8803,N_8922);
nor U9192 (N_9192,N_8969,N_8819);
or U9193 (N_9193,N_8889,N_8802);
nand U9194 (N_9194,N_8829,N_8806);
or U9195 (N_9195,N_8813,N_8822);
and U9196 (N_9196,N_8998,N_8914);
nand U9197 (N_9197,N_8920,N_8996);
nor U9198 (N_9198,N_8820,N_8893);
nand U9199 (N_9199,N_8854,N_8999);
nor U9200 (N_9200,N_9173,N_9105);
nor U9201 (N_9201,N_9057,N_9033);
nand U9202 (N_9202,N_9129,N_9083);
and U9203 (N_9203,N_9110,N_9195);
nand U9204 (N_9204,N_9066,N_9069);
nand U9205 (N_9205,N_9157,N_9048);
nand U9206 (N_9206,N_9043,N_9046);
xor U9207 (N_9207,N_9140,N_9184);
nor U9208 (N_9208,N_9049,N_9145);
xnor U9209 (N_9209,N_9005,N_9161);
nor U9210 (N_9210,N_9159,N_9116);
nor U9211 (N_9211,N_9016,N_9019);
and U9212 (N_9212,N_9119,N_9179);
and U9213 (N_9213,N_9030,N_9064);
xor U9214 (N_9214,N_9170,N_9176);
nor U9215 (N_9215,N_9172,N_9109);
and U9216 (N_9216,N_9012,N_9120);
nor U9217 (N_9217,N_9091,N_9090);
and U9218 (N_9218,N_9141,N_9187);
nor U9219 (N_9219,N_9058,N_9183);
nor U9220 (N_9220,N_9154,N_9039);
nand U9221 (N_9221,N_9135,N_9181);
nand U9222 (N_9222,N_9011,N_9113);
and U9223 (N_9223,N_9032,N_9193);
and U9224 (N_9224,N_9151,N_9102);
nand U9225 (N_9225,N_9054,N_9103);
nand U9226 (N_9226,N_9162,N_9021);
nor U9227 (N_9227,N_9188,N_9168);
or U9228 (N_9228,N_9017,N_9067);
and U9229 (N_9229,N_9084,N_9128);
nand U9230 (N_9230,N_9079,N_9190);
nor U9231 (N_9231,N_9106,N_9166);
nand U9232 (N_9232,N_9020,N_9078);
and U9233 (N_9233,N_9003,N_9042);
or U9234 (N_9234,N_9036,N_9028);
nand U9235 (N_9235,N_9185,N_9112);
or U9236 (N_9236,N_9004,N_9155);
nor U9237 (N_9237,N_9026,N_9062);
xor U9238 (N_9238,N_9010,N_9063);
xnor U9239 (N_9239,N_9094,N_9077);
nor U9240 (N_9240,N_9137,N_9055);
nand U9241 (N_9241,N_9070,N_9056);
nor U9242 (N_9242,N_9158,N_9038);
or U9243 (N_9243,N_9051,N_9047);
or U9244 (N_9244,N_9175,N_9198);
or U9245 (N_9245,N_9177,N_9008);
xnor U9246 (N_9246,N_9174,N_9138);
nor U9247 (N_9247,N_9147,N_9099);
or U9248 (N_9248,N_9018,N_9013);
nor U9249 (N_9249,N_9134,N_9133);
and U9250 (N_9250,N_9027,N_9023);
or U9251 (N_9251,N_9006,N_9098);
nor U9252 (N_9252,N_9178,N_9148);
nand U9253 (N_9253,N_9061,N_9100);
nand U9254 (N_9254,N_9059,N_9071);
and U9255 (N_9255,N_9080,N_9089);
xor U9256 (N_9256,N_9196,N_9085);
or U9257 (N_9257,N_9031,N_9040);
nand U9258 (N_9258,N_9081,N_9144);
nor U9259 (N_9259,N_9076,N_9192);
or U9260 (N_9260,N_9186,N_9024);
nand U9261 (N_9261,N_9035,N_9104);
or U9262 (N_9262,N_9045,N_9093);
nor U9263 (N_9263,N_9164,N_9136);
or U9264 (N_9264,N_9044,N_9111);
xnor U9265 (N_9265,N_9169,N_9115);
nand U9266 (N_9266,N_9180,N_9082);
or U9267 (N_9267,N_9124,N_9163);
nand U9268 (N_9268,N_9156,N_9125);
nand U9269 (N_9269,N_9101,N_9117);
xor U9270 (N_9270,N_9015,N_9122);
and U9271 (N_9271,N_9139,N_9052);
xnor U9272 (N_9272,N_9167,N_9199);
or U9273 (N_9273,N_9060,N_9171);
nand U9274 (N_9274,N_9118,N_9143);
or U9275 (N_9275,N_9150,N_9107);
nor U9276 (N_9276,N_9022,N_9127);
nor U9277 (N_9277,N_9041,N_9000);
nand U9278 (N_9278,N_9123,N_9108);
xor U9279 (N_9279,N_9087,N_9007);
nand U9280 (N_9280,N_9121,N_9130);
nand U9281 (N_9281,N_9037,N_9197);
xnor U9282 (N_9282,N_9034,N_9096);
nor U9283 (N_9283,N_9050,N_9025);
and U9284 (N_9284,N_9191,N_9068);
nand U9285 (N_9285,N_9074,N_9002);
and U9286 (N_9286,N_9088,N_9053);
nor U9287 (N_9287,N_9075,N_9029);
nand U9288 (N_9288,N_9001,N_9160);
nand U9289 (N_9289,N_9065,N_9009);
or U9290 (N_9290,N_9132,N_9073);
nand U9291 (N_9291,N_9182,N_9131);
or U9292 (N_9292,N_9152,N_9194);
nand U9293 (N_9293,N_9142,N_9189);
nor U9294 (N_9294,N_9149,N_9014);
xnor U9295 (N_9295,N_9097,N_9126);
nand U9296 (N_9296,N_9165,N_9072);
nor U9297 (N_9297,N_9092,N_9095);
nor U9298 (N_9298,N_9114,N_9146);
and U9299 (N_9299,N_9153,N_9086);
nor U9300 (N_9300,N_9121,N_9106);
nand U9301 (N_9301,N_9060,N_9019);
nand U9302 (N_9302,N_9001,N_9132);
nor U9303 (N_9303,N_9176,N_9080);
and U9304 (N_9304,N_9136,N_9181);
nand U9305 (N_9305,N_9003,N_9154);
nor U9306 (N_9306,N_9142,N_9144);
or U9307 (N_9307,N_9122,N_9157);
or U9308 (N_9308,N_9052,N_9025);
and U9309 (N_9309,N_9020,N_9177);
or U9310 (N_9310,N_9075,N_9084);
nand U9311 (N_9311,N_9017,N_9126);
or U9312 (N_9312,N_9101,N_9062);
and U9313 (N_9313,N_9181,N_9006);
or U9314 (N_9314,N_9001,N_9090);
and U9315 (N_9315,N_9121,N_9070);
and U9316 (N_9316,N_9109,N_9021);
and U9317 (N_9317,N_9090,N_9003);
nor U9318 (N_9318,N_9131,N_9195);
or U9319 (N_9319,N_9045,N_9160);
and U9320 (N_9320,N_9140,N_9072);
nor U9321 (N_9321,N_9152,N_9132);
or U9322 (N_9322,N_9190,N_9088);
or U9323 (N_9323,N_9172,N_9123);
nand U9324 (N_9324,N_9030,N_9097);
and U9325 (N_9325,N_9046,N_9020);
and U9326 (N_9326,N_9028,N_9120);
or U9327 (N_9327,N_9011,N_9009);
and U9328 (N_9328,N_9081,N_9061);
or U9329 (N_9329,N_9026,N_9141);
nor U9330 (N_9330,N_9187,N_9038);
and U9331 (N_9331,N_9110,N_9147);
nor U9332 (N_9332,N_9030,N_9093);
or U9333 (N_9333,N_9165,N_9177);
and U9334 (N_9334,N_9082,N_9019);
xnor U9335 (N_9335,N_9097,N_9123);
and U9336 (N_9336,N_9133,N_9087);
or U9337 (N_9337,N_9123,N_9022);
and U9338 (N_9338,N_9128,N_9199);
or U9339 (N_9339,N_9050,N_9158);
nand U9340 (N_9340,N_9092,N_9002);
nor U9341 (N_9341,N_9199,N_9005);
or U9342 (N_9342,N_9153,N_9176);
and U9343 (N_9343,N_9138,N_9153);
xor U9344 (N_9344,N_9115,N_9085);
nor U9345 (N_9345,N_9151,N_9048);
nand U9346 (N_9346,N_9068,N_9064);
and U9347 (N_9347,N_9140,N_9198);
xor U9348 (N_9348,N_9150,N_9093);
nor U9349 (N_9349,N_9179,N_9045);
and U9350 (N_9350,N_9156,N_9121);
and U9351 (N_9351,N_9018,N_9131);
nor U9352 (N_9352,N_9118,N_9096);
or U9353 (N_9353,N_9014,N_9106);
xor U9354 (N_9354,N_9048,N_9046);
nor U9355 (N_9355,N_9077,N_9048);
and U9356 (N_9356,N_9065,N_9170);
and U9357 (N_9357,N_9084,N_9189);
nor U9358 (N_9358,N_9014,N_9103);
and U9359 (N_9359,N_9189,N_9065);
or U9360 (N_9360,N_9127,N_9053);
nand U9361 (N_9361,N_9078,N_9039);
or U9362 (N_9362,N_9126,N_9100);
nand U9363 (N_9363,N_9066,N_9056);
and U9364 (N_9364,N_9020,N_9080);
nand U9365 (N_9365,N_9192,N_9085);
xor U9366 (N_9366,N_9072,N_9062);
nor U9367 (N_9367,N_9102,N_9121);
nand U9368 (N_9368,N_9123,N_9149);
nand U9369 (N_9369,N_9044,N_9014);
nor U9370 (N_9370,N_9045,N_9058);
or U9371 (N_9371,N_9126,N_9115);
nor U9372 (N_9372,N_9087,N_9126);
nor U9373 (N_9373,N_9062,N_9155);
xor U9374 (N_9374,N_9103,N_9077);
nor U9375 (N_9375,N_9065,N_9031);
and U9376 (N_9376,N_9027,N_9109);
and U9377 (N_9377,N_9031,N_9199);
xor U9378 (N_9378,N_9035,N_9064);
and U9379 (N_9379,N_9066,N_9110);
and U9380 (N_9380,N_9049,N_9188);
or U9381 (N_9381,N_9019,N_9161);
xor U9382 (N_9382,N_9022,N_9162);
nand U9383 (N_9383,N_9087,N_9111);
and U9384 (N_9384,N_9197,N_9120);
or U9385 (N_9385,N_9047,N_9003);
or U9386 (N_9386,N_9077,N_9186);
nand U9387 (N_9387,N_9090,N_9156);
nand U9388 (N_9388,N_9120,N_9092);
or U9389 (N_9389,N_9078,N_9195);
xor U9390 (N_9390,N_9161,N_9108);
nor U9391 (N_9391,N_9078,N_9140);
nand U9392 (N_9392,N_9137,N_9047);
xor U9393 (N_9393,N_9161,N_9079);
xnor U9394 (N_9394,N_9060,N_9035);
or U9395 (N_9395,N_9143,N_9117);
nor U9396 (N_9396,N_9037,N_9083);
nand U9397 (N_9397,N_9053,N_9141);
and U9398 (N_9398,N_9041,N_9031);
nand U9399 (N_9399,N_9062,N_9099);
nand U9400 (N_9400,N_9301,N_9367);
nand U9401 (N_9401,N_9315,N_9283);
nand U9402 (N_9402,N_9238,N_9365);
nand U9403 (N_9403,N_9320,N_9304);
and U9404 (N_9404,N_9252,N_9279);
nand U9405 (N_9405,N_9324,N_9352);
nor U9406 (N_9406,N_9363,N_9355);
nand U9407 (N_9407,N_9384,N_9319);
and U9408 (N_9408,N_9234,N_9359);
or U9409 (N_9409,N_9233,N_9397);
nor U9410 (N_9410,N_9378,N_9331);
nand U9411 (N_9411,N_9313,N_9248);
nor U9412 (N_9412,N_9326,N_9208);
or U9413 (N_9413,N_9338,N_9321);
nor U9414 (N_9414,N_9202,N_9206);
nor U9415 (N_9415,N_9366,N_9287);
and U9416 (N_9416,N_9204,N_9329);
xor U9417 (N_9417,N_9292,N_9229);
or U9418 (N_9418,N_9336,N_9246);
xor U9419 (N_9419,N_9368,N_9341);
and U9420 (N_9420,N_9225,N_9340);
xor U9421 (N_9421,N_9333,N_9286);
nor U9422 (N_9422,N_9226,N_9253);
nand U9423 (N_9423,N_9388,N_9269);
nand U9424 (N_9424,N_9330,N_9349);
or U9425 (N_9425,N_9380,N_9371);
xor U9426 (N_9426,N_9240,N_9219);
or U9427 (N_9427,N_9342,N_9213);
and U9428 (N_9428,N_9249,N_9255);
nand U9429 (N_9429,N_9360,N_9375);
nor U9430 (N_9430,N_9237,N_9241);
nor U9431 (N_9431,N_9227,N_9305);
nand U9432 (N_9432,N_9356,N_9210);
nand U9433 (N_9433,N_9242,N_9201);
nor U9434 (N_9434,N_9303,N_9372);
or U9435 (N_9435,N_9357,N_9258);
nand U9436 (N_9436,N_9231,N_9285);
nand U9437 (N_9437,N_9275,N_9256);
or U9438 (N_9438,N_9350,N_9362);
or U9439 (N_9439,N_9318,N_9392);
and U9440 (N_9440,N_9207,N_9254);
and U9441 (N_9441,N_9327,N_9383);
and U9442 (N_9442,N_9280,N_9284);
nand U9443 (N_9443,N_9312,N_9245);
nand U9444 (N_9444,N_9354,N_9224);
or U9445 (N_9445,N_9325,N_9391);
or U9446 (N_9446,N_9339,N_9369);
xnor U9447 (N_9447,N_9334,N_9209);
and U9448 (N_9448,N_9257,N_9273);
and U9449 (N_9449,N_9214,N_9260);
and U9450 (N_9450,N_9299,N_9200);
nor U9451 (N_9451,N_9382,N_9217);
nand U9452 (N_9452,N_9348,N_9394);
nand U9453 (N_9453,N_9259,N_9344);
and U9454 (N_9454,N_9374,N_9212);
xnor U9455 (N_9455,N_9393,N_9297);
nor U9456 (N_9456,N_9310,N_9223);
nor U9457 (N_9457,N_9220,N_9370);
or U9458 (N_9458,N_9239,N_9203);
nand U9459 (N_9459,N_9262,N_9236);
nor U9460 (N_9460,N_9265,N_9271);
nor U9461 (N_9461,N_9337,N_9300);
nor U9462 (N_9462,N_9316,N_9261);
and U9463 (N_9463,N_9345,N_9291);
xor U9464 (N_9464,N_9381,N_9263);
nand U9465 (N_9465,N_9364,N_9386);
and U9466 (N_9466,N_9222,N_9218);
nand U9467 (N_9467,N_9216,N_9288);
or U9468 (N_9468,N_9390,N_9289);
or U9469 (N_9469,N_9347,N_9235);
nor U9470 (N_9470,N_9244,N_9351);
nor U9471 (N_9471,N_9295,N_9395);
or U9472 (N_9472,N_9294,N_9398);
or U9473 (N_9473,N_9266,N_9290);
and U9474 (N_9474,N_9268,N_9247);
nand U9475 (N_9475,N_9278,N_9215);
or U9476 (N_9476,N_9232,N_9298);
nand U9477 (N_9477,N_9373,N_9385);
or U9478 (N_9478,N_9267,N_9322);
nor U9479 (N_9479,N_9387,N_9270);
nor U9480 (N_9480,N_9361,N_9250);
nand U9481 (N_9481,N_9272,N_9302);
and U9482 (N_9482,N_9281,N_9307);
xor U9483 (N_9483,N_9251,N_9205);
and U9484 (N_9484,N_9376,N_9308);
nand U9485 (N_9485,N_9309,N_9358);
nor U9486 (N_9486,N_9379,N_9211);
nor U9487 (N_9487,N_9323,N_9296);
nor U9488 (N_9488,N_9314,N_9277);
nand U9489 (N_9489,N_9230,N_9306);
nor U9490 (N_9490,N_9276,N_9264);
nor U9491 (N_9491,N_9311,N_9346);
xor U9492 (N_9492,N_9335,N_9377);
nor U9493 (N_9493,N_9243,N_9396);
xor U9494 (N_9494,N_9221,N_9343);
xnor U9495 (N_9495,N_9389,N_9293);
xnor U9496 (N_9496,N_9328,N_9399);
nor U9497 (N_9497,N_9282,N_9317);
and U9498 (N_9498,N_9274,N_9228);
or U9499 (N_9499,N_9353,N_9332);
nand U9500 (N_9500,N_9267,N_9365);
and U9501 (N_9501,N_9307,N_9379);
nor U9502 (N_9502,N_9228,N_9303);
and U9503 (N_9503,N_9231,N_9365);
nand U9504 (N_9504,N_9252,N_9223);
and U9505 (N_9505,N_9332,N_9394);
or U9506 (N_9506,N_9217,N_9290);
nand U9507 (N_9507,N_9390,N_9272);
nand U9508 (N_9508,N_9348,N_9266);
or U9509 (N_9509,N_9342,N_9327);
nand U9510 (N_9510,N_9205,N_9398);
or U9511 (N_9511,N_9343,N_9392);
and U9512 (N_9512,N_9298,N_9283);
or U9513 (N_9513,N_9287,N_9321);
or U9514 (N_9514,N_9254,N_9336);
nand U9515 (N_9515,N_9228,N_9273);
and U9516 (N_9516,N_9351,N_9350);
and U9517 (N_9517,N_9265,N_9313);
or U9518 (N_9518,N_9332,N_9312);
or U9519 (N_9519,N_9369,N_9351);
and U9520 (N_9520,N_9347,N_9274);
and U9521 (N_9521,N_9285,N_9240);
nor U9522 (N_9522,N_9363,N_9274);
nand U9523 (N_9523,N_9336,N_9259);
nor U9524 (N_9524,N_9286,N_9335);
or U9525 (N_9525,N_9235,N_9244);
nand U9526 (N_9526,N_9293,N_9364);
nand U9527 (N_9527,N_9306,N_9382);
and U9528 (N_9528,N_9290,N_9397);
or U9529 (N_9529,N_9250,N_9233);
and U9530 (N_9530,N_9372,N_9272);
xor U9531 (N_9531,N_9217,N_9201);
nand U9532 (N_9532,N_9225,N_9344);
and U9533 (N_9533,N_9249,N_9354);
nor U9534 (N_9534,N_9282,N_9337);
nor U9535 (N_9535,N_9362,N_9319);
and U9536 (N_9536,N_9295,N_9361);
nand U9537 (N_9537,N_9277,N_9238);
nand U9538 (N_9538,N_9225,N_9206);
or U9539 (N_9539,N_9208,N_9372);
or U9540 (N_9540,N_9339,N_9273);
or U9541 (N_9541,N_9245,N_9335);
or U9542 (N_9542,N_9363,N_9323);
nor U9543 (N_9543,N_9294,N_9248);
and U9544 (N_9544,N_9296,N_9398);
or U9545 (N_9545,N_9324,N_9383);
and U9546 (N_9546,N_9200,N_9300);
or U9547 (N_9547,N_9286,N_9227);
and U9548 (N_9548,N_9251,N_9347);
or U9549 (N_9549,N_9258,N_9312);
nor U9550 (N_9550,N_9350,N_9200);
and U9551 (N_9551,N_9276,N_9356);
nor U9552 (N_9552,N_9371,N_9276);
nor U9553 (N_9553,N_9323,N_9277);
nand U9554 (N_9554,N_9395,N_9214);
and U9555 (N_9555,N_9264,N_9354);
nor U9556 (N_9556,N_9228,N_9349);
nor U9557 (N_9557,N_9367,N_9256);
and U9558 (N_9558,N_9268,N_9358);
and U9559 (N_9559,N_9340,N_9211);
nor U9560 (N_9560,N_9310,N_9325);
and U9561 (N_9561,N_9300,N_9228);
and U9562 (N_9562,N_9331,N_9354);
nand U9563 (N_9563,N_9206,N_9238);
and U9564 (N_9564,N_9299,N_9393);
nor U9565 (N_9565,N_9298,N_9251);
and U9566 (N_9566,N_9363,N_9240);
or U9567 (N_9567,N_9373,N_9275);
xor U9568 (N_9568,N_9247,N_9287);
and U9569 (N_9569,N_9374,N_9341);
or U9570 (N_9570,N_9397,N_9243);
or U9571 (N_9571,N_9388,N_9241);
nand U9572 (N_9572,N_9233,N_9276);
and U9573 (N_9573,N_9202,N_9222);
or U9574 (N_9574,N_9210,N_9335);
or U9575 (N_9575,N_9208,N_9252);
nor U9576 (N_9576,N_9202,N_9361);
or U9577 (N_9577,N_9355,N_9342);
nand U9578 (N_9578,N_9276,N_9208);
or U9579 (N_9579,N_9259,N_9390);
and U9580 (N_9580,N_9309,N_9218);
xor U9581 (N_9581,N_9240,N_9394);
nor U9582 (N_9582,N_9257,N_9232);
or U9583 (N_9583,N_9233,N_9268);
xnor U9584 (N_9584,N_9261,N_9242);
nor U9585 (N_9585,N_9320,N_9201);
or U9586 (N_9586,N_9261,N_9324);
nor U9587 (N_9587,N_9331,N_9232);
nor U9588 (N_9588,N_9382,N_9374);
nor U9589 (N_9589,N_9287,N_9259);
and U9590 (N_9590,N_9270,N_9279);
and U9591 (N_9591,N_9272,N_9219);
nor U9592 (N_9592,N_9399,N_9381);
or U9593 (N_9593,N_9291,N_9305);
nor U9594 (N_9594,N_9346,N_9204);
nand U9595 (N_9595,N_9234,N_9209);
or U9596 (N_9596,N_9243,N_9216);
xor U9597 (N_9597,N_9234,N_9328);
xor U9598 (N_9598,N_9334,N_9363);
nor U9599 (N_9599,N_9263,N_9385);
or U9600 (N_9600,N_9511,N_9438);
nor U9601 (N_9601,N_9460,N_9579);
nor U9602 (N_9602,N_9561,N_9531);
nor U9603 (N_9603,N_9482,N_9426);
or U9604 (N_9604,N_9559,N_9530);
nand U9605 (N_9605,N_9543,N_9504);
xor U9606 (N_9606,N_9442,N_9501);
or U9607 (N_9607,N_9515,N_9425);
nor U9608 (N_9608,N_9469,N_9465);
or U9609 (N_9609,N_9509,N_9521);
xor U9610 (N_9610,N_9450,N_9410);
xnor U9611 (N_9611,N_9587,N_9514);
and U9612 (N_9612,N_9503,N_9599);
xnor U9613 (N_9613,N_9536,N_9506);
nor U9614 (N_9614,N_9516,N_9592);
and U9615 (N_9615,N_9492,N_9479);
nand U9616 (N_9616,N_9427,N_9443);
nor U9617 (N_9617,N_9597,N_9537);
nor U9618 (N_9618,N_9490,N_9459);
or U9619 (N_9619,N_9462,N_9452);
nand U9620 (N_9620,N_9575,N_9583);
or U9621 (N_9621,N_9508,N_9549);
or U9622 (N_9622,N_9567,N_9413);
xnor U9623 (N_9623,N_9447,N_9428);
nand U9624 (N_9624,N_9499,N_9591);
and U9625 (N_9625,N_9554,N_9580);
and U9626 (N_9626,N_9418,N_9403);
or U9627 (N_9627,N_9439,N_9457);
and U9628 (N_9628,N_9494,N_9540);
nor U9629 (N_9629,N_9491,N_9526);
nor U9630 (N_9630,N_9474,N_9545);
xor U9631 (N_9631,N_9585,N_9449);
and U9632 (N_9632,N_9404,N_9538);
nor U9633 (N_9633,N_9560,N_9402);
xnor U9634 (N_9634,N_9412,N_9434);
nor U9635 (N_9635,N_9467,N_9433);
or U9636 (N_9636,N_9502,N_9420);
nand U9637 (N_9637,N_9497,N_9400);
xnor U9638 (N_9638,N_9470,N_9568);
and U9639 (N_9639,N_9424,N_9436);
nor U9640 (N_9640,N_9464,N_9571);
nand U9641 (N_9641,N_9440,N_9444);
nor U9642 (N_9642,N_9417,N_9488);
nor U9643 (N_9643,N_9471,N_9525);
nor U9644 (N_9644,N_9505,N_9573);
or U9645 (N_9645,N_9586,N_9437);
nor U9646 (N_9646,N_9487,N_9510);
xor U9647 (N_9647,N_9553,N_9563);
xnor U9648 (N_9648,N_9546,N_9495);
or U9649 (N_9649,N_9408,N_9558);
or U9650 (N_9650,N_9445,N_9409);
nor U9651 (N_9651,N_9422,N_9527);
or U9652 (N_9652,N_9524,N_9411);
and U9653 (N_9653,N_9486,N_9578);
and U9654 (N_9654,N_9533,N_9528);
and U9655 (N_9655,N_9574,N_9453);
or U9656 (N_9656,N_9589,N_9565);
nor U9657 (N_9657,N_9596,N_9414);
xnor U9658 (N_9658,N_9522,N_9430);
nand U9659 (N_9659,N_9555,N_9466);
nor U9660 (N_9660,N_9419,N_9455);
nor U9661 (N_9661,N_9518,N_9406);
nor U9662 (N_9662,N_9519,N_9432);
xnor U9663 (N_9663,N_9456,N_9421);
or U9664 (N_9664,N_9542,N_9415);
nor U9665 (N_9665,N_9507,N_9454);
nor U9666 (N_9666,N_9562,N_9547);
nand U9667 (N_9667,N_9534,N_9557);
nand U9668 (N_9668,N_9463,N_9590);
nor U9669 (N_9669,N_9513,N_9481);
nor U9670 (N_9670,N_9480,N_9581);
nor U9671 (N_9671,N_9588,N_9435);
or U9672 (N_9672,N_9498,N_9539);
or U9673 (N_9673,N_9556,N_9576);
and U9674 (N_9674,N_9489,N_9551);
or U9675 (N_9675,N_9484,N_9569);
nor U9676 (N_9676,N_9401,N_9512);
nor U9677 (N_9677,N_9520,N_9416);
xor U9678 (N_9678,N_9458,N_9478);
nor U9679 (N_9679,N_9407,N_9582);
nor U9680 (N_9680,N_9441,N_9570);
nor U9681 (N_9681,N_9451,N_9532);
xnor U9682 (N_9682,N_9461,N_9493);
and U9683 (N_9683,N_9594,N_9598);
nor U9684 (N_9684,N_9548,N_9593);
nor U9685 (N_9685,N_9552,N_9544);
or U9686 (N_9686,N_9550,N_9529);
and U9687 (N_9687,N_9496,N_9473);
nor U9688 (N_9688,N_9483,N_9446);
nand U9689 (N_9689,N_9429,N_9595);
and U9690 (N_9690,N_9472,N_9485);
nand U9691 (N_9691,N_9541,N_9517);
and U9692 (N_9692,N_9423,N_9431);
nand U9693 (N_9693,N_9566,N_9475);
nand U9694 (N_9694,N_9584,N_9523);
and U9695 (N_9695,N_9476,N_9564);
and U9696 (N_9696,N_9448,N_9535);
nand U9697 (N_9697,N_9468,N_9577);
nand U9698 (N_9698,N_9405,N_9572);
nor U9699 (N_9699,N_9500,N_9477);
and U9700 (N_9700,N_9552,N_9490);
and U9701 (N_9701,N_9458,N_9520);
nand U9702 (N_9702,N_9586,N_9549);
and U9703 (N_9703,N_9414,N_9566);
or U9704 (N_9704,N_9563,N_9433);
nand U9705 (N_9705,N_9451,N_9530);
xnor U9706 (N_9706,N_9587,N_9456);
nand U9707 (N_9707,N_9577,N_9574);
or U9708 (N_9708,N_9492,N_9524);
nor U9709 (N_9709,N_9465,N_9429);
nor U9710 (N_9710,N_9592,N_9422);
and U9711 (N_9711,N_9510,N_9540);
nand U9712 (N_9712,N_9580,N_9548);
or U9713 (N_9713,N_9479,N_9569);
and U9714 (N_9714,N_9422,N_9499);
and U9715 (N_9715,N_9426,N_9524);
or U9716 (N_9716,N_9574,N_9499);
nand U9717 (N_9717,N_9524,N_9456);
nor U9718 (N_9718,N_9552,N_9455);
nor U9719 (N_9719,N_9407,N_9410);
and U9720 (N_9720,N_9422,N_9548);
nor U9721 (N_9721,N_9467,N_9457);
nand U9722 (N_9722,N_9499,N_9496);
and U9723 (N_9723,N_9439,N_9553);
or U9724 (N_9724,N_9426,N_9508);
and U9725 (N_9725,N_9450,N_9480);
xor U9726 (N_9726,N_9403,N_9566);
and U9727 (N_9727,N_9475,N_9524);
and U9728 (N_9728,N_9404,N_9456);
nor U9729 (N_9729,N_9576,N_9502);
xor U9730 (N_9730,N_9521,N_9412);
nand U9731 (N_9731,N_9514,N_9491);
nor U9732 (N_9732,N_9458,N_9416);
nor U9733 (N_9733,N_9505,N_9590);
nor U9734 (N_9734,N_9402,N_9435);
nand U9735 (N_9735,N_9551,N_9567);
and U9736 (N_9736,N_9591,N_9573);
and U9737 (N_9737,N_9403,N_9544);
nor U9738 (N_9738,N_9472,N_9548);
nand U9739 (N_9739,N_9477,N_9490);
nor U9740 (N_9740,N_9499,N_9462);
nand U9741 (N_9741,N_9420,N_9509);
nor U9742 (N_9742,N_9464,N_9401);
and U9743 (N_9743,N_9415,N_9512);
and U9744 (N_9744,N_9580,N_9413);
nand U9745 (N_9745,N_9461,N_9568);
nor U9746 (N_9746,N_9492,N_9438);
and U9747 (N_9747,N_9574,N_9518);
xnor U9748 (N_9748,N_9506,N_9483);
nand U9749 (N_9749,N_9432,N_9425);
xor U9750 (N_9750,N_9402,N_9554);
nand U9751 (N_9751,N_9465,N_9554);
or U9752 (N_9752,N_9454,N_9477);
nor U9753 (N_9753,N_9437,N_9524);
nor U9754 (N_9754,N_9451,N_9573);
nor U9755 (N_9755,N_9433,N_9590);
and U9756 (N_9756,N_9469,N_9433);
nand U9757 (N_9757,N_9472,N_9584);
nand U9758 (N_9758,N_9449,N_9454);
nand U9759 (N_9759,N_9537,N_9573);
xnor U9760 (N_9760,N_9463,N_9414);
or U9761 (N_9761,N_9416,N_9516);
or U9762 (N_9762,N_9571,N_9587);
and U9763 (N_9763,N_9430,N_9461);
and U9764 (N_9764,N_9417,N_9411);
nand U9765 (N_9765,N_9544,N_9535);
nor U9766 (N_9766,N_9428,N_9421);
nand U9767 (N_9767,N_9442,N_9553);
and U9768 (N_9768,N_9439,N_9568);
and U9769 (N_9769,N_9595,N_9541);
or U9770 (N_9770,N_9475,N_9541);
nand U9771 (N_9771,N_9475,N_9593);
xor U9772 (N_9772,N_9595,N_9590);
or U9773 (N_9773,N_9591,N_9538);
nand U9774 (N_9774,N_9537,N_9546);
and U9775 (N_9775,N_9405,N_9433);
nor U9776 (N_9776,N_9553,N_9437);
nand U9777 (N_9777,N_9462,N_9423);
and U9778 (N_9778,N_9521,N_9458);
or U9779 (N_9779,N_9433,N_9448);
or U9780 (N_9780,N_9586,N_9409);
xnor U9781 (N_9781,N_9438,N_9486);
or U9782 (N_9782,N_9503,N_9431);
nand U9783 (N_9783,N_9578,N_9520);
nor U9784 (N_9784,N_9563,N_9497);
or U9785 (N_9785,N_9415,N_9515);
nand U9786 (N_9786,N_9418,N_9587);
xor U9787 (N_9787,N_9537,N_9443);
nor U9788 (N_9788,N_9561,N_9414);
nand U9789 (N_9789,N_9577,N_9446);
nor U9790 (N_9790,N_9406,N_9555);
or U9791 (N_9791,N_9406,N_9571);
nor U9792 (N_9792,N_9547,N_9569);
nand U9793 (N_9793,N_9409,N_9530);
nand U9794 (N_9794,N_9467,N_9422);
and U9795 (N_9795,N_9576,N_9471);
xnor U9796 (N_9796,N_9503,N_9575);
or U9797 (N_9797,N_9472,N_9413);
or U9798 (N_9798,N_9472,N_9503);
or U9799 (N_9799,N_9428,N_9468);
or U9800 (N_9800,N_9627,N_9639);
and U9801 (N_9801,N_9794,N_9604);
nand U9802 (N_9802,N_9697,N_9773);
or U9803 (N_9803,N_9788,N_9700);
and U9804 (N_9804,N_9710,N_9612);
nand U9805 (N_9805,N_9667,N_9779);
or U9806 (N_9806,N_9753,N_9719);
or U9807 (N_9807,N_9643,N_9622);
nor U9808 (N_9808,N_9621,N_9786);
and U9809 (N_9809,N_9757,N_9775);
or U9810 (N_9810,N_9668,N_9664);
or U9811 (N_9811,N_9691,N_9646);
and U9812 (N_9812,N_9632,N_9698);
or U9813 (N_9813,N_9699,N_9688);
nor U9814 (N_9814,N_9704,N_9693);
and U9815 (N_9815,N_9716,N_9672);
nand U9816 (N_9816,N_9785,N_9746);
and U9817 (N_9817,N_9625,N_9745);
xor U9818 (N_9818,N_9790,N_9606);
and U9819 (N_9819,N_9791,N_9732);
nand U9820 (N_9820,N_9663,N_9651);
nand U9821 (N_9821,N_9647,N_9631);
nand U9822 (N_9822,N_9726,N_9692);
and U9823 (N_9823,N_9735,N_9637);
or U9824 (N_9824,N_9649,N_9644);
or U9825 (N_9825,N_9723,N_9706);
and U9826 (N_9826,N_9702,N_9680);
or U9827 (N_9827,N_9733,N_9736);
nor U9828 (N_9828,N_9721,N_9641);
and U9829 (N_9829,N_9707,N_9768);
and U9830 (N_9830,N_9728,N_9634);
and U9831 (N_9831,N_9795,N_9690);
nor U9832 (N_9832,N_9755,N_9626);
or U9833 (N_9833,N_9661,N_9769);
or U9834 (N_9834,N_9781,N_9765);
xnor U9835 (N_9835,N_9694,N_9615);
nor U9836 (N_9836,N_9659,N_9764);
nor U9837 (N_9837,N_9751,N_9756);
or U9838 (N_9838,N_9720,N_9616);
nor U9839 (N_9839,N_9743,N_9636);
and U9840 (N_9840,N_9617,N_9683);
and U9841 (N_9841,N_9684,N_9611);
and U9842 (N_9842,N_9608,N_9766);
and U9843 (N_9843,N_9650,N_9605);
nand U9844 (N_9844,N_9796,N_9749);
xnor U9845 (N_9845,N_9739,N_9747);
nor U9846 (N_9846,N_9703,N_9741);
or U9847 (N_9847,N_9799,N_9708);
and U9848 (N_9848,N_9673,N_9610);
and U9849 (N_9849,N_9687,N_9752);
or U9850 (N_9850,N_9714,N_9784);
or U9851 (N_9851,N_9628,N_9648);
nand U9852 (N_9852,N_9792,N_9638);
nor U9853 (N_9853,N_9725,N_9642);
nand U9854 (N_9854,N_9620,N_9653);
nor U9855 (N_9855,N_9629,N_9670);
or U9856 (N_9856,N_9624,N_9762);
or U9857 (N_9857,N_9718,N_9750);
and U9858 (N_9858,N_9686,N_9709);
and U9859 (N_9859,N_9798,N_9677);
nor U9860 (N_9860,N_9602,N_9731);
nand U9861 (N_9861,N_9685,N_9696);
or U9862 (N_9862,N_9759,N_9660);
and U9863 (N_9863,N_9609,N_9654);
nand U9864 (N_9864,N_9711,N_9678);
and U9865 (N_9865,N_9748,N_9776);
nor U9866 (N_9866,N_9763,N_9758);
xnor U9867 (N_9867,N_9774,N_9679);
or U9868 (N_9868,N_9740,N_9793);
xor U9869 (N_9869,N_9640,N_9712);
xnor U9870 (N_9870,N_9666,N_9713);
nor U9871 (N_9871,N_9630,N_9675);
nand U9872 (N_9872,N_9665,N_9652);
nand U9873 (N_9873,N_9645,N_9633);
nand U9874 (N_9874,N_9681,N_9600);
or U9875 (N_9875,N_9777,N_9744);
nor U9876 (N_9876,N_9782,N_9657);
xnor U9877 (N_9877,N_9724,N_9737);
or U9878 (N_9878,N_9730,N_9601);
nand U9879 (N_9879,N_9761,N_9674);
nand U9880 (N_9880,N_9701,N_9662);
nor U9881 (N_9881,N_9787,N_9671);
nor U9882 (N_9882,N_9780,N_9689);
and U9883 (N_9883,N_9717,N_9778);
nor U9884 (N_9884,N_9619,N_9734);
or U9885 (N_9885,N_9738,N_9655);
and U9886 (N_9886,N_9618,N_9607);
nor U9887 (N_9887,N_9658,N_9789);
and U9888 (N_9888,N_9722,N_9613);
and U9889 (N_9889,N_9705,N_9760);
and U9890 (N_9890,N_9727,N_9783);
nand U9891 (N_9891,N_9771,N_9695);
and U9892 (N_9892,N_9669,N_9656);
nor U9893 (N_9893,N_9772,N_9742);
and U9894 (N_9894,N_9676,N_9729);
xnor U9895 (N_9895,N_9770,N_9682);
or U9896 (N_9896,N_9614,N_9623);
and U9897 (N_9897,N_9635,N_9797);
nor U9898 (N_9898,N_9767,N_9603);
nand U9899 (N_9899,N_9715,N_9754);
and U9900 (N_9900,N_9799,N_9780);
or U9901 (N_9901,N_9664,N_9798);
or U9902 (N_9902,N_9604,N_9796);
or U9903 (N_9903,N_9697,N_9719);
nand U9904 (N_9904,N_9680,N_9676);
or U9905 (N_9905,N_9718,N_9652);
nand U9906 (N_9906,N_9631,N_9751);
nor U9907 (N_9907,N_9750,N_9632);
or U9908 (N_9908,N_9688,N_9698);
and U9909 (N_9909,N_9686,N_9703);
nor U9910 (N_9910,N_9710,N_9633);
or U9911 (N_9911,N_9794,N_9711);
or U9912 (N_9912,N_9681,N_9631);
nand U9913 (N_9913,N_9618,N_9685);
or U9914 (N_9914,N_9718,N_9654);
and U9915 (N_9915,N_9733,N_9750);
nand U9916 (N_9916,N_9700,N_9618);
or U9917 (N_9917,N_9678,N_9746);
nand U9918 (N_9918,N_9674,N_9751);
and U9919 (N_9919,N_9607,N_9692);
nand U9920 (N_9920,N_9632,N_9620);
and U9921 (N_9921,N_9641,N_9635);
xor U9922 (N_9922,N_9710,N_9606);
and U9923 (N_9923,N_9653,N_9797);
xor U9924 (N_9924,N_9667,N_9620);
nand U9925 (N_9925,N_9643,N_9649);
and U9926 (N_9926,N_9663,N_9699);
nand U9927 (N_9927,N_9733,N_9684);
nor U9928 (N_9928,N_9799,N_9650);
or U9929 (N_9929,N_9692,N_9790);
and U9930 (N_9930,N_9602,N_9630);
nand U9931 (N_9931,N_9618,N_9608);
or U9932 (N_9932,N_9740,N_9614);
or U9933 (N_9933,N_9633,N_9625);
and U9934 (N_9934,N_9684,N_9668);
and U9935 (N_9935,N_9645,N_9613);
or U9936 (N_9936,N_9742,N_9735);
nor U9937 (N_9937,N_9634,N_9773);
and U9938 (N_9938,N_9612,N_9633);
xnor U9939 (N_9939,N_9777,N_9646);
or U9940 (N_9940,N_9645,N_9693);
nor U9941 (N_9941,N_9784,N_9603);
and U9942 (N_9942,N_9704,N_9706);
nor U9943 (N_9943,N_9779,N_9624);
or U9944 (N_9944,N_9691,N_9649);
and U9945 (N_9945,N_9686,N_9706);
nor U9946 (N_9946,N_9694,N_9726);
or U9947 (N_9947,N_9756,N_9728);
and U9948 (N_9948,N_9719,N_9668);
nor U9949 (N_9949,N_9734,N_9661);
and U9950 (N_9950,N_9690,N_9640);
or U9951 (N_9951,N_9669,N_9744);
nand U9952 (N_9952,N_9641,N_9679);
and U9953 (N_9953,N_9776,N_9645);
and U9954 (N_9954,N_9608,N_9755);
or U9955 (N_9955,N_9738,N_9742);
or U9956 (N_9956,N_9666,N_9770);
or U9957 (N_9957,N_9713,N_9784);
xnor U9958 (N_9958,N_9747,N_9637);
or U9959 (N_9959,N_9622,N_9715);
nand U9960 (N_9960,N_9700,N_9738);
and U9961 (N_9961,N_9686,N_9662);
or U9962 (N_9962,N_9747,N_9667);
nor U9963 (N_9963,N_9745,N_9779);
and U9964 (N_9964,N_9738,N_9698);
nand U9965 (N_9965,N_9741,N_9761);
xnor U9966 (N_9966,N_9718,N_9723);
or U9967 (N_9967,N_9678,N_9608);
nor U9968 (N_9968,N_9605,N_9656);
or U9969 (N_9969,N_9611,N_9630);
nor U9970 (N_9970,N_9747,N_9632);
and U9971 (N_9971,N_9678,N_9776);
xor U9972 (N_9972,N_9758,N_9667);
nand U9973 (N_9973,N_9714,N_9663);
or U9974 (N_9974,N_9758,N_9770);
nor U9975 (N_9975,N_9725,N_9695);
nor U9976 (N_9976,N_9770,N_9689);
and U9977 (N_9977,N_9624,N_9649);
and U9978 (N_9978,N_9699,N_9680);
nand U9979 (N_9979,N_9707,N_9689);
nand U9980 (N_9980,N_9762,N_9789);
nor U9981 (N_9981,N_9614,N_9776);
nand U9982 (N_9982,N_9763,N_9699);
and U9983 (N_9983,N_9692,N_9688);
or U9984 (N_9984,N_9746,N_9791);
or U9985 (N_9985,N_9738,N_9635);
nor U9986 (N_9986,N_9690,N_9745);
nand U9987 (N_9987,N_9620,N_9742);
nand U9988 (N_9988,N_9720,N_9604);
nand U9989 (N_9989,N_9753,N_9672);
nand U9990 (N_9990,N_9691,N_9666);
nand U9991 (N_9991,N_9745,N_9766);
nor U9992 (N_9992,N_9660,N_9669);
or U9993 (N_9993,N_9659,N_9696);
nor U9994 (N_9994,N_9742,N_9653);
and U9995 (N_9995,N_9787,N_9788);
nor U9996 (N_9996,N_9617,N_9710);
or U9997 (N_9997,N_9626,N_9748);
or U9998 (N_9998,N_9730,N_9781);
nor U9999 (N_9999,N_9766,N_9637);
or UO_0 (O_0,N_9850,N_9937);
nand UO_1 (O_1,N_9845,N_9999);
and UO_2 (O_2,N_9854,N_9941);
or UO_3 (O_3,N_9907,N_9913);
and UO_4 (O_4,N_9932,N_9989);
or UO_5 (O_5,N_9953,N_9806);
and UO_6 (O_6,N_9873,N_9863);
nor UO_7 (O_7,N_9977,N_9990);
or UO_8 (O_8,N_9848,N_9800);
and UO_9 (O_9,N_9803,N_9819);
or UO_10 (O_10,N_9945,N_9991);
or UO_11 (O_11,N_9939,N_9986);
or UO_12 (O_12,N_9882,N_9843);
or UO_13 (O_13,N_9809,N_9983);
or UO_14 (O_14,N_9925,N_9971);
or UO_15 (O_15,N_9833,N_9846);
or UO_16 (O_16,N_9836,N_9914);
or UO_17 (O_17,N_9827,N_9830);
nand UO_18 (O_18,N_9974,N_9880);
nand UO_19 (O_19,N_9929,N_9852);
nand UO_20 (O_20,N_9958,N_9849);
and UO_21 (O_21,N_9912,N_9969);
or UO_22 (O_22,N_9968,N_9808);
or UO_23 (O_23,N_9928,N_9825);
and UO_24 (O_24,N_9804,N_9911);
or UO_25 (O_25,N_9935,N_9988);
nand UO_26 (O_26,N_9874,N_9970);
and UO_27 (O_27,N_9980,N_9896);
xnor UO_28 (O_28,N_9815,N_9998);
nand UO_29 (O_29,N_9859,N_9857);
and UO_30 (O_30,N_9834,N_9864);
xnor UO_31 (O_31,N_9842,N_9995);
nand UO_32 (O_32,N_9891,N_9975);
and UO_33 (O_33,N_9960,N_9877);
nand UO_34 (O_34,N_9818,N_9805);
nor UO_35 (O_35,N_9917,N_9868);
or UO_36 (O_36,N_9900,N_9853);
and UO_37 (O_37,N_9996,N_9839);
or UO_38 (O_38,N_9931,N_9940);
and UO_39 (O_39,N_9823,N_9963);
nor UO_40 (O_40,N_9910,N_9992);
nor UO_41 (O_41,N_9876,N_9878);
and UO_42 (O_42,N_9887,N_9812);
nor UO_43 (O_43,N_9898,N_9985);
and UO_44 (O_44,N_9817,N_9921);
nor UO_45 (O_45,N_9964,N_9875);
nor UO_46 (O_46,N_9856,N_9895);
nor UO_47 (O_47,N_9973,N_9813);
nand UO_48 (O_48,N_9903,N_9890);
xor UO_49 (O_49,N_9904,N_9872);
nand UO_50 (O_50,N_9909,N_9908);
nor UO_51 (O_51,N_9924,N_9889);
nand UO_52 (O_52,N_9905,N_9824);
and UO_53 (O_53,N_9810,N_9892);
and UO_54 (O_54,N_9918,N_9982);
nor UO_55 (O_55,N_9978,N_9916);
nor UO_56 (O_56,N_9906,N_9972);
or UO_57 (O_57,N_9922,N_9901);
nor UO_58 (O_58,N_9965,N_9984);
xnor UO_59 (O_59,N_9869,N_9851);
or UO_60 (O_60,N_9961,N_9862);
and UO_61 (O_61,N_9954,N_9884);
nor UO_62 (O_62,N_9976,N_9962);
or UO_63 (O_63,N_9811,N_9952);
or UO_64 (O_64,N_9950,N_9870);
nor UO_65 (O_65,N_9888,N_9816);
and UO_66 (O_66,N_9956,N_9879);
nand UO_67 (O_67,N_9923,N_9997);
nor UO_68 (O_68,N_9821,N_9936);
nand UO_69 (O_69,N_9981,N_9926);
nand UO_70 (O_70,N_9949,N_9919);
xor UO_71 (O_71,N_9814,N_9899);
or UO_72 (O_72,N_9927,N_9920);
nand UO_73 (O_73,N_9947,N_9847);
and UO_74 (O_74,N_9855,N_9807);
and UO_75 (O_75,N_9993,N_9897);
or UO_76 (O_76,N_9801,N_9943);
and UO_77 (O_77,N_9942,N_9841);
nor UO_78 (O_78,N_9885,N_9930);
nor UO_79 (O_79,N_9881,N_9865);
or UO_80 (O_80,N_9883,N_9957);
or UO_81 (O_81,N_9994,N_9829);
nand UO_82 (O_82,N_9835,N_9894);
nand UO_83 (O_83,N_9951,N_9893);
nor UO_84 (O_84,N_9955,N_9866);
and UO_85 (O_85,N_9967,N_9861);
and UO_86 (O_86,N_9934,N_9802);
nor UO_87 (O_87,N_9858,N_9820);
nand UO_88 (O_88,N_9831,N_9966);
nand UO_89 (O_89,N_9860,N_9840);
xnor UO_90 (O_90,N_9946,N_9944);
nor UO_91 (O_91,N_9915,N_9837);
nand UO_92 (O_92,N_9838,N_9902);
and UO_93 (O_93,N_9826,N_9938);
or UO_94 (O_94,N_9933,N_9822);
and UO_95 (O_95,N_9959,N_9979);
or UO_96 (O_96,N_9987,N_9871);
xor UO_97 (O_97,N_9948,N_9867);
nor UO_98 (O_98,N_9828,N_9832);
or UO_99 (O_99,N_9886,N_9844);
and UO_100 (O_100,N_9857,N_9891);
and UO_101 (O_101,N_9817,N_9943);
and UO_102 (O_102,N_9935,N_9814);
nand UO_103 (O_103,N_9906,N_9852);
nand UO_104 (O_104,N_9983,N_9891);
nand UO_105 (O_105,N_9819,N_9829);
or UO_106 (O_106,N_9881,N_9820);
or UO_107 (O_107,N_9902,N_9869);
and UO_108 (O_108,N_9809,N_9994);
or UO_109 (O_109,N_9850,N_9916);
or UO_110 (O_110,N_9967,N_9971);
nand UO_111 (O_111,N_9889,N_9944);
or UO_112 (O_112,N_9955,N_9895);
or UO_113 (O_113,N_9838,N_9821);
nor UO_114 (O_114,N_9972,N_9848);
nand UO_115 (O_115,N_9943,N_9904);
nand UO_116 (O_116,N_9861,N_9949);
nand UO_117 (O_117,N_9808,N_9902);
nor UO_118 (O_118,N_9913,N_9843);
and UO_119 (O_119,N_9846,N_9863);
nor UO_120 (O_120,N_9949,N_9905);
nor UO_121 (O_121,N_9839,N_9970);
or UO_122 (O_122,N_9967,N_9979);
xor UO_123 (O_123,N_9849,N_9959);
and UO_124 (O_124,N_9904,N_9841);
and UO_125 (O_125,N_9913,N_9871);
nor UO_126 (O_126,N_9858,N_9955);
or UO_127 (O_127,N_9842,N_9968);
nand UO_128 (O_128,N_9978,N_9808);
xor UO_129 (O_129,N_9804,N_9922);
nor UO_130 (O_130,N_9923,N_9994);
xnor UO_131 (O_131,N_9831,N_9994);
xor UO_132 (O_132,N_9998,N_9856);
xnor UO_133 (O_133,N_9959,N_9812);
nor UO_134 (O_134,N_9845,N_9932);
nor UO_135 (O_135,N_9930,N_9954);
or UO_136 (O_136,N_9830,N_9968);
and UO_137 (O_137,N_9932,N_9839);
xor UO_138 (O_138,N_9857,N_9831);
or UO_139 (O_139,N_9936,N_9858);
or UO_140 (O_140,N_9989,N_9816);
xor UO_141 (O_141,N_9902,N_9949);
nor UO_142 (O_142,N_9823,N_9884);
nor UO_143 (O_143,N_9859,N_9916);
and UO_144 (O_144,N_9834,N_9919);
xnor UO_145 (O_145,N_9832,N_9820);
or UO_146 (O_146,N_9891,N_9941);
or UO_147 (O_147,N_9889,N_9953);
and UO_148 (O_148,N_9933,N_9805);
or UO_149 (O_149,N_9966,N_9931);
or UO_150 (O_150,N_9986,N_9872);
or UO_151 (O_151,N_9956,N_9965);
nor UO_152 (O_152,N_9977,N_9901);
nor UO_153 (O_153,N_9997,N_9995);
xor UO_154 (O_154,N_9910,N_9908);
nor UO_155 (O_155,N_9952,N_9969);
or UO_156 (O_156,N_9832,N_9896);
and UO_157 (O_157,N_9846,N_9873);
nand UO_158 (O_158,N_9916,N_9857);
and UO_159 (O_159,N_9917,N_9903);
or UO_160 (O_160,N_9945,N_9962);
nand UO_161 (O_161,N_9917,N_9957);
nor UO_162 (O_162,N_9801,N_9972);
and UO_163 (O_163,N_9918,N_9883);
nand UO_164 (O_164,N_9851,N_9955);
and UO_165 (O_165,N_9840,N_9822);
and UO_166 (O_166,N_9972,N_9907);
nor UO_167 (O_167,N_9827,N_9915);
nor UO_168 (O_168,N_9805,N_9816);
xnor UO_169 (O_169,N_9996,N_9987);
and UO_170 (O_170,N_9920,N_9881);
or UO_171 (O_171,N_9932,N_9819);
nand UO_172 (O_172,N_9878,N_9953);
and UO_173 (O_173,N_9913,N_9811);
and UO_174 (O_174,N_9982,N_9985);
or UO_175 (O_175,N_9803,N_9876);
and UO_176 (O_176,N_9807,N_9903);
nand UO_177 (O_177,N_9984,N_9986);
xor UO_178 (O_178,N_9983,N_9940);
xor UO_179 (O_179,N_9979,N_9951);
nor UO_180 (O_180,N_9996,N_9937);
and UO_181 (O_181,N_9885,N_9816);
nor UO_182 (O_182,N_9933,N_9814);
or UO_183 (O_183,N_9958,N_9839);
nand UO_184 (O_184,N_9954,N_9874);
nor UO_185 (O_185,N_9972,N_9840);
nor UO_186 (O_186,N_9958,N_9994);
and UO_187 (O_187,N_9889,N_9856);
and UO_188 (O_188,N_9838,N_9895);
or UO_189 (O_189,N_9932,N_9946);
nand UO_190 (O_190,N_9804,N_9869);
or UO_191 (O_191,N_9821,N_9814);
nand UO_192 (O_192,N_9994,N_9821);
and UO_193 (O_193,N_9958,N_9911);
nor UO_194 (O_194,N_9826,N_9940);
or UO_195 (O_195,N_9902,N_9960);
nand UO_196 (O_196,N_9952,N_9899);
and UO_197 (O_197,N_9950,N_9821);
or UO_198 (O_198,N_9896,N_9947);
or UO_199 (O_199,N_9872,N_9976);
nand UO_200 (O_200,N_9909,N_9835);
nor UO_201 (O_201,N_9959,N_9860);
and UO_202 (O_202,N_9953,N_9805);
or UO_203 (O_203,N_9922,N_9818);
and UO_204 (O_204,N_9939,N_9874);
and UO_205 (O_205,N_9960,N_9837);
nor UO_206 (O_206,N_9807,N_9843);
or UO_207 (O_207,N_9855,N_9953);
and UO_208 (O_208,N_9874,N_9919);
and UO_209 (O_209,N_9913,N_9975);
nand UO_210 (O_210,N_9880,N_9933);
nor UO_211 (O_211,N_9877,N_9951);
nor UO_212 (O_212,N_9877,N_9862);
nand UO_213 (O_213,N_9937,N_9902);
xor UO_214 (O_214,N_9912,N_9834);
xor UO_215 (O_215,N_9972,N_9877);
nand UO_216 (O_216,N_9958,N_9967);
or UO_217 (O_217,N_9828,N_9960);
and UO_218 (O_218,N_9892,N_9909);
and UO_219 (O_219,N_9957,N_9807);
or UO_220 (O_220,N_9898,N_9906);
or UO_221 (O_221,N_9895,N_9925);
xor UO_222 (O_222,N_9934,N_9904);
nor UO_223 (O_223,N_9900,N_9815);
or UO_224 (O_224,N_9893,N_9972);
nor UO_225 (O_225,N_9908,N_9890);
or UO_226 (O_226,N_9856,N_9898);
and UO_227 (O_227,N_9818,N_9810);
nor UO_228 (O_228,N_9817,N_9941);
nand UO_229 (O_229,N_9898,N_9805);
nand UO_230 (O_230,N_9887,N_9914);
or UO_231 (O_231,N_9891,N_9971);
and UO_232 (O_232,N_9846,N_9990);
nor UO_233 (O_233,N_9937,N_9864);
nor UO_234 (O_234,N_9998,N_9957);
and UO_235 (O_235,N_9816,N_9819);
xnor UO_236 (O_236,N_9867,N_9952);
xnor UO_237 (O_237,N_9921,N_9951);
nor UO_238 (O_238,N_9817,N_9907);
xnor UO_239 (O_239,N_9952,N_9890);
nor UO_240 (O_240,N_9866,N_9868);
or UO_241 (O_241,N_9832,N_9956);
nand UO_242 (O_242,N_9983,N_9832);
nor UO_243 (O_243,N_9801,N_9946);
nand UO_244 (O_244,N_9823,N_9967);
nor UO_245 (O_245,N_9864,N_9808);
or UO_246 (O_246,N_9967,N_9936);
nor UO_247 (O_247,N_9932,N_9903);
and UO_248 (O_248,N_9900,N_9826);
or UO_249 (O_249,N_9971,N_9805);
and UO_250 (O_250,N_9801,N_9870);
xnor UO_251 (O_251,N_9942,N_9863);
or UO_252 (O_252,N_9998,N_9801);
nand UO_253 (O_253,N_9856,N_9814);
or UO_254 (O_254,N_9802,N_9849);
nor UO_255 (O_255,N_9900,N_9954);
nor UO_256 (O_256,N_9921,N_9834);
and UO_257 (O_257,N_9865,N_9912);
nor UO_258 (O_258,N_9999,N_9985);
nand UO_259 (O_259,N_9990,N_9964);
or UO_260 (O_260,N_9884,N_9941);
or UO_261 (O_261,N_9998,N_9858);
nor UO_262 (O_262,N_9801,N_9890);
nand UO_263 (O_263,N_9894,N_9826);
or UO_264 (O_264,N_9866,N_9920);
or UO_265 (O_265,N_9835,N_9991);
and UO_266 (O_266,N_9812,N_9910);
or UO_267 (O_267,N_9815,N_9910);
nor UO_268 (O_268,N_9930,N_9842);
nand UO_269 (O_269,N_9801,N_9854);
nor UO_270 (O_270,N_9848,N_9908);
nor UO_271 (O_271,N_9835,N_9860);
nor UO_272 (O_272,N_9805,N_9836);
xor UO_273 (O_273,N_9840,N_9862);
or UO_274 (O_274,N_9861,N_9966);
nor UO_275 (O_275,N_9990,N_9908);
nand UO_276 (O_276,N_9928,N_9803);
nor UO_277 (O_277,N_9917,N_9948);
and UO_278 (O_278,N_9988,N_9844);
or UO_279 (O_279,N_9958,N_9940);
nand UO_280 (O_280,N_9900,N_9890);
or UO_281 (O_281,N_9991,N_9872);
nand UO_282 (O_282,N_9967,N_9955);
or UO_283 (O_283,N_9875,N_9846);
and UO_284 (O_284,N_9942,N_9816);
nand UO_285 (O_285,N_9861,N_9886);
nor UO_286 (O_286,N_9903,N_9817);
nand UO_287 (O_287,N_9908,N_9823);
xnor UO_288 (O_288,N_9919,N_9806);
or UO_289 (O_289,N_9888,N_9902);
nand UO_290 (O_290,N_9810,N_9896);
and UO_291 (O_291,N_9873,N_9851);
nor UO_292 (O_292,N_9909,N_9977);
and UO_293 (O_293,N_9970,N_9922);
nor UO_294 (O_294,N_9815,N_9817);
nor UO_295 (O_295,N_9935,N_9948);
xor UO_296 (O_296,N_9998,N_9849);
xnor UO_297 (O_297,N_9917,N_9999);
nand UO_298 (O_298,N_9938,N_9929);
nand UO_299 (O_299,N_9974,N_9815);
and UO_300 (O_300,N_9844,N_9833);
and UO_301 (O_301,N_9960,N_9968);
nand UO_302 (O_302,N_9926,N_9944);
and UO_303 (O_303,N_9976,N_9883);
and UO_304 (O_304,N_9819,N_9855);
nand UO_305 (O_305,N_9997,N_9909);
and UO_306 (O_306,N_9872,N_9841);
or UO_307 (O_307,N_9860,N_9834);
and UO_308 (O_308,N_9808,N_9816);
nand UO_309 (O_309,N_9957,N_9914);
and UO_310 (O_310,N_9859,N_9877);
nor UO_311 (O_311,N_9826,N_9867);
or UO_312 (O_312,N_9834,N_9823);
or UO_313 (O_313,N_9911,N_9822);
xor UO_314 (O_314,N_9982,N_9911);
nor UO_315 (O_315,N_9967,N_9946);
or UO_316 (O_316,N_9828,N_9875);
or UO_317 (O_317,N_9845,N_9971);
and UO_318 (O_318,N_9824,N_9931);
xor UO_319 (O_319,N_9875,N_9804);
and UO_320 (O_320,N_9926,N_9967);
and UO_321 (O_321,N_9864,N_9843);
xnor UO_322 (O_322,N_9845,N_9897);
nor UO_323 (O_323,N_9856,N_9965);
and UO_324 (O_324,N_9918,N_9887);
or UO_325 (O_325,N_9888,N_9854);
nand UO_326 (O_326,N_9957,N_9825);
and UO_327 (O_327,N_9863,N_9859);
nor UO_328 (O_328,N_9955,N_9811);
nand UO_329 (O_329,N_9809,N_9866);
and UO_330 (O_330,N_9857,N_9952);
and UO_331 (O_331,N_9881,N_9838);
nand UO_332 (O_332,N_9948,N_9863);
and UO_333 (O_333,N_9867,N_9936);
nand UO_334 (O_334,N_9880,N_9879);
nor UO_335 (O_335,N_9905,N_9977);
nand UO_336 (O_336,N_9847,N_9979);
and UO_337 (O_337,N_9974,N_9881);
xnor UO_338 (O_338,N_9890,N_9893);
xnor UO_339 (O_339,N_9973,N_9971);
nor UO_340 (O_340,N_9826,N_9827);
or UO_341 (O_341,N_9951,N_9820);
xnor UO_342 (O_342,N_9824,N_9911);
nand UO_343 (O_343,N_9938,N_9960);
and UO_344 (O_344,N_9867,N_9962);
nor UO_345 (O_345,N_9931,N_9845);
nand UO_346 (O_346,N_9830,N_9936);
and UO_347 (O_347,N_9994,N_9999);
or UO_348 (O_348,N_9963,N_9828);
nor UO_349 (O_349,N_9963,N_9844);
nand UO_350 (O_350,N_9845,N_9861);
nor UO_351 (O_351,N_9924,N_9982);
xor UO_352 (O_352,N_9804,N_9865);
and UO_353 (O_353,N_9866,N_9965);
or UO_354 (O_354,N_9825,N_9940);
nor UO_355 (O_355,N_9887,N_9886);
or UO_356 (O_356,N_9894,N_9810);
nor UO_357 (O_357,N_9940,N_9882);
nor UO_358 (O_358,N_9827,N_9954);
nor UO_359 (O_359,N_9825,N_9898);
nand UO_360 (O_360,N_9942,N_9864);
or UO_361 (O_361,N_9899,N_9971);
nand UO_362 (O_362,N_9926,N_9984);
and UO_363 (O_363,N_9954,N_9828);
nor UO_364 (O_364,N_9921,N_9824);
nand UO_365 (O_365,N_9994,N_9814);
and UO_366 (O_366,N_9908,N_9885);
nor UO_367 (O_367,N_9873,N_9917);
and UO_368 (O_368,N_9967,N_9907);
nand UO_369 (O_369,N_9897,N_9855);
nor UO_370 (O_370,N_9983,N_9883);
xor UO_371 (O_371,N_9968,N_9852);
nand UO_372 (O_372,N_9996,N_9854);
nor UO_373 (O_373,N_9943,N_9873);
nor UO_374 (O_374,N_9901,N_9974);
or UO_375 (O_375,N_9918,N_9985);
nor UO_376 (O_376,N_9889,N_9822);
nor UO_377 (O_377,N_9921,N_9931);
and UO_378 (O_378,N_9939,N_9888);
nand UO_379 (O_379,N_9887,N_9895);
nand UO_380 (O_380,N_9953,N_9846);
and UO_381 (O_381,N_9950,N_9935);
nand UO_382 (O_382,N_9952,N_9992);
and UO_383 (O_383,N_9993,N_9934);
nor UO_384 (O_384,N_9892,N_9864);
nand UO_385 (O_385,N_9811,N_9808);
nor UO_386 (O_386,N_9965,N_9981);
nand UO_387 (O_387,N_9936,N_9845);
nor UO_388 (O_388,N_9979,N_9962);
and UO_389 (O_389,N_9910,N_9820);
xnor UO_390 (O_390,N_9873,N_9869);
nand UO_391 (O_391,N_9972,N_9800);
nor UO_392 (O_392,N_9922,N_9980);
or UO_393 (O_393,N_9885,N_9941);
and UO_394 (O_394,N_9812,N_9816);
or UO_395 (O_395,N_9997,N_9958);
nor UO_396 (O_396,N_9934,N_9902);
nand UO_397 (O_397,N_9976,N_9862);
or UO_398 (O_398,N_9833,N_9984);
and UO_399 (O_399,N_9876,N_9899);
and UO_400 (O_400,N_9820,N_9902);
or UO_401 (O_401,N_9972,N_9819);
nor UO_402 (O_402,N_9869,N_9942);
or UO_403 (O_403,N_9924,N_9879);
and UO_404 (O_404,N_9827,N_9805);
or UO_405 (O_405,N_9861,N_9991);
and UO_406 (O_406,N_9927,N_9876);
nor UO_407 (O_407,N_9997,N_9969);
or UO_408 (O_408,N_9810,N_9985);
or UO_409 (O_409,N_9842,N_9835);
or UO_410 (O_410,N_9886,N_9995);
or UO_411 (O_411,N_9863,N_9886);
or UO_412 (O_412,N_9845,N_9935);
nand UO_413 (O_413,N_9917,N_9955);
or UO_414 (O_414,N_9998,N_9966);
nor UO_415 (O_415,N_9884,N_9866);
and UO_416 (O_416,N_9802,N_9959);
nor UO_417 (O_417,N_9896,N_9801);
xor UO_418 (O_418,N_9930,N_9913);
and UO_419 (O_419,N_9878,N_9822);
and UO_420 (O_420,N_9890,N_9872);
or UO_421 (O_421,N_9995,N_9836);
and UO_422 (O_422,N_9942,N_9957);
and UO_423 (O_423,N_9926,N_9840);
or UO_424 (O_424,N_9911,N_9868);
nor UO_425 (O_425,N_9879,N_9827);
nand UO_426 (O_426,N_9834,N_9952);
or UO_427 (O_427,N_9815,N_9983);
nor UO_428 (O_428,N_9982,N_9855);
nor UO_429 (O_429,N_9841,N_9991);
and UO_430 (O_430,N_9938,N_9862);
or UO_431 (O_431,N_9823,N_9872);
nand UO_432 (O_432,N_9975,N_9828);
nor UO_433 (O_433,N_9873,N_9811);
or UO_434 (O_434,N_9822,N_9957);
nand UO_435 (O_435,N_9880,N_9837);
xnor UO_436 (O_436,N_9822,N_9821);
nor UO_437 (O_437,N_9803,N_9969);
or UO_438 (O_438,N_9945,N_9822);
or UO_439 (O_439,N_9813,N_9917);
or UO_440 (O_440,N_9967,N_9818);
nand UO_441 (O_441,N_9819,N_9912);
nand UO_442 (O_442,N_9990,N_9857);
or UO_443 (O_443,N_9937,N_9926);
nand UO_444 (O_444,N_9901,N_9944);
nor UO_445 (O_445,N_9913,N_9978);
and UO_446 (O_446,N_9890,N_9993);
nand UO_447 (O_447,N_9996,N_9819);
and UO_448 (O_448,N_9922,N_9906);
xor UO_449 (O_449,N_9985,N_9815);
nand UO_450 (O_450,N_9954,N_9866);
or UO_451 (O_451,N_9957,N_9922);
and UO_452 (O_452,N_9801,N_9981);
or UO_453 (O_453,N_9830,N_9817);
nand UO_454 (O_454,N_9892,N_9949);
nand UO_455 (O_455,N_9873,N_9972);
nor UO_456 (O_456,N_9897,N_9917);
and UO_457 (O_457,N_9819,N_9856);
nor UO_458 (O_458,N_9873,N_9864);
nor UO_459 (O_459,N_9861,N_9851);
or UO_460 (O_460,N_9859,N_9837);
or UO_461 (O_461,N_9919,N_9848);
and UO_462 (O_462,N_9986,N_9969);
and UO_463 (O_463,N_9840,N_9861);
or UO_464 (O_464,N_9840,N_9857);
and UO_465 (O_465,N_9814,N_9831);
and UO_466 (O_466,N_9969,N_9903);
and UO_467 (O_467,N_9857,N_9930);
nand UO_468 (O_468,N_9907,N_9881);
and UO_469 (O_469,N_9990,N_9910);
nor UO_470 (O_470,N_9884,N_9833);
nand UO_471 (O_471,N_9967,N_9999);
nor UO_472 (O_472,N_9906,N_9963);
and UO_473 (O_473,N_9929,N_9924);
nor UO_474 (O_474,N_9971,N_9893);
nand UO_475 (O_475,N_9908,N_9837);
and UO_476 (O_476,N_9908,N_9960);
xnor UO_477 (O_477,N_9873,N_9993);
and UO_478 (O_478,N_9832,N_9873);
nor UO_479 (O_479,N_9869,N_9909);
and UO_480 (O_480,N_9863,N_9999);
nor UO_481 (O_481,N_9892,N_9822);
or UO_482 (O_482,N_9992,N_9968);
nand UO_483 (O_483,N_9979,N_9957);
or UO_484 (O_484,N_9928,N_9977);
or UO_485 (O_485,N_9802,N_9808);
xor UO_486 (O_486,N_9941,N_9816);
nor UO_487 (O_487,N_9838,N_9811);
or UO_488 (O_488,N_9811,N_9885);
nand UO_489 (O_489,N_9803,N_9827);
xnor UO_490 (O_490,N_9985,N_9881);
or UO_491 (O_491,N_9854,N_9861);
nand UO_492 (O_492,N_9919,N_9990);
nand UO_493 (O_493,N_9817,N_9869);
nand UO_494 (O_494,N_9846,N_9869);
or UO_495 (O_495,N_9838,N_9853);
nand UO_496 (O_496,N_9957,N_9995);
nand UO_497 (O_497,N_9812,N_9886);
and UO_498 (O_498,N_9976,N_9850);
and UO_499 (O_499,N_9890,N_9899);
or UO_500 (O_500,N_9872,N_9843);
xor UO_501 (O_501,N_9843,N_9895);
nor UO_502 (O_502,N_9934,N_9807);
nor UO_503 (O_503,N_9810,N_9852);
xor UO_504 (O_504,N_9884,N_9975);
nor UO_505 (O_505,N_9885,N_9894);
or UO_506 (O_506,N_9827,N_9939);
or UO_507 (O_507,N_9960,N_9815);
and UO_508 (O_508,N_9817,N_9942);
nor UO_509 (O_509,N_9820,N_9965);
or UO_510 (O_510,N_9971,N_9886);
nand UO_511 (O_511,N_9976,N_9982);
nor UO_512 (O_512,N_9872,N_9990);
and UO_513 (O_513,N_9814,N_9893);
nor UO_514 (O_514,N_9911,N_9871);
nor UO_515 (O_515,N_9836,N_9909);
or UO_516 (O_516,N_9824,N_9853);
nor UO_517 (O_517,N_9928,N_9973);
nor UO_518 (O_518,N_9986,N_9925);
or UO_519 (O_519,N_9845,N_9802);
and UO_520 (O_520,N_9991,N_9912);
xnor UO_521 (O_521,N_9994,N_9897);
or UO_522 (O_522,N_9965,N_9810);
nand UO_523 (O_523,N_9993,N_9948);
and UO_524 (O_524,N_9850,N_9890);
nor UO_525 (O_525,N_9904,N_9961);
nor UO_526 (O_526,N_9953,N_9834);
and UO_527 (O_527,N_9821,N_9905);
and UO_528 (O_528,N_9879,N_9986);
nor UO_529 (O_529,N_9850,N_9834);
and UO_530 (O_530,N_9822,N_9897);
or UO_531 (O_531,N_9817,N_9969);
xnor UO_532 (O_532,N_9940,N_9979);
and UO_533 (O_533,N_9868,N_9828);
or UO_534 (O_534,N_9905,N_9913);
or UO_535 (O_535,N_9976,N_9847);
nand UO_536 (O_536,N_9971,N_9908);
and UO_537 (O_537,N_9925,N_9917);
xnor UO_538 (O_538,N_9926,N_9923);
xnor UO_539 (O_539,N_9954,N_9847);
nor UO_540 (O_540,N_9871,N_9872);
nand UO_541 (O_541,N_9982,N_9865);
nor UO_542 (O_542,N_9960,N_9981);
and UO_543 (O_543,N_9986,N_9821);
and UO_544 (O_544,N_9927,N_9892);
nand UO_545 (O_545,N_9954,N_9968);
nand UO_546 (O_546,N_9908,N_9969);
nor UO_547 (O_547,N_9927,N_9923);
nand UO_548 (O_548,N_9904,N_9939);
nor UO_549 (O_549,N_9967,N_9848);
or UO_550 (O_550,N_9854,N_9914);
and UO_551 (O_551,N_9900,N_9840);
and UO_552 (O_552,N_9866,N_9899);
nor UO_553 (O_553,N_9925,N_9913);
nor UO_554 (O_554,N_9949,N_9888);
xnor UO_555 (O_555,N_9840,N_9806);
or UO_556 (O_556,N_9996,N_9901);
or UO_557 (O_557,N_9853,N_9951);
nand UO_558 (O_558,N_9897,N_9850);
and UO_559 (O_559,N_9938,N_9865);
and UO_560 (O_560,N_9943,N_9869);
xor UO_561 (O_561,N_9917,N_9962);
and UO_562 (O_562,N_9939,N_9934);
and UO_563 (O_563,N_9925,N_9820);
or UO_564 (O_564,N_9952,N_9959);
xor UO_565 (O_565,N_9879,N_9819);
and UO_566 (O_566,N_9848,N_9929);
nor UO_567 (O_567,N_9865,N_9902);
xnor UO_568 (O_568,N_9831,N_9848);
nor UO_569 (O_569,N_9898,N_9970);
or UO_570 (O_570,N_9932,N_9886);
nand UO_571 (O_571,N_9820,N_9967);
nand UO_572 (O_572,N_9875,N_9931);
or UO_573 (O_573,N_9826,N_9964);
and UO_574 (O_574,N_9862,N_9844);
nor UO_575 (O_575,N_9812,N_9867);
xnor UO_576 (O_576,N_9907,N_9923);
or UO_577 (O_577,N_9903,N_9881);
nand UO_578 (O_578,N_9865,N_9871);
nor UO_579 (O_579,N_9938,N_9833);
nor UO_580 (O_580,N_9991,N_9892);
xor UO_581 (O_581,N_9825,N_9905);
nand UO_582 (O_582,N_9890,N_9974);
or UO_583 (O_583,N_9860,N_9821);
nor UO_584 (O_584,N_9979,N_9983);
or UO_585 (O_585,N_9803,N_9921);
xor UO_586 (O_586,N_9817,N_9884);
nand UO_587 (O_587,N_9936,N_9840);
nor UO_588 (O_588,N_9994,N_9826);
nor UO_589 (O_589,N_9987,N_9904);
and UO_590 (O_590,N_9931,N_9806);
or UO_591 (O_591,N_9900,N_9831);
nand UO_592 (O_592,N_9978,N_9986);
nor UO_593 (O_593,N_9886,N_9823);
or UO_594 (O_594,N_9843,N_9823);
nand UO_595 (O_595,N_9843,N_9973);
nand UO_596 (O_596,N_9995,N_9818);
xor UO_597 (O_597,N_9915,N_9853);
nand UO_598 (O_598,N_9830,N_9967);
and UO_599 (O_599,N_9982,N_9887);
nand UO_600 (O_600,N_9800,N_9828);
xor UO_601 (O_601,N_9910,N_9894);
nand UO_602 (O_602,N_9945,N_9820);
xor UO_603 (O_603,N_9805,N_9985);
nand UO_604 (O_604,N_9804,N_9960);
and UO_605 (O_605,N_9823,N_9891);
or UO_606 (O_606,N_9990,N_9823);
and UO_607 (O_607,N_9993,N_9917);
nand UO_608 (O_608,N_9852,N_9966);
and UO_609 (O_609,N_9935,N_9829);
and UO_610 (O_610,N_9881,N_9948);
and UO_611 (O_611,N_9888,N_9839);
nor UO_612 (O_612,N_9859,N_9850);
and UO_613 (O_613,N_9820,N_9803);
nor UO_614 (O_614,N_9842,N_9821);
nor UO_615 (O_615,N_9841,N_9974);
xor UO_616 (O_616,N_9988,N_9824);
nand UO_617 (O_617,N_9937,N_9805);
and UO_618 (O_618,N_9984,N_9983);
nand UO_619 (O_619,N_9816,N_9858);
nand UO_620 (O_620,N_9956,N_9977);
nor UO_621 (O_621,N_9957,N_9967);
nor UO_622 (O_622,N_9879,N_9824);
nand UO_623 (O_623,N_9969,N_9889);
xor UO_624 (O_624,N_9995,N_9879);
or UO_625 (O_625,N_9831,N_9903);
and UO_626 (O_626,N_9992,N_9939);
or UO_627 (O_627,N_9916,N_9815);
and UO_628 (O_628,N_9881,N_9941);
or UO_629 (O_629,N_9931,N_9850);
or UO_630 (O_630,N_9817,N_9915);
nand UO_631 (O_631,N_9848,N_9927);
and UO_632 (O_632,N_9989,N_9979);
nand UO_633 (O_633,N_9996,N_9867);
or UO_634 (O_634,N_9851,N_9911);
or UO_635 (O_635,N_9881,N_9822);
and UO_636 (O_636,N_9896,N_9816);
and UO_637 (O_637,N_9977,N_9957);
or UO_638 (O_638,N_9959,N_9856);
nand UO_639 (O_639,N_9875,N_9849);
and UO_640 (O_640,N_9835,N_9848);
nand UO_641 (O_641,N_9992,N_9882);
or UO_642 (O_642,N_9983,N_9870);
nor UO_643 (O_643,N_9842,N_9819);
or UO_644 (O_644,N_9957,N_9868);
and UO_645 (O_645,N_9951,N_9866);
nand UO_646 (O_646,N_9944,N_9985);
nand UO_647 (O_647,N_9800,N_9899);
or UO_648 (O_648,N_9928,N_9802);
nor UO_649 (O_649,N_9933,N_9894);
nand UO_650 (O_650,N_9993,N_9899);
or UO_651 (O_651,N_9959,N_9947);
or UO_652 (O_652,N_9870,N_9818);
nor UO_653 (O_653,N_9988,N_9889);
and UO_654 (O_654,N_9969,N_9841);
nor UO_655 (O_655,N_9933,N_9900);
or UO_656 (O_656,N_9831,N_9952);
or UO_657 (O_657,N_9866,N_9915);
and UO_658 (O_658,N_9888,N_9831);
nand UO_659 (O_659,N_9944,N_9891);
nor UO_660 (O_660,N_9875,N_9944);
and UO_661 (O_661,N_9950,N_9978);
nand UO_662 (O_662,N_9956,N_9970);
or UO_663 (O_663,N_9870,N_9922);
nand UO_664 (O_664,N_9996,N_9970);
and UO_665 (O_665,N_9951,N_9876);
xnor UO_666 (O_666,N_9940,N_9818);
and UO_667 (O_667,N_9833,N_9970);
or UO_668 (O_668,N_9981,N_9897);
nor UO_669 (O_669,N_9904,N_9906);
nor UO_670 (O_670,N_9925,N_9802);
nand UO_671 (O_671,N_9802,N_9969);
nand UO_672 (O_672,N_9992,N_9859);
and UO_673 (O_673,N_9950,N_9872);
nor UO_674 (O_674,N_9837,N_9887);
and UO_675 (O_675,N_9933,N_9891);
nor UO_676 (O_676,N_9942,N_9900);
and UO_677 (O_677,N_9955,N_9840);
and UO_678 (O_678,N_9949,N_9840);
xnor UO_679 (O_679,N_9921,N_9925);
or UO_680 (O_680,N_9919,N_9808);
and UO_681 (O_681,N_9905,N_9932);
nor UO_682 (O_682,N_9916,N_9935);
or UO_683 (O_683,N_9947,N_9804);
and UO_684 (O_684,N_9892,N_9989);
or UO_685 (O_685,N_9998,N_9816);
nand UO_686 (O_686,N_9839,N_9878);
and UO_687 (O_687,N_9927,N_9854);
nor UO_688 (O_688,N_9950,N_9842);
or UO_689 (O_689,N_9818,N_9996);
and UO_690 (O_690,N_9824,N_9934);
or UO_691 (O_691,N_9815,N_9903);
and UO_692 (O_692,N_9911,N_9976);
and UO_693 (O_693,N_9990,N_9972);
nand UO_694 (O_694,N_9816,N_9847);
xor UO_695 (O_695,N_9959,N_9934);
nor UO_696 (O_696,N_9898,N_9900);
nor UO_697 (O_697,N_9939,N_9800);
nand UO_698 (O_698,N_9824,N_9956);
nor UO_699 (O_699,N_9967,N_9944);
nor UO_700 (O_700,N_9881,N_9929);
nand UO_701 (O_701,N_9882,N_9894);
nand UO_702 (O_702,N_9859,N_9912);
nor UO_703 (O_703,N_9959,N_9996);
or UO_704 (O_704,N_9982,N_9854);
nand UO_705 (O_705,N_9965,N_9809);
nand UO_706 (O_706,N_9829,N_9925);
or UO_707 (O_707,N_9990,N_9924);
nand UO_708 (O_708,N_9896,N_9979);
or UO_709 (O_709,N_9932,N_9969);
and UO_710 (O_710,N_9962,N_9836);
and UO_711 (O_711,N_9917,N_9890);
nor UO_712 (O_712,N_9860,N_9944);
and UO_713 (O_713,N_9837,N_9961);
and UO_714 (O_714,N_9889,N_9977);
nor UO_715 (O_715,N_9854,N_9864);
or UO_716 (O_716,N_9971,N_9857);
nor UO_717 (O_717,N_9820,N_9898);
or UO_718 (O_718,N_9805,N_9941);
and UO_719 (O_719,N_9896,N_9967);
and UO_720 (O_720,N_9894,N_9825);
nand UO_721 (O_721,N_9980,N_9905);
or UO_722 (O_722,N_9841,N_9839);
nor UO_723 (O_723,N_9841,N_9820);
nand UO_724 (O_724,N_9940,N_9996);
nand UO_725 (O_725,N_9902,N_9896);
and UO_726 (O_726,N_9860,N_9978);
xor UO_727 (O_727,N_9975,N_9803);
nand UO_728 (O_728,N_9984,N_9933);
and UO_729 (O_729,N_9981,N_9859);
or UO_730 (O_730,N_9950,N_9861);
xor UO_731 (O_731,N_9881,N_9940);
nor UO_732 (O_732,N_9925,N_9827);
xor UO_733 (O_733,N_9872,N_9829);
or UO_734 (O_734,N_9888,N_9838);
and UO_735 (O_735,N_9991,N_9822);
xor UO_736 (O_736,N_9862,N_9824);
or UO_737 (O_737,N_9906,N_9921);
nor UO_738 (O_738,N_9802,N_9929);
or UO_739 (O_739,N_9816,N_9990);
nand UO_740 (O_740,N_9921,N_9879);
nand UO_741 (O_741,N_9880,N_9882);
and UO_742 (O_742,N_9869,N_9976);
or UO_743 (O_743,N_9961,N_9825);
nor UO_744 (O_744,N_9993,N_9823);
nand UO_745 (O_745,N_9983,N_9852);
nand UO_746 (O_746,N_9884,N_9934);
or UO_747 (O_747,N_9903,N_9965);
or UO_748 (O_748,N_9823,N_9934);
nor UO_749 (O_749,N_9906,N_9956);
nand UO_750 (O_750,N_9849,N_9851);
nand UO_751 (O_751,N_9809,N_9833);
nand UO_752 (O_752,N_9932,N_9863);
nor UO_753 (O_753,N_9806,N_9939);
or UO_754 (O_754,N_9818,N_9879);
or UO_755 (O_755,N_9813,N_9869);
nand UO_756 (O_756,N_9910,N_9917);
nand UO_757 (O_757,N_9937,N_9880);
xor UO_758 (O_758,N_9979,N_9960);
and UO_759 (O_759,N_9820,N_9852);
xnor UO_760 (O_760,N_9850,N_9840);
and UO_761 (O_761,N_9958,N_9837);
nand UO_762 (O_762,N_9977,N_9863);
and UO_763 (O_763,N_9866,N_9835);
or UO_764 (O_764,N_9985,N_9891);
or UO_765 (O_765,N_9812,N_9892);
and UO_766 (O_766,N_9916,N_9957);
xor UO_767 (O_767,N_9898,N_9813);
and UO_768 (O_768,N_9835,N_9979);
or UO_769 (O_769,N_9923,N_9939);
nor UO_770 (O_770,N_9800,N_9942);
and UO_771 (O_771,N_9962,N_9880);
nor UO_772 (O_772,N_9928,N_9981);
nand UO_773 (O_773,N_9994,N_9975);
or UO_774 (O_774,N_9944,N_9980);
and UO_775 (O_775,N_9892,N_9993);
nand UO_776 (O_776,N_9825,N_9987);
nand UO_777 (O_777,N_9803,N_9837);
nand UO_778 (O_778,N_9989,N_9803);
and UO_779 (O_779,N_9939,N_9802);
nand UO_780 (O_780,N_9806,N_9988);
nor UO_781 (O_781,N_9909,N_9878);
and UO_782 (O_782,N_9898,N_9976);
nor UO_783 (O_783,N_9803,N_9835);
or UO_784 (O_784,N_9956,N_9904);
and UO_785 (O_785,N_9949,N_9806);
xnor UO_786 (O_786,N_9985,N_9964);
nor UO_787 (O_787,N_9833,N_9966);
or UO_788 (O_788,N_9846,N_9832);
nor UO_789 (O_789,N_9921,N_9832);
or UO_790 (O_790,N_9924,N_9849);
or UO_791 (O_791,N_9933,N_9869);
or UO_792 (O_792,N_9976,N_9975);
or UO_793 (O_793,N_9912,N_9905);
nand UO_794 (O_794,N_9978,N_9889);
and UO_795 (O_795,N_9879,N_9972);
nor UO_796 (O_796,N_9993,N_9809);
nand UO_797 (O_797,N_9845,N_9938);
nor UO_798 (O_798,N_9833,N_9922);
and UO_799 (O_799,N_9971,N_9874);
xor UO_800 (O_800,N_9816,N_9943);
nor UO_801 (O_801,N_9930,N_9994);
xor UO_802 (O_802,N_9811,N_9940);
or UO_803 (O_803,N_9829,N_9831);
and UO_804 (O_804,N_9818,N_9924);
and UO_805 (O_805,N_9853,N_9942);
and UO_806 (O_806,N_9886,N_9910);
nor UO_807 (O_807,N_9968,N_9911);
nand UO_808 (O_808,N_9817,N_9965);
nand UO_809 (O_809,N_9803,N_9933);
nand UO_810 (O_810,N_9911,N_9855);
nand UO_811 (O_811,N_9863,N_9986);
nor UO_812 (O_812,N_9998,N_9870);
or UO_813 (O_813,N_9863,N_9801);
or UO_814 (O_814,N_9881,N_9925);
xnor UO_815 (O_815,N_9866,N_9814);
nand UO_816 (O_816,N_9972,N_9960);
xor UO_817 (O_817,N_9951,N_9900);
nand UO_818 (O_818,N_9917,N_9970);
or UO_819 (O_819,N_9903,N_9895);
nor UO_820 (O_820,N_9896,N_9963);
xor UO_821 (O_821,N_9874,N_9827);
nor UO_822 (O_822,N_9846,N_9834);
nand UO_823 (O_823,N_9853,N_9946);
xor UO_824 (O_824,N_9835,N_9930);
nor UO_825 (O_825,N_9915,N_9965);
nor UO_826 (O_826,N_9969,N_9916);
nand UO_827 (O_827,N_9828,N_9980);
or UO_828 (O_828,N_9845,N_9814);
nand UO_829 (O_829,N_9893,N_9815);
nand UO_830 (O_830,N_9883,N_9812);
or UO_831 (O_831,N_9847,N_9905);
nor UO_832 (O_832,N_9804,N_9932);
nand UO_833 (O_833,N_9924,N_9802);
or UO_834 (O_834,N_9835,N_9855);
nand UO_835 (O_835,N_9825,N_9851);
and UO_836 (O_836,N_9856,N_9980);
nor UO_837 (O_837,N_9814,N_9944);
nor UO_838 (O_838,N_9930,N_9952);
nand UO_839 (O_839,N_9981,N_9803);
or UO_840 (O_840,N_9925,N_9983);
or UO_841 (O_841,N_9857,N_9937);
or UO_842 (O_842,N_9957,N_9981);
and UO_843 (O_843,N_9858,N_9966);
nand UO_844 (O_844,N_9918,N_9834);
xor UO_845 (O_845,N_9986,N_9899);
xor UO_846 (O_846,N_9817,N_9868);
and UO_847 (O_847,N_9840,N_9919);
or UO_848 (O_848,N_9863,N_9938);
or UO_849 (O_849,N_9946,N_9841);
and UO_850 (O_850,N_9814,N_9979);
nand UO_851 (O_851,N_9818,N_9816);
nor UO_852 (O_852,N_9899,N_9822);
nand UO_853 (O_853,N_9844,N_9838);
nand UO_854 (O_854,N_9836,N_9817);
and UO_855 (O_855,N_9951,N_9954);
nor UO_856 (O_856,N_9930,N_9963);
or UO_857 (O_857,N_9811,N_9975);
or UO_858 (O_858,N_9898,N_9989);
nor UO_859 (O_859,N_9880,N_9894);
and UO_860 (O_860,N_9955,N_9951);
xnor UO_861 (O_861,N_9821,N_9901);
nor UO_862 (O_862,N_9824,N_9826);
nor UO_863 (O_863,N_9817,N_9838);
nor UO_864 (O_864,N_9919,N_9847);
or UO_865 (O_865,N_9939,N_9913);
nand UO_866 (O_866,N_9963,N_9997);
xnor UO_867 (O_867,N_9865,N_9963);
and UO_868 (O_868,N_9802,N_9858);
nor UO_869 (O_869,N_9994,N_9845);
or UO_870 (O_870,N_9809,N_9987);
and UO_871 (O_871,N_9970,N_9881);
and UO_872 (O_872,N_9931,N_9924);
and UO_873 (O_873,N_9850,N_9823);
and UO_874 (O_874,N_9924,N_9948);
or UO_875 (O_875,N_9817,N_9931);
and UO_876 (O_876,N_9837,N_9879);
nand UO_877 (O_877,N_9990,N_9943);
nor UO_878 (O_878,N_9833,N_9856);
nor UO_879 (O_879,N_9847,N_9912);
or UO_880 (O_880,N_9907,N_9920);
and UO_881 (O_881,N_9845,N_9837);
xor UO_882 (O_882,N_9847,N_9894);
and UO_883 (O_883,N_9902,N_9964);
nand UO_884 (O_884,N_9859,N_9814);
nand UO_885 (O_885,N_9986,N_9849);
or UO_886 (O_886,N_9822,N_9865);
nor UO_887 (O_887,N_9972,N_9825);
nor UO_888 (O_888,N_9826,N_9908);
nand UO_889 (O_889,N_9843,N_9874);
nand UO_890 (O_890,N_9881,N_9847);
nand UO_891 (O_891,N_9920,N_9838);
xnor UO_892 (O_892,N_9837,N_9964);
nor UO_893 (O_893,N_9803,N_9868);
nand UO_894 (O_894,N_9982,N_9997);
xor UO_895 (O_895,N_9834,N_9978);
nor UO_896 (O_896,N_9971,N_9927);
and UO_897 (O_897,N_9960,N_9966);
or UO_898 (O_898,N_9987,N_9830);
nor UO_899 (O_899,N_9854,N_9803);
and UO_900 (O_900,N_9963,N_9969);
and UO_901 (O_901,N_9940,N_9861);
or UO_902 (O_902,N_9877,N_9869);
nor UO_903 (O_903,N_9940,N_9845);
nor UO_904 (O_904,N_9916,N_9830);
xor UO_905 (O_905,N_9998,N_9818);
and UO_906 (O_906,N_9900,N_9883);
and UO_907 (O_907,N_9864,N_9943);
or UO_908 (O_908,N_9978,N_9873);
xor UO_909 (O_909,N_9913,N_9926);
nand UO_910 (O_910,N_9968,N_9820);
nand UO_911 (O_911,N_9937,N_9951);
and UO_912 (O_912,N_9837,N_9881);
xnor UO_913 (O_913,N_9938,N_9892);
nor UO_914 (O_914,N_9847,N_9987);
nor UO_915 (O_915,N_9845,N_9980);
and UO_916 (O_916,N_9817,N_9825);
or UO_917 (O_917,N_9963,N_9854);
or UO_918 (O_918,N_9917,N_9816);
nor UO_919 (O_919,N_9823,N_9964);
nor UO_920 (O_920,N_9968,N_9987);
xor UO_921 (O_921,N_9979,N_9976);
or UO_922 (O_922,N_9916,N_9909);
or UO_923 (O_923,N_9809,N_9812);
or UO_924 (O_924,N_9935,N_9952);
nor UO_925 (O_925,N_9914,N_9803);
and UO_926 (O_926,N_9875,N_9943);
nand UO_927 (O_927,N_9966,N_9969);
xor UO_928 (O_928,N_9912,N_9989);
nand UO_929 (O_929,N_9814,N_9884);
and UO_930 (O_930,N_9945,N_9903);
or UO_931 (O_931,N_9822,N_9867);
or UO_932 (O_932,N_9801,N_9987);
and UO_933 (O_933,N_9992,N_9880);
or UO_934 (O_934,N_9828,N_9843);
nand UO_935 (O_935,N_9996,N_9872);
or UO_936 (O_936,N_9807,N_9824);
and UO_937 (O_937,N_9864,N_9935);
and UO_938 (O_938,N_9970,N_9882);
or UO_939 (O_939,N_9965,N_9957);
and UO_940 (O_940,N_9834,N_9954);
and UO_941 (O_941,N_9946,N_9873);
and UO_942 (O_942,N_9942,N_9918);
xor UO_943 (O_943,N_9964,N_9829);
xnor UO_944 (O_944,N_9840,N_9826);
or UO_945 (O_945,N_9842,N_9974);
nand UO_946 (O_946,N_9922,N_9900);
and UO_947 (O_947,N_9866,N_9917);
and UO_948 (O_948,N_9955,N_9878);
or UO_949 (O_949,N_9977,N_9833);
nand UO_950 (O_950,N_9902,N_9946);
and UO_951 (O_951,N_9912,N_9894);
xnor UO_952 (O_952,N_9965,N_9933);
and UO_953 (O_953,N_9926,N_9861);
xnor UO_954 (O_954,N_9978,N_9906);
and UO_955 (O_955,N_9835,N_9839);
nand UO_956 (O_956,N_9949,N_9862);
nor UO_957 (O_957,N_9873,N_9815);
nand UO_958 (O_958,N_9949,N_9835);
xnor UO_959 (O_959,N_9827,N_9906);
nand UO_960 (O_960,N_9965,N_9822);
nor UO_961 (O_961,N_9862,N_9868);
nand UO_962 (O_962,N_9856,N_9823);
nand UO_963 (O_963,N_9811,N_9821);
and UO_964 (O_964,N_9847,N_9855);
nand UO_965 (O_965,N_9975,N_9974);
nand UO_966 (O_966,N_9864,N_9859);
nand UO_967 (O_967,N_9927,N_9998);
nand UO_968 (O_968,N_9818,N_9884);
nand UO_969 (O_969,N_9973,N_9834);
nand UO_970 (O_970,N_9983,N_9932);
xnor UO_971 (O_971,N_9822,N_9976);
xor UO_972 (O_972,N_9871,N_9982);
nor UO_973 (O_973,N_9858,N_9847);
or UO_974 (O_974,N_9997,N_9883);
nand UO_975 (O_975,N_9834,N_9877);
and UO_976 (O_976,N_9977,N_9986);
and UO_977 (O_977,N_9969,N_9953);
nor UO_978 (O_978,N_9927,N_9958);
nor UO_979 (O_979,N_9833,N_9875);
and UO_980 (O_980,N_9862,N_9954);
nor UO_981 (O_981,N_9871,N_9914);
nor UO_982 (O_982,N_9809,N_9957);
xnor UO_983 (O_983,N_9804,N_9810);
nand UO_984 (O_984,N_9939,N_9907);
or UO_985 (O_985,N_9922,N_9903);
and UO_986 (O_986,N_9825,N_9948);
or UO_987 (O_987,N_9974,N_9820);
nand UO_988 (O_988,N_9981,N_9864);
or UO_989 (O_989,N_9977,N_9859);
nand UO_990 (O_990,N_9975,N_9843);
nor UO_991 (O_991,N_9939,N_9915);
xor UO_992 (O_992,N_9802,N_9895);
and UO_993 (O_993,N_9882,N_9812);
nand UO_994 (O_994,N_9945,N_9844);
or UO_995 (O_995,N_9814,N_9800);
and UO_996 (O_996,N_9867,N_9814);
and UO_997 (O_997,N_9956,N_9816);
or UO_998 (O_998,N_9855,N_9978);
or UO_999 (O_999,N_9989,N_9873);
nand UO_1000 (O_1000,N_9882,N_9814);
nor UO_1001 (O_1001,N_9940,N_9976);
and UO_1002 (O_1002,N_9827,N_9897);
and UO_1003 (O_1003,N_9961,N_9966);
nand UO_1004 (O_1004,N_9984,N_9829);
nand UO_1005 (O_1005,N_9882,N_9851);
or UO_1006 (O_1006,N_9957,N_9961);
or UO_1007 (O_1007,N_9800,N_9962);
nor UO_1008 (O_1008,N_9899,N_9919);
nor UO_1009 (O_1009,N_9879,N_9959);
or UO_1010 (O_1010,N_9963,N_9900);
nor UO_1011 (O_1011,N_9962,N_9910);
nor UO_1012 (O_1012,N_9912,N_9829);
nor UO_1013 (O_1013,N_9893,N_9923);
nand UO_1014 (O_1014,N_9909,N_9923);
and UO_1015 (O_1015,N_9996,N_9957);
nand UO_1016 (O_1016,N_9871,N_9996);
xor UO_1017 (O_1017,N_9956,N_9911);
or UO_1018 (O_1018,N_9871,N_9948);
nand UO_1019 (O_1019,N_9838,N_9996);
nand UO_1020 (O_1020,N_9810,N_9955);
or UO_1021 (O_1021,N_9919,N_9978);
or UO_1022 (O_1022,N_9837,N_9939);
nor UO_1023 (O_1023,N_9842,N_9983);
or UO_1024 (O_1024,N_9937,N_9844);
xor UO_1025 (O_1025,N_9992,N_9967);
nor UO_1026 (O_1026,N_9927,N_9868);
and UO_1027 (O_1027,N_9959,N_9868);
and UO_1028 (O_1028,N_9931,N_9948);
xor UO_1029 (O_1029,N_9881,N_9813);
nor UO_1030 (O_1030,N_9949,N_9848);
and UO_1031 (O_1031,N_9968,N_9961);
nand UO_1032 (O_1032,N_9950,N_9840);
nor UO_1033 (O_1033,N_9893,N_9838);
nor UO_1034 (O_1034,N_9913,N_9898);
nand UO_1035 (O_1035,N_9978,N_9992);
xor UO_1036 (O_1036,N_9802,N_9833);
nor UO_1037 (O_1037,N_9872,N_9861);
nand UO_1038 (O_1038,N_9807,N_9847);
and UO_1039 (O_1039,N_9976,N_9922);
nand UO_1040 (O_1040,N_9938,N_9810);
or UO_1041 (O_1041,N_9856,N_9824);
nor UO_1042 (O_1042,N_9855,N_9999);
and UO_1043 (O_1043,N_9833,N_9910);
or UO_1044 (O_1044,N_9903,N_9835);
nand UO_1045 (O_1045,N_9994,N_9971);
and UO_1046 (O_1046,N_9937,N_9954);
or UO_1047 (O_1047,N_9998,N_9811);
nor UO_1048 (O_1048,N_9947,N_9952);
nand UO_1049 (O_1049,N_9963,N_9866);
or UO_1050 (O_1050,N_9886,N_9804);
nor UO_1051 (O_1051,N_9991,N_9890);
nand UO_1052 (O_1052,N_9855,N_9861);
and UO_1053 (O_1053,N_9951,N_9842);
xnor UO_1054 (O_1054,N_9943,N_9976);
nor UO_1055 (O_1055,N_9835,N_9990);
or UO_1056 (O_1056,N_9806,N_9970);
and UO_1057 (O_1057,N_9817,N_9991);
xnor UO_1058 (O_1058,N_9869,N_9823);
nor UO_1059 (O_1059,N_9921,N_9902);
or UO_1060 (O_1060,N_9898,N_9917);
and UO_1061 (O_1061,N_9859,N_9901);
nand UO_1062 (O_1062,N_9958,N_9960);
nor UO_1063 (O_1063,N_9992,N_9981);
or UO_1064 (O_1064,N_9832,N_9948);
nor UO_1065 (O_1065,N_9838,N_9900);
and UO_1066 (O_1066,N_9849,N_9868);
nor UO_1067 (O_1067,N_9983,N_9906);
nand UO_1068 (O_1068,N_9841,N_9958);
nand UO_1069 (O_1069,N_9928,N_9847);
nand UO_1070 (O_1070,N_9866,N_9927);
nand UO_1071 (O_1071,N_9816,N_9878);
or UO_1072 (O_1072,N_9928,N_9882);
or UO_1073 (O_1073,N_9990,N_9985);
or UO_1074 (O_1074,N_9985,N_9840);
nand UO_1075 (O_1075,N_9816,N_9965);
nand UO_1076 (O_1076,N_9813,N_9832);
nand UO_1077 (O_1077,N_9836,N_9944);
and UO_1078 (O_1078,N_9969,N_9975);
nor UO_1079 (O_1079,N_9852,N_9888);
nor UO_1080 (O_1080,N_9905,N_9803);
or UO_1081 (O_1081,N_9928,N_9941);
nand UO_1082 (O_1082,N_9981,N_9923);
or UO_1083 (O_1083,N_9944,N_9930);
and UO_1084 (O_1084,N_9903,N_9980);
or UO_1085 (O_1085,N_9838,N_9851);
nor UO_1086 (O_1086,N_9852,N_9885);
and UO_1087 (O_1087,N_9841,N_9956);
nor UO_1088 (O_1088,N_9964,N_9828);
nand UO_1089 (O_1089,N_9803,N_9948);
and UO_1090 (O_1090,N_9927,N_9930);
and UO_1091 (O_1091,N_9881,N_9967);
or UO_1092 (O_1092,N_9808,N_9959);
xor UO_1093 (O_1093,N_9945,N_9913);
or UO_1094 (O_1094,N_9959,N_9825);
nor UO_1095 (O_1095,N_9927,N_9887);
or UO_1096 (O_1096,N_9927,N_9991);
or UO_1097 (O_1097,N_9942,N_9904);
or UO_1098 (O_1098,N_9936,N_9950);
and UO_1099 (O_1099,N_9873,N_9962);
or UO_1100 (O_1100,N_9845,N_9834);
nor UO_1101 (O_1101,N_9832,N_9877);
or UO_1102 (O_1102,N_9837,N_9865);
nand UO_1103 (O_1103,N_9817,N_9999);
nand UO_1104 (O_1104,N_9856,N_9865);
or UO_1105 (O_1105,N_9842,N_9932);
nand UO_1106 (O_1106,N_9928,N_9817);
and UO_1107 (O_1107,N_9872,N_9881);
and UO_1108 (O_1108,N_9926,N_9849);
nand UO_1109 (O_1109,N_9880,N_9860);
and UO_1110 (O_1110,N_9903,N_9967);
nand UO_1111 (O_1111,N_9885,N_9998);
nor UO_1112 (O_1112,N_9959,N_9853);
nor UO_1113 (O_1113,N_9943,N_9977);
and UO_1114 (O_1114,N_9802,N_9898);
xor UO_1115 (O_1115,N_9893,N_9901);
nand UO_1116 (O_1116,N_9975,N_9973);
nand UO_1117 (O_1117,N_9835,N_9859);
nand UO_1118 (O_1118,N_9979,N_9859);
nor UO_1119 (O_1119,N_9977,N_9906);
nand UO_1120 (O_1120,N_9932,N_9826);
nand UO_1121 (O_1121,N_9968,N_9971);
or UO_1122 (O_1122,N_9839,N_9977);
nand UO_1123 (O_1123,N_9825,N_9918);
nand UO_1124 (O_1124,N_9954,N_9881);
or UO_1125 (O_1125,N_9885,N_9961);
and UO_1126 (O_1126,N_9808,N_9999);
xor UO_1127 (O_1127,N_9995,N_9859);
nand UO_1128 (O_1128,N_9903,N_9970);
or UO_1129 (O_1129,N_9833,N_9915);
nand UO_1130 (O_1130,N_9956,N_9811);
and UO_1131 (O_1131,N_9930,N_9874);
or UO_1132 (O_1132,N_9943,N_9958);
nor UO_1133 (O_1133,N_9945,N_9871);
xnor UO_1134 (O_1134,N_9850,N_9851);
xnor UO_1135 (O_1135,N_9983,N_9961);
nor UO_1136 (O_1136,N_9900,N_9913);
xor UO_1137 (O_1137,N_9832,N_9977);
nor UO_1138 (O_1138,N_9888,N_9980);
xnor UO_1139 (O_1139,N_9864,N_9911);
and UO_1140 (O_1140,N_9991,N_9929);
nand UO_1141 (O_1141,N_9905,N_9910);
or UO_1142 (O_1142,N_9891,N_9876);
or UO_1143 (O_1143,N_9909,N_9884);
and UO_1144 (O_1144,N_9960,N_9994);
or UO_1145 (O_1145,N_9820,N_9859);
nand UO_1146 (O_1146,N_9804,N_9978);
nor UO_1147 (O_1147,N_9955,N_9838);
xor UO_1148 (O_1148,N_9938,N_9877);
and UO_1149 (O_1149,N_9972,N_9969);
xor UO_1150 (O_1150,N_9900,N_9989);
and UO_1151 (O_1151,N_9985,N_9986);
xnor UO_1152 (O_1152,N_9925,N_9924);
nor UO_1153 (O_1153,N_9965,N_9998);
nand UO_1154 (O_1154,N_9904,N_9989);
nor UO_1155 (O_1155,N_9838,N_9983);
or UO_1156 (O_1156,N_9906,N_9803);
and UO_1157 (O_1157,N_9899,N_9904);
nand UO_1158 (O_1158,N_9902,N_9828);
nor UO_1159 (O_1159,N_9887,N_9934);
and UO_1160 (O_1160,N_9860,N_9846);
nor UO_1161 (O_1161,N_9971,N_9825);
or UO_1162 (O_1162,N_9999,N_9861);
and UO_1163 (O_1163,N_9833,N_9965);
and UO_1164 (O_1164,N_9938,N_9932);
and UO_1165 (O_1165,N_9810,N_9998);
nor UO_1166 (O_1166,N_9927,N_9886);
and UO_1167 (O_1167,N_9901,N_9924);
nor UO_1168 (O_1168,N_9803,N_9956);
nand UO_1169 (O_1169,N_9996,N_9945);
xnor UO_1170 (O_1170,N_9911,N_9893);
and UO_1171 (O_1171,N_9838,N_9967);
or UO_1172 (O_1172,N_9821,N_9815);
and UO_1173 (O_1173,N_9898,N_9954);
or UO_1174 (O_1174,N_9922,N_9823);
xor UO_1175 (O_1175,N_9816,N_9919);
and UO_1176 (O_1176,N_9896,N_9964);
nand UO_1177 (O_1177,N_9881,N_9979);
or UO_1178 (O_1178,N_9837,N_9902);
nor UO_1179 (O_1179,N_9904,N_9935);
nand UO_1180 (O_1180,N_9844,N_9837);
xnor UO_1181 (O_1181,N_9852,N_9813);
nand UO_1182 (O_1182,N_9819,N_9828);
nor UO_1183 (O_1183,N_9830,N_9932);
and UO_1184 (O_1184,N_9825,N_9992);
and UO_1185 (O_1185,N_9867,N_9810);
nand UO_1186 (O_1186,N_9973,N_9889);
nand UO_1187 (O_1187,N_9986,N_9866);
nor UO_1188 (O_1188,N_9889,N_9949);
nor UO_1189 (O_1189,N_9924,N_9894);
and UO_1190 (O_1190,N_9847,N_9985);
or UO_1191 (O_1191,N_9893,N_9899);
and UO_1192 (O_1192,N_9981,N_9891);
and UO_1193 (O_1193,N_9810,N_9986);
or UO_1194 (O_1194,N_9905,N_9916);
nor UO_1195 (O_1195,N_9877,N_9975);
and UO_1196 (O_1196,N_9997,N_9954);
nor UO_1197 (O_1197,N_9866,N_9994);
nand UO_1198 (O_1198,N_9806,N_9897);
nand UO_1199 (O_1199,N_9816,N_9908);
nor UO_1200 (O_1200,N_9825,N_9985);
nand UO_1201 (O_1201,N_9958,N_9934);
nand UO_1202 (O_1202,N_9956,N_9944);
nor UO_1203 (O_1203,N_9849,N_9981);
nand UO_1204 (O_1204,N_9821,N_9928);
and UO_1205 (O_1205,N_9992,N_9830);
and UO_1206 (O_1206,N_9981,N_9890);
nor UO_1207 (O_1207,N_9804,N_9953);
xnor UO_1208 (O_1208,N_9834,N_9869);
nor UO_1209 (O_1209,N_9997,N_9840);
nand UO_1210 (O_1210,N_9990,N_9918);
nand UO_1211 (O_1211,N_9988,N_9909);
nor UO_1212 (O_1212,N_9955,N_9983);
or UO_1213 (O_1213,N_9930,N_9868);
or UO_1214 (O_1214,N_9865,N_9825);
and UO_1215 (O_1215,N_9834,N_9841);
nand UO_1216 (O_1216,N_9824,N_9850);
nor UO_1217 (O_1217,N_9886,N_9900);
xor UO_1218 (O_1218,N_9826,N_9912);
or UO_1219 (O_1219,N_9825,N_9947);
and UO_1220 (O_1220,N_9820,N_9966);
or UO_1221 (O_1221,N_9859,N_9960);
xnor UO_1222 (O_1222,N_9884,N_9967);
or UO_1223 (O_1223,N_9900,N_9822);
or UO_1224 (O_1224,N_9849,N_9933);
nor UO_1225 (O_1225,N_9971,N_9818);
nor UO_1226 (O_1226,N_9901,N_9878);
nand UO_1227 (O_1227,N_9811,N_9992);
or UO_1228 (O_1228,N_9905,N_9873);
and UO_1229 (O_1229,N_9894,N_9873);
or UO_1230 (O_1230,N_9863,N_9940);
nand UO_1231 (O_1231,N_9898,N_9874);
and UO_1232 (O_1232,N_9906,N_9858);
nor UO_1233 (O_1233,N_9840,N_9945);
and UO_1234 (O_1234,N_9927,N_9963);
and UO_1235 (O_1235,N_9998,N_9956);
nand UO_1236 (O_1236,N_9945,N_9886);
nor UO_1237 (O_1237,N_9946,N_9866);
and UO_1238 (O_1238,N_9818,N_9982);
or UO_1239 (O_1239,N_9813,N_9942);
xor UO_1240 (O_1240,N_9891,N_9821);
and UO_1241 (O_1241,N_9902,N_9936);
nor UO_1242 (O_1242,N_9888,N_9820);
and UO_1243 (O_1243,N_9820,N_9863);
nor UO_1244 (O_1244,N_9886,N_9847);
xnor UO_1245 (O_1245,N_9948,N_9976);
and UO_1246 (O_1246,N_9947,N_9963);
xnor UO_1247 (O_1247,N_9842,N_9911);
nand UO_1248 (O_1248,N_9903,N_9885);
xor UO_1249 (O_1249,N_9993,N_9820);
nand UO_1250 (O_1250,N_9838,N_9944);
nor UO_1251 (O_1251,N_9837,N_9869);
and UO_1252 (O_1252,N_9823,N_9975);
or UO_1253 (O_1253,N_9928,N_9902);
nand UO_1254 (O_1254,N_9817,N_9806);
or UO_1255 (O_1255,N_9852,N_9911);
nand UO_1256 (O_1256,N_9995,N_9966);
nand UO_1257 (O_1257,N_9806,N_9847);
and UO_1258 (O_1258,N_9943,N_9981);
nand UO_1259 (O_1259,N_9869,N_9890);
nor UO_1260 (O_1260,N_9953,N_9803);
or UO_1261 (O_1261,N_9945,N_9810);
and UO_1262 (O_1262,N_9851,N_9901);
or UO_1263 (O_1263,N_9959,N_9836);
xnor UO_1264 (O_1264,N_9981,N_9873);
or UO_1265 (O_1265,N_9896,N_9885);
or UO_1266 (O_1266,N_9988,N_9962);
and UO_1267 (O_1267,N_9955,N_9890);
and UO_1268 (O_1268,N_9985,N_9812);
nand UO_1269 (O_1269,N_9907,N_9917);
nor UO_1270 (O_1270,N_9936,N_9906);
nand UO_1271 (O_1271,N_9948,N_9865);
nand UO_1272 (O_1272,N_9963,N_9911);
or UO_1273 (O_1273,N_9954,N_9814);
nor UO_1274 (O_1274,N_9993,N_9976);
xnor UO_1275 (O_1275,N_9971,N_9814);
nor UO_1276 (O_1276,N_9891,N_9845);
or UO_1277 (O_1277,N_9916,N_9823);
or UO_1278 (O_1278,N_9927,N_9870);
xor UO_1279 (O_1279,N_9958,N_9956);
or UO_1280 (O_1280,N_9908,N_9968);
xor UO_1281 (O_1281,N_9872,N_9877);
and UO_1282 (O_1282,N_9981,N_9819);
and UO_1283 (O_1283,N_9945,N_9926);
nor UO_1284 (O_1284,N_9807,N_9968);
nand UO_1285 (O_1285,N_9994,N_9859);
nor UO_1286 (O_1286,N_9934,N_9897);
or UO_1287 (O_1287,N_9981,N_9999);
nand UO_1288 (O_1288,N_9868,N_9916);
nor UO_1289 (O_1289,N_9825,N_9886);
nor UO_1290 (O_1290,N_9990,N_9809);
and UO_1291 (O_1291,N_9878,N_9830);
and UO_1292 (O_1292,N_9861,N_9811);
nand UO_1293 (O_1293,N_9821,N_9953);
xnor UO_1294 (O_1294,N_9816,N_9907);
nand UO_1295 (O_1295,N_9930,N_9880);
and UO_1296 (O_1296,N_9954,N_9932);
and UO_1297 (O_1297,N_9874,N_9812);
and UO_1298 (O_1298,N_9866,N_9852);
nor UO_1299 (O_1299,N_9839,N_9985);
nand UO_1300 (O_1300,N_9822,N_9880);
xor UO_1301 (O_1301,N_9876,N_9934);
nand UO_1302 (O_1302,N_9826,N_9859);
xnor UO_1303 (O_1303,N_9895,N_9833);
nor UO_1304 (O_1304,N_9953,N_9864);
and UO_1305 (O_1305,N_9985,N_9913);
and UO_1306 (O_1306,N_9935,N_9918);
xnor UO_1307 (O_1307,N_9893,N_9880);
nor UO_1308 (O_1308,N_9958,N_9987);
nor UO_1309 (O_1309,N_9818,N_9951);
and UO_1310 (O_1310,N_9806,N_9842);
and UO_1311 (O_1311,N_9963,N_9982);
nor UO_1312 (O_1312,N_9853,N_9809);
or UO_1313 (O_1313,N_9955,N_9961);
nand UO_1314 (O_1314,N_9918,N_9955);
or UO_1315 (O_1315,N_9865,N_9878);
and UO_1316 (O_1316,N_9877,N_9867);
nor UO_1317 (O_1317,N_9958,N_9904);
nor UO_1318 (O_1318,N_9863,N_9898);
xor UO_1319 (O_1319,N_9842,N_9800);
nand UO_1320 (O_1320,N_9888,N_9944);
nor UO_1321 (O_1321,N_9970,N_9822);
nand UO_1322 (O_1322,N_9899,N_9941);
or UO_1323 (O_1323,N_9882,N_9994);
and UO_1324 (O_1324,N_9976,N_9825);
or UO_1325 (O_1325,N_9891,N_9952);
or UO_1326 (O_1326,N_9909,N_9919);
xor UO_1327 (O_1327,N_9954,N_9891);
nor UO_1328 (O_1328,N_9841,N_9867);
nor UO_1329 (O_1329,N_9930,N_9941);
xor UO_1330 (O_1330,N_9825,N_9847);
nor UO_1331 (O_1331,N_9852,N_9923);
and UO_1332 (O_1332,N_9970,N_9980);
nor UO_1333 (O_1333,N_9816,N_9880);
or UO_1334 (O_1334,N_9872,N_9983);
or UO_1335 (O_1335,N_9931,N_9896);
and UO_1336 (O_1336,N_9822,N_9914);
nor UO_1337 (O_1337,N_9975,N_9892);
nor UO_1338 (O_1338,N_9826,N_9858);
or UO_1339 (O_1339,N_9805,N_9850);
xor UO_1340 (O_1340,N_9955,N_9891);
nor UO_1341 (O_1341,N_9847,N_9901);
nand UO_1342 (O_1342,N_9901,N_9823);
nand UO_1343 (O_1343,N_9973,N_9935);
or UO_1344 (O_1344,N_9883,N_9919);
and UO_1345 (O_1345,N_9912,N_9963);
nand UO_1346 (O_1346,N_9921,N_9935);
and UO_1347 (O_1347,N_9912,N_9857);
or UO_1348 (O_1348,N_9829,N_9998);
or UO_1349 (O_1349,N_9956,N_9908);
or UO_1350 (O_1350,N_9856,N_9888);
nand UO_1351 (O_1351,N_9929,N_9912);
or UO_1352 (O_1352,N_9947,N_9918);
nand UO_1353 (O_1353,N_9926,N_9800);
and UO_1354 (O_1354,N_9947,N_9879);
xor UO_1355 (O_1355,N_9855,N_9868);
and UO_1356 (O_1356,N_9961,N_9924);
xnor UO_1357 (O_1357,N_9861,N_9994);
and UO_1358 (O_1358,N_9968,N_9897);
and UO_1359 (O_1359,N_9943,N_9919);
nand UO_1360 (O_1360,N_9969,N_9940);
nand UO_1361 (O_1361,N_9858,N_9913);
nand UO_1362 (O_1362,N_9966,N_9893);
and UO_1363 (O_1363,N_9988,N_9859);
nor UO_1364 (O_1364,N_9836,N_9968);
xor UO_1365 (O_1365,N_9830,N_9872);
or UO_1366 (O_1366,N_9842,N_9848);
nor UO_1367 (O_1367,N_9994,N_9818);
nor UO_1368 (O_1368,N_9866,N_9820);
and UO_1369 (O_1369,N_9935,N_9841);
nand UO_1370 (O_1370,N_9971,N_9947);
nand UO_1371 (O_1371,N_9987,N_9983);
or UO_1372 (O_1372,N_9950,N_9957);
nor UO_1373 (O_1373,N_9995,N_9816);
nand UO_1374 (O_1374,N_9984,N_9988);
or UO_1375 (O_1375,N_9875,N_9880);
nor UO_1376 (O_1376,N_9985,N_9861);
and UO_1377 (O_1377,N_9964,N_9822);
nand UO_1378 (O_1378,N_9868,N_9935);
nand UO_1379 (O_1379,N_9905,N_9963);
and UO_1380 (O_1380,N_9900,N_9905);
nor UO_1381 (O_1381,N_9929,N_9878);
nor UO_1382 (O_1382,N_9976,N_9999);
or UO_1383 (O_1383,N_9875,N_9835);
nand UO_1384 (O_1384,N_9868,N_9824);
nor UO_1385 (O_1385,N_9837,N_9866);
or UO_1386 (O_1386,N_9892,N_9910);
xor UO_1387 (O_1387,N_9842,N_9956);
xor UO_1388 (O_1388,N_9971,N_9966);
and UO_1389 (O_1389,N_9958,N_9803);
and UO_1390 (O_1390,N_9986,N_9816);
nand UO_1391 (O_1391,N_9887,N_9975);
nor UO_1392 (O_1392,N_9901,N_9912);
or UO_1393 (O_1393,N_9971,N_9991);
and UO_1394 (O_1394,N_9890,N_9992);
nor UO_1395 (O_1395,N_9994,N_9939);
nand UO_1396 (O_1396,N_9903,N_9906);
nand UO_1397 (O_1397,N_9957,N_9920);
nor UO_1398 (O_1398,N_9989,N_9840);
xor UO_1399 (O_1399,N_9840,N_9966);
or UO_1400 (O_1400,N_9844,N_9985);
xor UO_1401 (O_1401,N_9916,N_9931);
nor UO_1402 (O_1402,N_9871,N_9828);
xnor UO_1403 (O_1403,N_9981,N_9935);
nor UO_1404 (O_1404,N_9975,N_9845);
xnor UO_1405 (O_1405,N_9940,N_9981);
xnor UO_1406 (O_1406,N_9997,N_9863);
nor UO_1407 (O_1407,N_9981,N_9894);
and UO_1408 (O_1408,N_9833,N_9908);
and UO_1409 (O_1409,N_9847,N_9868);
nand UO_1410 (O_1410,N_9943,N_9800);
nand UO_1411 (O_1411,N_9891,N_9811);
or UO_1412 (O_1412,N_9868,N_9851);
nand UO_1413 (O_1413,N_9947,N_9948);
nand UO_1414 (O_1414,N_9901,N_9850);
or UO_1415 (O_1415,N_9894,N_9871);
nor UO_1416 (O_1416,N_9987,N_9906);
and UO_1417 (O_1417,N_9811,N_9822);
and UO_1418 (O_1418,N_9813,N_9937);
nor UO_1419 (O_1419,N_9865,N_9870);
and UO_1420 (O_1420,N_9856,N_9977);
nor UO_1421 (O_1421,N_9878,N_9939);
nand UO_1422 (O_1422,N_9944,N_9988);
and UO_1423 (O_1423,N_9939,N_9949);
nor UO_1424 (O_1424,N_9950,N_9814);
nor UO_1425 (O_1425,N_9920,N_9837);
and UO_1426 (O_1426,N_9945,N_9958);
nand UO_1427 (O_1427,N_9966,N_9959);
nand UO_1428 (O_1428,N_9872,N_9998);
or UO_1429 (O_1429,N_9831,N_9872);
nand UO_1430 (O_1430,N_9882,N_9877);
xnor UO_1431 (O_1431,N_9954,N_9905);
or UO_1432 (O_1432,N_9931,N_9950);
and UO_1433 (O_1433,N_9992,N_9995);
nand UO_1434 (O_1434,N_9867,N_9838);
nand UO_1435 (O_1435,N_9852,N_9858);
nor UO_1436 (O_1436,N_9869,N_9821);
or UO_1437 (O_1437,N_9809,N_9966);
nand UO_1438 (O_1438,N_9866,N_9886);
nand UO_1439 (O_1439,N_9812,N_9962);
or UO_1440 (O_1440,N_9947,N_9821);
or UO_1441 (O_1441,N_9860,N_9947);
nor UO_1442 (O_1442,N_9887,N_9877);
or UO_1443 (O_1443,N_9902,N_9939);
or UO_1444 (O_1444,N_9822,N_9903);
nor UO_1445 (O_1445,N_9896,N_9986);
nor UO_1446 (O_1446,N_9922,N_9887);
nand UO_1447 (O_1447,N_9942,N_9856);
or UO_1448 (O_1448,N_9924,N_9809);
nand UO_1449 (O_1449,N_9959,N_9953);
and UO_1450 (O_1450,N_9971,N_9920);
nand UO_1451 (O_1451,N_9960,N_9990);
and UO_1452 (O_1452,N_9926,N_9998);
nand UO_1453 (O_1453,N_9919,N_9996);
and UO_1454 (O_1454,N_9996,N_9933);
and UO_1455 (O_1455,N_9964,N_9809);
or UO_1456 (O_1456,N_9982,N_9999);
and UO_1457 (O_1457,N_9953,N_9944);
or UO_1458 (O_1458,N_9872,N_9883);
nor UO_1459 (O_1459,N_9945,N_9934);
nor UO_1460 (O_1460,N_9901,N_9915);
nand UO_1461 (O_1461,N_9940,N_9915);
nor UO_1462 (O_1462,N_9835,N_9870);
and UO_1463 (O_1463,N_9825,N_9927);
or UO_1464 (O_1464,N_9964,N_9854);
and UO_1465 (O_1465,N_9973,N_9864);
nor UO_1466 (O_1466,N_9965,N_9857);
or UO_1467 (O_1467,N_9844,N_9911);
nor UO_1468 (O_1468,N_9883,N_9991);
and UO_1469 (O_1469,N_9983,N_9993);
and UO_1470 (O_1470,N_9907,N_9919);
and UO_1471 (O_1471,N_9979,N_9946);
nand UO_1472 (O_1472,N_9926,N_9949);
nand UO_1473 (O_1473,N_9952,N_9814);
nand UO_1474 (O_1474,N_9929,N_9996);
nor UO_1475 (O_1475,N_9983,N_9869);
or UO_1476 (O_1476,N_9834,N_9926);
nand UO_1477 (O_1477,N_9983,N_9996);
nand UO_1478 (O_1478,N_9963,N_9939);
and UO_1479 (O_1479,N_9926,N_9873);
or UO_1480 (O_1480,N_9885,N_9822);
nand UO_1481 (O_1481,N_9935,N_9855);
and UO_1482 (O_1482,N_9978,N_9963);
and UO_1483 (O_1483,N_9934,N_9840);
nand UO_1484 (O_1484,N_9806,N_9968);
nor UO_1485 (O_1485,N_9898,N_9897);
nand UO_1486 (O_1486,N_9836,N_9915);
nor UO_1487 (O_1487,N_9967,N_9840);
or UO_1488 (O_1488,N_9975,N_9920);
xor UO_1489 (O_1489,N_9905,N_9908);
nor UO_1490 (O_1490,N_9923,N_9878);
or UO_1491 (O_1491,N_9836,N_9977);
xor UO_1492 (O_1492,N_9924,N_9877);
nor UO_1493 (O_1493,N_9886,N_9870);
nand UO_1494 (O_1494,N_9864,N_9840);
nor UO_1495 (O_1495,N_9928,N_9810);
or UO_1496 (O_1496,N_9925,N_9803);
or UO_1497 (O_1497,N_9850,N_9856);
or UO_1498 (O_1498,N_9864,N_9806);
and UO_1499 (O_1499,N_9927,N_9982);
endmodule