module basic_1500_15000_2000_5_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_727,In_78);
nor U1 (N_1,In_1040,In_1055);
or U2 (N_2,In_598,In_620);
nand U3 (N_3,In_1098,In_1095);
and U4 (N_4,In_1247,In_130);
or U5 (N_5,In_1433,In_663);
or U6 (N_6,In_1071,In_1326);
nor U7 (N_7,In_329,In_760);
nor U8 (N_8,In_441,In_1005);
and U9 (N_9,In_770,In_1147);
nor U10 (N_10,In_761,In_84);
and U11 (N_11,In_641,In_1394);
nand U12 (N_12,In_1232,In_1466);
and U13 (N_13,In_605,In_37);
nor U14 (N_14,In_785,In_731);
nand U15 (N_15,In_29,In_295);
nor U16 (N_16,In_435,In_645);
and U17 (N_17,In_430,In_553);
nor U18 (N_18,In_1367,In_1408);
nand U19 (N_19,In_610,In_600);
and U20 (N_20,In_163,In_1180);
nand U21 (N_21,In_585,In_956);
or U22 (N_22,In_524,In_776);
nand U23 (N_23,In_642,In_789);
nor U24 (N_24,In_1077,In_1036);
and U25 (N_25,In_807,In_176);
or U26 (N_26,In_1245,In_955);
nor U27 (N_27,In_1457,In_380);
nand U28 (N_28,In_1151,In_570);
or U29 (N_29,In_364,In_1415);
or U30 (N_30,In_1134,In_243);
and U31 (N_31,In_710,In_1474);
and U32 (N_32,In_1109,In_285);
nor U33 (N_33,In_521,In_1168);
or U34 (N_34,In_816,In_1118);
or U35 (N_35,In_1460,In_1385);
nor U36 (N_36,In_874,In_260);
or U37 (N_37,In_103,In_1291);
nand U38 (N_38,In_879,In_766);
nor U39 (N_39,In_1099,In_274);
nand U40 (N_40,In_395,In_0);
and U41 (N_41,In_1398,In_286);
nand U42 (N_42,In_1288,In_1403);
nor U43 (N_43,In_1091,In_94);
or U44 (N_44,In_1366,In_7);
or U45 (N_45,In_1174,In_903);
nand U46 (N_46,In_520,In_5);
nor U47 (N_47,In_1268,In_1484);
and U48 (N_48,In_142,In_82);
nand U49 (N_49,In_1226,In_337);
nand U50 (N_50,In_222,In_530);
or U51 (N_51,In_930,In_450);
or U52 (N_52,In_999,In_775);
xor U53 (N_53,In_996,In_1271);
nor U54 (N_54,In_166,In_33);
and U55 (N_55,In_681,In_895);
or U56 (N_56,In_518,In_1383);
nor U57 (N_57,In_783,In_1315);
nor U58 (N_58,In_549,In_252);
or U59 (N_59,In_608,In_92);
nand U60 (N_60,In_348,In_59);
nor U61 (N_61,In_1356,In_250);
nand U62 (N_62,In_42,In_146);
and U63 (N_63,In_229,In_237);
nor U64 (N_64,In_793,In_193);
or U65 (N_65,In_230,In_1434);
or U66 (N_66,In_1453,In_1186);
or U67 (N_67,In_577,In_419);
or U68 (N_68,In_523,In_1331);
or U69 (N_69,In_898,In_1402);
or U70 (N_70,In_1250,In_343);
or U71 (N_71,In_556,In_1397);
and U72 (N_72,In_137,In_1489);
xnor U73 (N_73,In_601,In_110);
nor U74 (N_74,In_881,In_904);
and U75 (N_75,In_847,In_1208);
and U76 (N_76,In_932,In_648);
nand U77 (N_77,In_1204,In_637);
and U78 (N_78,In_2,In_519);
nor U79 (N_79,In_402,In_806);
nor U80 (N_80,In_1262,In_1035);
or U81 (N_81,In_1479,In_1449);
nor U82 (N_82,In_661,In_1308);
or U83 (N_83,In_671,In_1155);
nor U84 (N_84,In_496,In_583);
and U85 (N_85,In_13,In_246);
nand U86 (N_86,In_957,In_236);
and U87 (N_87,In_694,In_581);
or U88 (N_88,In_880,In_207);
nor U89 (N_89,In_1088,In_1381);
nand U90 (N_90,In_108,In_715);
and U91 (N_91,In_1336,In_1401);
and U92 (N_92,In_315,In_960);
nand U93 (N_93,In_1199,In_1297);
nand U94 (N_94,In_686,In_370);
nand U95 (N_95,In_249,In_1202);
nor U96 (N_96,In_862,In_1217);
nand U97 (N_97,In_1357,In_1476);
nor U98 (N_98,In_340,In_1253);
nor U99 (N_99,In_220,In_1019);
and U100 (N_100,In_836,In_358);
and U101 (N_101,In_772,In_414);
or U102 (N_102,In_672,In_309);
or U103 (N_103,In_1216,In_449);
nor U104 (N_104,In_385,In_680);
or U105 (N_105,In_532,In_1473);
and U106 (N_106,In_1221,In_1239);
nand U107 (N_107,In_1349,In_339);
and U108 (N_108,In_389,In_938);
or U109 (N_109,In_184,In_1122);
or U110 (N_110,In_203,In_80);
nand U111 (N_111,In_51,In_1079);
or U112 (N_112,In_363,In_1094);
nor U113 (N_113,In_1017,In_1175);
or U114 (N_114,In_354,In_705);
or U115 (N_115,In_1156,In_20);
nor U116 (N_116,In_704,In_526);
nor U117 (N_117,In_690,In_1465);
nand U118 (N_118,In_472,In_1007);
nand U119 (N_119,In_408,In_1126);
or U120 (N_120,In_683,In_452);
nor U121 (N_121,In_1264,In_1317);
nand U122 (N_122,In_1441,In_1076);
nor U123 (N_123,In_838,In_1013);
and U124 (N_124,In_759,In_1051);
nor U125 (N_125,In_390,In_1057);
nand U126 (N_126,In_1205,In_355);
or U127 (N_127,In_817,In_729);
and U128 (N_128,In_1439,In_706);
and U129 (N_129,In_1407,In_561);
or U130 (N_130,In_1133,In_3);
and U131 (N_131,In_1306,In_170);
nor U132 (N_132,In_225,In_811);
or U133 (N_133,In_349,In_1298);
and U134 (N_134,In_1000,In_1455);
nand U135 (N_135,In_1294,In_959);
and U136 (N_136,In_629,In_757);
and U137 (N_137,In_60,In_1060);
nand U138 (N_138,In_1283,In_981);
nand U139 (N_139,In_748,In_1376);
nor U140 (N_140,In_1259,In_311);
or U141 (N_141,In_739,In_1285);
nor U142 (N_142,In_937,In_278);
or U143 (N_143,In_599,In_201);
nor U144 (N_144,In_702,In_335);
or U145 (N_145,In_745,In_308);
or U146 (N_146,In_427,In_292);
nand U147 (N_147,In_1404,In_1072);
nor U148 (N_148,In_346,In_1364);
nand U149 (N_149,In_1260,In_438);
nor U150 (N_150,In_1276,In_56);
nand U151 (N_151,In_1018,In_1481);
and U152 (N_152,In_47,In_1448);
nor U153 (N_153,In_314,In_813);
nand U154 (N_154,In_1102,In_352);
nand U155 (N_155,In_91,In_187);
or U156 (N_156,In_651,In_525);
and U157 (N_157,In_474,In_189);
or U158 (N_158,In_1486,In_998);
nand U159 (N_159,In_1480,In_624);
or U160 (N_160,In_1379,In_49);
or U161 (N_161,In_801,In_782);
and U162 (N_162,In_1142,In_1444);
nor U163 (N_163,In_812,In_302);
or U164 (N_164,In_897,In_734);
nand U165 (N_165,In_963,In_635);
and U166 (N_166,In_587,In_386);
nor U167 (N_167,In_361,In_1209);
and U168 (N_168,In_1395,In_821);
nand U169 (N_169,In_893,In_799);
nand U170 (N_170,In_1496,In_1277);
nand U171 (N_171,In_1119,In_842);
and U172 (N_172,In_717,In_948);
or U173 (N_173,In_784,In_1124);
nor U174 (N_174,In_304,In_1422);
or U175 (N_175,In_463,In_915);
nand U176 (N_176,In_973,In_923);
nand U177 (N_177,In_211,In_462);
nand U178 (N_178,In_1413,In_646);
nand U179 (N_179,In_477,In_269);
or U180 (N_180,In_318,In_1137);
and U181 (N_181,In_120,In_437);
or U182 (N_182,In_1074,In_1488);
or U183 (N_183,In_535,In_136);
or U184 (N_184,In_30,In_953);
nand U185 (N_185,In_484,In_241);
or U186 (N_186,In_968,In_885);
nand U187 (N_187,In_822,In_928);
or U188 (N_188,In_1330,In_855);
nor U189 (N_189,In_351,In_1117);
nor U190 (N_190,In_1189,In_1140);
and U191 (N_191,In_1256,In_453);
nor U192 (N_192,In_342,In_721);
nor U193 (N_193,In_510,In_418);
nand U194 (N_194,In_367,In_962);
nor U195 (N_195,In_1445,In_678);
nand U196 (N_196,In_911,In_765);
and U197 (N_197,In_551,In_1046);
and U198 (N_198,In_1131,In_1062);
nor U199 (N_199,In_1196,In_53);
nand U200 (N_200,In_539,In_173);
or U201 (N_201,In_492,In_926);
and U202 (N_202,In_373,In_615);
nand U203 (N_203,In_567,In_144);
or U204 (N_204,In_914,In_270);
and U205 (N_205,In_448,In_735);
and U206 (N_206,In_147,In_1301);
nor U207 (N_207,In_1,In_612);
and U208 (N_208,In_1049,In_1375);
or U209 (N_209,In_1390,In_1108);
or U210 (N_210,In_1103,In_117);
nand U211 (N_211,In_906,In_1121);
nand U212 (N_212,In_1396,In_1083);
nand U213 (N_213,In_336,In_190);
or U214 (N_214,In_1106,In_1426);
nand U215 (N_215,In_98,In_954);
and U216 (N_216,In_1058,In_638);
or U217 (N_217,In_493,In_113);
xnor U218 (N_218,In_1206,In_436);
or U219 (N_219,In_22,In_1468);
or U220 (N_220,In_210,In_649);
nor U221 (N_221,In_1052,In_1311);
or U222 (N_222,In_212,In_974);
and U223 (N_223,In_1210,In_242);
nand U224 (N_224,In_321,In_296);
nor U225 (N_225,In_72,In_1258);
or U226 (N_226,In_899,In_548);
and U227 (N_227,In_623,In_1352);
or U228 (N_228,In_596,In_506);
nor U229 (N_229,In_997,In_1257);
or U230 (N_230,In_1010,In_1469);
or U231 (N_231,In_1490,In_133);
nor U232 (N_232,In_415,In_653);
nor U233 (N_233,In_982,In_347);
nand U234 (N_234,In_26,In_711);
nor U235 (N_235,In_413,In_79);
or U236 (N_236,In_559,In_67);
nor U237 (N_237,In_1037,In_21);
and U238 (N_238,In_140,In_1386);
and U239 (N_239,In_753,In_513);
and U240 (N_240,In_1167,In_1414);
or U241 (N_241,In_1327,In_540);
xor U242 (N_242,In_1201,In_543);
nand U243 (N_243,In_494,In_1370);
nand U244 (N_244,In_407,In_1345);
and U245 (N_245,In_165,In_428);
xnor U246 (N_246,In_1472,In_1498);
nand U247 (N_247,In_1190,In_57);
nand U248 (N_248,In_316,In_196);
and U249 (N_249,In_993,In_66);
and U250 (N_250,In_1358,In_95);
and U251 (N_251,In_183,In_970);
or U252 (N_252,In_1170,In_719);
nand U253 (N_253,In_485,In_1430);
xor U254 (N_254,In_618,In_823);
nand U255 (N_255,In_1406,In_185);
nor U256 (N_256,In_1361,In_1184);
and U257 (N_257,In_1123,In_353);
or U258 (N_258,In_383,In_1194);
nor U259 (N_259,In_394,In_1373);
and U260 (N_260,In_359,In_1063);
and U261 (N_261,In_668,In_289);
nor U262 (N_262,In_422,In_186);
nand U263 (N_263,In_856,In_247);
or U264 (N_264,In_476,In_268);
nor U265 (N_265,In_1159,In_1371);
or U266 (N_266,In_798,In_773);
and U267 (N_267,In_473,In_172);
nand U268 (N_268,In_168,In_1418);
or U269 (N_269,In_868,In_810);
and U270 (N_270,In_376,In_1387);
and U271 (N_271,In_1462,In_1176);
nor U272 (N_272,In_611,In_381);
and U273 (N_273,In_143,In_374);
or U274 (N_274,In_1061,In_1112);
xor U275 (N_275,In_416,In_490);
nand U276 (N_276,In_1319,In_1233);
or U277 (N_277,In_1429,In_213);
and U278 (N_278,In_1016,In_1127);
nand U279 (N_279,In_257,In_1200);
and U280 (N_280,In_554,In_1321);
or U281 (N_281,In_275,In_112);
and U282 (N_282,In_674,In_504);
and U283 (N_283,In_1343,In_126);
nand U284 (N_284,In_1038,In_277);
nand U285 (N_285,In_978,In_1014);
nor U286 (N_286,In_486,In_658);
nor U287 (N_287,In_946,In_1041);
nor U288 (N_288,In_1084,In_870);
nand U289 (N_289,In_182,In_1382);
nor U290 (N_290,In_118,In_896);
nor U291 (N_291,In_215,In_1341);
or U292 (N_292,In_319,In_1483);
nor U293 (N_293,In_890,In_105);
nor U294 (N_294,In_1064,In_1097);
or U295 (N_295,In_752,In_410);
nand U296 (N_296,In_68,In_746);
and U297 (N_297,In_1353,In_224);
nor U298 (N_298,In_457,In_440);
or U299 (N_299,In_259,In_1138);
nor U300 (N_300,In_1146,In_1089);
or U301 (N_301,In_104,In_167);
or U302 (N_302,In_876,In_1065);
and U303 (N_303,In_546,In_487);
and U304 (N_304,In_1183,In_708);
nor U305 (N_305,In_254,In_517);
nand U306 (N_306,In_1478,In_550);
or U307 (N_307,In_564,In_664);
nand U308 (N_308,In_1365,In_204);
nand U309 (N_309,In_1125,In_827);
and U310 (N_310,In_828,In_657);
and U311 (N_311,In_344,In_887);
nand U312 (N_312,In_279,In_50);
and U313 (N_313,In_912,In_209);
nor U314 (N_314,In_451,In_584);
and U315 (N_315,In_479,In_326);
nand U316 (N_316,In_423,In_1048);
and U317 (N_317,In_58,In_1244);
xor U318 (N_318,In_387,In_61);
and U319 (N_319,In_872,In_818);
or U320 (N_320,In_994,In_1399);
or U321 (N_321,In_826,In_1320);
and U322 (N_322,In_659,In_310);
nor U323 (N_323,In_294,In_677);
nand U324 (N_324,In_850,In_952);
nor U325 (N_325,In_399,In_1164);
nor U326 (N_326,In_161,In_465);
or U327 (N_327,In_398,In_155);
nand U328 (N_328,In_1464,In_431);
nand U329 (N_329,In_724,In_256);
nor U330 (N_330,In_421,In_1056);
or U331 (N_331,In_1001,In_778);
nand U332 (N_332,In_569,In_1192);
nor U333 (N_333,In_541,In_709);
nand U334 (N_334,In_71,In_616);
nand U335 (N_335,In_1181,In_18);
and U336 (N_336,In_1093,In_625);
or U337 (N_337,In_566,In_1458);
nor U338 (N_338,In_676,In_1372);
nor U339 (N_339,In_508,In_1463);
nand U340 (N_340,In_135,In_273);
nand U341 (N_341,In_334,In_1417);
and U342 (N_342,In_594,In_714);
or U343 (N_343,In_1020,In_258);
nand U344 (N_344,In_40,In_35);
or U345 (N_345,In_755,In_325);
and U346 (N_346,In_1274,In_1389);
nand U347 (N_347,In_889,In_634);
nor U348 (N_348,In_245,In_73);
or U349 (N_349,In_1293,In_1437);
or U350 (N_350,In_894,In_244);
nor U351 (N_351,In_927,In_89);
or U352 (N_352,In_803,In_1154);
nand U353 (N_353,In_533,In_1286);
nor U354 (N_354,In_703,In_820);
and U355 (N_355,In_164,In_497);
nand U356 (N_356,In_1350,In_1053);
or U357 (N_357,In_461,In_1235);
nand U358 (N_358,In_301,In_1270);
xnor U359 (N_359,In_684,In_439);
nor U360 (N_360,In_1114,In_281);
or U361 (N_361,In_1113,In_830);
nand U362 (N_362,In_988,In_454);
nor U363 (N_363,In_129,In_1299);
and U364 (N_364,In_1432,In_192);
and U365 (N_365,In_512,In_1169);
nor U366 (N_366,In_1185,In_432);
nor U367 (N_367,In_299,In_795);
nand U368 (N_368,In_666,In_65);
nand U369 (N_369,In_1494,In_989);
nand U370 (N_370,In_1220,In_580);
nor U371 (N_371,In_177,In_1165);
and U372 (N_372,In_206,In_633);
nand U373 (N_373,In_216,In_43);
and U374 (N_374,In_1360,In_97);
and U375 (N_375,In_1130,In_1380);
and U376 (N_376,In_1228,In_701);
or U377 (N_377,In_323,In_1024);
nand U378 (N_378,In_1369,In_1182);
nor U379 (N_379,In_1105,In_725);
and U380 (N_380,In_471,In_867);
or U381 (N_381,In_458,In_698);
or U382 (N_382,In_647,In_1028);
or U383 (N_383,In_986,In_1163);
nor U384 (N_384,In_489,In_825);
nor U385 (N_385,In_1240,In_280);
nor U386 (N_386,In_102,In_27);
nor U387 (N_387,In_1443,In_685);
nor U388 (N_388,In_969,In_1153);
or U389 (N_389,In_317,In_1116);
nand U390 (N_390,In_401,In_780);
or U391 (N_391,In_563,In_1197);
and U392 (N_392,In_1236,In_507);
nand U393 (N_393,In_511,In_829);
and U394 (N_394,In_796,In_443);
nand U395 (N_395,In_869,In_992);
nand U396 (N_396,In_699,In_1388);
and U397 (N_397,In_466,In_1251);
or U398 (N_398,In_199,In_264);
nor U399 (N_399,In_83,In_1447);
nor U400 (N_400,In_284,In_1042);
nand U401 (N_401,In_845,In_54);
nor U402 (N_402,In_1011,In_231);
nand U403 (N_403,In_758,In_682);
and U404 (N_404,In_1351,In_293);
nor U405 (N_405,In_1025,In_833);
nor U406 (N_406,In_1039,In_17);
and U407 (N_407,In_931,In_944);
nor U408 (N_408,In_901,In_905);
nand U409 (N_409,In_64,In_1081);
nand U410 (N_410,In_621,In_609);
or U411 (N_411,In_562,In_6);
nand U412 (N_412,In_188,In_1241);
nor U413 (N_413,In_1230,In_11);
or U414 (N_414,In_15,In_1323);
nor U415 (N_415,In_290,In_214);
nand U416 (N_416,In_498,In_769);
or U417 (N_417,In_716,In_400);
and U418 (N_418,In_636,In_854);
nand U419 (N_419,In_1325,In_1139);
or U420 (N_420,In_843,In_673);
and U421 (N_421,In_420,In_388);
or U422 (N_422,In_330,In_522);
and U423 (N_423,In_1150,In_300);
and U424 (N_424,In_1222,In_1442);
nand U425 (N_425,In_1284,In_1272);
nand U426 (N_426,In_1279,In_85);
nand U427 (N_427,In_990,In_1214);
and U428 (N_428,In_575,In_1289);
nor U429 (N_429,In_737,In_852);
or U430 (N_430,In_107,In_1290);
or U431 (N_431,In_1363,In_1374);
and U432 (N_432,In_1282,In_338);
nand U433 (N_433,In_1026,In_306);
or U434 (N_434,In_1440,In_839);
and U435 (N_435,In_819,In_670);
and U436 (N_436,In_1231,In_1045);
and U437 (N_437,In_69,In_883);
and U438 (N_438,In_205,In_469);
or U439 (N_439,In_425,In_536);
nor U440 (N_440,In_791,In_1188);
nand U441 (N_441,In_16,In_111);
or U442 (N_442,In_178,In_933);
nor U443 (N_443,In_62,In_145);
and U444 (N_444,In_327,In_669);
or U445 (N_445,In_483,In_712);
or U446 (N_446,In_426,In_468);
and U447 (N_447,In_1162,In_233);
nor U448 (N_448,In_1410,In_1459);
nor U449 (N_449,In_1400,In_654);
nand U450 (N_450,In_1033,In_916);
and U451 (N_451,In_573,In_1355);
or U452 (N_452,In_1292,In_579);
and U453 (N_453,In_764,In_1438);
nand U454 (N_454,In_831,In_360);
nor U455 (N_455,In_272,In_1431);
and U456 (N_456,In_689,In_350);
or U457 (N_457,In_1249,In_936);
xnor U458 (N_458,In_464,In_875);
nor U459 (N_459,In_943,In_1452);
and U460 (N_460,In_859,In_1029);
and U461 (N_461,In_202,In_495);
nor U462 (N_462,In_984,In_571);
nand U463 (N_463,In_1224,In_365);
nand U464 (N_464,In_125,In_1392);
and U465 (N_465,In_1339,In_195);
nand U466 (N_466,In_892,In_1225);
nand U467 (N_467,In_44,In_857);
or U468 (N_468,In_688,In_802);
and U469 (N_469,In_528,In_232);
or U470 (N_470,In_234,In_907);
nor U471 (N_471,In_626,In_1009);
nor U472 (N_472,In_267,In_980);
nor U473 (N_473,In_555,In_76);
nor U474 (N_474,In_499,In_48);
nand U475 (N_475,In_949,In_700);
nand U476 (N_476,In_283,In_55);
nand U477 (N_477,In_597,In_1477);
nor U478 (N_478,In_1173,In_405);
or U479 (N_479,In_1405,In_509);
nor U480 (N_480,In_1229,In_470);
nand U481 (N_481,In_751,In_1073);
nand U482 (N_482,In_1212,In_1090);
nor U483 (N_483,In_81,In_369);
nand U484 (N_484,In_1281,In_154);
nor U485 (N_485,In_1006,In_779);
and U486 (N_486,In_966,In_226);
nand U487 (N_487,In_101,In_1346);
nor U488 (N_488,In_742,In_1144);
nor U489 (N_489,In_832,In_1082);
nor U490 (N_490,In_1348,In_180);
nor U491 (N_491,In_514,In_261);
and U492 (N_492,In_603,In_1067);
or U493 (N_493,In_628,In_1149);
nand U494 (N_494,In_754,In_696);
or U495 (N_495,In_1303,In_707);
nor U496 (N_496,In_1207,In_1332);
nand U497 (N_497,In_662,In_500);
nand U498 (N_498,In_529,In_1419);
and U499 (N_499,In_667,In_809);
nand U500 (N_500,In_115,In_409);
nor U501 (N_501,In_119,In_1087);
or U502 (N_502,In_800,In_1409);
nor U503 (N_503,In_1435,In_922);
nand U504 (N_504,In_762,In_595);
nand U505 (N_505,In_491,In_781);
or U506 (N_506,In_24,In_920);
and U507 (N_507,In_1487,In_1096);
nand U508 (N_508,In_1110,In_860);
and U509 (N_509,In_945,In_198);
or U510 (N_510,In_287,In_1203);
or U511 (N_511,In_627,In_52);
nor U512 (N_512,In_866,In_767);
nor U513 (N_513,In_1027,In_1252);
and U514 (N_514,In_1316,In_977);
nor U515 (N_515,In_804,In_1344);
or U516 (N_516,In_565,In_378);
nor U517 (N_517,In_1068,In_1421);
nand U518 (N_518,In_961,In_1171);
and U519 (N_519,In_391,In_93);
nand U520 (N_520,In_1054,In_1302);
nand U521 (N_521,In_940,In_1255);
nand U522 (N_522,In_1492,In_1115);
nor U523 (N_523,In_74,In_1161);
and U524 (N_524,In_650,In_1309);
nand U525 (N_525,In_297,In_1377);
nor U526 (N_526,In_756,In_90);
xnor U527 (N_527,In_446,In_1314);
nand U528 (N_528,In_835,In_88);
or U529 (N_529,In_36,In_1135);
and U530 (N_530,In_768,In_732);
nor U531 (N_531,In_861,In_1008);
nand U532 (N_532,In_1347,In_1004);
or U533 (N_533,In_331,In_1211);
nor U534 (N_534,In_25,In_200);
nor U535 (N_535,In_1475,In_1266);
xnor U536 (N_536,In_444,In_46);
and U537 (N_537,In_771,In_86);
or U538 (N_538,In_333,In_223);
nor U539 (N_539,In_516,In_138);
nand U540 (N_540,In_77,In_1248);
nand U541 (N_541,In_790,In_1451);
and U542 (N_542,In_1342,In_298);
nor U543 (N_543,In_542,In_741);
nor U544 (N_544,In_687,In_592);
nor U545 (N_545,In_808,In_219);
and U546 (N_546,In_749,In_691);
nand U547 (N_547,In_844,In_877);
nand U548 (N_548,In_652,In_1378);
nor U549 (N_549,In_429,In_656);
nand U550 (N_550,In_891,In_1334);
nor U551 (N_551,In_1491,In_467);
nand U552 (N_552,In_1280,In_38);
nand U553 (N_553,In_1015,In_591);
and U554 (N_554,In_884,In_983);
nand U555 (N_555,In_14,In_307);
nor U556 (N_556,In_1107,In_160);
nor U557 (N_557,In_1043,In_263);
and U558 (N_558,In_197,In_538);
and U559 (N_559,In_697,In_1044);
and U560 (N_560,In_921,In_148);
or U561 (N_561,In_788,In_303);
nor U562 (N_562,In_1059,In_320);
nor U563 (N_563,In_552,In_1050);
nand U564 (N_564,In_99,In_1340);
nand U565 (N_565,In_693,In_851);
nor U566 (N_566,In_8,In_1104);
and U567 (N_567,In_31,In_312);
or U568 (N_568,In_547,In_1456);
nor U569 (N_569,In_871,In_96);
and U570 (N_570,In_723,In_1368);
nand U571 (N_571,In_1411,In_730);
and U572 (N_572,In_158,In_1295);
nand U573 (N_573,In_1499,In_39);
and U574 (N_574,In_1359,In_617);
nand U575 (N_575,In_985,In_750);
and U576 (N_576,In_834,In_1495);
and U577 (N_577,In_929,In_345);
or U578 (N_578,In_481,In_131);
nor U579 (N_579,In_1242,In_179);
and U580 (N_580,In_1269,In_313);
nand U581 (N_581,In_406,In_644);
nand U582 (N_582,In_1101,In_1354);
and U583 (N_583,In_175,In_1141);
nor U584 (N_584,In_480,In_695);
and U585 (N_585,In_574,In_1080);
nor U586 (N_586,In_1471,In_1446);
nor U587 (N_587,In_545,In_557);
nor U588 (N_588,In_578,In_606);
nor U589 (N_589,In_228,In_853);
or U590 (N_590,In_1300,In_675);
or U591 (N_591,In_858,In_534);
and U592 (N_592,In_459,In_488);
nand U593 (N_593,In_713,In_841);
and U594 (N_594,In_864,In_918);
and U595 (N_595,In_12,In_971);
and U596 (N_596,In_32,In_181);
and U597 (N_597,In_908,In_75);
nand U598 (N_598,In_362,In_10);
or U599 (N_599,In_478,In_774);
nand U600 (N_600,In_588,In_910);
or U601 (N_601,In_747,In_1310);
nor U602 (N_602,In_976,In_1412);
nor U603 (N_603,In_377,In_1425);
nand U604 (N_604,In_655,In_150);
or U605 (N_605,In_4,In_975);
nand U606 (N_606,In_941,In_1223);
or U607 (N_607,In_322,In_1070);
or U608 (N_608,In_1313,In_332);
and U609 (N_609,In_1254,In_153);
nand U610 (N_610,In_568,In_1215);
nor U611 (N_611,In_722,In_141);
or U612 (N_612,In_397,In_1287);
nand U613 (N_613,In_1069,In_404);
or U614 (N_614,In_805,In_1423);
or U615 (N_615,In_665,In_1075);
or U616 (N_616,In_1193,In_238);
and U617 (N_617,In_1304,In_604);
nor U618 (N_618,In_1362,In_1003);
nor U619 (N_619,In_777,In_116);
and U620 (N_620,In_1470,In_886);
nand U621 (N_621,In_271,In_1129);
nand U622 (N_622,In_157,In_840);
nor U623 (N_623,In_23,In_1296);
nand U624 (N_624,In_630,In_357);
xnor U625 (N_625,In_613,In_475);
nor U626 (N_626,In_643,In_128);
and U627 (N_627,In_455,In_947);
or U628 (N_628,In_282,In_726);
or U629 (N_629,In_434,In_743);
nor U630 (N_630,In_934,In_1047);
and U631 (N_631,In_127,In_1032);
and U632 (N_632,In_544,In_384);
nand U633 (N_633,In_1157,In_1132);
and U634 (N_634,In_939,In_1391);
and U635 (N_635,In_1318,In_1195);
or U636 (N_636,In_70,In_356);
and U637 (N_637,In_965,In_208);
and U638 (N_638,In_240,In_632);
nor U639 (N_639,In_614,In_909);
or U640 (N_640,In_572,In_121);
nand U641 (N_641,In_9,In_814);
nor U642 (N_642,In_679,In_660);
nand U643 (N_643,In_305,In_848);
nor U644 (N_644,In_156,In_124);
nor U645 (N_645,In_849,In_589);
nor U646 (N_646,In_942,In_1111);
or U647 (N_647,In_34,In_1166);
or U648 (N_648,In_692,In_1420);
or U649 (N_649,In_925,In_1136);
nand U650 (N_650,In_738,In_622);
nand U651 (N_651,In_1307,In_341);
and U652 (N_652,In_1172,In_935);
and U653 (N_653,In_139,In_560);
nand U654 (N_654,In_1333,In_537);
and U655 (N_655,In_1243,In_248);
nand U656 (N_656,In_763,In_151);
and U657 (N_657,In_1031,In_324);
or U658 (N_658,In_368,In_162);
nor U659 (N_659,In_728,In_863);
and U660 (N_660,In_718,In_1273);
nor U661 (N_661,In_445,In_882);
and U662 (N_662,In_379,In_19);
nand U663 (N_663,In_1305,In_433);
nor U664 (N_664,In_239,In_28);
and U665 (N_665,In_1145,In_1100);
and U666 (N_666,In_951,In_456);
and U667 (N_667,In_1227,In_619);
and U668 (N_668,In_815,In_1485);
nor U669 (N_669,In_586,In_460);
nor U670 (N_670,In_291,In_1263);
nand U671 (N_671,In_63,In_1384);
or U672 (N_672,In_593,In_1120);
nand U673 (N_673,In_527,In_288);
and U674 (N_674,In_950,In_964);
nor U675 (N_675,In_417,In_1092);
and U676 (N_676,In_1022,In_1312);
or U677 (N_677,In_1218,In_1497);
nand U678 (N_678,In_794,In_392);
or U679 (N_679,In_235,In_123);
nor U680 (N_680,In_590,In_917);
or U681 (N_681,In_1152,In_1329);
and U682 (N_682,In_191,In_45);
or U683 (N_683,In_262,In_900);
and U684 (N_684,In_979,In_967);
or U685 (N_685,In_1265,In_576);
nand U686 (N_686,In_1328,In_122);
nand U687 (N_687,In_134,In_1238);
nor U688 (N_688,In_328,In_396);
nand U689 (N_689,In_602,In_1237);
and U690 (N_690,In_1424,In_1002);
and U691 (N_691,In_1198,In_919);
and U692 (N_692,In_1338,In_1158);
nand U693 (N_693,In_227,In_1467);
nor U694 (N_694,In_1085,In_736);
and U695 (N_695,In_865,In_447);
or U696 (N_696,In_109,In_194);
nor U697 (N_697,In_132,In_639);
and U698 (N_698,In_1322,In_375);
nor U699 (N_699,In_502,In_888);
and U700 (N_700,In_913,In_1436);
nor U701 (N_701,In_837,In_1213);
nor U702 (N_702,In_1246,In_372);
nor U703 (N_703,In_442,In_1482);
nor U704 (N_704,In_1128,In_733);
or U705 (N_705,In_1261,In_1021);
and U706 (N_706,In_169,In_991);
nor U707 (N_707,In_824,In_106);
nor U708 (N_708,In_411,In_1461);
or U709 (N_709,In_640,In_1160);
and U710 (N_710,In_1335,In_482);
and U711 (N_711,In_1178,In_221);
nor U712 (N_712,In_253,In_114);
or U713 (N_713,In_744,In_366);
nor U714 (N_714,In_1012,In_786);
nand U715 (N_715,In_152,In_218);
nand U716 (N_716,In_1337,In_878);
nor U717 (N_717,In_1023,In_1324);
nand U718 (N_718,In_1493,In_217);
nor U719 (N_719,In_902,In_266);
or U720 (N_720,In_424,In_171);
and U721 (N_721,In_1267,In_174);
and U722 (N_722,In_558,In_403);
nor U723 (N_723,In_1191,In_159);
and U724 (N_724,In_995,In_100);
nor U725 (N_725,In_1086,In_607);
or U726 (N_726,In_505,In_1078);
nor U727 (N_727,In_255,In_265);
or U728 (N_728,In_972,In_276);
or U729 (N_729,In_924,In_846);
nand U730 (N_730,In_515,In_1148);
nand U731 (N_731,In_531,In_1066);
or U732 (N_732,In_1187,In_1450);
nand U733 (N_733,In_1416,In_1234);
or U734 (N_734,In_582,In_1454);
nor U735 (N_735,In_412,In_987);
and U736 (N_736,In_1143,In_1179);
or U737 (N_737,In_382,In_787);
or U738 (N_738,In_149,In_797);
nand U739 (N_739,In_873,In_1428);
nand U740 (N_740,In_631,In_1034);
nor U741 (N_741,In_41,In_1275);
nor U742 (N_742,In_87,In_740);
and U743 (N_743,In_1177,In_1393);
nor U744 (N_744,In_371,In_503);
and U745 (N_745,In_251,In_501);
nand U746 (N_746,In_393,In_1030);
nand U747 (N_747,In_720,In_958);
nor U748 (N_748,In_1427,In_792);
and U749 (N_749,In_1278,In_1219);
and U750 (N_750,In_1252,In_959);
nor U751 (N_751,In_159,In_80);
nand U752 (N_752,In_545,In_1484);
nand U753 (N_753,In_1044,In_312);
and U754 (N_754,In_1118,In_687);
or U755 (N_755,In_255,In_295);
and U756 (N_756,In_505,In_1);
or U757 (N_757,In_424,In_1207);
nand U758 (N_758,In_48,In_1196);
and U759 (N_759,In_1002,In_1230);
nand U760 (N_760,In_93,In_892);
and U761 (N_761,In_884,In_137);
and U762 (N_762,In_1245,In_381);
and U763 (N_763,In_1104,In_1430);
nor U764 (N_764,In_138,In_47);
nand U765 (N_765,In_814,In_78);
nor U766 (N_766,In_804,In_261);
or U767 (N_767,In_453,In_1261);
or U768 (N_768,In_21,In_285);
nand U769 (N_769,In_669,In_37);
nand U770 (N_770,In_962,In_1148);
and U771 (N_771,In_750,In_146);
or U772 (N_772,In_1245,In_1098);
nand U773 (N_773,In_505,In_240);
nand U774 (N_774,In_816,In_1261);
nand U775 (N_775,In_1441,In_1087);
nand U776 (N_776,In_1330,In_747);
and U777 (N_777,In_450,In_1053);
and U778 (N_778,In_572,In_882);
nand U779 (N_779,In_1010,In_996);
nand U780 (N_780,In_969,In_833);
nor U781 (N_781,In_236,In_1253);
nor U782 (N_782,In_754,In_924);
and U783 (N_783,In_659,In_355);
and U784 (N_784,In_362,In_660);
nand U785 (N_785,In_1206,In_457);
nor U786 (N_786,In_583,In_1239);
and U787 (N_787,In_1485,In_1077);
nand U788 (N_788,In_77,In_929);
nor U789 (N_789,In_1123,In_947);
or U790 (N_790,In_325,In_911);
nand U791 (N_791,In_916,In_161);
or U792 (N_792,In_940,In_1014);
and U793 (N_793,In_717,In_174);
or U794 (N_794,In_369,In_594);
or U795 (N_795,In_623,In_965);
nor U796 (N_796,In_519,In_1173);
and U797 (N_797,In_811,In_923);
xor U798 (N_798,In_1372,In_956);
nor U799 (N_799,In_1380,In_818);
nor U800 (N_800,In_939,In_538);
nand U801 (N_801,In_208,In_1286);
nand U802 (N_802,In_988,In_787);
and U803 (N_803,In_245,In_575);
nand U804 (N_804,In_329,In_1191);
and U805 (N_805,In_1278,In_1418);
nand U806 (N_806,In_395,In_161);
and U807 (N_807,In_504,In_1477);
nor U808 (N_808,In_216,In_1120);
and U809 (N_809,In_1263,In_99);
or U810 (N_810,In_1260,In_1432);
nand U811 (N_811,In_1296,In_373);
nand U812 (N_812,In_1451,In_355);
or U813 (N_813,In_218,In_1076);
nor U814 (N_814,In_779,In_288);
and U815 (N_815,In_348,In_750);
nand U816 (N_816,In_430,In_981);
nand U817 (N_817,In_1037,In_782);
nand U818 (N_818,In_1467,In_1053);
and U819 (N_819,In_593,In_457);
nand U820 (N_820,In_807,In_839);
and U821 (N_821,In_631,In_26);
nor U822 (N_822,In_563,In_1283);
or U823 (N_823,In_1047,In_590);
nand U824 (N_824,In_319,In_682);
and U825 (N_825,In_8,In_1498);
nand U826 (N_826,In_894,In_887);
nand U827 (N_827,In_1045,In_64);
or U828 (N_828,In_480,In_1163);
nor U829 (N_829,In_1499,In_635);
xor U830 (N_830,In_1425,In_304);
and U831 (N_831,In_1267,In_403);
nand U832 (N_832,In_746,In_1477);
and U833 (N_833,In_1159,In_1482);
or U834 (N_834,In_1348,In_672);
or U835 (N_835,In_184,In_1106);
or U836 (N_836,In_388,In_308);
and U837 (N_837,In_67,In_320);
nor U838 (N_838,In_449,In_1132);
nor U839 (N_839,In_826,In_864);
nor U840 (N_840,In_1470,In_1093);
nand U841 (N_841,In_810,In_515);
nor U842 (N_842,In_382,In_1259);
nand U843 (N_843,In_1008,In_440);
and U844 (N_844,In_1480,In_1359);
nor U845 (N_845,In_278,In_726);
and U846 (N_846,In_951,In_602);
or U847 (N_847,In_105,In_906);
or U848 (N_848,In_1251,In_237);
and U849 (N_849,In_474,In_158);
nor U850 (N_850,In_1296,In_349);
nand U851 (N_851,In_1200,In_1193);
nor U852 (N_852,In_872,In_1422);
or U853 (N_853,In_779,In_1425);
nor U854 (N_854,In_200,In_386);
or U855 (N_855,In_1389,In_601);
nand U856 (N_856,In_1280,In_1205);
and U857 (N_857,In_290,In_339);
nor U858 (N_858,In_1217,In_685);
nor U859 (N_859,In_1424,In_1468);
nand U860 (N_860,In_1433,In_842);
or U861 (N_861,In_254,In_729);
or U862 (N_862,In_250,In_897);
or U863 (N_863,In_99,In_1152);
or U864 (N_864,In_1063,In_835);
and U865 (N_865,In_1009,In_67);
or U866 (N_866,In_1165,In_1274);
or U867 (N_867,In_107,In_978);
and U868 (N_868,In_859,In_1038);
nand U869 (N_869,In_170,In_1321);
and U870 (N_870,In_945,In_129);
or U871 (N_871,In_498,In_593);
and U872 (N_872,In_248,In_296);
and U873 (N_873,In_430,In_1318);
or U874 (N_874,In_610,In_1441);
nand U875 (N_875,In_835,In_653);
or U876 (N_876,In_795,In_346);
or U877 (N_877,In_554,In_1408);
or U878 (N_878,In_805,In_852);
and U879 (N_879,In_776,In_639);
or U880 (N_880,In_1464,In_1404);
xor U881 (N_881,In_441,In_81);
nor U882 (N_882,In_1138,In_1118);
nand U883 (N_883,In_1193,In_926);
or U884 (N_884,In_895,In_116);
or U885 (N_885,In_1152,In_224);
nand U886 (N_886,In_1237,In_1131);
and U887 (N_887,In_789,In_819);
and U888 (N_888,In_1370,In_1328);
or U889 (N_889,In_1036,In_1123);
nand U890 (N_890,In_340,In_937);
and U891 (N_891,In_247,In_1193);
or U892 (N_892,In_1481,In_722);
and U893 (N_893,In_491,In_170);
nor U894 (N_894,In_99,In_1270);
nor U895 (N_895,In_1374,In_708);
nor U896 (N_896,In_1105,In_1087);
nand U897 (N_897,In_450,In_953);
and U898 (N_898,In_1403,In_1260);
and U899 (N_899,In_572,In_1236);
and U900 (N_900,In_750,In_235);
nand U901 (N_901,In_710,In_1246);
or U902 (N_902,In_1031,In_95);
nor U903 (N_903,In_926,In_1011);
xor U904 (N_904,In_330,In_1296);
or U905 (N_905,In_641,In_1368);
nor U906 (N_906,In_892,In_624);
nand U907 (N_907,In_792,In_1251);
and U908 (N_908,In_1233,In_244);
nor U909 (N_909,In_1004,In_1403);
nand U910 (N_910,In_1045,In_417);
and U911 (N_911,In_1285,In_554);
and U912 (N_912,In_83,In_485);
nor U913 (N_913,In_1176,In_127);
or U914 (N_914,In_119,In_68);
and U915 (N_915,In_191,In_239);
or U916 (N_916,In_284,In_595);
and U917 (N_917,In_1289,In_758);
and U918 (N_918,In_748,In_749);
and U919 (N_919,In_415,In_359);
or U920 (N_920,In_126,In_838);
or U921 (N_921,In_1328,In_1192);
and U922 (N_922,In_1217,In_1213);
or U923 (N_923,In_817,In_1465);
nand U924 (N_924,In_1370,In_216);
or U925 (N_925,In_1191,In_769);
and U926 (N_926,In_1341,In_1356);
nor U927 (N_927,In_409,In_1256);
or U928 (N_928,In_1396,In_18);
or U929 (N_929,In_22,In_626);
xnor U930 (N_930,In_907,In_1187);
nor U931 (N_931,In_298,In_1284);
nor U932 (N_932,In_422,In_645);
nand U933 (N_933,In_1393,In_591);
nor U934 (N_934,In_496,In_970);
or U935 (N_935,In_232,In_1468);
and U936 (N_936,In_343,In_1278);
nand U937 (N_937,In_1412,In_1144);
and U938 (N_938,In_807,In_1397);
nor U939 (N_939,In_1107,In_387);
nand U940 (N_940,In_734,In_500);
or U941 (N_941,In_966,In_781);
xnor U942 (N_942,In_1257,In_1003);
and U943 (N_943,In_535,In_892);
and U944 (N_944,In_668,In_419);
or U945 (N_945,In_1374,In_614);
or U946 (N_946,In_1442,In_213);
or U947 (N_947,In_938,In_369);
nor U948 (N_948,In_954,In_515);
nand U949 (N_949,In_191,In_1472);
nand U950 (N_950,In_151,In_472);
nand U951 (N_951,In_263,In_115);
and U952 (N_952,In_233,In_1257);
nand U953 (N_953,In_503,In_781);
nand U954 (N_954,In_672,In_1441);
and U955 (N_955,In_1046,In_927);
nor U956 (N_956,In_1389,In_483);
or U957 (N_957,In_1433,In_367);
nor U958 (N_958,In_113,In_1010);
and U959 (N_959,In_143,In_563);
nand U960 (N_960,In_491,In_52);
nand U961 (N_961,In_1482,In_1334);
or U962 (N_962,In_486,In_518);
nor U963 (N_963,In_1385,In_1326);
and U964 (N_964,In_462,In_468);
or U965 (N_965,In_1298,In_1448);
nor U966 (N_966,In_102,In_528);
and U967 (N_967,In_199,In_590);
nand U968 (N_968,In_305,In_156);
xor U969 (N_969,In_942,In_748);
nor U970 (N_970,In_135,In_54);
or U971 (N_971,In_1106,In_122);
and U972 (N_972,In_1305,In_624);
nand U973 (N_973,In_932,In_580);
nand U974 (N_974,In_572,In_697);
or U975 (N_975,In_300,In_265);
nor U976 (N_976,In_127,In_1194);
and U977 (N_977,In_232,In_1220);
nand U978 (N_978,In_261,In_502);
or U979 (N_979,In_1264,In_677);
and U980 (N_980,In_674,In_393);
nand U981 (N_981,In_794,In_895);
nand U982 (N_982,In_1367,In_532);
nor U983 (N_983,In_1014,In_1008);
and U984 (N_984,In_664,In_607);
and U985 (N_985,In_1177,In_156);
and U986 (N_986,In_302,In_1417);
and U987 (N_987,In_83,In_565);
or U988 (N_988,In_424,In_168);
nand U989 (N_989,In_971,In_123);
and U990 (N_990,In_1446,In_746);
nor U991 (N_991,In_885,In_1030);
nor U992 (N_992,In_1364,In_1157);
or U993 (N_993,In_1404,In_415);
nand U994 (N_994,In_632,In_952);
and U995 (N_995,In_590,In_50);
nand U996 (N_996,In_165,In_1346);
and U997 (N_997,In_1499,In_851);
or U998 (N_998,In_1055,In_906);
and U999 (N_999,In_915,In_813);
and U1000 (N_1000,In_782,In_552);
and U1001 (N_1001,In_673,In_652);
and U1002 (N_1002,In_761,In_1021);
nand U1003 (N_1003,In_922,In_1472);
nor U1004 (N_1004,In_365,In_591);
nor U1005 (N_1005,In_382,In_1018);
and U1006 (N_1006,In_292,In_683);
and U1007 (N_1007,In_176,In_649);
nor U1008 (N_1008,In_1002,In_1430);
or U1009 (N_1009,In_1021,In_0);
and U1010 (N_1010,In_792,In_850);
and U1011 (N_1011,In_991,In_836);
or U1012 (N_1012,In_423,In_941);
or U1013 (N_1013,In_717,In_1239);
nand U1014 (N_1014,In_1433,In_1359);
nand U1015 (N_1015,In_102,In_747);
nand U1016 (N_1016,In_443,In_867);
nor U1017 (N_1017,In_1181,In_210);
or U1018 (N_1018,In_1223,In_1253);
nand U1019 (N_1019,In_1047,In_803);
or U1020 (N_1020,In_803,In_1386);
nor U1021 (N_1021,In_448,In_70);
nand U1022 (N_1022,In_314,In_361);
xnor U1023 (N_1023,In_1335,In_583);
or U1024 (N_1024,In_44,In_541);
nand U1025 (N_1025,In_164,In_912);
and U1026 (N_1026,In_1044,In_1077);
nor U1027 (N_1027,In_1289,In_1268);
and U1028 (N_1028,In_120,In_631);
nand U1029 (N_1029,In_894,In_1409);
or U1030 (N_1030,In_1209,In_1022);
nand U1031 (N_1031,In_1360,In_281);
and U1032 (N_1032,In_540,In_655);
nand U1033 (N_1033,In_573,In_520);
nand U1034 (N_1034,In_1103,In_1129);
nor U1035 (N_1035,In_999,In_1201);
or U1036 (N_1036,In_966,In_464);
or U1037 (N_1037,In_111,In_1189);
or U1038 (N_1038,In_304,In_151);
nand U1039 (N_1039,In_97,In_569);
and U1040 (N_1040,In_363,In_1263);
and U1041 (N_1041,In_1423,In_1279);
nand U1042 (N_1042,In_794,In_515);
nor U1043 (N_1043,In_1492,In_527);
nand U1044 (N_1044,In_868,In_575);
nand U1045 (N_1045,In_349,In_1046);
or U1046 (N_1046,In_768,In_256);
and U1047 (N_1047,In_447,In_248);
nor U1048 (N_1048,In_134,In_346);
or U1049 (N_1049,In_340,In_889);
and U1050 (N_1050,In_405,In_1057);
or U1051 (N_1051,In_1032,In_1371);
nor U1052 (N_1052,In_1372,In_1300);
nor U1053 (N_1053,In_1413,In_239);
nor U1054 (N_1054,In_1009,In_380);
nor U1055 (N_1055,In_693,In_1251);
nand U1056 (N_1056,In_1145,In_1154);
and U1057 (N_1057,In_1046,In_477);
nor U1058 (N_1058,In_909,In_538);
nor U1059 (N_1059,In_990,In_454);
and U1060 (N_1060,In_644,In_352);
and U1061 (N_1061,In_993,In_702);
or U1062 (N_1062,In_969,In_478);
xnor U1063 (N_1063,In_1347,In_738);
nor U1064 (N_1064,In_774,In_580);
nor U1065 (N_1065,In_1101,In_556);
or U1066 (N_1066,In_1429,In_387);
and U1067 (N_1067,In_255,In_172);
or U1068 (N_1068,In_17,In_1195);
nor U1069 (N_1069,In_96,In_339);
and U1070 (N_1070,In_1364,In_784);
and U1071 (N_1071,In_654,In_838);
and U1072 (N_1072,In_254,In_1045);
and U1073 (N_1073,In_911,In_906);
nand U1074 (N_1074,In_668,In_522);
and U1075 (N_1075,In_393,In_1269);
nor U1076 (N_1076,In_1464,In_607);
nor U1077 (N_1077,In_488,In_815);
and U1078 (N_1078,In_1345,In_885);
and U1079 (N_1079,In_826,In_60);
and U1080 (N_1080,In_594,In_993);
nand U1081 (N_1081,In_1349,In_1427);
and U1082 (N_1082,In_760,In_1342);
nor U1083 (N_1083,In_1260,In_27);
nand U1084 (N_1084,In_357,In_689);
nand U1085 (N_1085,In_665,In_1051);
and U1086 (N_1086,In_1218,In_558);
nor U1087 (N_1087,In_1066,In_425);
and U1088 (N_1088,In_330,In_179);
or U1089 (N_1089,In_41,In_1039);
nand U1090 (N_1090,In_1121,In_150);
or U1091 (N_1091,In_1143,In_687);
and U1092 (N_1092,In_1190,In_365);
nand U1093 (N_1093,In_222,In_152);
and U1094 (N_1094,In_197,In_1140);
and U1095 (N_1095,In_532,In_1402);
and U1096 (N_1096,In_254,In_946);
or U1097 (N_1097,In_1031,In_1183);
nand U1098 (N_1098,In_406,In_1224);
and U1099 (N_1099,In_730,In_657);
or U1100 (N_1100,In_1364,In_521);
or U1101 (N_1101,In_1347,In_532);
and U1102 (N_1102,In_1182,In_337);
and U1103 (N_1103,In_1201,In_1311);
and U1104 (N_1104,In_1100,In_805);
and U1105 (N_1105,In_229,In_1192);
nand U1106 (N_1106,In_517,In_437);
nor U1107 (N_1107,In_884,In_1173);
xnor U1108 (N_1108,In_520,In_1179);
nand U1109 (N_1109,In_343,In_696);
nor U1110 (N_1110,In_708,In_1056);
and U1111 (N_1111,In_1471,In_188);
and U1112 (N_1112,In_1083,In_1041);
nand U1113 (N_1113,In_565,In_1158);
nor U1114 (N_1114,In_1381,In_664);
nand U1115 (N_1115,In_553,In_294);
nor U1116 (N_1116,In_38,In_847);
nand U1117 (N_1117,In_544,In_925);
or U1118 (N_1118,In_762,In_1476);
nor U1119 (N_1119,In_1229,In_1329);
nor U1120 (N_1120,In_1025,In_1104);
and U1121 (N_1121,In_1149,In_1124);
and U1122 (N_1122,In_436,In_755);
nand U1123 (N_1123,In_572,In_1229);
nor U1124 (N_1124,In_1149,In_964);
nand U1125 (N_1125,In_404,In_915);
nor U1126 (N_1126,In_662,In_362);
nand U1127 (N_1127,In_781,In_347);
or U1128 (N_1128,In_1002,In_460);
nand U1129 (N_1129,In_876,In_686);
and U1130 (N_1130,In_1408,In_581);
nor U1131 (N_1131,In_247,In_1184);
nor U1132 (N_1132,In_184,In_1324);
or U1133 (N_1133,In_1177,In_874);
or U1134 (N_1134,In_1442,In_751);
nor U1135 (N_1135,In_824,In_1351);
xnor U1136 (N_1136,In_1402,In_1391);
nand U1137 (N_1137,In_1334,In_1263);
and U1138 (N_1138,In_839,In_498);
nor U1139 (N_1139,In_618,In_1139);
or U1140 (N_1140,In_1083,In_914);
and U1141 (N_1141,In_939,In_413);
nand U1142 (N_1142,In_49,In_1394);
and U1143 (N_1143,In_1182,In_1153);
xnor U1144 (N_1144,In_669,In_111);
nor U1145 (N_1145,In_210,In_1424);
and U1146 (N_1146,In_129,In_640);
nand U1147 (N_1147,In_1116,In_1178);
nor U1148 (N_1148,In_1393,In_440);
nand U1149 (N_1149,In_988,In_1363);
or U1150 (N_1150,In_197,In_797);
or U1151 (N_1151,In_1241,In_999);
or U1152 (N_1152,In_905,In_1313);
nor U1153 (N_1153,In_563,In_1039);
nor U1154 (N_1154,In_226,In_506);
and U1155 (N_1155,In_850,In_1169);
nand U1156 (N_1156,In_707,In_443);
xnor U1157 (N_1157,In_911,In_274);
nor U1158 (N_1158,In_117,In_738);
nand U1159 (N_1159,In_407,In_279);
nor U1160 (N_1160,In_446,In_216);
nand U1161 (N_1161,In_512,In_1433);
nor U1162 (N_1162,In_188,In_960);
nand U1163 (N_1163,In_1020,In_579);
nor U1164 (N_1164,In_224,In_621);
nand U1165 (N_1165,In_770,In_830);
and U1166 (N_1166,In_742,In_347);
nand U1167 (N_1167,In_326,In_768);
nor U1168 (N_1168,In_925,In_662);
nand U1169 (N_1169,In_957,In_847);
nand U1170 (N_1170,In_1470,In_245);
nand U1171 (N_1171,In_1407,In_690);
and U1172 (N_1172,In_1430,In_179);
nor U1173 (N_1173,In_862,In_1205);
or U1174 (N_1174,In_252,In_1462);
or U1175 (N_1175,In_1116,In_219);
and U1176 (N_1176,In_435,In_534);
nand U1177 (N_1177,In_1102,In_1176);
nand U1178 (N_1178,In_1029,In_157);
nand U1179 (N_1179,In_1493,In_1035);
nor U1180 (N_1180,In_330,In_1483);
nor U1181 (N_1181,In_880,In_610);
and U1182 (N_1182,In_391,In_596);
and U1183 (N_1183,In_874,In_1062);
or U1184 (N_1184,In_833,In_980);
or U1185 (N_1185,In_899,In_1353);
nor U1186 (N_1186,In_1041,In_38);
xnor U1187 (N_1187,In_503,In_352);
nor U1188 (N_1188,In_1012,In_529);
nor U1189 (N_1189,In_1320,In_1138);
nand U1190 (N_1190,In_550,In_1150);
and U1191 (N_1191,In_537,In_1406);
nand U1192 (N_1192,In_141,In_483);
or U1193 (N_1193,In_55,In_480);
or U1194 (N_1194,In_83,In_618);
or U1195 (N_1195,In_1031,In_956);
xnor U1196 (N_1196,In_1284,In_661);
nand U1197 (N_1197,In_347,In_1199);
nand U1198 (N_1198,In_572,In_649);
nand U1199 (N_1199,In_945,In_779);
or U1200 (N_1200,In_858,In_481);
or U1201 (N_1201,In_634,In_214);
nor U1202 (N_1202,In_82,In_549);
nand U1203 (N_1203,In_355,In_1493);
nor U1204 (N_1204,In_1456,In_1498);
nor U1205 (N_1205,In_311,In_1091);
nor U1206 (N_1206,In_742,In_682);
or U1207 (N_1207,In_235,In_377);
nand U1208 (N_1208,In_443,In_300);
and U1209 (N_1209,In_609,In_206);
or U1210 (N_1210,In_906,In_1011);
nand U1211 (N_1211,In_4,In_804);
nor U1212 (N_1212,In_88,In_773);
or U1213 (N_1213,In_1443,In_890);
nand U1214 (N_1214,In_1201,In_905);
nand U1215 (N_1215,In_866,In_346);
or U1216 (N_1216,In_1389,In_940);
nand U1217 (N_1217,In_640,In_1369);
nor U1218 (N_1218,In_1105,In_9);
or U1219 (N_1219,In_903,In_1103);
nor U1220 (N_1220,In_395,In_1346);
or U1221 (N_1221,In_248,In_786);
nor U1222 (N_1222,In_914,In_641);
nand U1223 (N_1223,In_71,In_68);
nor U1224 (N_1224,In_188,In_904);
and U1225 (N_1225,In_29,In_995);
and U1226 (N_1226,In_315,In_169);
and U1227 (N_1227,In_251,In_1205);
and U1228 (N_1228,In_697,In_1214);
nor U1229 (N_1229,In_533,In_485);
and U1230 (N_1230,In_1090,In_1027);
or U1231 (N_1231,In_1354,In_1128);
and U1232 (N_1232,In_346,In_1251);
nor U1233 (N_1233,In_1110,In_985);
nand U1234 (N_1234,In_516,In_698);
or U1235 (N_1235,In_80,In_1482);
nor U1236 (N_1236,In_786,In_776);
and U1237 (N_1237,In_377,In_165);
and U1238 (N_1238,In_1268,In_1320);
nand U1239 (N_1239,In_894,In_219);
nand U1240 (N_1240,In_768,In_910);
nand U1241 (N_1241,In_440,In_1476);
and U1242 (N_1242,In_980,In_696);
and U1243 (N_1243,In_572,In_1148);
nor U1244 (N_1244,In_97,In_1371);
nor U1245 (N_1245,In_841,In_1052);
or U1246 (N_1246,In_823,In_1120);
nor U1247 (N_1247,In_145,In_1398);
nor U1248 (N_1248,In_550,In_1056);
and U1249 (N_1249,In_180,In_1016);
nand U1250 (N_1250,In_6,In_237);
and U1251 (N_1251,In_1452,In_601);
nor U1252 (N_1252,In_738,In_869);
and U1253 (N_1253,In_1210,In_919);
nand U1254 (N_1254,In_135,In_389);
nor U1255 (N_1255,In_342,In_498);
or U1256 (N_1256,In_1166,In_345);
nor U1257 (N_1257,In_351,In_1237);
nor U1258 (N_1258,In_294,In_1137);
nand U1259 (N_1259,In_451,In_1087);
nand U1260 (N_1260,In_254,In_1186);
or U1261 (N_1261,In_734,In_1069);
nor U1262 (N_1262,In_843,In_854);
nand U1263 (N_1263,In_265,In_112);
and U1264 (N_1264,In_1234,In_69);
nand U1265 (N_1265,In_1106,In_202);
or U1266 (N_1266,In_606,In_408);
nand U1267 (N_1267,In_651,In_400);
or U1268 (N_1268,In_576,In_505);
nand U1269 (N_1269,In_1389,In_960);
and U1270 (N_1270,In_905,In_1226);
or U1271 (N_1271,In_70,In_1179);
nand U1272 (N_1272,In_1235,In_145);
or U1273 (N_1273,In_1356,In_206);
xnor U1274 (N_1274,In_839,In_355);
nor U1275 (N_1275,In_399,In_259);
nand U1276 (N_1276,In_970,In_376);
or U1277 (N_1277,In_903,In_1402);
and U1278 (N_1278,In_921,In_63);
nand U1279 (N_1279,In_978,In_601);
nor U1280 (N_1280,In_224,In_104);
and U1281 (N_1281,In_1379,In_275);
and U1282 (N_1282,In_1015,In_715);
nor U1283 (N_1283,In_1428,In_377);
and U1284 (N_1284,In_1470,In_591);
nand U1285 (N_1285,In_435,In_414);
or U1286 (N_1286,In_1291,In_324);
and U1287 (N_1287,In_1292,In_1300);
nor U1288 (N_1288,In_130,In_783);
nor U1289 (N_1289,In_462,In_928);
nand U1290 (N_1290,In_558,In_1163);
and U1291 (N_1291,In_926,In_1069);
nand U1292 (N_1292,In_1264,In_534);
or U1293 (N_1293,In_11,In_840);
nand U1294 (N_1294,In_1186,In_187);
nand U1295 (N_1295,In_320,In_908);
and U1296 (N_1296,In_1342,In_435);
nand U1297 (N_1297,In_1375,In_1003);
and U1298 (N_1298,In_946,In_259);
nor U1299 (N_1299,In_236,In_33);
nor U1300 (N_1300,In_1372,In_866);
nor U1301 (N_1301,In_762,In_1291);
or U1302 (N_1302,In_60,In_1261);
nor U1303 (N_1303,In_261,In_784);
or U1304 (N_1304,In_190,In_121);
and U1305 (N_1305,In_203,In_1053);
or U1306 (N_1306,In_9,In_1070);
and U1307 (N_1307,In_322,In_942);
and U1308 (N_1308,In_360,In_648);
or U1309 (N_1309,In_880,In_1004);
nor U1310 (N_1310,In_1176,In_81);
nand U1311 (N_1311,In_15,In_843);
or U1312 (N_1312,In_1270,In_205);
nor U1313 (N_1313,In_1376,In_594);
and U1314 (N_1314,In_1348,In_89);
or U1315 (N_1315,In_59,In_1463);
nand U1316 (N_1316,In_122,In_1369);
and U1317 (N_1317,In_1271,In_1207);
nor U1318 (N_1318,In_589,In_102);
or U1319 (N_1319,In_1112,In_119);
nand U1320 (N_1320,In_473,In_1393);
nand U1321 (N_1321,In_370,In_1497);
or U1322 (N_1322,In_1316,In_662);
or U1323 (N_1323,In_1123,In_452);
or U1324 (N_1324,In_1097,In_950);
and U1325 (N_1325,In_71,In_913);
nor U1326 (N_1326,In_1059,In_683);
nor U1327 (N_1327,In_353,In_645);
or U1328 (N_1328,In_821,In_2);
nand U1329 (N_1329,In_1346,In_1143);
nor U1330 (N_1330,In_668,In_1256);
nand U1331 (N_1331,In_879,In_134);
or U1332 (N_1332,In_1209,In_867);
or U1333 (N_1333,In_1206,In_1012);
and U1334 (N_1334,In_77,In_555);
or U1335 (N_1335,In_1037,In_1286);
nand U1336 (N_1336,In_498,In_1348);
or U1337 (N_1337,In_1165,In_572);
or U1338 (N_1338,In_421,In_520);
nor U1339 (N_1339,In_894,In_261);
or U1340 (N_1340,In_173,In_813);
and U1341 (N_1341,In_573,In_568);
and U1342 (N_1342,In_103,In_350);
xnor U1343 (N_1343,In_68,In_35);
nor U1344 (N_1344,In_804,In_90);
or U1345 (N_1345,In_667,In_16);
nand U1346 (N_1346,In_1424,In_946);
and U1347 (N_1347,In_1497,In_1267);
nor U1348 (N_1348,In_700,In_584);
and U1349 (N_1349,In_561,In_382);
nand U1350 (N_1350,In_167,In_1339);
nor U1351 (N_1351,In_1132,In_841);
nor U1352 (N_1352,In_535,In_1217);
and U1353 (N_1353,In_565,In_696);
nor U1354 (N_1354,In_112,In_327);
nand U1355 (N_1355,In_192,In_472);
and U1356 (N_1356,In_1138,In_47);
and U1357 (N_1357,In_199,In_389);
or U1358 (N_1358,In_274,In_1411);
or U1359 (N_1359,In_57,In_933);
nand U1360 (N_1360,In_231,In_960);
and U1361 (N_1361,In_823,In_254);
xor U1362 (N_1362,In_259,In_62);
or U1363 (N_1363,In_158,In_1047);
and U1364 (N_1364,In_353,In_339);
or U1365 (N_1365,In_1456,In_1452);
nand U1366 (N_1366,In_1482,In_249);
and U1367 (N_1367,In_314,In_1082);
nand U1368 (N_1368,In_156,In_966);
or U1369 (N_1369,In_95,In_682);
nor U1370 (N_1370,In_556,In_1047);
nor U1371 (N_1371,In_226,In_410);
nor U1372 (N_1372,In_381,In_179);
or U1373 (N_1373,In_152,In_200);
nand U1374 (N_1374,In_969,In_1147);
nand U1375 (N_1375,In_902,In_1015);
and U1376 (N_1376,In_626,In_4);
or U1377 (N_1377,In_595,In_1093);
or U1378 (N_1378,In_303,In_138);
nor U1379 (N_1379,In_520,In_780);
and U1380 (N_1380,In_267,In_1334);
nand U1381 (N_1381,In_9,In_1143);
or U1382 (N_1382,In_870,In_1247);
nand U1383 (N_1383,In_862,In_585);
xor U1384 (N_1384,In_392,In_925);
nand U1385 (N_1385,In_225,In_924);
nor U1386 (N_1386,In_766,In_982);
nand U1387 (N_1387,In_1382,In_642);
nand U1388 (N_1388,In_1313,In_542);
xnor U1389 (N_1389,In_1127,In_1179);
or U1390 (N_1390,In_1022,In_892);
and U1391 (N_1391,In_150,In_574);
nor U1392 (N_1392,In_1382,In_1131);
or U1393 (N_1393,In_150,In_384);
nor U1394 (N_1394,In_546,In_276);
nor U1395 (N_1395,In_589,In_756);
and U1396 (N_1396,In_1111,In_1363);
and U1397 (N_1397,In_1323,In_1429);
or U1398 (N_1398,In_145,In_727);
and U1399 (N_1399,In_661,In_763);
nand U1400 (N_1400,In_98,In_632);
and U1401 (N_1401,In_690,In_944);
and U1402 (N_1402,In_1355,In_1257);
and U1403 (N_1403,In_901,In_1431);
nand U1404 (N_1404,In_600,In_501);
or U1405 (N_1405,In_602,In_806);
nor U1406 (N_1406,In_697,In_110);
nor U1407 (N_1407,In_611,In_1206);
nand U1408 (N_1408,In_424,In_906);
nand U1409 (N_1409,In_205,In_1434);
and U1410 (N_1410,In_892,In_640);
or U1411 (N_1411,In_266,In_437);
nor U1412 (N_1412,In_649,In_881);
nor U1413 (N_1413,In_414,In_312);
nor U1414 (N_1414,In_814,In_1496);
or U1415 (N_1415,In_382,In_62);
or U1416 (N_1416,In_1196,In_770);
and U1417 (N_1417,In_88,In_263);
nor U1418 (N_1418,In_738,In_1290);
and U1419 (N_1419,In_281,In_1191);
nand U1420 (N_1420,In_1463,In_864);
nor U1421 (N_1421,In_176,In_374);
and U1422 (N_1422,In_1314,In_937);
nor U1423 (N_1423,In_1305,In_1354);
nor U1424 (N_1424,In_137,In_771);
nand U1425 (N_1425,In_1325,In_1204);
and U1426 (N_1426,In_80,In_1026);
or U1427 (N_1427,In_580,In_712);
or U1428 (N_1428,In_95,In_1020);
nor U1429 (N_1429,In_17,In_340);
and U1430 (N_1430,In_1318,In_162);
nor U1431 (N_1431,In_459,In_26);
or U1432 (N_1432,In_484,In_409);
and U1433 (N_1433,In_1108,In_911);
and U1434 (N_1434,In_95,In_126);
and U1435 (N_1435,In_722,In_1073);
and U1436 (N_1436,In_1046,In_707);
or U1437 (N_1437,In_232,In_688);
nor U1438 (N_1438,In_95,In_880);
and U1439 (N_1439,In_1409,In_833);
nor U1440 (N_1440,In_972,In_743);
or U1441 (N_1441,In_221,In_526);
nand U1442 (N_1442,In_1060,In_267);
or U1443 (N_1443,In_1194,In_125);
nand U1444 (N_1444,In_548,In_991);
nor U1445 (N_1445,In_1364,In_279);
nand U1446 (N_1446,In_1294,In_887);
and U1447 (N_1447,In_1350,In_1384);
nand U1448 (N_1448,In_1001,In_194);
or U1449 (N_1449,In_1223,In_1090);
nor U1450 (N_1450,In_1072,In_906);
and U1451 (N_1451,In_924,In_1115);
nand U1452 (N_1452,In_573,In_389);
nand U1453 (N_1453,In_494,In_880);
and U1454 (N_1454,In_1310,In_478);
and U1455 (N_1455,In_123,In_672);
and U1456 (N_1456,In_866,In_1095);
xnor U1457 (N_1457,In_148,In_1421);
and U1458 (N_1458,In_404,In_162);
nor U1459 (N_1459,In_366,In_497);
or U1460 (N_1460,In_132,In_596);
and U1461 (N_1461,In_208,In_31);
and U1462 (N_1462,In_588,In_141);
or U1463 (N_1463,In_231,In_515);
nand U1464 (N_1464,In_327,In_408);
nor U1465 (N_1465,In_547,In_1006);
nor U1466 (N_1466,In_969,In_720);
nand U1467 (N_1467,In_492,In_1268);
nor U1468 (N_1468,In_702,In_667);
nand U1469 (N_1469,In_1324,In_947);
nor U1470 (N_1470,In_956,In_46);
and U1471 (N_1471,In_974,In_327);
or U1472 (N_1472,In_240,In_1023);
nor U1473 (N_1473,In_913,In_1125);
nand U1474 (N_1474,In_1371,In_378);
nand U1475 (N_1475,In_1356,In_774);
or U1476 (N_1476,In_463,In_1001);
or U1477 (N_1477,In_1104,In_1082);
and U1478 (N_1478,In_1107,In_638);
nor U1479 (N_1479,In_1282,In_562);
xor U1480 (N_1480,In_1335,In_832);
nand U1481 (N_1481,In_8,In_1050);
xor U1482 (N_1482,In_4,In_1463);
or U1483 (N_1483,In_1069,In_49);
or U1484 (N_1484,In_1192,In_637);
or U1485 (N_1485,In_832,In_430);
and U1486 (N_1486,In_42,In_1141);
or U1487 (N_1487,In_563,In_350);
or U1488 (N_1488,In_738,In_181);
or U1489 (N_1489,In_670,In_1197);
nor U1490 (N_1490,In_1094,In_1121);
and U1491 (N_1491,In_715,In_1458);
and U1492 (N_1492,In_471,In_605);
nand U1493 (N_1493,In_780,In_933);
or U1494 (N_1494,In_178,In_637);
nand U1495 (N_1495,In_139,In_317);
or U1496 (N_1496,In_131,In_636);
xnor U1497 (N_1497,In_505,In_756);
and U1498 (N_1498,In_1009,In_1081);
nor U1499 (N_1499,In_92,In_1251);
and U1500 (N_1500,In_1298,In_923);
and U1501 (N_1501,In_461,In_1491);
nand U1502 (N_1502,In_937,In_109);
nor U1503 (N_1503,In_1415,In_760);
nand U1504 (N_1504,In_1062,In_597);
nand U1505 (N_1505,In_1284,In_216);
nand U1506 (N_1506,In_586,In_726);
nor U1507 (N_1507,In_940,In_36);
and U1508 (N_1508,In_1099,In_1233);
nand U1509 (N_1509,In_1263,In_1336);
and U1510 (N_1510,In_744,In_839);
and U1511 (N_1511,In_685,In_651);
or U1512 (N_1512,In_1262,In_25);
nor U1513 (N_1513,In_27,In_543);
or U1514 (N_1514,In_1410,In_1087);
or U1515 (N_1515,In_256,In_850);
or U1516 (N_1516,In_1379,In_405);
and U1517 (N_1517,In_608,In_510);
nor U1518 (N_1518,In_216,In_1227);
and U1519 (N_1519,In_68,In_692);
nor U1520 (N_1520,In_152,In_495);
or U1521 (N_1521,In_777,In_1180);
or U1522 (N_1522,In_392,In_872);
nor U1523 (N_1523,In_54,In_1348);
nand U1524 (N_1524,In_1426,In_1383);
nand U1525 (N_1525,In_491,In_439);
and U1526 (N_1526,In_173,In_1483);
nor U1527 (N_1527,In_110,In_536);
nor U1528 (N_1528,In_423,In_650);
or U1529 (N_1529,In_509,In_1219);
nand U1530 (N_1530,In_53,In_917);
and U1531 (N_1531,In_1050,In_1248);
nor U1532 (N_1532,In_1156,In_17);
nor U1533 (N_1533,In_668,In_935);
or U1534 (N_1534,In_118,In_1120);
nand U1535 (N_1535,In_726,In_698);
or U1536 (N_1536,In_333,In_686);
nand U1537 (N_1537,In_518,In_1033);
nand U1538 (N_1538,In_967,In_460);
and U1539 (N_1539,In_365,In_173);
or U1540 (N_1540,In_1251,In_862);
nand U1541 (N_1541,In_284,In_479);
nor U1542 (N_1542,In_713,In_1350);
nor U1543 (N_1543,In_263,In_68);
nor U1544 (N_1544,In_16,In_294);
or U1545 (N_1545,In_858,In_1229);
nor U1546 (N_1546,In_648,In_711);
nand U1547 (N_1547,In_1105,In_1422);
or U1548 (N_1548,In_701,In_538);
nand U1549 (N_1549,In_278,In_246);
nor U1550 (N_1550,In_822,In_482);
or U1551 (N_1551,In_1376,In_1300);
nor U1552 (N_1552,In_572,In_1337);
and U1553 (N_1553,In_989,In_943);
or U1554 (N_1554,In_870,In_1285);
or U1555 (N_1555,In_219,In_597);
and U1556 (N_1556,In_545,In_603);
nand U1557 (N_1557,In_1184,In_557);
and U1558 (N_1558,In_1089,In_471);
and U1559 (N_1559,In_1065,In_1343);
and U1560 (N_1560,In_420,In_822);
nor U1561 (N_1561,In_1132,In_961);
nor U1562 (N_1562,In_788,In_400);
or U1563 (N_1563,In_882,In_1174);
and U1564 (N_1564,In_1327,In_1494);
or U1565 (N_1565,In_414,In_388);
nor U1566 (N_1566,In_310,In_296);
and U1567 (N_1567,In_1046,In_84);
or U1568 (N_1568,In_1124,In_332);
nand U1569 (N_1569,In_1042,In_1321);
or U1570 (N_1570,In_49,In_235);
and U1571 (N_1571,In_949,In_40);
nor U1572 (N_1572,In_1177,In_922);
xor U1573 (N_1573,In_1353,In_833);
or U1574 (N_1574,In_522,In_752);
and U1575 (N_1575,In_771,In_398);
nor U1576 (N_1576,In_1446,In_713);
nand U1577 (N_1577,In_285,In_970);
nor U1578 (N_1578,In_619,In_1460);
and U1579 (N_1579,In_631,In_1170);
or U1580 (N_1580,In_973,In_401);
nand U1581 (N_1581,In_34,In_732);
and U1582 (N_1582,In_389,In_19);
nand U1583 (N_1583,In_608,In_1262);
or U1584 (N_1584,In_1386,In_1340);
or U1585 (N_1585,In_512,In_261);
or U1586 (N_1586,In_978,In_1259);
or U1587 (N_1587,In_56,In_94);
or U1588 (N_1588,In_1181,In_173);
and U1589 (N_1589,In_380,In_48);
or U1590 (N_1590,In_1125,In_11);
or U1591 (N_1591,In_1211,In_718);
xor U1592 (N_1592,In_808,In_1496);
nand U1593 (N_1593,In_1442,In_211);
and U1594 (N_1594,In_675,In_1265);
or U1595 (N_1595,In_1350,In_1377);
nand U1596 (N_1596,In_131,In_1295);
and U1597 (N_1597,In_1154,In_894);
nand U1598 (N_1598,In_909,In_1446);
nor U1599 (N_1599,In_455,In_552);
or U1600 (N_1600,In_808,In_1080);
nand U1601 (N_1601,In_1000,In_517);
nand U1602 (N_1602,In_247,In_782);
and U1603 (N_1603,In_646,In_1032);
and U1604 (N_1604,In_1342,In_1183);
or U1605 (N_1605,In_34,In_61);
and U1606 (N_1606,In_1278,In_134);
nand U1607 (N_1607,In_341,In_160);
nor U1608 (N_1608,In_1237,In_1197);
nand U1609 (N_1609,In_395,In_322);
nand U1610 (N_1610,In_1046,In_1302);
nand U1611 (N_1611,In_1366,In_602);
and U1612 (N_1612,In_388,In_148);
nor U1613 (N_1613,In_1393,In_920);
nand U1614 (N_1614,In_1483,In_371);
nand U1615 (N_1615,In_901,In_422);
nand U1616 (N_1616,In_930,In_913);
xnor U1617 (N_1617,In_1460,In_685);
or U1618 (N_1618,In_1312,In_785);
nor U1619 (N_1619,In_1355,In_194);
and U1620 (N_1620,In_1138,In_1189);
nand U1621 (N_1621,In_1188,In_181);
nor U1622 (N_1622,In_403,In_1415);
and U1623 (N_1623,In_650,In_1122);
and U1624 (N_1624,In_459,In_1312);
or U1625 (N_1625,In_860,In_29);
nand U1626 (N_1626,In_536,In_772);
and U1627 (N_1627,In_991,In_665);
nor U1628 (N_1628,In_340,In_1008);
nor U1629 (N_1629,In_181,In_501);
nand U1630 (N_1630,In_831,In_17);
or U1631 (N_1631,In_309,In_1402);
or U1632 (N_1632,In_889,In_308);
nand U1633 (N_1633,In_1143,In_1382);
or U1634 (N_1634,In_705,In_11);
nand U1635 (N_1635,In_167,In_511);
nand U1636 (N_1636,In_385,In_866);
and U1637 (N_1637,In_1175,In_1102);
nand U1638 (N_1638,In_138,In_248);
nand U1639 (N_1639,In_1101,In_953);
and U1640 (N_1640,In_1237,In_144);
and U1641 (N_1641,In_934,In_807);
and U1642 (N_1642,In_1254,In_439);
nor U1643 (N_1643,In_818,In_1082);
and U1644 (N_1644,In_864,In_911);
and U1645 (N_1645,In_273,In_85);
or U1646 (N_1646,In_1421,In_468);
nand U1647 (N_1647,In_42,In_509);
nor U1648 (N_1648,In_553,In_823);
and U1649 (N_1649,In_256,In_628);
or U1650 (N_1650,In_267,In_944);
and U1651 (N_1651,In_794,In_1042);
nor U1652 (N_1652,In_1324,In_149);
and U1653 (N_1653,In_621,In_1471);
or U1654 (N_1654,In_653,In_807);
and U1655 (N_1655,In_1124,In_422);
and U1656 (N_1656,In_191,In_1128);
or U1657 (N_1657,In_739,In_802);
and U1658 (N_1658,In_8,In_76);
and U1659 (N_1659,In_117,In_1363);
nand U1660 (N_1660,In_1477,In_474);
and U1661 (N_1661,In_367,In_1416);
nor U1662 (N_1662,In_696,In_1109);
nor U1663 (N_1663,In_658,In_466);
or U1664 (N_1664,In_253,In_543);
nand U1665 (N_1665,In_833,In_1461);
or U1666 (N_1666,In_1455,In_383);
or U1667 (N_1667,In_1479,In_745);
nand U1668 (N_1668,In_673,In_634);
or U1669 (N_1669,In_719,In_703);
nand U1670 (N_1670,In_1438,In_958);
nand U1671 (N_1671,In_149,In_87);
nand U1672 (N_1672,In_900,In_1457);
nor U1673 (N_1673,In_1197,In_1109);
and U1674 (N_1674,In_1125,In_107);
nor U1675 (N_1675,In_1020,In_1191);
or U1676 (N_1676,In_454,In_1176);
or U1677 (N_1677,In_660,In_691);
and U1678 (N_1678,In_1054,In_264);
and U1679 (N_1679,In_1400,In_743);
nor U1680 (N_1680,In_1386,In_1217);
or U1681 (N_1681,In_266,In_1206);
nand U1682 (N_1682,In_1266,In_401);
or U1683 (N_1683,In_954,In_480);
or U1684 (N_1684,In_1473,In_1189);
or U1685 (N_1685,In_664,In_1357);
or U1686 (N_1686,In_1034,In_149);
or U1687 (N_1687,In_1132,In_808);
nor U1688 (N_1688,In_598,In_1107);
nand U1689 (N_1689,In_46,In_505);
nor U1690 (N_1690,In_489,In_964);
and U1691 (N_1691,In_1378,In_453);
or U1692 (N_1692,In_150,In_55);
or U1693 (N_1693,In_304,In_1209);
nor U1694 (N_1694,In_660,In_120);
nor U1695 (N_1695,In_1047,In_95);
nor U1696 (N_1696,In_364,In_1306);
nor U1697 (N_1697,In_418,In_1329);
nand U1698 (N_1698,In_223,In_1125);
nand U1699 (N_1699,In_307,In_1152);
and U1700 (N_1700,In_1408,In_351);
nand U1701 (N_1701,In_697,In_1450);
or U1702 (N_1702,In_1044,In_1331);
nand U1703 (N_1703,In_1331,In_624);
nor U1704 (N_1704,In_614,In_290);
nand U1705 (N_1705,In_159,In_803);
nand U1706 (N_1706,In_947,In_700);
nand U1707 (N_1707,In_1075,In_179);
nand U1708 (N_1708,In_3,In_615);
nand U1709 (N_1709,In_793,In_1334);
nor U1710 (N_1710,In_262,In_610);
nor U1711 (N_1711,In_562,In_1060);
nor U1712 (N_1712,In_127,In_240);
nand U1713 (N_1713,In_995,In_102);
or U1714 (N_1714,In_731,In_1051);
and U1715 (N_1715,In_1159,In_1446);
and U1716 (N_1716,In_787,In_1377);
or U1717 (N_1717,In_823,In_945);
and U1718 (N_1718,In_552,In_12);
and U1719 (N_1719,In_290,In_417);
nor U1720 (N_1720,In_841,In_134);
and U1721 (N_1721,In_540,In_844);
or U1722 (N_1722,In_342,In_1156);
and U1723 (N_1723,In_1117,In_3);
nor U1724 (N_1724,In_310,In_501);
and U1725 (N_1725,In_1279,In_106);
nor U1726 (N_1726,In_53,In_648);
and U1727 (N_1727,In_233,In_808);
nand U1728 (N_1728,In_548,In_1376);
nor U1729 (N_1729,In_45,In_348);
or U1730 (N_1730,In_1479,In_1093);
nor U1731 (N_1731,In_1039,In_1379);
nand U1732 (N_1732,In_655,In_445);
and U1733 (N_1733,In_565,In_1212);
and U1734 (N_1734,In_642,In_29);
or U1735 (N_1735,In_910,In_306);
nor U1736 (N_1736,In_1159,In_1379);
nor U1737 (N_1737,In_810,In_920);
nand U1738 (N_1738,In_827,In_403);
and U1739 (N_1739,In_1293,In_95);
nand U1740 (N_1740,In_928,In_1063);
nor U1741 (N_1741,In_498,In_1260);
nor U1742 (N_1742,In_180,In_278);
nand U1743 (N_1743,In_537,In_267);
nor U1744 (N_1744,In_250,In_1001);
nand U1745 (N_1745,In_534,In_1465);
and U1746 (N_1746,In_530,In_642);
and U1747 (N_1747,In_1284,In_44);
and U1748 (N_1748,In_70,In_189);
nand U1749 (N_1749,In_23,In_39);
nand U1750 (N_1750,In_1321,In_891);
nor U1751 (N_1751,In_1182,In_1187);
nor U1752 (N_1752,In_191,In_1433);
and U1753 (N_1753,In_638,In_1345);
and U1754 (N_1754,In_1375,In_79);
or U1755 (N_1755,In_167,In_693);
and U1756 (N_1756,In_567,In_512);
and U1757 (N_1757,In_428,In_484);
and U1758 (N_1758,In_1476,In_465);
nand U1759 (N_1759,In_1436,In_1403);
or U1760 (N_1760,In_280,In_1335);
or U1761 (N_1761,In_1193,In_1389);
nand U1762 (N_1762,In_1217,In_117);
and U1763 (N_1763,In_319,In_1412);
nand U1764 (N_1764,In_442,In_1406);
or U1765 (N_1765,In_242,In_1367);
nand U1766 (N_1766,In_1355,In_979);
and U1767 (N_1767,In_333,In_373);
and U1768 (N_1768,In_623,In_1155);
nand U1769 (N_1769,In_431,In_384);
nor U1770 (N_1770,In_304,In_337);
or U1771 (N_1771,In_1269,In_66);
nand U1772 (N_1772,In_1236,In_630);
or U1773 (N_1773,In_1405,In_1078);
or U1774 (N_1774,In_481,In_26);
nor U1775 (N_1775,In_154,In_585);
and U1776 (N_1776,In_752,In_1460);
or U1777 (N_1777,In_308,In_3);
nor U1778 (N_1778,In_433,In_695);
or U1779 (N_1779,In_1395,In_362);
and U1780 (N_1780,In_1302,In_676);
or U1781 (N_1781,In_1244,In_73);
nand U1782 (N_1782,In_557,In_75);
nand U1783 (N_1783,In_247,In_1080);
and U1784 (N_1784,In_934,In_1054);
or U1785 (N_1785,In_803,In_207);
nor U1786 (N_1786,In_136,In_66);
and U1787 (N_1787,In_1269,In_606);
nand U1788 (N_1788,In_1256,In_841);
and U1789 (N_1789,In_503,In_379);
nand U1790 (N_1790,In_1396,In_1116);
or U1791 (N_1791,In_305,In_1340);
nand U1792 (N_1792,In_246,In_1138);
nand U1793 (N_1793,In_907,In_1195);
nor U1794 (N_1794,In_115,In_1279);
and U1795 (N_1795,In_919,In_1036);
nand U1796 (N_1796,In_1110,In_765);
and U1797 (N_1797,In_659,In_1046);
and U1798 (N_1798,In_934,In_1123);
or U1799 (N_1799,In_1433,In_1016);
and U1800 (N_1800,In_56,In_1);
or U1801 (N_1801,In_1162,In_1038);
nand U1802 (N_1802,In_1047,In_345);
or U1803 (N_1803,In_1342,In_535);
nor U1804 (N_1804,In_1285,In_734);
or U1805 (N_1805,In_821,In_1422);
and U1806 (N_1806,In_1387,In_1233);
nor U1807 (N_1807,In_504,In_1403);
and U1808 (N_1808,In_437,In_1037);
and U1809 (N_1809,In_265,In_869);
nor U1810 (N_1810,In_165,In_283);
or U1811 (N_1811,In_441,In_890);
nor U1812 (N_1812,In_793,In_396);
or U1813 (N_1813,In_363,In_1131);
and U1814 (N_1814,In_976,In_809);
nand U1815 (N_1815,In_760,In_488);
and U1816 (N_1816,In_1157,In_218);
nand U1817 (N_1817,In_229,In_496);
nor U1818 (N_1818,In_269,In_1130);
and U1819 (N_1819,In_524,In_1421);
and U1820 (N_1820,In_938,In_944);
nand U1821 (N_1821,In_722,In_983);
nor U1822 (N_1822,In_743,In_1413);
and U1823 (N_1823,In_528,In_274);
nand U1824 (N_1824,In_140,In_923);
or U1825 (N_1825,In_67,In_1061);
or U1826 (N_1826,In_1121,In_829);
nor U1827 (N_1827,In_32,In_1390);
or U1828 (N_1828,In_839,In_516);
or U1829 (N_1829,In_352,In_534);
nor U1830 (N_1830,In_61,In_1288);
nor U1831 (N_1831,In_1140,In_457);
or U1832 (N_1832,In_434,In_819);
or U1833 (N_1833,In_980,In_626);
and U1834 (N_1834,In_426,In_1488);
nor U1835 (N_1835,In_715,In_117);
and U1836 (N_1836,In_9,In_531);
nand U1837 (N_1837,In_647,In_681);
and U1838 (N_1838,In_1231,In_807);
nand U1839 (N_1839,In_500,In_1379);
nand U1840 (N_1840,In_349,In_1453);
or U1841 (N_1841,In_1104,In_862);
nand U1842 (N_1842,In_329,In_765);
nor U1843 (N_1843,In_338,In_725);
or U1844 (N_1844,In_1452,In_752);
and U1845 (N_1845,In_1116,In_82);
nor U1846 (N_1846,In_870,In_1000);
and U1847 (N_1847,In_865,In_1069);
nand U1848 (N_1848,In_51,In_1314);
and U1849 (N_1849,In_1220,In_1343);
nand U1850 (N_1850,In_460,In_1078);
xor U1851 (N_1851,In_1410,In_254);
nor U1852 (N_1852,In_535,In_929);
nor U1853 (N_1853,In_780,In_457);
or U1854 (N_1854,In_1002,In_940);
and U1855 (N_1855,In_749,In_466);
nor U1856 (N_1856,In_651,In_0);
nand U1857 (N_1857,In_857,In_1340);
or U1858 (N_1858,In_1466,In_1139);
nand U1859 (N_1859,In_666,In_1176);
and U1860 (N_1860,In_15,In_1148);
or U1861 (N_1861,In_77,In_1306);
and U1862 (N_1862,In_1308,In_1076);
or U1863 (N_1863,In_1361,In_1207);
or U1864 (N_1864,In_289,In_785);
nor U1865 (N_1865,In_28,In_852);
or U1866 (N_1866,In_388,In_997);
and U1867 (N_1867,In_345,In_1207);
nor U1868 (N_1868,In_96,In_857);
nand U1869 (N_1869,In_1043,In_1439);
and U1870 (N_1870,In_1224,In_1362);
or U1871 (N_1871,In_544,In_1002);
nand U1872 (N_1872,In_152,In_1005);
or U1873 (N_1873,In_512,In_975);
nor U1874 (N_1874,In_746,In_1015);
nor U1875 (N_1875,In_164,In_754);
or U1876 (N_1876,In_273,In_674);
nor U1877 (N_1877,In_1229,In_320);
nand U1878 (N_1878,In_144,In_580);
nor U1879 (N_1879,In_442,In_364);
or U1880 (N_1880,In_533,In_686);
or U1881 (N_1881,In_786,In_1226);
nand U1882 (N_1882,In_367,In_1066);
or U1883 (N_1883,In_459,In_54);
and U1884 (N_1884,In_1296,In_701);
nor U1885 (N_1885,In_447,In_314);
nand U1886 (N_1886,In_376,In_676);
nor U1887 (N_1887,In_537,In_672);
nor U1888 (N_1888,In_1149,In_621);
nor U1889 (N_1889,In_1180,In_1062);
nor U1890 (N_1890,In_43,In_446);
nand U1891 (N_1891,In_1306,In_1070);
nand U1892 (N_1892,In_791,In_428);
nand U1893 (N_1893,In_976,In_234);
or U1894 (N_1894,In_487,In_129);
nand U1895 (N_1895,In_570,In_540);
nor U1896 (N_1896,In_1103,In_693);
or U1897 (N_1897,In_189,In_1226);
nor U1898 (N_1898,In_1030,In_639);
nand U1899 (N_1899,In_1385,In_1243);
nor U1900 (N_1900,In_316,In_888);
nor U1901 (N_1901,In_117,In_267);
nand U1902 (N_1902,In_55,In_165);
and U1903 (N_1903,In_1356,In_146);
nand U1904 (N_1904,In_585,In_59);
and U1905 (N_1905,In_1079,In_1284);
nor U1906 (N_1906,In_390,In_1355);
or U1907 (N_1907,In_488,In_642);
nor U1908 (N_1908,In_666,In_1032);
and U1909 (N_1909,In_1385,In_1420);
or U1910 (N_1910,In_594,In_606);
nand U1911 (N_1911,In_561,In_1217);
nor U1912 (N_1912,In_1240,In_699);
nand U1913 (N_1913,In_992,In_219);
nor U1914 (N_1914,In_192,In_1037);
and U1915 (N_1915,In_1033,In_879);
or U1916 (N_1916,In_865,In_884);
or U1917 (N_1917,In_1309,In_439);
or U1918 (N_1918,In_538,In_549);
nor U1919 (N_1919,In_1381,In_167);
nand U1920 (N_1920,In_125,In_1264);
nand U1921 (N_1921,In_1432,In_1114);
and U1922 (N_1922,In_1379,In_810);
or U1923 (N_1923,In_407,In_194);
or U1924 (N_1924,In_352,In_568);
nand U1925 (N_1925,In_1196,In_657);
nand U1926 (N_1926,In_1343,In_251);
nor U1927 (N_1927,In_32,In_1405);
nand U1928 (N_1928,In_1392,In_1014);
nand U1929 (N_1929,In_1440,In_82);
nor U1930 (N_1930,In_65,In_205);
nor U1931 (N_1931,In_1324,In_555);
or U1932 (N_1932,In_815,In_1306);
nand U1933 (N_1933,In_63,In_674);
nand U1934 (N_1934,In_202,In_328);
or U1935 (N_1935,In_510,In_973);
nand U1936 (N_1936,In_570,In_1113);
nand U1937 (N_1937,In_1355,In_254);
nand U1938 (N_1938,In_331,In_254);
nand U1939 (N_1939,In_903,In_213);
nand U1940 (N_1940,In_1094,In_863);
nor U1941 (N_1941,In_1227,In_44);
nand U1942 (N_1942,In_865,In_1078);
or U1943 (N_1943,In_1261,In_748);
nand U1944 (N_1944,In_1156,In_1010);
or U1945 (N_1945,In_82,In_1100);
nand U1946 (N_1946,In_527,In_558);
nor U1947 (N_1947,In_75,In_1486);
nand U1948 (N_1948,In_951,In_579);
nor U1949 (N_1949,In_1449,In_946);
nand U1950 (N_1950,In_1299,In_193);
and U1951 (N_1951,In_214,In_1461);
and U1952 (N_1952,In_809,In_907);
nand U1953 (N_1953,In_144,In_275);
nor U1954 (N_1954,In_684,In_955);
or U1955 (N_1955,In_384,In_787);
nand U1956 (N_1956,In_313,In_817);
nor U1957 (N_1957,In_524,In_574);
or U1958 (N_1958,In_1133,In_1054);
nor U1959 (N_1959,In_1408,In_259);
and U1960 (N_1960,In_873,In_1021);
or U1961 (N_1961,In_1497,In_735);
and U1962 (N_1962,In_474,In_736);
and U1963 (N_1963,In_152,In_370);
and U1964 (N_1964,In_1184,In_29);
nand U1965 (N_1965,In_304,In_669);
nand U1966 (N_1966,In_1370,In_1080);
nand U1967 (N_1967,In_920,In_1102);
or U1968 (N_1968,In_58,In_45);
and U1969 (N_1969,In_494,In_917);
nand U1970 (N_1970,In_720,In_465);
nor U1971 (N_1971,In_1010,In_65);
or U1972 (N_1972,In_1151,In_589);
or U1973 (N_1973,In_1412,In_1291);
or U1974 (N_1974,In_50,In_727);
and U1975 (N_1975,In_784,In_1154);
nand U1976 (N_1976,In_177,In_9);
nand U1977 (N_1977,In_418,In_452);
nand U1978 (N_1978,In_380,In_745);
or U1979 (N_1979,In_1417,In_1310);
nand U1980 (N_1980,In_565,In_851);
and U1981 (N_1981,In_1012,In_1101);
nor U1982 (N_1982,In_1307,In_648);
nand U1983 (N_1983,In_219,In_1354);
and U1984 (N_1984,In_487,In_1284);
nor U1985 (N_1985,In_423,In_944);
and U1986 (N_1986,In_360,In_1000);
or U1987 (N_1987,In_994,In_1157);
and U1988 (N_1988,In_1244,In_802);
nor U1989 (N_1989,In_278,In_1334);
nand U1990 (N_1990,In_273,In_114);
nand U1991 (N_1991,In_114,In_830);
and U1992 (N_1992,In_1149,In_1431);
nor U1993 (N_1993,In_700,In_1122);
or U1994 (N_1994,In_467,In_864);
nor U1995 (N_1995,In_1021,In_1243);
nand U1996 (N_1996,In_226,In_1191);
and U1997 (N_1997,In_138,In_162);
nand U1998 (N_1998,In_733,In_1025);
nand U1999 (N_1999,In_1340,In_408);
nor U2000 (N_2000,In_653,In_1402);
and U2001 (N_2001,In_40,In_45);
or U2002 (N_2002,In_75,In_1096);
and U2003 (N_2003,In_615,In_1217);
or U2004 (N_2004,In_932,In_869);
and U2005 (N_2005,In_227,In_220);
and U2006 (N_2006,In_132,In_851);
or U2007 (N_2007,In_262,In_1325);
nand U2008 (N_2008,In_561,In_167);
or U2009 (N_2009,In_631,In_380);
nand U2010 (N_2010,In_1349,In_1068);
nand U2011 (N_2011,In_737,In_476);
nand U2012 (N_2012,In_1279,In_1446);
and U2013 (N_2013,In_445,In_1026);
nor U2014 (N_2014,In_95,In_19);
nor U2015 (N_2015,In_1221,In_356);
or U2016 (N_2016,In_117,In_787);
nand U2017 (N_2017,In_1056,In_383);
nand U2018 (N_2018,In_259,In_162);
and U2019 (N_2019,In_159,In_1138);
and U2020 (N_2020,In_762,In_11);
nand U2021 (N_2021,In_1407,In_1016);
nor U2022 (N_2022,In_1161,In_1430);
nand U2023 (N_2023,In_887,In_293);
nor U2024 (N_2024,In_975,In_1187);
nand U2025 (N_2025,In_1432,In_1268);
and U2026 (N_2026,In_1018,In_78);
nor U2027 (N_2027,In_696,In_678);
and U2028 (N_2028,In_149,In_1087);
or U2029 (N_2029,In_333,In_954);
and U2030 (N_2030,In_26,In_986);
or U2031 (N_2031,In_1367,In_959);
and U2032 (N_2032,In_1139,In_1165);
nand U2033 (N_2033,In_379,In_965);
and U2034 (N_2034,In_989,In_875);
and U2035 (N_2035,In_856,In_246);
nand U2036 (N_2036,In_274,In_1446);
or U2037 (N_2037,In_958,In_1397);
and U2038 (N_2038,In_1210,In_307);
or U2039 (N_2039,In_211,In_1012);
nor U2040 (N_2040,In_946,In_1432);
and U2041 (N_2041,In_114,In_235);
nand U2042 (N_2042,In_408,In_305);
nand U2043 (N_2043,In_1467,In_496);
or U2044 (N_2044,In_305,In_236);
or U2045 (N_2045,In_481,In_250);
and U2046 (N_2046,In_1108,In_1448);
nor U2047 (N_2047,In_790,In_626);
and U2048 (N_2048,In_122,In_242);
nand U2049 (N_2049,In_80,In_232);
and U2050 (N_2050,In_1291,In_1457);
nor U2051 (N_2051,In_973,In_364);
or U2052 (N_2052,In_1483,In_68);
or U2053 (N_2053,In_1003,In_246);
nand U2054 (N_2054,In_1491,In_241);
and U2055 (N_2055,In_753,In_721);
and U2056 (N_2056,In_215,In_1289);
and U2057 (N_2057,In_617,In_65);
or U2058 (N_2058,In_579,In_633);
and U2059 (N_2059,In_730,In_987);
nand U2060 (N_2060,In_1361,In_1166);
nor U2061 (N_2061,In_700,In_1261);
or U2062 (N_2062,In_474,In_525);
or U2063 (N_2063,In_939,In_1299);
and U2064 (N_2064,In_242,In_703);
nand U2065 (N_2065,In_515,In_1248);
nand U2066 (N_2066,In_483,In_509);
and U2067 (N_2067,In_427,In_1460);
and U2068 (N_2068,In_1346,In_1244);
nand U2069 (N_2069,In_1030,In_1145);
nand U2070 (N_2070,In_910,In_302);
nor U2071 (N_2071,In_1049,In_1179);
nor U2072 (N_2072,In_171,In_1267);
and U2073 (N_2073,In_31,In_1116);
and U2074 (N_2074,In_100,In_860);
nor U2075 (N_2075,In_412,In_97);
and U2076 (N_2076,In_430,In_1040);
nor U2077 (N_2077,In_838,In_1066);
nand U2078 (N_2078,In_1302,In_172);
or U2079 (N_2079,In_107,In_1384);
or U2080 (N_2080,In_918,In_1301);
nand U2081 (N_2081,In_282,In_629);
nor U2082 (N_2082,In_1160,In_834);
and U2083 (N_2083,In_248,In_1129);
nand U2084 (N_2084,In_45,In_625);
nor U2085 (N_2085,In_1386,In_888);
nor U2086 (N_2086,In_754,In_1004);
nand U2087 (N_2087,In_374,In_662);
and U2088 (N_2088,In_688,In_218);
nor U2089 (N_2089,In_801,In_856);
and U2090 (N_2090,In_683,In_445);
and U2091 (N_2091,In_271,In_736);
or U2092 (N_2092,In_305,In_88);
or U2093 (N_2093,In_162,In_453);
and U2094 (N_2094,In_922,In_498);
or U2095 (N_2095,In_429,In_1024);
or U2096 (N_2096,In_929,In_1384);
nand U2097 (N_2097,In_1129,In_438);
nor U2098 (N_2098,In_563,In_957);
nand U2099 (N_2099,In_806,In_997);
nor U2100 (N_2100,In_1038,In_819);
nand U2101 (N_2101,In_851,In_1175);
and U2102 (N_2102,In_535,In_446);
xor U2103 (N_2103,In_554,In_587);
and U2104 (N_2104,In_68,In_619);
nand U2105 (N_2105,In_624,In_1110);
nand U2106 (N_2106,In_767,In_1266);
nand U2107 (N_2107,In_211,In_1035);
nand U2108 (N_2108,In_957,In_1156);
or U2109 (N_2109,In_1464,In_549);
and U2110 (N_2110,In_572,In_1062);
and U2111 (N_2111,In_748,In_1159);
nand U2112 (N_2112,In_717,In_759);
and U2113 (N_2113,In_85,In_930);
or U2114 (N_2114,In_865,In_580);
nor U2115 (N_2115,In_742,In_1059);
nand U2116 (N_2116,In_385,In_847);
or U2117 (N_2117,In_689,In_1413);
xnor U2118 (N_2118,In_318,In_880);
and U2119 (N_2119,In_499,In_1166);
nor U2120 (N_2120,In_1374,In_1297);
nor U2121 (N_2121,In_255,In_922);
and U2122 (N_2122,In_496,In_646);
nor U2123 (N_2123,In_1333,In_827);
nand U2124 (N_2124,In_1434,In_1177);
xnor U2125 (N_2125,In_1343,In_1405);
and U2126 (N_2126,In_1420,In_588);
nor U2127 (N_2127,In_1143,In_1374);
nor U2128 (N_2128,In_882,In_205);
nand U2129 (N_2129,In_501,In_1340);
nand U2130 (N_2130,In_1217,In_651);
nand U2131 (N_2131,In_1356,In_519);
nand U2132 (N_2132,In_184,In_1238);
nor U2133 (N_2133,In_1096,In_224);
nand U2134 (N_2134,In_1120,In_1339);
or U2135 (N_2135,In_391,In_769);
or U2136 (N_2136,In_227,In_242);
or U2137 (N_2137,In_95,In_316);
nand U2138 (N_2138,In_1079,In_366);
or U2139 (N_2139,In_1364,In_68);
or U2140 (N_2140,In_630,In_1055);
nor U2141 (N_2141,In_343,In_1102);
and U2142 (N_2142,In_874,In_1253);
nand U2143 (N_2143,In_838,In_1140);
or U2144 (N_2144,In_1071,In_1101);
or U2145 (N_2145,In_1314,In_478);
nor U2146 (N_2146,In_690,In_176);
nor U2147 (N_2147,In_234,In_46);
nand U2148 (N_2148,In_916,In_931);
and U2149 (N_2149,In_1260,In_1106);
nand U2150 (N_2150,In_575,In_1418);
nand U2151 (N_2151,In_1300,In_63);
nand U2152 (N_2152,In_201,In_318);
and U2153 (N_2153,In_831,In_239);
or U2154 (N_2154,In_1444,In_368);
and U2155 (N_2155,In_664,In_486);
and U2156 (N_2156,In_901,In_1085);
nor U2157 (N_2157,In_619,In_111);
nor U2158 (N_2158,In_693,In_908);
nand U2159 (N_2159,In_151,In_339);
nor U2160 (N_2160,In_1277,In_969);
and U2161 (N_2161,In_291,In_1133);
nand U2162 (N_2162,In_1476,In_1491);
or U2163 (N_2163,In_151,In_950);
nor U2164 (N_2164,In_465,In_873);
or U2165 (N_2165,In_418,In_130);
nand U2166 (N_2166,In_835,In_192);
nand U2167 (N_2167,In_143,In_1242);
nor U2168 (N_2168,In_1315,In_492);
and U2169 (N_2169,In_454,In_1430);
nand U2170 (N_2170,In_1431,In_743);
or U2171 (N_2171,In_97,In_1437);
or U2172 (N_2172,In_959,In_705);
or U2173 (N_2173,In_105,In_273);
nand U2174 (N_2174,In_785,In_614);
nand U2175 (N_2175,In_1426,In_1174);
or U2176 (N_2176,In_1332,In_556);
or U2177 (N_2177,In_710,In_567);
or U2178 (N_2178,In_1,In_597);
and U2179 (N_2179,In_842,In_33);
and U2180 (N_2180,In_700,In_882);
nand U2181 (N_2181,In_425,In_888);
nand U2182 (N_2182,In_1378,In_716);
nor U2183 (N_2183,In_1067,In_396);
or U2184 (N_2184,In_521,In_1411);
nor U2185 (N_2185,In_28,In_175);
nand U2186 (N_2186,In_394,In_925);
nor U2187 (N_2187,In_585,In_495);
and U2188 (N_2188,In_269,In_1489);
nor U2189 (N_2189,In_8,In_1333);
or U2190 (N_2190,In_992,In_1496);
or U2191 (N_2191,In_1333,In_1046);
or U2192 (N_2192,In_832,In_58);
nor U2193 (N_2193,In_323,In_927);
nand U2194 (N_2194,In_1161,In_947);
or U2195 (N_2195,In_235,In_212);
nor U2196 (N_2196,In_1364,In_1400);
nand U2197 (N_2197,In_424,In_754);
or U2198 (N_2198,In_89,In_42);
or U2199 (N_2199,In_58,In_1003);
or U2200 (N_2200,In_540,In_1000);
nand U2201 (N_2201,In_271,In_651);
or U2202 (N_2202,In_415,In_1186);
nand U2203 (N_2203,In_683,In_594);
or U2204 (N_2204,In_1031,In_323);
nand U2205 (N_2205,In_890,In_33);
nand U2206 (N_2206,In_405,In_1462);
nor U2207 (N_2207,In_1346,In_902);
or U2208 (N_2208,In_191,In_701);
or U2209 (N_2209,In_1154,In_951);
and U2210 (N_2210,In_310,In_777);
nor U2211 (N_2211,In_134,In_1053);
nor U2212 (N_2212,In_1218,In_1085);
and U2213 (N_2213,In_937,In_106);
nand U2214 (N_2214,In_1035,In_354);
nand U2215 (N_2215,In_743,In_1232);
xnor U2216 (N_2216,In_884,In_615);
and U2217 (N_2217,In_1443,In_1132);
nand U2218 (N_2218,In_133,In_731);
or U2219 (N_2219,In_232,In_978);
nand U2220 (N_2220,In_375,In_417);
nor U2221 (N_2221,In_1193,In_191);
nor U2222 (N_2222,In_1098,In_1468);
or U2223 (N_2223,In_335,In_548);
and U2224 (N_2224,In_1147,In_725);
or U2225 (N_2225,In_1260,In_483);
and U2226 (N_2226,In_1343,In_52);
or U2227 (N_2227,In_311,In_137);
and U2228 (N_2228,In_609,In_1339);
or U2229 (N_2229,In_1225,In_409);
or U2230 (N_2230,In_59,In_667);
nand U2231 (N_2231,In_562,In_429);
or U2232 (N_2232,In_1249,In_275);
nor U2233 (N_2233,In_1486,In_679);
nand U2234 (N_2234,In_675,In_948);
nand U2235 (N_2235,In_405,In_1201);
or U2236 (N_2236,In_1479,In_1237);
and U2237 (N_2237,In_1386,In_1124);
nand U2238 (N_2238,In_1389,In_194);
xnor U2239 (N_2239,In_523,In_1382);
nor U2240 (N_2240,In_547,In_1020);
and U2241 (N_2241,In_726,In_949);
or U2242 (N_2242,In_634,In_287);
and U2243 (N_2243,In_1130,In_126);
nand U2244 (N_2244,In_1283,In_1379);
or U2245 (N_2245,In_1252,In_729);
or U2246 (N_2246,In_1184,In_69);
nor U2247 (N_2247,In_520,In_217);
nor U2248 (N_2248,In_260,In_666);
or U2249 (N_2249,In_1288,In_613);
and U2250 (N_2250,In_532,In_150);
nor U2251 (N_2251,In_226,In_561);
nor U2252 (N_2252,In_1320,In_740);
or U2253 (N_2253,In_169,In_361);
nand U2254 (N_2254,In_273,In_1098);
and U2255 (N_2255,In_1164,In_262);
nand U2256 (N_2256,In_969,In_899);
xnor U2257 (N_2257,In_1147,In_889);
and U2258 (N_2258,In_1389,In_1310);
nor U2259 (N_2259,In_1313,In_409);
and U2260 (N_2260,In_1169,In_1104);
nand U2261 (N_2261,In_1304,In_259);
nand U2262 (N_2262,In_1119,In_1245);
nand U2263 (N_2263,In_231,In_964);
nor U2264 (N_2264,In_828,In_386);
nand U2265 (N_2265,In_124,In_77);
and U2266 (N_2266,In_314,In_1326);
or U2267 (N_2267,In_13,In_255);
nor U2268 (N_2268,In_556,In_20);
or U2269 (N_2269,In_208,In_926);
or U2270 (N_2270,In_251,In_1022);
or U2271 (N_2271,In_285,In_487);
nand U2272 (N_2272,In_360,In_334);
nand U2273 (N_2273,In_471,In_1491);
nand U2274 (N_2274,In_835,In_1166);
nand U2275 (N_2275,In_810,In_837);
and U2276 (N_2276,In_220,In_600);
and U2277 (N_2277,In_1116,In_1237);
nand U2278 (N_2278,In_1329,In_827);
nand U2279 (N_2279,In_1375,In_1387);
nand U2280 (N_2280,In_155,In_578);
xor U2281 (N_2281,In_1173,In_645);
or U2282 (N_2282,In_1459,In_463);
or U2283 (N_2283,In_191,In_1146);
or U2284 (N_2284,In_324,In_826);
and U2285 (N_2285,In_296,In_220);
nand U2286 (N_2286,In_889,In_71);
nor U2287 (N_2287,In_474,In_524);
or U2288 (N_2288,In_702,In_1369);
nor U2289 (N_2289,In_1028,In_705);
nor U2290 (N_2290,In_241,In_831);
or U2291 (N_2291,In_1030,In_76);
nor U2292 (N_2292,In_537,In_181);
and U2293 (N_2293,In_542,In_543);
or U2294 (N_2294,In_675,In_789);
nor U2295 (N_2295,In_94,In_286);
and U2296 (N_2296,In_1382,In_25);
nand U2297 (N_2297,In_649,In_183);
or U2298 (N_2298,In_226,In_1494);
or U2299 (N_2299,In_1058,In_814);
and U2300 (N_2300,In_1099,In_670);
or U2301 (N_2301,In_1452,In_575);
nor U2302 (N_2302,In_222,In_639);
nand U2303 (N_2303,In_1196,In_960);
nor U2304 (N_2304,In_1182,In_881);
nor U2305 (N_2305,In_73,In_485);
or U2306 (N_2306,In_1298,In_1339);
or U2307 (N_2307,In_250,In_874);
or U2308 (N_2308,In_1389,In_179);
and U2309 (N_2309,In_880,In_1481);
nor U2310 (N_2310,In_455,In_958);
nor U2311 (N_2311,In_673,In_1428);
or U2312 (N_2312,In_1062,In_898);
nor U2313 (N_2313,In_1143,In_210);
nor U2314 (N_2314,In_499,In_977);
and U2315 (N_2315,In_733,In_145);
nand U2316 (N_2316,In_1259,In_798);
or U2317 (N_2317,In_1141,In_1053);
or U2318 (N_2318,In_772,In_47);
and U2319 (N_2319,In_1042,In_1284);
nor U2320 (N_2320,In_56,In_619);
nand U2321 (N_2321,In_1400,In_1121);
or U2322 (N_2322,In_125,In_804);
nand U2323 (N_2323,In_1132,In_399);
and U2324 (N_2324,In_1384,In_1270);
and U2325 (N_2325,In_1172,In_475);
nor U2326 (N_2326,In_926,In_946);
and U2327 (N_2327,In_1335,In_804);
or U2328 (N_2328,In_895,In_882);
nor U2329 (N_2329,In_188,In_448);
nand U2330 (N_2330,In_662,In_1089);
nor U2331 (N_2331,In_1482,In_296);
or U2332 (N_2332,In_811,In_1010);
nor U2333 (N_2333,In_593,In_458);
nor U2334 (N_2334,In_954,In_542);
nand U2335 (N_2335,In_352,In_291);
and U2336 (N_2336,In_161,In_680);
and U2337 (N_2337,In_1434,In_930);
and U2338 (N_2338,In_360,In_1142);
and U2339 (N_2339,In_1047,In_269);
nand U2340 (N_2340,In_1465,In_793);
nor U2341 (N_2341,In_1378,In_1362);
nor U2342 (N_2342,In_12,In_1074);
nor U2343 (N_2343,In_304,In_425);
nand U2344 (N_2344,In_1044,In_57);
nor U2345 (N_2345,In_1188,In_570);
or U2346 (N_2346,In_127,In_1180);
or U2347 (N_2347,In_1185,In_809);
nor U2348 (N_2348,In_1033,In_91);
and U2349 (N_2349,In_638,In_246);
nand U2350 (N_2350,In_598,In_116);
nand U2351 (N_2351,In_438,In_1274);
and U2352 (N_2352,In_730,In_622);
or U2353 (N_2353,In_505,In_65);
nor U2354 (N_2354,In_1016,In_721);
and U2355 (N_2355,In_1495,In_299);
nand U2356 (N_2356,In_284,In_1353);
or U2357 (N_2357,In_961,In_555);
or U2358 (N_2358,In_1329,In_1084);
or U2359 (N_2359,In_120,In_1088);
or U2360 (N_2360,In_965,In_977);
or U2361 (N_2361,In_822,In_1237);
or U2362 (N_2362,In_165,In_642);
nor U2363 (N_2363,In_773,In_256);
nand U2364 (N_2364,In_790,In_730);
nand U2365 (N_2365,In_658,In_281);
or U2366 (N_2366,In_277,In_161);
nor U2367 (N_2367,In_24,In_660);
or U2368 (N_2368,In_717,In_80);
nor U2369 (N_2369,In_1432,In_196);
or U2370 (N_2370,In_1388,In_675);
or U2371 (N_2371,In_1059,In_1363);
nand U2372 (N_2372,In_351,In_1288);
and U2373 (N_2373,In_960,In_786);
nand U2374 (N_2374,In_189,In_693);
and U2375 (N_2375,In_1241,In_110);
or U2376 (N_2376,In_1120,In_1008);
or U2377 (N_2377,In_94,In_1034);
or U2378 (N_2378,In_727,In_1361);
and U2379 (N_2379,In_294,In_742);
and U2380 (N_2380,In_724,In_360);
nand U2381 (N_2381,In_558,In_1190);
and U2382 (N_2382,In_300,In_500);
nand U2383 (N_2383,In_1144,In_1002);
nand U2384 (N_2384,In_307,In_313);
nand U2385 (N_2385,In_999,In_435);
and U2386 (N_2386,In_527,In_1287);
nor U2387 (N_2387,In_1409,In_616);
or U2388 (N_2388,In_1039,In_641);
or U2389 (N_2389,In_803,In_402);
and U2390 (N_2390,In_305,In_1495);
nor U2391 (N_2391,In_1031,In_153);
and U2392 (N_2392,In_1124,In_92);
nand U2393 (N_2393,In_941,In_746);
nor U2394 (N_2394,In_775,In_6);
and U2395 (N_2395,In_1091,In_618);
nor U2396 (N_2396,In_1102,In_987);
nand U2397 (N_2397,In_827,In_27);
and U2398 (N_2398,In_1201,In_1374);
nor U2399 (N_2399,In_1168,In_595);
nand U2400 (N_2400,In_680,In_1082);
nand U2401 (N_2401,In_771,In_436);
and U2402 (N_2402,In_362,In_391);
nor U2403 (N_2403,In_1319,In_1244);
nand U2404 (N_2404,In_692,In_316);
nor U2405 (N_2405,In_1079,In_697);
and U2406 (N_2406,In_892,In_654);
or U2407 (N_2407,In_1199,In_324);
and U2408 (N_2408,In_1370,In_194);
or U2409 (N_2409,In_641,In_1407);
or U2410 (N_2410,In_1040,In_1146);
and U2411 (N_2411,In_1383,In_11);
nand U2412 (N_2412,In_115,In_257);
or U2413 (N_2413,In_567,In_401);
nand U2414 (N_2414,In_1403,In_672);
and U2415 (N_2415,In_1176,In_1016);
nand U2416 (N_2416,In_762,In_499);
or U2417 (N_2417,In_669,In_1088);
nor U2418 (N_2418,In_664,In_584);
nor U2419 (N_2419,In_264,In_542);
nor U2420 (N_2420,In_1105,In_501);
nand U2421 (N_2421,In_132,In_1241);
or U2422 (N_2422,In_349,In_1086);
and U2423 (N_2423,In_1493,In_367);
nor U2424 (N_2424,In_20,In_678);
or U2425 (N_2425,In_783,In_121);
or U2426 (N_2426,In_1097,In_802);
or U2427 (N_2427,In_187,In_121);
or U2428 (N_2428,In_1401,In_1497);
and U2429 (N_2429,In_922,In_1481);
xnor U2430 (N_2430,In_264,In_997);
or U2431 (N_2431,In_827,In_84);
or U2432 (N_2432,In_1396,In_1391);
nand U2433 (N_2433,In_709,In_39);
nor U2434 (N_2434,In_880,In_1251);
nand U2435 (N_2435,In_1085,In_210);
and U2436 (N_2436,In_13,In_890);
and U2437 (N_2437,In_1204,In_1072);
and U2438 (N_2438,In_781,In_1478);
nand U2439 (N_2439,In_2,In_871);
and U2440 (N_2440,In_155,In_200);
and U2441 (N_2441,In_437,In_1315);
and U2442 (N_2442,In_428,In_859);
nand U2443 (N_2443,In_310,In_753);
or U2444 (N_2444,In_1023,In_823);
nand U2445 (N_2445,In_1147,In_177);
or U2446 (N_2446,In_257,In_1213);
nor U2447 (N_2447,In_1316,In_1182);
and U2448 (N_2448,In_998,In_33);
nand U2449 (N_2449,In_126,In_682);
and U2450 (N_2450,In_1014,In_1407);
nor U2451 (N_2451,In_334,In_116);
nand U2452 (N_2452,In_519,In_616);
nor U2453 (N_2453,In_872,In_1038);
nor U2454 (N_2454,In_1356,In_782);
nand U2455 (N_2455,In_1440,In_1210);
or U2456 (N_2456,In_1205,In_1413);
and U2457 (N_2457,In_1390,In_528);
or U2458 (N_2458,In_1408,In_1436);
xor U2459 (N_2459,In_944,In_91);
and U2460 (N_2460,In_1257,In_64);
nand U2461 (N_2461,In_174,In_1407);
nor U2462 (N_2462,In_708,In_184);
nand U2463 (N_2463,In_813,In_121);
nor U2464 (N_2464,In_213,In_874);
nand U2465 (N_2465,In_32,In_692);
and U2466 (N_2466,In_1382,In_362);
nor U2467 (N_2467,In_620,In_614);
and U2468 (N_2468,In_947,In_1247);
nor U2469 (N_2469,In_269,In_690);
or U2470 (N_2470,In_885,In_598);
or U2471 (N_2471,In_719,In_1352);
nor U2472 (N_2472,In_267,In_855);
nand U2473 (N_2473,In_699,In_882);
nand U2474 (N_2474,In_813,In_1174);
and U2475 (N_2475,In_608,In_696);
nand U2476 (N_2476,In_716,In_1479);
or U2477 (N_2477,In_990,In_1302);
nand U2478 (N_2478,In_596,In_664);
nor U2479 (N_2479,In_56,In_770);
nor U2480 (N_2480,In_345,In_1297);
or U2481 (N_2481,In_681,In_637);
nand U2482 (N_2482,In_257,In_967);
nor U2483 (N_2483,In_1201,In_1428);
and U2484 (N_2484,In_1080,In_101);
nor U2485 (N_2485,In_949,In_970);
and U2486 (N_2486,In_1233,In_853);
nand U2487 (N_2487,In_1173,In_1407);
nand U2488 (N_2488,In_1192,In_376);
or U2489 (N_2489,In_349,In_941);
and U2490 (N_2490,In_1242,In_1439);
or U2491 (N_2491,In_440,In_698);
or U2492 (N_2492,In_166,In_665);
or U2493 (N_2493,In_47,In_99);
nand U2494 (N_2494,In_1277,In_1225);
and U2495 (N_2495,In_1462,In_466);
nand U2496 (N_2496,In_813,In_101);
and U2497 (N_2497,In_941,In_1381);
nand U2498 (N_2498,In_903,In_679);
nand U2499 (N_2499,In_351,In_1373);
nor U2500 (N_2500,In_844,In_1444);
nor U2501 (N_2501,In_579,In_626);
nor U2502 (N_2502,In_1239,In_597);
or U2503 (N_2503,In_976,In_1007);
nand U2504 (N_2504,In_1235,In_788);
and U2505 (N_2505,In_1131,In_936);
and U2506 (N_2506,In_1211,In_1361);
nand U2507 (N_2507,In_386,In_59);
or U2508 (N_2508,In_1479,In_764);
and U2509 (N_2509,In_863,In_913);
nand U2510 (N_2510,In_1273,In_593);
nand U2511 (N_2511,In_1420,In_43);
nor U2512 (N_2512,In_704,In_453);
nand U2513 (N_2513,In_1329,In_1346);
or U2514 (N_2514,In_515,In_146);
nor U2515 (N_2515,In_1365,In_776);
nor U2516 (N_2516,In_830,In_583);
nor U2517 (N_2517,In_1388,In_371);
nor U2518 (N_2518,In_1143,In_982);
nor U2519 (N_2519,In_455,In_866);
and U2520 (N_2520,In_96,In_1478);
and U2521 (N_2521,In_1115,In_841);
nand U2522 (N_2522,In_654,In_240);
and U2523 (N_2523,In_246,In_180);
nand U2524 (N_2524,In_207,In_1025);
and U2525 (N_2525,In_416,In_12);
xor U2526 (N_2526,In_1080,In_403);
nor U2527 (N_2527,In_15,In_740);
nand U2528 (N_2528,In_622,In_1424);
nor U2529 (N_2529,In_1150,In_1347);
or U2530 (N_2530,In_337,In_961);
or U2531 (N_2531,In_898,In_1073);
or U2532 (N_2532,In_1264,In_18);
and U2533 (N_2533,In_1185,In_39);
xnor U2534 (N_2534,In_1224,In_879);
or U2535 (N_2535,In_1358,In_215);
or U2536 (N_2536,In_146,In_783);
nand U2537 (N_2537,In_1151,In_603);
or U2538 (N_2538,In_1059,In_326);
or U2539 (N_2539,In_909,In_988);
xor U2540 (N_2540,In_1129,In_37);
and U2541 (N_2541,In_421,In_969);
nand U2542 (N_2542,In_1407,In_1059);
nand U2543 (N_2543,In_1409,In_57);
or U2544 (N_2544,In_1008,In_912);
nand U2545 (N_2545,In_671,In_144);
nand U2546 (N_2546,In_357,In_780);
and U2547 (N_2547,In_1173,In_990);
nor U2548 (N_2548,In_1012,In_6);
or U2549 (N_2549,In_606,In_1390);
nand U2550 (N_2550,In_922,In_586);
or U2551 (N_2551,In_1028,In_610);
nand U2552 (N_2552,In_957,In_502);
nand U2553 (N_2553,In_253,In_669);
nand U2554 (N_2554,In_716,In_879);
or U2555 (N_2555,In_398,In_782);
nand U2556 (N_2556,In_1106,In_700);
and U2557 (N_2557,In_1075,In_102);
or U2558 (N_2558,In_29,In_1017);
or U2559 (N_2559,In_482,In_1267);
nor U2560 (N_2560,In_789,In_856);
nand U2561 (N_2561,In_1410,In_17);
nand U2562 (N_2562,In_130,In_440);
nand U2563 (N_2563,In_128,In_802);
and U2564 (N_2564,In_429,In_1008);
and U2565 (N_2565,In_311,In_582);
nand U2566 (N_2566,In_835,In_957);
or U2567 (N_2567,In_782,In_370);
or U2568 (N_2568,In_102,In_416);
nor U2569 (N_2569,In_484,In_694);
nor U2570 (N_2570,In_787,In_778);
nor U2571 (N_2571,In_903,In_365);
nor U2572 (N_2572,In_1311,In_775);
nor U2573 (N_2573,In_64,In_627);
nand U2574 (N_2574,In_1486,In_692);
nand U2575 (N_2575,In_1441,In_582);
and U2576 (N_2576,In_564,In_1316);
nand U2577 (N_2577,In_563,In_623);
nor U2578 (N_2578,In_1434,In_589);
nor U2579 (N_2579,In_353,In_1468);
or U2580 (N_2580,In_1142,In_48);
nor U2581 (N_2581,In_1033,In_635);
nand U2582 (N_2582,In_1215,In_1111);
and U2583 (N_2583,In_233,In_12);
or U2584 (N_2584,In_23,In_790);
nand U2585 (N_2585,In_191,In_132);
nand U2586 (N_2586,In_1222,In_663);
and U2587 (N_2587,In_834,In_1215);
nand U2588 (N_2588,In_991,In_91);
nand U2589 (N_2589,In_969,In_1139);
nor U2590 (N_2590,In_1481,In_297);
nand U2591 (N_2591,In_1443,In_551);
or U2592 (N_2592,In_173,In_1393);
nand U2593 (N_2593,In_369,In_1377);
nor U2594 (N_2594,In_986,In_608);
nor U2595 (N_2595,In_1170,In_482);
nor U2596 (N_2596,In_342,In_486);
nor U2597 (N_2597,In_833,In_1236);
and U2598 (N_2598,In_325,In_453);
or U2599 (N_2599,In_1124,In_984);
and U2600 (N_2600,In_1398,In_1397);
and U2601 (N_2601,In_253,In_521);
nor U2602 (N_2602,In_747,In_998);
nor U2603 (N_2603,In_643,In_180);
and U2604 (N_2604,In_691,In_177);
nor U2605 (N_2605,In_894,In_270);
xnor U2606 (N_2606,In_1328,In_265);
or U2607 (N_2607,In_1081,In_908);
nor U2608 (N_2608,In_1150,In_227);
or U2609 (N_2609,In_104,In_1355);
nand U2610 (N_2610,In_312,In_884);
or U2611 (N_2611,In_512,In_842);
nand U2612 (N_2612,In_324,In_632);
or U2613 (N_2613,In_295,In_792);
or U2614 (N_2614,In_299,In_1052);
and U2615 (N_2615,In_1366,In_466);
and U2616 (N_2616,In_20,In_1178);
or U2617 (N_2617,In_1126,In_1244);
or U2618 (N_2618,In_1215,In_1033);
nor U2619 (N_2619,In_164,In_1014);
and U2620 (N_2620,In_83,In_1409);
nor U2621 (N_2621,In_393,In_264);
nor U2622 (N_2622,In_1284,In_443);
or U2623 (N_2623,In_1215,In_1079);
or U2624 (N_2624,In_619,In_991);
nor U2625 (N_2625,In_97,In_964);
and U2626 (N_2626,In_688,In_293);
nand U2627 (N_2627,In_198,In_546);
and U2628 (N_2628,In_1251,In_137);
nor U2629 (N_2629,In_905,In_255);
nand U2630 (N_2630,In_590,In_4);
nand U2631 (N_2631,In_657,In_252);
or U2632 (N_2632,In_1289,In_1494);
and U2633 (N_2633,In_421,In_1327);
nand U2634 (N_2634,In_60,In_798);
and U2635 (N_2635,In_340,In_249);
or U2636 (N_2636,In_1121,In_468);
or U2637 (N_2637,In_1104,In_951);
nand U2638 (N_2638,In_1087,In_604);
nand U2639 (N_2639,In_726,In_206);
and U2640 (N_2640,In_779,In_765);
nand U2641 (N_2641,In_875,In_543);
or U2642 (N_2642,In_828,In_343);
nand U2643 (N_2643,In_39,In_128);
and U2644 (N_2644,In_402,In_324);
or U2645 (N_2645,In_61,In_1258);
and U2646 (N_2646,In_648,In_696);
or U2647 (N_2647,In_147,In_148);
nor U2648 (N_2648,In_757,In_1259);
and U2649 (N_2649,In_1019,In_1354);
nand U2650 (N_2650,In_923,In_900);
and U2651 (N_2651,In_1378,In_95);
or U2652 (N_2652,In_1114,In_153);
nor U2653 (N_2653,In_661,In_357);
nor U2654 (N_2654,In_664,In_416);
nand U2655 (N_2655,In_411,In_1404);
and U2656 (N_2656,In_533,In_247);
nor U2657 (N_2657,In_358,In_668);
nand U2658 (N_2658,In_1483,In_1072);
nor U2659 (N_2659,In_1497,In_485);
and U2660 (N_2660,In_670,In_874);
nor U2661 (N_2661,In_1156,In_700);
and U2662 (N_2662,In_461,In_10);
nand U2663 (N_2663,In_976,In_953);
or U2664 (N_2664,In_420,In_412);
and U2665 (N_2665,In_1101,In_527);
nor U2666 (N_2666,In_283,In_323);
and U2667 (N_2667,In_571,In_743);
and U2668 (N_2668,In_1181,In_1282);
and U2669 (N_2669,In_1200,In_645);
nor U2670 (N_2670,In_1016,In_1);
or U2671 (N_2671,In_352,In_100);
nor U2672 (N_2672,In_1480,In_854);
or U2673 (N_2673,In_720,In_1322);
and U2674 (N_2674,In_329,In_451);
nand U2675 (N_2675,In_748,In_1375);
nor U2676 (N_2676,In_1193,In_475);
nand U2677 (N_2677,In_243,In_812);
nand U2678 (N_2678,In_99,In_1134);
nor U2679 (N_2679,In_753,In_1342);
and U2680 (N_2680,In_307,In_983);
nand U2681 (N_2681,In_977,In_1287);
nand U2682 (N_2682,In_457,In_381);
or U2683 (N_2683,In_987,In_280);
nand U2684 (N_2684,In_466,In_553);
and U2685 (N_2685,In_875,In_70);
nand U2686 (N_2686,In_153,In_578);
and U2687 (N_2687,In_248,In_64);
nand U2688 (N_2688,In_144,In_614);
nand U2689 (N_2689,In_785,In_1176);
and U2690 (N_2690,In_416,In_815);
nor U2691 (N_2691,In_1126,In_957);
nand U2692 (N_2692,In_211,In_972);
nand U2693 (N_2693,In_1189,In_597);
nand U2694 (N_2694,In_499,In_1070);
or U2695 (N_2695,In_1103,In_1348);
or U2696 (N_2696,In_767,In_302);
nand U2697 (N_2697,In_1235,In_640);
or U2698 (N_2698,In_566,In_918);
and U2699 (N_2699,In_488,In_134);
and U2700 (N_2700,In_1325,In_489);
or U2701 (N_2701,In_97,In_1126);
or U2702 (N_2702,In_1323,In_467);
nor U2703 (N_2703,In_1414,In_1190);
or U2704 (N_2704,In_454,In_743);
and U2705 (N_2705,In_728,In_1263);
and U2706 (N_2706,In_443,In_378);
and U2707 (N_2707,In_398,In_452);
nand U2708 (N_2708,In_273,In_82);
or U2709 (N_2709,In_902,In_369);
or U2710 (N_2710,In_1393,In_325);
and U2711 (N_2711,In_291,In_1081);
nand U2712 (N_2712,In_1341,In_1230);
nand U2713 (N_2713,In_1481,In_866);
nor U2714 (N_2714,In_682,In_240);
nor U2715 (N_2715,In_489,In_401);
nor U2716 (N_2716,In_1210,In_440);
nor U2717 (N_2717,In_1193,In_264);
or U2718 (N_2718,In_1163,In_357);
or U2719 (N_2719,In_435,In_843);
nand U2720 (N_2720,In_1072,In_111);
nor U2721 (N_2721,In_1006,In_940);
nand U2722 (N_2722,In_490,In_1215);
nand U2723 (N_2723,In_1338,In_1349);
nand U2724 (N_2724,In_911,In_535);
nand U2725 (N_2725,In_68,In_1226);
nor U2726 (N_2726,In_93,In_1012);
and U2727 (N_2727,In_2,In_1248);
or U2728 (N_2728,In_1299,In_1086);
and U2729 (N_2729,In_334,In_654);
nor U2730 (N_2730,In_262,In_1170);
and U2731 (N_2731,In_549,In_110);
and U2732 (N_2732,In_33,In_159);
or U2733 (N_2733,In_923,In_372);
or U2734 (N_2734,In_1068,In_720);
and U2735 (N_2735,In_614,In_1407);
nor U2736 (N_2736,In_874,In_970);
or U2737 (N_2737,In_29,In_1080);
and U2738 (N_2738,In_916,In_673);
or U2739 (N_2739,In_985,In_230);
nor U2740 (N_2740,In_120,In_243);
and U2741 (N_2741,In_1000,In_494);
nand U2742 (N_2742,In_630,In_1395);
nand U2743 (N_2743,In_1477,In_1051);
xnor U2744 (N_2744,In_22,In_970);
or U2745 (N_2745,In_190,In_28);
nand U2746 (N_2746,In_823,In_571);
nand U2747 (N_2747,In_116,In_151);
nor U2748 (N_2748,In_1377,In_1379);
and U2749 (N_2749,In_1238,In_1292);
nand U2750 (N_2750,In_964,In_158);
nor U2751 (N_2751,In_1304,In_2);
nand U2752 (N_2752,In_1235,In_802);
and U2753 (N_2753,In_1096,In_27);
and U2754 (N_2754,In_888,In_825);
and U2755 (N_2755,In_88,In_1229);
xnor U2756 (N_2756,In_830,In_309);
nand U2757 (N_2757,In_226,In_212);
nor U2758 (N_2758,In_712,In_1286);
nor U2759 (N_2759,In_801,In_1065);
nand U2760 (N_2760,In_367,In_226);
or U2761 (N_2761,In_1263,In_1052);
nor U2762 (N_2762,In_1032,In_1233);
and U2763 (N_2763,In_1020,In_655);
and U2764 (N_2764,In_1193,In_57);
nand U2765 (N_2765,In_160,In_1038);
nor U2766 (N_2766,In_560,In_1303);
nand U2767 (N_2767,In_246,In_1399);
or U2768 (N_2768,In_110,In_1316);
nand U2769 (N_2769,In_595,In_1127);
nand U2770 (N_2770,In_662,In_820);
or U2771 (N_2771,In_85,In_1085);
and U2772 (N_2772,In_887,In_189);
and U2773 (N_2773,In_144,In_452);
or U2774 (N_2774,In_1376,In_597);
nor U2775 (N_2775,In_1453,In_1059);
or U2776 (N_2776,In_76,In_390);
or U2777 (N_2777,In_787,In_1346);
nor U2778 (N_2778,In_647,In_129);
and U2779 (N_2779,In_420,In_1061);
nor U2780 (N_2780,In_249,In_824);
nand U2781 (N_2781,In_1268,In_1489);
or U2782 (N_2782,In_1208,In_174);
or U2783 (N_2783,In_422,In_987);
or U2784 (N_2784,In_584,In_654);
or U2785 (N_2785,In_1305,In_191);
nand U2786 (N_2786,In_940,In_556);
nor U2787 (N_2787,In_1420,In_388);
nand U2788 (N_2788,In_1173,In_27);
or U2789 (N_2789,In_1081,In_372);
and U2790 (N_2790,In_768,In_76);
or U2791 (N_2791,In_467,In_592);
or U2792 (N_2792,In_747,In_603);
nand U2793 (N_2793,In_1405,In_747);
or U2794 (N_2794,In_16,In_922);
and U2795 (N_2795,In_521,In_404);
nor U2796 (N_2796,In_901,In_1274);
or U2797 (N_2797,In_373,In_582);
nand U2798 (N_2798,In_45,In_877);
or U2799 (N_2799,In_346,In_1296);
and U2800 (N_2800,In_796,In_104);
nand U2801 (N_2801,In_662,In_1131);
nand U2802 (N_2802,In_1146,In_1302);
and U2803 (N_2803,In_235,In_1440);
nor U2804 (N_2804,In_625,In_1158);
or U2805 (N_2805,In_270,In_62);
nor U2806 (N_2806,In_124,In_511);
nor U2807 (N_2807,In_1398,In_1138);
nor U2808 (N_2808,In_1467,In_423);
nor U2809 (N_2809,In_351,In_1370);
or U2810 (N_2810,In_408,In_13);
nor U2811 (N_2811,In_1121,In_879);
and U2812 (N_2812,In_545,In_786);
or U2813 (N_2813,In_260,In_1036);
and U2814 (N_2814,In_1009,In_1100);
nand U2815 (N_2815,In_1456,In_1489);
nand U2816 (N_2816,In_1468,In_812);
nand U2817 (N_2817,In_260,In_126);
and U2818 (N_2818,In_1139,In_1026);
nand U2819 (N_2819,In_1224,In_626);
nor U2820 (N_2820,In_579,In_1093);
nor U2821 (N_2821,In_735,In_253);
nor U2822 (N_2822,In_656,In_83);
nor U2823 (N_2823,In_568,In_845);
nor U2824 (N_2824,In_591,In_499);
nor U2825 (N_2825,In_732,In_975);
or U2826 (N_2826,In_1307,In_1338);
or U2827 (N_2827,In_67,In_825);
nor U2828 (N_2828,In_1010,In_296);
or U2829 (N_2829,In_1020,In_15);
nor U2830 (N_2830,In_317,In_760);
nor U2831 (N_2831,In_432,In_903);
and U2832 (N_2832,In_958,In_1213);
nand U2833 (N_2833,In_1280,In_1174);
or U2834 (N_2834,In_955,In_451);
or U2835 (N_2835,In_1382,In_955);
nand U2836 (N_2836,In_335,In_755);
nor U2837 (N_2837,In_832,In_1);
nor U2838 (N_2838,In_316,In_944);
or U2839 (N_2839,In_1428,In_811);
and U2840 (N_2840,In_744,In_1106);
nand U2841 (N_2841,In_218,In_284);
and U2842 (N_2842,In_1242,In_864);
nand U2843 (N_2843,In_335,In_807);
or U2844 (N_2844,In_1083,In_377);
or U2845 (N_2845,In_1379,In_1094);
nor U2846 (N_2846,In_7,In_1107);
nor U2847 (N_2847,In_124,In_1192);
nor U2848 (N_2848,In_294,In_278);
nand U2849 (N_2849,In_724,In_736);
nor U2850 (N_2850,In_1440,In_124);
and U2851 (N_2851,In_1196,In_83);
nor U2852 (N_2852,In_414,In_754);
nor U2853 (N_2853,In_16,In_1056);
nor U2854 (N_2854,In_573,In_594);
nor U2855 (N_2855,In_610,In_475);
nor U2856 (N_2856,In_1101,In_167);
nand U2857 (N_2857,In_915,In_477);
xor U2858 (N_2858,In_1116,In_141);
nand U2859 (N_2859,In_993,In_1386);
nand U2860 (N_2860,In_939,In_1042);
and U2861 (N_2861,In_1359,In_1443);
nor U2862 (N_2862,In_1014,In_1142);
nand U2863 (N_2863,In_231,In_1251);
nand U2864 (N_2864,In_875,In_766);
nor U2865 (N_2865,In_1126,In_1342);
nand U2866 (N_2866,In_1026,In_672);
nand U2867 (N_2867,In_69,In_182);
nor U2868 (N_2868,In_414,In_1388);
nor U2869 (N_2869,In_1012,In_1211);
nor U2870 (N_2870,In_950,In_388);
and U2871 (N_2871,In_171,In_1431);
or U2872 (N_2872,In_116,In_192);
and U2873 (N_2873,In_1341,In_741);
and U2874 (N_2874,In_1037,In_851);
nand U2875 (N_2875,In_199,In_180);
and U2876 (N_2876,In_152,In_663);
or U2877 (N_2877,In_222,In_319);
nor U2878 (N_2878,In_393,In_364);
nand U2879 (N_2879,In_1494,In_604);
or U2880 (N_2880,In_1465,In_6);
nor U2881 (N_2881,In_322,In_841);
and U2882 (N_2882,In_1420,In_137);
nor U2883 (N_2883,In_1394,In_217);
nor U2884 (N_2884,In_681,In_1069);
nand U2885 (N_2885,In_574,In_243);
nand U2886 (N_2886,In_1368,In_767);
nand U2887 (N_2887,In_1145,In_1331);
or U2888 (N_2888,In_1086,In_67);
nor U2889 (N_2889,In_1102,In_1471);
and U2890 (N_2890,In_1237,In_1315);
or U2891 (N_2891,In_54,In_440);
nor U2892 (N_2892,In_1035,In_742);
nand U2893 (N_2893,In_972,In_309);
nand U2894 (N_2894,In_1182,In_909);
nand U2895 (N_2895,In_1168,In_1224);
nor U2896 (N_2896,In_23,In_111);
nor U2897 (N_2897,In_257,In_551);
nand U2898 (N_2898,In_1436,In_746);
or U2899 (N_2899,In_950,In_1022);
or U2900 (N_2900,In_1025,In_297);
nand U2901 (N_2901,In_419,In_756);
and U2902 (N_2902,In_1141,In_73);
nand U2903 (N_2903,In_845,In_1474);
and U2904 (N_2904,In_1231,In_947);
and U2905 (N_2905,In_158,In_1265);
and U2906 (N_2906,In_366,In_1345);
or U2907 (N_2907,In_806,In_700);
and U2908 (N_2908,In_345,In_1468);
nor U2909 (N_2909,In_844,In_25);
nor U2910 (N_2910,In_1141,In_1483);
nor U2911 (N_2911,In_82,In_808);
or U2912 (N_2912,In_876,In_1460);
and U2913 (N_2913,In_1037,In_1281);
nand U2914 (N_2914,In_1445,In_466);
or U2915 (N_2915,In_824,In_1027);
xor U2916 (N_2916,In_1331,In_841);
nand U2917 (N_2917,In_422,In_981);
and U2918 (N_2918,In_254,In_579);
or U2919 (N_2919,In_27,In_553);
nand U2920 (N_2920,In_915,In_794);
or U2921 (N_2921,In_133,In_1254);
nor U2922 (N_2922,In_1100,In_1317);
nand U2923 (N_2923,In_1430,In_932);
nor U2924 (N_2924,In_878,In_1119);
nand U2925 (N_2925,In_1129,In_1128);
or U2926 (N_2926,In_1267,In_237);
and U2927 (N_2927,In_1276,In_767);
nor U2928 (N_2928,In_973,In_1362);
and U2929 (N_2929,In_914,In_121);
and U2930 (N_2930,In_599,In_547);
and U2931 (N_2931,In_440,In_973);
and U2932 (N_2932,In_581,In_599);
or U2933 (N_2933,In_1311,In_717);
nand U2934 (N_2934,In_408,In_809);
or U2935 (N_2935,In_241,In_1476);
and U2936 (N_2936,In_1325,In_1406);
nor U2937 (N_2937,In_1237,In_905);
and U2938 (N_2938,In_1018,In_1002);
or U2939 (N_2939,In_71,In_1253);
nor U2940 (N_2940,In_1398,In_1442);
nand U2941 (N_2941,In_183,In_121);
and U2942 (N_2942,In_1214,In_549);
or U2943 (N_2943,In_1103,In_616);
or U2944 (N_2944,In_1180,In_411);
nand U2945 (N_2945,In_428,In_1182);
and U2946 (N_2946,In_62,In_776);
or U2947 (N_2947,In_67,In_227);
or U2948 (N_2948,In_301,In_218);
or U2949 (N_2949,In_192,In_1173);
nand U2950 (N_2950,In_534,In_1342);
or U2951 (N_2951,In_424,In_213);
nor U2952 (N_2952,In_989,In_1115);
and U2953 (N_2953,In_973,In_1058);
and U2954 (N_2954,In_135,In_544);
nand U2955 (N_2955,In_792,In_556);
xor U2956 (N_2956,In_264,In_62);
nand U2957 (N_2957,In_1128,In_1477);
nand U2958 (N_2958,In_654,In_753);
nand U2959 (N_2959,In_446,In_409);
or U2960 (N_2960,In_1182,In_1214);
and U2961 (N_2961,In_930,In_888);
nand U2962 (N_2962,In_1313,In_351);
or U2963 (N_2963,In_1002,In_90);
nor U2964 (N_2964,In_472,In_1295);
or U2965 (N_2965,In_704,In_1118);
and U2966 (N_2966,In_984,In_820);
nor U2967 (N_2967,In_754,In_1487);
nor U2968 (N_2968,In_1422,In_1205);
xnor U2969 (N_2969,In_126,In_119);
and U2970 (N_2970,In_984,In_610);
and U2971 (N_2971,In_382,In_1343);
nor U2972 (N_2972,In_325,In_1377);
nand U2973 (N_2973,In_131,In_1101);
or U2974 (N_2974,In_1140,In_756);
nor U2975 (N_2975,In_318,In_1420);
nor U2976 (N_2976,In_464,In_1293);
nand U2977 (N_2977,In_607,In_1279);
and U2978 (N_2978,In_1448,In_127);
nand U2979 (N_2979,In_811,In_801);
and U2980 (N_2980,In_934,In_1457);
nand U2981 (N_2981,In_701,In_69);
and U2982 (N_2982,In_12,In_675);
or U2983 (N_2983,In_485,In_559);
nor U2984 (N_2984,In_926,In_280);
or U2985 (N_2985,In_616,In_947);
or U2986 (N_2986,In_876,In_1483);
nand U2987 (N_2987,In_954,In_1294);
or U2988 (N_2988,In_173,In_824);
nand U2989 (N_2989,In_446,In_253);
or U2990 (N_2990,In_626,In_958);
and U2991 (N_2991,In_126,In_262);
nor U2992 (N_2992,In_1215,In_213);
or U2993 (N_2993,In_834,In_927);
or U2994 (N_2994,In_214,In_733);
nor U2995 (N_2995,In_568,In_1232);
nor U2996 (N_2996,In_302,In_274);
nor U2997 (N_2997,In_1188,In_815);
nand U2998 (N_2998,In_1000,In_850);
and U2999 (N_2999,In_1480,In_1129);
and U3000 (N_3000,N_1673,N_2533);
nand U3001 (N_3001,N_39,N_1996);
and U3002 (N_3002,N_2317,N_2487);
and U3003 (N_3003,N_796,N_1310);
or U3004 (N_3004,N_2051,N_1038);
or U3005 (N_3005,N_1056,N_426);
nand U3006 (N_3006,N_1409,N_1121);
nand U3007 (N_3007,N_1457,N_2062);
or U3008 (N_3008,N_776,N_265);
nor U3009 (N_3009,N_1302,N_2682);
or U3010 (N_3010,N_821,N_230);
and U3011 (N_3011,N_2718,N_1988);
nor U3012 (N_3012,N_1877,N_1526);
and U3013 (N_3013,N_2626,N_1437);
and U3014 (N_3014,N_843,N_2233);
or U3015 (N_3015,N_2764,N_1402);
and U3016 (N_3016,N_2929,N_2484);
and U3017 (N_3017,N_1290,N_342);
nor U3018 (N_3018,N_177,N_1636);
nand U3019 (N_3019,N_1954,N_2958);
nand U3020 (N_3020,N_636,N_1284);
and U3021 (N_3021,N_1461,N_1130);
and U3022 (N_3022,N_2504,N_863);
or U3023 (N_3023,N_217,N_1514);
and U3024 (N_3024,N_460,N_38);
nor U3025 (N_3025,N_473,N_364);
nor U3026 (N_3026,N_2596,N_6);
or U3027 (N_3027,N_1032,N_12);
nand U3028 (N_3028,N_1852,N_1582);
and U3029 (N_3029,N_2066,N_2361);
or U3030 (N_3030,N_405,N_1239);
nand U3031 (N_3031,N_1875,N_2890);
nand U3032 (N_3032,N_2425,N_2878);
or U3033 (N_3033,N_541,N_2831);
or U3034 (N_3034,N_206,N_2248);
or U3035 (N_3035,N_714,N_2825);
or U3036 (N_3036,N_2386,N_2580);
or U3037 (N_3037,N_706,N_1844);
nand U3038 (N_3038,N_648,N_463);
or U3039 (N_3039,N_2086,N_2658);
and U3040 (N_3040,N_1640,N_2981);
nor U3041 (N_3041,N_1772,N_1676);
and U3042 (N_3042,N_25,N_995);
nand U3043 (N_3043,N_1707,N_2799);
nor U3044 (N_3044,N_2968,N_1412);
nor U3045 (N_3045,N_2322,N_1986);
and U3046 (N_3046,N_2664,N_2901);
or U3047 (N_3047,N_2720,N_2624);
nand U3048 (N_3048,N_2360,N_654);
nand U3049 (N_3049,N_1458,N_886);
nor U3050 (N_3050,N_1712,N_1711);
or U3051 (N_3051,N_1492,N_2429);
or U3052 (N_3052,N_2252,N_2090);
or U3053 (N_3053,N_2659,N_808);
nand U3054 (N_3054,N_2368,N_44);
and U3055 (N_3055,N_2271,N_539);
nor U3056 (N_3056,N_1648,N_2044);
nand U3057 (N_3057,N_170,N_2065);
nor U3058 (N_3058,N_2685,N_1163);
nor U3059 (N_3059,N_1721,N_2809);
nor U3060 (N_3060,N_1420,N_2542);
or U3061 (N_3061,N_2163,N_2672);
or U3062 (N_3062,N_2514,N_2103);
or U3063 (N_3063,N_961,N_826);
or U3064 (N_3064,N_1775,N_1375);
and U3065 (N_3065,N_2148,N_2781);
nand U3066 (N_3066,N_2684,N_178);
and U3067 (N_3067,N_1730,N_1235);
and U3068 (N_3068,N_1500,N_1270);
and U3069 (N_3069,N_2644,N_1899);
or U3070 (N_3070,N_1802,N_2378);
xnor U3071 (N_3071,N_1479,N_1311);
and U3072 (N_3072,N_453,N_1685);
xor U3073 (N_3073,N_2022,N_359);
and U3074 (N_3074,N_1193,N_2620);
nand U3075 (N_3075,N_13,N_1631);
or U3076 (N_3076,N_391,N_2277);
and U3077 (N_3077,N_978,N_2587);
nand U3078 (N_3078,N_896,N_1984);
or U3079 (N_3079,N_731,N_350);
or U3080 (N_3080,N_1401,N_2858);
or U3081 (N_3081,N_1735,N_1745);
nor U3082 (N_3082,N_2641,N_2920);
or U3083 (N_3083,N_2333,N_1814);
and U3084 (N_3084,N_2773,N_2670);
nand U3085 (N_3085,N_2726,N_2228);
nor U3086 (N_3086,N_2030,N_2731);
or U3087 (N_3087,N_2679,N_428);
nor U3088 (N_3088,N_2350,N_2199);
nor U3089 (N_3089,N_79,N_542);
or U3090 (N_3090,N_990,N_374);
nand U3091 (N_3091,N_3,N_1429);
or U3092 (N_3092,N_1257,N_410);
or U3093 (N_3093,N_2141,N_472);
or U3094 (N_3094,N_300,N_2238);
nand U3095 (N_3095,N_518,N_2394);
or U3096 (N_3096,N_2883,N_2375);
nand U3097 (N_3097,N_2827,N_1929);
and U3098 (N_3098,N_1366,N_1334);
and U3099 (N_3099,N_1450,N_640);
and U3100 (N_3100,N_2717,N_1157);
and U3101 (N_3101,N_833,N_591);
or U3102 (N_3102,N_976,N_573);
or U3103 (N_3103,N_1358,N_1556);
and U3104 (N_3104,N_2536,N_1258);
and U3105 (N_3105,N_1050,N_2565);
and U3106 (N_3106,N_256,N_432);
nor U3107 (N_3107,N_1190,N_2857);
or U3108 (N_3108,N_2205,N_127);
nor U3109 (N_3109,N_1424,N_214);
or U3110 (N_3110,N_2554,N_2454);
and U3111 (N_3111,N_2107,N_1759);
nor U3112 (N_3112,N_2266,N_2772);
or U3113 (N_3113,N_302,N_313);
or U3114 (N_3114,N_1435,N_2492);
and U3115 (N_3115,N_132,N_2821);
and U3116 (N_3116,N_1460,N_799);
or U3117 (N_3117,N_2982,N_1590);
nand U3118 (N_3118,N_1100,N_682);
nand U3119 (N_3119,N_1603,N_162);
and U3120 (N_3120,N_1208,N_2358);
or U3121 (N_3121,N_2275,N_27);
nand U3122 (N_3122,N_119,N_890);
nand U3123 (N_3123,N_114,N_2519);
and U3124 (N_3124,N_2192,N_257);
and U3125 (N_3125,N_694,N_348);
nor U3126 (N_3126,N_229,N_1166);
or U3127 (N_3127,N_1770,N_1389);
nand U3128 (N_3128,N_2026,N_946);
nor U3129 (N_3129,N_2295,N_2558);
and U3130 (N_3130,N_771,N_2279);
nor U3131 (N_3131,N_150,N_2509);
nand U3132 (N_3132,N_1146,N_1548);
and U3133 (N_3133,N_1584,N_1626);
or U3134 (N_3134,N_2833,N_2222);
or U3135 (N_3135,N_829,N_1055);
or U3136 (N_3136,N_2045,N_2769);
nand U3137 (N_3137,N_1906,N_2435);
or U3138 (N_3138,N_1918,N_2278);
nand U3139 (N_3139,N_1850,N_2806);
and U3140 (N_3140,N_567,N_1635);
xnor U3141 (N_3141,N_7,N_2481);
nand U3142 (N_3142,N_637,N_2410);
or U3143 (N_3143,N_226,N_1849);
or U3144 (N_3144,N_669,N_1233);
and U3145 (N_3145,N_2572,N_2354);
nor U3146 (N_3146,N_2113,N_400);
nor U3147 (N_3147,N_622,N_1671);
nor U3148 (N_3148,N_1755,N_2521);
and U3149 (N_3149,N_901,N_225);
or U3150 (N_3150,N_91,N_543);
nand U3151 (N_3151,N_813,N_23);
nand U3152 (N_3152,N_155,N_112);
nand U3153 (N_3153,N_739,N_2064);
or U3154 (N_3154,N_2715,N_1566);
nor U3155 (N_3155,N_1507,N_1224);
or U3156 (N_3156,N_2013,N_2910);
nor U3157 (N_3157,N_1292,N_1154);
and U3158 (N_3158,N_2766,N_2153);
nand U3159 (N_3159,N_2227,N_2170);
or U3160 (N_3160,N_1240,N_1252);
and U3161 (N_3161,N_1728,N_1747);
and U3162 (N_3162,N_371,N_2143);
nor U3163 (N_3163,N_1997,N_1909);
or U3164 (N_3164,N_2181,N_2486);
or U3165 (N_3165,N_17,N_219);
nand U3166 (N_3166,N_1612,N_2609);
or U3167 (N_3167,N_515,N_2853);
nor U3168 (N_3168,N_503,N_19);
nand U3169 (N_3169,N_152,N_1405);
nor U3170 (N_3170,N_1710,N_2423);
and U3171 (N_3171,N_2891,N_2699);
and U3172 (N_3172,N_1131,N_2401);
nand U3173 (N_3173,N_2031,N_1957);
nor U3174 (N_3174,N_1777,N_1897);
and U3175 (N_3175,N_656,N_2735);
or U3176 (N_3176,N_2837,N_1790);
nand U3177 (N_3177,N_1729,N_1468);
or U3178 (N_3178,N_420,N_22);
nand U3179 (N_3179,N_1168,N_2144);
nand U3180 (N_3180,N_2125,N_2852);
nor U3181 (N_3181,N_2357,N_1451);
nand U3182 (N_3182,N_1244,N_2632);
nand U3183 (N_3183,N_1427,N_2232);
nor U3184 (N_3184,N_1567,N_245);
and U3185 (N_3185,N_1783,N_2424);
nor U3186 (N_3186,N_282,N_171);
nor U3187 (N_3187,N_1953,N_958);
nor U3188 (N_3188,N_1198,N_1016);
nand U3189 (N_3189,N_234,N_1894);
and U3190 (N_3190,N_1000,N_14);
xnor U3191 (N_3191,N_384,N_2560);
and U3192 (N_3192,N_183,N_271);
and U3193 (N_3193,N_1336,N_956);
and U3194 (N_3194,N_766,N_811);
nand U3195 (N_3195,N_2804,N_687);
and U3196 (N_3196,N_2421,N_1028);
nand U3197 (N_3197,N_2615,N_2420);
and U3198 (N_3198,N_1717,N_2269);
nor U3199 (N_3199,N_2352,N_1051);
nand U3200 (N_3200,N_2897,N_2246);
and U3201 (N_3201,N_815,N_1335);
or U3202 (N_3202,N_1810,N_2921);
nand U3203 (N_3203,N_2527,N_2184);
nand U3204 (N_3204,N_1091,N_1364);
or U3205 (N_3205,N_2476,N_200);
and U3206 (N_3206,N_2261,N_2540);
and U3207 (N_3207,N_2061,N_2941);
nor U3208 (N_3208,N_1384,N_643);
nor U3209 (N_3209,N_467,N_1749);
nand U3210 (N_3210,N_1554,N_1155);
and U3211 (N_3211,N_729,N_2577);
nor U3212 (N_3212,N_1985,N_1162);
or U3213 (N_3213,N_1312,N_576);
and U3214 (N_3214,N_923,N_1250);
nor U3215 (N_3215,N_1023,N_2588);
nor U3216 (N_3216,N_1101,N_2946);
nor U3217 (N_3217,N_2365,N_1515);
and U3218 (N_3218,N_1724,N_2077);
and U3219 (N_3219,N_1062,N_2604);
or U3220 (N_3220,N_2256,N_2330);
nand U3221 (N_3221,N_382,N_1394);
and U3222 (N_3222,N_827,N_2979);
or U3223 (N_3223,N_1714,N_2899);
nand U3224 (N_3224,N_1498,N_2346);
nand U3225 (N_3225,N_491,N_1553);
or U3226 (N_3226,N_209,N_1277);
nor U3227 (N_3227,N_1396,N_2653);
nand U3228 (N_3228,N_2307,N_238);
nor U3229 (N_3229,N_129,N_1604);
nor U3230 (N_3230,N_1560,N_1592);
nor U3231 (N_3231,N_1605,N_2348);
nor U3232 (N_3232,N_2447,N_446);
nor U3233 (N_3233,N_2282,N_1078);
nor U3234 (N_3234,N_1361,N_1610);
and U3235 (N_3235,N_2612,N_1170);
and U3236 (N_3236,N_1977,N_508);
nand U3237 (N_3237,N_1496,N_2057);
and U3238 (N_3238,N_1187,N_1891);
or U3239 (N_3239,N_89,N_2250);
nand U3240 (N_3240,N_1314,N_2902);
and U3241 (N_3241,N_2943,N_1008);
or U3242 (N_3242,N_2241,N_149);
nand U3243 (N_3243,N_207,N_1029);
nor U3244 (N_3244,N_2950,N_2513);
nor U3245 (N_3245,N_660,N_1669);
or U3246 (N_3246,N_2725,N_969);
and U3247 (N_3247,N_1150,N_2006);
and U3248 (N_3248,N_727,N_2570);
or U3249 (N_3249,N_719,N_1663);
or U3250 (N_3250,N_2099,N_1249);
or U3251 (N_3251,N_233,N_1332);
nor U3252 (N_3252,N_2647,N_476);
or U3253 (N_3253,N_2582,N_699);
nor U3254 (N_3254,N_2089,N_980);
nor U3255 (N_3255,N_2854,N_1666);
nand U3256 (N_3256,N_488,N_2996);
nor U3257 (N_3257,N_2067,N_318);
or U3258 (N_3258,N_942,N_2004);
or U3259 (N_3259,N_2473,N_1818);
and U3260 (N_3260,N_101,N_2529);
nor U3261 (N_3261,N_2997,N_1944);
nor U3262 (N_3262,N_2888,N_2047);
nand U3263 (N_3263,N_2614,N_1768);
or U3264 (N_3264,N_659,N_2092);
nor U3265 (N_3265,N_370,N_2984);
or U3266 (N_3266,N_1497,N_565);
nand U3267 (N_3267,N_666,N_1319);
or U3268 (N_3268,N_1153,N_2942);
nor U3269 (N_3269,N_871,N_1992);
or U3270 (N_3270,N_560,N_2539);
nor U3271 (N_3271,N_2200,N_639);
nand U3272 (N_3272,N_2505,N_2722);
nor U3273 (N_3273,N_509,N_1798);
nor U3274 (N_3274,N_298,N_592);
xnor U3275 (N_3275,N_2127,N_1732);
nor U3276 (N_3276,N_145,N_1385);
or U3277 (N_3277,N_2312,N_2347);
and U3278 (N_3278,N_224,N_55);
or U3279 (N_3279,N_2571,N_2165);
nor U3280 (N_3280,N_1737,N_1822);
and U3281 (N_3281,N_2616,N_2801);
nor U3282 (N_3282,N_250,N_450);
and U3283 (N_3283,N_1423,N_2060);
or U3284 (N_3284,N_2007,N_981);
and U3285 (N_3285,N_605,N_2733);
nand U3286 (N_3286,N_2151,N_2563);
and U3287 (N_3287,N_803,N_2071);
or U3288 (N_3288,N_2448,N_1120);
or U3289 (N_3289,N_1439,N_1159);
nor U3290 (N_3290,N_293,N_1134);
nand U3291 (N_3291,N_1718,N_1328);
and U3292 (N_3292,N_33,N_1539);
nor U3293 (N_3293,N_2585,N_1585);
and U3294 (N_3294,N_545,N_75);
and U3295 (N_3295,N_2353,N_2972);
nor U3296 (N_3296,N_1709,N_1470);
and U3297 (N_3297,N_1386,N_1081);
nor U3298 (N_3298,N_1327,N_2290);
nand U3299 (N_3299,N_667,N_1246);
or U3300 (N_3300,N_1620,N_1045);
or U3301 (N_3301,N_2667,N_54);
nor U3302 (N_3302,N_710,N_435);
nor U3303 (N_3303,N_2705,N_661);
nor U3304 (N_3304,N_2270,N_2046);
nor U3305 (N_3305,N_1180,N_2948);
nand U3306 (N_3306,N_303,N_1473);
nor U3307 (N_3307,N_2373,N_2191);
and U3308 (N_3308,N_421,N_1531);
nand U3309 (N_3309,N_239,N_1148);
nor U3310 (N_3310,N_1693,N_103);
nor U3311 (N_3311,N_1086,N_236);
nand U3312 (N_3312,N_201,N_2074);
or U3313 (N_3313,N_126,N_764);
nor U3314 (N_3314,N_1015,N_2597);
nor U3315 (N_3315,N_2157,N_1882);
nor U3316 (N_3316,N_1880,N_903);
and U3317 (N_3317,N_2146,N_2754);
nor U3318 (N_3318,N_2818,N_2247);
nand U3319 (N_3319,N_470,N_1917);
or U3320 (N_3320,N_1087,N_1811);
and U3321 (N_3321,N_1521,N_1670);
or U3322 (N_3322,N_154,N_865);
and U3323 (N_3323,N_2949,N_35);
nand U3324 (N_3324,N_1762,N_1268);
or U3325 (N_3325,N_1456,N_1549);
nand U3326 (N_3326,N_153,N_212);
nor U3327 (N_3327,N_1807,N_2311);
or U3328 (N_3328,N_1065,N_2055);
or U3329 (N_3329,N_862,N_235);
or U3330 (N_3330,N_1757,N_1504);
nor U3331 (N_3331,N_2223,N_320);
nor U3332 (N_3332,N_2712,N_2161);
and U3333 (N_3333,N_418,N_736);
or U3334 (N_3334,N_2656,N_2121);
nand U3335 (N_3335,N_1483,N_1588);
nor U3336 (N_3336,N_1939,N_1838);
and U3337 (N_3337,N_2477,N_2914);
and U3338 (N_3338,N_423,N_1408);
nand U3339 (N_3339,N_2328,N_276);
nor U3340 (N_3340,N_1994,N_383);
nand U3341 (N_3341,N_2633,N_357);
or U3342 (N_3342,N_1524,N_2169);
nor U3343 (N_3343,N_1647,N_1191);
nor U3344 (N_3344,N_417,N_671);
and U3345 (N_3345,N_959,N_1188);
and U3346 (N_3346,N_46,N_2072);
nor U3347 (N_3347,N_895,N_2451);
or U3348 (N_3348,N_2440,N_294);
nand U3349 (N_3349,N_629,N_2158);
and U3350 (N_3350,N_452,N_1021);
nor U3351 (N_3351,N_864,N_1383);
and U3352 (N_3352,N_2384,N_1975);
nand U3353 (N_3353,N_603,N_787);
nand U3354 (N_3354,N_1934,N_1967);
nor U3355 (N_3355,N_1534,N_1726);
nand U3356 (N_3356,N_1309,N_1214);
or U3357 (N_3357,N_1202,N_952);
and U3358 (N_3358,N_1002,N_2042);
nor U3359 (N_3359,N_2627,N_1067);
nand U3360 (N_3360,N_2048,N_602);
and U3361 (N_3361,N_2452,N_1700);
and U3362 (N_3362,N_819,N_451);
nand U3363 (N_3363,N_692,N_1981);
nand U3364 (N_3364,N_1758,N_621);
or U3365 (N_3365,N_477,N_2172);
nor U3366 (N_3366,N_1307,N_2418);
and U3367 (N_3367,N_273,N_1990);
xnor U3368 (N_3368,N_697,N_93);
and U3369 (N_3369,N_1184,N_850);
and U3370 (N_3370,N_1893,N_8);
nand U3371 (N_3371,N_63,N_1158);
nor U3372 (N_3372,N_2276,N_1106);
nor U3373 (N_3373,N_2376,N_1847);
and U3374 (N_3374,N_2613,N_984);
or U3375 (N_3375,N_2651,N_809);
nand U3376 (N_3376,N_1491,N_193);
nand U3377 (N_3377,N_2525,N_2027);
nand U3378 (N_3378,N_386,N_2990);
and U3379 (N_3379,N_544,N_2518);
nand U3380 (N_3380,N_2498,N_2009);
nand U3381 (N_3381,N_2245,N_760);
and U3382 (N_3382,N_802,N_1010);
or U3383 (N_3383,N_2324,N_1020);
or U3384 (N_3384,N_1857,N_2075);
and U3385 (N_3385,N_994,N_2268);
or U3386 (N_3386,N_572,N_1256);
and U3387 (N_3387,N_498,N_242);
or U3388 (N_3388,N_689,N_98);
nor U3389 (N_3389,N_2218,N_1704);
and U3390 (N_3390,N_2339,N_2267);
nand U3391 (N_3391,N_354,N_454);
and U3392 (N_3392,N_2621,N_480);
and U3393 (N_3393,N_2532,N_2868);
nor U3394 (N_3394,N_2584,N_204);
or U3395 (N_3395,N_2016,N_2922);
and U3396 (N_3396,N_1708,N_1097);
or U3397 (N_3397,N_2224,N_1035);
nand U3398 (N_3398,N_1506,N_2931);
and U3399 (N_3399,N_2162,N_389);
nand U3400 (N_3400,N_2342,N_2412);
nand U3401 (N_3401,N_1831,N_199);
and U3402 (N_3402,N_74,N_168);
or U3403 (N_3403,N_2179,N_2955);
or U3404 (N_3404,N_2872,N_50);
or U3405 (N_3405,N_249,N_810);
or U3406 (N_3406,N_2230,N_254);
and U3407 (N_3407,N_1776,N_1200);
nor U3408 (N_3408,N_156,N_2713);
nor U3409 (N_3409,N_1641,N_2916);
or U3410 (N_3410,N_823,N_381);
nand U3411 (N_3411,N_2895,N_324);
nand U3412 (N_3412,N_392,N_1574);
and U3413 (N_3413,N_2742,N_1616);
or U3414 (N_3414,N_1298,N_1487);
nor U3415 (N_3415,N_2093,N_322);
nand U3416 (N_3416,N_2028,N_48);
and U3417 (N_3417,N_2344,N_1551);
nor U3418 (N_3418,N_1446,N_1808);
or U3419 (N_3419,N_1699,N_1733);
nand U3420 (N_3420,N_2262,N_71);
and U3421 (N_3421,N_2041,N_311);
nor U3422 (N_3422,N_30,N_2973);
and U3423 (N_3423,N_2779,N_161);
and U3424 (N_3424,N_2555,N_1681);
or U3425 (N_3425,N_1901,N_1922);
nand U3426 (N_3426,N_2810,N_2195);
or U3427 (N_3427,N_2874,N_2839);
or U3428 (N_3428,N_613,N_2683);
or U3429 (N_3429,N_1508,N_1895);
or U3430 (N_3430,N_1480,N_241);
nand U3431 (N_3431,N_2755,N_992);
xnor U3432 (N_3432,N_828,N_676);
or U3433 (N_3433,N_2272,N_2650);
nand U3434 (N_3434,N_1927,N_1443);
or U3435 (N_3435,N_1340,N_712);
nand U3436 (N_3436,N_2194,N_705);
nand U3437 (N_3437,N_1675,N_2496);
and U3438 (N_3438,N_1436,N_2130);
or U3439 (N_3439,N_1825,N_847);
and U3440 (N_3440,N_741,N_1377);
and U3441 (N_3441,N_1305,N_2636);
and U3442 (N_3442,N_1824,N_2419);
and U3443 (N_3443,N_2300,N_1474);
nand U3444 (N_3444,N_2574,N_2017);
or U3445 (N_3445,N_2945,N_938);
nor U3446 (N_3446,N_1668,N_1122);
and U3447 (N_3447,N_1274,N_921);
or U3448 (N_3448,N_2673,N_1528);
and U3449 (N_3449,N_1318,N_558);
or U3450 (N_3450,N_910,N_2594);
nor U3451 (N_3451,N_1189,N_2782);
nand U3452 (N_3452,N_1611,N_1090);
or U3453 (N_3453,N_2649,N_2428);
or U3454 (N_3454,N_465,N_1989);
nor U3455 (N_3455,N_936,N_385);
and U3456 (N_3456,N_1207,N_1085);
nand U3457 (N_3457,N_610,N_2033);
xor U3458 (N_3458,N_1209,N_596);
nand U3459 (N_3459,N_606,N_29);
nor U3460 (N_3460,N_1232,N_28);
or U3461 (N_3461,N_2315,N_335);
or U3462 (N_3462,N_718,N_562);
nor U3463 (N_3463,N_120,N_1978);
nor U3464 (N_3464,N_587,N_2349);
and U3465 (N_3465,N_2434,N_2078);
and U3466 (N_3466,N_1452,N_180);
or U3467 (N_3467,N_2020,N_340);
nand U3468 (N_3468,N_1837,N_550);
nor U3469 (N_3469,N_931,N_534);
nand U3470 (N_3470,N_2959,N_1255);
nand U3471 (N_3471,N_1476,N_1112);
or U3472 (N_3472,N_1805,N_447);
nand U3473 (N_3473,N_2770,N_1971);
nor U3474 (N_3474,N_36,N_2953);
nand U3475 (N_3475,N_2204,N_1784);
nor U3476 (N_3476,N_1260,N_1963);
nor U3477 (N_3477,N_2453,N_0);
nand U3478 (N_3478,N_272,N_2912);
nor U3479 (N_3479,N_1321,N_569);
nand U3480 (N_3480,N_2791,N_379);
nor U3481 (N_3481,N_1806,N_2038);
and U3482 (N_3482,N_41,N_2557);
and U3483 (N_3483,N_1475,N_678);
and U3484 (N_3484,N_2431,N_554);
and U3485 (N_3485,N_1127,N_619);
nor U3486 (N_3486,N_2135,N_2925);
or U3487 (N_3487,N_116,N_975);
and U3488 (N_3488,N_685,N_11);
and U3489 (N_3489,N_944,N_970);
and U3490 (N_3490,N_1195,N_582);
nand U3491 (N_3491,N_1471,N_1980);
or U3492 (N_3492,N_1650,N_2965);
nor U3493 (N_3493,N_1621,N_1441);
nand U3494 (N_3494,N_1734,N_1013);
nand U3495 (N_3495,N_2466,N_2550);
and U3496 (N_3496,N_2189,N_2383);
nor U3497 (N_3497,N_726,N_1564);
and U3498 (N_3498,N_2652,N_1835);
or U3499 (N_3499,N_2108,N_547);
and U3500 (N_3500,N_1266,N_2904);
nor U3501 (N_3501,N_2395,N_424);
nor U3502 (N_3502,N_1522,N_1279);
and U3503 (N_3503,N_2390,N_60);
and U3504 (N_3504,N_128,N_2178);
or U3505 (N_3505,N_1464,N_1596);
or U3506 (N_3506,N_844,N_873);
nor U3507 (N_3507,N_1365,N_485);
nor U3508 (N_3508,N_2927,N_504);
nand U3509 (N_3509,N_2744,N_1046);
and U3510 (N_3510,N_2019,N_2721);
nor U3511 (N_3511,N_2701,N_1890);
xor U3512 (N_3512,N_722,N_927);
nand U3513 (N_3513,N_1296,N_1581);
or U3514 (N_3514,N_2050,N_1501);
or U3515 (N_3515,N_2214,N_577);
and U3516 (N_3516,N_2828,N_872);
nand U3517 (N_3517,N_1855,N_775);
or U3518 (N_3518,N_1892,N_2171);
and U3519 (N_3519,N_2678,N_306);
nand U3520 (N_3520,N_941,N_1915);
and U3521 (N_3521,N_2906,N_1813);
and U3522 (N_3522,N_1819,N_1294);
or U3523 (N_3523,N_59,N_247);
and U3524 (N_3524,N_2082,N_651);
nor U3525 (N_3525,N_2399,N_2287);
and U3526 (N_3526,N_2080,N_1623);
nand U3527 (N_3527,N_2759,N_548);
nand U3528 (N_3528,N_2882,N_1902);
and U3529 (N_3529,N_1799,N_2302);
nor U3530 (N_3530,N_2102,N_213);
nand U3531 (N_3531,N_1943,N_1143);
or U3532 (N_3532,N_260,N_1466);
nand U3533 (N_3533,N_2296,N_716);
nand U3534 (N_3534,N_494,N_1525);
nand U3535 (N_3535,N_2217,N_2154);
nand U3536 (N_3536,N_877,N_2562);
and U3537 (N_3537,N_695,N_2559);
nand U3538 (N_3538,N_2928,N_1215);
nand U3539 (N_3539,N_2417,N_1686);
or U3540 (N_3540,N_96,N_763);
nor U3541 (N_3541,N_100,N_1791);
and U3542 (N_3542,N_174,N_1025);
and U3543 (N_3543,N_1779,N_2689);
nand U3544 (N_3544,N_1126,N_1469);
or U3545 (N_3545,N_2193,N_1039);
and U3546 (N_3546,N_1337,N_1371);
and U3547 (N_3547,N_1058,N_1493);
or U3548 (N_3548,N_1628,N_2793);
and U3549 (N_3549,N_2483,N_1350);
nor U3550 (N_3550,N_2124,N_2128);
nor U3551 (N_3551,N_1118,N_626);
or U3552 (N_3552,N_797,N_85);
and U3553 (N_3553,N_2131,N_90);
and U3554 (N_3554,N_1921,N_2085);
nor U3555 (N_3555,N_1467,N_2001);
nor U3556 (N_3556,N_1826,N_2599);
or U3557 (N_3557,N_402,N_1653);
and U3558 (N_3558,N_590,N_1961);
nand U3559 (N_3559,N_2589,N_31);
and U3560 (N_3560,N_474,N_2601);
or U3561 (N_3561,N_268,N_2364);
or U3562 (N_3562,N_595,N_1459);
nand U3563 (N_3563,N_861,N_1731);
nor U3564 (N_3564,N_1346,N_986);
and U3565 (N_3565,N_1253,N_2011);
or U3566 (N_3566,N_1027,N_701);
and U3567 (N_3567,N_2538,N_880);
and U3568 (N_3568,N_1173,N_2894);
or U3569 (N_3569,N_713,N_367);
nor U3570 (N_3570,N_918,N_2905);
or U3571 (N_3571,N_2441,N_684);
nand U3572 (N_3572,N_1177,N_917);
nand U3573 (N_3573,N_468,N_1786);
nor U3574 (N_3574,N_658,N_2933);
and U3575 (N_3575,N_2700,N_2511);
nand U3576 (N_3576,N_2993,N_793);
nor U3577 (N_3577,N_691,N_1833);
and U3578 (N_3578,N_1341,N_2416);
or U3579 (N_3579,N_778,N_1715);
and U3580 (N_3580,N_618,N_1012);
or U3581 (N_3581,N_2002,N_1949);
and U3582 (N_3582,N_2753,N_1651);
and U3583 (N_3583,N_1804,N_407);
nand U3584 (N_3584,N_1387,N_274);
nor U3585 (N_3585,N_2788,N_2219);
and U3586 (N_3586,N_507,N_72);
or U3587 (N_3587,N_1503,N_502);
or U3588 (N_3588,N_2260,N_2152);
and U3589 (N_3589,N_1739,N_223);
or U3590 (N_3590,N_1904,N_593);
or U3591 (N_3591,N_1511,N_1391);
and U3592 (N_3592,N_1428,N_1555);
nand U3593 (N_3593,N_1049,N_777);
and U3594 (N_3594,N_939,N_2243);
and U3595 (N_3595,N_2457,N_2859);
nand U3596 (N_3596,N_814,N_1164);
nor U3597 (N_3597,N_1956,N_909);
or U3598 (N_3598,N_1933,N_1014);
and U3599 (N_3599,N_773,N_2708);
and U3600 (N_3600,N_2635,N_2526);
nor U3601 (N_3601,N_2400,N_2462);
and U3602 (N_3602,N_1006,N_1059);
and U3603 (N_3603,N_1455,N_172);
or U3604 (N_3604,N_2063,N_2472);
and U3605 (N_3605,N_277,N_589);
nor U3606 (N_3606,N_356,N_540);
nor U3607 (N_3607,N_645,N_2114);
nand U3608 (N_3608,N_1499,N_2798);
nand U3609 (N_3609,N_2710,N_954);
nor U3610 (N_3610,N_1238,N_2992);
and U3611 (N_3611,N_831,N_1218);
nor U3612 (N_3612,N_1317,N_2807);
or U3613 (N_3613,N_326,N_1950);
nor U3614 (N_3614,N_86,N_2388);
or U3615 (N_3615,N_1286,N_1823);
nand U3616 (N_3616,N_2284,N_2379);
nor U3617 (N_3617,N_738,N_1787);
nor U3618 (N_3618,N_1231,N_523);
xor U3619 (N_3619,N_1970,N_2617);
nand U3620 (N_3620,N_94,N_967);
or U3621 (N_3621,N_2355,N_2479);
xnor U3622 (N_3622,N_2321,N_1174);
or U3623 (N_3623,N_2639,N_425);
nor U3624 (N_3624,N_905,N_2334);
nor U3625 (N_3625,N_2593,N_840);
nand U3626 (N_3626,N_1987,N_611);
or U3627 (N_3627,N_788,N_993);
and U3628 (N_3628,N_533,N_1264);
nor U3629 (N_3629,N_1338,N_1472);
xnor U3630 (N_3630,N_538,N_1416);
nand U3631 (N_3631,N_856,N_2414);
or U3632 (N_3632,N_2187,N_1430);
or U3633 (N_3633,N_757,N_2787);
or U3634 (N_3634,N_1932,N_1293);
or U3635 (N_3635,N_2814,N_1754);
nand U3636 (N_3636,N_513,N_1107);
nor U3637 (N_3637,N_1178,N_1597);
nor U3638 (N_3638,N_588,N_316);
nand U3639 (N_3639,N_2698,N_702);
nand U3640 (N_3640,N_372,N_2029);
or U3641 (N_3641,N_1962,N_2693);
and U3642 (N_3642,N_1969,N_1397);
nor U3643 (N_3643,N_434,N_1854);
or U3644 (N_3644,N_309,N_1414);
or U3645 (N_3645,N_499,N_1517);
or U3646 (N_3646,N_144,N_279);
xor U3647 (N_3647,N_1518,N_117);
or U3648 (N_3648,N_2785,N_1089);
nand U3649 (N_3649,N_1509,N_2748);
nand U3650 (N_3650,N_1952,N_1354);
and U3651 (N_3651,N_2966,N_2547);
and U3652 (N_3652,N_529,N_1259);
and U3653 (N_3653,N_1053,N_1339);
and U3654 (N_3654,N_743,N_369);
or U3655 (N_3655,N_2215,N_1692);
and U3656 (N_3656,N_937,N_2797);
nor U3657 (N_3657,N_1993,N_1353);
nor U3658 (N_3658,N_1868,N_2081);
nand U3659 (N_3659,N_1613,N_283);
nand U3660 (N_3660,N_1194,N_1165);
and U3661 (N_3661,N_1516,N_1746);
and U3662 (N_3662,N_1236,N_2520);
nor U3663 (N_3663,N_2319,N_734);
and U3664 (N_3664,N_1017,N_2129);
nand U3665 (N_3665,N_974,N_2449);
and U3666 (N_3666,N_390,N_950);
or U3667 (N_3667,N_263,N_1716);
nor U3668 (N_3668,N_1774,N_1068);
and U3669 (N_3669,N_1672,N_377);
nand U3670 (N_3670,N_1440,N_780);
nor U3671 (N_3671,N_2913,N_1966);
nand U3672 (N_3672,N_49,N_1362);
and U3673 (N_3673,N_2727,N_674);
nor U3674 (N_3674,N_563,N_478);
or U3675 (N_3675,N_1513,N_1767);
nor U3676 (N_3676,N_1325,N_1713);
or U3677 (N_3677,N_2091,N_908);
and U3678 (N_3678,N_662,N_1009);
nand U3679 (N_3679,N_1282,N_210);
nand U3680 (N_3680,N_2734,N_960);
and U3681 (N_3681,N_2991,N_848);
nand U3682 (N_3682,N_730,N_1976);
and U3683 (N_3683,N_2488,N_2654);
nor U3684 (N_3684,N_395,N_80);
nor U3685 (N_3685,N_339,N_2567);
nor U3686 (N_3686,N_527,N_2908);
nand U3687 (N_3687,N_216,N_52);
nor U3688 (N_3688,N_2323,N_2024);
nand U3689 (N_3689,N_2954,N_2776);
or U3690 (N_3690,N_2490,N_1948);
nand U3691 (N_3691,N_1689,N_2778);
and U3692 (N_3692,N_299,N_1829);
nor U3693 (N_3693,N_786,N_414);
or U3694 (N_3694,N_2808,N_1182);
or U3695 (N_3695,N_222,N_1679);
and U3696 (N_3696,N_2335,N_1481);
or U3697 (N_3697,N_487,N_2625);
or U3698 (N_3698,N_2889,N_148);
or U3699 (N_3699,N_1557,N_2264);
nor U3700 (N_3700,N_1351,N_1222);
nand U3701 (N_3701,N_345,N_262);
nand U3702 (N_3702,N_2122,N_526);
nand U3703 (N_3703,N_1109,N_124);
nor U3704 (N_3704,N_438,N_1372);
and U3705 (N_3705,N_69,N_1761);
nor U3706 (N_3706,N_1304,N_2068);
and U3707 (N_3707,N_2815,N_1660);
nor U3708 (N_3708,N_583,N_2543);
or U3709 (N_3709,N_436,N_655);
and U3710 (N_3710,N_1789,N_1349);
and U3711 (N_3711,N_1907,N_999);
xnor U3712 (N_3712,N_2464,N_1579);
nor U3713 (N_3713,N_920,N_769);
and U3714 (N_3714,N_2745,N_2840);
nor U3715 (N_3715,N_1167,N_2283);
and U3716 (N_3716,N_2254,N_2470);
nand U3717 (N_3717,N_141,N_1295);
and U3718 (N_3718,N_581,N_1937);
nand U3719 (N_3719,N_9,N_982);
nand U3720 (N_3720,N_416,N_2919);
nor U3721 (N_3721,N_2917,N_2012);
nor U3722 (N_3722,N_900,N_2716);
and U3723 (N_3723,N_2608,N_1380);
nor U3724 (N_3724,N_388,N_2957);
or U3725 (N_3725,N_1599,N_2677);
nor U3726 (N_3726,N_882,N_612);
nor U3727 (N_3727,N_2740,N_1417);
xor U3728 (N_3728,N_800,N_1465);
and U3729 (N_3729,N_830,N_2098);
nand U3730 (N_3730,N_744,N_922);
nor U3731 (N_3731,N_57,N_2049);
and U3732 (N_3732,N_1546,N_1129);
and U3733 (N_3733,N_586,N_789);
nor U3734 (N_3734,N_2054,N_2611);
or U3735 (N_3735,N_2499,N_987);
and U3736 (N_3736,N_2474,N_1869);
or U3737 (N_3737,N_2497,N_1771);
xnor U3738 (N_3738,N_1422,N_2149);
xnor U3739 (N_3739,N_1103,N_1931);
nor U3740 (N_3740,N_2478,N_2320);
nand U3741 (N_3741,N_2073,N_2834);
nand U3742 (N_3742,N_1145,N_4);
or U3743 (N_3743,N_2010,N_1186);
nand U3744 (N_3744,N_2036,N_107);
or U3745 (N_3745,N_1541,N_1830);
nand U3746 (N_3746,N_1690,N_1703);
nand U3747 (N_3747,N_2747,N_1520);
and U3748 (N_3748,N_2545,N_1096);
nand U3749 (N_3749,N_663,N_794);
and U3750 (N_3750,N_2095,N_289);
and U3751 (N_3751,N_2468,N_1269);
nor U3752 (N_3752,N_2824,N_568);
and U3753 (N_3753,N_2396,N_798);
nor U3754 (N_3754,N_243,N_1098);
and U3755 (N_3755,N_146,N_2578);
nor U3756 (N_3756,N_1617,N_867);
xnor U3757 (N_3757,N_105,N_715);
or U3758 (N_3758,N_1695,N_2869);
and U3759 (N_3759,N_1645,N_2535);
and U3760 (N_3760,N_185,N_73);
nor U3761 (N_3761,N_1535,N_1723);
and U3762 (N_3762,N_1303,N_2469);
and U3763 (N_3763,N_1076,N_1054);
or U3764 (N_3764,N_2226,N_894);
or U3765 (N_3765,N_849,N_1743);
or U3766 (N_3766,N_2591,N_1543);
or U3767 (N_3767,N_208,N_1530);
or U3768 (N_3768,N_2553,N_1495);
and U3769 (N_3769,N_2281,N_1225);
xnor U3770 (N_3770,N_1324,N_2998);
nor U3771 (N_3771,N_2823,N_244);
or U3772 (N_3772,N_1860,N_160);
nor U3773 (N_3773,N_679,N_2768);
or U3774 (N_3774,N_2690,N_1320);
and U3775 (N_3775,N_1674,N_1356);
nor U3776 (N_3776,N_1552,N_68);
nor U3777 (N_3777,N_1136,N_1742);
nand U3778 (N_3778,N_1821,N_904);
nor U3779 (N_3779,N_2325,N_18);
nor U3780 (N_3780,N_1661,N_2637);
and U3781 (N_3781,N_1572,N_2021);
nand U3782 (N_3782,N_142,N_912);
nand U3783 (N_3783,N_448,N_2147);
xnor U3784 (N_3784,N_2995,N_373);
nor U3785 (N_3785,N_2491,N_1418);
or U3786 (N_3786,N_1586,N_2739);
and U3787 (N_3787,N_58,N_475);
or U3788 (N_3788,N_1580,N_2628);
nand U3789 (N_3789,N_228,N_2963);
nand U3790 (N_3790,N_2746,N_1803);
xnor U3791 (N_3791,N_2164,N_624);
nand U3792 (N_3792,N_2871,N_2777);
nand U3793 (N_3793,N_2409,N_2887);
and U3794 (N_3794,N_887,N_1179);
nor U3795 (N_3795,N_653,N_1433);
or U3796 (N_3796,N_2829,N_638);
and U3797 (N_3797,N_211,N_2926);
and U3798 (N_3798,N_881,N_761);
or U3799 (N_3799,N_412,N_792);
or U3800 (N_3800,N_1449,N_66);
or U3801 (N_3801,N_1910,N_2475);
or U3802 (N_3802,N_2789,N_147);
or U3803 (N_3803,N_319,N_2456);
nor U3804 (N_3804,N_2534,N_1896);
nand U3805 (N_3805,N_2439,N_329);
and U3806 (N_3806,N_1840,N_1308);
and U3807 (N_3807,N_1602,N_1979);
nor U3808 (N_3808,N_623,N_968);
or U3809 (N_3809,N_615,N_102);
nor U3810 (N_3810,N_735,N_1958);
nand U3811 (N_3811,N_403,N_2573);
nand U3812 (N_3812,N_1221,N_753);
nand U3813 (N_3813,N_2035,N_2502);
nand U3814 (N_3814,N_1884,N_2079);
nor U3815 (N_3815,N_1741,N_2730);
or U3816 (N_3816,N_1001,N_396);
and U3817 (N_3817,N_2728,N_394);
or U3818 (N_3818,N_2059,N_1033);
nor U3819 (N_3819,N_361,N_2372);
nand U3820 (N_3820,N_195,N_988);
or U3821 (N_3821,N_2552,N_297);
nor U3822 (N_3822,N_884,N_1390);
and U3823 (N_3823,N_21,N_1593);
or U3824 (N_3824,N_681,N_2706);
and U3825 (N_3825,N_2155,N_442);
nand U3826 (N_3826,N_879,N_5);
nor U3827 (N_3827,N_1928,N_1359);
nor U3828 (N_3828,N_437,N_2971);
or U3829 (N_3829,N_2118,N_2522);
or U3830 (N_3830,N_2643,N_2115);
or U3831 (N_3831,N_288,N_1267);
nand U3832 (N_3832,N_1750,N_2516);
or U3833 (N_3833,N_269,N_500);
nor U3834 (N_3834,N_2326,N_834);
nor U3835 (N_3835,N_205,N_125);
nor U3836 (N_3836,N_2835,N_2316);
nand U3837 (N_3837,N_580,N_431);
nor U3838 (N_3838,N_2318,N_947);
nand U3839 (N_3839,N_2210,N_2738);
or U3840 (N_3840,N_2900,N_1614);
nor U3841 (N_3841,N_1348,N_883);
nor U3842 (N_3842,N_358,N_331);
nor U3843 (N_3843,N_341,N_1099);
nor U3844 (N_3844,N_2736,N_1242);
or U3845 (N_3845,N_88,N_1773);
xnor U3846 (N_3846,N_2314,N_1316);
and U3847 (N_3847,N_1425,N_1889);
nand U3848 (N_3848,N_2743,N_854);
or U3849 (N_3849,N_1919,N_139);
and U3850 (N_3850,N_675,N_2397);
and U3851 (N_3851,N_2084,N_2803);
or U3852 (N_3852,N_307,N_644);
or U3853 (N_3853,N_16,N_330);
and U3854 (N_3854,N_115,N_2458);
or U3855 (N_3855,N_37,N_1908);
xor U3856 (N_3856,N_511,N_2579);
nand U3857 (N_3857,N_2980,N_248);
nand U3858 (N_3858,N_259,N_747);
and U3859 (N_3859,N_2236,N_2911);
and U3860 (N_3860,N_1071,N_1633);
nor U3861 (N_3861,N_855,N_551);
nor U3862 (N_3862,N_1486,N_1760);
nor U3863 (N_3863,N_2583,N_2947);
nand U3864 (N_3864,N_2240,N_1228);
or U3865 (N_3865,N_258,N_1344);
and U3866 (N_3866,N_2805,N_783);
nor U3867 (N_3867,N_2263,N_700);
and U3868 (N_3868,N_665,N_346);
and U3869 (N_3869,N_686,N_1945);
nor U3870 (N_3870,N_77,N_1756);
nand U3871 (N_3871,N_444,N_585);
nand U3872 (N_3872,N_1550,N_2817);
nand U3873 (N_3873,N_1083,N_1104);
nand U3874 (N_3874,N_1538,N_1662);
and U3875 (N_3875,N_2438,N_167);
xnor U3876 (N_3876,N_1769,N_2251);
nor U3877 (N_3877,N_1227,N_1237);
or U3878 (N_3878,N_2413,N_971);
and U3879 (N_3879,N_360,N_2043);
nor U3880 (N_3880,N_600,N_190);
nor U3881 (N_3881,N_1637,N_2640);
and U3882 (N_3882,N_1738,N_740);
or U3883 (N_3883,N_123,N_1080);
and U3884 (N_3884,N_1780,N_1748);
and U3885 (N_3885,N_1141,N_2123);
and U3886 (N_3886,N_720,N_176);
or U3887 (N_3887,N_181,N_2568);
and U3888 (N_3888,N_492,N_2999);
and U3889 (N_3889,N_1084,N_1419);
or U3890 (N_3890,N_1871,N_2402);
and U3891 (N_3891,N_2802,N_1094);
or U3892 (N_3892,N_1935,N_1982);
nand U3893 (N_3893,N_275,N_721);
nor U3894 (N_3894,N_1665,N_221);
or U3895 (N_3895,N_1794,N_2259);
nand U3896 (N_3896,N_165,N_220);
and U3897 (N_3897,N_1478,N_2544);
nor U3898 (N_3898,N_2120,N_584);
or U3899 (N_3899,N_532,N_2209);
and U3900 (N_3900,N_1911,N_1589);
and U3901 (N_3901,N_62,N_996);
or U3902 (N_3902,N_1367,N_2737);
nor U3903 (N_3903,N_496,N_1697);
nand U3904 (N_3904,N_943,N_1138);
or U3905 (N_3905,N_1370,N_2489);
or U3906 (N_3906,N_1477,N_2436);
or U3907 (N_3907,N_198,N_1876);
nand U3908 (N_3908,N_707,N_443);
or U3909 (N_3909,N_404,N_1034);
nand U3910 (N_3910,N_2437,N_1037);
and U3911 (N_3911,N_688,N_2935);
or U3912 (N_3912,N_1569,N_312);
nand U3913 (N_3913,N_1151,N_2934);
nor U3914 (N_3914,N_709,N_64);
nand U3915 (N_3915,N_2687,N_698);
or U3916 (N_3916,N_599,N_1415);
or U3917 (N_3917,N_2212,N_1974);
nand U3918 (N_3918,N_1275,N_2106);
and U3919 (N_3919,N_2630,N_2918);
nor U3920 (N_3920,N_774,N_2337);
nand U3921 (N_3921,N_2830,N_2188);
nor U3922 (N_3922,N_1485,N_1658);
nor U3923 (N_3923,N_2105,N_925);
nor U3924 (N_3924,N_868,N_724);
and U3925 (N_3925,N_1859,N_1800);
xnor U3926 (N_3926,N_2197,N_67);
or U3927 (N_3927,N_2308,N_2694);
nor U3928 (N_3928,N_1542,N_805);
nor U3929 (N_3929,N_649,N_1115);
or U3930 (N_3930,N_732,N_1752);
nor U3931 (N_3931,N_164,N_752);
nand U3932 (N_3932,N_859,N_1639);
and U3933 (N_3933,N_2239,N_2676);
nor U3934 (N_3934,N_2600,N_20);
or U3935 (N_3935,N_2903,N_2592);
and U3936 (N_3936,N_2253,N_2367);
nand U3937 (N_3937,N_2750,N_2138);
and U3938 (N_3938,N_106,N_1706);
and U3939 (N_3939,N_34,N_2763);
and U3940 (N_3940,N_888,N_490);
nor U3941 (N_3941,N_1537,N_1271);
or U3942 (N_3942,N_255,N_525);
nand U3943 (N_3943,N_2634,N_2618);
nor U3944 (N_3944,N_1842,N_1866);
nor U3945 (N_3945,N_1156,N_1627);
and U3946 (N_3946,N_842,N_2382);
nor U3947 (N_3947,N_2967,N_528);
and U3948 (N_3948,N_2303,N_1152);
nand U3949 (N_3949,N_1297,N_2752);
nor U3950 (N_3950,N_824,N_2174);
or U3951 (N_3951,N_1413,N_459);
nand U3952 (N_3952,N_1357,N_703);
nor U3953 (N_3953,N_189,N_159);
nor U3954 (N_3954,N_1036,N_111);
nand U3955 (N_3955,N_1108,N_2000);
and U3956 (N_3956,N_2976,N_2363);
nor U3957 (N_3957,N_693,N_2359);
or U3958 (N_3958,N_991,N_192);
nor U3959 (N_3959,N_2341,N_945);
or U3960 (N_3960,N_2696,N_1204);
nor U3961 (N_3961,N_1815,N_1070);
or U3962 (N_3962,N_338,N_24);
nand U3963 (N_3963,N_1959,N_1360);
nand U3964 (N_3964,N_2711,N_1226);
nand U3965 (N_3965,N_1870,N_135);
or U3966 (N_3966,N_1533,N_930);
nand U3967 (N_3967,N_985,N_2761);
nor U3968 (N_3968,N_1374,N_630);
or U3969 (N_3969,N_2724,N_1463);
nand U3970 (N_3970,N_2225,N_2765);
nor U3971 (N_3971,N_1914,N_246);
xor U3972 (N_3972,N_566,N_791);
nor U3973 (N_3973,N_604,N_1846);
and U3974 (N_3974,N_2951,N_2668);
nand U3975 (N_3975,N_304,N_1659);
nand U3976 (N_3976,N_2465,N_1117);
and U3977 (N_3977,N_32,N_484);
and U3978 (N_3978,N_1848,N_1657);
and U3979 (N_3979,N_151,N_2843);
nand U3980 (N_3980,N_439,N_61);
or U3981 (N_3981,N_2756,N_2896);
or U3982 (N_3982,N_121,N_804);
nand U3983 (N_3983,N_2847,N_1171);
and U3984 (N_3984,N_2480,N_2964);
nand U3985 (N_3985,N_728,N_427);
or U3986 (N_3986,N_399,N_1388);
nor U3987 (N_3987,N_926,N_2485);
or U3988 (N_3988,N_1393,N_2168);
and U3989 (N_3989,N_1400,N_578);
nor U3990 (N_3990,N_2493,N_2732);
nand U3991 (N_3991,N_2660,N_1287);
nor U3992 (N_3992,N_1694,N_1041);
or U3993 (N_3993,N_2096,N_2723);
and U3994 (N_3994,N_1562,N_2666);
nor U3995 (N_3995,N_1925,N_913);
nor U3996 (N_3996,N_1778,N_2288);
nand U3997 (N_3997,N_2607,N_1203);
or U3998 (N_3998,N_2229,N_1392);
or U3999 (N_3999,N_413,N_278);
nand U4000 (N_4000,N_1061,N_1278);
nand U4001 (N_4001,N_1432,N_2280);
nand U4002 (N_4002,N_1793,N_2796);
and U4003 (N_4003,N_1410,N_782);
or U4004 (N_4004,N_2622,N_2780);
or U4005 (N_4005,N_2977,N_1619);
nor U4006 (N_4006,N_2052,N_1047);
and U4007 (N_4007,N_2867,N_1795);
nor U4008 (N_4008,N_2885,N_2551);
and U4009 (N_4009,N_1140,N_1095);
and U4010 (N_4010,N_1792,N_2862);
and U4011 (N_4011,N_1867,N_2056);
and U4012 (N_4012,N_531,N_2602);
or U4013 (N_4013,N_495,N_2855);
and U4014 (N_4014,N_2494,N_1861);
nand U4015 (N_4015,N_1395,N_1705);
and U4016 (N_4016,N_65,N_553);
and U4017 (N_4017,N_742,N_1625);
nor U4018 (N_4018,N_1212,N_2603);
or U4019 (N_4019,N_1563,N_387);
or U4020 (N_4020,N_1024,N_1241);
and U4021 (N_4021,N_1220,N_765);
or U4022 (N_4022,N_352,N_97);
nor U4023 (N_4023,N_899,N_2669);
nor U4024 (N_4024,N_1352,N_1816);
and U4025 (N_4025,N_1128,N_574);
nor U4026 (N_4026,N_1139,N_284);
nand U4027 (N_4027,N_368,N_2863);
nor U4028 (N_4028,N_1630,N_2975);
nor U4029 (N_4029,N_429,N_2595);
xnor U4030 (N_4030,N_40,N_1088);
nand U4031 (N_4031,N_1048,N_1333);
nor U4032 (N_4032,N_2566,N_1598);
and U4033 (N_4033,N_2537,N_2177);
nand U4034 (N_4034,N_2886,N_785);
nor U4035 (N_4035,N_1568,N_1251);
or U4036 (N_4036,N_1075,N_1853);
nand U4037 (N_4037,N_1764,N_768);
nand U4038 (N_4038,N_2757,N_1862);
nand U4039 (N_4039,N_2032,N_2674);
or U4040 (N_4040,N_1135,N_1594);
nand U4041 (N_4041,N_2983,N_301);
and U4042 (N_4042,N_2203,N_1941);
nor U4043 (N_4043,N_1570,N_2117);
and U4044 (N_4044,N_1147,N_571);
or U4045 (N_4045,N_1864,N_1331);
or U4046 (N_4046,N_1968,N_1300);
and U4047 (N_4047,N_1608,N_1540);
nand U4048 (N_4048,N_898,N_2304);
or U4049 (N_4049,N_2111,N_672);
and U4050 (N_4050,N_1057,N_2671);
and U4051 (N_4051,N_1820,N_1229);
nand U4052 (N_4052,N_1677,N_1691);
or U4053 (N_4053,N_524,N_670);
xnor U4054 (N_4054,N_1797,N_1736);
nand U4055 (N_4055,N_2495,N_2988);
nand U4056 (N_4056,N_1313,N_2463);
and U4057 (N_4057,N_1347,N_745);
and U4058 (N_4058,N_169,N_2083);
nand U4059 (N_4059,N_92,N_2850);
or U4060 (N_4060,N_949,N_175);
or U4061 (N_4061,N_157,N_449);
and U4062 (N_4062,N_2208,N_415);
nand U4063 (N_4063,N_1753,N_1898);
or U4064 (N_4064,N_2309,N_2156);
nand U4065 (N_4065,N_1872,N_535);
and U4066 (N_4066,N_784,N_1601);
nor U4067 (N_4067,N_767,N_2249);
or U4068 (N_4068,N_1210,N_2783);
and U4069 (N_4069,N_2569,N_1995);
nand U4070 (N_4070,N_817,N_983);
or U4071 (N_4071,N_445,N_1638);
nor U4072 (N_4072,N_1766,N_2792);
and U4073 (N_4073,N_1378,N_2183);
or U4074 (N_4074,N_934,N_1326);
or U4075 (N_4075,N_2939,N_2590);
and U4076 (N_4076,N_310,N_1403);
nand U4077 (N_4077,N_998,N_2446);
nor U4078 (N_4078,N_2235,N_530);
or U4079 (N_4079,N_375,N_1161);
or U4080 (N_4080,N_2185,N_2610);
and U4081 (N_4081,N_2258,N_2969);
and U4082 (N_4082,N_1030,N_853);
or U4083 (N_4083,N_512,N_118);
nand U4084 (N_4084,N_2956,N_517);
nor U4085 (N_4085,N_570,N_466);
and U4086 (N_4086,N_2500,N_1206);
nand U4087 (N_4087,N_892,N_902);
and U4088 (N_4088,N_822,N_2003);
or U4089 (N_4089,N_53,N_1248);
xnor U4090 (N_4090,N_2134,N_2015);
xor U4091 (N_4091,N_838,N_2729);
nand U4092 (N_4092,N_683,N_1573);
or U4093 (N_4093,N_579,N_2297);
or U4094 (N_4094,N_2619,N_1018);
nand U4095 (N_4095,N_755,N_264);
nor U4096 (N_4096,N_1196,N_252);
or U4097 (N_4097,N_1183,N_1972);
and U4098 (N_4098,N_138,N_42);
nor U4099 (N_4099,N_1719,N_1411);
or U4100 (N_4100,N_790,N_1453);
nor U4101 (N_4101,N_296,N_1856);
or U4102 (N_4102,N_1512,N_1688);
nor U4103 (N_4103,N_2291,N_1114);
nand U4104 (N_4104,N_816,N_2707);
and U4105 (N_4105,N_1074,N_2274);
nand U4106 (N_4106,N_1649,N_2237);
nand U4107 (N_4107,N_501,N_471);
nor U4108 (N_4108,N_1622,N_1431);
nand U4109 (N_4109,N_1119,N_1079);
and U4110 (N_4110,N_2507,N_2811);
or U4111 (N_4111,N_1607,N_2286);
and U4112 (N_4112,N_1421,N_1510);
or U4113 (N_4113,N_1276,N_2182);
and U4114 (N_4114,N_2207,N_696);
and U4115 (N_4115,N_557,N_140);
and U4116 (N_4116,N_2515,N_1124);
nand U4117 (N_4117,N_889,N_1376);
or U4118 (N_4118,N_2289,N_594);
or U4119 (N_4119,N_2025,N_520);
nor U4120 (N_4120,N_1368,N_2132);
nand U4121 (N_4121,N_1247,N_2377);
nand U4122 (N_4122,N_2784,N_845);
and U4123 (N_4123,N_1494,N_852);
and U4124 (N_4124,N_2631,N_955);
and U4125 (N_4125,N_2758,N_2936);
nand U4126 (N_4126,N_627,N_935);
nand U4127 (N_4127,N_1832,N_751);
or U4128 (N_4128,N_1373,N_2692);
nor U4129 (N_4129,N_608,N_2404);
and U4130 (N_4130,N_758,N_1575);
or U4131 (N_4131,N_1069,N_2257);
or U4132 (N_4132,N_635,N_1632);
nor U4133 (N_4133,N_469,N_1137);
or U4134 (N_4134,N_2586,N_182);
and U4135 (N_4135,N_2907,N_1217);
or U4136 (N_4136,N_2875,N_1022);
nand U4137 (N_4137,N_81,N_2695);
nand U4138 (N_4138,N_1920,N_143);
or U4139 (N_4139,N_1482,N_2380);
and U4140 (N_4140,N_957,N_2655);
nand U4141 (N_4141,N_1684,N_2037);
nand U4142 (N_4142,N_2697,N_2159);
nand U4143 (N_4143,N_458,N_2014);
or U4144 (N_4144,N_2528,N_1102);
nor U4145 (N_4145,N_1587,N_1082);
nor U4146 (N_4146,N_1060,N_1565);
or U4147 (N_4147,N_2370,N_2255);
and U4148 (N_4148,N_1199,N_196);
or U4149 (N_4149,N_2196,N_1133);
nand U4150 (N_4150,N_2094,N_1272);
and U4151 (N_4151,N_2285,N_641);
nor U4152 (N_4152,N_1442,N_108);
or U4153 (N_4153,N_188,N_907);
nor U4154 (N_4154,N_336,N_2432);
and U4155 (N_4155,N_2675,N_2842);
nand U4156 (N_4156,N_2813,N_2008);
or U4157 (N_4157,N_1142,N_45);
or U4158 (N_4158,N_1629,N_2820);
nand U4159 (N_4159,N_1940,N_1812);
and U4160 (N_4160,N_2512,N_2430);
nor U4161 (N_4161,N_1329,N_851);
or U4162 (N_4162,N_411,N_1323);
and U4163 (N_4163,N_194,N_841);
and U4164 (N_4164,N_2467,N_184);
nand U4165 (N_4165,N_837,N_290);
or U4166 (N_4166,N_556,N_2866);
nor U4167 (N_4167,N_1545,N_2293);
and U4168 (N_4168,N_15,N_43);
nor U4169 (N_4169,N_2392,N_1263);
or U4170 (N_4170,N_1144,N_166);
or U4171 (N_4171,N_1484,N_1342);
and U4172 (N_4172,N_1113,N_327);
nand U4173 (N_4173,N_456,N_2663);
nor U4174 (N_4174,N_325,N_1315);
nand U4175 (N_4175,N_401,N_1398);
nand U4176 (N_4176,N_202,N_1216);
nand U4177 (N_4177,N_2415,N_514);
and U4178 (N_4178,N_1680,N_748);
and U4179 (N_4179,N_2301,N_625);
and U4180 (N_4180,N_634,N_628);
and U4181 (N_4181,N_1381,N_1863);
nand U4182 (N_4182,N_2145,N_1973);
nor U4183 (N_4183,N_440,N_876);
or U4184 (N_4184,N_136,N_76);
nor U4185 (N_4185,N_2166,N_506);
or U4186 (N_4186,N_1281,N_323);
nor U4187 (N_4187,N_2471,N_2053);
or U4188 (N_4188,N_493,N_197);
nor U4189 (N_4189,N_1291,N_1092);
nor U4190 (N_4190,N_305,N_2391);
nor U4191 (N_4191,N_1701,N_2069);
and U4192 (N_4192,N_84,N_187);
nor U4193 (N_4193,N_1558,N_2206);
nand U4194 (N_4194,N_2832,N_2556);
nand U4195 (N_4195,N_2305,N_1176);
nand U4196 (N_4196,N_2180,N_2893);
nand U4197 (N_4197,N_1682,N_355);
and U4198 (N_4198,N_2,N_1438);
or U4199 (N_4199,N_2856,N_1197);
and U4200 (N_4200,N_133,N_1123);
nor U4201 (N_4201,N_891,N_2657);
nor U4202 (N_4202,N_1093,N_2444);
and U4203 (N_4203,N_516,N_1817);
nand U4204 (N_4204,N_1285,N_2985);
nor U4205 (N_4205,N_1544,N_1900);
or U4206 (N_4206,N_2741,N_2508);
or U4207 (N_4207,N_1160,N_2299);
nand U4208 (N_4208,N_779,N_397);
or U4209 (N_4209,N_1843,N_2548);
xnor U4210 (N_4210,N_2332,N_2242);
and U4211 (N_4211,N_2629,N_99);
nor U4212 (N_4212,N_2648,N_266);
nor U4213 (N_4213,N_315,N_87);
or U4214 (N_4214,N_1185,N_2442);
nand U4215 (N_4215,N_2909,N_287);
nor U4216 (N_4216,N_878,N_1606);
nor U4217 (N_4217,N_1678,N_1801);
and U4218 (N_4218,N_781,N_915);
nand U4219 (N_4219,N_1211,N_2864);
nand U4220 (N_4220,N_1865,N_409);
nor U4221 (N_4221,N_857,N_607);
or U4222 (N_4222,N_966,N_807);
and U4223 (N_4223,N_137,N_2058);
nand U4224 (N_4224,N_321,N_858);
and U4225 (N_4225,N_179,N_617);
nor U4226 (N_4226,N_2459,N_646);
and U4227 (N_4227,N_1169,N_1946);
and U4228 (N_4228,N_1265,N_972);
nor U4229 (N_4229,N_2865,N_353);
nor U4230 (N_4230,N_2345,N_1727);
nor U4231 (N_4231,N_2018,N_2104);
or U4232 (N_4232,N_365,N_1447);
and U4233 (N_4233,N_2070,N_351);
nor U4234 (N_4234,N_1523,N_2327);
nand U4235 (N_4235,N_2987,N_932);
or U4236 (N_4236,N_1609,N_1382);
or U4237 (N_4237,N_2749,N_575);
nand U4238 (N_4238,N_869,N_1529);
nor U4239 (N_4239,N_347,N_680);
nor U4240 (N_4240,N_481,N_924);
nand U4241 (N_4241,N_1654,N_2944);
xnor U4242 (N_4242,N_772,N_26);
and U4243 (N_4243,N_2786,N_1751);
nand U4244 (N_4244,N_1489,N_2940);
and U4245 (N_4245,N_1448,N_2771);
nand U4246 (N_4246,N_134,N_1003);
nand U4247 (N_4247,N_2411,N_1044);
xnor U4248 (N_4248,N_2795,N_1063);
nor U4249 (N_4249,N_378,N_362);
and U4250 (N_4250,N_2646,N_2406);
and U4251 (N_4251,N_2445,N_237);
nand U4252 (N_4252,N_717,N_314);
nand U4253 (N_4253,N_1172,N_1841);
or U4254 (N_4254,N_2898,N_1615);
and U4255 (N_4255,N_479,N_1879);
nand U4256 (N_4256,N_292,N_2023);
and U4257 (N_4257,N_1110,N_10);
nor U4258 (N_4258,N_1883,N_1744);
or U4259 (N_4259,N_497,N_2994);
nor U4260 (N_4260,N_1634,N_1042);
nor U4261 (N_4261,N_2530,N_2638);
and U4262 (N_4262,N_2097,N_642);
nand U4263 (N_4263,N_2501,N_1289);
or U4264 (N_4264,N_113,N_408);
nor U4265 (N_4265,N_1288,N_2362);
or U4266 (N_4266,N_1445,N_536);
nand U4267 (N_4267,N_1019,N_632);
nand U4268 (N_4268,N_1243,N_2142);
nor U4269 (N_4269,N_614,N_1624);
and U4270 (N_4270,N_1132,N_332);
or U4271 (N_4271,N_2819,N_893);
nor U4272 (N_4272,N_2952,N_2116);
nor U4273 (N_4273,N_1505,N_2702);
or U4274 (N_4274,N_1926,N_1664);
nand U4275 (N_4275,N_2306,N_1667);
nor U4276 (N_4276,N_1527,N_308);
or U4277 (N_4277,N_2974,N_616);
nor U4278 (N_4278,N_770,N_2623);
nand U4279 (N_4279,N_1213,N_56);
nor U4280 (N_4280,N_2374,N_158);
and U4281 (N_4281,N_2510,N_846);
nor U4282 (N_4282,N_2930,N_929);
and U4283 (N_4283,N_1404,N_1702);
or U4284 (N_4284,N_866,N_1571);
nor U4285 (N_4285,N_836,N_2338);
nor U4286 (N_4286,N_2680,N_1643);
nor U4287 (N_4287,N_2662,N_997);
and U4288 (N_4288,N_2549,N_2150);
and U4289 (N_4289,N_1125,N_1454);
nor U4290 (N_4290,N_70,N_2836);
nand U4291 (N_4291,N_2751,N_218);
or U4292 (N_4292,N_489,N_1105);
nand U4293 (N_4293,N_1519,N_1576);
and U4294 (N_4294,N_1947,N_1618);
nor U4295 (N_4295,N_1796,N_1583);
and U4296 (N_4296,N_2137,N_1836);
or U4297 (N_4297,N_2407,N_1192);
xnor U4298 (N_4298,N_2292,N_977);
or U4299 (N_4299,N_227,N_940);
nor U4300 (N_4300,N_2336,N_1683);
nand U4301 (N_4301,N_2076,N_2100);
and U4302 (N_4302,N_2691,N_1254);
nor U4303 (N_4303,N_519,N_1924);
nand U4304 (N_4304,N_2329,N_82);
and U4305 (N_4305,N_933,N_1426);
nor U4306 (N_4306,N_2167,N_1245);
and U4307 (N_4307,N_875,N_1936);
and U4308 (N_4308,N_337,N_812);
and U4309 (N_4309,N_1066,N_2160);
nand U4310 (N_4310,N_2762,N_2443);
or U4311 (N_4311,N_2201,N_870);
and U4312 (N_4312,N_2381,N_1262);
nand U4313 (N_4313,N_232,N_2861);
or U4314 (N_4314,N_2546,N_2978);
nor U4315 (N_4315,N_215,N_1965);
nand U4316 (N_4316,N_725,N_737);
nor U4317 (N_4317,N_1887,N_1283);
and U4318 (N_4318,N_251,N_130);
or U4319 (N_4319,N_1077,N_2175);
nor U4320 (N_4320,N_1073,N_2190);
nor U4321 (N_4321,N_559,N_2220);
and U4322 (N_4322,N_2645,N_2426);
nand U4323 (N_4323,N_2719,N_1072);
nand U4324 (N_4324,N_1916,N_203);
nand U4325 (N_4325,N_1839,N_240);
nor U4326 (N_4326,N_2506,N_1004);
and U4327 (N_4327,N_2760,N_2366);
nor U4328 (N_4328,N_2541,N_2393);
or U4329 (N_4329,N_759,N_2216);
or U4330 (N_4330,N_2405,N_989);
nor U4331 (N_4331,N_2039,N_979);
and U4332 (N_4332,N_825,N_334);
and U4333 (N_4333,N_2849,N_2433);
or U4334 (N_4334,N_2575,N_1559);
nor U4335 (N_4335,N_1273,N_620);
or U4336 (N_4336,N_2101,N_2176);
nor U4337 (N_4337,N_2703,N_673);
and U4338 (N_4338,N_1111,N_270);
or U4339 (N_4339,N_2564,N_2351);
nor U4340 (N_4340,N_1532,N_2665);
or U4341 (N_4341,N_963,N_552);
or U4342 (N_4342,N_2576,N_1201);
and U4343 (N_4343,N_647,N_2503);
nand U4344 (N_4344,N_1399,N_2387);
or U4345 (N_4345,N_2460,N_1547);
or U4346 (N_4346,N_455,N_1656);
and U4347 (N_4347,N_1040,N_2213);
and U4348 (N_4348,N_2126,N_83);
and U4349 (N_4349,N_2450,N_380);
nand U4350 (N_4350,N_951,N_2681);
nor U4351 (N_4351,N_832,N_2989);
nand U4352 (N_4352,N_1912,N_914);
or U4353 (N_4353,N_1991,N_2340);
nand U4354 (N_4354,N_1960,N_2841);
or U4355 (N_4355,N_2133,N_690);
nand U4356 (N_4356,N_1951,N_2087);
and U4357 (N_4357,N_537,N_2598);
and U4358 (N_4358,N_1652,N_2517);
nand U4359 (N_4359,N_2482,N_1407);
and U4360 (N_4360,N_1219,N_839);
and U4361 (N_4361,N_835,N_1299);
and U4362 (N_4362,N_1834,N_317);
and U4363 (N_4363,N_122,N_708);
or U4364 (N_4364,N_860,N_795);
or U4365 (N_4365,N_2331,N_2767);
and U4366 (N_4366,N_1845,N_1577);
nand U4367 (N_4367,N_163,N_51);
and U4368 (N_4368,N_1828,N_2686);
and U4369 (N_4369,N_2136,N_2186);
nand U4370 (N_4370,N_1363,N_2173);
or U4371 (N_4371,N_131,N_1873);
and U4372 (N_4372,N_874,N_2915);
and U4373 (N_4373,N_95,N_1591);
and U4374 (N_4374,N_1234,N_1785);
nor U4375 (N_4375,N_2356,N_1301);
nand U4376 (N_4376,N_419,N_1379);
nor U4377 (N_4377,N_2873,N_285);
nand U4378 (N_4378,N_1788,N_1026);
nor U4379 (N_4379,N_2606,N_1781);
nand U4380 (N_4380,N_295,N_953);
and U4381 (N_4381,N_1646,N_820);
nor U4382 (N_4382,N_801,N_1698);
nor U4383 (N_4383,N_483,N_631);
or U4384 (N_4384,N_2845,N_1905);
or U4385 (N_4385,N_2844,N_2877);
nor U4386 (N_4386,N_2221,N_2310);
nor U4387 (N_4387,N_1642,N_1052);
nor U4388 (N_4388,N_1011,N_2880);
and U4389 (N_4389,N_422,N_1007);
nand U4390 (N_4390,N_750,N_78);
nand U4391 (N_4391,N_2313,N_746);
nor U4392 (N_4392,N_1998,N_965);
nand U4393 (N_4393,N_2389,N_1031);
and U4394 (N_4394,N_2775,N_2343);
nor U4395 (N_4395,N_561,N_2932);
and U4396 (N_4396,N_2846,N_110);
nand U4397 (N_4397,N_2704,N_885);
or U4398 (N_4398,N_2455,N_1561);
nand U4399 (N_4399,N_2139,N_2986);
nand U4400 (N_4400,N_2822,N_1322);
or U4401 (N_4401,N_462,N_1886);
nand U4402 (N_4402,N_546,N_2119);
and U4403 (N_4403,N_47,N_398);
or U4404 (N_4404,N_2294,N_1763);
and U4405 (N_4405,N_2202,N_2892);
nor U4406 (N_4406,N_2211,N_754);
and U4407 (N_4407,N_267,N_1502);
and U4408 (N_4408,N_1230,N_1306);
and U4409 (N_4409,N_1851,N_733);
nand U4410 (N_4410,N_2403,N_911);
nor U4411 (N_4411,N_457,N_1330);
nand U4412 (N_4412,N_1345,N_2198);
and U4413 (N_4413,N_1955,N_1881);
nor U4414 (N_4414,N_2923,N_1874);
or U4415 (N_4415,N_2879,N_756);
and U4416 (N_4416,N_762,N_1434);
or U4417 (N_4417,N_2109,N_521);
nand U4418 (N_4418,N_430,N_723);
or U4419 (N_4419,N_1858,N_2273);
and U4420 (N_4420,N_1064,N_650);
nand U4421 (N_4421,N_2040,N_286);
or U4422 (N_4422,N_906,N_344);
or U4423 (N_4423,N_2884,N_376);
nand U4424 (N_4424,N_2812,N_2523);
and U4425 (N_4425,N_2265,N_1930);
nor U4426 (N_4426,N_2398,N_2605);
nor U4427 (N_4427,N_1149,N_2661);
and U4428 (N_4428,N_2826,N_2851);
nand U4429 (N_4429,N_964,N_657);
and U4430 (N_4430,N_505,N_1205);
nor U4431 (N_4431,N_2937,N_2924);
and U4432 (N_4432,N_522,N_2860);
nor U4433 (N_4433,N_1369,N_291);
nand U4434 (N_4434,N_1600,N_948);
xor U4435 (N_4435,N_818,N_2800);
and U4436 (N_4436,N_555,N_2005);
nor U4437 (N_4437,N_1687,N_2524);
nor U4438 (N_4438,N_109,N_2088);
or U4439 (N_4439,N_1720,N_1488);
nand U4440 (N_4440,N_597,N_1878);
and U4441 (N_4441,N_2244,N_1);
nand U4442 (N_4442,N_2034,N_668);
nand U4443 (N_4443,N_1938,N_1343);
nor U4444 (N_4444,N_549,N_1888);
nor U4445 (N_4445,N_1913,N_664);
nor U4446 (N_4446,N_104,N_1999);
nand U4447 (N_4447,N_2112,N_962);
nand U4448 (N_4448,N_1444,N_564);
nand U4449 (N_4449,N_2960,N_441);
or U4450 (N_4450,N_1942,N_806);
or U4451 (N_4451,N_253,N_231);
and U4452 (N_4452,N_186,N_333);
nand U4453 (N_4453,N_2422,N_433);
nor U4454 (N_4454,N_2427,N_1223);
or U4455 (N_4455,N_2408,N_2848);
or U4456 (N_4456,N_366,N_464);
nand U4457 (N_4457,N_2774,N_2790);
or U4458 (N_4458,N_1578,N_2794);
and U4459 (N_4459,N_1644,N_328);
nand U4460 (N_4460,N_461,N_2461);
and U4461 (N_4461,N_191,N_2970);
and U4462 (N_4462,N_343,N_2876);
and U4463 (N_4463,N_2140,N_349);
nand U4464 (N_4464,N_1983,N_601);
and U4465 (N_4465,N_2962,N_2298);
and U4466 (N_4466,N_1462,N_2938);
nand U4467 (N_4467,N_1406,N_2581);
nand U4468 (N_4468,N_1116,N_482);
and U4469 (N_4469,N_2688,N_2371);
nand U4470 (N_4470,N_1280,N_1809);
nor U4471 (N_4471,N_510,N_1595);
nor U4472 (N_4472,N_1005,N_393);
nand U4473 (N_4473,N_1903,N_486);
nor U4474 (N_4474,N_677,N_1655);
and U4475 (N_4475,N_1536,N_919);
and U4476 (N_4476,N_2709,N_2385);
nor U4477 (N_4477,N_1782,N_1923);
nand U4478 (N_4478,N_1696,N_281);
and U4479 (N_4479,N_1765,N_2561);
and U4480 (N_4480,N_1885,N_897);
or U4481 (N_4481,N_928,N_711);
nand U4482 (N_4482,N_2234,N_280);
and U4483 (N_4483,N_2531,N_916);
nor U4484 (N_4484,N_2369,N_1827);
and U4485 (N_4485,N_1964,N_1175);
nor U4486 (N_4486,N_973,N_609);
and U4487 (N_4487,N_1261,N_2231);
or U4488 (N_4488,N_173,N_406);
xor U4489 (N_4489,N_749,N_1355);
nand U4490 (N_4490,N_2110,N_2642);
nand U4491 (N_4491,N_1740,N_2881);
nand U4492 (N_4492,N_1043,N_1722);
nand U4493 (N_4493,N_633,N_1181);
nor U4494 (N_4494,N_2714,N_704);
and U4495 (N_4495,N_652,N_1490);
nor U4496 (N_4496,N_1725,N_2838);
and U4497 (N_4497,N_2961,N_2870);
and U4498 (N_4498,N_2816,N_261);
and U4499 (N_4499,N_598,N_363);
or U4500 (N_4500,N_69,N_1476);
nand U4501 (N_4501,N_2809,N_592);
nor U4502 (N_4502,N_750,N_1550);
nand U4503 (N_4503,N_237,N_2374);
and U4504 (N_4504,N_1201,N_1149);
or U4505 (N_4505,N_2715,N_353);
nor U4506 (N_4506,N_965,N_451);
nand U4507 (N_4507,N_520,N_2802);
nand U4508 (N_4508,N_542,N_891);
and U4509 (N_4509,N_470,N_113);
or U4510 (N_4510,N_2486,N_2227);
and U4511 (N_4511,N_2278,N_909);
and U4512 (N_4512,N_2285,N_2595);
nand U4513 (N_4513,N_1621,N_858);
nand U4514 (N_4514,N_2645,N_149);
or U4515 (N_4515,N_2804,N_1705);
and U4516 (N_4516,N_307,N_2226);
and U4517 (N_4517,N_2788,N_1508);
nor U4518 (N_4518,N_2744,N_186);
and U4519 (N_4519,N_1814,N_2558);
nor U4520 (N_4520,N_2754,N_2374);
nand U4521 (N_4521,N_784,N_1024);
or U4522 (N_4522,N_2359,N_2170);
or U4523 (N_4523,N_2806,N_608);
nand U4524 (N_4524,N_92,N_191);
or U4525 (N_4525,N_276,N_821);
and U4526 (N_4526,N_481,N_426);
nor U4527 (N_4527,N_1488,N_811);
nand U4528 (N_4528,N_1842,N_857);
and U4529 (N_4529,N_1797,N_2042);
and U4530 (N_4530,N_777,N_2468);
or U4531 (N_4531,N_36,N_774);
and U4532 (N_4532,N_1038,N_2949);
or U4533 (N_4533,N_1309,N_15);
and U4534 (N_4534,N_808,N_2959);
nor U4535 (N_4535,N_1764,N_1245);
and U4536 (N_4536,N_1719,N_1747);
nand U4537 (N_4537,N_339,N_115);
and U4538 (N_4538,N_2774,N_593);
nand U4539 (N_4539,N_33,N_809);
or U4540 (N_4540,N_1709,N_1341);
nand U4541 (N_4541,N_1646,N_72);
or U4542 (N_4542,N_624,N_2864);
and U4543 (N_4543,N_2807,N_2101);
xnor U4544 (N_4544,N_2616,N_1540);
and U4545 (N_4545,N_2093,N_1942);
nand U4546 (N_4546,N_523,N_1232);
nand U4547 (N_4547,N_732,N_2914);
or U4548 (N_4548,N_341,N_955);
and U4549 (N_4549,N_43,N_579);
and U4550 (N_4550,N_355,N_2184);
and U4551 (N_4551,N_913,N_2592);
nand U4552 (N_4552,N_136,N_1655);
or U4553 (N_4553,N_1360,N_1925);
or U4554 (N_4554,N_2855,N_1025);
or U4555 (N_4555,N_1571,N_1053);
nor U4556 (N_4556,N_2635,N_186);
nand U4557 (N_4557,N_159,N_2562);
or U4558 (N_4558,N_2883,N_1381);
nor U4559 (N_4559,N_1364,N_2654);
nand U4560 (N_4560,N_2586,N_363);
and U4561 (N_4561,N_1263,N_2756);
or U4562 (N_4562,N_2669,N_2884);
nand U4563 (N_4563,N_1310,N_2953);
nand U4564 (N_4564,N_669,N_182);
nand U4565 (N_4565,N_856,N_845);
and U4566 (N_4566,N_1602,N_2243);
and U4567 (N_4567,N_2483,N_2177);
and U4568 (N_4568,N_1471,N_1489);
or U4569 (N_4569,N_534,N_2967);
or U4570 (N_4570,N_1184,N_12);
nand U4571 (N_4571,N_1517,N_1071);
and U4572 (N_4572,N_2180,N_2949);
nand U4573 (N_4573,N_2309,N_2216);
nand U4574 (N_4574,N_2012,N_325);
and U4575 (N_4575,N_410,N_2691);
nand U4576 (N_4576,N_624,N_332);
and U4577 (N_4577,N_247,N_1958);
nor U4578 (N_4578,N_1674,N_851);
nor U4579 (N_4579,N_2969,N_869);
or U4580 (N_4580,N_2563,N_1201);
nor U4581 (N_4581,N_2445,N_2006);
nor U4582 (N_4582,N_1504,N_1500);
or U4583 (N_4583,N_1143,N_1676);
nor U4584 (N_4584,N_1781,N_1460);
nor U4585 (N_4585,N_1610,N_505);
nand U4586 (N_4586,N_1416,N_872);
or U4587 (N_4587,N_1898,N_2356);
or U4588 (N_4588,N_1741,N_842);
nand U4589 (N_4589,N_1984,N_949);
and U4590 (N_4590,N_2600,N_1266);
nand U4591 (N_4591,N_870,N_679);
or U4592 (N_4592,N_2192,N_2526);
nand U4593 (N_4593,N_2391,N_684);
nand U4594 (N_4594,N_189,N_2725);
or U4595 (N_4595,N_1231,N_2515);
or U4596 (N_4596,N_1507,N_469);
nand U4597 (N_4597,N_2717,N_2174);
or U4598 (N_4598,N_2465,N_1224);
or U4599 (N_4599,N_436,N_2186);
or U4600 (N_4600,N_2603,N_1928);
nor U4601 (N_4601,N_524,N_1084);
or U4602 (N_4602,N_2537,N_2606);
xor U4603 (N_4603,N_2978,N_2352);
or U4604 (N_4604,N_1288,N_1374);
nor U4605 (N_4605,N_1741,N_2744);
or U4606 (N_4606,N_2668,N_541);
nand U4607 (N_4607,N_1276,N_519);
nor U4608 (N_4608,N_1559,N_2813);
nor U4609 (N_4609,N_94,N_2155);
or U4610 (N_4610,N_2937,N_1702);
nand U4611 (N_4611,N_338,N_2223);
nand U4612 (N_4612,N_644,N_2618);
and U4613 (N_4613,N_1304,N_14);
nand U4614 (N_4614,N_1536,N_1679);
and U4615 (N_4615,N_301,N_2851);
nand U4616 (N_4616,N_2680,N_2342);
and U4617 (N_4617,N_228,N_370);
or U4618 (N_4618,N_198,N_432);
nand U4619 (N_4619,N_1358,N_149);
or U4620 (N_4620,N_2742,N_883);
or U4621 (N_4621,N_1253,N_2522);
or U4622 (N_4622,N_2339,N_251);
nor U4623 (N_4623,N_1973,N_1819);
and U4624 (N_4624,N_1909,N_149);
and U4625 (N_4625,N_339,N_2282);
and U4626 (N_4626,N_2911,N_195);
nor U4627 (N_4627,N_1923,N_2108);
and U4628 (N_4628,N_2582,N_1894);
or U4629 (N_4629,N_2466,N_2638);
nor U4630 (N_4630,N_1343,N_2642);
nor U4631 (N_4631,N_1474,N_1126);
nor U4632 (N_4632,N_2179,N_737);
or U4633 (N_4633,N_2540,N_2040);
or U4634 (N_4634,N_303,N_2726);
nor U4635 (N_4635,N_429,N_2235);
nor U4636 (N_4636,N_93,N_1252);
nor U4637 (N_4637,N_2133,N_1216);
nand U4638 (N_4638,N_722,N_666);
nor U4639 (N_4639,N_858,N_810);
xnor U4640 (N_4640,N_2908,N_2752);
or U4641 (N_4641,N_2536,N_1431);
nor U4642 (N_4642,N_1818,N_1664);
nor U4643 (N_4643,N_325,N_1567);
nand U4644 (N_4644,N_943,N_1463);
and U4645 (N_4645,N_2648,N_634);
and U4646 (N_4646,N_2521,N_2805);
nor U4647 (N_4647,N_1578,N_861);
nor U4648 (N_4648,N_2513,N_1023);
or U4649 (N_4649,N_900,N_810);
nand U4650 (N_4650,N_123,N_125);
or U4651 (N_4651,N_69,N_294);
nor U4652 (N_4652,N_1029,N_2257);
or U4653 (N_4653,N_706,N_1900);
nor U4654 (N_4654,N_325,N_2574);
nor U4655 (N_4655,N_1839,N_2828);
xor U4656 (N_4656,N_842,N_1364);
nor U4657 (N_4657,N_869,N_2034);
nor U4658 (N_4658,N_1303,N_1419);
nor U4659 (N_4659,N_25,N_1106);
nand U4660 (N_4660,N_51,N_432);
and U4661 (N_4661,N_908,N_159);
and U4662 (N_4662,N_1124,N_2752);
nor U4663 (N_4663,N_145,N_2028);
or U4664 (N_4664,N_1417,N_2455);
or U4665 (N_4665,N_859,N_54);
or U4666 (N_4666,N_252,N_936);
nand U4667 (N_4667,N_168,N_537);
nor U4668 (N_4668,N_2527,N_1729);
and U4669 (N_4669,N_1338,N_1107);
or U4670 (N_4670,N_2071,N_1181);
or U4671 (N_4671,N_1264,N_622);
nand U4672 (N_4672,N_1786,N_1258);
or U4673 (N_4673,N_364,N_419);
nand U4674 (N_4674,N_379,N_1074);
and U4675 (N_4675,N_1808,N_2084);
nand U4676 (N_4676,N_1617,N_1840);
nand U4677 (N_4677,N_282,N_2749);
nor U4678 (N_4678,N_1605,N_1860);
or U4679 (N_4679,N_2920,N_2044);
nor U4680 (N_4680,N_123,N_1149);
and U4681 (N_4681,N_2397,N_2650);
nand U4682 (N_4682,N_2304,N_1261);
nor U4683 (N_4683,N_324,N_2346);
and U4684 (N_4684,N_1443,N_1650);
or U4685 (N_4685,N_2042,N_2926);
and U4686 (N_4686,N_2008,N_1463);
nor U4687 (N_4687,N_623,N_2444);
or U4688 (N_4688,N_1757,N_2599);
and U4689 (N_4689,N_1301,N_660);
or U4690 (N_4690,N_1202,N_2084);
nor U4691 (N_4691,N_1172,N_1245);
nand U4692 (N_4692,N_2457,N_1230);
nor U4693 (N_4693,N_2885,N_1463);
and U4694 (N_4694,N_22,N_2092);
or U4695 (N_4695,N_784,N_538);
nor U4696 (N_4696,N_1102,N_462);
and U4697 (N_4697,N_2624,N_2194);
and U4698 (N_4698,N_2672,N_317);
nand U4699 (N_4699,N_2213,N_248);
or U4700 (N_4700,N_2740,N_861);
and U4701 (N_4701,N_443,N_1128);
nand U4702 (N_4702,N_1710,N_2655);
nor U4703 (N_4703,N_950,N_1509);
nor U4704 (N_4704,N_2121,N_2941);
and U4705 (N_4705,N_2117,N_54);
or U4706 (N_4706,N_1731,N_804);
and U4707 (N_4707,N_1182,N_1604);
and U4708 (N_4708,N_2515,N_1876);
or U4709 (N_4709,N_1796,N_29);
and U4710 (N_4710,N_2814,N_1452);
nand U4711 (N_4711,N_293,N_2855);
nand U4712 (N_4712,N_2431,N_1167);
and U4713 (N_4713,N_826,N_1356);
nand U4714 (N_4714,N_2080,N_1362);
or U4715 (N_4715,N_2484,N_216);
and U4716 (N_4716,N_45,N_1760);
nand U4717 (N_4717,N_622,N_1514);
or U4718 (N_4718,N_354,N_2921);
or U4719 (N_4719,N_1455,N_2036);
nand U4720 (N_4720,N_605,N_2185);
or U4721 (N_4721,N_1013,N_295);
and U4722 (N_4722,N_2630,N_2254);
nor U4723 (N_4723,N_1721,N_81);
nor U4724 (N_4724,N_399,N_310);
or U4725 (N_4725,N_557,N_164);
and U4726 (N_4726,N_1396,N_866);
and U4727 (N_4727,N_2145,N_1031);
and U4728 (N_4728,N_2017,N_1050);
or U4729 (N_4729,N_2632,N_1303);
nand U4730 (N_4730,N_2325,N_168);
and U4731 (N_4731,N_1760,N_1677);
and U4732 (N_4732,N_2269,N_1137);
and U4733 (N_4733,N_1844,N_518);
or U4734 (N_4734,N_235,N_2201);
nand U4735 (N_4735,N_1748,N_261);
nor U4736 (N_4736,N_2090,N_1361);
or U4737 (N_4737,N_1053,N_2372);
or U4738 (N_4738,N_2947,N_2701);
nand U4739 (N_4739,N_1500,N_1912);
or U4740 (N_4740,N_1592,N_1122);
or U4741 (N_4741,N_10,N_1584);
nor U4742 (N_4742,N_1278,N_2518);
nor U4743 (N_4743,N_2402,N_2285);
nand U4744 (N_4744,N_2326,N_2324);
or U4745 (N_4745,N_285,N_2479);
and U4746 (N_4746,N_2243,N_596);
xor U4747 (N_4747,N_934,N_457);
nand U4748 (N_4748,N_1067,N_1655);
nand U4749 (N_4749,N_1457,N_1300);
or U4750 (N_4750,N_1915,N_776);
nand U4751 (N_4751,N_1647,N_721);
or U4752 (N_4752,N_606,N_194);
nor U4753 (N_4753,N_1263,N_805);
and U4754 (N_4754,N_1299,N_1730);
nand U4755 (N_4755,N_1709,N_1435);
nand U4756 (N_4756,N_1483,N_2554);
nor U4757 (N_4757,N_1956,N_1399);
nor U4758 (N_4758,N_396,N_1644);
nor U4759 (N_4759,N_2304,N_1189);
nand U4760 (N_4760,N_2550,N_296);
nor U4761 (N_4761,N_2274,N_46);
and U4762 (N_4762,N_2123,N_1293);
nand U4763 (N_4763,N_238,N_724);
nand U4764 (N_4764,N_2715,N_901);
and U4765 (N_4765,N_1377,N_2386);
or U4766 (N_4766,N_67,N_1500);
or U4767 (N_4767,N_1482,N_167);
and U4768 (N_4768,N_2101,N_1850);
or U4769 (N_4769,N_449,N_247);
nand U4770 (N_4770,N_1387,N_1812);
or U4771 (N_4771,N_1404,N_1598);
or U4772 (N_4772,N_1376,N_1953);
and U4773 (N_4773,N_632,N_2236);
and U4774 (N_4774,N_360,N_1260);
nor U4775 (N_4775,N_1276,N_1731);
nand U4776 (N_4776,N_2830,N_1695);
nand U4777 (N_4777,N_2537,N_1897);
or U4778 (N_4778,N_342,N_2491);
and U4779 (N_4779,N_521,N_2605);
nand U4780 (N_4780,N_207,N_1677);
nor U4781 (N_4781,N_1766,N_1808);
and U4782 (N_4782,N_2781,N_2795);
nor U4783 (N_4783,N_1328,N_132);
nand U4784 (N_4784,N_2098,N_2599);
and U4785 (N_4785,N_2496,N_2755);
or U4786 (N_4786,N_2877,N_2773);
nand U4787 (N_4787,N_773,N_164);
or U4788 (N_4788,N_1321,N_1181);
nor U4789 (N_4789,N_653,N_2104);
nand U4790 (N_4790,N_1374,N_1868);
xnor U4791 (N_4791,N_445,N_2615);
or U4792 (N_4792,N_1857,N_2798);
or U4793 (N_4793,N_1578,N_1994);
and U4794 (N_4794,N_262,N_1411);
nand U4795 (N_4795,N_1242,N_2826);
and U4796 (N_4796,N_1319,N_1951);
and U4797 (N_4797,N_588,N_1532);
or U4798 (N_4798,N_1932,N_2204);
or U4799 (N_4799,N_2598,N_731);
or U4800 (N_4800,N_2873,N_296);
nand U4801 (N_4801,N_2080,N_2883);
and U4802 (N_4802,N_178,N_837);
or U4803 (N_4803,N_2616,N_1255);
nor U4804 (N_4804,N_2671,N_818);
nor U4805 (N_4805,N_1053,N_263);
or U4806 (N_4806,N_2138,N_2080);
nand U4807 (N_4807,N_2489,N_1523);
nor U4808 (N_4808,N_2229,N_879);
or U4809 (N_4809,N_1631,N_2673);
and U4810 (N_4810,N_2843,N_1314);
or U4811 (N_4811,N_1151,N_1166);
nor U4812 (N_4812,N_870,N_402);
and U4813 (N_4813,N_385,N_2790);
and U4814 (N_4814,N_2699,N_2818);
nand U4815 (N_4815,N_548,N_2580);
and U4816 (N_4816,N_1417,N_1413);
or U4817 (N_4817,N_2647,N_1205);
and U4818 (N_4818,N_2694,N_1114);
nor U4819 (N_4819,N_701,N_129);
nand U4820 (N_4820,N_322,N_313);
nor U4821 (N_4821,N_2169,N_1248);
or U4822 (N_4822,N_2311,N_2100);
nor U4823 (N_4823,N_1151,N_109);
or U4824 (N_4824,N_447,N_824);
or U4825 (N_4825,N_1935,N_697);
or U4826 (N_4826,N_233,N_1208);
nor U4827 (N_4827,N_2193,N_945);
or U4828 (N_4828,N_2384,N_649);
nor U4829 (N_4829,N_1008,N_1012);
or U4830 (N_4830,N_1385,N_768);
nor U4831 (N_4831,N_1889,N_2969);
nor U4832 (N_4832,N_2727,N_2443);
and U4833 (N_4833,N_399,N_2688);
nand U4834 (N_4834,N_745,N_2495);
and U4835 (N_4835,N_697,N_2637);
nand U4836 (N_4836,N_859,N_866);
or U4837 (N_4837,N_2034,N_762);
xor U4838 (N_4838,N_2567,N_2876);
or U4839 (N_4839,N_2180,N_1970);
and U4840 (N_4840,N_2358,N_1326);
and U4841 (N_4841,N_1570,N_2874);
and U4842 (N_4842,N_138,N_237);
and U4843 (N_4843,N_1125,N_2383);
nor U4844 (N_4844,N_2582,N_2473);
nor U4845 (N_4845,N_849,N_2150);
nor U4846 (N_4846,N_2238,N_191);
or U4847 (N_4847,N_1230,N_1108);
and U4848 (N_4848,N_2130,N_2864);
or U4849 (N_4849,N_1837,N_32);
or U4850 (N_4850,N_1022,N_476);
nand U4851 (N_4851,N_1394,N_561);
or U4852 (N_4852,N_115,N_975);
and U4853 (N_4853,N_1688,N_109);
and U4854 (N_4854,N_2272,N_1184);
nor U4855 (N_4855,N_1284,N_1364);
nand U4856 (N_4856,N_1138,N_313);
nand U4857 (N_4857,N_2796,N_100);
and U4858 (N_4858,N_849,N_1091);
nand U4859 (N_4859,N_1293,N_952);
or U4860 (N_4860,N_372,N_1808);
xor U4861 (N_4861,N_1345,N_987);
nor U4862 (N_4862,N_1551,N_1123);
nand U4863 (N_4863,N_661,N_1791);
nor U4864 (N_4864,N_1353,N_995);
and U4865 (N_4865,N_1663,N_950);
and U4866 (N_4866,N_2381,N_2583);
or U4867 (N_4867,N_807,N_520);
or U4868 (N_4868,N_516,N_2608);
or U4869 (N_4869,N_1484,N_1288);
nand U4870 (N_4870,N_1578,N_2802);
and U4871 (N_4871,N_2053,N_2640);
and U4872 (N_4872,N_2646,N_284);
or U4873 (N_4873,N_578,N_1655);
nand U4874 (N_4874,N_1827,N_1120);
nand U4875 (N_4875,N_1095,N_2766);
nor U4876 (N_4876,N_281,N_1905);
or U4877 (N_4877,N_762,N_1288);
nor U4878 (N_4878,N_1741,N_1029);
nor U4879 (N_4879,N_1745,N_1734);
and U4880 (N_4880,N_324,N_2482);
nor U4881 (N_4881,N_1930,N_1397);
or U4882 (N_4882,N_2602,N_982);
and U4883 (N_4883,N_1882,N_2034);
or U4884 (N_4884,N_2887,N_2501);
nor U4885 (N_4885,N_1925,N_2051);
nand U4886 (N_4886,N_1324,N_2799);
and U4887 (N_4887,N_2085,N_2422);
nand U4888 (N_4888,N_138,N_27);
and U4889 (N_4889,N_1175,N_105);
and U4890 (N_4890,N_974,N_852);
nand U4891 (N_4891,N_48,N_544);
or U4892 (N_4892,N_2833,N_334);
nor U4893 (N_4893,N_553,N_982);
nor U4894 (N_4894,N_282,N_295);
nor U4895 (N_4895,N_445,N_1759);
or U4896 (N_4896,N_2423,N_2368);
and U4897 (N_4897,N_2403,N_781);
nor U4898 (N_4898,N_2298,N_1036);
or U4899 (N_4899,N_2225,N_1448);
and U4900 (N_4900,N_2718,N_2420);
nand U4901 (N_4901,N_788,N_2216);
and U4902 (N_4902,N_696,N_2551);
or U4903 (N_4903,N_2810,N_407);
and U4904 (N_4904,N_683,N_313);
and U4905 (N_4905,N_432,N_2903);
nor U4906 (N_4906,N_1441,N_2602);
nand U4907 (N_4907,N_2,N_428);
nor U4908 (N_4908,N_1859,N_454);
nand U4909 (N_4909,N_1918,N_2131);
nor U4910 (N_4910,N_1082,N_1215);
nand U4911 (N_4911,N_462,N_334);
or U4912 (N_4912,N_2399,N_2230);
and U4913 (N_4913,N_2471,N_133);
and U4914 (N_4914,N_2364,N_1071);
or U4915 (N_4915,N_2698,N_1845);
nor U4916 (N_4916,N_1519,N_1223);
or U4917 (N_4917,N_2884,N_1493);
nand U4918 (N_4918,N_2682,N_1014);
nor U4919 (N_4919,N_2809,N_1645);
nor U4920 (N_4920,N_513,N_1842);
and U4921 (N_4921,N_1610,N_1104);
and U4922 (N_4922,N_1251,N_1509);
nor U4923 (N_4923,N_476,N_1314);
nor U4924 (N_4924,N_2791,N_2947);
and U4925 (N_4925,N_2355,N_2806);
nand U4926 (N_4926,N_1776,N_484);
nor U4927 (N_4927,N_1580,N_2273);
nor U4928 (N_4928,N_1652,N_1515);
nand U4929 (N_4929,N_507,N_1533);
or U4930 (N_4930,N_713,N_2430);
nand U4931 (N_4931,N_1912,N_505);
nand U4932 (N_4932,N_2010,N_1661);
or U4933 (N_4933,N_1899,N_1366);
nand U4934 (N_4934,N_1275,N_217);
and U4935 (N_4935,N_2723,N_199);
nor U4936 (N_4936,N_1657,N_691);
xnor U4937 (N_4937,N_586,N_2468);
nand U4938 (N_4938,N_1794,N_337);
and U4939 (N_4939,N_88,N_376);
nor U4940 (N_4940,N_2964,N_2707);
and U4941 (N_4941,N_1864,N_2244);
nor U4942 (N_4942,N_1931,N_2778);
or U4943 (N_4943,N_2344,N_424);
nor U4944 (N_4944,N_2271,N_2588);
or U4945 (N_4945,N_655,N_513);
and U4946 (N_4946,N_2491,N_2742);
nor U4947 (N_4947,N_1956,N_2157);
nand U4948 (N_4948,N_1490,N_2923);
nor U4949 (N_4949,N_1354,N_938);
nor U4950 (N_4950,N_2414,N_1886);
nor U4951 (N_4951,N_2762,N_1770);
or U4952 (N_4952,N_2349,N_601);
and U4953 (N_4953,N_421,N_2007);
nand U4954 (N_4954,N_1375,N_2010);
and U4955 (N_4955,N_1100,N_47);
nand U4956 (N_4956,N_2372,N_1352);
and U4957 (N_4957,N_112,N_2678);
or U4958 (N_4958,N_2487,N_687);
nor U4959 (N_4959,N_2172,N_2243);
nand U4960 (N_4960,N_2625,N_2839);
or U4961 (N_4961,N_2350,N_2152);
nor U4962 (N_4962,N_1172,N_1913);
nand U4963 (N_4963,N_985,N_823);
nor U4964 (N_4964,N_2744,N_676);
and U4965 (N_4965,N_1888,N_18);
nand U4966 (N_4966,N_2758,N_1454);
nand U4967 (N_4967,N_2804,N_2702);
and U4968 (N_4968,N_2208,N_2873);
or U4969 (N_4969,N_1977,N_1992);
and U4970 (N_4970,N_2318,N_1619);
nor U4971 (N_4971,N_2254,N_904);
and U4972 (N_4972,N_671,N_1797);
and U4973 (N_4973,N_1103,N_1131);
nor U4974 (N_4974,N_337,N_2229);
nand U4975 (N_4975,N_353,N_1196);
nand U4976 (N_4976,N_1989,N_176);
nor U4977 (N_4977,N_2736,N_2759);
nor U4978 (N_4978,N_1238,N_1126);
nand U4979 (N_4979,N_145,N_1277);
and U4980 (N_4980,N_63,N_2228);
and U4981 (N_4981,N_2604,N_2028);
nor U4982 (N_4982,N_2628,N_2147);
and U4983 (N_4983,N_786,N_990);
and U4984 (N_4984,N_2201,N_828);
or U4985 (N_4985,N_1395,N_228);
and U4986 (N_4986,N_230,N_2225);
nand U4987 (N_4987,N_2365,N_802);
or U4988 (N_4988,N_147,N_831);
nand U4989 (N_4989,N_2912,N_370);
xor U4990 (N_4990,N_2081,N_1539);
nand U4991 (N_4991,N_2911,N_2185);
or U4992 (N_4992,N_2605,N_2151);
nor U4993 (N_4993,N_785,N_1316);
and U4994 (N_4994,N_160,N_2156);
or U4995 (N_4995,N_2879,N_1640);
nor U4996 (N_4996,N_2585,N_606);
and U4997 (N_4997,N_362,N_351);
or U4998 (N_4998,N_532,N_1952);
nand U4999 (N_4999,N_1643,N_1148);
or U5000 (N_5000,N_1906,N_1328);
and U5001 (N_5001,N_2991,N_2595);
nor U5002 (N_5002,N_1614,N_461);
and U5003 (N_5003,N_1534,N_938);
nor U5004 (N_5004,N_1162,N_730);
nor U5005 (N_5005,N_1370,N_1820);
nand U5006 (N_5006,N_903,N_1123);
or U5007 (N_5007,N_1755,N_500);
and U5008 (N_5008,N_2658,N_2824);
nor U5009 (N_5009,N_1141,N_1743);
nand U5010 (N_5010,N_399,N_171);
xor U5011 (N_5011,N_2319,N_1884);
nor U5012 (N_5012,N_1428,N_2559);
and U5013 (N_5013,N_1700,N_1547);
nor U5014 (N_5014,N_1238,N_1849);
nand U5015 (N_5015,N_888,N_253);
or U5016 (N_5016,N_1784,N_2514);
or U5017 (N_5017,N_2500,N_1110);
and U5018 (N_5018,N_586,N_1054);
and U5019 (N_5019,N_2567,N_2242);
and U5020 (N_5020,N_2158,N_1921);
or U5021 (N_5021,N_1303,N_1059);
nand U5022 (N_5022,N_700,N_1589);
nand U5023 (N_5023,N_2392,N_207);
nor U5024 (N_5024,N_537,N_1762);
nand U5025 (N_5025,N_842,N_2913);
and U5026 (N_5026,N_129,N_1270);
and U5027 (N_5027,N_957,N_901);
nor U5028 (N_5028,N_1626,N_2185);
or U5029 (N_5029,N_399,N_2165);
nand U5030 (N_5030,N_55,N_138);
and U5031 (N_5031,N_1004,N_383);
or U5032 (N_5032,N_852,N_2999);
nor U5033 (N_5033,N_1120,N_974);
or U5034 (N_5034,N_2280,N_214);
nand U5035 (N_5035,N_2670,N_2662);
nor U5036 (N_5036,N_2879,N_1815);
nor U5037 (N_5037,N_1347,N_1911);
nor U5038 (N_5038,N_2584,N_2353);
and U5039 (N_5039,N_832,N_1409);
nor U5040 (N_5040,N_2929,N_105);
nor U5041 (N_5041,N_1067,N_501);
nor U5042 (N_5042,N_630,N_1652);
or U5043 (N_5043,N_2474,N_108);
nor U5044 (N_5044,N_1866,N_1909);
or U5045 (N_5045,N_1673,N_437);
or U5046 (N_5046,N_1288,N_2282);
nand U5047 (N_5047,N_1385,N_1607);
nor U5048 (N_5048,N_1663,N_2);
nor U5049 (N_5049,N_2668,N_1291);
and U5050 (N_5050,N_51,N_1447);
nor U5051 (N_5051,N_2175,N_2903);
nand U5052 (N_5052,N_160,N_422);
and U5053 (N_5053,N_1220,N_34);
nor U5054 (N_5054,N_2769,N_2543);
or U5055 (N_5055,N_40,N_2879);
or U5056 (N_5056,N_156,N_1623);
or U5057 (N_5057,N_1131,N_69);
and U5058 (N_5058,N_2421,N_1439);
and U5059 (N_5059,N_1389,N_1138);
or U5060 (N_5060,N_869,N_2863);
or U5061 (N_5061,N_2602,N_2428);
nand U5062 (N_5062,N_2293,N_248);
and U5063 (N_5063,N_245,N_657);
nor U5064 (N_5064,N_1721,N_1372);
nor U5065 (N_5065,N_2982,N_1392);
nor U5066 (N_5066,N_1342,N_1500);
nor U5067 (N_5067,N_196,N_1040);
and U5068 (N_5068,N_2973,N_2880);
and U5069 (N_5069,N_1421,N_937);
nor U5070 (N_5070,N_722,N_1386);
and U5071 (N_5071,N_970,N_1775);
and U5072 (N_5072,N_1037,N_1017);
and U5073 (N_5073,N_1532,N_2294);
nor U5074 (N_5074,N_2958,N_2286);
nor U5075 (N_5075,N_1539,N_2632);
nand U5076 (N_5076,N_2474,N_2385);
nand U5077 (N_5077,N_610,N_369);
and U5078 (N_5078,N_45,N_2856);
nor U5079 (N_5079,N_2776,N_1368);
and U5080 (N_5080,N_196,N_1175);
or U5081 (N_5081,N_509,N_1109);
nand U5082 (N_5082,N_230,N_825);
nand U5083 (N_5083,N_2359,N_2761);
nand U5084 (N_5084,N_873,N_2092);
nand U5085 (N_5085,N_2689,N_2921);
nor U5086 (N_5086,N_1460,N_2472);
nand U5087 (N_5087,N_981,N_101);
and U5088 (N_5088,N_686,N_2751);
and U5089 (N_5089,N_2636,N_341);
or U5090 (N_5090,N_783,N_1882);
nand U5091 (N_5091,N_979,N_1603);
or U5092 (N_5092,N_588,N_2707);
and U5093 (N_5093,N_138,N_2121);
and U5094 (N_5094,N_702,N_294);
nand U5095 (N_5095,N_1369,N_545);
or U5096 (N_5096,N_1863,N_1057);
or U5097 (N_5097,N_2166,N_1448);
nand U5098 (N_5098,N_1008,N_1660);
nand U5099 (N_5099,N_1644,N_2542);
or U5100 (N_5100,N_1140,N_2500);
nand U5101 (N_5101,N_1602,N_2080);
and U5102 (N_5102,N_606,N_1509);
and U5103 (N_5103,N_219,N_1530);
and U5104 (N_5104,N_2228,N_1008);
nor U5105 (N_5105,N_1418,N_2658);
and U5106 (N_5106,N_559,N_730);
and U5107 (N_5107,N_1861,N_2318);
nand U5108 (N_5108,N_807,N_1262);
and U5109 (N_5109,N_225,N_2238);
xor U5110 (N_5110,N_1472,N_2940);
nor U5111 (N_5111,N_2651,N_1474);
or U5112 (N_5112,N_2485,N_873);
nor U5113 (N_5113,N_922,N_2826);
nand U5114 (N_5114,N_2886,N_1302);
nand U5115 (N_5115,N_1048,N_1339);
nand U5116 (N_5116,N_2666,N_997);
nor U5117 (N_5117,N_2033,N_648);
or U5118 (N_5118,N_1385,N_1574);
nand U5119 (N_5119,N_162,N_2612);
and U5120 (N_5120,N_563,N_1531);
nor U5121 (N_5121,N_1422,N_260);
or U5122 (N_5122,N_2635,N_2672);
xnor U5123 (N_5123,N_1841,N_89);
nand U5124 (N_5124,N_1403,N_1504);
and U5125 (N_5125,N_2009,N_639);
nand U5126 (N_5126,N_986,N_2685);
nand U5127 (N_5127,N_269,N_952);
and U5128 (N_5128,N_960,N_1104);
nand U5129 (N_5129,N_1813,N_1233);
nor U5130 (N_5130,N_716,N_703);
nand U5131 (N_5131,N_1269,N_1827);
or U5132 (N_5132,N_2664,N_1750);
or U5133 (N_5133,N_1873,N_551);
nor U5134 (N_5134,N_660,N_1899);
or U5135 (N_5135,N_2099,N_1683);
or U5136 (N_5136,N_66,N_811);
nor U5137 (N_5137,N_360,N_2279);
or U5138 (N_5138,N_1562,N_2295);
or U5139 (N_5139,N_233,N_175);
nor U5140 (N_5140,N_1512,N_301);
or U5141 (N_5141,N_423,N_224);
nor U5142 (N_5142,N_479,N_2582);
or U5143 (N_5143,N_817,N_1512);
nor U5144 (N_5144,N_1058,N_2218);
nor U5145 (N_5145,N_359,N_1190);
nor U5146 (N_5146,N_831,N_2319);
nor U5147 (N_5147,N_2865,N_2687);
or U5148 (N_5148,N_1551,N_2551);
nor U5149 (N_5149,N_544,N_2877);
nand U5150 (N_5150,N_112,N_784);
and U5151 (N_5151,N_218,N_2646);
or U5152 (N_5152,N_1719,N_222);
and U5153 (N_5153,N_2035,N_571);
nor U5154 (N_5154,N_2497,N_1024);
nor U5155 (N_5155,N_2645,N_2147);
nand U5156 (N_5156,N_1006,N_2003);
nor U5157 (N_5157,N_1521,N_1590);
or U5158 (N_5158,N_2264,N_960);
nand U5159 (N_5159,N_1346,N_2301);
and U5160 (N_5160,N_175,N_1647);
nand U5161 (N_5161,N_2654,N_2217);
and U5162 (N_5162,N_2336,N_2354);
or U5163 (N_5163,N_22,N_1641);
nor U5164 (N_5164,N_2429,N_17);
nand U5165 (N_5165,N_2800,N_214);
nor U5166 (N_5166,N_832,N_1178);
or U5167 (N_5167,N_256,N_282);
or U5168 (N_5168,N_2973,N_805);
and U5169 (N_5169,N_180,N_910);
or U5170 (N_5170,N_263,N_939);
and U5171 (N_5171,N_450,N_730);
or U5172 (N_5172,N_2241,N_132);
nor U5173 (N_5173,N_2843,N_1182);
or U5174 (N_5174,N_343,N_905);
nor U5175 (N_5175,N_2603,N_1351);
and U5176 (N_5176,N_2132,N_320);
and U5177 (N_5177,N_2791,N_2862);
and U5178 (N_5178,N_1071,N_801);
nand U5179 (N_5179,N_1920,N_1449);
xnor U5180 (N_5180,N_2913,N_2130);
or U5181 (N_5181,N_2544,N_571);
xor U5182 (N_5182,N_1356,N_454);
nand U5183 (N_5183,N_15,N_2963);
or U5184 (N_5184,N_1855,N_1478);
or U5185 (N_5185,N_13,N_309);
nor U5186 (N_5186,N_341,N_2728);
and U5187 (N_5187,N_926,N_2634);
or U5188 (N_5188,N_1243,N_2683);
or U5189 (N_5189,N_375,N_1881);
nor U5190 (N_5190,N_465,N_698);
nand U5191 (N_5191,N_901,N_2605);
and U5192 (N_5192,N_1538,N_1339);
or U5193 (N_5193,N_505,N_469);
nor U5194 (N_5194,N_2932,N_1261);
and U5195 (N_5195,N_1683,N_2188);
nor U5196 (N_5196,N_564,N_2778);
nand U5197 (N_5197,N_1571,N_2955);
nor U5198 (N_5198,N_253,N_1038);
or U5199 (N_5199,N_2659,N_2070);
nand U5200 (N_5200,N_1841,N_1365);
nor U5201 (N_5201,N_2780,N_1474);
and U5202 (N_5202,N_2439,N_1092);
and U5203 (N_5203,N_1724,N_1051);
nor U5204 (N_5204,N_1741,N_2214);
and U5205 (N_5205,N_1193,N_1720);
nor U5206 (N_5206,N_128,N_2327);
and U5207 (N_5207,N_811,N_1151);
nor U5208 (N_5208,N_580,N_2429);
and U5209 (N_5209,N_1042,N_281);
nand U5210 (N_5210,N_74,N_2772);
and U5211 (N_5211,N_422,N_875);
nand U5212 (N_5212,N_2084,N_42);
and U5213 (N_5213,N_1025,N_2962);
nand U5214 (N_5214,N_1258,N_1931);
and U5215 (N_5215,N_2839,N_2332);
nand U5216 (N_5216,N_1558,N_2106);
and U5217 (N_5217,N_1909,N_2113);
nand U5218 (N_5218,N_2786,N_1832);
or U5219 (N_5219,N_776,N_1080);
and U5220 (N_5220,N_1146,N_2123);
nand U5221 (N_5221,N_2574,N_2381);
nor U5222 (N_5222,N_1631,N_2016);
nor U5223 (N_5223,N_860,N_2993);
and U5224 (N_5224,N_1406,N_1951);
or U5225 (N_5225,N_774,N_1477);
or U5226 (N_5226,N_434,N_2876);
nand U5227 (N_5227,N_1665,N_2211);
or U5228 (N_5228,N_2355,N_1856);
and U5229 (N_5229,N_2953,N_1793);
nand U5230 (N_5230,N_1141,N_1295);
and U5231 (N_5231,N_353,N_1403);
and U5232 (N_5232,N_2307,N_1784);
or U5233 (N_5233,N_2640,N_1597);
nor U5234 (N_5234,N_255,N_1559);
or U5235 (N_5235,N_2666,N_531);
nand U5236 (N_5236,N_366,N_665);
and U5237 (N_5237,N_1876,N_717);
and U5238 (N_5238,N_451,N_2206);
nand U5239 (N_5239,N_1280,N_1615);
or U5240 (N_5240,N_751,N_1955);
nand U5241 (N_5241,N_1999,N_351);
or U5242 (N_5242,N_1940,N_1227);
nand U5243 (N_5243,N_2242,N_361);
or U5244 (N_5244,N_2920,N_936);
and U5245 (N_5245,N_2936,N_2533);
or U5246 (N_5246,N_196,N_174);
or U5247 (N_5247,N_1777,N_1147);
or U5248 (N_5248,N_2584,N_329);
nor U5249 (N_5249,N_2238,N_88);
nand U5250 (N_5250,N_396,N_2191);
and U5251 (N_5251,N_1487,N_2381);
nor U5252 (N_5252,N_1950,N_1631);
nand U5253 (N_5253,N_1116,N_2108);
nor U5254 (N_5254,N_1110,N_2932);
and U5255 (N_5255,N_2259,N_2045);
and U5256 (N_5256,N_873,N_1324);
nor U5257 (N_5257,N_1167,N_2847);
nor U5258 (N_5258,N_1083,N_2048);
and U5259 (N_5259,N_804,N_1519);
and U5260 (N_5260,N_979,N_1140);
and U5261 (N_5261,N_1924,N_590);
nand U5262 (N_5262,N_38,N_1259);
nand U5263 (N_5263,N_1020,N_708);
or U5264 (N_5264,N_1564,N_2341);
nor U5265 (N_5265,N_2558,N_1302);
nor U5266 (N_5266,N_191,N_920);
nand U5267 (N_5267,N_2697,N_955);
nand U5268 (N_5268,N_94,N_826);
nor U5269 (N_5269,N_1454,N_209);
or U5270 (N_5270,N_697,N_917);
and U5271 (N_5271,N_2736,N_2161);
nor U5272 (N_5272,N_471,N_2341);
nand U5273 (N_5273,N_744,N_591);
or U5274 (N_5274,N_2194,N_2517);
nor U5275 (N_5275,N_364,N_2790);
nor U5276 (N_5276,N_219,N_231);
or U5277 (N_5277,N_325,N_693);
or U5278 (N_5278,N_2256,N_1616);
or U5279 (N_5279,N_1765,N_2349);
nand U5280 (N_5280,N_1541,N_2951);
or U5281 (N_5281,N_1829,N_2587);
nand U5282 (N_5282,N_2066,N_399);
nand U5283 (N_5283,N_1306,N_75);
nor U5284 (N_5284,N_2141,N_1418);
or U5285 (N_5285,N_1073,N_395);
and U5286 (N_5286,N_124,N_1687);
nor U5287 (N_5287,N_1625,N_1569);
nand U5288 (N_5288,N_2208,N_131);
nand U5289 (N_5289,N_106,N_2766);
and U5290 (N_5290,N_1472,N_106);
nor U5291 (N_5291,N_1833,N_403);
nor U5292 (N_5292,N_2621,N_984);
and U5293 (N_5293,N_2917,N_2009);
nor U5294 (N_5294,N_458,N_2263);
or U5295 (N_5295,N_319,N_1448);
and U5296 (N_5296,N_1803,N_774);
and U5297 (N_5297,N_2396,N_258);
or U5298 (N_5298,N_520,N_1222);
nand U5299 (N_5299,N_1406,N_533);
and U5300 (N_5300,N_121,N_256);
nor U5301 (N_5301,N_577,N_62);
nand U5302 (N_5302,N_2093,N_433);
and U5303 (N_5303,N_2235,N_917);
nor U5304 (N_5304,N_1975,N_1623);
nand U5305 (N_5305,N_235,N_232);
or U5306 (N_5306,N_2492,N_2292);
nand U5307 (N_5307,N_696,N_385);
nand U5308 (N_5308,N_1426,N_2231);
and U5309 (N_5309,N_342,N_1391);
and U5310 (N_5310,N_587,N_2296);
and U5311 (N_5311,N_1556,N_2650);
nor U5312 (N_5312,N_2563,N_1488);
or U5313 (N_5313,N_1123,N_1709);
nor U5314 (N_5314,N_2036,N_1576);
nand U5315 (N_5315,N_74,N_2505);
nor U5316 (N_5316,N_2324,N_1339);
nor U5317 (N_5317,N_684,N_12);
nor U5318 (N_5318,N_2428,N_110);
or U5319 (N_5319,N_1570,N_2446);
or U5320 (N_5320,N_1543,N_2651);
nand U5321 (N_5321,N_2557,N_1843);
or U5322 (N_5322,N_1585,N_396);
or U5323 (N_5323,N_982,N_2902);
or U5324 (N_5324,N_369,N_41);
nand U5325 (N_5325,N_2257,N_155);
xor U5326 (N_5326,N_188,N_8);
and U5327 (N_5327,N_1648,N_545);
nor U5328 (N_5328,N_1008,N_1018);
and U5329 (N_5329,N_838,N_1163);
and U5330 (N_5330,N_1053,N_437);
and U5331 (N_5331,N_2575,N_1045);
nand U5332 (N_5332,N_2276,N_2156);
nor U5333 (N_5333,N_629,N_1657);
nand U5334 (N_5334,N_2628,N_2329);
nand U5335 (N_5335,N_2601,N_2567);
nor U5336 (N_5336,N_2646,N_2741);
nand U5337 (N_5337,N_1222,N_2872);
nor U5338 (N_5338,N_625,N_674);
and U5339 (N_5339,N_1309,N_1240);
nand U5340 (N_5340,N_1859,N_2424);
nand U5341 (N_5341,N_2030,N_260);
nor U5342 (N_5342,N_2793,N_2680);
or U5343 (N_5343,N_2279,N_2410);
nor U5344 (N_5344,N_2438,N_2858);
or U5345 (N_5345,N_308,N_2533);
nor U5346 (N_5346,N_1995,N_1332);
or U5347 (N_5347,N_706,N_1668);
nand U5348 (N_5348,N_937,N_2593);
or U5349 (N_5349,N_59,N_2186);
or U5350 (N_5350,N_1796,N_66);
nand U5351 (N_5351,N_787,N_278);
xor U5352 (N_5352,N_2222,N_1471);
and U5353 (N_5353,N_411,N_2472);
and U5354 (N_5354,N_2185,N_47);
or U5355 (N_5355,N_667,N_262);
or U5356 (N_5356,N_1145,N_1884);
or U5357 (N_5357,N_390,N_2644);
and U5358 (N_5358,N_730,N_2441);
nand U5359 (N_5359,N_1651,N_1189);
or U5360 (N_5360,N_2381,N_2886);
and U5361 (N_5361,N_1168,N_2606);
nand U5362 (N_5362,N_751,N_2937);
nand U5363 (N_5363,N_2645,N_1185);
nand U5364 (N_5364,N_119,N_1327);
nand U5365 (N_5365,N_768,N_1537);
nand U5366 (N_5366,N_2521,N_789);
or U5367 (N_5367,N_1813,N_2516);
nand U5368 (N_5368,N_2523,N_2332);
nand U5369 (N_5369,N_367,N_2220);
or U5370 (N_5370,N_722,N_1801);
nand U5371 (N_5371,N_1046,N_2423);
or U5372 (N_5372,N_625,N_2852);
and U5373 (N_5373,N_2924,N_1251);
nand U5374 (N_5374,N_1745,N_227);
nor U5375 (N_5375,N_2507,N_2375);
and U5376 (N_5376,N_896,N_2614);
nor U5377 (N_5377,N_2241,N_2507);
and U5378 (N_5378,N_2487,N_1947);
and U5379 (N_5379,N_1987,N_2711);
nor U5380 (N_5380,N_2097,N_1585);
nand U5381 (N_5381,N_603,N_795);
nand U5382 (N_5382,N_650,N_1285);
and U5383 (N_5383,N_557,N_2659);
or U5384 (N_5384,N_431,N_2903);
xor U5385 (N_5385,N_1661,N_282);
and U5386 (N_5386,N_2758,N_1062);
nor U5387 (N_5387,N_1692,N_1535);
or U5388 (N_5388,N_2461,N_364);
nand U5389 (N_5389,N_1529,N_932);
and U5390 (N_5390,N_389,N_925);
and U5391 (N_5391,N_2066,N_367);
nor U5392 (N_5392,N_426,N_803);
and U5393 (N_5393,N_885,N_584);
and U5394 (N_5394,N_2329,N_399);
and U5395 (N_5395,N_907,N_1160);
or U5396 (N_5396,N_1563,N_2763);
nor U5397 (N_5397,N_2509,N_623);
or U5398 (N_5398,N_2251,N_1576);
nor U5399 (N_5399,N_2363,N_484);
nor U5400 (N_5400,N_1809,N_1340);
nor U5401 (N_5401,N_920,N_2027);
nand U5402 (N_5402,N_1302,N_324);
or U5403 (N_5403,N_1358,N_1044);
nand U5404 (N_5404,N_2599,N_939);
nand U5405 (N_5405,N_1557,N_2499);
nand U5406 (N_5406,N_1162,N_1804);
nand U5407 (N_5407,N_2539,N_1451);
and U5408 (N_5408,N_1403,N_2174);
nor U5409 (N_5409,N_808,N_1143);
nand U5410 (N_5410,N_1835,N_1896);
nand U5411 (N_5411,N_885,N_1453);
and U5412 (N_5412,N_2695,N_181);
or U5413 (N_5413,N_2492,N_934);
or U5414 (N_5414,N_2266,N_1122);
nand U5415 (N_5415,N_2045,N_1628);
nand U5416 (N_5416,N_2052,N_1356);
or U5417 (N_5417,N_2716,N_1894);
nor U5418 (N_5418,N_323,N_2072);
nand U5419 (N_5419,N_2404,N_537);
xnor U5420 (N_5420,N_1853,N_2843);
nand U5421 (N_5421,N_2462,N_264);
nand U5422 (N_5422,N_2980,N_1151);
nor U5423 (N_5423,N_39,N_2826);
and U5424 (N_5424,N_2351,N_1810);
xnor U5425 (N_5425,N_1333,N_73);
nor U5426 (N_5426,N_2052,N_13);
nand U5427 (N_5427,N_99,N_1681);
nor U5428 (N_5428,N_1498,N_167);
or U5429 (N_5429,N_1590,N_2736);
or U5430 (N_5430,N_1272,N_2866);
or U5431 (N_5431,N_698,N_2657);
nand U5432 (N_5432,N_1313,N_1114);
or U5433 (N_5433,N_708,N_1516);
or U5434 (N_5434,N_2214,N_2149);
nand U5435 (N_5435,N_2825,N_588);
or U5436 (N_5436,N_846,N_1571);
nand U5437 (N_5437,N_1722,N_1841);
and U5438 (N_5438,N_2528,N_13);
and U5439 (N_5439,N_63,N_65);
and U5440 (N_5440,N_2309,N_2332);
xnor U5441 (N_5441,N_640,N_401);
and U5442 (N_5442,N_2344,N_1927);
and U5443 (N_5443,N_2931,N_2831);
nand U5444 (N_5444,N_2389,N_538);
nand U5445 (N_5445,N_2936,N_387);
and U5446 (N_5446,N_1975,N_2265);
nand U5447 (N_5447,N_1404,N_2407);
nor U5448 (N_5448,N_796,N_451);
or U5449 (N_5449,N_2224,N_183);
nand U5450 (N_5450,N_2064,N_1412);
nand U5451 (N_5451,N_1930,N_1105);
or U5452 (N_5452,N_1911,N_435);
and U5453 (N_5453,N_1991,N_560);
or U5454 (N_5454,N_2059,N_252);
nand U5455 (N_5455,N_1027,N_331);
nand U5456 (N_5456,N_728,N_892);
and U5457 (N_5457,N_126,N_1478);
or U5458 (N_5458,N_1338,N_387);
nand U5459 (N_5459,N_785,N_2465);
or U5460 (N_5460,N_1298,N_284);
and U5461 (N_5461,N_2658,N_103);
nor U5462 (N_5462,N_1740,N_1308);
nand U5463 (N_5463,N_1801,N_821);
nand U5464 (N_5464,N_825,N_2394);
nor U5465 (N_5465,N_1245,N_1481);
or U5466 (N_5466,N_243,N_295);
nor U5467 (N_5467,N_2992,N_1064);
nor U5468 (N_5468,N_2257,N_2933);
nand U5469 (N_5469,N_1047,N_1764);
or U5470 (N_5470,N_2544,N_1502);
nor U5471 (N_5471,N_2197,N_1011);
nand U5472 (N_5472,N_1437,N_1697);
or U5473 (N_5473,N_2936,N_1182);
nor U5474 (N_5474,N_2133,N_2411);
and U5475 (N_5475,N_2321,N_1189);
nor U5476 (N_5476,N_763,N_180);
nand U5477 (N_5477,N_1217,N_1227);
or U5478 (N_5478,N_2306,N_2926);
and U5479 (N_5479,N_853,N_468);
or U5480 (N_5480,N_188,N_2957);
and U5481 (N_5481,N_951,N_2577);
nor U5482 (N_5482,N_1805,N_2336);
or U5483 (N_5483,N_1956,N_220);
nand U5484 (N_5484,N_568,N_2224);
nand U5485 (N_5485,N_408,N_2808);
nand U5486 (N_5486,N_490,N_2776);
nor U5487 (N_5487,N_306,N_2146);
or U5488 (N_5488,N_1113,N_307);
and U5489 (N_5489,N_307,N_1907);
nand U5490 (N_5490,N_1247,N_1386);
or U5491 (N_5491,N_2133,N_860);
or U5492 (N_5492,N_2750,N_963);
nor U5493 (N_5493,N_831,N_97);
nand U5494 (N_5494,N_1438,N_341);
nor U5495 (N_5495,N_2125,N_1311);
nor U5496 (N_5496,N_1489,N_1613);
and U5497 (N_5497,N_2619,N_1594);
or U5498 (N_5498,N_96,N_1979);
and U5499 (N_5499,N_1579,N_299);
and U5500 (N_5500,N_2638,N_304);
nor U5501 (N_5501,N_2551,N_1732);
nand U5502 (N_5502,N_2206,N_2801);
and U5503 (N_5503,N_2587,N_2217);
and U5504 (N_5504,N_1065,N_2528);
nor U5505 (N_5505,N_2688,N_224);
or U5506 (N_5506,N_481,N_1188);
or U5507 (N_5507,N_520,N_411);
or U5508 (N_5508,N_280,N_1517);
and U5509 (N_5509,N_1434,N_1108);
and U5510 (N_5510,N_2701,N_792);
and U5511 (N_5511,N_86,N_2880);
nand U5512 (N_5512,N_2324,N_1401);
and U5513 (N_5513,N_2222,N_1707);
nor U5514 (N_5514,N_2794,N_1888);
and U5515 (N_5515,N_2451,N_2254);
or U5516 (N_5516,N_623,N_900);
nor U5517 (N_5517,N_747,N_1463);
nand U5518 (N_5518,N_486,N_1981);
nor U5519 (N_5519,N_52,N_2263);
and U5520 (N_5520,N_1883,N_2705);
xor U5521 (N_5521,N_2210,N_592);
nand U5522 (N_5522,N_1332,N_2428);
or U5523 (N_5523,N_2663,N_1947);
nand U5524 (N_5524,N_890,N_42);
or U5525 (N_5525,N_2737,N_1739);
or U5526 (N_5526,N_529,N_1786);
or U5527 (N_5527,N_1686,N_295);
and U5528 (N_5528,N_1820,N_2103);
or U5529 (N_5529,N_1137,N_2692);
and U5530 (N_5530,N_1278,N_823);
or U5531 (N_5531,N_732,N_89);
and U5532 (N_5532,N_2323,N_789);
nand U5533 (N_5533,N_321,N_584);
nand U5534 (N_5534,N_2932,N_2459);
nand U5535 (N_5535,N_1423,N_1330);
nand U5536 (N_5536,N_1601,N_678);
nor U5537 (N_5537,N_1181,N_316);
nor U5538 (N_5538,N_424,N_104);
nand U5539 (N_5539,N_1093,N_2501);
and U5540 (N_5540,N_222,N_389);
or U5541 (N_5541,N_86,N_738);
and U5542 (N_5542,N_46,N_986);
nand U5543 (N_5543,N_1459,N_2373);
nand U5544 (N_5544,N_2493,N_940);
nand U5545 (N_5545,N_959,N_1123);
nor U5546 (N_5546,N_1142,N_774);
nor U5547 (N_5547,N_1179,N_2925);
nor U5548 (N_5548,N_1076,N_1867);
nand U5549 (N_5549,N_2105,N_593);
and U5550 (N_5550,N_1981,N_1901);
and U5551 (N_5551,N_1052,N_2080);
nor U5552 (N_5552,N_1883,N_1150);
nor U5553 (N_5553,N_65,N_1977);
xnor U5554 (N_5554,N_2590,N_2247);
nor U5555 (N_5555,N_1246,N_574);
and U5556 (N_5556,N_248,N_1262);
or U5557 (N_5557,N_1240,N_2454);
xnor U5558 (N_5558,N_657,N_2474);
nor U5559 (N_5559,N_2736,N_980);
or U5560 (N_5560,N_2672,N_2037);
or U5561 (N_5561,N_2333,N_136);
and U5562 (N_5562,N_1004,N_674);
and U5563 (N_5563,N_1877,N_1825);
or U5564 (N_5564,N_2410,N_1999);
or U5565 (N_5565,N_507,N_1918);
nor U5566 (N_5566,N_2243,N_2016);
nor U5567 (N_5567,N_245,N_2321);
nor U5568 (N_5568,N_1193,N_2546);
or U5569 (N_5569,N_2416,N_2778);
nand U5570 (N_5570,N_478,N_2175);
and U5571 (N_5571,N_15,N_2417);
or U5572 (N_5572,N_2510,N_799);
nand U5573 (N_5573,N_898,N_1009);
or U5574 (N_5574,N_1464,N_1862);
or U5575 (N_5575,N_1700,N_2654);
or U5576 (N_5576,N_414,N_1349);
nand U5577 (N_5577,N_2028,N_780);
or U5578 (N_5578,N_1429,N_450);
nor U5579 (N_5579,N_234,N_406);
nand U5580 (N_5580,N_1595,N_1283);
nand U5581 (N_5581,N_61,N_392);
and U5582 (N_5582,N_1330,N_1855);
nand U5583 (N_5583,N_2072,N_1168);
and U5584 (N_5584,N_597,N_970);
nand U5585 (N_5585,N_2391,N_1696);
nand U5586 (N_5586,N_2977,N_1621);
or U5587 (N_5587,N_2938,N_2067);
nand U5588 (N_5588,N_1738,N_2562);
or U5589 (N_5589,N_1968,N_1736);
nor U5590 (N_5590,N_2759,N_2304);
nand U5591 (N_5591,N_457,N_2496);
and U5592 (N_5592,N_152,N_668);
nor U5593 (N_5593,N_756,N_278);
nor U5594 (N_5594,N_2722,N_1812);
or U5595 (N_5595,N_920,N_713);
nand U5596 (N_5596,N_911,N_380);
or U5597 (N_5597,N_2867,N_2926);
or U5598 (N_5598,N_2396,N_2697);
nand U5599 (N_5599,N_1738,N_808);
nand U5600 (N_5600,N_667,N_1012);
nor U5601 (N_5601,N_843,N_649);
nor U5602 (N_5602,N_984,N_1749);
and U5603 (N_5603,N_780,N_153);
nor U5604 (N_5604,N_330,N_350);
nand U5605 (N_5605,N_755,N_940);
and U5606 (N_5606,N_2242,N_1528);
nand U5607 (N_5607,N_2275,N_1673);
and U5608 (N_5608,N_403,N_837);
or U5609 (N_5609,N_2422,N_141);
or U5610 (N_5610,N_2658,N_702);
nand U5611 (N_5611,N_1897,N_2126);
and U5612 (N_5612,N_1896,N_338);
nand U5613 (N_5613,N_1384,N_1766);
nor U5614 (N_5614,N_1716,N_515);
nor U5615 (N_5615,N_2304,N_2207);
or U5616 (N_5616,N_440,N_1653);
nand U5617 (N_5617,N_2260,N_933);
nand U5618 (N_5618,N_2741,N_157);
or U5619 (N_5619,N_2036,N_1943);
nand U5620 (N_5620,N_2749,N_1212);
nand U5621 (N_5621,N_1980,N_1544);
nor U5622 (N_5622,N_106,N_2013);
nand U5623 (N_5623,N_780,N_2489);
nand U5624 (N_5624,N_984,N_1367);
and U5625 (N_5625,N_1333,N_1269);
and U5626 (N_5626,N_987,N_620);
or U5627 (N_5627,N_2765,N_1728);
or U5628 (N_5628,N_619,N_2583);
nand U5629 (N_5629,N_733,N_1072);
nor U5630 (N_5630,N_839,N_1056);
and U5631 (N_5631,N_2996,N_220);
or U5632 (N_5632,N_2039,N_558);
nand U5633 (N_5633,N_664,N_1076);
nand U5634 (N_5634,N_177,N_1006);
nand U5635 (N_5635,N_2046,N_732);
or U5636 (N_5636,N_1337,N_2855);
or U5637 (N_5637,N_439,N_242);
and U5638 (N_5638,N_739,N_817);
and U5639 (N_5639,N_2082,N_1724);
or U5640 (N_5640,N_2497,N_2020);
nor U5641 (N_5641,N_598,N_1339);
or U5642 (N_5642,N_1061,N_669);
and U5643 (N_5643,N_873,N_422);
xor U5644 (N_5644,N_2994,N_2082);
nand U5645 (N_5645,N_2378,N_2533);
nor U5646 (N_5646,N_344,N_308);
nor U5647 (N_5647,N_107,N_6);
and U5648 (N_5648,N_1112,N_2685);
nor U5649 (N_5649,N_2504,N_91);
or U5650 (N_5650,N_2826,N_923);
and U5651 (N_5651,N_1110,N_2119);
and U5652 (N_5652,N_1795,N_206);
and U5653 (N_5653,N_2111,N_2320);
or U5654 (N_5654,N_1348,N_355);
or U5655 (N_5655,N_980,N_2092);
xnor U5656 (N_5656,N_2534,N_2863);
nor U5657 (N_5657,N_1897,N_115);
or U5658 (N_5658,N_1870,N_144);
nand U5659 (N_5659,N_1297,N_2472);
nor U5660 (N_5660,N_1700,N_2833);
nor U5661 (N_5661,N_568,N_1333);
nor U5662 (N_5662,N_977,N_2928);
nor U5663 (N_5663,N_2586,N_236);
nor U5664 (N_5664,N_1707,N_2742);
nand U5665 (N_5665,N_1008,N_1174);
or U5666 (N_5666,N_2514,N_1849);
nor U5667 (N_5667,N_1021,N_866);
and U5668 (N_5668,N_214,N_915);
nand U5669 (N_5669,N_620,N_2291);
nand U5670 (N_5670,N_1856,N_1426);
and U5671 (N_5671,N_1494,N_998);
nor U5672 (N_5672,N_1091,N_1024);
or U5673 (N_5673,N_1717,N_2504);
nor U5674 (N_5674,N_1965,N_2608);
and U5675 (N_5675,N_2810,N_2246);
or U5676 (N_5676,N_2904,N_1280);
nand U5677 (N_5677,N_604,N_1036);
nor U5678 (N_5678,N_2565,N_286);
and U5679 (N_5679,N_427,N_405);
and U5680 (N_5680,N_1416,N_2708);
or U5681 (N_5681,N_1228,N_1844);
nand U5682 (N_5682,N_2751,N_1476);
and U5683 (N_5683,N_746,N_1640);
or U5684 (N_5684,N_2678,N_821);
and U5685 (N_5685,N_370,N_1643);
or U5686 (N_5686,N_592,N_2221);
or U5687 (N_5687,N_2625,N_2113);
and U5688 (N_5688,N_1155,N_267);
or U5689 (N_5689,N_2139,N_751);
nor U5690 (N_5690,N_2447,N_899);
nor U5691 (N_5691,N_1541,N_1505);
and U5692 (N_5692,N_2752,N_277);
nand U5693 (N_5693,N_1114,N_194);
nand U5694 (N_5694,N_2554,N_528);
and U5695 (N_5695,N_2802,N_1170);
nand U5696 (N_5696,N_2225,N_1800);
xor U5697 (N_5697,N_713,N_712);
nor U5698 (N_5698,N_1813,N_1223);
nand U5699 (N_5699,N_818,N_563);
and U5700 (N_5700,N_2059,N_2915);
nand U5701 (N_5701,N_1199,N_2231);
or U5702 (N_5702,N_521,N_2413);
and U5703 (N_5703,N_1583,N_1279);
and U5704 (N_5704,N_1705,N_482);
nor U5705 (N_5705,N_1676,N_1032);
or U5706 (N_5706,N_2959,N_790);
nor U5707 (N_5707,N_173,N_419);
and U5708 (N_5708,N_898,N_494);
nand U5709 (N_5709,N_1123,N_1011);
or U5710 (N_5710,N_1408,N_2438);
nor U5711 (N_5711,N_2052,N_1499);
or U5712 (N_5712,N_2503,N_2110);
and U5713 (N_5713,N_2620,N_1110);
and U5714 (N_5714,N_1442,N_246);
and U5715 (N_5715,N_2316,N_437);
or U5716 (N_5716,N_991,N_1257);
nand U5717 (N_5717,N_140,N_2844);
or U5718 (N_5718,N_1780,N_2155);
nor U5719 (N_5719,N_2842,N_790);
nor U5720 (N_5720,N_618,N_2848);
nor U5721 (N_5721,N_106,N_1834);
or U5722 (N_5722,N_754,N_70);
nor U5723 (N_5723,N_2250,N_1437);
nor U5724 (N_5724,N_1903,N_1587);
nor U5725 (N_5725,N_1944,N_86);
and U5726 (N_5726,N_2691,N_2142);
or U5727 (N_5727,N_1126,N_1986);
nand U5728 (N_5728,N_2201,N_2823);
nor U5729 (N_5729,N_541,N_2741);
nand U5730 (N_5730,N_406,N_1624);
nor U5731 (N_5731,N_1425,N_2936);
and U5732 (N_5732,N_1683,N_2546);
or U5733 (N_5733,N_2928,N_747);
or U5734 (N_5734,N_779,N_2862);
nor U5735 (N_5735,N_1206,N_311);
or U5736 (N_5736,N_1627,N_1196);
and U5737 (N_5737,N_2862,N_1366);
nor U5738 (N_5738,N_1510,N_1959);
nor U5739 (N_5739,N_2707,N_2669);
nand U5740 (N_5740,N_210,N_1323);
or U5741 (N_5741,N_1980,N_1661);
nand U5742 (N_5742,N_2689,N_2462);
or U5743 (N_5743,N_399,N_1685);
and U5744 (N_5744,N_2073,N_2136);
nor U5745 (N_5745,N_937,N_1508);
nand U5746 (N_5746,N_564,N_1688);
nand U5747 (N_5747,N_2693,N_2199);
nor U5748 (N_5748,N_1184,N_2650);
nand U5749 (N_5749,N_2704,N_416);
nor U5750 (N_5750,N_397,N_193);
or U5751 (N_5751,N_2214,N_2493);
nor U5752 (N_5752,N_2425,N_2302);
nand U5753 (N_5753,N_1554,N_356);
nand U5754 (N_5754,N_1855,N_1167);
or U5755 (N_5755,N_1308,N_2956);
or U5756 (N_5756,N_2999,N_2895);
and U5757 (N_5757,N_1880,N_1110);
or U5758 (N_5758,N_990,N_1087);
nor U5759 (N_5759,N_678,N_821);
and U5760 (N_5760,N_418,N_2061);
or U5761 (N_5761,N_2851,N_1103);
nand U5762 (N_5762,N_1039,N_2535);
and U5763 (N_5763,N_1236,N_414);
nand U5764 (N_5764,N_2642,N_2846);
nor U5765 (N_5765,N_1194,N_71);
nand U5766 (N_5766,N_1891,N_2777);
or U5767 (N_5767,N_1277,N_948);
nand U5768 (N_5768,N_949,N_887);
nor U5769 (N_5769,N_737,N_2173);
nor U5770 (N_5770,N_2384,N_999);
or U5771 (N_5771,N_1044,N_89);
and U5772 (N_5772,N_2027,N_1150);
nor U5773 (N_5773,N_1642,N_470);
and U5774 (N_5774,N_1696,N_2797);
or U5775 (N_5775,N_1557,N_1680);
nor U5776 (N_5776,N_875,N_142);
nor U5777 (N_5777,N_2492,N_90);
and U5778 (N_5778,N_505,N_1442);
nor U5779 (N_5779,N_189,N_2913);
or U5780 (N_5780,N_1540,N_1846);
or U5781 (N_5781,N_2542,N_2708);
and U5782 (N_5782,N_173,N_1252);
and U5783 (N_5783,N_1532,N_2081);
nand U5784 (N_5784,N_983,N_125);
nand U5785 (N_5785,N_771,N_1485);
nor U5786 (N_5786,N_460,N_2579);
nor U5787 (N_5787,N_2758,N_1987);
or U5788 (N_5788,N_2721,N_1459);
nand U5789 (N_5789,N_2313,N_2757);
nand U5790 (N_5790,N_2686,N_1056);
nand U5791 (N_5791,N_1842,N_811);
nor U5792 (N_5792,N_432,N_735);
and U5793 (N_5793,N_1445,N_720);
and U5794 (N_5794,N_93,N_441);
or U5795 (N_5795,N_1748,N_2095);
or U5796 (N_5796,N_2295,N_2377);
nand U5797 (N_5797,N_1959,N_816);
and U5798 (N_5798,N_1821,N_43);
or U5799 (N_5799,N_873,N_1269);
and U5800 (N_5800,N_2785,N_2665);
nor U5801 (N_5801,N_2834,N_2982);
and U5802 (N_5802,N_1803,N_1040);
and U5803 (N_5803,N_1653,N_836);
nand U5804 (N_5804,N_810,N_2426);
nand U5805 (N_5805,N_960,N_1091);
or U5806 (N_5806,N_1858,N_863);
or U5807 (N_5807,N_104,N_269);
or U5808 (N_5808,N_2193,N_737);
nand U5809 (N_5809,N_1260,N_2552);
and U5810 (N_5810,N_1205,N_2626);
nor U5811 (N_5811,N_149,N_1101);
nor U5812 (N_5812,N_1922,N_1281);
nand U5813 (N_5813,N_2621,N_2362);
and U5814 (N_5814,N_2419,N_771);
nand U5815 (N_5815,N_1694,N_2764);
nand U5816 (N_5816,N_573,N_376);
nand U5817 (N_5817,N_710,N_2802);
and U5818 (N_5818,N_1638,N_2191);
and U5819 (N_5819,N_2067,N_2924);
or U5820 (N_5820,N_2272,N_348);
nand U5821 (N_5821,N_698,N_2805);
xnor U5822 (N_5822,N_2393,N_2322);
or U5823 (N_5823,N_2087,N_1583);
and U5824 (N_5824,N_2074,N_108);
and U5825 (N_5825,N_2439,N_1642);
nand U5826 (N_5826,N_1480,N_1454);
or U5827 (N_5827,N_2648,N_1486);
nand U5828 (N_5828,N_2464,N_2688);
nand U5829 (N_5829,N_1625,N_114);
or U5830 (N_5830,N_2840,N_2474);
nand U5831 (N_5831,N_458,N_2731);
and U5832 (N_5832,N_2363,N_2125);
and U5833 (N_5833,N_2625,N_2572);
nand U5834 (N_5834,N_1820,N_437);
or U5835 (N_5835,N_1127,N_1838);
or U5836 (N_5836,N_2512,N_2807);
and U5837 (N_5837,N_674,N_1687);
nor U5838 (N_5838,N_714,N_2458);
nand U5839 (N_5839,N_1226,N_463);
and U5840 (N_5840,N_2121,N_2103);
or U5841 (N_5841,N_638,N_666);
or U5842 (N_5842,N_969,N_2111);
nor U5843 (N_5843,N_1802,N_2906);
nand U5844 (N_5844,N_1758,N_1091);
or U5845 (N_5845,N_517,N_1821);
and U5846 (N_5846,N_1344,N_2474);
nor U5847 (N_5847,N_81,N_2727);
nor U5848 (N_5848,N_2566,N_2834);
nand U5849 (N_5849,N_1683,N_340);
and U5850 (N_5850,N_1304,N_638);
xor U5851 (N_5851,N_1617,N_2192);
nor U5852 (N_5852,N_2228,N_60);
or U5853 (N_5853,N_2558,N_1298);
or U5854 (N_5854,N_1093,N_1176);
nand U5855 (N_5855,N_613,N_827);
and U5856 (N_5856,N_2748,N_1070);
nor U5857 (N_5857,N_1907,N_2038);
nor U5858 (N_5858,N_2340,N_261);
and U5859 (N_5859,N_1636,N_1457);
or U5860 (N_5860,N_459,N_970);
or U5861 (N_5861,N_905,N_1261);
nor U5862 (N_5862,N_593,N_2670);
nor U5863 (N_5863,N_405,N_472);
xnor U5864 (N_5864,N_1363,N_289);
nor U5865 (N_5865,N_2645,N_713);
and U5866 (N_5866,N_1789,N_543);
nor U5867 (N_5867,N_2038,N_842);
and U5868 (N_5868,N_1207,N_1374);
and U5869 (N_5869,N_2893,N_2322);
nor U5870 (N_5870,N_2031,N_2223);
nor U5871 (N_5871,N_2679,N_1314);
and U5872 (N_5872,N_1148,N_251);
or U5873 (N_5873,N_492,N_650);
nor U5874 (N_5874,N_1292,N_2630);
nor U5875 (N_5875,N_2454,N_1715);
or U5876 (N_5876,N_1423,N_1999);
and U5877 (N_5877,N_1590,N_1024);
and U5878 (N_5878,N_455,N_874);
nand U5879 (N_5879,N_843,N_1442);
nand U5880 (N_5880,N_534,N_516);
and U5881 (N_5881,N_2447,N_490);
and U5882 (N_5882,N_1270,N_1750);
nor U5883 (N_5883,N_2971,N_1214);
and U5884 (N_5884,N_2508,N_2194);
nand U5885 (N_5885,N_1253,N_2465);
nand U5886 (N_5886,N_1458,N_106);
nand U5887 (N_5887,N_243,N_565);
or U5888 (N_5888,N_1271,N_1059);
and U5889 (N_5889,N_2791,N_1099);
or U5890 (N_5890,N_2173,N_2423);
nand U5891 (N_5891,N_1974,N_1625);
or U5892 (N_5892,N_1089,N_2750);
or U5893 (N_5893,N_2799,N_345);
xor U5894 (N_5894,N_972,N_2829);
or U5895 (N_5895,N_125,N_2543);
and U5896 (N_5896,N_1115,N_2874);
or U5897 (N_5897,N_1604,N_1411);
or U5898 (N_5898,N_2909,N_2256);
nand U5899 (N_5899,N_780,N_55);
nor U5900 (N_5900,N_1510,N_2297);
or U5901 (N_5901,N_34,N_924);
and U5902 (N_5902,N_1754,N_781);
nor U5903 (N_5903,N_1226,N_1895);
or U5904 (N_5904,N_996,N_1458);
or U5905 (N_5905,N_124,N_1021);
or U5906 (N_5906,N_1611,N_1515);
nand U5907 (N_5907,N_217,N_921);
nor U5908 (N_5908,N_1563,N_2122);
nor U5909 (N_5909,N_1698,N_2780);
nand U5910 (N_5910,N_974,N_1226);
and U5911 (N_5911,N_105,N_2287);
and U5912 (N_5912,N_526,N_2344);
and U5913 (N_5913,N_2969,N_1973);
or U5914 (N_5914,N_185,N_320);
nor U5915 (N_5915,N_1445,N_158);
and U5916 (N_5916,N_1853,N_2463);
or U5917 (N_5917,N_53,N_171);
nor U5918 (N_5918,N_7,N_2048);
nand U5919 (N_5919,N_123,N_756);
nor U5920 (N_5920,N_545,N_197);
or U5921 (N_5921,N_1712,N_2238);
and U5922 (N_5922,N_1513,N_2032);
or U5923 (N_5923,N_1817,N_2949);
nand U5924 (N_5924,N_1729,N_2321);
or U5925 (N_5925,N_2567,N_1514);
nor U5926 (N_5926,N_852,N_2763);
xnor U5927 (N_5927,N_1927,N_105);
and U5928 (N_5928,N_540,N_1781);
nor U5929 (N_5929,N_1248,N_1861);
nor U5930 (N_5930,N_2137,N_1091);
and U5931 (N_5931,N_1993,N_2316);
and U5932 (N_5932,N_2037,N_1232);
or U5933 (N_5933,N_1233,N_1758);
or U5934 (N_5934,N_2122,N_42);
nand U5935 (N_5935,N_1225,N_1771);
nor U5936 (N_5936,N_1311,N_2467);
and U5937 (N_5937,N_2027,N_2176);
or U5938 (N_5938,N_1107,N_2937);
nand U5939 (N_5939,N_2684,N_2673);
nand U5940 (N_5940,N_1104,N_1771);
and U5941 (N_5941,N_632,N_1547);
nor U5942 (N_5942,N_1965,N_1934);
or U5943 (N_5943,N_267,N_2485);
or U5944 (N_5944,N_236,N_1973);
or U5945 (N_5945,N_587,N_2297);
and U5946 (N_5946,N_2705,N_1207);
or U5947 (N_5947,N_375,N_2869);
and U5948 (N_5948,N_2916,N_1060);
and U5949 (N_5949,N_1156,N_771);
nor U5950 (N_5950,N_1218,N_465);
nand U5951 (N_5951,N_472,N_2038);
nor U5952 (N_5952,N_2176,N_1065);
or U5953 (N_5953,N_2228,N_598);
or U5954 (N_5954,N_1299,N_1287);
nand U5955 (N_5955,N_843,N_219);
and U5956 (N_5956,N_331,N_1968);
nor U5957 (N_5957,N_897,N_1164);
and U5958 (N_5958,N_1248,N_1042);
or U5959 (N_5959,N_569,N_2684);
and U5960 (N_5960,N_1946,N_204);
nor U5961 (N_5961,N_2894,N_225);
or U5962 (N_5962,N_1265,N_1744);
or U5963 (N_5963,N_2506,N_1069);
nor U5964 (N_5964,N_2744,N_278);
nand U5965 (N_5965,N_172,N_2393);
nor U5966 (N_5966,N_772,N_2650);
and U5967 (N_5967,N_1578,N_1764);
or U5968 (N_5968,N_2663,N_350);
nand U5969 (N_5969,N_2849,N_2874);
nor U5970 (N_5970,N_2494,N_2648);
or U5971 (N_5971,N_2695,N_1144);
nor U5972 (N_5972,N_2839,N_1104);
nand U5973 (N_5973,N_2032,N_1893);
or U5974 (N_5974,N_2158,N_706);
nor U5975 (N_5975,N_193,N_488);
nor U5976 (N_5976,N_1458,N_351);
and U5977 (N_5977,N_903,N_909);
or U5978 (N_5978,N_786,N_2495);
and U5979 (N_5979,N_1674,N_89);
or U5980 (N_5980,N_2006,N_604);
or U5981 (N_5981,N_2779,N_2773);
nand U5982 (N_5982,N_795,N_1011);
nor U5983 (N_5983,N_2851,N_353);
nand U5984 (N_5984,N_1280,N_2443);
or U5985 (N_5985,N_2751,N_478);
nand U5986 (N_5986,N_1125,N_1019);
nand U5987 (N_5987,N_2603,N_2009);
and U5988 (N_5988,N_2689,N_1913);
and U5989 (N_5989,N_2507,N_711);
nand U5990 (N_5990,N_1053,N_2142);
nor U5991 (N_5991,N_2557,N_297);
and U5992 (N_5992,N_2426,N_2651);
nand U5993 (N_5993,N_2929,N_2057);
nor U5994 (N_5994,N_448,N_1954);
nand U5995 (N_5995,N_2187,N_16);
nor U5996 (N_5996,N_2845,N_2501);
or U5997 (N_5997,N_2185,N_1555);
or U5998 (N_5998,N_38,N_2686);
or U5999 (N_5999,N_740,N_2784);
nor U6000 (N_6000,N_4732,N_3462);
or U6001 (N_6001,N_3902,N_5123);
nand U6002 (N_6002,N_3921,N_5108);
nand U6003 (N_6003,N_4437,N_3154);
and U6004 (N_6004,N_5142,N_3246);
or U6005 (N_6005,N_4675,N_4332);
or U6006 (N_6006,N_5521,N_5444);
xor U6007 (N_6007,N_4508,N_3693);
and U6008 (N_6008,N_5164,N_4449);
and U6009 (N_6009,N_4703,N_3074);
or U6010 (N_6010,N_4409,N_5564);
nor U6011 (N_6011,N_4917,N_5978);
and U6012 (N_6012,N_5220,N_3495);
nand U6013 (N_6013,N_3493,N_5203);
or U6014 (N_6014,N_3285,N_4073);
nand U6015 (N_6015,N_4210,N_3291);
and U6016 (N_6016,N_5171,N_4289);
nor U6017 (N_6017,N_4140,N_3317);
nand U6018 (N_6018,N_3164,N_5163);
or U6019 (N_6019,N_4300,N_4813);
or U6020 (N_6020,N_4785,N_3449);
nor U6021 (N_6021,N_5532,N_5561);
nor U6022 (N_6022,N_4514,N_3406);
nand U6023 (N_6023,N_4923,N_4493);
or U6024 (N_6024,N_4781,N_4528);
or U6025 (N_6025,N_3894,N_4924);
nand U6026 (N_6026,N_3679,N_5659);
nor U6027 (N_6027,N_4033,N_5594);
xor U6028 (N_6028,N_5362,N_4836);
and U6029 (N_6029,N_3520,N_5194);
nand U6030 (N_6030,N_5461,N_5156);
nand U6031 (N_6031,N_5317,N_5051);
nor U6032 (N_6032,N_3436,N_5145);
or U6033 (N_6033,N_3990,N_3818);
or U6034 (N_6034,N_5871,N_4476);
and U6035 (N_6035,N_4318,N_4240);
and U6036 (N_6036,N_5588,N_5650);
or U6037 (N_6037,N_4253,N_4797);
and U6038 (N_6038,N_3985,N_3701);
or U6039 (N_6039,N_5700,N_4420);
or U6040 (N_6040,N_3724,N_3116);
nor U6041 (N_6041,N_4987,N_5434);
nand U6042 (N_6042,N_5961,N_4749);
and U6043 (N_6043,N_3385,N_3880);
and U6044 (N_6044,N_3260,N_5718);
or U6045 (N_6045,N_5773,N_3381);
and U6046 (N_6046,N_4855,N_5223);
nor U6047 (N_6047,N_5986,N_4395);
or U6048 (N_6048,N_4618,N_3720);
nor U6049 (N_6049,N_3315,N_3937);
and U6050 (N_6050,N_5404,N_3202);
or U6051 (N_6051,N_4990,N_5204);
nor U6052 (N_6052,N_4683,N_4358);
nand U6053 (N_6053,N_4879,N_4060);
nor U6054 (N_6054,N_3283,N_3755);
nand U6055 (N_6055,N_5852,N_5620);
nor U6056 (N_6056,N_3425,N_4739);
nor U6057 (N_6057,N_4848,N_3275);
nand U6058 (N_6058,N_5684,N_5769);
or U6059 (N_6059,N_3007,N_5116);
and U6060 (N_6060,N_5130,N_3564);
nand U6061 (N_6061,N_4662,N_3120);
or U6062 (N_6062,N_3538,N_5392);
or U6063 (N_6063,N_4901,N_5335);
nor U6064 (N_6064,N_3354,N_3587);
nand U6065 (N_6065,N_5431,N_5968);
nor U6066 (N_6066,N_3732,N_3307);
or U6067 (N_6067,N_5360,N_3253);
nor U6068 (N_6068,N_5936,N_3267);
nand U6069 (N_6069,N_3103,N_4546);
or U6070 (N_6070,N_3544,N_3515);
nand U6071 (N_6071,N_5102,N_4559);
nand U6072 (N_6072,N_3150,N_3930);
and U6073 (N_6073,N_4277,N_4203);
nor U6074 (N_6074,N_4489,N_4249);
or U6075 (N_6075,N_5579,N_4564);
and U6076 (N_6076,N_5008,N_3015);
nand U6077 (N_6077,N_3438,N_5315);
nor U6078 (N_6078,N_4650,N_3663);
nor U6079 (N_6079,N_4767,N_4267);
nor U6080 (N_6080,N_5613,N_5029);
and U6081 (N_6081,N_5602,N_4973);
or U6082 (N_6082,N_3613,N_5880);
nor U6083 (N_6083,N_4750,N_4204);
nand U6084 (N_6084,N_4666,N_5424);
nor U6085 (N_6085,N_4578,N_4967);
nor U6086 (N_6086,N_5664,N_4936);
nand U6087 (N_6087,N_4371,N_3974);
and U6088 (N_6088,N_4932,N_5001);
nor U6089 (N_6089,N_3736,N_4524);
nor U6090 (N_6090,N_5405,N_5074);
or U6091 (N_6091,N_3960,N_3459);
or U6092 (N_6092,N_4628,N_4684);
nand U6093 (N_6093,N_3813,N_3026);
or U6094 (N_6094,N_4688,N_3376);
or U6095 (N_6095,N_5550,N_4343);
xnor U6096 (N_6096,N_4174,N_3797);
xor U6097 (N_6097,N_3398,N_3653);
and U6098 (N_6098,N_3696,N_4895);
nand U6099 (N_6099,N_3888,N_3829);
nor U6100 (N_6100,N_4063,N_5635);
nand U6101 (N_6101,N_4101,N_3591);
and U6102 (N_6102,N_3590,N_3200);
or U6103 (N_6103,N_5776,N_3940);
nor U6104 (N_6104,N_5722,N_4560);
nand U6105 (N_6105,N_4036,N_5258);
and U6106 (N_6106,N_4758,N_3992);
or U6107 (N_6107,N_5125,N_5435);
nor U6108 (N_6108,N_3130,N_4288);
and U6109 (N_6109,N_3805,N_4861);
or U6110 (N_6110,N_4342,N_4893);
nand U6111 (N_6111,N_4606,N_4283);
or U6112 (N_6112,N_5436,N_3874);
nand U6113 (N_6113,N_3440,N_5349);
nor U6114 (N_6114,N_4229,N_5511);
and U6115 (N_6115,N_3656,N_3968);
or U6116 (N_6116,N_3830,N_5732);
nor U6117 (N_6117,N_4974,N_5144);
and U6118 (N_6118,N_5334,N_3109);
and U6119 (N_6119,N_5672,N_5980);
nand U6120 (N_6120,N_4028,N_5834);
nand U6121 (N_6121,N_4245,N_3083);
or U6122 (N_6122,N_3337,N_3999);
nand U6123 (N_6123,N_4513,N_4226);
or U6124 (N_6124,N_4287,N_5420);
or U6125 (N_6125,N_5823,N_5807);
nand U6126 (N_6126,N_4867,N_4935);
or U6127 (N_6127,N_4760,N_5158);
nor U6128 (N_6128,N_4580,N_5985);
nor U6129 (N_6129,N_5843,N_5239);
or U6130 (N_6130,N_3356,N_3110);
and U6131 (N_6131,N_3197,N_4938);
nor U6132 (N_6132,N_5497,N_3998);
nand U6133 (N_6133,N_5294,N_4573);
and U6134 (N_6134,N_3382,N_5378);
or U6135 (N_6135,N_3262,N_5046);
nand U6136 (N_6136,N_3734,N_5249);
nand U6137 (N_6137,N_4059,N_4829);
and U6138 (N_6138,N_5087,N_4875);
or U6139 (N_6139,N_3100,N_3251);
and U6140 (N_6140,N_5548,N_3121);
and U6141 (N_6141,N_5311,N_5148);
or U6142 (N_6142,N_3205,N_5669);
nor U6143 (N_6143,N_5296,N_3394);
nor U6144 (N_6144,N_3667,N_5456);
nand U6145 (N_6145,N_5831,N_5792);
and U6146 (N_6146,N_3136,N_4016);
or U6147 (N_6147,N_3081,N_3966);
nor U6148 (N_6148,N_4756,N_4706);
and U6149 (N_6149,N_5056,N_4160);
and U6150 (N_6150,N_3391,N_5339);
or U6151 (N_6151,N_4219,N_3692);
and U6152 (N_6152,N_5066,N_3341);
and U6153 (N_6153,N_4214,N_4223);
nand U6154 (N_6154,N_5887,N_5821);
or U6155 (N_6155,N_3632,N_3107);
nand U6156 (N_6156,N_4152,N_4091);
and U6157 (N_6157,N_5925,N_5332);
or U6158 (N_6158,N_4379,N_4693);
xnor U6159 (N_6159,N_5859,N_4215);
and U6160 (N_6160,N_4045,N_3240);
nand U6161 (N_6161,N_4362,N_3627);
and U6162 (N_6162,N_5288,N_3957);
or U6163 (N_6163,N_5581,N_3188);
and U6164 (N_6164,N_4029,N_3129);
nand U6165 (N_6165,N_3481,N_5812);
nor U6166 (N_6166,N_3997,N_3365);
and U6167 (N_6167,N_3645,N_5643);
or U6168 (N_6168,N_4090,N_5027);
nor U6169 (N_6169,N_4579,N_4419);
or U6170 (N_6170,N_5297,N_5896);
or U6171 (N_6171,N_3155,N_5313);
and U6172 (N_6172,N_3447,N_5055);
or U6173 (N_6173,N_4122,N_4525);
nor U6174 (N_6174,N_3383,N_4238);
and U6175 (N_6175,N_3794,N_5729);
and U6176 (N_6176,N_4327,N_4868);
or U6177 (N_6177,N_5445,N_5942);
nor U6178 (N_6178,N_5146,N_5777);
nand U6179 (N_6179,N_5480,N_3118);
nor U6180 (N_6180,N_3640,N_5566);
nor U6181 (N_6181,N_3361,N_4657);
nor U6182 (N_6182,N_4046,N_4507);
nand U6183 (N_6183,N_5844,N_5440);
nand U6184 (N_6184,N_3045,N_3994);
nor U6185 (N_6185,N_4412,N_4772);
nand U6186 (N_6186,N_3924,N_3507);
and U6187 (N_6187,N_5582,N_5346);
nor U6188 (N_6188,N_3835,N_3745);
nand U6189 (N_6189,N_5500,N_5540);
nand U6190 (N_6190,N_3738,N_4164);
xor U6191 (N_6191,N_3423,N_5610);
and U6192 (N_6192,N_4766,N_5873);
nand U6193 (N_6193,N_3841,N_3056);
and U6194 (N_6194,N_4891,N_5067);
nor U6195 (N_6195,N_5916,N_5685);
nand U6196 (N_6196,N_4558,N_3752);
nor U6197 (N_6197,N_4190,N_4506);
nor U6198 (N_6198,N_3928,N_4143);
and U6199 (N_6199,N_5592,N_4926);
nor U6200 (N_6200,N_5257,N_3411);
nand U6201 (N_6201,N_3198,N_3542);
nor U6202 (N_6202,N_5463,N_4397);
nor U6203 (N_6203,N_3364,N_5675);
or U6204 (N_6204,N_5817,N_5671);
nand U6205 (N_6205,N_5121,N_4236);
or U6206 (N_6206,N_5260,N_4451);
and U6207 (N_6207,N_4070,N_3788);
and U6208 (N_6208,N_5374,N_5907);
nand U6209 (N_6209,N_5606,N_5176);
nand U6210 (N_6210,N_3525,N_4312);
and U6211 (N_6211,N_5923,N_3360);
nor U6212 (N_6212,N_5356,N_4414);
and U6213 (N_6213,N_5959,N_4590);
nand U6214 (N_6214,N_5960,N_4039);
or U6215 (N_6215,N_3430,N_5997);
and U6216 (N_6216,N_4316,N_5818);
or U6217 (N_6217,N_3869,N_3967);
or U6218 (N_6218,N_5273,N_3000);
or U6219 (N_6219,N_5202,N_5282);
nor U6220 (N_6220,N_3404,N_5353);
nand U6221 (N_6221,N_5251,N_3153);
nand U6222 (N_6222,N_5231,N_4784);
and U6223 (N_6223,N_3670,N_4697);
nand U6224 (N_6224,N_4981,N_4268);
nor U6225 (N_6225,N_4716,N_5167);
or U6226 (N_6226,N_5133,N_4272);
nor U6227 (N_6227,N_5028,N_5612);
nand U6228 (N_6228,N_3102,N_4297);
nor U6229 (N_6229,N_5169,N_5198);
and U6230 (N_6230,N_5652,N_3798);
or U6231 (N_6231,N_4888,N_4290);
nand U6232 (N_6232,N_3088,N_5963);
and U6233 (N_6233,N_5229,N_5021);
nand U6234 (N_6234,N_4357,N_4156);
or U6235 (N_6235,N_5357,N_3929);
nand U6236 (N_6236,N_4771,N_5319);
nor U6237 (N_6237,N_5882,N_4299);
nand U6238 (N_6238,N_5484,N_4361);
or U6239 (N_6239,N_3393,N_5149);
or U6240 (N_6240,N_4481,N_5023);
and U6241 (N_6241,N_3823,N_4882);
or U6242 (N_6242,N_5017,N_4149);
or U6243 (N_6243,N_3846,N_3223);
or U6244 (N_6244,N_4824,N_4473);
and U6245 (N_6245,N_4687,N_5003);
and U6246 (N_6246,N_5721,N_3889);
or U6247 (N_6247,N_3470,N_5250);
xor U6248 (N_6248,N_3886,N_3655);
nand U6249 (N_6249,N_4814,N_4776);
or U6250 (N_6250,N_3221,N_5478);
or U6251 (N_6251,N_3322,N_4334);
and U6252 (N_6252,N_5479,N_4609);
and U6253 (N_6253,N_5651,N_3375);
nor U6254 (N_6254,N_3858,N_4890);
nor U6255 (N_6255,N_5798,N_5979);
or U6256 (N_6256,N_3479,N_5944);
nand U6257 (N_6257,N_4341,N_3292);
nor U6258 (N_6258,N_5838,N_3448);
nor U6259 (N_6259,N_3592,N_3731);
and U6260 (N_6260,N_5900,N_3066);
or U6261 (N_6261,N_4040,N_4542);
nor U6262 (N_6262,N_5795,N_5004);
nor U6263 (N_6263,N_3139,N_5302);
or U6264 (N_6264,N_3638,N_4443);
xnor U6265 (N_6265,N_3560,N_5941);
or U6266 (N_6266,N_4761,N_5926);
nor U6267 (N_6267,N_4945,N_5493);
nor U6268 (N_6268,N_4920,N_4900);
nand U6269 (N_6269,N_4872,N_4404);
nand U6270 (N_6270,N_3913,N_4589);
or U6271 (N_6271,N_4155,N_3273);
or U6272 (N_6272,N_4595,N_3137);
nor U6273 (N_6273,N_3089,N_4479);
nand U6274 (N_6274,N_4636,N_5030);
nor U6275 (N_6275,N_3885,N_3218);
or U6276 (N_6276,N_3134,N_5967);
nand U6277 (N_6277,N_3023,N_4241);
and U6278 (N_6278,N_3201,N_5965);
and U6279 (N_6279,N_5530,N_5165);
and U6280 (N_6280,N_3467,N_4392);
and U6281 (N_6281,N_3789,N_5050);
or U6282 (N_6282,N_4584,N_4025);
nand U6283 (N_6283,N_4637,N_4077);
nand U6284 (N_6284,N_5553,N_3384);
or U6285 (N_6285,N_5499,N_5457);
or U6286 (N_6286,N_5212,N_3568);
nand U6287 (N_6287,N_4411,N_3122);
nor U6288 (N_6288,N_5869,N_3780);
nand U6289 (N_6289,N_3219,N_4458);
and U6290 (N_6290,N_5233,N_3511);
and U6291 (N_6291,N_4531,N_5574);
nor U6292 (N_6292,N_5932,N_5059);
and U6293 (N_6293,N_5832,N_3435);
nand U6294 (N_6294,N_4220,N_3485);
or U6295 (N_6295,N_3643,N_3681);
or U6296 (N_6296,N_5623,N_3242);
nand U6297 (N_6297,N_5136,N_5597);
or U6298 (N_6298,N_3625,N_3257);
nor U6299 (N_6299,N_3238,N_4218);
and U6300 (N_6300,N_4802,N_5438);
and U6301 (N_6301,N_5731,N_5062);
and U6302 (N_6302,N_3141,N_5042);
nand U6303 (N_6303,N_4992,N_4660);
nor U6304 (N_6304,N_3917,N_3977);
and U6305 (N_6305,N_5803,N_3417);
nand U6306 (N_6306,N_4496,N_5641);
nor U6307 (N_6307,N_4355,N_3502);
and U6308 (N_6308,N_5575,N_3003);
nor U6309 (N_6309,N_5006,N_5549);
and U6310 (N_6310,N_5510,N_5019);
xor U6311 (N_6311,N_5201,N_3397);
nand U6312 (N_6312,N_4423,N_4654);
or U6313 (N_6313,N_3464,N_5507);
and U6314 (N_6314,N_5426,N_4398);
and U6315 (N_6315,N_4511,N_5611);
and U6316 (N_6316,N_4344,N_4642);
nand U6317 (N_6317,N_4625,N_5089);
nor U6318 (N_6318,N_4087,N_5138);
nand U6319 (N_6319,N_5088,N_3595);
nand U6320 (N_6320,N_4723,N_5767);
or U6321 (N_6321,N_5232,N_5536);
nor U6322 (N_6322,N_5236,N_4141);
nand U6323 (N_6323,N_3688,N_4259);
and U6324 (N_6324,N_3490,N_5793);
or U6325 (N_6325,N_4158,N_3804);
or U6326 (N_6326,N_4533,N_5488);
nand U6327 (N_6327,N_3708,N_5477);
and U6328 (N_6328,N_3290,N_5902);
nor U6329 (N_6329,N_3105,N_5955);
nand U6330 (N_6330,N_4535,N_4971);
nand U6331 (N_6331,N_5207,N_3882);
or U6332 (N_6332,N_5556,N_5780);
nand U6333 (N_6333,N_3896,N_3092);
nor U6334 (N_6334,N_3875,N_4770);
or U6335 (N_6335,N_5318,N_5157);
nand U6336 (N_6336,N_5054,N_4322);
nor U6337 (N_6337,N_4233,N_4425);
nor U6338 (N_6338,N_4186,N_3450);
nor U6339 (N_6339,N_4934,N_4474);
xnor U6340 (N_6340,N_3048,N_3282);
nand U6341 (N_6341,N_5235,N_4517);
nor U6342 (N_6342,N_3060,N_4389);
and U6343 (N_6343,N_5244,N_4258);
and U6344 (N_6344,N_5390,N_5962);
or U6345 (N_6345,N_4187,N_5337);
nand U6346 (N_6346,N_3304,N_3578);
nand U6347 (N_6347,N_5515,N_4664);
and U6348 (N_6348,N_4747,N_3849);
and U6349 (N_6349,N_4231,N_3582);
or U6350 (N_6350,N_3543,N_3715);
or U6351 (N_6351,N_5712,N_3265);
nand U6352 (N_6352,N_4178,N_5376);
nand U6353 (N_6353,N_4250,N_4588);
nand U6354 (N_6354,N_3842,N_5211);
and U6355 (N_6355,N_5421,N_5654);
or U6356 (N_6356,N_3839,N_3621);
and U6357 (N_6357,N_3635,N_3295);
nor U6358 (N_6358,N_5576,N_4892);
nand U6359 (N_6359,N_3451,N_3801);
and U6360 (N_6360,N_4899,N_3539);
nand U6361 (N_6361,N_4448,N_3503);
and U6362 (N_6362,N_5016,N_3348);
nor U6363 (N_6363,N_3009,N_3687);
and U6364 (N_6364,N_4224,N_3949);
and U6365 (N_6365,N_5455,N_3445);
nor U6366 (N_6366,N_4189,N_3766);
or U6367 (N_6367,N_3526,N_4541);
nand U6368 (N_6368,N_4969,N_4304);
nand U6369 (N_6369,N_5482,N_4646);
nand U6370 (N_6370,N_4720,N_3575);
or U6371 (N_6371,N_3099,N_5987);
and U6372 (N_6372,N_5316,N_4366);
nand U6373 (N_6373,N_4310,N_4175);
nor U6374 (N_6374,N_3334,N_3871);
nand U6375 (N_6375,N_5905,N_5913);
and U6376 (N_6376,N_4594,N_5632);
or U6377 (N_6377,N_4939,N_5662);
or U6378 (N_6378,N_4490,N_4275);
nand U6379 (N_6379,N_5185,N_4865);
and U6380 (N_6380,N_3729,N_5783);
nor U6381 (N_6381,N_3236,N_4007);
and U6382 (N_6382,N_3837,N_3243);
nand U6383 (N_6383,N_5143,N_4375);
and U6384 (N_6384,N_4738,N_3025);
or U6385 (N_6385,N_3303,N_5881);
nor U6386 (N_6386,N_5551,N_4799);
nor U6387 (N_6387,N_4078,N_3561);
nor U6388 (N_6388,N_4418,N_3194);
or U6389 (N_6389,N_4031,N_5763);
nand U6390 (N_6390,N_3831,N_4196);
or U6391 (N_6391,N_5155,N_5544);
nor U6392 (N_6392,N_3697,N_5329);
nor U6393 (N_6393,N_4922,N_5765);
or U6394 (N_6394,N_5183,N_4575);
nor U6395 (N_6395,N_5772,N_5717);
and U6396 (N_6396,N_4012,N_3821);
nand U6397 (N_6397,N_3085,N_5940);
nand U6398 (N_6398,N_3714,N_4096);
or U6399 (N_6399,N_5104,N_4326);
and U6400 (N_6400,N_3313,N_4577);
or U6401 (N_6401,N_3603,N_3138);
nand U6402 (N_6402,N_3234,N_5490);
nor U6403 (N_6403,N_5846,N_5888);
and U6404 (N_6404,N_4886,N_5071);
nand U6405 (N_6405,N_3021,N_4377);
nand U6406 (N_6406,N_5206,N_5636);
nor U6407 (N_6407,N_3353,N_3115);
or U6408 (N_6408,N_3328,N_3702);
nor U6409 (N_6409,N_5724,N_3864);
or U6410 (N_6410,N_4921,N_5058);
xnor U6411 (N_6411,N_4555,N_3387);
and U6412 (N_6412,N_3735,N_5147);
nor U6413 (N_6413,N_4370,N_4933);
nand U6414 (N_6414,N_5072,N_5689);
xnor U6415 (N_6415,N_4736,N_3605);
nand U6416 (N_6416,N_3860,N_4906);
and U6417 (N_6417,N_4024,N_5366);
and U6418 (N_6418,N_3647,N_5922);
nor U6419 (N_6419,N_5842,N_5467);
and U6420 (N_6420,N_3634,N_5061);
nand U6421 (N_6421,N_5523,N_4500);
nor U6422 (N_6422,N_5808,N_3458);
xor U6423 (N_6423,N_3898,N_4094);
nand U6424 (N_6424,N_5683,N_3787);
nand U6425 (N_6425,N_4167,N_5190);
and U6426 (N_6426,N_5214,N_4305);
nand U6427 (N_6427,N_4438,N_3807);
and U6428 (N_6428,N_5791,N_4058);
nand U6429 (N_6429,N_5603,N_4957);
and U6430 (N_6430,N_4616,N_3817);
nand U6431 (N_6431,N_3877,N_5991);
and U6432 (N_6432,N_5278,N_5084);
nand U6433 (N_6433,N_5753,N_5973);
and U6434 (N_6434,N_4393,N_4453);
and U6435 (N_6435,N_5310,N_4126);
nor U6436 (N_6436,N_3711,N_3456);
and U6437 (N_6437,N_3019,N_3895);
and U6438 (N_6438,N_4503,N_5928);
nor U6439 (N_6439,N_3927,N_5835);
or U6440 (N_6440,N_4896,N_5075);
nor U6441 (N_6441,N_5172,N_5441);
or U6442 (N_6442,N_4842,N_3565);
nor U6443 (N_6443,N_4192,N_5934);
and U6444 (N_6444,N_3707,N_5999);
nor U6445 (N_6445,N_4837,N_4498);
or U6446 (N_6446,N_3017,N_5953);
nor U6447 (N_6447,N_4242,N_5267);
nor U6448 (N_6448,N_3727,N_5387);
nor U6449 (N_6449,N_3832,N_3691);
nor U6450 (N_6450,N_4796,N_3466);
and U6451 (N_6451,N_4884,N_5646);
nor U6452 (N_6452,N_4860,N_3016);
and U6453 (N_6453,N_3596,N_3989);
or U6454 (N_6454,N_3649,N_4043);
nand U6455 (N_6455,N_4424,N_4047);
nor U6456 (N_6456,N_4733,N_4839);
nor U6457 (N_6457,N_3043,N_3547);
and U6458 (N_6458,N_5741,N_5414);
or U6459 (N_6459,N_4455,N_5118);
or U6460 (N_6460,N_3710,N_4599);
or U6461 (N_6461,N_3359,N_5674);
nor U6462 (N_6462,N_5680,N_4819);
nor U6463 (N_6463,N_5621,N_4112);
and U6464 (N_6464,N_3269,N_4456);
nand U6465 (N_6465,N_4937,N_4661);
nand U6466 (N_6466,N_4432,N_4308);
and U6467 (N_6467,N_5520,N_5789);
nor U6468 (N_6468,N_5264,N_4365);
nand U6469 (N_6469,N_5425,N_3601);
and U6470 (N_6470,N_4065,N_5697);
nor U6471 (N_6471,N_3271,N_5868);
nand U6472 (N_6472,N_4116,N_5344);
and U6473 (N_6473,N_3712,N_4543);
nand U6474 (N_6474,N_5607,N_4572);
and U6475 (N_6475,N_4009,N_4124);
or U6476 (N_6476,N_5415,N_4041);
and U6477 (N_6477,N_3733,N_4339);
nand U6478 (N_6478,N_4347,N_5759);
nand U6479 (N_6479,N_4279,N_4742);
nand U6480 (N_6480,N_3824,N_4569);
or U6481 (N_6481,N_3344,N_4880);
nor U6482 (N_6482,N_5644,N_5633);
or U6483 (N_6483,N_3469,N_3132);
and U6484 (N_6484,N_5982,N_3244);
and U6485 (N_6485,N_3220,N_4519);
and U6486 (N_6486,N_4821,N_3576);
nor U6487 (N_6487,N_5041,N_4144);
nor U6488 (N_6488,N_4239,N_5320);
nand U6489 (N_6489,N_3222,N_5738);
nor U6490 (N_6490,N_3075,N_5129);
nor U6491 (N_6491,N_4908,N_3577);
nand U6492 (N_6492,N_4306,N_5901);
or U6493 (N_6493,N_4185,N_3033);
or U6494 (N_6494,N_5095,N_5906);
nor U6495 (N_6495,N_4658,N_3339);
nand U6496 (N_6496,N_5625,N_3029);
and U6497 (N_6497,N_5449,N_5383);
nor U6498 (N_6498,N_4360,N_3551);
nor U6499 (N_6499,N_3918,N_3604);
or U6500 (N_6500,N_5252,N_5281);
nand U6501 (N_6501,N_3190,N_5528);
or U6502 (N_6502,N_5292,N_3465);
nand U6503 (N_6503,N_3623,N_3996);
and U6504 (N_6504,N_3529,N_5598);
or U6505 (N_6505,N_5043,N_4296);
and U6506 (N_6506,N_4367,N_3501);
nor U6507 (N_6507,N_4777,N_4261);
nand U6508 (N_6508,N_3333,N_5326);
nand U6509 (N_6509,N_3975,N_5083);
nand U6510 (N_6510,N_4368,N_3408);
nor U6511 (N_6511,N_3644,N_3034);
nor U6512 (N_6512,N_4273,N_3619);
nand U6513 (N_6513,N_3747,N_4930);
nor U6514 (N_6514,N_5723,N_5430);
nand U6515 (N_6515,N_3174,N_4102);
nand U6516 (N_6516,N_4916,N_5860);
or U6517 (N_6517,N_5411,N_4006);
or U6518 (N_6518,N_3915,N_3810);
or U6519 (N_6519,N_5498,N_3528);
or U6520 (N_6520,N_3047,N_5401);
nor U6521 (N_6521,N_5305,N_5538);
and U6522 (N_6522,N_3719,N_4913);
and U6523 (N_6523,N_3855,N_4851);
nand U6524 (N_6524,N_5663,N_3239);
nand U6525 (N_6525,N_5673,N_5175);
and U6526 (N_6526,N_3757,N_4051);
nand U6527 (N_6527,N_3177,N_4833);
xor U6528 (N_6528,N_5847,N_4812);
or U6529 (N_6529,N_3053,N_5048);
xor U6530 (N_6530,N_3487,N_3002);
and U6531 (N_6531,N_4176,N_3216);
nand U6532 (N_6532,N_5943,N_5178);
and U6533 (N_6533,N_4406,N_4807);
nor U6534 (N_6534,N_5580,N_4044);
nand U6535 (N_6535,N_4972,N_4105);
and U6536 (N_6536,N_3598,N_3452);
nor U6537 (N_6537,N_5693,N_3039);
and U6538 (N_6538,N_3617,N_4056);
nand U6539 (N_6539,N_4447,N_3453);
and U6540 (N_6540,N_3434,N_5708);
or U6541 (N_6541,N_3978,N_5716);
nor U6542 (N_6542,N_4854,N_3897);
nor U6543 (N_6543,N_5891,N_3148);
nand U6544 (N_6544,N_5745,N_3211);
nand U6545 (N_6545,N_4399,N_5395);
nor U6546 (N_6546,N_5475,N_4165);
or U6547 (N_6547,N_4243,N_3159);
and U6548 (N_6548,N_4670,N_3294);
and U6549 (N_6549,N_5168,N_3004);
or U6550 (N_6550,N_3351,N_4137);
and U6551 (N_6551,N_3834,N_3133);
or U6552 (N_6552,N_5757,N_5454);
and U6553 (N_6553,N_5892,N_4602);
and U6554 (N_6554,N_3983,N_3883);
nand U6555 (N_6555,N_4717,N_3076);
and U6556 (N_6556,N_3600,N_4597);
and U6557 (N_6557,N_5166,N_5849);
nor U6558 (N_6558,N_5851,N_5487);
nor U6559 (N_6559,N_4857,N_4801);
and U6560 (N_6560,N_3210,N_5830);
or U6561 (N_6561,N_3633,N_3400);
or U6562 (N_6562,N_5393,N_5241);
nor U6563 (N_6563,N_3666,N_4004);
nand U6564 (N_6564,N_4991,N_4125);
nor U6565 (N_6565,N_3293,N_5492);
nand U6566 (N_6566,N_5195,N_3626);
nor U6567 (N_6567,N_5245,N_4128);
nand U6568 (N_6568,N_4260,N_5555);
or U6569 (N_6569,N_3683,N_5174);
nor U6570 (N_6570,N_5801,N_3852);
nor U6571 (N_6571,N_4545,N_5964);
and U6572 (N_6572,N_4098,N_4198);
xor U6573 (N_6573,N_3163,N_3296);
nor U6574 (N_6574,N_3028,N_4446);
nor U6575 (N_6575,N_3609,N_5379);
and U6576 (N_6576,N_3051,N_5694);
and U6577 (N_6577,N_3248,N_5117);
and U6578 (N_6578,N_4707,N_4831);
and U6579 (N_6579,N_3119,N_5197);
or U6580 (N_6580,N_5151,N_5287);
or U6581 (N_6581,N_3815,N_3209);
or U6582 (N_6582,N_5221,N_5501);
or U6583 (N_6583,N_3995,N_5954);
nor U6584 (N_6584,N_5453,N_3052);
and U6585 (N_6585,N_5272,N_5111);
nand U6586 (N_6586,N_5766,N_4858);
nand U6587 (N_6587,N_3455,N_5746);
or U6588 (N_6588,N_5726,N_3444);
nor U6589 (N_6589,N_3767,N_3581);
or U6590 (N_6590,N_4632,N_3549);
nand U6591 (N_6591,N_5275,N_3488);
and U6592 (N_6592,N_4433,N_5737);
and U6593 (N_6593,N_4416,N_5587);
nand U6594 (N_6594,N_4975,N_4369);
and U6595 (N_6595,N_4017,N_4169);
or U6596 (N_6596,N_5112,N_4083);
or U6597 (N_6597,N_5824,N_3703);
nor U6598 (N_6598,N_4337,N_4581);
or U6599 (N_6599,N_4053,N_3368);
or U6600 (N_6600,N_5542,N_3607);
or U6601 (N_6601,N_3756,N_4764);
or U6602 (N_6602,N_5184,N_4551);
and U6603 (N_6603,N_4909,N_5914);
nor U6604 (N_6604,N_4346,N_4015);
and U6605 (N_6605,N_5740,N_4526);
and U6606 (N_6606,N_4475,N_4894);
nor U6607 (N_6607,N_5866,N_4844);
and U6608 (N_6608,N_5503,N_5090);
and U6609 (N_6609,N_4235,N_3094);
nor U6610 (N_6610,N_3737,N_3660);
or U6611 (N_6611,N_5248,N_5910);
or U6612 (N_6612,N_5085,N_5571);
nand U6613 (N_6613,N_5351,N_3776);
nor U6614 (N_6614,N_5715,N_3784);
and U6615 (N_6615,N_3800,N_4131);
nor U6616 (N_6616,N_5947,N_5369);
or U6617 (N_6617,N_5170,N_5841);
or U6618 (N_6618,N_5890,N_4672);
and U6619 (N_6619,N_5591,N_5626);
nand U6620 (N_6620,N_4069,N_3147);
nor U6621 (N_6621,N_5569,N_4107);
nor U6622 (N_6622,N_3329,N_4881);
or U6623 (N_6623,N_4834,N_5800);
or U6624 (N_6624,N_5097,N_5018);
nand U6625 (N_6625,N_5047,N_5764);
and U6626 (N_6626,N_4005,N_5779);
nand U6627 (N_6627,N_5274,N_3217);
and U6628 (N_6628,N_5076,N_3559);
nor U6629 (N_6629,N_5327,N_4724);
and U6630 (N_6630,N_5988,N_5312);
nand U6631 (N_6631,N_5416,N_5898);
or U6632 (N_6632,N_5573,N_4265);
nand U6633 (N_6633,N_5702,N_5234);
nor U6634 (N_6634,N_4391,N_5984);
nor U6635 (N_6635,N_5246,N_5086);
nand U6636 (N_6636,N_5589,N_3149);
or U6637 (N_6637,N_5781,N_4074);
nand U6638 (N_6638,N_5375,N_4527);
and U6639 (N_6639,N_5537,N_4151);
or U6640 (N_6640,N_3254,N_4488);
nor U6641 (N_6641,N_3527,N_4790);
or U6642 (N_6642,N_4325,N_5188);
nor U6643 (N_6643,N_3268,N_5929);
nand U6644 (N_6644,N_5295,N_4626);
or U6645 (N_6645,N_5209,N_5862);
nor U6646 (N_6646,N_4568,N_3206);
nor U6647 (N_6647,N_4832,N_4008);
or U6648 (N_6648,N_3680,N_4212);
or U6649 (N_6649,N_5744,N_5787);
nand U6650 (N_6650,N_5971,N_4252);
nor U6651 (N_6651,N_4410,N_4313);
nand U6652 (N_6652,N_5711,N_4097);
and U6653 (N_6653,N_4194,N_4032);
nor U6654 (N_6654,N_3428,N_5080);
nand U6655 (N_6655,N_3324,N_5939);
or U6656 (N_6656,N_5568,N_3441);
or U6657 (N_6657,N_4586,N_3785);
and U6658 (N_6658,N_5396,N_3372);
and U6659 (N_6659,N_3758,N_5469);
nand U6660 (N_6660,N_3027,N_5804);
and U6661 (N_6661,N_3524,N_3557);
or U6662 (N_6662,N_5418,N_5079);
or U6663 (N_6663,N_4811,N_3854);
nor U6664 (N_6664,N_5931,N_4088);
and U6665 (N_6665,N_4826,N_3820);
or U6666 (N_6666,N_4284,N_5915);
and U6667 (N_6667,N_5552,N_5687);
or U6668 (N_6668,N_5382,N_3969);
nand U6669 (N_6669,N_4787,N_4695);
nand U6670 (N_6670,N_4014,N_5439);
or U6671 (N_6671,N_3552,N_3851);
or U6672 (N_6672,N_3233,N_3868);
or U6673 (N_6673,N_3084,N_5466);
and U6674 (N_6674,N_4381,N_4282);
nor U6675 (N_6675,N_4269,N_4708);
or U6676 (N_6676,N_4563,N_5945);
and U6677 (N_6677,N_5354,N_3405);
and U6678 (N_6678,N_5825,N_4741);
and U6679 (N_6679,N_4690,N_4548);
nor U6680 (N_6680,N_5409,N_5619);
and U6681 (N_6681,N_4057,N_5998);
and U6682 (N_6682,N_5060,N_3091);
nor U6683 (N_6683,N_3970,N_5210);
nand U6684 (N_6684,N_4591,N_4351);
and U6685 (N_6685,N_3370,N_3742);
or U6686 (N_6686,N_5350,N_5014);
and U6687 (N_6687,N_4390,N_4352);
xnor U6688 (N_6688,N_5254,N_3641);
nor U6689 (N_6689,N_3208,N_3176);
or U6690 (N_6690,N_5114,N_3297);
nand U6691 (N_6691,N_3224,N_3049);
or U6692 (N_6692,N_3584,N_5417);
nor U6693 (N_6693,N_3672,N_3887);
or U6694 (N_6694,N_3090,N_3765);
nor U6695 (N_6695,N_4213,N_3532);
and U6696 (N_6696,N_3232,N_4232);
nor U6697 (N_6697,N_4768,N_3836);
nor U6698 (N_6698,N_5630,N_3059);
and U6699 (N_6699,N_5486,N_3170);
nand U6700 (N_6700,N_3536,N_3064);
or U6701 (N_6701,N_3347,N_5864);
nand U6702 (N_6702,N_5394,N_3349);
nand U6703 (N_6703,N_4207,N_4775);
and U6704 (N_6704,N_4949,N_3463);
or U6705 (N_6705,N_4955,N_5301);
nand U6706 (N_6706,N_4740,N_4959);
nor U6707 (N_6707,N_3192,N_3816);
nor U6708 (N_6708,N_3537,N_4540);
nand U6709 (N_6709,N_5560,N_3908);
and U6710 (N_6710,N_3320,N_3790);
nor U6711 (N_6711,N_5022,N_5343);
nor U6712 (N_6712,N_3827,N_5806);
nand U6713 (N_6713,N_3358,N_3981);
xor U6714 (N_6714,N_4999,N_5736);
nand U6715 (N_6715,N_5352,N_3332);
and U6716 (N_6716,N_3588,N_5811);
and U6717 (N_6717,N_3247,N_3069);
nand U6718 (N_6718,N_5969,N_4436);
or U6719 (N_6719,N_3437,N_5255);
xnor U6720 (N_6720,N_5078,N_5321);
nand U6721 (N_6721,N_5531,N_4671);
nor U6722 (N_6722,N_5427,N_4394);
nand U6723 (N_6723,N_5972,N_4003);
and U6724 (N_6724,N_3157,N_4038);
or U6725 (N_6725,N_3097,N_4735);
nor U6726 (N_6726,N_4721,N_5154);
nand U6727 (N_6727,N_3080,N_4307);
or U6728 (N_6728,N_3389,N_3316);
or U6729 (N_6729,N_4828,N_4440);
or U6730 (N_6730,N_3899,N_3279);
or U6731 (N_6731,N_4638,N_5433);
and U6732 (N_6732,N_4385,N_3579);
nand U6733 (N_6733,N_4887,N_4281);
and U6734 (N_6734,N_4593,N_3700);
and U6735 (N_6735,N_4669,N_4782);
nand U6736 (N_6736,N_4608,N_4464);
nand U6737 (N_6737,N_4997,N_3558);
nand U6738 (N_6738,N_3414,N_4954);
nand U6739 (N_6739,N_3117,N_4072);
nor U6740 (N_6740,N_4792,N_5661);
and U6741 (N_6741,N_3648,N_4100);
or U6742 (N_6742,N_3012,N_3345);
nand U6743 (N_6743,N_5750,N_3144);
and U6744 (N_6744,N_3775,N_4401);
and U6745 (N_6745,N_5705,N_5299);
or U6746 (N_6746,N_3948,N_4345);
nor U6747 (N_6747,N_5213,N_4980);
nor U6748 (N_6748,N_3230,N_4222);
nand U6749 (N_6749,N_3572,N_5518);
or U6750 (N_6750,N_4019,N_4904);
nand U6751 (N_6751,N_5309,N_3250);
nor U6752 (N_6752,N_3610,N_5460);
nor U6753 (N_6753,N_4134,N_3597);
nor U6754 (N_6754,N_5472,N_4677);
or U6755 (N_6755,N_5140,N_4989);
or U6756 (N_6756,N_3857,N_3682);
and U6757 (N_6757,N_5527,N_3357);
or U6758 (N_6758,N_3113,N_3843);
or U6759 (N_6759,N_4138,N_5010);
or U6760 (N_6760,N_3678,N_5159);
nor U6761 (N_6761,N_4820,N_5897);
and U6762 (N_6762,N_4679,N_3958);
nand U6763 (N_6763,N_3096,N_3363);
and U6764 (N_6764,N_4499,N_3694);
and U6765 (N_6765,N_5120,N_3070);
or U6766 (N_6766,N_4270,N_4309);
nand U6767 (N_6767,N_5489,N_5037);
nor U6768 (N_6768,N_3646,N_5364);
nor U6769 (N_6769,N_4791,N_3276);
and U6770 (N_6770,N_3366,N_5381);
nand U6771 (N_6771,N_3228,N_4817);
and U6772 (N_6772,N_3439,N_5494);
nand U6773 (N_6773,N_4228,N_3225);
and U6774 (N_6774,N_4179,N_3395);
or U6775 (N_6775,N_5794,N_3569);
nor U6776 (N_6776,N_5863,N_3010);
or U6777 (N_6777,N_4311,N_3373);
nor U6778 (N_6778,N_5385,N_3773);
nor U6779 (N_6779,N_3124,N_4353);
or U6780 (N_6780,N_3753,N_4536);
or U6781 (N_6781,N_3278,N_3778);
or U6782 (N_6782,N_3331,N_5649);
and U6783 (N_6783,N_5884,N_4292);
or U6784 (N_6784,N_5713,N_3743);
and U6785 (N_6785,N_5878,N_3593);
and U6786 (N_6786,N_3971,N_5228);
or U6787 (N_6787,N_4567,N_4504);
or U6788 (N_6788,N_5728,N_5782);
and U6789 (N_6789,N_5380,N_5033);
or U6790 (N_6790,N_3151,N_5408);
nor U6791 (N_6791,N_3865,N_4510);
or U6792 (N_6792,N_3169,N_3073);
and U6793 (N_6793,N_3284,N_4133);
and U6794 (N_6794,N_3803,N_5622);
nor U6795 (N_6795,N_3468,N_5595);
and U6796 (N_6796,N_4566,N_3904);
nor U6797 (N_6797,N_4633,N_5270);
nand U6798 (N_6798,N_5367,N_3312);
or U6799 (N_6799,N_3741,N_5082);
or U6800 (N_6800,N_4704,N_5132);
nor U6801 (N_6801,N_5373,N_4001);
nand U6802 (N_6802,N_3460,N_3723);
nor U6803 (N_6803,N_4434,N_3934);
nand U6804 (N_6804,N_5572,N_4678);
and U6805 (N_6805,N_5268,N_4788);
or U6806 (N_6806,N_5771,N_3942);
nor U6807 (N_6807,N_4356,N_3416);
or U6808 (N_6808,N_4139,N_4627);
and U6809 (N_6809,N_4000,N_3926);
nor U6810 (N_6810,N_5161,N_5735);
or U6811 (N_6811,N_5946,N_4208);
nand U6812 (N_6812,N_4319,N_4274);
or U6813 (N_6813,N_5372,N_3665);
or U6814 (N_6814,N_4929,N_3497);
nand U6815 (N_6815,N_5856,N_5845);
nand U6816 (N_6816,N_3214,N_4089);
or U6817 (N_6817,N_5285,N_5665);
or U6818 (N_6818,N_4728,N_3690);
nand U6819 (N_6819,N_5015,N_4520);
and U6820 (N_6820,N_5570,N_4387);
nand U6821 (N_6821,N_3879,N_5966);
nor U6822 (N_6822,N_4010,N_5247);
and U6823 (N_6823,N_4491,N_4180);
and U6824 (N_6824,N_4382,N_4869);
nor U6825 (N_6825,N_5578,N_4745);
and U6826 (N_6826,N_4686,N_5522);
and U6827 (N_6827,N_5468,N_4092);
and U6828 (N_6828,N_5917,N_4136);
nand U6829 (N_6829,N_3699,N_4603);
xor U6830 (N_6830,N_4132,N_5432);
nand U6831 (N_6831,N_5596,N_4853);
nand U6832 (N_6832,N_3306,N_5879);
nand U6833 (N_6833,N_4960,N_3654);
nor U6834 (N_6834,N_4719,N_4104);
and U6835 (N_6835,N_3401,N_5323);
and U6836 (N_6836,N_4639,N_4478);
or U6837 (N_6837,N_5458,N_3892);
and U6838 (N_6838,N_4759,N_5052);
nand U6839 (N_6839,N_3522,N_5217);
and U6840 (N_6840,N_4943,N_3057);
and U6841 (N_6841,N_5586,N_5730);
and U6842 (N_6842,N_3792,N_4629);
nand U6843 (N_6843,N_5977,N_4330);
or U6844 (N_6844,N_4075,N_3396);
and U6845 (N_6845,N_4209,N_5514);
or U6846 (N_6846,N_5107,N_3477);
nor U6847 (N_6847,N_4847,N_3160);
and U6848 (N_6848,N_5872,N_3369);
nand U6849 (N_6849,N_4617,N_4246);
nor U6850 (N_6850,N_3862,N_4495);
and U6851 (N_6851,N_3553,N_4952);
nor U6852 (N_6852,N_5359,N_4630);
nor U6853 (N_6853,N_5877,N_5819);
nor U6854 (N_6854,N_4976,N_3698);
nand U6855 (N_6855,N_4685,N_5152);
nand U6856 (N_6856,N_3041,N_3054);
nor U6857 (N_6857,N_5100,N_3947);
and U6858 (N_6858,N_4953,N_4314);
and U6859 (N_6859,N_3386,N_5240);
or U6860 (N_6860,N_4465,N_4786);
nor U6861 (N_6861,N_5437,N_5677);
nand U6862 (N_6862,N_3965,N_3311);
or U6863 (N_6863,N_3943,N_3005);
nor U6864 (N_6864,N_3042,N_3162);
nor U6865 (N_6865,N_5557,N_5371);
and U6866 (N_6866,N_5893,N_3615);
or U6867 (N_6867,N_5828,N_3718);
or U6868 (N_6868,N_3288,N_4020);
nand U6869 (N_6869,N_3082,N_3878);
nand U6870 (N_6870,N_4753,N_5786);
and U6871 (N_6871,N_3457,N_3237);
nor U6872 (N_6872,N_4444,N_5280);
or U6873 (N_6873,N_5009,N_3563);
nand U6874 (N_6874,N_5617,N_5822);
xnor U6875 (N_6875,N_3227,N_4783);
or U6876 (N_6876,N_3550,N_4940);
nor U6877 (N_6877,N_3079,N_5338);
nor U6878 (N_6878,N_4644,N_4744);
nand U6879 (N_6879,N_3750,N_3172);
nand U6880 (N_6880,N_4754,N_3475);
or U6881 (N_6881,N_5098,N_5698);
nand U6882 (N_6882,N_5827,N_4614);
nand U6883 (N_6883,N_5608,N_5706);
and U6884 (N_6884,N_5336,N_4765);
nor U6885 (N_6885,N_3891,N_4623);
and U6886 (N_6886,N_5224,N_4052);
nor U6887 (N_6887,N_5068,N_3779);
nor U6888 (N_6888,N_3146,N_4324);
or U6889 (N_6889,N_3309,N_4794);
and U6890 (N_6890,N_4068,N_5034);
and U6891 (N_6891,N_3825,N_3442);
nor U6892 (N_6892,N_3922,N_3628);
nor U6893 (N_6893,N_5126,N_3104);
or U6894 (N_6894,N_4011,N_4328);
and U6895 (N_6895,N_5957,N_3510);
or U6896 (N_6896,N_4266,N_4701);
or U6897 (N_6897,N_5124,N_3760);
and U6898 (N_6898,N_3953,N_4166);
and U6899 (N_6899,N_4964,N_3809);
or U6900 (N_6900,N_5853,N_3838);
nand U6901 (N_6901,N_4565,N_5304);
nand U6902 (N_6902,N_5948,N_5912);
and U6903 (N_6903,N_3182,N_4849);
or U6904 (N_6904,N_3762,N_3319);
nand U6905 (N_6905,N_3705,N_3226);
nand U6906 (N_6906,N_4435,N_4752);
nand U6907 (N_6907,N_5476,N_3131);
nor U6908 (N_6908,N_3945,N_4376);
nor U6909 (N_6909,N_5935,N_3008);
nor U6910 (N_6910,N_4968,N_4217);
and U6911 (N_6911,N_4726,N_4876);
or U6912 (N_6912,N_3193,N_4905);
nor U6913 (N_6913,N_5565,N_5243);
and U6914 (N_6914,N_4206,N_4722);
nor U6915 (N_6915,N_3986,N_3483);
or U6916 (N_6916,N_3061,N_3108);
or U6917 (N_6917,N_4878,N_3772);
and U6918 (N_6918,N_5631,N_3336);
nor U6919 (N_6919,N_3814,N_4417);
or U6920 (N_6920,N_4454,N_4022);
nand U6921 (N_6921,N_3454,N_5748);
nor U6922 (N_6922,N_4202,N_5865);
nand U6923 (N_6923,N_4995,N_3388);
nor U6924 (N_6924,N_5081,N_5495);
and U6925 (N_6925,N_3095,N_4883);
or U6926 (N_6926,N_3939,N_3920);
or U6927 (N_6927,N_4191,N_5347);
and U6928 (N_6928,N_5180,N_4117);
nand U6929 (N_6929,N_4378,N_4518);
nand U6930 (N_6930,N_4532,N_5547);
or U6931 (N_6931,N_3717,N_3287);
nand U6932 (N_6932,N_4110,N_5413);
nand U6933 (N_6933,N_4729,N_3472);
or U6934 (N_6934,N_5720,N_3199);
or U6935 (N_6935,N_3327,N_3876);
nor U6936 (N_6936,N_4114,N_5911);
xor U6937 (N_6937,N_4681,N_4845);
nor U6938 (N_6938,N_4715,N_4713);
and U6939 (N_6939,N_3326,N_3338);
nand U6940 (N_6940,N_3018,N_4225);
nand U6941 (N_6941,N_5465,N_4383);
nor U6942 (N_6942,N_5690,N_5237);
and U6943 (N_6943,N_5341,N_5035);
nand U6944 (N_6944,N_3793,N_3759);
nor U6945 (N_6945,N_4430,N_5749);
nand U6946 (N_6946,N_5727,N_5242);
or U6947 (N_6947,N_4711,N_5271);
nor U6948 (N_6948,N_4280,N_3305);
nand U6949 (N_6949,N_5857,N_3196);
and U6950 (N_6950,N_5615,N_3637);
nor U6951 (N_6951,N_4181,N_4184);
or U6952 (N_6952,N_4205,N_3175);
nor U6953 (N_6953,N_5192,N_3740);
and U6954 (N_6954,N_5448,N_3739);
nand U6955 (N_6955,N_4109,N_4317);
and U6956 (N_6956,N_4769,N_3668);
nor U6957 (N_6957,N_5218,N_5403);
nand U6958 (N_6958,N_5647,N_3420);
xnor U6959 (N_6959,N_3342,N_5291);
and U6960 (N_6960,N_5820,N_5069);
and U6961 (N_6961,N_4815,N_3030);
xnor U6962 (N_6962,N_5115,N_5002);
and U6963 (N_6963,N_4431,N_4350);
nand U6964 (N_6964,N_5284,N_5013);
nand U6965 (N_6965,N_3191,N_3721);
and U6966 (N_6966,N_3443,N_5040);
nor U6967 (N_6967,N_3861,N_5496);
nor U6968 (N_6968,N_5815,N_4822);
nor U6969 (N_6969,N_3746,N_4619);
nand U6970 (N_6970,N_4408,N_3932);
nor U6971 (N_6971,N_3806,N_4838);
nor U6972 (N_6972,N_5227,N_4247);
and U6973 (N_6973,N_4427,N_4659);
nor U6974 (N_6974,N_4470,N_4562);
and U6975 (N_6975,N_4374,N_3355);
nand U6976 (N_6976,N_5670,N_4426);
and U6977 (N_6977,N_5363,N_4537);
and U6978 (N_6978,N_5096,N_4561);
nand U6979 (N_6979,N_5259,N_4081);
and U6980 (N_6980,N_4944,N_3972);
nand U6981 (N_6981,N_5927,N_5109);
nand U6982 (N_6982,N_3474,N_3585);
nand U6983 (N_6983,N_5419,N_3726);
or U6984 (N_6984,N_5848,N_5049);
or U6985 (N_6985,N_4947,N_5110);
nor U6986 (N_6986,N_3662,N_3611);
nor U6987 (N_6987,N_5797,N_3931);
or U6988 (N_6988,N_5585,N_3521);
or U6989 (N_6989,N_5219,N_4778);
nor U6990 (N_6990,N_4668,N_4583);
nand U6991 (N_6991,N_3944,N_5676);
nor U6992 (N_6992,N_5837,N_4027);
and U6993 (N_6993,N_3629,N_3255);
and U6994 (N_6994,N_3044,N_3893);
nor U6995 (N_6995,N_3586,N_5545);
nor U6996 (N_6996,N_5921,N_5951);
nand U6997 (N_6997,N_5225,N_5025);
xnor U6998 (N_6998,N_3125,N_4871);
nor U6999 (N_6999,N_3013,N_5920);
nand U7000 (N_7000,N_4648,N_3517);
or U7001 (N_7001,N_5629,N_3642);
nand U7002 (N_7002,N_4018,N_4873);
xor U7003 (N_7003,N_4201,N_4585);
or U7004 (N_7004,N_5279,N_5289);
and U7005 (N_7005,N_4466,N_3936);
and U7006 (N_7006,N_3046,N_5814);
or U7007 (N_7007,N_4468,N_5355);
or U7008 (N_7008,N_3901,N_5263);
nand U7009 (N_7009,N_5026,N_3709);
nand U7010 (N_7010,N_3555,N_3352);
nand U7011 (N_7011,N_5981,N_5443);
nand U7012 (N_7012,N_3377,N_3433);
and U7013 (N_7013,N_5345,N_4710);
or U7014 (N_7014,N_3811,N_4544);
nor U7015 (N_7015,N_5874,N_4755);
or U7016 (N_7016,N_3424,N_3301);
and U7017 (N_7017,N_5628,N_4612);
nor U7018 (N_7018,N_5044,N_3713);
nand U7019 (N_7019,N_4271,N_5655);
or U7020 (N_7020,N_4956,N_5996);
and U7021 (N_7021,N_5639,N_5397);
or U7022 (N_7022,N_4647,N_3961);
nor U7023 (N_7023,N_5919,N_4998);
nor U7024 (N_7024,N_4172,N_3791);
and U7025 (N_7025,N_3514,N_5975);
nor U7026 (N_7026,N_3371,N_4631);
or U7027 (N_7027,N_5885,N_3286);
nor U7028 (N_7028,N_5634,N_4363);
or U7029 (N_7029,N_3554,N_5805);
nand U7030 (N_7030,N_5648,N_3826);
or U7031 (N_7031,N_5840,N_3689);
nand U7032 (N_7032,N_5775,N_4197);
and U7033 (N_7033,N_5153,N_5230);
nor U7034 (N_7034,N_3180,N_4295);
nand U7035 (N_7035,N_4803,N_3128);
nand U7036 (N_7036,N_3402,N_5502);
or U7037 (N_7037,N_3606,N_4147);
nor U7038 (N_7038,N_3987,N_4948);
nand U7039 (N_7039,N_5609,N_4680);
nor U7040 (N_7040,N_4148,N_3916);
nor U7041 (N_7041,N_4624,N_3764);
and U7042 (N_7042,N_4830,N_3181);
nor U7043 (N_7043,N_3777,N_5325);
and U7044 (N_7044,N_3770,N_4700);
nor U7045 (N_7045,N_3796,N_5191);
or U7046 (N_7046,N_3264,N_5386);
nor U7047 (N_7047,N_4994,N_5134);
nor U7048 (N_7048,N_4064,N_3909);
nand U7049 (N_7049,N_5829,N_3346);
nand U7050 (N_7050,N_3959,N_3599);
or U7051 (N_7051,N_5314,N_5131);
and U7052 (N_7052,N_5508,N_3300);
or U7053 (N_7053,N_3845,N_3991);
nor U7054 (N_7054,N_4663,N_3270);
or U7055 (N_7055,N_4115,N_3905);
and U7056 (N_7056,N_5870,N_3594);
nor U7057 (N_7057,N_3566,N_4705);
or U7058 (N_7058,N_3768,N_3658);
nor U7059 (N_7059,N_3101,N_3379);
and U7060 (N_7060,N_4712,N_4509);
and U7061 (N_7061,N_4651,N_5286);
nor U7062 (N_7062,N_4286,N_3751);
and U7063 (N_7063,N_5370,N_5983);
nand U7064 (N_7064,N_3078,N_3266);
and U7065 (N_7065,N_5790,N_4146);
and U7066 (N_7066,N_5642,N_3933);
or U7067 (N_7067,N_5504,N_4985);
nand U7068 (N_7068,N_3795,N_3390);
nor U7069 (N_7069,N_5322,N_5719);
nor U7070 (N_7070,N_5714,N_5701);
nand U7071 (N_7071,N_3614,N_4689);
and U7072 (N_7072,N_3754,N_4257);
and U7073 (N_7073,N_3982,N_3272);
nor U7074 (N_7074,N_3516,N_5861);
nand U7075 (N_7075,N_4301,N_4512);
and U7076 (N_7076,N_3489,N_4071);
or U7077 (N_7077,N_5599,N_5459);
nand U7078 (N_7078,N_4965,N_3020);
nand U7079 (N_7079,N_3186,N_3245);
xor U7080 (N_7080,N_5330,N_5407);
nor U7081 (N_7081,N_5624,N_3189);
and U7082 (N_7082,N_3847,N_4622);
and U7083 (N_7083,N_4699,N_3031);
and U7084 (N_7084,N_5293,N_4026);
nor U7085 (N_7085,N_5113,N_5091);
xor U7086 (N_7086,N_5742,N_5876);
and U7087 (N_7087,N_3675,N_4911);
and U7088 (N_7088,N_5491,N_5276);
and U7089 (N_7089,N_4958,N_3541);
nor U7090 (N_7090,N_3509,N_4255);
and U7091 (N_7091,N_4667,N_4649);
nor U7092 (N_7092,N_5839,N_3413);
and U7093 (N_7093,N_3608,N_4984);
and U7094 (N_7094,N_5193,N_5524);
nand U7095 (N_7095,N_5696,N_4472);
nor U7096 (N_7096,N_5036,N_4996);
nor U7097 (N_7097,N_5005,N_5020);
nor U7098 (N_7098,N_3261,N_4862);
nand U7099 (N_7099,N_4730,N_3716);
and U7100 (N_7100,N_3213,N_5645);
nor U7101 (N_7101,N_4413,N_3252);
nor U7102 (N_7102,N_3231,N_4294);
nand U7103 (N_7103,N_5703,N_4574);
and U7104 (N_7104,N_4034,N_3914);
nand U7105 (N_7105,N_4674,N_4113);
nand U7106 (N_7106,N_3556,N_4177);
nand U7107 (N_7107,N_4634,N_3492);
nor U7108 (N_7108,N_4161,N_5546);
and U7109 (N_7109,N_3856,N_4037);
nor U7110 (N_7110,N_5653,N_5106);
nor U7111 (N_7111,N_5543,N_4462);
nand U7112 (N_7112,N_5640,N_3919);
nand U7113 (N_7113,N_4497,N_3427);
or U7114 (N_7114,N_5473,N_5562);
nand U7115 (N_7115,N_5517,N_4823);
and U7116 (N_7116,N_3840,N_3158);
or U7117 (N_7117,N_3062,N_5899);
nor U7118 (N_7118,N_5451,N_3867);
or U7119 (N_7119,N_5761,N_5308);
and U7120 (N_7120,N_5796,N_4734);
nand U7121 (N_7121,N_5253,N_3014);
nor U7122 (N_7122,N_3432,N_3548);
nand U7123 (N_7123,N_4457,N_3380);
and U7124 (N_7124,N_5563,N_4093);
nand U7125 (N_7125,N_4793,N_3024);
and U7126 (N_7126,N_5452,N_4482);
and U7127 (N_7127,N_5930,N_4570);
nor U7128 (N_7128,N_3167,N_5389);
nor U7129 (N_7129,N_3631,N_5908);
and U7130 (N_7130,N_3040,N_5045);
or U7131 (N_7131,N_4171,N_3491);
or U7132 (N_7132,N_5993,N_4441);
nor U7133 (N_7133,N_5162,N_4538);
or U7134 (N_7134,N_4013,N_5918);
nand U7135 (N_7135,N_4380,N_4359);
or U7136 (N_7136,N_4988,N_4970);
and U7137 (N_7137,N_3446,N_5331);
nand U7138 (N_7138,N_5513,N_4977);
nand U7139 (N_7139,N_4620,N_3098);
or U7140 (N_7140,N_3979,N_3330);
or U7141 (N_7141,N_3988,N_4106);
or U7142 (N_7142,N_3574,N_3412);
and U7143 (N_7143,N_5222,N_4336);
nand U7144 (N_7144,N_5826,N_4762);
nor U7145 (N_7145,N_4635,N_4592);
or U7146 (N_7146,N_5119,N_4841);
nor U7147 (N_7147,N_4655,N_4903);
nor U7148 (N_7148,N_5215,N_4656);
and U7149 (N_7149,N_3212,N_3274);
nor U7150 (N_7150,N_3618,N_4331);
nand U7151 (N_7151,N_3499,N_5529);
nor U7152 (N_7152,N_4746,N_5784);
or U7153 (N_7153,N_3704,N_4459);
and U7154 (N_7154,N_4515,N_4076);
nor U7155 (N_7155,N_3500,N_5638);
nor U7156 (N_7156,N_5614,N_5751);
or U7157 (N_7157,N_5368,N_4652);
nand U7158 (N_7158,N_5135,N_5516);
nand U7159 (N_7159,N_4914,N_4885);
and U7160 (N_7160,N_4129,N_5785);
or U7161 (N_7161,N_3077,N_4471);
nor U7162 (N_7162,N_4168,N_3923);
nand U7163 (N_7163,N_4086,N_4576);
nand U7164 (N_7164,N_5412,N_4095);
or U7165 (N_7165,N_5593,N_5342);
and U7166 (N_7166,N_5601,N_3494);
and U7167 (N_7167,N_5127,N_3249);
or U7168 (N_7168,N_5762,N_5778);
and U7169 (N_7169,N_4556,N_4061);
and U7170 (N_7170,N_5681,N_5189);
nand U7171 (N_7171,N_4682,N_4338);
nand U7172 (N_7172,N_3407,N_4276);
nand U7173 (N_7173,N_4993,N_5937);
nand U7174 (N_7174,N_3258,N_5238);
nor U7175 (N_7175,N_3850,N_5577);
or U7176 (N_7176,N_5186,N_4445);
or U7177 (N_7177,N_4963,N_4870);
nor U7178 (N_7178,N_3639,N_3298);
nand U7179 (N_7179,N_3037,N_5699);
and U7180 (N_7180,N_3461,N_5590);
or U7181 (N_7181,N_4877,N_5216);
nand U7182 (N_7182,N_4264,N_5428);
and U7183 (N_7183,N_4262,N_4643);
nand U7184 (N_7184,N_3744,N_4918);
nor U7185 (N_7185,N_3962,N_5854);
or U7186 (N_7186,N_3038,N_4702);
nand U7187 (N_7187,N_4354,N_3321);
nand U7188 (N_7188,N_5442,N_3318);
nor U7189 (N_7189,N_5995,N_5604);
nor U7190 (N_7190,N_4827,N_3473);
or U7191 (N_7191,N_3976,N_4157);
nand U7192 (N_7192,N_3093,N_5889);
or U7193 (N_7193,N_4698,N_3409);
or U7194 (N_7194,N_4931,N_5012);
or U7195 (N_7195,N_5182,N_4248);
or U7196 (N_7196,N_3471,N_3263);
or U7197 (N_7197,N_5760,N_3822);
nor U7198 (N_7198,N_4084,N_4477);
nor U7199 (N_7199,N_5567,N_5031);
and U7200 (N_7200,N_4810,N_4494);
nand U7201 (N_7201,N_4554,N_4159);
nor U7202 (N_7202,N_5388,N_5303);
and U7203 (N_7203,N_3722,N_4806);
nor U7204 (N_7204,N_3674,N_3032);
nor U7205 (N_7205,N_4534,N_5688);
or U7206 (N_7206,N_4789,N_3410);
nand U7207 (N_7207,N_3530,N_3506);
nor U7208 (N_7208,N_5402,N_3392);
nor U7209 (N_7209,N_3763,N_4291);
nor U7210 (N_7210,N_5391,N_5474);
nor U7211 (N_7211,N_3399,N_5298);
nor U7212 (N_7212,N_4062,N_5541);
xor U7213 (N_7213,N_3168,N_3022);
nor U7214 (N_7214,N_4641,N_3482);
and U7215 (N_7215,N_3504,N_4961);
nor U7216 (N_7216,N_5340,N_5682);
nor U7217 (N_7217,N_5205,N_5208);
and U7218 (N_7218,N_4200,N_5173);
or U7219 (N_7219,N_5752,N_5958);
nand U7220 (N_7220,N_3589,N_3035);
nand U7221 (N_7221,N_4329,N_4604);
nor U7222 (N_7222,N_3870,N_3938);
nand U7223 (N_7223,N_3676,N_3235);
nand U7224 (N_7224,N_5384,N_4323);
or U7225 (N_7225,N_4085,N_3616);
or U7226 (N_7226,N_5410,N_5101);
nor U7227 (N_7227,N_4621,N_3229);
nor U7228 (N_7228,N_4795,N_5094);
nor U7229 (N_7229,N_4547,N_4486);
or U7230 (N_7230,N_5160,N_3661);
and U7231 (N_7231,N_4298,N_3519);
nand U7232 (N_7232,N_4121,N_4763);
or U7233 (N_7233,N_3204,N_5141);
nand U7234 (N_7234,N_5137,N_4485);
nor U7235 (N_7235,N_5949,N_4227);
nand U7236 (N_7236,N_5533,N_3171);
nand U7237 (N_7237,N_4460,N_4874);
or U7238 (N_7238,N_3956,N_4645);
and U7239 (N_7239,N_5103,N_4030);
nor U7240 (N_7240,N_5994,N_5464);
nand U7241 (N_7241,N_4234,N_3415);
nor U7242 (N_7242,N_4349,N_4600);
and U7243 (N_7243,N_3802,N_4962);
or U7244 (N_7244,N_4315,N_5584);
nand U7245 (N_7245,N_5535,N_4372);
nand U7246 (N_7246,N_4067,N_5756);
and U7247 (N_7247,N_5471,N_5105);
nor U7248 (N_7248,N_3562,N_3184);
and U7249 (N_7249,N_4863,N_3872);
or U7250 (N_7250,N_4653,N_5057);
and U7251 (N_7251,N_5092,N_5558);
nand U7252 (N_7252,N_3695,N_4320);
nand U7253 (N_7253,N_3580,N_5833);
nand U7254 (N_7254,N_4718,N_5266);
nand U7255 (N_7255,N_3955,N_4193);
and U7256 (N_7256,N_3935,N_5950);
and U7257 (N_7257,N_4400,N_3669);
nand U7258 (N_7258,N_5450,N_4800);
or U7259 (N_7259,N_3636,N_3911);
and U7260 (N_7260,N_4082,N_3925);
or U7261 (N_7261,N_3145,N_3859);
nand U7262 (N_7262,N_4521,N_4571);
xnor U7263 (N_7263,N_3508,N_5989);
nor U7264 (N_7264,N_4230,N_3912);
and U7265 (N_7265,N_4557,N_4889);
nand U7266 (N_7266,N_4864,N_4405);
or U7267 (N_7267,N_3535,N_4415);
or U7268 (N_7268,N_5904,N_5361);
nor U7269 (N_7269,N_5667,N_5855);
nor U7270 (N_7270,N_3308,N_5070);
or U7271 (N_7271,N_5658,N_4244);
nor U7272 (N_7272,N_3071,N_5788);
nor U7273 (N_7273,N_3853,N_3664);
and U7274 (N_7274,N_3819,N_4278);
and U7275 (N_7275,N_3622,N_4694);
nor U7276 (N_7276,N_5269,N_4120);
nor U7277 (N_7277,N_4691,N_5063);
and U7278 (N_7278,N_4386,N_4928);
and U7279 (N_7279,N_3828,N_4505);
or U7280 (N_7280,N_5328,N_4665);
nor U7281 (N_7281,N_4502,N_5024);
or U7282 (N_7282,N_3950,N_3112);
and U7283 (N_7283,N_4550,N_5128);
nor U7284 (N_7284,N_5802,N_3166);
and U7285 (N_7285,N_3299,N_4021);
and U7286 (N_7286,N_4035,N_4373);
nor U7287 (N_7287,N_3518,N_5754);
or U7288 (N_7288,N_5065,N_4135);
nand U7289 (N_7289,N_4263,N_4727);
or U7290 (N_7290,N_4483,N_3403);
or U7291 (N_7291,N_3277,N_4852);
and U7292 (N_7292,N_5758,N_3781);
and U7293 (N_7293,N_4605,N_5734);
nor U7294 (N_7294,N_4731,N_3980);
nor U7295 (N_7295,N_5064,N_4066);
nor U7296 (N_7296,N_3067,N_4335);
nand U7297 (N_7297,N_5836,N_3748);
nor U7298 (N_7298,N_4850,N_3783);
nand U7299 (N_7299,N_5660,N_3050);
and U7300 (N_7300,N_4402,N_3730);
nor U7301 (N_7301,N_4897,N_3812);
nand U7302 (N_7302,N_4188,N_3546);
nand U7303 (N_7303,N_3310,N_4950);
nand U7304 (N_7304,N_5199,N_5990);
nand U7305 (N_7305,N_4773,N_3419);
and U7306 (N_7306,N_3624,N_4048);
nor U7307 (N_7307,N_3505,N_4613);
and U7308 (N_7308,N_4054,N_3374);
and U7309 (N_7309,N_4774,N_5774);
and U7310 (N_7310,N_5032,N_3152);
and U7311 (N_7311,N_4256,N_4450);
nand U7312 (N_7312,N_3848,N_3156);
and U7313 (N_7313,N_3135,N_5554);
and U7314 (N_7314,N_4484,N_3659);
or U7315 (N_7315,N_4982,N_4582);
nor U7316 (N_7316,N_5616,N_3946);
or U7317 (N_7317,N_5447,N_3954);
or U7318 (N_7318,N_3183,N_5534);
or U7319 (N_7319,N_3484,N_5695);
xnor U7320 (N_7320,N_3123,N_4780);
and U7321 (N_7321,N_5725,N_4403);
or U7322 (N_7322,N_3540,N_4002);
nor U7323 (N_7323,N_4348,N_4692);
or U7324 (N_7324,N_3993,N_4907);
and U7325 (N_7325,N_5053,N_3072);
or U7326 (N_7326,N_4979,N_3323);
nor U7327 (N_7327,N_3289,N_3106);
nor U7328 (N_7328,N_4170,N_4587);
and U7329 (N_7329,N_3006,N_5290);
or U7330 (N_7330,N_5077,N_5539);
or U7331 (N_7331,N_5970,N_4023);
or U7332 (N_7332,N_3161,N_3378);
nand U7333 (N_7333,N_3512,N_5637);
or U7334 (N_7334,N_5813,N_4340);
or U7335 (N_7335,N_5300,N_3065);
nand U7336 (N_7336,N_4050,N_3421);
nand U7337 (N_7337,N_3652,N_3881);
nor U7338 (N_7338,N_4183,N_5011);
or U7339 (N_7339,N_4601,N_3063);
or U7340 (N_7340,N_5692,N_5226);
nor U7341 (N_7341,N_3761,N_3087);
and U7342 (N_7342,N_5768,N_4856);
nand U7343 (N_7343,N_3178,N_4452);
and U7344 (N_7344,N_4941,N_4529);
nor U7345 (N_7345,N_4919,N_4846);
nor U7346 (N_7346,N_3259,N_5000);
nor U7347 (N_7347,N_3651,N_5583);
nand U7348 (N_7348,N_4816,N_3833);
nand U7349 (N_7349,N_5039,N_3429);
or U7350 (N_7350,N_3749,N_5883);
and U7351 (N_7351,N_4986,N_5399);
and U7352 (N_7352,N_3431,N_5809);
nor U7353 (N_7353,N_4321,N_3058);
or U7354 (N_7354,N_4553,N_3486);
and U7355 (N_7355,N_4615,N_4714);
and U7356 (N_7356,N_4467,N_5200);
nor U7357 (N_7357,N_3903,N_4103);
nor U7358 (N_7358,N_4195,N_3884);
nor U7359 (N_7359,N_3362,N_5099);
nand U7360 (N_7360,N_5406,N_5187);
nor U7361 (N_7361,N_5139,N_3215);
and U7362 (N_7362,N_3728,N_5974);
or U7363 (N_7363,N_5377,N_5512);
or U7364 (N_7364,N_3630,N_3602);
nor U7365 (N_7365,N_5657,N_4966);
and U7366 (N_7366,N_5519,N_4743);
nor U7367 (N_7367,N_3280,N_5007);
nand U7368 (N_7368,N_5627,N_3534);
or U7369 (N_7369,N_4673,N_3195);
nor U7370 (N_7370,N_3799,N_4818);
or U7371 (N_7371,N_5333,N_4798);
and U7372 (N_7372,N_3786,N_3671);
and U7373 (N_7373,N_5707,N_5952);
nor U7374 (N_7374,N_4123,N_5150);
nor U7375 (N_7375,N_4199,N_5992);
nor U7376 (N_7376,N_3620,N_4859);
nand U7377 (N_7377,N_4469,N_4388);
or U7378 (N_7378,N_5525,N_5938);
nand U7379 (N_7379,N_3673,N_3571);
and U7380 (N_7380,N_4211,N_5306);
nor U7381 (N_7381,N_3523,N_3808);
or U7382 (N_7382,N_3496,N_4835);
or U7383 (N_7383,N_5903,N_3281);
nand U7384 (N_7384,N_5816,N_5600);
and U7385 (N_7385,N_4422,N_3774);
or U7386 (N_7386,N_3706,N_4442);
nand U7387 (N_7387,N_4163,N_3907);
nand U7388 (N_7388,N_3203,N_4737);
nor U7389 (N_7389,N_4480,N_3335);
or U7390 (N_7390,N_3686,N_5446);
and U7391 (N_7391,N_5733,N_4080);
and U7392 (N_7392,N_3173,N_3127);
nor U7393 (N_7393,N_5483,N_5358);
and U7394 (N_7394,N_3725,N_5277);
nor U7395 (N_7395,N_4293,N_4162);
nor U7396 (N_7396,N_3142,N_5348);
and U7397 (N_7397,N_3964,N_5770);
and U7398 (N_7398,N_4364,N_5177);
or U7399 (N_7399,N_5429,N_4676);
nor U7400 (N_7400,N_4254,N_5400);
or U7401 (N_7401,N_3241,N_4607);
or U7402 (N_7402,N_5256,N_4912);
and U7403 (N_7403,N_3498,N_5691);
nand U7404 (N_7404,N_3478,N_3011);
and U7405 (N_7405,N_4983,N_4333);
nand U7406 (N_7406,N_5747,N_5924);
nand U7407 (N_7407,N_3350,N_4946);
nor U7408 (N_7408,N_3126,N_4552);
and U7409 (N_7409,N_3256,N_5122);
nor U7410 (N_7410,N_5307,N_4119);
nand U7411 (N_7411,N_3165,N_4118);
nor U7412 (N_7412,N_5422,N_5755);
and U7413 (N_7413,N_4902,N_4925);
and U7414 (N_7414,N_3873,N_4725);
and U7415 (N_7415,N_4804,N_3343);
nor U7416 (N_7416,N_5875,N_3179);
nand U7417 (N_7417,N_4910,N_4463);
nand U7418 (N_7418,N_4978,N_3863);
nand U7419 (N_7419,N_4779,N_5867);
nor U7420 (N_7420,N_4915,N_3650);
nor U7421 (N_7421,N_5799,N_5858);
nor U7422 (N_7422,N_3900,N_5605);
xor U7423 (N_7423,N_5073,N_4866);
or U7424 (N_7424,N_5485,N_4302);
and U7425 (N_7425,N_5181,N_4598);
or U7426 (N_7426,N_4145,N_3340);
nor U7427 (N_7427,N_5365,N_3001);
and U7428 (N_7428,N_3302,N_5704);
and U7429 (N_7429,N_3426,N_3068);
nand U7430 (N_7430,N_5261,N_5470);
nor U7431 (N_7431,N_4809,N_4428);
nor U7432 (N_7432,N_4154,N_5810);
nand U7433 (N_7433,N_3657,N_5506);
and U7434 (N_7434,N_5283,N_3910);
or U7435 (N_7435,N_3567,N_3984);
and U7436 (N_7436,N_3782,N_3906);
nand U7437 (N_7437,N_4610,N_4099);
nor U7438 (N_7438,N_4808,N_5038);
nor U7439 (N_7439,N_3844,N_5678);
and U7440 (N_7440,N_4150,N_4942);
and U7441 (N_7441,N_4108,N_4492);
nand U7442 (N_7442,N_3951,N_4751);
nor U7443 (N_7443,N_5956,N_5262);
nand U7444 (N_7444,N_3583,N_4951);
nor U7445 (N_7445,N_3114,N_4111);
nor U7446 (N_7446,N_5886,N_4709);
and U7447 (N_7447,N_5656,N_4501);
or U7448 (N_7448,N_4216,N_3140);
nand U7449 (N_7449,N_5894,N_4429);
and U7450 (N_7450,N_4748,N_3513);
or U7451 (N_7451,N_5976,N_4221);
or U7452 (N_7452,N_4640,N_5505);
nand U7453 (N_7453,N_3533,N_5850);
or U7454 (N_7454,N_5895,N_5423);
nand U7455 (N_7455,N_4153,N_3314);
nor U7456 (N_7456,N_4251,N_4549);
and U7457 (N_7457,N_3941,N_4127);
nor U7458 (N_7458,N_4596,N_3367);
nand U7459 (N_7459,N_3111,N_3143);
or U7460 (N_7460,N_5093,N_5909);
nor U7461 (N_7461,N_4055,N_3684);
nand U7462 (N_7462,N_3187,N_3036);
nor U7463 (N_7463,N_4898,N_4757);
nor U7464 (N_7464,N_4439,N_3771);
and U7465 (N_7465,N_4825,N_4843);
nand U7466 (N_7466,N_5481,N_3476);
nand U7467 (N_7467,N_5509,N_3685);
nor U7468 (N_7468,N_3866,N_4142);
or U7469 (N_7469,N_4805,N_5668);
nor U7470 (N_7470,N_4530,N_4130);
nor U7471 (N_7471,N_3573,N_4927);
and U7472 (N_7472,N_4840,N_3207);
and U7473 (N_7473,N_5739,N_3963);
or U7474 (N_7474,N_4384,N_3055);
or U7475 (N_7475,N_4516,N_4523);
or U7476 (N_7476,N_3325,N_3890);
nand U7477 (N_7477,N_5686,N_5709);
and U7478 (N_7478,N_4303,N_4611);
nand U7479 (N_7479,N_4539,N_4237);
and U7480 (N_7480,N_5666,N_4461);
nand U7481 (N_7481,N_4396,N_3086);
and U7482 (N_7482,N_5398,N_3531);
nand U7483 (N_7483,N_5559,N_3422);
nand U7484 (N_7484,N_3570,N_5679);
nand U7485 (N_7485,N_5179,N_5526);
and U7486 (N_7486,N_3769,N_5462);
nand U7487 (N_7487,N_4042,N_3677);
and U7488 (N_7488,N_3185,N_4522);
nor U7489 (N_7489,N_5743,N_3612);
or U7490 (N_7490,N_3480,N_5196);
nor U7491 (N_7491,N_4079,N_4696);
nand U7492 (N_7492,N_3545,N_5324);
and U7493 (N_7493,N_5265,N_4487);
nand U7494 (N_7494,N_3418,N_4421);
and U7495 (N_7495,N_5933,N_3952);
nand U7496 (N_7496,N_3973,N_4285);
nor U7497 (N_7497,N_4407,N_5710);
or U7498 (N_7498,N_4049,N_4182);
and U7499 (N_7499,N_4173,N_5618);
or U7500 (N_7500,N_5295,N_4423);
nand U7501 (N_7501,N_3410,N_4806);
and U7502 (N_7502,N_5667,N_5164);
or U7503 (N_7503,N_5702,N_4561);
nor U7504 (N_7504,N_3090,N_5708);
and U7505 (N_7505,N_3090,N_4661);
nor U7506 (N_7506,N_5340,N_3611);
nand U7507 (N_7507,N_4306,N_3180);
nand U7508 (N_7508,N_4272,N_3586);
nor U7509 (N_7509,N_3738,N_3888);
and U7510 (N_7510,N_4239,N_4765);
nor U7511 (N_7511,N_4637,N_3928);
nand U7512 (N_7512,N_4090,N_5934);
nand U7513 (N_7513,N_5772,N_4027);
or U7514 (N_7514,N_3961,N_4852);
and U7515 (N_7515,N_5567,N_3571);
and U7516 (N_7516,N_4152,N_3250);
and U7517 (N_7517,N_4005,N_4625);
or U7518 (N_7518,N_4671,N_4340);
and U7519 (N_7519,N_4663,N_5250);
nor U7520 (N_7520,N_4745,N_4432);
nand U7521 (N_7521,N_3307,N_5224);
or U7522 (N_7522,N_3751,N_5272);
nand U7523 (N_7523,N_5465,N_3898);
nand U7524 (N_7524,N_4538,N_5817);
nor U7525 (N_7525,N_3953,N_5975);
nand U7526 (N_7526,N_4147,N_5387);
or U7527 (N_7527,N_5500,N_3925);
nand U7528 (N_7528,N_5468,N_4775);
or U7529 (N_7529,N_4968,N_3151);
or U7530 (N_7530,N_5687,N_3740);
nor U7531 (N_7531,N_4241,N_3515);
and U7532 (N_7532,N_4832,N_4686);
and U7533 (N_7533,N_5407,N_5283);
nor U7534 (N_7534,N_3871,N_5688);
nor U7535 (N_7535,N_3097,N_5904);
xnor U7536 (N_7536,N_5974,N_4179);
or U7537 (N_7537,N_3778,N_5340);
nand U7538 (N_7538,N_3676,N_5669);
nor U7539 (N_7539,N_3464,N_5171);
nand U7540 (N_7540,N_3482,N_3935);
and U7541 (N_7541,N_5042,N_5639);
and U7542 (N_7542,N_3126,N_4806);
nand U7543 (N_7543,N_5679,N_5865);
and U7544 (N_7544,N_5868,N_5613);
xnor U7545 (N_7545,N_5642,N_4340);
or U7546 (N_7546,N_4125,N_3199);
nor U7547 (N_7547,N_4434,N_4589);
nor U7548 (N_7548,N_5051,N_3181);
nand U7549 (N_7549,N_5483,N_3043);
nand U7550 (N_7550,N_4441,N_4889);
or U7551 (N_7551,N_3490,N_5402);
and U7552 (N_7552,N_5029,N_3982);
nor U7553 (N_7553,N_4217,N_3702);
nand U7554 (N_7554,N_4957,N_5447);
nor U7555 (N_7555,N_4108,N_4535);
or U7556 (N_7556,N_5547,N_5430);
nor U7557 (N_7557,N_4898,N_3296);
nor U7558 (N_7558,N_3724,N_4181);
or U7559 (N_7559,N_5742,N_4976);
nor U7560 (N_7560,N_4999,N_5477);
nor U7561 (N_7561,N_4976,N_3961);
nor U7562 (N_7562,N_5037,N_4183);
and U7563 (N_7563,N_3959,N_4704);
nand U7564 (N_7564,N_3871,N_5444);
or U7565 (N_7565,N_4382,N_5636);
and U7566 (N_7566,N_5391,N_4916);
nand U7567 (N_7567,N_4536,N_3462);
or U7568 (N_7568,N_5192,N_5187);
or U7569 (N_7569,N_3953,N_4870);
or U7570 (N_7570,N_4539,N_3119);
nor U7571 (N_7571,N_4161,N_3273);
nand U7572 (N_7572,N_3986,N_5546);
nand U7573 (N_7573,N_4121,N_5665);
nand U7574 (N_7574,N_5621,N_5774);
or U7575 (N_7575,N_3123,N_5662);
xor U7576 (N_7576,N_4109,N_3322);
nand U7577 (N_7577,N_5679,N_5701);
nand U7578 (N_7578,N_3493,N_5064);
and U7579 (N_7579,N_3374,N_3627);
or U7580 (N_7580,N_5377,N_3921);
nand U7581 (N_7581,N_5684,N_5340);
or U7582 (N_7582,N_3102,N_3416);
and U7583 (N_7583,N_5709,N_4542);
and U7584 (N_7584,N_3371,N_4261);
nor U7585 (N_7585,N_3410,N_5311);
nand U7586 (N_7586,N_5938,N_5577);
nand U7587 (N_7587,N_4225,N_3296);
and U7588 (N_7588,N_5014,N_5579);
nand U7589 (N_7589,N_5900,N_4102);
or U7590 (N_7590,N_3633,N_4682);
and U7591 (N_7591,N_5999,N_4535);
and U7592 (N_7592,N_5427,N_5094);
nand U7593 (N_7593,N_4051,N_4196);
nor U7594 (N_7594,N_3036,N_4341);
and U7595 (N_7595,N_5727,N_5259);
nor U7596 (N_7596,N_5154,N_3003);
nor U7597 (N_7597,N_4293,N_3092);
or U7598 (N_7598,N_3964,N_3769);
and U7599 (N_7599,N_5020,N_3425);
nand U7600 (N_7600,N_5719,N_3102);
and U7601 (N_7601,N_4627,N_4145);
nand U7602 (N_7602,N_3627,N_3144);
nor U7603 (N_7603,N_3008,N_5609);
nor U7604 (N_7604,N_5022,N_5607);
nand U7605 (N_7605,N_4272,N_3150);
nor U7606 (N_7606,N_5410,N_3929);
nor U7607 (N_7607,N_3317,N_3827);
or U7608 (N_7608,N_3749,N_4820);
nor U7609 (N_7609,N_4853,N_4609);
and U7610 (N_7610,N_3108,N_5184);
nand U7611 (N_7611,N_4201,N_5082);
or U7612 (N_7612,N_4548,N_3229);
or U7613 (N_7613,N_5435,N_5340);
and U7614 (N_7614,N_5305,N_3313);
and U7615 (N_7615,N_3661,N_4523);
or U7616 (N_7616,N_4148,N_3352);
or U7617 (N_7617,N_3002,N_3757);
or U7618 (N_7618,N_4056,N_5330);
nor U7619 (N_7619,N_4873,N_3214);
nand U7620 (N_7620,N_3164,N_4520);
and U7621 (N_7621,N_3534,N_5116);
and U7622 (N_7622,N_3714,N_3487);
nor U7623 (N_7623,N_4015,N_4485);
nand U7624 (N_7624,N_4672,N_3291);
nand U7625 (N_7625,N_5758,N_4309);
or U7626 (N_7626,N_4889,N_5367);
nand U7627 (N_7627,N_4674,N_3601);
nand U7628 (N_7628,N_3971,N_3593);
nor U7629 (N_7629,N_5189,N_5067);
or U7630 (N_7630,N_5742,N_3187);
or U7631 (N_7631,N_4295,N_3540);
nor U7632 (N_7632,N_4151,N_3397);
and U7633 (N_7633,N_5869,N_3320);
and U7634 (N_7634,N_3032,N_3806);
nand U7635 (N_7635,N_4486,N_5276);
nand U7636 (N_7636,N_5518,N_4477);
nor U7637 (N_7637,N_4032,N_3459);
nor U7638 (N_7638,N_4550,N_4148);
and U7639 (N_7639,N_4650,N_4093);
nor U7640 (N_7640,N_3463,N_4370);
nand U7641 (N_7641,N_4545,N_5179);
or U7642 (N_7642,N_4332,N_3479);
or U7643 (N_7643,N_3615,N_3693);
nor U7644 (N_7644,N_3396,N_4352);
nor U7645 (N_7645,N_4934,N_4662);
nand U7646 (N_7646,N_4332,N_3478);
or U7647 (N_7647,N_3699,N_5775);
nand U7648 (N_7648,N_5510,N_5444);
nor U7649 (N_7649,N_3481,N_4212);
nor U7650 (N_7650,N_3654,N_4912);
and U7651 (N_7651,N_5910,N_5376);
nor U7652 (N_7652,N_4118,N_3190);
or U7653 (N_7653,N_4187,N_3426);
nor U7654 (N_7654,N_5159,N_3894);
and U7655 (N_7655,N_4976,N_3769);
nor U7656 (N_7656,N_3237,N_5179);
nand U7657 (N_7657,N_5611,N_5998);
nand U7658 (N_7658,N_5848,N_4910);
and U7659 (N_7659,N_5217,N_3808);
nor U7660 (N_7660,N_3945,N_4630);
nor U7661 (N_7661,N_5712,N_3322);
nand U7662 (N_7662,N_5040,N_4186);
nand U7663 (N_7663,N_3300,N_4150);
nand U7664 (N_7664,N_5110,N_4423);
nand U7665 (N_7665,N_3354,N_4565);
or U7666 (N_7666,N_5724,N_3506);
nand U7667 (N_7667,N_5140,N_4487);
nor U7668 (N_7668,N_4753,N_5189);
or U7669 (N_7669,N_4234,N_4670);
nand U7670 (N_7670,N_3153,N_3376);
nand U7671 (N_7671,N_4526,N_4811);
or U7672 (N_7672,N_5512,N_4633);
and U7673 (N_7673,N_3403,N_5358);
nor U7674 (N_7674,N_3136,N_4325);
or U7675 (N_7675,N_5018,N_5323);
or U7676 (N_7676,N_3213,N_5101);
nor U7677 (N_7677,N_3745,N_3749);
nor U7678 (N_7678,N_4619,N_3302);
or U7679 (N_7679,N_3378,N_4765);
nor U7680 (N_7680,N_5584,N_3462);
nand U7681 (N_7681,N_4686,N_3790);
and U7682 (N_7682,N_3350,N_4227);
nand U7683 (N_7683,N_4996,N_3625);
or U7684 (N_7684,N_3620,N_4839);
nor U7685 (N_7685,N_5249,N_3816);
nand U7686 (N_7686,N_5318,N_4748);
nand U7687 (N_7687,N_4296,N_5451);
nor U7688 (N_7688,N_3553,N_5507);
and U7689 (N_7689,N_3409,N_4763);
or U7690 (N_7690,N_5703,N_3244);
or U7691 (N_7691,N_3452,N_5391);
or U7692 (N_7692,N_4404,N_5492);
nor U7693 (N_7693,N_5134,N_5768);
nand U7694 (N_7694,N_4137,N_3919);
nor U7695 (N_7695,N_3685,N_3285);
or U7696 (N_7696,N_3585,N_5796);
nand U7697 (N_7697,N_3688,N_5759);
or U7698 (N_7698,N_4435,N_3922);
or U7699 (N_7699,N_3106,N_5288);
and U7700 (N_7700,N_3816,N_4160);
or U7701 (N_7701,N_3420,N_5594);
xnor U7702 (N_7702,N_3845,N_3123);
nor U7703 (N_7703,N_4863,N_4176);
nand U7704 (N_7704,N_4173,N_5306);
nor U7705 (N_7705,N_5451,N_3052);
or U7706 (N_7706,N_3579,N_4597);
nand U7707 (N_7707,N_3160,N_5796);
or U7708 (N_7708,N_3523,N_5062);
nor U7709 (N_7709,N_4427,N_4789);
nor U7710 (N_7710,N_3297,N_3387);
or U7711 (N_7711,N_5377,N_5535);
and U7712 (N_7712,N_5883,N_4273);
and U7713 (N_7713,N_3623,N_5532);
nor U7714 (N_7714,N_4553,N_3029);
nor U7715 (N_7715,N_5382,N_5638);
nand U7716 (N_7716,N_3479,N_3160);
and U7717 (N_7717,N_4890,N_4994);
nor U7718 (N_7718,N_4330,N_5882);
and U7719 (N_7719,N_5996,N_4180);
nand U7720 (N_7720,N_3543,N_4652);
and U7721 (N_7721,N_4896,N_5371);
or U7722 (N_7722,N_5288,N_3207);
nor U7723 (N_7723,N_5197,N_5133);
nand U7724 (N_7724,N_3517,N_5129);
or U7725 (N_7725,N_3881,N_4226);
nor U7726 (N_7726,N_4009,N_5660);
or U7727 (N_7727,N_5472,N_3733);
or U7728 (N_7728,N_4831,N_3015);
nor U7729 (N_7729,N_4959,N_5353);
nand U7730 (N_7730,N_5832,N_3116);
nor U7731 (N_7731,N_5799,N_4027);
or U7732 (N_7732,N_5899,N_3242);
nand U7733 (N_7733,N_3880,N_3315);
nand U7734 (N_7734,N_5336,N_3804);
or U7735 (N_7735,N_5869,N_4273);
nor U7736 (N_7736,N_5065,N_4863);
or U7737 (N_7737,N_4673,N_5233);
nand U7738 (N_7738,N_3165,N_4384);
and U7739 (N_7739,N_3663,N_3590);
nand U7740 (N_7740,N_3491,N_4638);
nor U7741 (N_7741,N_4146,N_4684);
and U7742 (N_7742,N_4800,N_3016);
nor U7743 (N_7743,N_4541,N_4356);
and U7744 (N_7744,N_3016,N_3010);
nand U7745 (N_7745,N_4316,N_4781);
nand U7746 (N_7746,N_5243,N_5203);
or U7747 (N_7747,N_3106,N_4149);
or U7748 (N_7748,N_5151,N_4644);
and U7749 (N_7749,N_3663,N_4673);
nand U7750 (N_7750,N_4372,N_5312);
or U7751 (N_7751,N_4579,N_4881);
and U7752 (N_7752,N_3233,N_5358);
nor U7753 (N_7753,N_4491,N_3601);
nor U7754 (N_7754,N_5513,N_3989);
or U7755 (N_7755,N_5989,N_5844);
and U7756 (N_7756,N_3329,N_3497);
and U7757 (N_7757,N_4560,N_3230);
nand U7758 (N_7758,N_3610,N_5840);
or U7759 (N_7759,N_5640,N_5019);
nand U7760 (N_7760,N_3380,N_4246);
nand U7761 (N_7761,N_4237,N_4544);
and U7762 (N_7762,N_5132,N_4560);
or U7763 (N_7763,N_3433,N_3238);
and U7764 (N_7764,N_5547,N_5494);
nor U7765 (N_7765,N_4410,N_3555);
nand U7766 (N_7766,N_5731,N_4983);
and U7767 (N_7767,N_3515,N_5130);
nor U7768 (N_7768,N_4433,N_4973);
and U7769 (N_7769,N_5109,N_5850);
nand U7770 (N_7770,N_4534,N_4561);
nor U7771 (N_7771,N_5115,N_5327);
nand U7772 (N_7772,N_3444,N_3150);
or U7773 (N_7773,N_4544,N_3222);
and U7774 (N_7774,N_3661,N_4391);
nand U7775 (N_7775,N_3014,N_4395);
and U7776 (N_7776,N_3999,N_5482);
nand U7777 (N_7777,N_4117,N_3553);
and U7778 (N_7778,N_5587,N_4776);
nor U7779 (N_7779,N_5098,N_5136);
and U7780 (N_7780,N_4342,N_5292);
nand U7781 (N_7781,N_3650,N_4948);
or U7782 (N_7782,N_5968,N_5719);
and U7783 (N_7783,N_3190,N_5128);
nand U7784 (N_7784,N_4921,N_5968);
xnor U7785 (N_7785,N_5998,N_4205);
nor U7786 (N_7786,N_3246,N_5425);
or U7787 (N_7787,N_3188,N_4474);
and U7788 (N_7788,N_4763,N_4641);
or U7789 (N_7789,N_5171,N_4750);
or U7790 (N_7790,N_5936,N_3760);
or U7791 (N_7791,N_4353,N_3746);
nor U7792 (N_7792,N_5319,N_3928);
nor U7793 (N_7793,N_3033,N_5197);
nor U7794 (N_7794,N_5029,N_3260);
and U7795 (N_7795,N_4970,N_4558);
nor U7796 (N_7796,N_3755,N_4765);
and U7797 (N_7797,N_4234,N_3759);
nand U7798 (N_7798,N_4709,N_5391);
and U7799 (N_7799,N_4675,N_4246);
nand U7800 (N_7800,N_3404,N_5243);
and U7801 (N_7801,N_4190,N_4456);
nor U7802 (N_7802,N_4304,N_4224);
nor U7803 (N_7803,N_3094,N_3213);
and U7804 (N_7804,N_4804,N_3461);
or U7805 (N_7805,N_4409,N_4510);
and U7806 (N_7806,N_3265,N_5635);
and U7807 (N_7807,N_4606,N_4766);
or U7808 (N_7808,N_5415,N_5231);
nor U7809 (N_7809,N_5286,N_4930);
and U7810 (N_7810,N_5527,N_4703);
and U7811 (N_7811,N_5953,N_3820);
and U7812 (N_7812,N_5691,N_5104);
or U7813 (N_7813,N_4613,N_3629);
nand U7814 (N_7814,N_3748,N_3694);
or U7815 (N_7815,N_5174,N_5710);
nor U7816 (N_7816,N_4074,N_4108);
or U7817 (N_7817,N_5233,N_3738);
nor U7818 (N_7818,N_4088,N_3122);
and U7819 (N_7819,N_5391,N_4146);
or U7820 (N_7820,N_4763,N_3225);
or U7821 (N_7821,N_5572,N_3564);
or U7822 (N_7822,N_3026,N_3078);
nor U7823 (N_7823,N_5820,N_3224);
and U7824 (N_7824,N_4044,N_4026);
and U7825 (N_7825,N_4352,N_4414);
or U7826 (N_7826,N_3951,N_5880);
or U7827 (N_7827,N_5285,N_4708);
nand U7828 (N_7828,N_3271,N_5398);
nor U7829 (N_7829,N_3885,N_5808);
or U7830 (N_7830,N_4525,N_4156);
or U7831 (N_7831,N_3535,N_5095);
or U7832 (N_7832,N_5440,N_4875);
nor U7833 (N_7833,N_3528,N_5794);
nand U7834 (N_7834,N_4720,N_4575);
nand U7835 (N_7835,N_5409,N_5728);
nor U7836 (N_7836,N_3364,N_3997);
nand U7837 (N_7837,N_5632,N_3464);
nand U7838 (N_7838,N_3039,N_4576);
and U7839 (N_7839,N_3743,N_5628);
or U7840 (N_7840,N_5800,N_5076);
nand U7841 (N_7841,N_5546,N_3009);
or U7842 (N_7842,N_3180,N_3299);
nand U7843 (N_7843,N_3103,N_3829);
nor U7844 (N_7844,N_5272,N_3577);
nand U7845 (N_7845,N_4808,N_5414);
or U7846 (N_7846,N_5943,N_3715);
nor U7847 (N_7847,N_3877,N_4739);
nand U7848 (N_7848,N_5779,N_3368);
nor U7849 (N_7849,N_4334,N_4139);
or U7850 (N_7850,N_5797,N_5473);
or U7851 (N_7851,N_5982,N_4853);
nand U7852 (N_7852,N_3054,N_4983);
nor U7853 (N_7853,N_5862,N_4674);
nand U7854 (N_7854,N_4976,N_5514);
and U7855 (N_7855,N_4306,N_3819);
or U7856 (N_7856,N_3585,N_5718);
and U7857 (N_7857,N_4315,N_4463);
or U7858 (N_7858,N_3223,N_3617);
and U7859 (N_7859,N_5820,N_5615);
nor U7860 (N_7860,N_4595,N_3196);
nand U7861 (N_7861,N_4287,N_4623);
nand U7862 (N_7862,N_4104,N_4804);
or U7863 (N_7863,N_3684,N_3465);
nand U7864 (N_7864,N_4582,N_5991);
or U7865 (N_7865,N_4237,N_3838);
nor U7866 (N_7866,N_5918,N_3981);
or U7867 (N_7867,N_4758,N_3840);
or U7868 (N_7868,N_4485,N_5970);
or U7869 (N_7869,N_3966,N_4853);
nor U7870 (N_7870,N_5774,N_5001);
nand U7871 (N_7871,N_4785,N_5977);
nor U7872 (N_7872,N_4329,N_4451);
or U7873 (N_7873,N_3995,N_3839);
and U7874 (N_7874,N_4333,N_4756);
nor U7875 (N_7875,N_3753,N_5790);
nor U7876 (N_7876,N_3547,N_3085);
nand U7877 (N_7877,N_4398,N_5726);
nand U7878 (N_7878,N_5554,N_5045);
nor U7879 (N_7879,N_3457,N_5924);
or U7880 (N_7880,N_3698,N_4552);
or U7881 (N_7881,N_5951,N_3702);
nand U7882 (N_7882,N_3249,N_3789);
and U7883 (N_7883,N_4870,N_5380);
nor U7884 (N_7884,N_3985,N_3261);
nor U7885 (N_7885,N_5968,N_4909);
nand U7886 (N_7886,N_3480,N_3172);
nor U7887 (N_7887,N_5180,N_3316);
nand U7888 (N_7888,N_4089,N_4978);
nor U7889 (N_7889,N_5613,N_4997);
nand U7890 (N_7890,N_4268,N_4454);
xor U7891 (N_7891,N_4595,N_3214);
or U7892 (N_7892,N_4756,N_4694);
and U7893 (N_7893,N_5680,N_5263);
or U7894 (N_7894,N_3005,N_4035);
or U7895 (N_7895,N_3310,N_3759);
and U7896 (N_7896,N_3726,N_5395);
nor U7897 (N_7897,N_4020,N_4829);
or U7898 (N_7898,N_4786,N_3613);
nor U7899 (N_7899,N_5321,N_3443);
nor U7900 (N_7900,N_5223,N_4832);
and U7901 (N_7901,N_3686,N_4068);
or U7902 (N_7902,N_5616,N_5594);
and U7903 (N_7903,N_5876,N_3631);
or U7904 (N_7904,N_3390,N_5836);
nand U7905 (N_7905,N_3406,N_3038);
or U7906 (N_7906,N_4531,N_5152);
nand U7907 (N_7907,N_5967,N_3445);
and U7908 (N_7908,N_5543,N_3154);
or U7909 (N_7909,N_4878,N_5426);
nor U7910 (N_7910,N_4513,N_4672);
or U7911 (N_7911,N_3491,N_3679);
nand U7912 (N_7912,N_3029,N_5823);
nor U7913 (N_7913,N_3811,N_3135);
and U7914 (N_7914,N_3262,N_4916);
and U7915 (N_7915,N_4140,N_5303);
xnor U7916 (N_7916,N_5610,N_4768);
and U7917 (N_7917,N_3299,N_5980);
nor U7918 (N_7918,N_5535,N_3532);
and U7919 (N_7919,N_4466,N_4496);
nor U7920 (N_7920,N_3875,N_5574);
nand U7921 (N_7921,N_4519,N_4054);
nand U7922 (N_7922,N_5651,N_3568);
nand U7923 (N_7923,N_5707,N_3821);
nor U7924 (N_7924,N_3541,N_5899);
or U7925 (N_7925,N_5251,N_4424);
nand U7926 (N_7926,N_3886,N_5962);
nor U7927 (N_7927,N_3942,N_3214);
and U7928 (N_7928,N_3225,N_3942);
nor U7929 (N_7929,N_3634,N_3154);
or U7930 (N_7930,N_3904,N_4090);
nand U7931 (N_7931,N_5467,N_4254);
xor U7932 (N_7932,N_3366,N_4151);
nor U7933 (N_7933,N_5126,N_5886);
and U7934 (N_7934,N_3787,N_5082);
or U7935 (N_7935,N_3565,N_5591);
or U7936 (N_7936,N_5060,N_5890);
nand U7937 (N_7937,N_4544,N_5114);
and U7938 (N_7938,N_3380,N_3760);
nor U7939 (N_7939,N_3842,N_4200);
and U7940 (N_7940,N_3383,N_3778);
nand U7941 (N_7941,N_5607,N_3036);
or U7942 (N_7942,N_3081,N_4193);
or U7943 (N_7943,N_5648,N_3957);
or U7944 (N_7944,N_5780,N_3579);
or U7945 (N_7945,N_3682,N_5570);
or U7946 (N_7946,N_4880,N_5523);
or U7947 (N_7947,N_5450,N_4093);
nand U7948 (N_7948,N_4130,N_5886);
nand U7949 (N_7949,N_5817,N_3769);
and U7950 (N_7950,N_3339,N_3620);
and U7951 (N_7951,N_3053,N_5753);
nand U7952 (N_7952,N_5879,N_5185);
nor U7953 (N_7953,N_3395,N_4376);
nor U7954 (N_7954,N_5820,N_4575);
or U7955 (N_7955,N_4751,N_5582);
nand U7956 (N_7956,N_3720,N_3818);
and U7957 (N_7957,N_3820,N_5087);
or U7958 (N_7958,N_3115,N_3039);
or U7959 (N_7959,N_5030,N_5107);
or U7960 (N_7960,N_3244,N_3490);
and U7961 (N_7961,N_3274,N_4451);
or U7962 (N_7962,N_5181,N_3023);
or U7963 (N_7963,N_4729,N_5913);
nand U7964 (N_7964,N_3587,N_4442);
or U7965 (N_7965,N_4987,N_5885);
nor U7966 (N_7966,N_5496,N_3034);
and U7967 (N_7967,N_5891,N_5139);
nor U7968 (N_7968,N_4197,N_4580);
nand U7969 (N_7969,N_3527,N_3394);
and U7970 (N_7970,N_3141,N_3037);
or U7971 (N_7971,N_3440,N_5877);
nand U7972 (N_7972,N_3449,N_4931);
nor U7973 (N_7973,N_3488,N_5316);
nand U7974 (N_7974,N_4716,N_5675);
nand U7975 (N_7975,N_4850,N_4323);
or U7976 (N_7976,N_3603,N_5017);
nor U7977 (N_7977,N_3353,N_5028);
nor U7978 (N_7978,N_3699,N_5807);
and U7979 (N_7979,N_3415,N_5343);
nand U7980 (N_7980,N_5522,N_4438);
nor U7981 (N_7981,N_3196,N_5433);
nand U7982 (N_7982,N_3245,N_5380);
and U7983 (N_7983,N_3350,N_3393);
nand U7984 (N_7984,N_5493,N_5324);
nand U7985 (N_7985,N_3831,N_4759);
nand U7986 (N_7986,N_4248,N_4697);
or U7987 (N_7987,N_3073,N_4502);
or U7988 (N_7988,N_5163,N_3435);
nor U7989 (N_7989,N_5384,N_5773);
and U7990 (N_7990,N_3253,N_5663);
and U7991 (N_7991,N_5803,N_4411);
nand U7992 (N_7992,N_4798,N_4324);
nand U7993 (N_7993,N_3594,N_4724);
nor U7994 (N_7994,N_5375,N_3094);
nor U7995 (N_7995,N_4629,N_3246);
or U7996 (N_7996,N_4046,N_3486);
nor U7997 (N_7997,N_4993,N_5727);
nor U7998 (N_7998,N_4641,N_4027);
and U7999 (N_7999,N_3410,N_3325);
nand U8000 (N_8000,N_4293,N_4646);
or U8001 (N_8001,N_4197,N_4841);
nor U8002 (N_8002,N_4387,N_4220);
or U8003 (N_8003,N_3074,N_4895);
nor U8004 (N_8004,N_3820,N_3931);
or U8005 (N_8005,N_5214,N_3340);
nand U8006 (N_8006,N_3951,N_4184);
or U8007 (N_8007,N_5299,N_3330);
and U8008 (N_8008,N_5863,N_5670);
nor U8009 (N_8009,N_3441,N_3990);
nand U8010 (N_8010,N_3197,N_5637);
nor U8011 (N_8011,N_3045,N_4282);
and U8012 (N_8012,N_4782,N_5663);
nand U8013 (N_8013,N_3191,N_3823);
nand U8014 (N_8014,N_5451,N_3397);
or U8015 (N_8015,N_3366,N_4383);
and U8016 (N_8016,N_4187,N_4473);
nor U8017 (N_8017,N_4858,N_3054);
or U8018 (N_8018,N_4365,N_5845);
or U8019 (N_8019,N_4473,N_3016);
and U8020 (N_8020,N_5627,N_4738);
and U8021 (N_8021,N_3453,N_4649);
and U8022 (N_8022,N_5272,N_5733);
or U8023 (N_8023,N_5933,N_3932);
or U8024 (N_8024,N_3490,N_5879);
nor U8025 (N_8025,N_4557,N_4801);
and U8026 (N_8026,N_5705,N_4745);
nand U8027 (N_8027,N_4825,N_5731);
nand U8028 (N_8028,N_3817,N_4870);
nand U8029 (N_8029,N_4305,N_4266);
nor U8030 (N_8030,N_5314,N_3794);
nand U8031 (N_8031,N_4302,N_3118);
nand U8032 (N_8032,N_5155,N_3979);
nor U8033 (N_8033,N_3832,N_5538);
nand U8034 (N_8034,N_3555,N_3605);
or U8035 (N_8035,N_3497,N_3861);
nand U8036 (N_8036,N_3340,N_3770);
or U8037 (N_8037,N_4679,N_3331);
or U8038 (N_8038,N_5350,N_4362);
nor U8039 (N_8039,N_3438,N_3656);
and U8040 (N_8040,N_5347,N_5651);
nor U8041 (N_8041,N_3528,N_5890);
nor U8042 (N_8042,N_3058,N_5549);
and U8043 (N_8043,N_5542,N_3133);
and U8044 (N_8044,N_5710,N_3441);
or U8045 (N_8045,N_3864,N_4393);
or U8046 (N_8046,N_4445,N_4475);
nand U8047 (N_8047,N_4835,N_4874);
nor U8048 (N_8048,N_5380,N_4103);
nor U8049 (N_8049,N_4081,N_5457);
or U8050 (N_8050,N_4910,N_5377);
or U8051 (N_8051,N_5966,N_3165);
nor U8052 (N_8052,N_3664,N_5959);
nand U8053 (N_8053,N_4009,N_5966);
or U8054 (N_8054,N_3749,N_3892);
or U8055 (N_8055,N_3092,N_5197);
nand U8056 (N_8056,N_5950,N_3291);
nor U8057 (N_8057,N_5860,N_3758);
nand U8058 (N_8058,N_4971,N_4226);
nor U8059 (N_8059,N_4824,N_5442);
nor U8060 (N_8060,N_5454,N_4810);
nand U8061 (N_8061,N_4264,N_4352);
or U8062 (N_8062,N_5113,N_4986);
and U8063 (N_8063,N_5397,N_3639);
and U8064 (N_8064,N_5429,N_4611);
nor U8065 (N_8065,N_4877,N_4555);
nand U8066 (N_8066,N_3974,N_3365);
or U8067 (N_8067,N_4894,N_5764);
or U8068 (N_8068,N_5730,N_3266);
and U8069 (N_8069,N_3879,N_3561);
or U8070 (N_8070,N_3556,N_5924);
nand U8071 (N_8071,N_5600,N_5141);
nand U8072 (N_8072,N_4221,N_4264);
nor U8073 (N_8073,N_3351,N_5328);
and U8074 (N_8074,N_3509,N_3620);
nor U8075 (N_8075,N_4046,N_3583);
nor U8076 (N_8076,N_5636,N_4493);
and U8077 (N_8077,N_4671,N_3011);
or U8078 (N_8078,N_4683,N_5130);
nand U8079 (N_8079,N_3591,N_4589);
xor U8080 (N_8080,N_3721,N_4903);
or U8081 (N_8081,N_5263,N_4280);
and U8082 (N_8082,N_5878,N_3984);
or U8083 (N_8083,N_5118,N_4197);
or U8084 (N_8084,N_5543,N_3388);
or U8085 (N_8085,N_5019,N_4737);
and U8086 (N_8086,N_5091,N_5161);
nand U8087 (N_8087,N_5361,N_3149);
or U8088 (N_8088,N_4070,N_4289);
or U8089 (N_8089,N_4467,N_5069);
and U8090 (N_8090,N_3489,N_4118);
or U8091 (N_8091,N_5427,N_3213);
nand U8092 (N_8092,N_5576,N_4862);
nor U8093 (N_8093,N_5696,N_4229);
nand U8094 (N_8094,N_3018,N_3595);
xnor U8095 (N_8095,N_4204,N_3114);
nand U8096 (N_8096,N_3385,N_3826);
nand U8097 (N_8097,N_3985,N_5083);
or U8098 (N_8098,N_5820,N_4462);
or U8099 (N_8099,N_5203,N_3762);
and U8100 (N_8100,N_5080,N_5458);
nand U8101 (N_8101,N_3338,N_5170);
nand U8102 (N_8102,N_3434,N_4246);
nand U8103 (N_8103,N_4085,N_4839);
and U8104 (N_8104,N_3032,N_3704);
nor U8105 (N_8105,N_4705,N_5469);
and U8106 (N_8106,N_4066,N_3467);
and U8107 (N_8107,N_3265,N_3211);
nor U8108 (N_8108,N_3610,N_4077);
nor U8109 (N_8109,N_4647,N_3341);
or U8110 (N_8110,N_5569,N_3256);
nor U8111 (N_8111,N_4027,N_4026);
or U8112 (N_8112,N_5102,N_4658);
nand U8113 (N_8113,N_5540,N_5048);
and U8114 (N_8114,N_4239,N_5877);
and U8115 (N_8115,N_4089,N_4331);
nand U8116 (N_8116,N_4593,N_3521);
nor U8117 (N_8117,N_5770,N_3282);
nor U8118 (N_8118,N_5021,N_5429);
or U8119 (N_8119,N_5369,N_5927);
and U8120 (N_8120,N_4729,N_5757);
nand U8121 (N_8121,N_3117,N_4619);
nand U8122 (N_8122,N_5914,N_4452);
nand U8123 (N_8123,N_5516,N_4331);
nand U8124 (N_8124,N_3878,N_5278);
nand U8125 (N_8125,N_4509,N_3335);
nor U8126 (N_8126,N_5537,N_4127);
nor U8127 (N_8127,N_5452,N_5283);
nor U8128 (N_8128,N_4821,N_5844);
nand U8129 (N_8129,N_3485,N_3098);
nand U8130 (N_8130,N_3947,N_5820);
nand U8131 (N_8131,N_3969,N_5275);
or U8132 (N_8132,N_5983,N_5527);
or U8133 (N_8133,N_3761,N_4962);
nand U8134 (N_8134,N_4129,N_5027);
nand U8135 (N_8135,N_5048,N_3879);
and U8136 (N_8136,N_5428,N_4795);
nand U8137 (N_8137,N_5230,N_4071);
and U8138 (N_8138,N_3038,N_4250);
or U8139 (N_8139,N_4004,N_4990);
nor U8140 (N_8140,N_3964,N_4664);
nor U8141 (N_8141,N_3480,N_5130);
nor U8142 (N_8142,N_5844,N_3261);
nand U8143 (N_8143,N_5808,N_5044);
nor U8144 (N_8144,N_4362,N_5037);
or U8145 (N_8145,N_5277,N_3926);
or U8146 (N_8146,N_4843,N_4484);
and U8147 (N_8147,N_4902,N_4798);
and U8148 (N_8148,N_5219,N_4239);
nor U8149 (N_8149,N_3243,N_3093);
and U8150 (N_8150,N_4392,N_5138);
nand U8151 (N_8151,N_3578,N_4102);
or U8152 (N_8152,N_5278,N_5685);
and U8153 (N_8153,N_4565,N_3591);
and U8154 (N_8154,N_3494,N_3781);
nor U8155 (N_8155,N_3095,N_5885);
or U8156 (N_8156,N_3624,N_5197);
and U8157 (N_8157,N_4424,N_5811);
nor U8158 (N_8158,N_3704,N_4375);
nand U8159 (N_8159,N_4074,N_4037);
and U8160 (N_8160,N_3698,N_5409);
nand U8161 (N_8161,N_5208,N_4473);
or U8162 (N_8162,N_5001,N_3990);
nand U8163 (N_8163,N_5407,N_3757);
and U8164 (N_8164,N_5663,N_3152);
and U8165 (N_8165,N_3376,N_4198);
nand U8166 (N_8166,N_4540,N_5083);
nor U8167 (N_8167,N_4165,N_4029);
and U8168 (N_8168,N_3021,N_5940);
nor U8169 (N_8169,N_4444,N_5795);
or U8170 (N_8170,N_4176,N_5805);
and U8171 (N_8171,N_4770,N_4790);
and U8172 (N_8172,N_5911,N_3534);
or U8173 (N_8173,N_4110,N_3396);
and U8174 (N_8174,N_4997,N_4259);
or U8175 (N_8175,N_4457,N_3300);
nand U8176 (N_8176,N_4650,N_3155);
or U8177 (N_8177,N_5509,N_4582);
or U8178 (N_8178,N_4017,N_5052);
and U8179 (N_8179,N_3306,N_3905);
nand U8180 (N_8180,N_3584,N_4357);
and U8181 (N_8181,N_4525,N_5119);
nand U8182 (N_8182,N_5587,N_5284);
nand U8183 (N_8183,N_5748,N_5011);
or U8184 (N_8184,N_5112,N_4511);
nand U8185 (N_8185,N_4924,N_3111);
nand U8186 (N_8186,N_4873,N_4940);
nand U8187 (N_8187,N_3444,N_3460);
and U8188 (N_8188,N_4962,N_3663);
nor U8189 (N_8189,N_5438,N_3048);
nor U8190 (N_8190,N_5410,N_4862);
xor U8191 (N_8191,N_4503,N_3919);
nor U8192 (N_8192,N_4557,N_5828);
or U8193 (N_8193,N_3869,N_4864);
nor U8194 (N_8194,N_5509,N_3681);
and U8195 (N_8195,N_5558,N_3418);
and U8196 (N_8196,N_3492,N_4955);
or U8197 (N_8197,N_5051,N_5781);
and U8198 (N_8198,N_3479,N_3551);
nand U8199 (N_8199,N_4696,N_3987);
nand U8200 (N_8200,N_4596,N_5045);
nand U8201 (N_8201,N_5290,N_3147);
nand U8202 (N_8202,N_4487,N_3637);
nor U8203 (N_8203,N_4284,N_5163);
nand U8204 (N_8204,N_3530,N_4461);
and U8205 (N_8205,N_4128,N_5484);
nor U8206 (N_8206,N_5481,N_4529);
nand U8207 (N_8207,N_5770,N_3617);
nor U8208 (N_8208,N_3662,N_5679);
and U8209 (N_8209,N_4082,N_3416);
nand U8210 (N_8210,N_5747,N_5632);
nand U8211 (N_8211,N_4461,N_5235);
and U8212 (N_8212,N_5303,N_5614);
or U8213 (N_8213,N_5581,N_5240);
and U8214 (N_8214,N_5463,N_4009);
nand U8215 (N_8215,N_3924,N_3973);
nor U8216 (N_8216,N_3363,N_4598);
or U8217 (N_8217,N_4698,N_5782);
and U8218 (N_8218,N_5587,N_3326);
nor U8219 (N_8219,N_4161,N_5258);
nand U8220 (N_8220,N_4441,N_4679);
and U8221 (N_8221,N_4743,N_4341);
nor U8222 (N_8222,N_3559,N_3055);
nor U8223 (N_8223,N_5267,N_3384);
nor U8224 (N_8224,N_3874,N_4718);
and U8225 (N_8225,N_5876,N_3714);
nor U8226 (N_8226,N_5995,N_3902);
and U8227 (N_8227,N_3161,N_3282);
nor U8228 (N_8228,N_5978,N_3912);
nand U8229 (N_8229,N_4062,N_5274);
and U8230 (N_8230,N_5355,N_3568);
nand U8231 (N_8231,N_3542,N_3162);
nand U8232 (N_8232,N_4258,N_3211);
or U8233 (N_8233,N_5838,N_4656);
or U8234 (N_8234,N_4338,N_4395);
and U8235 (N_8235,N_5845,N_5038);
nand U8236 (N_8236,N_5537,N_4675);
or U8237 (N_8237,N_3840,N_5132);
and U8238 (N_8238,N_5807,N_3360);
nand U8239 (N_8239,N_4802,N_3260);
and U8240 (N_8240,N_5753,N_5942);
and U8241 (N_8241,N_4547,N_5186);
and U8242 (N_8242,N_4652,N_3070);
nor U8243 (N_8243,N_3880,N_5439);
or U8244 (N_8244,N_4485,N_5105);
nor U8245 (N_8245,N_3507,N_3504);
or U8246 (N_8246,N_4189,N_5900);
nand U8247 (N_8247,N_4654,N_4293);
xor U8248 (N_8248,N_4938,N_4382);
and U8249 (N_8249,N_5842,N_4153);
nand U8250 (N_8250,N_5229,N_3070);
and U8251 (N_8251,N_5996,N_5262);
or U8252 (N_8252,N_3262,N_3407);
xnor U8253 (N_8253,N_5936,N_3247);
nand U8254 (N_8254,N_4441,N_3370);
and U8255 (N_8255,N_3281,N_4860);
or U8256 (N_8256,N_5846,N_3210);
nand U8257 (N_8257,N_3841,N_5342);
and U8258 (N_8258,N_3476,N_3715);
or U8259 (N_8259,N_5044,N_3794);
and U8260 (N_8260,N_3418,N_4828);
and U8261 (N_8261,N_4622,N_3627);
and U8262 (N_8262,N_5646,N_3230);
nand U8263 (N_8263,N_3085,N_5181);
or U8264 (N_8264,N_4077,N_3551);
and U8265 (N_8265,N_3013,N_5137);
and U8266 (N_8266,N_5388,N_3865);
or U8267 (N_8267,N_3703,N_4433);
nand U8268 (N_8268,N_4894,N_4934);
nor U8269 (N_8269,N_4507,N_4544);
or U8270 (N_8270,N_5623,N_5310);
nor U8271 (N_8271,N_4544,N_4038);
and U8272 (N_8272,N_4959,N_3683);
nand U8273 (N_8273,N_5909,N_4031);
nand U8274 (N_8274,N_4682,N_3069);
and U8275 (N_8275,N_4292,N_5529);
nor U8276 (N_8276,N_4566,N_3066);
nand U8277 (N_8277,N_4871,N_3821);
and U8278 (N_8278,N_5835,N_5010);
and U8279 (N_8279,N_5057,N_5602);
or U8280 (N_8280,N_5355,N_4420);
nor U8281 (N_8281,N_5342,N_3922);
nor U8282 (N_8282,N_3493,N_5495);
and U8283 (N_8283,N_5459,N_4799);
and U8284 (N_8284,N_3284,N_5638);
and U8285 (N_8285,N_5206,N_3908);
nand U8286 (N_8286,N_5449,N_5379);
and U8287 (N_8287,N_5765,N_5374);
nand U8288 (N_8288,N_4154,N_3044);
nand U8289 (N_8289,N_4577,N_3843);
and U8290 (N_8290,N_3884,N_3483);
or U8291 (N_8291,N_3749,N_5748);
nor U8292 (N_8292,N_3874,N_4806);
and U8293 (N_8293,N_3800,N_5693);
and U8294 (N_8294,N_4131,N_5561);
nor U8295 (N_8295,N_3450,N_4248);
and U8296 (N_8296,N_3415,N_5659);
and U8297 (N_8297,N_5829,N_3904);
nor U8298 (N_8298,N_4683,N_3952);
nand U8299 (N_8299,N_5499,N_3867);
nor U8300 (N_8300,N_4744,N_3340);
and U8301 (N_8301,N_5762,N_4217);
or U8302 (N_8302,N_5211,N_4425);
and U8303 (N_8303,N_3585,N_4209);
or U8304 (N_8304,N_5157,N_5661);
or U8305 (N_8305,N_4520,N_3436);
or U8306 (N_8306,N_5999,N_3241);
or U8307 (N_8307,N_5912,N_4432);
nand U8308 (N_8308,N_5107,N_3767);
nor U8309 (N_8309,N_5276,N_4616);
or U8310 (N_8310,N_4999,N_5490);
nor U8311 (N_8311,N_5063,N_4858);
nor U8312 (N_8312,N_4288,N_4750);
nor U8313 (N_8313,N_3019,N_3806);
or U8314 (N_8314,N_5314,N_4113);
nor U8315 (N_8315,N_4967,N_5504);
xor U8316 (N_8316,N_5172,N_5956);
nand U8317 (N_8317,N_4136,N_3933);
nand U8318 (N_8318,N_5253,N_4033);
nand U8319 (N_8319,N_3947,N_3935);
or U8320 (N_8320,N_4928,N_3294);
or U8321 (N_8321,N_3413,N_3055);
nand U8322 (N_8322,N_3073,N_3975);
and U8323 (N_8323,N_3470,N_5354);
nor U8324 (N_8324,N_5928,N_4468);
and U8325 (N_8325,N_5133,N_4896);
nand U8326 (N_8326,N_4523,N_4287);
nand U8327 (N_8327,N_3714,N_4008);
or U8328 (N_8328,N_3478,N_3823);
and U8329 (N_8329,N_3473,N_4774);
nand U8330 (N_8330,N_4668,N_5288);
or U8331 (N_8331,N_5887,N_4888);
nand U8332 (N_8332,N_5952,N_4525);
nor U8333 (N_8333,N_4013,N_5205);
or U8334 (N_8334,N_4248,N_3906);
or U8335 (N_8335,N_3540,N_4499);
and U8336 (N_8336,N_4491,N_5102);
or U8337 (N_8337,N_4203,N_4581);
and U8338 (N_8338,N_4995,N_5867);
or U8339 (N_8339,N_4384,N_4386);
and U8340 (N_8340,N_5591,N_5975);
nand U8341 (N_8341,N_5968,N_4520);
nand U8342 (N_8342,N_3952,N_4092);
nor U8343 (N_8343,N_4723,N_3602);
and U8344 (N_8344,N_4309,N_4415);
xnor U8345 (N_8345,N_5726,N_4164);
nand U8346 (N_8346,N_4632,N_4440);
nor U8347 (N_8347,N_5074,N_4848);
and U8348 (N_8348,N_5347,N_3570);
nand U8349 (N_8349,N_3873,N_4871);
nor U8350 (N_8350,N_4070,N_4749);
and U8351 (N_8351,N_3761,N_5919);
and U8352 (N_8352,N_4798,N_5988);
nor U8353 (N_8353,N_5549,N_4560);
nand U8354 (N_8354,N_3512,N_5174);
and U8355 (N_8355,N_5101,N_5816);
nor U8356 (N_8356,N_5909,N_5340);
and U8357 (N_8357,N_5283,N_4639);
nor U8358 (N_8358,N_3552,N_4821);
and U8359 (N_8359,N_4441,N_3987);
and U8360 (N_8360,N_4904,N_3149);
or U8361 (N_8361,N_5757,N_3876);
and U8362 (N_8362,N_4335,N_4306);
and U8363 (N_8363,N_3292,N_4087);
or U8364 (N_8364,N_4823,N_3475);
and U8365 (N_8365,N_4943,N_3823);
or U8366 (N_8366,N_3452,N_3904);
and U8367 (N_8367,N_5332,N_5942);
nor U8368 (N_8368,N_4906,N_3069);
or U8369 (N_8369,N_5922,N_5493);
nand U8370 (N_8370,N_5189,N_4932);
or U8371 (N_8371,N_3167,N_5316);
and U8372 (N_8372,N_5959,N_5257);
or U8373 (N_8373,N_5656,N_4835);
or U8374 (N_8374,N_3068,N_3482);
and U8375 (N_8375,N_5133,N_4624);
nand U8376 (N_8376,N_4406,N_5233);
nor U8377 (N_8377,N_5311,N_3453);
nor U8378 (N_8378,N_4375,N_3404);
or U8379 (N_8379,N_5559,N_4651);
nand U8380 (N_8380,N_5856,N_3238);
xnor U8381 (N_8381,N_4083,N_4804);
and U8382 (N_8382,N_3827,N_3253);
and U8383 (N_8383,N_3738,N_5051);
or U8384 (N_8384,N_5873,N_4155);
and U8385 (N_8385,N_5495,N_3211);
nand U8386 (N_8386,N_4994,N_5980);
or U8387 (N_8387,N_5995,N_4237);
and U8388 (N_8388,N_3663,N_4764);
nand U8389 (N_8389,N_3018,N_4924);
or U8390 (N_8390,N_3735,N_4895);
nor U8391 (N_8391,N_3349,N_3772);
or U8392 (N_8392,N_5935,N_5242);
and U8393 (N_8393,N_5306,N_3071);
or U8394 (N_8394,N_3876,N_5072);
and U8395 (N_8395,N_3079,N_5267);
or U8396 (N_8396,N_4571,N_4156);
nor U8397 (N_8397,N_3638,N_4876);
and U8398 (N_8398,N_4375,N_4199);
or U8399 (N_8399,N_5836,N_3739);
and U8400 (N_8400,N_3787,N_5650);
and U8401 (N_8401,N_4302,N_4724);
and U8402 (N_8402,N_3604,N_4853);
nor U8403 (N_8403,N_5254,N_4707);
nor U8404 (N_8404,N_5107,N_3670);
nand U8405 (N_8405,N_5165,N_3744);
or U8406 (N_8406,N_4551,N_5400);
nor U8407 (N_8407,N_4860,N_3076);
or U8408 (N_8408,N_5640,N_3017);
and U8409 (N_8409,N_3722,N_5023);
nor U8410 (N_8410,N_4855,N_4438);
nand U8411 (N_8411,N_4468,N_3940);
nor U8412 (N_8412,N_3087,N_5960);
nand U8413 (N_8413,N_5924,N_5782);
and U8414 (N_8414,N_3402,N_4567);
and U8415 (N_8415,N_5070,N_5264);
and U8416 (N_8416,N_4155,N_3473);
and U8417 (N_8417,N_5970,N_4177);
and U8418 (N_8418,N_4595,N_5695);
nand U8419 (N_8419,N_4157,N_4498);
and U8420 (N_8420,N_4641,N_5569);
and U8421 (N_8421,N_3277,N_5537);
nand U8422 (N_8422,N_3990,N_3891);
nor U8423 (N_8423,N_5543,N_3253);
nand U8424 (N_8424,N_3937,N_4248);
nand U8425 (N_8425,N_3469,N_3880);
and U8426 (N_8426,N_4223,N_5096);
nor U8427 (N_8427,N_5655,N_3014);
and U8428 (N_8428,N_4764,N_5290);
nor U8429 (N_8429,N_4171,N_5019);
nand U8430 (N_8430,N_5926,N_5802);
nor U8431 (N_8431,N_5256,N_3658);
and U8432 (N_8432,N_4209,N_4576);
and U8433 (N_8433,N_3180,N_4475);
and U8434 (N_8434,N_4981,N_4396);
nand U8435 (N_8435,N_3785,N_5667);
or U8436 (N_8436,N_5182,N_5583);
nand U8437 (N_8437,N_3514,N_5136);
or U8438 (N_8438,N_3040,N_5360);
or U8439 (N_8439,N_3948,N_4212);
nor U8440 (N_8440,N_3217,N_5825);
or U8441 (N_8441,N_4735,N_4320);
and U8442 (N_8442,N_3412,N_5809);
and U8443 (N_8443,N_5973,N_5119);
nor U8444 (N_8444,N_3546,N_4175);
or U8445 (N_8445,N_5962,N_5047);
nand U8446 (N_8446,N_5833,N_5884);
nor U8447 (N_8447,N_5831,N_4568);
or U8448 (N_8448,N_3789,N_5439);
nor U8449 (N_8449,N_4055,N_4572);
and U8450 (N_8450,N_5770,N_5513);
nor U8451 (N_8451,N_3357,N_3374);
and U8452 (N_8452,N_3905,N_4720);
and U8453 (N_8453,N_5598,N_3082);
and U8454 (N_8454,N_3317,N_5215);
nor U8455 (N_8455,N_3765,N_3971);
or U8456 (N_8456,N_5945,N_5000);
and U8457 (N_8457,N_4528,N_3058);
or U8458 (N_8458,N_5907,N_3297);
nor U8459 (N_8459,N_3039,N_3521);
nand U8460 (N_8460,N_5486,N_4751);
nor U8461 (N_8461,N_4811,N_3463);
nor U8462 (N_8462,N_3130,N_4184);
nor U8463 (N_8463,N_4846,N_5837);
nor U8464 (N_8464,N_3876,N_3095);
nand U8465 (N_8465,N_5017,N_5041);
nand U8466 (N_8466,N_4053,N_4359);
or U8467 (N_8467,N_5186,N_5625);
nor U8468 (N_8468,N_3856,N_4974);
nand U8469 (N_8469,N_5267,N_3202);
or U8470 (N_8470,N_3560,N_4041);
and U8471 (N_8471,N_5005,N_4039);
nor U8472 (N_8472,N_3122,N_3269);
and U8473 (N_8473,N_3470,N_4532);
xor U8474 (N_8474,N_3189,N_4452);
and U8475 (N_8475,N_5690,N_3092);
and U8476 (N_8476,N_4419,N_5154);
nand U8477 (N_8477,N_3087,N_3484);
or U8478 (N_8478,N_3483,N_3831);
or U8479 (N_8479,N_5568,N_5049);
or U8480 (N_8480,N_3087,N_5814);
and U8481 (N_8481,N_5949,N_4089);
nand U8482 (N_8482,N_4598,N_5875);
or U8483 (N_8483,N_4764,N_3919);
nor U8484 (N_8484,N_3758,N_4427);
nor U8485 (N_8485,N_3803,N_4319);
nor U8486 (N_8486,N_3432,N_4254);
or U8487 (N_8487,N_4268,N_3083);
nor U8488 (N_8488,N_4325,N_5227);
nor U8489 (N_8489,N_3963,N_3949);
nor U8490 (N_8490,N_5975,N_5134);
or U8491 (N_8491,N_4585,N_4949);
and U8492 (N_8492,N_5729,N_5517);
and U8493 (N_8493,N_4855,N_4490);
or U8494 (N_8494,N_3660,N_3335);
or U8495 (N_8495,N_4159,N_5435);
nand U8496 (N_8496,N_5298,N_5951);
and U8497 (N_8497,N_4286,N_4920);
or U8498 (N_8498,N_5035,N_4227);
or U8499 (N_8499,N_4878,N_5858);
nand U8500 (N_8500,N_4440,N_4475);
nand U8501 (N_8501,N_3534,N_3581);
nand U8502 (N_8502,N_5816,N_5210);
nor U8503 (N_8503,N_5560,N_3642);
or U8504 (N_8504,N_4823,N_3013);
nor U8505 (N_8505,N_5555,N_5657);
nand U8506 (N_8506,N_4525,N_3541);
nand U8507 (N_8507,N_3150,N_3269);
and U8508 (N_8508,N_3192,N_5003);
nand U8509 (N_8509,N_3301,N_3217);
and U8510 (N_8510,N_5081,N_3508);
or U8511 (N_8511,N_3985,N_3486);
or U8512 (N_8512,N_3885,N_4385);
nand U8513 (N_8513,N_4509,N_4850);
nor U8514 (N_8514,N_5366,N_5515);
nand U8515 (N_8515,N_3991,N_5616);
or U8516 (N_8516,N_3910,N_4693);
or U8517 (N_8517,N_4757,N_3406);
nor U8518 (N_8518,N_3978,N_3931);
xor U8519 (N_8519,N_3786,N_3443);
and U8520 (N_8520,N_4752,N_5407);
or U8521 (N_8521,N_3731,N_3966);
or U8522 (N_8522,N_4498,N_5553);
and U8523 (N_8523,N_3933,N_3873);
and U8524 (N_8524,N_3879,N_4781);
and U8525 (N_8525,N_4912,N_3216);
nand U8526 (N_8526,N_5342,N_4486);
nand U8527 (N_8527,N_4645,N_5633);
nand U8528 (N_8528,N_5889,N_3848);
nand U8529 (N_8529,N_5479,N_4344);
or U8530 (N_8530,N_5550,N_4895);
nand U8531 (N_8531,N_3660,N_4005);
or U8532 (N_8532,N_5253,N_5193);
nand U8533 (N_8533,N_4735,N_4318);
or U8534 (N_8534,N_4442,N_3690);
nand U8535 (N_8535,N_3030,N_4513);
nand U8536 (N_8536,N_5733,N_4887);
or U8537 (N_8537,N_4545,N_3866);
nand U8538 (N_8538,N_4159,N_3439);
nand U8539 (N_8539,N_4444,N_5239);
and U8540 (N_8540,N_4563,N_3675);
and U8541 (N_8541,N_5942,N_3707);
nand U8542 (N_8542,N_5066,N_4347);
nand U8543 (N_8543,N_4937,N_3295);
nor U8544 (N_8544,N_3875,N_4549);
and U8545 (N_8545,N_3778,N_4522);
nor U8546 (N_8546,N_3818,N_4941);
or U8547 (N_8547,N_3353,N_4211);
nand U8548 (N_8548,N_5410,N_4219);
nand U8549 (N_8549,N_5649,N_5343);
or U8550 (N_8550,N_3332,N_5125);
or U8551 (N_8551,N_4348,N_5588);
or U8552 (N_8552,N_3794,N_3294);
nand U8553 (N_8553,N_5065,N_5524);
or U8554 (N_8554,N_5764,N_5268);
nor U8555 (N_8555,N_3998,N_4758);
nor U8556 (N_8556,N_3298,N_5199);
or U8557 (N_8557,N_3746,N_3007);
nor U8558 (N_8558,N_3890,N_5263);
or U8559 (N_8559,N_3627,N_5367);
and U8560 (N_8560,N_3565,N_3895);
or U8561 (N_8561,N_3400,N_3326);
or U8562 (N_8562,N_4555,N_4393);
or U8563 (N_8563,N_4175,N_5167);
nand U8564 (N_8564,N_3609,N_3873);
nor U8565 (N_8565,N_3702,N_3784);
nand U8566 (N_8566,N_4167,N_3874);
and U8567 (N_8567,N_4343,N_3998);
nor U8568 (N_8568,N_5736,N_3260);
or U8569 (N_8569,N_3803,N_3552);
and U8570 (N_8570,N_4601,N_4718);
nand U8571 (N_8571,N_5573,N_4025);
nor U8572 (N_8572,N_5264,N_4867);
and U8573 (N_8573,N_5385,N_5531);
nor U8574 (N_8574,N_3198,N_4489);
nand U8575 (N_8575,N_4922,N_4044);
or U8576 (N_8576,N_4263,N_3137);
nand U8577 (N_8577,N_4300,N_4042);
nand U8578 (N_8578,N_4645,N_3178);
nand U8579 (N_8579,N_3774,N_4622);
nor U8580 (N_8580,N_4151,N_4465);
and U8581 (N_8581,N_5235,N_3504);
xnor U8582 (N_8582,N_4972,N_3992);
nor U8583 (N_8583,N_4300,N_3410);
or U8584 (N_8584,N_5113,N_3699);
nand U8585 (N_8585,N_5371,N_5729);
nor U8586 (N_8586,N_4501,N_5606);
xnor U8587 (N_8587,N_5491,N_4901);
and U8588 (N_8588,N_4549,N_5842);
xnor U8589 (N_8589,N_4911,N_5160);
or U8590 (N_8590,N_3479,N_3588);
nor U8591 (N_8591,N_4613,N_4172);
nor U8592 (N_8592,N_4690,N_3329);
or U8593 (N_8593,N_5949,N_3128);
and U8594 (N_8594,N_5579,N_5857);
and U8595 (N_8595,N_4153,N_4739);
or U8596 (N_8596,N_5740,N_4346);
and U8597 (N_8597,N_4826,N_4494);
nor U8598 (N_8598,N_3903,N_4074);
or U8599 (N_8599,N_5006,N_4143);
nand U8600 (N_8600,N_4546,N_4626);
nand U8601 (N_8601,N_5579,N_3678);
nor U8602 (N_8602,N_4977,N_5376);
and U8603 (N_8603,N_4105,N_4373);
and U8604 (N_8604,N_3180,N_4312);
and U8605 (N_8605,N_5821,N_5994);
or U8606 (N_8606,N_5568,N_4157);
and U8607 (N_8607,N_5152,N_5281);
nor U8608 (N_8608,N_4857,N_4781);
and U8609 (N_8609,N_5425,N_3963);
and U8610 (N_8610,N_5739,N_3998);
or U8611 (N_8611,N_5990,N_5855);
and U8612 (N_8612,N_4817,N_5907);
and U8613 (N_8613,N_5089,N_4807);
nand U8614 (N_8614,N_5756,N_3024);
or U8615 (N_8615,N_3161,N_5559);
nand U8616 (N_8616,N_3568,N_3030);
nand U8617 (N_8617,N_3038,N_3947);
nand U8618 (N_8618,N_3193,N_5636);
and U8619 (N_8619,N_3683,N_3758);
or U8620 (N_8620,N_5938,N_3463);
and U8621 (N_8621,N_3179,N_4188);
or U8622 (N_8622,N_4737,N_5844);
nor U8623 (N_8623,N_5053,N_5584);
or U8624 (N_8624,N_3323,N_3325);
and U8625 (N_8625,N_4231,N_4258);
and U8626 (N_8626,N_5828,N_3750);
nor U8627 (N_8627,N_4112,N_5377);
and U8628 (N_8628,N_3573,N_5681);
or U8629 (N_8629,N_5104,N_3462);
nand U8630 (N_8630,N_4348,N_3001);
or U8631 (N_8631,N_4477,N_5162);
or U8632 (N_8632,N_5187,N_4650);
and U8633 (N_8633,N_4071,N_4822);
or U8634 (N_8634,N_4042,N_5741);
and U8635 (N_8635,N_5260,N_4966);
nand U8636 (N_8636,N_4756,N_5267);
or U8637 (N_8637,N_3550,N_5601);
nand U8638 (N_8638,N_4785,N_5320);
or U8639 (N_8639,N_5968,N_4780);
nand U8640 (N_8640,N_5135,N_4152);
or U8641 (N_8641,N_4233,N_5303);
and U8642 (N_8642,N_3535,N_3773);
or U8643 (N_8643,N_3197,N_5995);
and U8644 (N_8644,N_5858,N_4480);
nand U8645 (N_8645,N_4479,N_3217);
nand U8646 (N_8646,N_3975,N_5714);
nand U8647 (N_8647,N_4530,N_5731);
or U8648 (N_8648,N_4486,N_5520);
or U8649 (N_8649,N_3210,N_3174);
and U8650 (N_8650,N_4733,N_3667);
or U8651 (N_8651,N_3395,N_5074);
nand U8652 (N_8652,N_3106,N_3887);
nor U8653 (N_8653,N_4747,N_5127);
or U8654 (N_8654,N_5308,N_3288);
and U8655 (N_8655,N_3863,N_4557);
and U8656 (N_8656,N_5145,N_4921);
and U8657 (N_8657,N_4619,N_4510);
nor U8658 (N_8658,N_4396,N_4405);
nand U8659 (N_8659,N_4179,N_5833);
or U8660 (N_8660,N_4694,N_5406);
or U8661 (N_8661,N_5922,N_4385);
nor U8662 (N_8662,N_4219,N_5369);
nor U8663 (N_8663,N_5447,N_4871);
nor U8664 (N_8664,N_3823,N_4635);
nor U8665 (N_8665,N_4999,N_5798);
nand U8666 (N_8666,N_3449,N_4135);
nand U8667 (N_8667,N_3563,N_4775);
nand U8668 (N_8668,N_4629,N_4771);
and U8669 (N_8669,N_5845,N_4257);
or U8670 (N_8670,N_3113,N_3111);
nand U8671 (N_8671,N_4767,N_5904);
and U8672 (N_8672,N_4709,N_3843);
nand U8673 (N_8673,N_4013,N_4671);
nor U8674 (N_8674,N_3847,N_3661);
nand U8675 (N_8675,N_3053,N_5871);
nor U8676 (N_8676,N_5400,N_5844);
and U8677 (N_8677,N_5922,N_4096);
nor U8678 (N_8678,N_5511,N_5005);
or U8679 (N_8679,N_3117,N_5047);
or U8680 (N_8680,N_3358,N_5375);
or U8681 (N_8681,N_4757,N_4626);
and U8682 (N_8682,N_5997,N_3507);
or U8683 (N_8683,N_5707,N_5701);
nand U8684 (N_8684,N_4062,N_5305);
or U8685 (N_8685,N_5847,N_3322);
nor U8686 (N_8686,N_3204,N_3780);
or U8687 (N_8687,N_3539,N_3657);
nor U8688 (N_8688,N_3795,N_3780);
nand U8689 (N_8689,N_5517,N_4324);
nor U8690 (N_8690,N_4479,N_3625);
nor U8691 (N_8691,N_3034,N_5066);
nor U8692 (N_8692,N_3110,N_4609);
and U8693 (N_8693,N_3616,N_4788);
and U8694 (N_8694,N_3701,N_4063);
nor U8695 (N_8695,N_5910,N_5126);
or U8696 (N_8696,N_4521,N_5888);
and U8697 (N_8697,N_3544,N_3299);
nand U8698 (N_8698,N_5572,N_5027);
nand U8699 (N_8699,N_3897,N_5876);
and U8700 (N_8700,N_3634,N_3819);
or U8701 (N_8701,N_3941,N_4547);
nand U8702 (N_8702,N_3927,N_3007);
or U8703 (N_8703,N_3186,N_5153);
and U8704 (N_8704,N_5012,N_4474);
and U8705 (N_8705,N_3002,N_4527);
nor U8706 (N_8706,N_4684,N_5478);
xnor U8707 (N_8707,N_5992,N_4777);
nand U8708 (N_8708,N_3120,N_4467);
nand U8709 (N_8709,N_5541,N_5355);
nor U8710 (N_8710,N_5895,N_3804);
or U8711 (N_8711,N_4741,N_3963);
or U8712 (N_8712,N_5565,N_4522);
nor U8713 (N_8713,N_4127,N_4046);
xnor U8714 (N_8714,N_3149,N_4163);
xor U8715 (N_8715,N_4606,N_3535);
or U8716 (N_8716,N_5472,N_3856);
nor U8717 (N_8717,N_3203,N_5955);
nand U8718 (N_8718,N_4145,N_4929);
and U8719 (N_8719,N_5648,N_3979);
and U8720 (N_8720,N_5435,N_5129);
nor U8721 (N_8721,N_5512,N_5450);
or U8722 (N_8722,N_5747,N_5696);
and U8723 (N_8723,N_4372,N_3197);
and U8724 (N_8724,N_3167,N_5011);
nand U8725 (N_8725,N_5998,N_5637);
nor U8726 (N_8726,N_4224,N_3335);
or U8727 (N_8727,N_5333,N_4668);
nand U8728 (N_8728,N_3075,N_4353);
or U8729 (N_8729,N_4771,N_4943);
and U8730 (N_8730,N_5391,N_5927);
nand U8731 (N_8731,N_4090,N_4630);
nor U8732 (N_8732,N_5589,N_3343);
nand U8733 (N_8733,N_5300,N_5533);
nand U8734 (N_8734,N_5659,N_5067);
or U8735 (N_8735,N_5461,N_3978);
or U8736 (N_8736,N_4930,N_5791);
and U8737 (N_8737,N_5415,N_5377);
or U8738 (N_8738,N_5090,N_4488);
nor U8739 (N_8739,N_3719,N_3817);
or U8740 (N_8740,N_4929,N_5893);
nor U8741 (N_8741,N_4729,N_4250);
or U8742 (N_8742,N_5298,N_3479);
nor U8743 (N_8743,N_5476,N_3251);
and U8744 (N_8744,N_5531,N_5999);
or U8745 (N_8745,N_3975,N_3895);
nor U8746 (N_8746,N_3548,N_4165);
nand U8747 (N_8747,N_4198,N_4921);
nor U8748 (N_8748,N_4930,N_5388);
and U8749 (N_8749,N_4236,N_4107);
nand U8750 (N_8750,N_3722,N_5339);
and U8751 (N_8751,N_5369,N_5274);
nor U8752 (N_8752,N_5852,N_4635);
and U8753 (N_8753,N_4621,N_3925);
and U8754 (N_8754,N_4121,N_5632);
nand U8755 (N_8755,N_3146,N_4373);
and U8756 (N_8756,N_5237,N_5322);
or U8757 (N_8757,N_5522,N_3764);
or U8758 (N_8758,N_5341,N_4262);
nor U8759 (N_8759,N_3348,N_3299);
and U8760 (N_8760,N_4763,N_3742);
and U8761 (N_8761,N_3832,N_5970);
nor U8762 (N_8762,N_4785,N_3532);
nor U8763 (N_8763,N_4655,N_4196);
nor U8764 (N_8764,N_3665,N_4833);
nand U8765 (N_8765,N_5346,N_5347);
nand U8766 (N_8766,N_5006,N_3348);
nor U8767 (N_8767,N_5719,N_5409);
nand U8768 (N_8768,N_3458,N_5436);
and U8769 (N_8769,N_3751,N_3519);
or U8770 (N_8770,N_5223,N_4717);
nor U8771 (N_8771,N_4663,N_4513);
nor U8772 (N_8772,N_3852,N_5773);
and U8773 (N_8773,N_5073,N_3680);
xor U8774 (N_8774,N_5514,N_3665);
and U8775 (N_8775,N_4998,N_5087);
or U8776 (N_8776,N_4307,N_3694);
nor U8777 (N_8777,N_3994,N_3925);
nor U8778 (N_8778,N_5526,N_3957);
or U8779 (N_8779,N_5504,N_3326);
xnor U8780 (N_8780,N_5226,N_3456);
nand U8781 (N_8781,N_4611,N_5575);
or U8782 (N_8782,N_3022,N_4747);
nor U8783 (N_8783,N_4857,N_4807);
nor U8784 (N_8784,N_3236,N_4525);
or U8785 (N_8785,N_5882,N_3837);
and U8786 (N_8786,N_3945,N_5814);
nand U8787 (N_8787,N_5274,N_4101);
and U8788 (N_8788,N_3607,N_4363);
nor U8789 (N_8789,N_4386,N_3043);
and U8790 (N_8790,N_3406,N_5657);
and U8791 (N_8791,N_3579,N_4696);
and U8792 (N_8792,N_4835,N_4222);
and U8793 (N_8793,N_5664,N_3335);
nor U8794 (N_8794,N_5006,N_4711);
and U8795 (N_8795,N_3671,N_3489);
or U8796 (N_8796,N_3404,N_3690);
nand U8797 (N_8797,N_4500,N_4659);
nand U8798 (N_8798,N_4932,N_4830);
or U8799 (N_8799,N_3305,N_3616);
and U8800 (N_8800,N_3600,N_3672);
nor U8801 (N_8801,N_4827,N_4724);
or U8802 (N_8802,N_4455,N_3005);
nor U8803 (N_8803,N_5062,N_4434);
or U8804 (N_8804,N_4830,N_4544);
and U8805 (N_8805,N_5562,N_5446);
or U8806 (N_8806,N_5808,N_4462);
nor U8807 (N_8807,N_5499,N_3745);
and U8808 (N_8808,N_4093,N_5834);
nand U8809 (N_8809,N_4450,N_3651);
nand U8810 (N_8810,N_4929,N_4532);
nor U8811 (N_8811,N_5701,N_3903);
or U8812 (N_8812,N_4980,N_5759);
nor U8813 (N_8813,N_3082,N_3761);
and U8814 (N_8814,N_3004,N_5164);
or U8815 (N_8815,N_4992,N_5484);
and U8816 (N_8816,N_4501,N_3396);
or U8817 (N_8817,N_4069,N_5244);
nor U8818 (N_8818,N_4219,N_4624);
or U8819 (N_8819,N_3256,N_5216);
nor U8820 (N_8820,N_4445,N_3832);
nor U8821 (N_8821,N_5388,N_5661);
nand U8822 (N_8822,N_3607,N_3473);
and U8823 (N_8823,N_4864,N_4812);
nor U8824 (N_8824,N_4157,N_5496);
or U8825 (N_8825,N_4684,N_4745);
nand U8826 (N_8826,N_3099,N_4858);
and U8827 (N_8827,N_4746,N_5617);
and U8828 (N_8828,N_5888,N_4607);
or U8829 (N_8829,N_5974,N_5723);
or U8830 (N_8830,N_5891,N_5657);
and U8831 (N_8831,N_3518,N_3445);
or U8832 (N_8832,N_4027,N_4651);
or U8833 (N_8833,N_3928,N_5685);
nand U8834 (N_8834,N_3814,N_4563);
nor U8835 (N_8835,N_4905,N_5402);
nand U8836 (N_8836,N_4169,N_4603);
nor U8837 (N_8837,N_5932,N_3164);
nor U8838 (N_8838,N_5144,N_4050);
nor U8839 (N_8839,N_4260,N_4524);
nand U8840 (N_8840,N_4245,N_3944);
nor U8841 (N_8841,N_5543,N_5523);
nor U8842 (N_8842,N_4833,N_4100);
and U8843 (N_8843,N_3871,N_3766);
nand U8844 (N_8844,N_5865,N_5311);
nor U8845 (N_8845,N_5340,N_3718);
nand U8846 (N_8846,N_5185,N_3672);
nor U8847 (N_8847,N_4560,N_3233);
nor U8848 (N_8848,N_4518,N_4652);
nor U8849 (N_8849,N_4784,N_5082);
or U8850 (N_8850,N_4877,N_5223);
nand U8851 (N_8851,N_5023,N_3663);
nand U8852 (N_8852,N_5046,N_5525);
nand U8853 (N_8853,N_5410,N_3595);
nor U8854 (N_8854,N_5513,N_4606);
or U8855 (N_8855,N_3060,N_3079);
nor U8856 (N_8856,N_5969,N_3795);
nand U8857 (N_8857,N_5595,N_4901);
and U8858 (N_8858,N_5876,N_4321);
nand U8859 (N_8859,N_4167,N_4734);
or U8860 (N_8860,N_5337,N_5734);
xnor U8861 (N_8861,N_4967,N_5536);
or U8862 (N_8862,N_3734,N_5643);
nor U8863 (N_8863,N_4923,N_5222);
and U8864 (N_8864,N_3577,N_5625);
nor U8865 (N_8865,N_4835,N_5649);
nand U8866 (N_8866,N_3452,N_5491);
and U8867 (N_8867,N_3066,N_5864);
nand U8868 (N_8868,N_5530,N_3730);
or U8869 (N_8869,N_3952,N_5535);
or U8870 (N_8870,N_4201,N_3209);
or U8871 (N_8871,N_5649,N_3213);
nor U8872 (N_8872,N_3381,N_5751);
and U8873 (N_8873,N_5513,N_4637);
nor U8874 (N_8874,N_4262,N_5238);
and U8875 (N_8875,N_3747,N_5784);
nand U8876 (N_8876,N_4118,N_5902);
nor U8877 (N_8877,N_5934,N_3248);
or U8878 (N_8878,N_5765,N_3836);
nor U8879 (N_8879,N_3212,N_3432);
nand U8880 (N_8880,N_5412,N_5700);
nor U8881 (N_8881,N_4037,N_5834);
nor U8882 (N_8882,N_5337,N_4204);
and U8883 (N_8883,N_3561,N_3805);
nand U8884 (N_8884,N_4696,N_3117);
nand U8885 (N_8885,N_3357,N_3836);
or U8886 (N_8886,N_3616,N_4911);
or U8887 (N_8887,N_3752,N_5192);
and U8888 (N_8888,N_4329,N_5265);
and U8889 (N_8889,N_4041,N_3458);
nor U8890 (N_8890,N_4732,N_5387);
and U8891 (N_8891,N_5747,N_3666);
and U8892 (N_8892,N_5940,N_4452);
or U8893 (N_8893,N_5520,N_4096);
nor U8894 (N_8894,N_5042,N_3506);
and U8895 (N_8895,N_3209,N_5055);
nor U8896 (N_8896,N_4734,N_3872);
and U8897 (N_8897,N_4032,N_3511);
or U8898 (N_8898,N_3837,N_5586);
or U8899 (N_8899,N_4155,N_4768);
nand U8900 (N_8900,N_4989,N_3937);
nor U8901 (N_8901,N_4860,N_4397);
nand U8902 (N_8902,N_3953,N_4707);
and U8903 (N_8903,N_4881,N_3701);
nand U8904 (N_8904,N_4152,N_4844);
xnor U8905 (N_8905,N_5553,N_3728);
and U8906 (N_8906,N_4056,N_5107);
nor U8907 (N_8907,N_3924,N_5509);
or U8908 (N_8908,N_4077,N_4372);
nor U8909 (N_8909,N_5738,N_5043);
and U8910 (N_8910,N_3952,N_4699);
nand U8911 (N_8911,N_3712,N_5659);
or U8912 (N_8912,N_4384,N_4352);
or U8913 (N_8913,N_4546,N_4662);
nor U8914 (N_8914,N_4866,N_3319);
and U8915 (N_8915,N_4238,N_5156);
nand U8916 (N_8916,N_4601,N_5554);
and U8917 (N_8917,N_4065,N_5945);
nand U8918 (N_8918,N_5480,N_5373);
and U8919 (N_8919,N_3042,N_3902);
and U8920 (N_8920,N_3214,N_3361);
nor U8921 (N_8921,N_3882,N_3855);
and U8922 (N_8922,N_5847,N_5124);
or U8923 (N_8923,N_5119,N_4600);
or U8924 (N_8924,N_3186,N_4865);
nand U8925 (N_8925,N_5058,N_3248);
nand U8926 (N_8926,N_5880,N_3080);
xor U8927 (N_8927,N_5941,N_3562);
and U8928 (N_8928,N_5274,N_3925);
nor U8929 (N_8929,N_5196,N_4500);
nand U8930 (N_8930,N_3978,N_4717);
or U8931 (N_8931,N_4668,N_4558);
or U8932 (N_8932,N_4625,N_3248);
or U8933 (N_8933,N_5441,N_4666);
or U8934 (N_8934,N_4146,N_3723);
nand U8935 (N_8935,N_5900,N_5998);
or U8936 (N_8936,N_3103,N_3381);
or U8937 (N_8937,N_3847,N_4492);
nand U8938 (N_8938,N_3111,N_3238);
or U8939 (N_8939,N_3139,N_4283);
and U8940 (N_8940,N_4911,N_3144);
nor U8941 (N_8941,N_4634,N_3999);
and U8942 (N_8942,N_3075,N_3739);
or U8943 (N_8943,N_4309,N_3067);
or U8944 (N_8944,N_4515,N_4579);
nand U8945 (N_8945,N_4436,N_4257);
and U8946 (N_8946,N_4209,N_5920);
and U8947 (N_8947,N_3858,N_4108);
nor U8948 (N_8948,N_5119,N_3528);
or U8949 (N_8949,N_3654,N_5221);
nand U8950 (N_8950,N_5790,N_5430);
nor U8951 (N_8951,N_4779,N_4455);
nand U8952 (N_8952,N_5790,N_5312);
or U8953 (N_8953,N_5773,N_3371);
or U8954 (N_8954,N_5692,N_3165);
nand U8955 (N_8955,N_5296,N_5960);
nor U8956 (N_8956,N_4208,N_4641);
nor U8957 (N_8957,N_5922,N_5190);
nand U8958 (N_8958,N_5000,N_4020);
nor U8959 (N_8959,N_3677,N_3192);
xor U8960 (N_8960,N_3752,N_4493);
nor U8961 (N_8961,N_3584,N_5745);
and U8962 (N_8962,N_3753,N_5684);
nor U8963 (N_8963,N_4394,N_5066);
nor U8964 (N_8964,N_5039,N_4658);
nand U8965 (N_8965,N_3372,N_5464);
nor U8966 (N_8966,N_5435,N_5468);
and U8967 (N_8967,N_4442,N_4502);
and U8968 (N_8968,N_3935,N_4071);
and U8969 (N_8969,N_3996,N_5901);
or U8970 (N_8970,N_4219,N_3222);
nand U8971 (N_8971,N_5509,N_4116);
and U8972 (N_8972,N_5724,N_4215);
or U8973 (N_8973,N_4319,N_5753);
or U8974 (N_8974,N_3054,N_5614);
and U8975 (N_8975,N_4582,N_3677);
nor U8976 (N_8976,N_5163,N_5045);
and U8977 (N_8977,N_3385,N_3599);
or U8978 (N_8978,N_4296,N_5632);
nor U8979 (N_8979,N_5950,N_5504);
nor U8980 (N_8980,N_5296,N_4879);
or U8981 (N_8981,N_4005,N_5155);
or U8982 (N_8982,N_5388,N_4513);
nor U8983 (N_8983,N_3529,N_5323);
and U8984 (N_8984,N_4441,N_4163);
and U8985 (N_8985,N_5376,N_4350);
nor U8986 (N_8986,N_5368,N_5518);
and U8987 (N_8987,N_5940,N_4700);
or U8988 (N_8988,N_3886,N_5483);
and U8989 (N_8989,N_3468,N_4272);
or U8990 (N_8990,N_5159,N_3188);
nor U8991 (N_8991,N_3581,N_4692);
nand U8992 (N_8992,N_5576,N_3175);
nand U8993 (N_8993,N_5625,N_5657);
or U8994 (N_8994,N_3276,N_3844);
nand U8995 (N_8995,N_5639,N_5860);
or U8996 (N_8996,N_3913,N_4096);
nand U8997 (N_8997,N_3246,N_4060);
nor U8998 (N_8998,N_4635,N_5279);
and U8999 (N_8999,N_5539,N_3515);
nor U9000 (N_9000,N_8676,N_7469);
nor U9001 (N_9001,N_8183,N_7557);
or U9002 (N_9002,N_6993,N_6059);
nor U9003 (N_9003,N_6356,N_8873);
and U9004 (N_9004,N_7994,N_6101);
or U9005 (N_9005,N_8947,N_6047);
and U9006 (N_9006,N_8352,N_6032);
nand U9007 (N_9007,N_8263,N_6697);
and U9008 (N_9008,N_7555,N_7827);
or U9009 (N_9009,N_8006,N_6541);
nand U9010 (N_9010,N_7166,N_7013);
and U9011 (N_9011,N_8554,N_6397);
and U9012 (N_9012,N_8719,N_7476);
or U9013 (N_9013,N_7628,N_7489);
and U9014 (N_9014,N_7864,N_7097);
or U9015 (N_9015,N_7137,N_8570);
nand U9016 (N_9016,N_7958,N_6870);
nor U9017 (N_9017,N_8555,N_8191);
nand U9018 (N_9018,N_8730,N_6358);
nand U9019 (N_9019,N_7580,N_6796);
and U9020 (N_9020,N_6269,N_7216);
nor U9021 (N_9021,N_7867,N_8951);
and U9022 (N_9022,N_6716,N_7033);
or U9023 (N_9023,N_7724,N_7534);
or U9024 (N_9024,N_7665,N_6134);
or U9025 (N_9025,N_6316,N_7548);
nand U9026 (N_9026,N_6312,N_7083);
nor U9027 (N_9027,N_8445,N_6942);
nor U9028 (N_9028,N_8435,N_7089);
nand U9029 (N_9029,N_7700,N_7487);
xnor U9030 (N_9030,N_6086,N_7415);
nor U9031 (N_9031,N_8962,N_7505);
nand U9032 (N_9032,N_8330,N_7587);
xnor U9033 (N_9033,N_6749,N_7894);
and U9034 (N_9034,N_7854,N_6744);
or U9035 (N_9035,N_8140,N_8997);
nor U9036 (N_9036,N_6394,N_7046);
nand U9037 (N_9037,N_6966,N_6897);
or U9038 (N_9038,N_6343,N_6932);
nand U9039 (N_9039,N_7132,N_7825);
and U9040 (N_9040,N_6490,N_8147);
and U9041 (N_9041,N_8159,N_6708);
nor U9042 (N_9042,N_6309,N_7733);
or U9043 (N_9043,N_8866,N_8920);
nor U9044 (N_9044,N_8833,N_7435);
nor U9045 (N_9045,N_7511,N_6165);
and U9046 (N_9046,N_8747,N_6650);
nand U9047 (N_9047,N_6843,N_8665);
nand U9048 (N_9048,N_8662,N_7103);
nand U9049 (N_9049,N_8046,N_6042);
nor U9050 (N_9050,N_8444,N_8313);
nand U9051 (N_9051,N_8639,N_7217);
nor U9052 (N_9052,N_8457,N_8891);
nor U9053 (N_9053,N_8706,N_7093);
nor U9054 (N_9054,N_6694,N_6637);
nor U9055 (N_9055,N_6570,N_6132);
and U9056 (N_9056,N_6168,N_8825);
or U9057 (N_9057,N_8704,N_8558);
nor U9058 (N_9058,N_7831,N_8057);
and U9059 (N_9059,N_7621,N_7065);
or U9060 (N_9060,N_6430,N_8656);
nor U9061 (N_9061,N_6439,N_7997);
nor U9062 (N_9062,N_8212,N_8083);
and U9063 (N_9063,N_8561,N_7053);
nand U9064 (N_9064,N_6040,N_8168);
and U9065 (N_9065,N_8431,N_6767);
or U9066 (N_9066,N_6543,N_7535);
and U9067 (N_9067,N_8996,N_6863);
and U9068 (N_9068,N_6894,N_7481);
and U9069 (N_9069,N_7357,N_8848);
or U9070 (N_9070,N_8139,N_6081);
and U9071 (N_9071,N_6948,N_7752);
and U9072 (N_9072,N_6636,N_6555);
nor U9073 (N_9073,N_6135,N_6520);
and U9074 (N_9074,N_7992,N_7637);
nand U9075 (N_9075,N_8312,N_6099);
and U9076 (N_9076,N_6146,N_7664);
and U9077 (N_9077,N_8541,N_6917);
nand U9078 (N_9078,N_6869,N_6061);
nand U9079 (N_9079,N_7183,N_8889);
and U9080 (N_9080,N_8539,N_6437);
nand U9081 (N_9081,N_6803,N_6524);
nor U9082 (N_9082,N_6922,N_8577);
or U9083 (N_9083,N_8478,N_8852);
and U9084 (N_9084,N_7066,N_7638);
and U9085 (N_9085,N_8547,N_6734);
nor U9086 (N_9086,N_8290,N_7988);
and U9087 (N_9087,N_6362,N_8520);
and U9088 (N_9088,N_7869,N_7981);
or U9089 (N_9089,N_7881,N_7903);
or U9090 (N_9090,N_8461,N_7510);
and U9091 (N_9091,N_8247,N_6409);
nand U9092 (N_9092,N_8724,N_7188);
or U9093 (N_9093,N_7552,N_7165);
or U9094 (N_9094,N_7084,N_6652);
nor U9095 (N_9095,N_7015,N_7687);
nand U9096 (N_9096,N_6185,N_8750);
and U9097 (N_9097,N_7815,N_6581);
xor U9098 (N_9098,N_6895,N_7373);
or U9099 (N_9099,N_6314,N_7719);
nand U9100 (N_9100,N_8632,N_7159);
nor U9101 (N_9101,N_7214,N_7937);
nand U9102 (N_9102,N_6308,N_7744);
nor U9103 (N_9103,N_7675,N_8772);
or U9104 (N_9104,N_7797,N_6190);
and U9105 (N_9105,N_6002,N_7443);
or U9106 (N_9106,N_7883,N_6600);
nand U9107 (N_9107,N_7351,N_7227);
and U9108 (N_9108,N_7960,N_6363);
nand U9109 (N_9109,N_8036,N_8427);
or U9110 (N_9110,N_8583,N_6423);
and U9111 (N_9111,N_7269,N_6022);
and U9112 (N_9112,N_7512,N_6635);
or U9113 (N_9113,N_7905,N_6984);
nor U9114 (N_9114,N_7353,N_7800);
or U9115 (N_9115,N_6127,N_7394);
nor U9116 (N_9116,N_8945,N_8801);
nand U9117 (N_9117,N_7769,N_8766);
and U9118 (N_9118,N_7514,N_7829);
and U9119 (N_9119,N_6854,N_8410);
or U9120 (N_9120,N_7395,N_7418);
xnor U9121 (N_9121,N_6735,N_7316);
nand U9122 (N_9122,N_6189,N_8409);
nand U9123 (N_9123,N_6727,N_8213);
or U9124 (N_9124,N_6176,N_8818);
and U9125 (N_9125,N_8783,N_8118);
or U9126 (N_9126,N_8727,N_6859);
and U9127 (N_9127,N_6242,N_8879);
nand U9128 (N_9128,N_8636,N_8426);
and U9129 (N_9129,N_8005,N_8549);
nand U9130 (N_9130,N_8963,N_8720);
nand U9131 (N_9131,N_8507,N_7276);
nand U9132 (N_9132,N_6221,N_7725);
xor U9133 (N_9133,N_8862,N_6286);
and U9134 (N_9134,N_7895,N_6526);
or U9135 (N_9135,N_8565,N_6017);
or U9136 (N_9136,N_6462,N_8019);
and U9137 (N_9137,N_6631,N_7948);
nor U9138 (N_9138,N_7100,N_7607);
nor U9139 (N_9139,N_6626,N_8047);
nand U9140 (N_9140,N_6045,N_6724);
and U9141 (N_9141,N_6407,N_6043);
nand U9142 (N_9142,N_6172,N_7402);
or U9143 (N_9143,N_8530,N_6392);
nor U9144 (N_9144,N_7757,N_6512);
nor U9145 (N_9145,N_8420,N_8712);
nor U9146 (N_9146,N_7080,N_6569);
and U9147 (N_9147,N_6780,N_7537);
or U9148 (N_9148,N_6548,N_8128);
nor U9149 (N_9149,N_6740,N_6949);
or U9150 (N_9150,N_6274,N_7925);
or U9151 (N_9151,N_7658,N_7691);
nand U9152 (N_9152,N_6074,N_6317);
nand U9153 (N_9153,N_7283,N_6436);
and U9154 (N_9154,N_8543,N_6521);
and U9155 (N_9155,N_7078,N_6050);
and U9156 (N_9156,N_8514,N_8796);
nand U9157 (N_9157,N_7244,N_7285);
nand U9158 (N_9158,N_6239,N_7626);
and U9159 (N_9159,N_7866,N_7914);
nand U9160 (N_9160,N_7023,N_7301);
nor U9161 (N_9161,N_6339,N_8707);
nor U9162 (N_9162,N_7966,N_6464);
and U9163 (N_9163,N_6479,N_7462);
nor U9164 (N_9164,N_8396,N_6641);
or U9165 (N_9165,N_7693,N_7671);
and U9166 (N_9166,N_6206,N_8193);
nor U9167 (N_9167,N_8200,N_8517);
or U9168 (N_9168,N_6055,N_7928);
or U9169 (N_9169,N_7554,N_6240);
nand U9170 (N_9170,N_8575,N_8936);
nand U9171 (N_9171,N_7528,N_8279);
nand U9172 (N_9172,N_7531,N_8844);
nor U9173 (N_9173,N_7593,N_8782);
and U9174 (N_9174,N_7375,N_6842);
and U9175 (N_9175,N_7323,N_8502);
and U9176 (N_9176,N_6654,N_8902);
and U9177 (N_9177,N_7899,N_7906);
nand U9178 (N_9178,N_6044,N_6179);
or U9179 (N_9179,N_7965,N_8276);
nor U9180 (N_9180,N_6372,N_8692);
or U9181 (N_9181,N_6364,N_8949);
and U9182 (N_9182,N_6933,N_7119);
nor U9183 (N_9183,N_6324,N_7796);
or U9184 (N_9184,N_6277,N_8806);
nor U9185 (N_9185,N_8999,N_7943);
nand U9186 (N_9186,N_6784,N_7525);
and U9187 (N_9187,N_7245,N_7047);
nand U9188 (N_9188,N_6878,N_8081);
or U9189 (N_9189,N_8967,N_6927);
or U9190 (N_9190,N_8856,N_8850);
nor U9191 (N_9191,N_6881,N_6910);
nor U9192 (N_9192,N_7211,N_7989);
nand U9193 (N_9193,N_8647,N_6432);
nor U9194 (N_9194,N_8122,N_8232);
nor U9195 (N_9195,N_8425,N_8474);
nor U9196 (N_9196,N_7057,N_7001);
or U9197 (N_9197,N_7616,N_6589);
nor U9198 (N_9198,N_6906,N_8485);
or U9199 (N_9199,N_8983,N_6338);
or U9200 (N_9200,N_7926,N_8239);
nor U9201 (N_9201,N_7924,N_7884);
and U9202 (N_9202,N_8469,N_7496);
and U9203 (N_9203,N_7542,N_7758);
or U9204 (N_9204,N_6429,N_8815);
and U9205 (N_9205,N_6300,N_7314);
nor U9206 (N_9206,N_7967,N_6331);
or U9207 (N_9207,N_8436,N_6728);
and U9208 (N_9208,N_7972,N_8791);
or U9209 (N_9209,N_6578,N_7911);
and U9210 (N_9210,N_6396,N_6427);
or U9211 (N_9211,N_8695,N_8799);
nand U9212 (N_9212,N_7399,N_7169);
nor U9213 (N_9213,N_6198,N_8854);
nand U9214 (N_9214,N_6835,N_6037);
nand U9215 (N_9215,N_6930,N_6504);
or U9216 (N_9216,N_6875,N_6388);
nor U9217 (N_9217,N_7729,N_8380);
nand U9218 (N_9218,N_8370,N_8939);
nand U9219 (N_9219,N_7684,N_7378);
or U9220 (N_9220,N_6700,N_7203);
nor U9221 (N_9221,N_8131,N_7425);
or U9222 (N_9222,N_7356,N_6455);
nor U9223 (N_9223,N_6545,N_6272);
nor U9224 (N_9224,N_8817,N_7319);
nor U9225 (N_9225,N_6169,N_7857);
or U9226 (N_9226,N_6511,N_8402);
or U9227 (N_9227,N_6561,N_7986);
and U9228 (N_9228,N_6264,N_6826);
and U9229 (N_9229,N_6162,N_7061);
and U9230 (N_9230,N_6689,N_6610);
or U9231 (N_9231,N_8600,N_8120);
or U9232 (N_9232,N_8816,N_8762);
nand U9233 (N_9233,N_8986,N_7980);
or U9234 (N_9234,N_8744,N_7030);
nor U9235 (N_9235,N_6790,N_8702);
nor U9236 (N_9236,N_8125,N_7673);
and U9237 (N_9237,N_7265,N_8065);
and U9238 (N_9238,N_8767,N_7458);
and U9239 (N_9239,N_6173,N_7662);
nand U9240 (N_9240,N_6270,N_8830);
nor U9241 (N_9241,N_8397,N_7212);
and U9242 (N_9242,N_7320,N_8339);
xor U9243 (N_9243,N_7742,N_7472);
or U9244 (N_9244,N_6742,N_6143);
or U9245 (N_9245,N_8864,N_6380);
nand U9246 (N_9246,N_6608,N_8738);
xor U9247 (N_9247,N_8883,N_8977);
nor U9248 (N_9248,N_6766,N_7803);
and U9249 (N_9249,N_8596,N_6885);
nor U9250 (N_9250,N_8364,N_8984);
and U9251 (N_9251,N_7408,N_8433);
and U9252 (N_9252,N_8172,N_6214);
or U9253 (N_9253,N_8228,N_7674);
nand U9254 (N_9254,N_8287,N_8351);
or U9255 (N_9255,N_8871,N_7368);
nand U9256 (N_9256,N_8980,N_7748);
and U9257 (N_9257,N_6757,N_8466);
nand U9258 (N_9258,N_6690,N_7010);
or U9259 (N_9259,N_8569,N_7920);
or U9260 (N_9260,N_6282,N_6605);
or U9261 (N_9261,N_6473,N_6152);
nand U9262 (N_9262,N_6585,N_6497);
or U9263 (N_9263,N_6874,N_8302);
and U9264 (N_9264,N_8413,N_7241);
nor U9265 (N_9265,N_6295,N_7727);
nand U9266 (N_9266,N_6819,N_6112);
nand U9267 (N_9267,N_6000,N_7467);
or U9268 (N_9268,N_8821,N_6730);
nand U9269 (N_9269,N_8089,N_8211);
or U9270 (N_9270,N_8359,N_8462);
and U9271 (N_9271,N_8576,N_6258);
nand U9272 (N_9272,N_7562,N_8216);
and U9273 (N_9273,N_7694,N_6691);
or U9274 (N_9274,N_8145,N_8226);
and U9275 (N_9275,N_6831,N_6120);
nor U9276 (N_9276,N_8333,N_6913);
nand U9277 (N_9277,N_6213,N_8646);
and U9278 (N_9278,N_6255,N_8257);
or U9279 (N_9279,N_8690,N_8925);
nand U9280 (N_9280,N_8785,N_7627);
or U9281 (N_9281,N_7450,N_6904);
nor U9282 (N_9282,N_6568,N_7776);
nand U9283 (N_9283,N_6092,N_8367);
nor U9284 (N_9284,N_8079,N_8971);
nor U9285 (N_9285,N_8752,N_6711);
nor U9286 (N_9286,N_7309,N_8499);
or U9287 (N_9287,N_7655,N_6514);
nor U9288 (N_9288,N_7915,N_6571);
and U9289 (N_9289,N_7363,N_8115);
nor U9290 (N_9290,N_7515,N_8628);
xor U9291 (N_9291,N_6953,N_6212);
and U9292 (N_9292,N_8749,N_8255);
nor U9293 (N_9293,N_8360,N_6964);
and U9294 (N_9294,N_7336,N_7077);
or U9295 (N_9295,N_6257,N_8519);
or U9296 (N_9296,N_7365,N_7792);
nor U9297 (N_9297,N_7569,N_6911);
and U9298 (N_9298,N_8236,N_8698);
nand U9299 (N_9299,N_7974,N_8614);
or U9300 (N_9300,N_8373,N_6484);
and U9301 (N_9301,N_7377,N_7358);
or U9302 (N_9302,N_6077,N_7584);
and U9303 (N_9303,N_6801,N_6961);
or U9304 (N_9304,N_6719,N_7781);
nor U9305 (N_9305,N_8523,N_8340);
and U9306 (N_9306,N_6013,N_7848);
nand U9307 (N_9307,N_7107,N_7279);
nor U9308 (N_9308,N_7063,N_7016);
nor U9309 (N_9309,N_7788,N_8553);
and U9310 (N_9310,N_6475,N_8432);
or U9311 (N_9311,N_6684,N_7412);
and U9312 (N_9312,N_6829,N_6415);
nor U9313 (N_9313,N_6915,N_7297);
or U9314 (N_9314,N_8099,N_6124);
nand U9315 (N_9315,N_6402,N_6737);
and U9316 (N_9316,N_7303,N_6035);
nor U9317 (N_9317,N_6651,N_7955);
nor U9318 (N_9318,N_7631,N_8044);
or U9319 (N_9319,N_7110,N_8898);
nor U9320 (N_9320,N_6603,N_6108);
nand U9321 (N_9321,N_8197,N_7254);
nand U9322 (N_9322,N_8002,N_6144);
or U9323 (N_9323,N_6063,N_6852);
nand U9324 (N_9324,N_6187,N_7381);
or U9325 (N_9325,N_6688,N_6725);
and U9326 (N_9326,N_8497,N_7613);
or U9327 (N_9327,N_7238,N_8016);
nor U9328 (N_9328,N_7712,N_7386);
or U9329 (N_9329,N_8717,N_6098);
nand U9330 (N_9330,N_7052,N_8733);
nand U9331 (N_9331,N_8477,N_7518);
xor U9332 (N_9332,N_8107,N_7036);
nor U9333 (N_9333,N_7657,N_6088);
nor U9334 (N_9334,N_6816,N_8696);
nand U9335 (N_9335,N_8774,N_8886);
and U9336 (N_9336,N_6003,N_8138);
nand U9337 (N_9337,N_8989,N_6290);
and U9338 (N_9338,N_8347,N_8500);
nand U9339 (N_9339,N_8937,N_7460);
nand U9340 (N_9340,N_6623,N_6739);
or U9341 (N_9341,N_8531,N_6887);
and U9342 (N_9342,N_7186,N_6547);
nor U9343 (N_9343,N_8878,N_7162);
and U9344 (N_9344,N_7793,N_6007);
and U9345 (N_9345,N_7993,N_6425);
or U9346 (N_9346,N_8298,N_8195);
nand U9347 (N_9347,N_8742,N_8948);
nand U9348 (N_9348,N_6921,N_7201);
or U9349 (N_9349,N_6068,N_6136);
or U9350 (N_9350,N_8293,N_7286);
or U9351 (N_9351,N_6487,N_7181);
and U9352 (N_9352,N_8096,N_6049);
nand U9353 (N_9353,N_7221,N_8379);
or U9354 (N_9354,N_6268,N_8108);
or U9355 (N_9355,N_8437,N_6588);
and U9356 (N_9356,N_7886,N_6294);
nand U9357 (N_9357,N_8880,N_6667);
or U9358 (N_9358,N_6025,N_7455);
nand U9359 (N_9359,N_7660,N_6865);
nand U9360 (N_9360,N_8011,N_7661);
nor U9361 (N_9361,N_6232,N_6699);
and U9362 (N_9362,N_7233,N_7979);
and U9363 (N_9363,N_8231,N_8024);
nand U9364 (N_9364,N_8875,N_6909);
nand U9365 (N_9365,N_6544,N_6642);
nor U9366 (N_9366,N_8981,N_7017);
or U9367 (N_9367,N_7753,N_7076);
nand U9368 (N_9368,N_8486,N_7086);
nor U9369 (N_9369,N_7290,N_8181);
nor U9370 (N_9370,N_7038,N_8222);
or U9371 (N_9371,N_8641,N_7274);
nor U9372 (N_9372,N_6238,N_7713);
nand U9373 (N_9373,N_6955,N_8224);
nor U9374 (N_9374,N_7440,N_8771);
nand U9375 (N_9375,N_7987,N_7374);
or U9376 (N_9376,N_6115,N_6898);
and U9377 (N_9377,N_7600,N_7260);
or U9378 (N_9378,N_6093,N_6813);
and U9379 (N_9379,N_7605,N_8770);
and U9380 (N_9380,N_8516,N_6539);
or U9381 (N_9381,N_6582,N_7819);
and U9382 (N_9382,N_8853,N_6029);
nand U9383 (N_9383,N_7208,N_7456);
nand U9384 (N_9384,N_8826,N_7324);
and U9385 (N_9385,N_7642,N_6791);
nor U9386 (N_9386,N_6122,N_7405);
and U9387 (N_9387,N_7666,N_8084);
nand U9388 (N_9388,N_8192,N_8753);
nand U9389 (N_9389,N_8709,N_6401);
or U9390 (N_9390,N_8905,N_6998);
or U9391 (N_9391,N_8185,N_6387);
nor U9392 (N_9392,N_8847,N_6271);
nor U9393 (N_9393,N_8025,N_7114);
and U9394 (N_9394,N_7651,N_7182);
nand U9395 (N_9395,N_6593,N_6982);
nor U9396 (N_9396,N_8130,N_8617);
or U9397 (N_9397,N_8526,N_7092);
nand U9398 (N_9398,N_6460,N_8580);
nor U9399 (N_9399,N_6208,N_6104);
or U9400 (N_9400,N_6556,N_7098);
or U9401 (N_9401,N_7344,N_6428);
or U9402 (N_9402,N_7816,N_8321);
nor U9403 (N_9403,N_8759,N_7704);
xor U9404 (N_9404,N_7619,N_6260);
and U9405 (N_9405,N_7633,N_8388);
nand U9406 (N_9406,N_6211,N_8412);
nand U9407 (N_9407,N_8974,N_6024);
or U9408 (N_9408,N_6702,N_8304);
nand U9409 (N_9409,N_7766,N_6023);
and U9410 (N_9410,N_6969,N_8106);
or U9411 (N_9411,N_6782,N_7292);
nor U9412 (N_9412,N_8043,N_7723);
and U9413 (N_9413,N_8215,N_7861);
nand U9414 (N_9414,N_7205,N_7442);
and U9415 (N_9415,N_8054,N_8537);
nand U9416 (N_9416,N_7945,N_8545);
nor U9417 (N_9417,N_6970,N_6330);
nor U9418 (N_9418,N_6795,N_6550);
nand U9419 (N_9419,N_6515,N_6178);
nand U9420 (N_9420,N_6171,N_6789);
or U9421 (N_9421,N_8094,N_7207);
nand U9422 (N_9422,N_8327,N_7000);
nand U9423 (N_9423,N_7951,N_7659);
and U9424 (N_9424,N_8325,N_6351);
nor U9425 (N_9425,N_6778,N_7291);
and U9426 (N_9426,N_8885,N_6070);
nand U9427 (N_9427,N_8266,N_7983);
and U9428 (N_9428,N_6977,N_6762);
nand U9429 (N_9429,N_6718,N_7270);
and U9430 (N_9430,N_7751,N_6458);
nand U9431 (N_9431,N_7689,N_8001);
and U9432 (N_9432,N_8722,N_8863);
or U9433 (N_9433,N_8955,N_6553);
and U9434 (N_9434,N_8104,N_7722);
nor U9435 (N_9435,N_6233,N_7597);
nand U9436 (N_9436,N_7773,N_8559);
nor U9437 (N_9437,N_6518,N_6618);
nor U9438 (N_9438,N_6194,N_8095);
nand U9439 (N_9439,N_8563,N_6450);
nand U9440 (N_9440,N_7088,N_8322);
and U9441 (N_9441,N_8992,N_6454);
or U9442 (N_9442,N_7230,N_6659);
nand U9443 (N_9443,N_6466,N_8059);
nand U9444 (N_9444,N_7503,N_8842);
or U9445 (N_9445,N_6346,N_8303);
nor U9446 (N_9446,N_7759,N_6102);
or U9447 (N_9447,N_8672,N_6313);
and U9448 (N_9448,N_7498,N_7573);
and U9449 (N_9449,N_6564,N_6157);
nor U9450 (N_9450,N_7389,N_7040);
and U9451 (N_9451,N_7714,N_8438);
and U9452 (N_9452,N_7240,N_8010);
or U9453 (N_9453,N_6661,N_7954);
and U9454 (N_9454,N_7005,N_6918);
and U9455 (N_9455,N_7591,N_6525);
nor U9456 (N_9456,N_6884,N_8184);
nor U9457 (N_9457,N_7497,N_6530);
and U9458 (N_9458,N_7916,N_8912);
or U9459 (N_9459,N_6595,N_8270);
nand U9460 (N_9460,N_8417,N_8209);
or U9461 (N_9461,N_7822,N_6950);
or U9462 (N_9462,N_6328,N_6041);
nand U9463 (N_9463,N_6109,N_6249);
or U9464 (N_9464,N_8376,N_6573);
and U9465 (N_9465,N_7148,N_7438);
nand U9466 (N_9466,N_8418,N_8611);
nor U9467 (N_9467,N_7109,N_6720);
nor U9468 (N_9468,N_7117,N_7200);
and U9469 (N_9469,N_6442,N_7012);
and U9470 (N_9470,N_8103,N_8126);
or U9471 (N_9471,N_8355,N_6732);
nand U9472 (N_9472,N_6096,N_6301);
or U9473 (N_9473,N_7982,N_6685);
and U9474 (N_9474,N_6936,N_8392);
nor U9475 (N_9475,N_6783,N_6371);
nor U9476 (N_9476,N_6523,N_8341);
nor U9477 (N_9477,N_6203,N_7170);
nand U9478 (N_9478,N_7859,N_6847);
or U9479 (N_9479,N_8009,N_8943);
or U9480 (N_9480,N_8015,N_8916);
and U9481 (N_9481,N_8336,N_7404);
and U9482 (N_9482,N_7553,N_8495);
nand U9483 (N_9483,N_6599,N_8071);
nor U9484 (N_9484,N_8252,N_6147);
or U9485 (N_9485,N_6446,N_6644);
and U9486 (N_9486,N_6137,N_6360);
nand U9487 (N_9487,N_7820,N_6471);
nor U9488 (N_9488,N_7738,N_7006);
nor U9489 (N_9489,N_8451,N_6731);
nand U9490 (N_9490,N_8259,N_8729);
or U9491 (N_9491,N_6195,N_7024);
nand U9492 (N_9492,N_8242,N_6532);
and U9493 (N_9493,N_7736,N_7037);
nor U9494 (N_9494,N_7896,N_7508);
nor U9495 (N_9495,N_6072,N_6155);
and U9496 (N_9496,N_6758,N_7403);
and U9497 (N_9497,N_6225,N_7846);
and U9498 (N_9498,N_8278,N_8697);
and U9499 (N_9499,N_6704,N_8182);
and U9500 (N_9500,N_8876,N_6733);
and U9501 (N_9501,N_6990,N_6598);
nor U9502 (N_9502,N_8283,N_8204);
and U9503 (N_9503,N_6975,N_7635);
nand U9504 (N_9504,N_6337,N_8154);
and U9505 (N_9505,N_6498,N_7176);
nor U9506 (N_9506,N_8795,N_7681);
and U9507 (N_9507,N_6892,N_7042);
or U9508 (N_9508,N_6449,N_6840);
nand U9509 (N_9509,N_8112,N_6075);
nand U9510 (N_9510,N_6748,N_6891);
nand U9511 (N_9511,N_8487,N_7191);
nand U9512 (N_9512,N_6105,N_7225);
and U9513 (N_9513,N_8346,N_7343);
or U9514 (N_9514,N_8538,N_6496);
or U9515 (N_9515,N_7087,N_7457);
or U9516 (N_9516,N_8299,N_6400);
nand U9517 (N_9517,N_8217,N_7294);
and U9518 (N_9518,N_6995,N_8055);
nand U9519 (N_9519,N_6151,N_7009);
nor U9520 (N_9520,N_7544,N_6634);
nor U9521 (N_9521,N_6193,N_6914);
or U9522 (N_9522,N_8721,N_7774);
and U9523 (N_9523,N_6763,N_7502);
nand U9524 (N_9524,N_8615,N_8845);
and U9525 (N_9525,N_8329,N_8053);
nor U9526 (N_9526,N_6119,N_6237);
nand U9527 (N_9527,N_7501,N_7026);
or U9528 (N_9528,N_8394,N_8887);
and U9529 (N_9529,N_6528,N_6770);
nand U9530 (N_9530,N_7810,N_6129);
nor U9531 (N_9531,N_8160,N_6321);
and U9532 (N_9532,N_6067,N_6551);
nand U9533 (N_9533,N_6786,N_8513);
or U9534 (N_9534,N_6494,N_8711);
nand U9535 (N_9535,N_7008,N_8165);
and U9536 (N_9536,N_6296,N_6849);
and U9537 (N_9537,N_7807,N_7546);
nand U9538 (N_9538,N_8448,N_7224);
or U9539 (N_9539,N_8718,N_8603);
or U9540 (N_9540,N_8268,N_7519);
nand U9541 (N_9541,N_8756,N_6161);
or U9542 (N_9542,N_6389,N_8076);
and U9543 (N_9543,N_8870,N_7787);
nand U9544 (N_9544,N_8331,N_7454);
or U9545 (N_9545,N_7091,N_7145);
nand U9546 (N_9546,N_8802,N_7430);
and U9547 (N_9547,N_6645,N_7004);
or U9548 (N_9548,N_7174,N_8174);
nand U9549 (N_9549,N_7620,N_8369);
nand U9550 (N_9550,N_8528,N_6750);
and U9551 (N_9551,N_7478,N_8033);
nand U9552 (N_9552,N_8384,N_6846);
and U9553 (N_9553,N_7206,N_7865);
xor U9554 (N_9554,N_8828,N_8052);
nand U9555 (N_9555,N_6615,N_8244);
nand U9556 (N_9556,N_6489,N_8930);
nand U9557 (N_9557,N_7589,N_8901);
nor U9558 (N_9558,N_8743,N_8913);
and U9559 (N_9559,N_8631,N_6591);
and U9560 (N_9560,N_7175,N_8703);
or U9561 (N_9561,N_8368,N_7171);
or U9562 (N_9562,N_6584,N_6499);
and U9563 (N_9563,N_6170,N_7255);
nor U9564 (N_9564,N_8798,N_6792);
nand U9565 (N_9565,N_7603,N_6174);
and U9566 (N_9566,N_6678,N_8868);
nor U9567 (N_9567,N_8097,N_7161);
nor U9568 (N_9568,N_7461,N_6148);
nor U9569 (N_9569,N_7420,N_6039);
and U9570 (N_9570,N_8291,N_7594);
and U9571 (N_9571,N_6369,N_8088);
and U9572 (N_9572,N_7708,N_8365);
and U9573 (N_9573,N_6386,N_6996);
nand U9574 (N_9574,N_6121,N_7090);
nor U9575 (N_9575,N_7326,N_7124);
nand U9576 (N_9576,N_6492,N_7789);
nor U9577 (N_9577,N_7898,N_8423);
xnor U9578 (N_9578,N_8503,N_7801);
nor U9579 (N_9579,N_7147,N_7976);
nand U9580 (N_9580,N_7141,N_6417);
or U9581 (N_9581,N_8452,N_7588);
or U9582 (N_9582,N_6243,N_7180);
nand U9583 (N_9583,N_7778,N_7720);
or U9584 (N_9584,N_8143,N_7625);
nor U9585 (N_9585,N_8900,N_6929);
or U9586 (N_9586,N_7877,N_6663);
or U9587 (N_9587,N_6827,N_7130);
nor U9588 (N_9588,N_7602,N_7812);
and U9589 (N_9589,N_8383,N_6721);
and U9590 (N_9590,N_8246,N_7464);
and U9591 (N_9591,N_7650,N_8858);
and U9592 (N_9592,N_6540,N_6633);
nor U9593 (N_9593,N_7592,N_7385);
or U9594 (N_9594,N_8998,N_8619);
nand U9595 (N_9595,N_7718,N_7728);
nor U9596 (N_9596,N_7685,N_8401);
or U9597 (N_9597,N_6992,N_8841);
nand U9598 (N_9598,N_8642,N_6601);
and U9599 (N_9599,N_6114,N_7818);
and U9600 (N_9600,N_7178,N_6421);
and U9601 (N_9601,N_7539,N_8080);
nor U9602 (N_9602,N_6131,N_6756);
nand U9603 (N_9603,N_8620,N_8789);
nand U9604 (N_9604,N_7608,N_7990);
or U9605 (N_9605,N_8443,N_8377);
nor U9606 (N_9606,N_8621,N_8823);
nor U9607 (N_9607,N_7298,N_8350);
and U9608 (N_9608,N_8150,N_6278);
nand U9609 (N_9609,N_8429,N_6201);
and U9610 (N_9610,N_6920,N_8966);
and U9611 (N_9611,N_7977,N_6299);
and U9612 (N_9612,N_6834,N_7134);
and U9613 (N_9613,N_8540,N_7105);
and U9614 (N_9614,N_7599,N_7901);
or U9615 (N_9615,N_7832,N_7376);
nor U9616 (N_9616,N_6513,N_7287);
nand U9617 (N_9617,N_8610,N_8430);
nand U9618 (N_9618,N_6452,N_6416);
nand U9619 (N_9619,N_8245,N_8419);
or U9620 (N_9620,N_6639,N_8403);
and U9621 (N_9621,N_7209,N_8907);
xnor U9622 (N_9622,N_7471,N_7841);
nand U9623 (N_9623,N_8190,N_6247);
nor U9624 (N_9624,N_6246,N_7910);
or U9625 (N_9625,N_7253,N_8896);
or U9626 (N_9626,N_8155,N_8110);
or U9627 (N_9627,N_7222,N_6329);
or U9628 (N_9628,N_7734,N_8969);
nor U9629 (N_9629,N_6310,N_6004);
or U9630 (N_9630,N_7882,N_8651);
nand U9631 (N_9631,N_6046,N_7571);
nand U9632 (N_9632,N_6962,N_6680);
nor U9633 (N_9633,N_6315,N_8146);
and U9634 (N_9634,N_6375,N_7880);
nand U9635 (N_9635,N_8658,N_6987);
and U9636 (N_9636,N_6753,N_6188);
nor U9637 (N_9637,N_7187,N_7814);
nand U9638 (N_9638,N_7839,N_8127);
nand U9639 (N_9639,N_8085,N_8157);
or U9640 (N_9640,N_6785,N_6062);
and U9641 (N_9641,N_6307,N_8758);
or U9642 (N_9642,N_8748,N_8454);
nor U9643 (N_9643,N_7071,N_8685);
nand U9644 (N_9644,N_6769,N_8116);
or U9645 (N_9645,N_8787,N_6056);
and U9646 (N_9646,N_6776,N_6283);
or U9647 (N_9647,N_7889,N_6297);
and U9648 (N_9648,N_6226,N_8295);
and U9649 (N_9649,N_6717,N_8311);
or U9650 (N_9650,N_6705,N_8300);
and U9651 (N_9651,N_8070,N_7561);
or U9652 (N_9652,N_6860,N_7850);
nor U9653 (N_9653,N_6926,N_6937);
and U9654 (N_9654,N_7022,N_8170);
nand U9655 (N_9655,N_7407,N_7530);
nor U9656 (N_9656,N_8923,N_8194);
nand U9657 (N_9657,N_6111,N_7237);
nor U9658 (N_9658,N_6587,N_8189);
nand U9659 (N_9659,N_6822,N_7449);
and U9660 (N_9660,N_8488,N_8834);
nor U9661 (N_9661,N_7654,N_6177);
nand U9662 (N_9662,N_7513,N_8203);
and U9663 (N_9663,N_8532,N_6646);
and U9664 (N_9664,N_6230,N_7721);
and U9665 (N_9665,N_6158,N_7551);
nand U9666 (N_9666,N_8221,N_6261);
or U9667 (N_9667,N_6787,N_7784);
nor U9668 (N_9668,N_8637,N_6657);
nand U9669 (N_9669,N_7785,N_6845);
nand U9670 (N_9670,N_8700,N_7428);
or U9671 (N_9671,N_6542,N_6818);
nand U9672 (N_9672,N_8038,N_7261);
or U9673 (N_9673,N_7572,N_7434);
and U9674 (N_9674,N_7731,N_7695);
or U9675 (N_9675,N_7463,N_8414);
and U9676 (N_9676,N_8725,N_8904);
or U9677 (N_9677,N_7582,N_6420);
or U9678 (N_9678,N_6590,N_8320);
and U9679 (N_9679,N_8550,N_8684);
or U9680 (N_9680,N_7823,N_7649);
nand U9681 (N_9681,N_6621,N_7996);
or U9682 (N_9682,N_7964,N_6729);
nor U9683 (N_9683,N_8612,N_7872);
and U9684 (N_9684,N_7433,N_8965);
or U9685 (N_9685,N_6668,N_7830);
nand U9686 (N_9686,N_7179,N_7640);
nand U9687 (N_9687,N_7334,N_8578);
or U9688 (N_9688,N_8018,N_6882);
nor U9689 (N_9689,N_6200,N_6311);
and U9690 (N_9690,N_8661,N_8308);
nand U9691 (N_9691,N_7900,N_7874);
nand U9692 (N_9692,N_8098,N_8249);
nor U9693 (N_9693,N_8353,N_6896);
nor U9694 (N_9694,N_8564,N_6106);
nand U9695 (N_9695,N_8958,N_7413);
nand U9696 (N_9696,N_8093,N_8942);
nor U9697 (N_9697,N_6527,N_7570);
or U9698 (N_9698,N_6139,N_7581);
or U9699 (N_9699,N_8400,N_8807);
nor U9700 (N_9700,N_8769,N_6010);
or U9701 (N_9701,N_8666,N_7645);
nor U9702 (N_9702,N_8214,N_8472);
nand U9703 (N_9703,N_6113,N_6900);
or U9704 (N_9704,N_8827,N_7128);
and U9705 (N_9705,N_6622,N_7550);
nand U9706 (N_9706,N_8917,N_7735);
nor U9707 (N_9707,N_8358,N_8129);
nand U9708 (N_9708,N_7150,N_6957);
nor U9709 (N_9709,N_8393,N_7909);
or U9710 (N_9710,N_8835,N_8069);
nand U9711 (N_9711,N_6447,N_7223);
nor U9712 (N_9712,N_8483,N_8133);
or U9713 (N_9713,N_7887,N_8994);
or U9714 (N_9714,N_6838,N_6231);
or U9715 (N_9715,N_7676,N_6537);
or U9716 (N_9716,N_7963,N_6347);
nand U9717 (N_9717,N_6435,N_6060);
nor U9718 (N_9718,N_6284,N_8316);
nor U9719 (N_9719,N_7095,N_7577);
nor U9720 (N_9720,N_7969,N_7172);
or U9721 (N_9721,N_8306,N_7538);
nor U9722 (N_9722,N_8229,N_8933);
and U9723 (N_9723,N_8186,N_7229);
nand U9724 (N_9724,N_7629,N_6620);
and U9725 (N_9725,N_7422,N_8679);
and U9726 (N_9726,N_7406,N_7772);
nor U9727 (N_9727,N_8525,N_7509);
xor U9728 (N_9728,N_7249,N_8114);
and U9729 (N_9729,N_6531,N_6383);
and U9730 (N_9730,N_8288,N_8471);
nor U9731 (N_9731,N_7780,N_8381);
or U9732 (N_9732,N_6519,N_7913);
or U9733 (N_9733,N_7393,N_7575);
nand U9734 (N_9734,N_7384,N_6412);
nor U9735 (N_9735,N_6501,N_8225);
or U9736 (N_9736,N_6609,N_7690);
and U9737 (N_9737,N_6026,N_8465);
nor U9738 (N_9738,N_8456,N_8349);
nand U9739 (N_9739,N_6305,N_7540);
nor U9740 (N_9740,N_7590,N_8223);
nor U9741 (N_9741,N_7232,N_7424);
nor U9742 (N_9742,N_8374,N_6794);
or U9743 (N_9743,N_6303,N_8382);
nor U9744 (N_9744,N_6128,N_6456);
and U9745 (N_9745,N_6125,N_8344);
or U9746 (N_9746,N_7907,N_8064);
or U9747 (N_9747,N_7198,N_8701);
nand U9748 (N_9748,N_7099,N_6746);
and U9749 (N_9749,N_7429,N_8585);
nand U9750 (N_9750,N_6883,N_8968);
or U9751 (N_9751,N_7940,N_6095);
nand U9752 (N_9752,N_7398,N_8027);
or U9753 (N_9753,N_6919,N_8136);
or U9754 (N_9754,N_6474,N_8567);
nor U9755 (N_9755,N_8045,N_8371);
nor U9756 (N_9756,N_6981,N_6805);
nand U9757 (N_9757,N_7112,N_7474);
nor U9758 (N_9758,N_6722,N_7275);
nor U9759 (N_9759,N_7014,N_7257);
and U9760 (N_9760,N_8775,N_6419);
and U9761 (N_9761,N_6850,N_8979);
nand U9762 (N_9762,N_6516,N_6967);
or U9763 (N_9763,N_8793,N_7447);
and U9764 (N_9764,N_6752,N_6710);
nor U9765 (N_9765,N_7939,N_6679);
and U9766 (N_9766,N_8275,N_6482);
nor U9767 (N_9767,N_6107,N_8473);
or U9768 (N_9768,N_8305,N_6916);
nor U9769 (N_9769,N_7614,N_6985);
nand U9770 (N_9770,N_6559,N_8476);
nand U9771 (N_9771,N_6319,N_6485);
nor U9772 (N_9772,N_7189,N_8688);
nand U9773 (N_9773,N_6138,N_6325);
nand U9774 (N_9774,N_7018,N_8613);
or U9775 (N_9775,N_7504,N_6433);
or U9776 (N_9776,N_7444,N_8493);
nand U9777 (N_9777,N_6451,N_6159);
nand U9778 (N_9778,N_6335,N_8261);
or U9779 (N_9779,N_6828,N_6069);
nor U9780 (N_9780,N_6839,N_8294);
nor U9781 (N_9781,N_7946,N_8586);
or U9782 (N_9782,N_8623,N_8634);
and U9783 (N_9783,N_7045,N_6648);
nor U9784 (N_9784,N_6788,N_8135);
nand U9785 (N_9785,N_6229,N_7596);
nand U9786 (N_9786,N_6989,N_7258);
or U9787 (N_9787,N_6858,N_7416);
and U9788 (N_9788,N_7871,N_8664);
nand U9789 (N_9789,N_6265,N_7745);
or U9790 (N_9790,N_7388,N_8241);
and U9791 (N_9791,N_6160,N_7419);
nand U9792 (N_9792,N_8238,N_8092);
nor U9793 (N_9793,N_7085,N_6592);
and U9794 (N_9794,N_8285,N_8468);
and U9795 (N_9795,N_7056,N_6085);
nor U9796 (N_9796,N_6087,N_7154);
nor U9797 (N_9797,N_7563,N_7299);
nor U9798 (N_9798,N_6676,N_8062);
nand U9799 (N_9799,N_7029,N_8056);
and U9800 (N_9800,N_7401,N_7934);
nor U9801 (N_9801,N_8023,N_7195);
nor U9802 (N_9802,N_6653,N_7342);
nor U9803 (N_9803,N_6465,N_6627);
or U9804 (N_9804,N_8233,N_8256);
or U9805 (N_9805,N_6535,N_8843);
nor U9806 (N_9806,N_7436,N_8601);
nand U9807 (N_9807,N_8897,N_6481);
xor U9808 (N_9808,N_6097,N_7931);
or U9809 (N_9809,N_7824,N_8978);
nor U9810 (N_9810,N_7585,N_6745);
or U9811 (N_9811,N_8004,N_7267);
and U9812 (N_9812,N_7521,N_7360);
nand U9813 (N_9813,N_6677,N_7400);
nand U9814 (N_9814,N_6228,N_8398);
nor U9815 (N_9815,N_6326,N_6281);
nand U9816 (N_9816,N_7680,N_8188);
or U9817 (N_9817,N_7337,N_6761);
nand U9818 (N_9818,N_6398,N_8041);
nand U9819 (N_9819,N_6480,N_6814);
or U9820 (N_9820,N_8101,N_6191);
or U9821 (N_9821,N_7248,N_6538);
and U9822 (N_9822,N_8334,N_7242);
nand U9823 (N_9823,N_7122,N_7157);
and U9824 (N_9824,N_8909,N_6666);
or U9825 (N_9825,N_6972,N_6457);
nand U9826 (N_9826,N_7228,N_8218);
or U9827 (N_9827,N_6476,N_6304);
nand U9828 (N_9828,N_8987,N_6954);
and U9829 (N_9829,N_7192,N_8940);
nand U9830 (N_9830,N_6488,N_6500);
nand U9831 (N_9831,N_8319,N_8482);
and U9832 (N_9832,N_6015,N_8645);
nand U9833 (N_9833,N_7892,N_7794);
nor U9834 (N_9834,N_7707,N_7764);
nand U9835 (N_9835,N_6759,N_6202);
and U9836 (N_9836,N_7295,N_8490);
and U9837 (N_9837,N_6712,N_8797);
or U9838 (N_9838,N_6974,N_8134);
nand U9839 (N_9839,N_8741,N_8995);
nand U9840 (N_9840,N_8492,N_6709);
nand U9841 (N_9841,N_6660,N_6886);
nor U9842 (N_9842,N_8511,N_7641);
nand U9843 (N_9843,N_8582,N_6692);
nor U9844 (N_9844,N_6800,N_7484);
or U9845 (N_9845,N_6332,N_6640);
nor U9846 (N_9846,N_7311,N_6505);
nand U9847 (N_9847,N_8424,N_7851);
nand U9848 (N_9848,N_6552,N_7579);
nor U9849 (N_9849,N_6406,N_8906);
and U9850 (N_9850,N_7329,N_8102);
nand U9851 (N_9851,N_8020,N_8985);
nor U9852 (N_9852,N_7397,N_7069);
or U9853 (N_9853,N_8142,N_8144);
or U9854 (N_9854,N_7396,N_8768);
or U9855 (N_9855,N_8464,N_6873);
nand U9856 (N_9856,N_8599,N_8618);
nor U9857 (N_9857,N_7574,N_7480);
nand U9858 (N_9858,N_7204,N_8952);
nand U9859 (N_9859,N_7506,N_8404);
and U9860 (N_9860,N_8993,N_7220);
nand U9861 (N_9861,N_6033,N_8505);
and U9862 (N_9862,N_7379,N_7606);
xor U9863 (N_9863,N_7153,N_7806);
nand U9864 (N_9864,N_8235,N_8180);
nor U9865 (N_9865,N_7074,N_8003);
nor U9866 (N_9866,N_7417,N_6868);
and U9867 (N_9867,N_7558,N_6510);
or U9868 (N_9868,N_7636,N_6293);
and U9869 (N_9869,N_7485,N_7717);
nand U9870 (N_9870,N_6793,N_6244);
nor U9871 (N_9871,N_6566,N_6110);
and U9872 (N_9872,N_8363,N_8077);
nor U9873 (N_9873,N_8924,N_8663);
and U9874 (N_9874,N_7490,N_8824);
nand U9875 (N_9875,N_8177,N_7125);
xor U9876 (N_9876,N_6872,N_8988);
nor U9877 (N_9877,N_7533,N_7055);
or U9878 (N_9878,N_8021,N_8441);
nand U9879 (N_9879,N_7421,N_6765);
or U9880 (N_9880,N_7043,N_7507);
nor U9881 (N_9881,N_7120,N_8447);
or U9882 (N_9882,N_7139,N_7843);
and U9883 (N_9883,N_8812,N_8029);
nand U9884 (N_9884,N_7372,N_8608);
nand U9885 (N_9885,N_8048,N_7760);
nor U9886 (N_9886,N_8669,N_7317);
or U9887 (N_9887,N_7361,N_6945);
or U9888 (N_9888,N_8345,N_8338);
nor U9889 (N_9889,N_8292,N_7330);
nand U9890 (N_9890,N_7348,N_6563);
nand U9891 (N_9891,N_7470,N_8683);
or U9892 (N_9892,N_6254,N_7683);
and U9893 (N_9893,N_7643,N_7885);
and U9894 (N_9894,N_7984,N_6851);
and U9895 (N_9895,N_6811,N_8362);
or U9896 (N_9896,N_6083,N_8975);
and U9897 (N_9897,N_6262,N_8957);
nand U9898 (N_9898,N_7352,N_6289);
nor U9899 (N_9899,N_8786,N_8882);
nand U9900 (N_9900,N_6825,N_6391);
or U9901 (N_9901,N_7219,N_6560);
or U9902 (N_9902,N_7500,N_7362);
and U9903 (N_9903,N_6291,N_6643);
nor U9904 (N_9904,N_7366,N_7798);
nand U9905 (N_9905,N_6880,N_6754);
and U9906 (N_9906,N_7493,N_6123);
or U9907 (N_9907,N_6145,N_7335);
nand U9908 (N_9908,N_7264,N_6901);
nand U9909 (N_9909,N_6889,N_7699);
nand U9910 (N_9910,N_8391,N_6422);
or U9911 (N_9911,N_7073,N_6001);
nand U9912 (N_9912,N_8202,N_7517);
and U9913 (N_9913,N_6799,N_8594);
and U9914 (N_9914,N_6844,N_7019);
and U9915 (N_9915,N_7639,N_6073);
and U9916 (N_9916,N_8522,N_8638);
and U9917 (N_9917,N_7338,N_7536);
nand U9918 (N_9918,N_8670,N_6772);
nor U9919 (N_9919,N_8489,N_8699);
nor U9920 (N_9920,N_6771,N_6773);
and U9921 (N_9921,N_7155,N_7210);
or U9922 (N_9922,N_7060,N_7138);
and U9923 (N_9923,N_8946,N_6267);
or U9924 (N_9924,N_7051,N_8574);
nor U9925 (N_9925,N_8794,N_8809);
nand U9926 (N_9926,N_6978,N_7475);
and U9927 (N_9927,N_7709,N_7160);
nand U9928 (N_9928,N_7663,N_7529);
xnor U9929 (N_9929,N_8518,N_6820);
nor U9930 (N_9930,N_7947,N_8091);
nand U9931 (N_9931,N_6036,N_8595);
and U9932 (N_9932,N_6166,N_6506);
or U9933 (N_9933,N_6747,N_7115);
and U9934 (N_9934,N_6164,N_8328);
or U9935 (N_9935,N_7312,N_7131);
or U9936 (N_9936,N_6628,N_6963);
nand U9937 (N_9937,N_7564,N_8982);
and U9938 (N_9938,N_7096,N_7252);
nor U9939 (N_9939,N_8406,N_6344);
nor U9940 (N_9940,N_7541,N_8008);
and U9941 (N_9941,N_6939,N_7834);
nor U9942 (N_9942,N_7761,N_7215);
nand U9943 (N_9943,N_7786,N_6440);
or U9944 (N_9944,N_7956,N_7321);
nand U9945 (N_9945,N_8764,N_8529);
and U9946 (N_9946,N_6577,N_7904);
nor U9947 (N_9947,N_6459,N_8141);
nor U9948 (N_9948,N_8199,N_6888);
or U9949 (N_9949,N_6118,N_6522);
nand U9950 (N_9950,N_6279,N_7838);
and U9951 (N_9951,N_7218,N_6495);
or U9952 (N_9952,N_7300,N_6673);
and U9953 (N_9953,N_8686,N_8449);
and U9954 (N_9954,N_6463,N_7064);
nor U9955 (N_9955,N_8169,N_8932);
or U9956 (N_9956,N_6812,N_7243);
and U9957 (N_9957,N_8039,N_6935);
nand U9958 (N_9958,N_8357,N_7879);
and U9959 (N_9959,N_7711,N_8148);
and U9960 (N_9960,N_8678,N_8544);
or U9961 (N_9961,N_8874,N_6382);
nand U9962 (N_9962,N_7236,N_8277);
nand U9963 (N_9963,N_7325,N_6091);
nor U9964 (N_9964,N_6234,N_8475);
and U9965 (N_9965,N_7118,N_7646);
and U9966 (N_9966,N_7094,N_8361);
nor U9967 (N_9967,N_6965,N_7146);
and U9968 (N_9968,N_6210,N_8680);
and U9969 (N_9969,N_6616,N_8395);
nand U9970 (N_9970,N_8149,N_8571);
nor U9971 (N_9971,N_8167,N_6052);
nor U9972 (N_9972,N_6681,N_7545);
nor U9973 (N_9973,N_6245,N_6438);
nor U9974 (N_9974,N_8100,N_6248);
nor U9975 (N_9975,N_7754,N_7281);
nand U9976 (N_9976,N_6669,N_8919);
and U9977 (N_9977,N_8479,N_8761);
nand U9978 (N_9978,N_8230,N_8390);
nand U9979 (N_9979,N_7520,N_8072);
nor U9980 (N_9980,N_6012,N_7345);
nand U9981 (N_9981,N_8440,N_6486);
nand U9982 (N_9982,N_6378,N_7196);
nor U9983 (N_9983,N_6629,N_6695);
nand U9984 (N_9984,N_8058,N_7266);
nand U9985 (N_9985,N_7847,N_6817);
nor U9986 (N_9986,N_8137,N_7383);
nor U9987 (N_9987,N_7855,N_8271);
or U9988 (N_9988,N_8579,N_8746);
or U9989 (N_9989,N_7692,N_7853);
or U9990 (N_9990,N_7364,N_7998);
nor U9991 (N_9991,N_7426,N_6302);
nand U9992 (N_9992,N_8416,N_7938);
and U9993 (N_9993,N_8314,N_8124);
or U9994 (N_9994,N_7048,N_6403);
nand U9995 (N_9995,N_8872,N_8282);
nor U9996 (N_9996,N_8593,N_7523);
nand U9997 (N_9997,N_7282,N_8627);
and U9998 (N_9998,N_7893,N_7876);
nor U9999 (N_9999,N_6986,N_8446);
or U10000 (N_10000,N_6938,N_7604);
nand U10001 (N_10001,N_8839,N_8163);
or U10002 (N_10002,N_6855,N_7268);
nor U10003 (N_10003,N_6028,N_8808);
nor U10004 (N_10004,N_8587,N_8407);
nand U10005 (N_10005,N_8307,N_8309);
nand U10006 (N_10006,N_8534,N_8504);
nor U10007 (N_10007,N_7067,N_7653);
nor U10008 (N_10008,N_6285,N_8649);
xnor U10009 (N_10009,N_6130,N_6768);
nor U10010 (N_10010,N_6367,N_6924);
nand U10011 (N_10011,N_8557,N_8310);
or U10012 (N_10012,N_8175,N_7486);
nor U10013 (N_10013,N_6053,N_8467);
and U10014 (N_10014,N_7985,N_6833);
nand U10015 (N_10015,N_8861,N_6625);
nand U10016 (N_10016,N_7483,N_7246);
nor U10017 (N_10017,N_7058,N_8941);
and U10018 (N_10018,N_6876,N_8708);
and U10019 (N_10019,N_8173,N_7870);
nand U10020 (N_10020,N_7328,N_6508);
or U10021 (N_10021,N_7644,N_8090);
or U10022 (N_10022,N_7669,N_8755);
and U10023 (N_10023,N_8535,N_6810);
nor U10024 (N_10024,N_8822,N_6205);
nand U10025 (N_10025,N_7556,N_8778);
and U10026 (N_10026,N_6071,N_7262);
and U10027 (N_10027,N_6156,N_8026);
and U10028 (N_10028,N_6365,N_6076);
nand U10029 (N_10029,N_6142,N_7973);
and U10030 (N_10030,N_7747,N_8675);
nor U10031 (N_10031,N_7354,N_6019);
and U10032 (N_10032,N_8713,N_7035);
nand U10033 (N_10033,N_7696,N_8012);
or U10034 (N_10034,N_8899,N_7912);
nor U10035 (N_10035,N_6517,N_6395);
and U10036 (N_10036,N_8687,N_6557);
and U10037 (N_10037,N_8542,N_8682);
and U10038 (N_10038,N_6674,N_7868);
and U10039 (N_10039,N_7367,N_6477);
or U10040 (N_10040,N_7341,N_6453);
nand U10041 (N_10041,N_6089,N_7031);
nor U10042 (N_10042,N_8066,N_7488);
or U10043 (N_10043,N_7932,N_8415);
nor U10044 (N_10044,N_6370,N_6209);
nand U10045 (N_10045,N_7716,N_6005);
or U10046 (N_10046,N_6241,N_6971);
nand U10047 (N_10047,N_7802,N_8857);
nor U10048 (N_10048,N_8991,N_8805);
nor U10049 (N_10049,N_7173,N_8196);
and U10050 (N_10050,N_8068,N_6443);
and U10051 (N_10051,N_8028,N_8840);
or U10052 (N_10052,N_8337,N_7897);
and U10053 (N_10053,N_6084,N_8859);
nand U10054 (N_10054,N_7809,N_8105);
and U10055 (N_10055,N_7235,N_7102);
or U10056 (N_10056,N_7331,N_6856);
or U10057 (N_10057,N_8515,N_8660);
or U10058 (N_10058,N_8207,N_7050);
nand U10059 (N_10059,N_7284,N_6686);
and U10060 (N_10060,N_8042,N_8735);
or U10061 (N_10061,N_8591,N_6988);
nor U10062 (N_10062,N_8366,N_7836);
nor U10063 (N_10063,N_7813,N_7027);
or U10064 (N_10064,N_7020,N_8605);
or U10065 (N_10065,N_6979,N_6366);
or U10066 (N_10066,N_7340,N_6871);
nor U10067 (N_10067,N_7492,N_7479);
nand U10068 (N_10068,N_8644,N_7840);
or U10069 (N_10069,N_8198,N_8434);
nor U10070 (N_10070,N_7908,N_6256);
nor U10071 (N_10071,N_6809,N_6764);
nand U10072 (N_10072,N_7740,N_6861);
and U10073 (N_10073,N_6292,N_6038);
nor U10074 (N_10074,N_6057,N_7583);
nor U10075 (N_10075,N_6064,N_8855);
or U10076 (N_10076,N_6502,N_7559);
or U10077 (N_10077,N_8022,N_7247);
or U10078 (N_10078,N_6879,N_8014);
and U10079 (N_10079,N_7927,N_8286);
nor U10080 (N_10080,N_6617,N_8598);
or U10081 (N_10081,N_8671,N_8264);
and U10082 (N_10082,N_6807,N_7231);
nor U10083 (N_10083,N_8655,N_7380);
xnor U10084 (N_10084,N_6802,N_8653);
nor U10085 (N_10085,N_6361,N_8031);
and U10086 (N_10086,N_6672,N_7768);
nor U10087 (N_10087,N_6952,N_6065);
nand U10088 (N_10088,N_7902,N_6217);
nand U10089 (N_10089,N_6665,N_8918);
or U10090 (N_10090,N_8243,N_6696);
or U10091 (N_10091,N_7250,N_7202);
nor U10092 (N_10092,N_6774,N_6192);
nand U10093 (N_10093,N_8773,N_8606);
nor U10094 (N_10094,N_8740,N_7158);
or U10095 (N_10095,N_7567,N_8691);
nor U10096 (N_10096,N_7482,N_6509);
and U10097 (N_10097,N_8086,N_7678);
or U10098 (N_10098,N_6655,N_8654);
nor U10099 (N_10099,N_6682,N_8908);
nand U10100 (N_10100,N_8356,N_6912);
or U10101 (N_10101,N_6334,N_8934);
nor U10102 (N_10102,N_8629,N_7059);
and U10103 (N_10103,N_6222,N_6751);
or U10104 (N_10104,N_8556,N_7423);
nand U10105 (N_10105,N_6687,N_6385);
or U10106 (N_10106,N_7962,N_6020);
or U10107 (N_10107,N_8113,N_8630);
nand U10108 (N_10108,N_8332,N_6931);
nand U10109 (N_10109,N_7890,N_7970);
and U10110 (N_10110,N_6958,N_6675);
or U10111 (N_10111,N_7844,N_6701);
nand U10112 (N_10112,N_7477,N_6140);
or U10113 (N_10113,N_6048,N_6777);
or U10114 (N_10114,N_6153,N_6549);
or U10115 (N_10115,N_7116,N_7526);
or U10116 (N_10116,N_8067,N_7568);
xor U10117 (N_10117,N_6204,N_6944);
nor U10118 (N_10118,N_8552,N_8757);
or U10119 (N_10119,N_8652,N_7856);
xor U10120 (N_10120,N_7686,N_7156);
nor U10121 (N_10121,N_7011,N_7041);
and U10122 (N_10122,N_6078,N_6478);
nor U10123 (N_10123,N_7790,N_8121);
nor U10124 (N_10124,N_6943,N_8508);
or U10125 (N_10125,N_8481,N_7875);
nand U10126 (N_10126,N_8378,N_6960);
nand U10127 (N_10127,N_8964,N_7448);
nand U10128 (N_10128,N_8248,N_7318);
nor U10129 (N_10129,N_6715,N_7278);
nand U10130 (N_10130,N_7762,N_6445);
nand U10131 (N_10131,N_6597,N_7755);
and U10132 (N_10132,N_6399,N_7136);
nand U10133 (N_10133,N_8422,N_8533);
nand U10134 (N_10134,N_7313,N_6253);
or U10135 (N_10135,N_7516,N_8109);
and U10136 (N_10136,N_8342,N_7127);
nor U10137 (N_10137,N_6862,N_7756);
and U10138 (N_10138,N_7028,N_8710);
and U10139 (N_10139,N_8950,N_6054);
nand U10140 (N_10140,N_8944,N_7411);
and U10141 (N_10141,N_7135,N_7634);
nand U10142 (N_10142,N_7524,N_8931);
nand U10143 (N_10143,N_6322,N_6723);
nand U10144 (N_10144,N_8078,N_8411);
and U10145 (N_10145,N_7226,N_7306);
nor U10146 (N_10146,N_6133,N_8790);
or U10147 (N_10147,N_6034,N_7167);
and U10148 (N_10148,N_8810,N_7359);
and U10149 (N_10149,N_7609,N_8935);
nand U10150 (N_10150,N_8877,N_7630);
or U10151 (N_10151,N_7070,N_6126);
and U10152 (N_10152,N_7239,N_7427);
and U10153 (N_10153,N_6815,N_6596);
or U10154 (N_10154,N_6219,N_8956);
and U10155 (N_10155,N_6624,N_6841);
nor U10156 (N_10156,N_7339,N_6444);
nand U10157 (N_10157,N_6117,N_7177);
or U10158 (N_10158,N_6184,N_6252);
nor U10159 (N_10159,N_6341,N_8354);
or U10160 (N_10160,N_8408,N_8650);
or U10161 (N_10161,N_7730,N_6377);
nand U10162 (N_10162,N_8450,N_7441);
nor U10163 (N_10163,N_7369,N_6804);
and U10164 (N_10164,N_8037,N_7739);
nand U10165 (N_10165,N_7197,N_6223);
and U10166 (N_10166,N_6066,N_7961);
nor U10167 (N_10167,N_8524,N_8609);
or U10168 (N_10168,N_7271,N_7670);
nand U10169 (N_10169,N_6298,N_7817);
nand U10170 (N_10170,N_6656,N_7277);
or U10171 (N_10171,N_7346,N_8439);
nor U10172 (N_10172,N_7322,N_6434);
xnor U10173 (N_10173,N_7332,N_8496);
nand U10174 (N_10174,N_8734,N_6276);
nor U10175 (N_10175,N_7251,N_7072);
nor U10176 (N_10176,N_7770,N_8739);
nor U10177 (N_10177,N_6405,N_8051);
or U10178 (N_10178,N_6736,N_6664);
nor U10179 (N_10179,N_6956,N_8927);
and U10180 (N_10180,N_7032,N_8903);
nand U10181 (N_10181,N_8289,N_7667);
or U10182 (N_10182,N_8075,N_7878);
and U10183 (N_10183,N_7710,N_6263);
nor U10184 (N_10184,N_8227,N_8562);
and U10185 (N_10185,N_7873,N_6959);
and U10186 (N_10186,N_7293,N_8811);
and U10187 (N_10187,N_8273,N_7082);
and U10188 (N_10188,N_6368,N_7862);
and U10189 (N_10189,N_8324,N_6726);
and U10190 (N_10190,N_6630,N_7808);
nand U10191 (N_10191,N_8677,N_8237);
or U10192 (N_10192,N_7715,N_6604);
nand U10193 (N_10193,N_6355,N_6348);
and U10194 (N_10194,N_7891,N_8208);
nand U10195 (N_10195,N_7439,N_6779);
and U10196 (N_10196,N_7075,N_6662);
nand U10197 (N_10197,N_7113,N_7495);
nand U10198 (N_10198,N_8881,N_7194);
and U10199 (N_10199,N_7799,N_7168);
or U10200 (N_10200,N_6899,N_6009);
or U10201 (N_10201,N_8087,N_6404);
nand U10202 (N_10202,N_6215,N_6016);
and U10203 (N_10203,N_7975,N_7370);
nor U10204 (N_10204,N_6483,N_7466);
and U10205 (N_10205,N_6418,N_7852);
or U10206 (N_10206,N_7193,N_7632);
nand U10207 (N_10207,N_8590,N_8032);
nor U10208 (N_10208,N_7144,N_7978);
or U10209 (N_10209,N_6797,N_6288);
nor U10210 (N_10210,N_8234,N_7763);
and U10211 (N_10211,N_6340,N_7950);
or U10212 (N_10212,N_8745,N_8800);
nor U10213 (N_10213,N_8588,N_7304);
nand U10214 (N_10214,N_8990,N_7804);
and U10215 (N_10215,N_6529,N_7152);
nand U10216 (N_10216,N_8494,N_6469);
nor U10217 (N_10217,N_8272,N_6374);
or U10218 (N_10218,N_8803,N_8281);
or U10219 (N_10219,N_6923,N_6546);
xnor U10220 (N_10220,N_6908,N_8187);
nand U10221 (N_10221,N_8219,N_8017);
and U10222 (N_10222,N_7003,N_8061);
nor U10223 (N_10223,N_8681,N_8258);
nand U10224 (N_10224,N_7560,N_6390);
and U10225 (N_10225,N_6259,N_7921);
or U10226 (N_10226,N_7923,N_6180);
nand U10227 (N_10227,N_7791,N_6755);
or U10228 (N_10228,N_7410,N_7826);
nand U10229 (N_10229,N_8498,N_6461);
nand U10230 (N_10230,N_7142,N_6614);
nor U10231 (N_10231,N_8892,N_6994);
xor U10232 (N_10232,N_7543,N_8171);
and U10233 (N_10233,N_6218,N_8893);
and U10234 (N_10234,N_7953,N_6632);
nand U10235 (N_10235,N_6823,N_8668);
and U10236 (N_10236,N_6877,N_7811);
nand U10237 (N_10237,N_7310,N_8792);
and U10238 (N_10238,N_8648,N_8164);
xnor U10239 (N_10239,N_7453,N_8780);
and U10240 (N_10240,N_8253,N_7701);
and U10241 (N_10241,N_7918,N_6533);
nand U10242 (N_10242,N_8581,N_7108);
or U10243 (N_10243,N_6080,N_6836);
and U10244 (N_10244,N_6349,N_8938);
and U10245 (N_10245,N_6345,N_6014);
xor U10246 (N_10246,N_8251,N_6116);
or U10247 (N_10247,N_7566,N_6079);
and U10248 (N_10248,N_8693,N_8667);
nand U10249 (N_10249,N_7922,N_8250);
or U10250 (N_10250,N_7598,N_8117);
nor U10251 (N_10251,N_8501,N_7705);
nor U10252 (N_10252,N_6441,N_6554);
nand U10253 (N_10253,N_8297,N_8597);
nor U10254 (N_10254,N_6713,N_8723);
nand U10255 (N_10255,N_8458,N_7234);
nor U10256 (N_10256,N_7842,N_7296);
or U10257 (N_10257,N_6100,N_8776);
or U10258 (N_10258,N_8512,N_8265);
or U10259 (N_10259,N_6227,N_8860);
and U10260 (N_10260,N_6318,N_7333);
and U10261 (N_10261,N_6414,N_8626);
nor U10262 (N_10262,N_8715,N_8929);
nand U10263 (N_10263,N_8829,N_8260);
and U10264 (N_10264,N_7111,N_7668);
or U10265 (N_10265,N_6866,N_7703);
nand U10266 (N_10266,N_8536,N_6821);
or U10267 (N_10267,N_6798,N_8030);
nor U10268 (N_10268,N_7126,N_6167);
nor U10269 (N_10269,N_6612,N_6006);
or U10270 (N_10270,N_7289,N_6867);
nor U10271 (N_10271,N_8317,N_6968);
nor U10272 (N_10272,N_7795,N_6583);
or U10273 (N_10273,N_8694,N_8584);
nand U10274 (N_10274,N_7468,N_6030);
or U10275 (N_10275,N_6853,N_6706);
nor U10276 (N_10276,N_7624,N_6507);
and U10277 (N_10277,N_7688,N_7452);
nor U10278 (N_10278,N_7821,N_6670);
nor U10279 (N_10279,N_6051,N_7382);
or U10280 (N_10280,N_8814,N_7995);
or U10281 (N_10281,N_8049,N_7648);
and U10282 (N_10282,N_8819,N_8166);
nand U10283 (N_10283,N_7750,N_8274);
nand U10284 (N_10284,N_6094,N_7652);
or U10285 (N_10285,N_6613,N_7390);
nand U10286 (N_10286,N_7835,N_8779);
or U10287 (N_10287,N_6336,N_8836);
xnor U10288 (N_10288,N_6607,N_8119);
nor U10289 (N_10289,N_8867,N_6027);
nor U10290 (N_10290,N_7959,N_8111);
or U10291 (N_10291,N_7783,N_6379);
nand U10292 (N_10292,N_6575,N_6359);
or U10293 (N_10293,N_8491,N_6426);
nand U10294 (N_10294,N_8178,N_7732);
and U10295 (N_10295,N_8602,N_7347);
nand U10296 (N_10296,N_7288,N_7414);
or U10297 (N_10297,N_8161,N_8463);
nand U10298 (N_10298,N_6342,N_6196);
nor U10299 (N_10299,N_8428,N_6940);
nand U10300 (N_10300,N_6638,N_7933);
nor U10301 (N_10301,N_6658,N_6902);
nor U10302 (N_10302,N_6760,N_6572);
and U10303 (N_10303,N_7272,N_6150);
nor U10304 (N_10304,N_8914,N_8421);
or U10305 (N_10305,N_7129,N_7350);
nor U10306 (N_10306,N_7054,N_8210);
or U10307 (N_10307,N_7837,N_8082);
and U10308 (N_10308,N_7610,N_8922);
nand U10309 (N_10309,N_6503,N_8459);
nand U10310 (N_10310,N_6408,N_6320);
nand U10311 (N_10311,N_7371,N_6393);
nor U10312 (N_10312,N_6472,N_6287);
nor U10313 (N_10313,N_7387,N_7936);
or U10314 (N_10314,N_8510,N_7622);
or U10315 (N_10315,N_8013,N_6266);
nor U10316 (N_10316,N_7749,N_7256);
nand U10317 (N_10317,N_7935,N_8754);
nand U10318 (N_10318,N_6103,N_8673);
nand U10319 (N_10319,N_7079,N_7349);
nand U10320 (N_10320,N_7746,N_7863);
nor U10321 (N_10321,N_6163,N_7140);
nor U10322 (N_10322,N_7919,N_7949);
and U10323 (N_10323,N_6576,N_6357);
nand U10324 (N_10324,N_8714,N_7133);
and U10325 (N_10325,N_8521,N_6333);
or U10326 (N_10326,N_7775,N_8280);
xor U10327 (N_10327,N_7565,N_8201);
or U10328 (N_10328,N_7741,N_6743);
or U10329 (N_10329,N_7611,N_8915);
nand U10330 (N_10330,N_6973,N_6586);
nor U10331 (N_10331,N_7315,N_6183);
nor U10332 (N_10332,N_6925,N_8162);
and U10333 (N_10333,N_8399,N_6574);
and U10334 (N_10334,N_6602,N_8953);
nor U10335 (N_10335,N_6141,N_8837);
and U10336 (N_10336,N_8972,N_7942);
and U10337 (N_10337,N_8405,N_8152);
nor U10338 (N_10338,N_6431,N_7929);
nor U10339 (N_10339,N_6619,N_7957);
nor U10340 (N_10340,N_7532,N_8387);
nand U10341 (N_10341,N_8884,N_8592);
or U10342 (N_10342,N_6323,N_6216);
or U10343 (N_10343,N_6468,N_7143);
nor U10344 (N_10344,N_8732,N_8326);
nor U10345 (N_10345,N_6275,N_6235);
or U10346 (N_10346,N_7767,N_6448);
nand U10347 (N_10347,N_8566,N_7432);
nand U10348 (N_10348,N_7327,N_6934);
and U10349 (N_10349,N_7499,N_7068);
and U10350 (N_10350,N_8643,N_6671);
or U10351 (N_10351,N_6893,N_7782);
or U10352 (N_10352,N_8132,N_8335);
xor U10353 (N_10353,N_7833,N_6207);
nor U10354 (N_10354,N_8689,N_8760);
or U10355 (N_10355,N_7578,N_6175);
and U10356 (N_10356,N_8954,N_8659);
and U10357 (N_10357,N_7586,N_8674);
and U10358 (N_10358,N_8060,N_8737);
or U10359 (N_10359,N_8926,N_7849);
nand U10360 (N_10360,N_8386,N_7049);
nor U10361 (N_10361,N_7623,N_6594);
or U10362 (N_10362,N_7930,N_6082);
nand U10363 (N_10363,N_8442,N_6580);
and U10364 (N_10364,N_7944,N_7451);
and U10365 (N_10365,N_6251,N_8705);
nor U10366 (N_10366,N_8220,N_6008);
or U10367 (N_10367,N_8206,N_6018);
nor U10368 (N_10368,N_7617,N_8888);
and U10369 (N_10369,N_8851,N_7081);
or U10370 (N_10370,N_6021,N_7391);
and U10371 (N_10371,N_8460,N_7845);
nand U10372 (N_10372,N_7021,N_6154);
nor U10373 (N_10373,N_6306,N_6197);
nand U10374 (N_10374,N_6683,N_6714);
or U10375 (N_10375,N_6350,N_6903);
or U10376 (N_10376,N_7917,N_6384);
nand U10377 (N_10377,N_7615,N_8960);
nor U10378 (N_10378,N_8831,N_6558);
nand U10379 (N_10379,N_6890,N_8269);
or U10380 (N_10380,N_7465,N_8961);
nand U10381 (N_10381,N_7991,N_6562);
nor U10382 (N_10382,N_8548,N_8911);
and U10383 (N_10383,N_7547,N_8343);
nand U10384 (N_10384,N_8726,N_6951);
nor U10385 (N_10385,N_8731,N_7952);
nor U10386 (N_10386,N_8063,N_7779);
and U10387 (N_10387,N_6947,N_6327);
or U10388 (N_10388,N_7677,N_8007);
nor U10389 (N_10389,N_8318,N_8040);
nand U10390 (N_10390,N_7494,N_7445);
and U10391 (N_10391,N_7656,N_7104);
nand U10392 (N_10392,N_7184,N_7706);
or U10393 (N_10393,N_7149,N_7941);
or U10394 (N_10394,N_7698,N_7527);
nand U10395 (N_10395,N_8589,N_8551);
nor U10396 (N_10396,N_6848,N_6905);
nor U10397 (N_10397,N_6250,N_7151);
nor U10398 (N_10398,N_6181,N_8976);
and U10399 (N_10399,N_6536,N_7647);
nand U10400 (N_10400,N_6280,N_6649);
nand U10401 (N_10401,N_7190,N_8254);
nand U10402 (N_10402,N_7199,N_8455);
and U10403 (N_10403,N_6703,N_8625);
nand U10404 (N_10404,N_8372,N_6830);
nand U10405 (N_10405,N_6354,N_8959);
or U10406 (N_10406,N_8763,N_6273);
nand U10407 (N_10407,N_6031,N_6090);
nand U10408 (N_10408,N_7164,N_6857);
or U10409 (N_10409,N_8151,N_8894);
and U10410 (N_10410,N_7062,N_8205);
and U10411 (N_10411,N_6491,N_6410);
or U10412 (N_10412,N_7355,N_8921);
or U10413 (N_10413,N_6976,N_8050);
or U10414 (N_10414,N_8240,N_6352);
and U10415 (N_10415,N_7549,N_6411);
nand U10416 (N_10416,N_6224,N_7765);
and U10417 (N_10417,N_8777,N_8153);
and U10418 (N_10418,N_8284,N_8034);
nand U10419 (N_10419,N_7679,N_7828);
nand U10420 (N_10420,N_8716,N_8657);
nand U10421 (N_10421,N_8728,N_6611);
nand U10422 (N_10422,N_8573,N_8604);
or U10423 (N_10423,N_8849,N_7308);
nand U10424 (N_10424,N_8865,N_6983);
and U10425 (N_10425,N_7971,N_7446);
and U10426 (N_10426,N_8074,N_8262);
and U10427 (N_10427,N_7185,N_6946);
or U10428 (N_10428,N_8765,N_8635);
nor U10429 (N_10429,N_7392,N_7697);
or U10430 (N_10430,N_7576,N_7034);
nand U10431 (N_10431,N_8910,N_7431);
or U10432 (N_10432,N_7409,N_6808);
nand U10433 (N_10433,N_8846,N_8781);
or U10434 (N_10434,N_7259,N_7601);
nor U10435 (N_10435,N_8820,N_8869);
or U10436 (N_10436,N_8973,N_8624);
nor U10437 (N_10437,N_7612,N_7123);
or U10438 (N_10438,N_7858,N_8813);
nand U10439 (N_10439,N_8622,N_6376);
and U10440 (N_10440,N_8267,N_8470);
or U10441 (N_10441,N_8179,N_8000);
or U10442 (N_10442,N_8506,N_7522);
nor U10443 (N_10443,N_8572,N_8375);
nand U10444 (N_10444,N_7726,N_8560);
and U10445 (N_10445,N_8484,N_6493);
or U10446 (N_10446,N_8315,N_7002);
nor U10447 (N_10447,N_7491,N_8633);
nand U10448 (N_10448,N_8480,N_6424);
nand U10449 (N_10449,N_8546,N_6832);
and U10450 (N_10450,N_8176,N_6997);
or U10451 (N_10451,N_7777,N_7263);
nor U10452 (N_10452,N_6353,N_7007);
or U10453 (N_10453,N_6824,N_6199);
and U10454 (N_10454,N_6698,N_6413);
nand U10455 (N_10455,N_6381,N_6606);
or U10456 (N_10456,N_7437,N_8385);
and U10457 (N_10457,N_6991,N_7307);
and U10458 (N_10458,N_8784,N_8073);
nand U10459 (N_10459,N_8970,N_6980);
or U10460 (N_10460,N_6907,N_6182);
and U10461 (N_10461,N_8736,N_7805);
and U10462 (N_10462,N_6806,N_7888);
and U10463 (N_10463,N_7025,N_6467);
and U10464 (N_10464,N_8156,N_6837);
or U10465 (N_10465,N_6999,N_8928);
nand U10466 (N_10466,N_8751,N_8895);
and U10467 (N_10467,N_8788,N_7968);
and U10468 (N_10468,N_7044,N_7273);
nand U10469 (N_10469,N_7305,N_8035);
or U10470 (N_10470,N_7280,N_8158);
or U10471 (N_10471,N_8509,N_7163);
nand U10472 (N_10472,N_6011,N_7702);
or U10473 (N_10473,N_7473,N_7672);
nor U10474 (N_10474,N_6775,N_7459);
xor U10475 (N_10475,N_6781,N_6373);
and U10476 (N_10476,N_8453,N_8348);
and U10477 (N_10477,N_7106,N_7682);
nand U10478 (N_10478,N_8838,N_6236);
nor U10479 (N_10479,N_6186,N_7771);
or U10480 (N_10480,N_6941,N_8832);
and U10481 (N_10481,N_6928,N_7039);
nor U10482 (N_10482,N_8296,N_6565);
and U10483 (N_10483,N_7860,N_8389);
or U10484 (N_10484,N_6579,N_6647);
or U10485 (N_10485,N_6741,N_8640);
nor U10486 (N_10486,N_7743,N_8616);
nand U10487 (N_10487,N_8323,N_7595);
or U10488 (N_10488,N_8123,N_6534);
nor U10489 (N_10489,N_6149,N_8804);
and U10490 (N_10490,N_7121,N_6567);
or U10491 (N_10491,N_6738,N_7737);
and U10492 (N_10492,N_6864,N_8301);
or U10493 (N_10493,N_8568,N_6470);
xnor U10494 (N_10494,N_7302,N_6220);
or U10495 (N_10495,N_6707,N_8607);
or U10496 (N_10496,N_7213,N_7999);
or U10497 (N_10497,N_8890,N_6058);
or U10498 (N_10498,N_7101,N_6693);
nor U10499 (N_10499,N_7618,N_8527);
and U10500 (N_10500,N_8009,N_8107);
and U10501 (N_10501,N_6142,N_7960);
nand U10502 (N_10502,N_7911,N_8319);
nand U10503 (N_10503,N_7138,N_7184);
and U10504 (N_10504,N_6923,N_8046);
or U10505 (N_10505,N_8785,N_6655);
nor U10506 (N_10506,N_7810,N_8874);
and U10507 (N_10507,N_7045,N_8994);
nand U10508 (N_10508,N_7872,N_8609);
and U10509 (N_10509,N_7588,N_6246);
or U10510 (N_10510,N_6874,N_7168);
or U10511 (N_10511,N_7767,N_8427);
nand U10512 (N_10512,N_7198,N_8549);
nand U10513 (N_10513,N_8553,N_8042);
and U10514 (N_10514,N_8368,N_7136);
or U10515 (N_10515,N_8208,N_6742);
and U10516 (N_10516,N_7435,N_8714);
or U10517 (N_10517,N_8863,N_8293);
or U10518 (N_10518,N_8276,N_7751);
and U10519 (N_10519,N_8235,N_8782);
nor U10520 (N_10520,N_6084,N_6424);
or U10521 (N_10521,N_8528,N_8441);
and U10522 (N_10522,N_6487,N_6704);
or U10523 (N_10523,N_6485,N_7066);
nor U10524 (N_10524,N_8777,N_8060);
nand U10525 (N_10525,N_6500,N_8614);
or U10526 (N_10526,N_8399,N_7777);
and U10527 (N_10527,N_8391,N_7299);
nor U10528 (N_10528,N_6230,N_7088);
nand U10529 (N_10529,N_8415,N_7006);
nand U10530 (N_10530,N_6438,N_6937);
nor U10531 (N_10531,N_8403,N_6285);
and U10532 (N_10532,N_6293,N_7611);
nand U10533 (N_10533,N_8423,N_8589);
nor U10534 (N_10534,N_8103,N_6944);
nor U10535 (N_10535,N_8975,N_7182);
nand U10536 (N_10536,N_6748,N_8406);
xnor U10537 (N_10537,N_8881,N_7644);
nor U10538 (N_10538,N_6176,N_8042);
and U10539 (N_10539,N_7900,N_8199);
nand U10540 (N_10540,N_7801,N_6232);
nor U10541 (N_10541,N_8975,N_6489);
nor U10542 (N_10542,N_6577,N_7325);
nor U10543 (N_10543,N_6098,N_7064);
and U10544 (N_10544,N_7999,N_6174);
and U10545 (N_10545,N_8539,N_6313);
and U10546 (N_10546,N_7198,N_8645);
nor U10547 (N_10547,N_8434,N_6821);
nand U10548 (N_10548,N_6291,N_7057);
or U10549 (N_10549,N_7178,N_6731);
and U10550 (N_10550,N_6906,N_8273);
nor U10551 (N_10551,N_7574,N_6828);
and U10552 (N_10552,N_7841,N_6932);
nand U10553 (N_10553,N_7639,N_7760);
or U10554 (N_10554,N_7106,N_7351);
nor U10555 (N_10555,N_8526,N_6425);
or U10556 (N_10556,N_6104,N_7013);
or U10557 (N_10557,N_6969,N_7059);
or U10558 (N_10558,N_8112,N_7876);
and U10559 (N_10559,N_8324,N_8266);
nand U10560 (N_10560,N_6646,N_8363);
and U10561 (N_10561,N_6995,N_8017);
nand U10562 (N_10562,N_6809,N_6772);
or U10563 (N_10563,N_8586,N_8968);
nand U10564 (N_10564,N_6000,N_7092);
or U10565 (N_10565,N_8099,N_6016);
nand U10566 (N_10566,N_6566,N_6316);
or U10567 (N_10567,N_6687,N_7285);
and U10568 (N_10568,N_7750,N_8245);
and U10569 (N_10569,N_6923,N_8969);
and U10570 (N_10570,N_7424,N_7256);
nor U10571 (N_10571,N_7226,N_6448);
and U10572 (N_10572,N_6207,N_8747);
or U10573 (N_10573,N_7245,N_8752);
or U10574 (N_10574,N_8947,N_8187);
and U10575 (N_10575,N_6823,N_8143);
and U10576 (N_10576,N_7236,N_7957);
nor U10577 (N_10577,N_6415,N_7447);
or U10578 (N_10578,N_6553,N_8990);
or U10579 (N_10579,N_8539,N_8627);
nand U10580 (N_10580,N_8213,N_6341);
or U10581 (N_10581,N_7068,N_7161);
and U10582 (N_10582,N_7597,N_8394);
nor U10583 (N_10583,N_8573,N_7896);
and U10584 (N_10584,N_6297,N_6247);
nand U10585 (N_10585,N_7989,N_6633);
nor U10586 (N_10586,N_7280,N_7311);
and U10587 (N_10587,N_6839,N_8688);
nor U10588 (N_10588,N_8270,N_7618);
and U10589 (N_10589,N_8444,N_7357);
and U10590 (N_10590,N_7498,N_6915);
or U10591 (N_10591,N_7333,N_7750);
and U10592 (N_10592,N_8827,N_6939);
nor U10593 (N_10593,N_7751,N_7957);
or U10594 (N_10594,N_6013,N_8896);
nor U10595 (N_10595,N_6895,N_6429);
nor U10596 (N_10596,N_6213,N_6375);
nand U10597 (N_10597,N_7809,N_6931);
nor U10598 (N_10598,N_8364,N_8912);
nand U10599 (N_10599,N_7057,N_7683);
nand U10600 (N_10600,N_7031,N_8109);
and U10601 (N_10601,N_7028,N_8451);
nand U10602 (N_10602,N_8334,N_7236);
nand U10603 (N_10603,N_8468,N_7237);
and U10604 (N_10604,N_8912,N_7884);
xnor U10605 (N_10605,N_8279,N_6286);
nor U10606 (N_10606,N_7075,N_8538);
and U10607 (N_10607,N_8152,N_6329);
nor U10608 (N_10608,N_7053,N_6823);
or U10609 (N_10609,N_8771,N_6071);
or U10610 (N_10610,N_7946,N_8504);
or U10611 (N_10611,N_7554,N_8112);
and U10612 (N_10612,N_8021,N_6137);
nand U10613 (N_10613,N_8206,N_6604);
nor U10614 (N_10614,N_6656,N_6804);
or U10615 (N_10615,N_6747,N_7355);
nand U10616 (N_10616,N_7555,N_8122);
nor U10617 (N_10617,N_8155,N_8877);
nor U10618 (N_10618,N_6063,N_7536);
nand U10619 (N_10619,N_7917,N_8432);
and U10620 (N_10620,N_7104,N_8373);
nand U10621 (N_10621,N_8973,N_6671);
nor U10622 (N_10622,N_6186,N_7243);
and U10623 (N_10623,N_7579,N_8758);
or U10624 (N_10624,N_7034,N_7944);
nor U10625 (N_10625,N_8911,N_8967);
and U10626 (N_10626,N_8533,N_7916);
nor U10627 (N_10627,N_6636,N_6919);
or U10628 (N_10628,N_6643,N_8189);
nand U10629 (N_10629,N_7978,N_6843);
and U10630 (N_10630,N_6693,N_6210);
and U10631 (N_10631,N_7112,N_7785);
nand U10632 (N_10632,N_8959,N_8244);
nor U10633 (N_10633,N_7111,N_6831);
and U10634 (N_10634,N_8577,N_6921);
or U10635 (N_10635,N_8950,N_7259);
and U10636 (N_10636,N_8355,N_8713);
nand U10637 (N_10637,N_7246,N_8396);
nor U10638 (N_10638,N_7894,N_6449);
and U10639 (N_10639,N_7916,N_6733);
nor U10640 (N_10640,N_8725,N_8802);
xor U10641 (N_10641,N_6996,N_7478);
and U10642 (N_10642,N_8042,N_7014);
nor U10643 (N_10643,N_8410,N_7551);
or U10644 (N_10644,N_8938,N_8351);
nand U10645 (N_10645,N_6470,N_8320);
nand U10646 (N_10646,N_7966,N_6985);
nor U10647 (N_10647,N_8532,N_6743);
or U10648 (N_10648,N_7705,N_8753);
or U10649 (N_10649,N_7655,N_6930);
and U10650 (N_10650,N_6272,N_8117);
nand U10651 (N_10651,N_7052,N_8428);
nand U10652 (N_10652,N_8276,N_7868);
nand U10653 (N_10653,N_6851,N_6383);
and U10654 (N_10654,N_7551,N_6474);
or U10655 (N_10655,N_8448,N_7278);
nand U10656 (N_10656,N_6437,N_6811);
nand U10657 (N_10657,N_7008,N_7566);
or U10658 (N_10658,N_7525,N_6671);
or U10659 (N_10659,N_6748,N_6578);
nand U10660 (N_10660,N_7059,N_8577);
and U10661 (N_10661,N_7030,N_6339);
nor U10662 (N_10662,N_7613,N_8414);
or U10663 (N_10663,N_7554,N_6741);
and U10664 (N_10664,N_6658,N_6484);
nor U10665 (N_10665,N_8549,N_7634);
and U10666 (N_10666,N_8071,N_7195);
or U10667 (N_10667,N_8232,N_7007);
nor U10668 (N_10668,N_6341,N_7105);
and U10669 (N_10669,N_8290,N_7367);
nor U10670 (N_10670,N_7337,N_7526);
nor U10671 (N_10671,N_6512,N_8862);
nand U10672 (N_10672,N_6542,N_7190);
or U10673 (N_10673,N_7349,N_8972);
and U10674 (N_10674,N_6792,N_8462);
nand U10675 (N_10675,N_8781,N_6914);
and U10676 (N_10676,N_7767,N_8144);
or U10677 (N_10677,N_8088,N_6504);
and U10678 (N_10678,N_6188,N_7759);
nand U10679 (N_10679,N_8242,N_8238);
and U10680 (N_10680,N_8155,N_6365);
nand U10681 (N_10681,N_8775,N_6748);
nand U10682 (N_10682,N_6909,N_6546);
and U10683 (N_10683,N_6304,N_6842);
and U10684 (N_10684,N_8558,N_6152);
and U10685 (N_10685,N_6077,N_6456);
or U10686 (N_10686,N_6231,N_6449);
nor U10687 (N_10687,N_8302,N_8090);
or U10688 (N_10688,N_6547,N_6755);
or U10689 (N_10689,N_8306,N_6456);
nand U10690 (N_10690,N_6716,N_8864);
and U10691 (N_10691,N_7160,N_8918);
and U10692 (N_10692,N_8050,N_8409);
and U10693 (N_10693,N_7861,N_7060);
nand U10694 (N_10694,N_8777,N_8469);
or U10695 (N_10695,N_7199,N_7859);
or U10696 (N_10696,N_6805,N_6963);
nor U10697 (N_10697,N_8694,N_6155);
or U10698 (N_10698,N_8785,N_6529);
or U10699 (N_10699,N_6880,N_8332);
nor U10700 (N_10700,N_8881,N_6917);
or U10701 (N_10701,N_8023,N_8448);
nand U10702 (N_10702,N_8155,N_8724);
nand U10703 (N_10703,N_6266,N_6958);
and U10704 (N_10704,N_6100,N_8442);
and U10705 (N_10705,N_8998,N_8793);
and U10706 (N_10706,N_7441,N_8041);
nand U10707 (N_10707,N_7023,N_7951);
nand U10708 (N_10708,N_7795,N_7471);
xnor U10709 (N_10709,N_7145,N_8043);
nand U10710 (N_10710,N_8210,N_6408);
and U10711 (N_10711,N_6112,N_6970);
nor U10712 (N_10712,N_8950,N_6648);
nand U10713 (N_10713,N_6982,N_7763);
and U10714 (N_10714,N_7669,N_7075);
and U10715 (N_10715,N_8215,N_6494);
nor U10716 (N_10716,N_7355,N_6289);
nand U10717 (N_10717,N_8710,N_7036);
nand U10718 (N_10718,N_8992,N_6079);
nand U10719 (N_10719,N_6498,N_6820);
nor U10720 (N_10720,N_6393,N_6610);
or U10721 (N_10721,N_8861,N_7492);
nand U10722 (N_10722,N_8355,N_7178);
nand U10723 (N_10723,N_8542,N_7923);
or U10724 (N_10724,N_6262,N_8628);
or U10725 (N_10725,N_6424,N_6899);
and U10726 (N_10726,N_7188,N_7927);
nand U10727 (N_10727,N_6828,N_7597);
nand U10728 (N_10728,N_8029,N_6720);
nor U10729 (N_10729,N_6805,N_7580);
and U10730 (N_10730,N_6290,N_7385);
nand U10731 (N_10731,N_7529,N_7605);
nor U10732 (N_10732,N_8970,N_7795);
and U10733 (N_10733,N_7870,N_7022);
or U10734 (N_10734,N_8728,N_7658);
nor U10735 (N_10735,N_8417,N_8574);
nand U10736 (N_10736,N_7795,N_7972);
nand U10737 (N_10737,N_8261,N_7426);
or U10738 (N_10738,N_8981,N_7312);
nand U10739 (N_10739,N_8338,N_8436);
or U10740 (N_10740,N_6380,N_6302);
and U10741 (N_10741,N_7971,N_7833);
or U10742 (N_10742,N_8295,N_6290);
nor U10743 (N_10743,N_8610,N_7418);
nand U10744 (N_10744,N_7774,N_7541);
and U10745 (N_10745,N_7746,N_8630);
nor U10746 (N_10746,N_6313,N_6701);
nand U10747 (N_10747,N_6597,N_7969);
nor U10748 (N_10748,N_7197,N_7967);
nand U10749 (N_10749,N_8917,N_6726);
nor U10750 (N_10750,N_8330,N_6684);
and U10751 (N_10751,N_7980,N_7509);
or U10752 (N_10752,N_7514,N_7866);
or U10753 (N_10753,N_6968,N_7488);
or U10754 (N_10754,N_7960,N_8081);
and U10755 (N_10755,N_7921,N_8255);
nor U10756 (N_10756,N_6731,N_6340);
and U10757 (N_10757,N_8182,N_8274);
or U10758 (N_10758,N_6683,N_8188);
nor U10759 (N_10759,N_6940,N_6047);
or U10760 (N_10760,N_6494,N_7770);
nand U10761 (N_10761,N_6063,N_7986);
nor U10762 (N_10762,N_8264,N_8919);
nand U10763 (N_10763,N_6979,N_8572);
nor U10764 (N_10764,N_6273,N_6831);
and U10765 (N_10765,N_6175,N_6858);
nand U10766 (N_10766,N_8155,N_8766);
or U10767 (N_10767,N_8321,N_7129);
nand U10768 (N_10768,N_8822,N_6828);
and U10769 (N_10769,N_7529,N_7553);
nor U10770 (N_10770,N_7382,N_6755);
nor U10771 (N_10771,N_6601,N_8721);
and U10772 (N_10772,N_7266,N_7760);
nor U10773 (N_10773,N_6072,N_7711);
nor U10774 (N_10774,N_8578,N_8523);
and U10775 (N_10775,N_7997,N_6456);
nor U10776 (N_10776,N_6296,N_7754);
nor U10777 (N_10777,N_8043,N_7558);
and U10778 (N_10778,N_7936,N_8867);
or U10779 (N_10779,N_8789,N_7320);
nand U10780 (N_10780,N_6534,N_7862);
nand U10781 (N_10781,N_8324,N_7663);
or U10782 (N_10782,N_6092,N_8085);
or U10783 (N_10783,N_6543,N_7237);
and U10784 (N_10784,N_6427,N_6366);
nor U10785 (N_10785,N_8732,N_8418);
or U10786 (N_10786,N_6488,N_8689);
nand U10787 (N_10787,N_6395,N_7354);
nor U10788 (N_10788,N_8679,N_7288);
nor U10789 (N_10789,N_7071,N_8612);
nand U10790 (N_10790,N_7742,N_7475);
or U10791 (N_10791,N_7911,N_7018);
nand U10792 (N_10792,N_8972,N_8050);
nand U10793 (N_10793,N_6729,N_6517);
xor U10794 (N_10794,N_8781,N_6741);
nand U10795 (N_10795,N_7050,N_7381);
nand U10796 (N_10796,N_7249,N_7267);
or U10797 (N_10797,N_8430,N_7836);
or U10798 (N_10798,N_7952,N_6158);
or U10799 (N_10799,N_7599,N_6464);
nand U10800 (N_10800,N_8812,N_6164);
nor U10801 (N_10801,N_7395,N_8626);
and U10802 (N_10802,N_7166,N_6557);
nor U10803 (N_10803,N_6198,N_6852);
and U10804 (N_10804,N_8881,N_7121);
nand U10805 (N_10805,N_6179,N_6861);
and U10806 (N_10806,N_8108,N_6053);
or U10807 (N_10807,N_6491,N_8228);
or U10808 (N_10808,N_7426,N_6943);
nor U10809 (N_10809,N_7613,N_6205);
nand U10810 (N_10810,N_7690,N_7402);
xor U10811 (N_10811,N_8079,N_7506);
or U10812 (N_10812,N_6145,N_7780);
nand U10813 (N_10813,N_8159,N_8611);
nand U10814 (N_10814,N_6134,N_7957);
nand U10815 (N_10815,N_7665,N_8099);
and U10816 (N_10816,N_6773,N_7767);
or U10817 (N_10817,N_7198,N_7358);
and U10818 (N_10818,N_7484,N_8950);
or U10819 (N_10819,N_7406,N_7381);
or U10820 (N_10820,N_8051,N_7963);
nor U10821 (N_10821,N_7805,N_7793);
and U10822 (N_10822,N_8935,N_7689);
nor U10823 (N_10823,N_6364,N_8155);
and U10824 (N_10824,N_7364,N_6983);
or U10825 (N_10825,N_7776,N_7522);
and U10826 (N_10826,N_6368,N_8387);
and U10827 (N_10827,N_7754,N_8140);
nor U10828 (N_10828,N_6722,N_7395);
nand U10829 (N_10829,N_7566,N_7823);
nand U10830 (N_10830,N_7888,N_8225);
or U10831 (N_10831,N_8897,N_8940);
nand U10832 (N_10832,N_8611,N_7956);
nand U10833 (N_10833,N_8736,N_7697);
or U10834 (N_10834,N_7913,N_8955);
nor U10835 (N_10835,N_7678,N_8484);
or U10836 (N_10836,N_6087,N_8017);
nand U10837 (N_10837,N_6631,N_8750);
nand U10838 (N_10838,N_7783,N_8271);
or U10839 (N_10839,N_7888,N_7165);
nor U10840 (N_10840,N_6874,N_8222);
or U10841 (N_10841,N_6221,N_7699);
nor U10842 (N_10842,N_6969,N_8351);
nand U10843 (N_10843,N_6489,N_6615);
or U10844 (N_10844,N_6999,N_7684);
nor U10845 (N_10845,N_7061,N_6338);
or U10846 (N_10846,N_8546,N_7484);
nor U10847 (N_10847,N_6341,N_8925);
nand U10848 (N_10848,N_6731,N_6508);
or U10849 (N_10849,N_6097,N_7718);
nand U10850 (N_10850,N_8111,N_7507);
or U10851 (N_10851,N_8311,N_6476);
and U10852 (N_10852,N_8740,N_7074);
nand U10853 (N_10853,N_8402,N_8427);
nand U10854 (N_10854,N_8256,N_7848);
nand U10855 (N_10855,N_7470,N_8743);
or U10856 (N_10856,N_8623,N_8730);
nor U10857 (N_10857,N_6250,N_8879);
nor U10858 (N_10858,N_7180,N_8012);
nand U10859 (N_10859,N_8236,N_6911);
nand U10860 (N_10860,N_7767,N_6192);
nand U10861 (N_10861,N_7577,N_7328);
or U10862 (N_10862,N_6744,N_8387);
nor U10863 (N_10863,N_6612,N_6646);
nand U10864 (N_10864,N_7295,N_8334);
or U10865 (N_10865,N_7034,N_7262);
or U10866 (N_10866,N_7926,N_6471);
and U10867 (N_10867,N_8175,N_7592);
nand U10868 (N_10868,N_8465,N_7819);
nor U10869 (N_10869,N_7601,N_6078);
and U10870 (N_10870,N_8366,N_7496);
nor U10871 (N_10871,N_6555,N_7518);
nor U10872 (N_10872,N_7008,N_7813);
and U10873 (N_10873,N_6421,N_6088);
and U10874 (N_10874,N_8957,N_6147);
nand U10875 (N_10875,N_7265,N_6188);
nand U10876 (N_10876,N_7125,N_6981);
nor U10877 (N_10877,N_8983,N_8272);
or U10878 (N_10878,N_7142,N_7621);
or U10879 (N_10879,N_7783,N_7869);
or U10880 (N_10880,N_8210,N_6659);
or U10881 (N_10881,N_6211,N_6432);
nand U10882 (N_10882,N_6022,N_8259);
or U10883 (N_10883,N_7717,N_6746);
or U10884 (N_10884,N_7769,N_8916);
or U10885 (N_10885,N_8945,N_8488);
nand U10886 (N_10886,N_8240,N_7470);
and U10887 (N_10887,N_6831,N_7941);
or U10888 (N_10888,N_6019,N_8074);
nor U10889 (N_10889,N_8503,N_7320);
and U10890 (N_10890,N_7225,N_6237);
and U10891 (N_10891,N_7625,N_8809);
nor U10892 (N_10892,N_6925,N_7426);
and U10893 (N_10893,N_7472,N_7707);
nand U10894 (N_10894,N_6306,N_7428);
or U10895 (N_10895,N_8686,N_8438);
nor U10896 (N_10896,N_7285,N_8850);
xor U10897 (N_10897,N_7710,N_8304);
nor U10898 (N_10898,N_8757,N_8330);
nand U10899 (N_10899,N_8959,N_6675);
or U10900 (N_10900,N_7134,N_7428);
nand U10901 (N_10901,N_6102,N_7242);
or U10902 (N_10902,N_6263,N_8726);
nand U10903 (N_10903,N_7696,N_8258);
and U10904 (N_10904,N_8380,N_8500);
or U10905 (N_10905,N_7017,N_8131);
nand U10906 (N_10906,N_8337,N_8785);
or U10907 (N_10907,N_8149,N_6809);
nand U10908 (N_10908,N_6751,N_7016);
or U10909 (N_10909,N_8925,N_7475);
or U10910 (N_10910,N_7570,N_6197);
and U10911 (N_10911,N_8640,N_6342);
nor U10912 (N_10912,N_8570,N_7759);
or U10913 (N_10913,N_8955,N_7282);
and U10914 (N_10914,N_8563,N_6852);
nand U10915 (N_10915,N_6832,N_8566);
nand U10916 (N_10916,N_6703,N_8965);
or U10917 (N_10917,N_7370,N_6704);
and U10918 (N_10918,N_6819,N_7863);
or U10919 (N_10919,N_8738,N_8482);
nor U10920 (N_10920,N_7845,N_8235);
xor U10921 (N_10921,N_7960,N_7086);
and U10922 (N_10922,N_7087,N_6044);
nor U10923 (N_10923,N_8258,N_8767);
nand U10924 (N_10924,N_7476,N_6868);
or U10925 (N_10925,N_8862,N_8385);
nand U10926 (N_10926,N_8850,N_8673);
nor U10927 (N_10927,N_6203,N_7022);
and U10928 (N_10928,N_7162,N_7540);
nand U10929 (N_10929,N_8101,N_8316);
nand U10930 (N_10930,N_7381,N_7481);
nor U10931 (N_10931,N_7147,N_8960);
nor U10932 (N_10932,N_7073,N_7525);
nor U10933 (N_10933,N_7211,N_7164);
or U10934 (N_10934,N_6794,N_7740);
nor U10935 (N_10935,N_8504,N_8489);
and U10936 (N_10936,N_6500,N_6522);
nand U10937 (N_10937,N_8860,N_8763);
and U10938 (N_10938,N_6045,N_8836);
and U10939 (N_10939,N_7731,N_7747);
nor U10940 (N_10940,N_8987,N_7498);
nand U10941 (N_10941,N_6524,N_6312);
or U10942 (N_10942,N_8973,N_6776);
or U10943 (N_10943,N_8659,N_8334);
and U10944 (N_10944,N_7619,N_6135);
and U10945 (N_10945,N_7005,N_8846);
nand U10946 (N_10946,N_8011,N_7419);
nor U10947 (N_10947,N_7652,N_7300);
nand U10948 (N_10948,N_8638,N_6651);
nor U10949 (N_10949,N_7492,N_8235);
nand U10950 (N_10950,N_7889,N_7091);
nand U10951 (N_10951,N_8718,N_8307);
or U10952 (N_10952,N_7993,N_6298);
nor U10953 (N_10953,N_8106,N_7415);
nand U10954 (N_10954,N_8778,N_7108);
nor U10955 (N_10955,N_8561,N_8429);
and U10956 (N_10956,N_7883,N_6367);
or U10957 (N_10957,N_8761,N_8539);
or U10958 (N_10958,N_7141,N_7814);
nand U10959 (N_10959,N_6952,N_8245);
or U10960 (N_10960,N_7842,N_7565);
or U10961 (N_10961,N_8349,N_7738);
or U10962 (N_10962,N_6880,N_8794);
or U10963 (N_10963,N_8814,N_8508);
nor U10964 (N_10964,N_6067,N_7174);
nand U10965 (N_10965,N_6933,N_7153);
or U10966 (N_10966,N_8018,N_6697);
or U10967 (N_10967,N_7532,N_6790);
nand U10968 (N_10968,N_8195,N_7452);
nand U10969 (N_10969,N_6286,N_8221);
or U10970 (N_10970,N_7466,N_7745);
nor U10971 (N_10971,N_6686,N_6495);
and U10972 (N_10972,N_6212,N_8397);
or U10973 (N_10973,N_7027,N_8242);
nor U10974 (N_10974,N_7990,N_6325);
and U10975 (N_10975,N_7195,N_6884);
nor U10976 (N_10976,N_7381,N_7205);
nor U10977 (N_10977,N_8686,N_6742);
or U10978 (N_10978,N_6979,N_6870);
and U10979 (N_10979,N_6911,N_7202);
nor U10980 (N_10980,N_6589,N_7383);
nor U10981 (N_10981,N_7869,N_7030);
or U10982 (N_10982,N_8231,N_8235);
nor U10983 (N_10983,N_8569,N_7537);
nor U10984 (N_10984,N_7039,N_7282);
and U10985 (N_10985,N_7795,N_7946);
and U10986 (N_10986,N_6384,N_6765);
nor U10987 (N_10987,N_8098,N_6983);
or U10988 (N_10988,N_8001,N_6682);
nand U10989 (N_10989,N_8958,N_6714);
nor U10990 (N_10990,N_8613,N_8231);
or U10991 (N_10991,N_6931,N_6272);
nand U10992 (N_10992,N_7325,N_7612);
nand U10993 (N_10993,N_7592,N_6665);
nor U10994 (N_10994,N_8753,N_8292);
nand U10995 (N_10995,N_8647,N_7019);
and U10996 (N_10996,N_8051,N_7631);
nor U10997 (N_10997,N_7380,N_8109);
or U10998 (N_10998,N_6250,N_6003);
nand U10999 (N_10999,N_7049,N_7835);
nor U11000 (N_11000,N_6206,N_7767);
nand U11001 (N_11001,N_8292,N_7357);
or U11002 (N_11002,N_7466,N_6298);
and U11003 (N_11003,N_6687,N_7804);
nor U11004 (N_11004,N_6246,N_8204);
nor U11005 (N_11005,N_8134,N_6821);
nand U11006 (N_11006,N_6585,N_7188);
nor U11007 (N_11007,N_6606,N_8444);
nand U11008 (N_11008,N_8364,N_8884);
and U11009 (N_11009,N_6274,N_6726);
nand U11010 (N_11010,N_6832,N_8918);
nor U11011 (N_11011,N_7920,N_7963);
nand U11012 (N_11012,N_6176,N_7296);
nor U11013 (N_11013,N_8699,N_8998);
nand U11014 (N_11014,N_6801,N_6856);
and U11015 (N_11015,N_8411,N_6797);
or U11016 (N_11016,N_8978,N_8569);
nor U11017 (N_11017,N_6058,N_6582);
and U11018 (N_11018,N_6547,N_7969);
and U11019 (N_11019,N_8773,N_8949);
or U11020 (N_11020,N_7103,N_8743);
nor U11021 (N_11021,N_8500,N_7927);
or U11022 (N_11022,N_8019,N_8650);
nor U11023 (N_11023,N_7110,N_7119);
and U11024 (N_11024,N_8182,N_6301);
or U11025 (N_11025,N_6901,N_6990);
nand U11026 (N_11026,N_8099,N_7164);
or U11027 (N_11027,N_7540,N_8098);
and U11028 (N_11028,N_8444,N_6695);
nand U11029 (N_11029,N_8181,N_6780);
nand U11030 (N_11030,N_8906,N_8813);
nor U11031 (N_11031,N_8199,N_8576);
nand U11032 (N_11032,N_8873,N_7850);
nand U11033 (N_11033,N_8801,N_6802);
nand U11034 (N_11034,N_8699,N_8312);
and U11035 (N_11035,N_8021,N_7421);
nor U11036 (N_11036,N_7430,N_7488);
or U11037 (N_11037,N_6728,N_7173);
and U11038 (N_11038,N_6972,N_8337);
nor U11039 (N_11039,N_7568,N_6288);
and U11040 (N_11040,N_8281,N_7253);
or U11041 (N_11041,N_8928,N_6789);
or U11042 (N_11042,N_6298,N_8333);
nand U11043 (N_11043,N_6634,N_6319);
or U11044 (N_11044,N_7806,N_7372);
nor U11045 (N_11045,N_7608,N_7901);
and U11046 (N_11046,N_6066,N_7979);
nor U11047 (N_11047,N_6621,N_6745);
nand U11048 (N_11048,N_7525,N_6482);
nand U11049 (N_11049,N_7130,N_7308);
nand U11050 (N_11050,N_6960,N_6870);
or U11051 (N_11051,N_8714,N_8306);
nand U11052 (N_11052,N_6450,N_8036);
nand U11053 (N_11053,N_7030,N_8342);
or U11054 (N_11054,N_8429,N_6904);
and U11055 (N_11055,N_8593,N_6039);
nand U11056 (N_11056,N_8535,N_8802);
nor U11057 (N_11057,N_6667,N_8128);
nand U11058 (N_11058,N_8154,N_7308);
nand U11059 (N_11059,N_7450,N_7972);
nor U11060 (N_11060,N_7384,N_7117);
nor U11061 (N_11061,N_8429,N_8738);
xnor U11062 (N_11062,N_6914,N_7287);
nand U11063 (N_11063,N_8970,N_8205);
or U11064 (N_11064,N_6921,N_6051);
or U11065 (N_11065,N_7898,N_6994);
or U11066 (N_11066,N_6508,N_6342);
nor U11067 (N_11067,N_7026,N_8388);
nand U11068 (N_11068,N_6011,N_7178);
nand U11069 (N_11069,N_7488,N_8608);
and U11070 (N_11070,N_8934,N_8618);
or U11071 (N_11071,N_7524,N_8847);
or U11072 (N_11072,N_6627,N_7301);
nor U11073 (N_11073,N_6860,N_8960);
and U11074 (N_11074,N_8123,N_8623);
nand U11075 (N_11075,N_7632,N_6555);
nor U11076 (N_11076,N_6574,N_7455);
or U11077 (N_11077,N_8859,N_6195);
or U11078 (N_11078,N_7054,N_6292);
or U11079 (N_11079,N_8549,N_6308);
and U11080 (N_11080,N_6373,N_7692);
or U11081 (N_11081,N_8589,N_7716);
nor U11082 (N_11082,N_8809,N_8526);
or U11083 (N_11083,N_8171,N_7608);
and U11084 (N_11084,N_6069,N_7556);
nand U11085 (N_11085,N_8741,N_8458);
and U11086 (N_11086,N_6186,N_7401);
nor U11087 (N_11087,N_8577,N_7294);
and U11088 (N_11088,N_7731,N_7627);
or U11089 (N_11089,N_6005,N_8884);
or U11090 (N_11090,N_6940,N_8901);
or U11091 (N_11091,N_6818,N_7567);
and U11092 (N_11092,N_6603,N_6452);
nand U11093 (N_11093,N_7256,N_7699);
and U11094 (N_11094,N_7523,N_8260);
nor U11095 (N_11095,N_7652,N_8806);
xnor U11096 (N_11096,N_8196,N_8973);
xor U11097 (N_11097,N_8734,N_8235);
and U11098 (N_11098,N_8085,N_8199);
nand U11099 (N_11099,N_7049,N_7305);
nand U11100 (N_11100,N_6510,N_6576);
nand U11101 (N_11101,N_8261,N_7292);
nor U11102 (N_11102,N_8683,N_8681);
or U11103 (N_11103,N_7783,N_7899);
and U11104 (N_11104,N_7734,N_8697);
or U11105 (N_11105,N_8905,N_7992);
and U11106 (N_11106,N_6395,N_7659);
nand U11107 (N_11107,N_7273,N_7318);
or U11108 (N_11108,N_8198,N_7498);
nand U11109 (N_11109,N_7357,N_7865);
or U11110 (N_11110,N_8902,N_6121);
nand U11111 (N_11111,N_7081,N_7226);
nor U11112 (N_11112,N_7275,N_7424);
nand U11113 (N_11113,N_8836,N_7360);
or U11114 (N_11114,N_6127,N_8237);
nand U11115 (N_11115,N_6725,N_7712);
nor U11116 (N_11116,N_7900,N_8103);
nand U11117 (N_11117,N_8337,N_6312);
or U11118 (N_11118,N_8684,N_8946);
nor U11119 (N_11119,N_6367,N_7784);
nand U11120 (N_11120,N_7710,N_6632);
or U11121 (N_11121,N_8033,N_7444);
nor U11122 (N_11122,N_6567,N_6854);
nor U11123 (N_11123,N_6462,N_6997);
nand U11124 (N_11124,N_7673,N_6329);
nand U11125 (N_11125,N_8232,N_7446);
and U11126 (N_11126,N_6792,N_6028);
nand U11127 (N_11127,N_7442,N_8226);
nor U11128 (N_11128,N_6250,N_7557);
nand U11129 (N_11129,N_8235,N_7140);
nand U11130 (N_11130,N_7974,N_8741);
and U11131 (N_11131,N_8309,N_7754);
and U11132 (N_11132,N_8358,N_6481);
nand U11133 (N_11133,N_8229,N_8303);
or U11134 (N_11134,N_8286,N_7711);
and U11135 (N_11135,N_7170,N_7730);
nand U11136 (N_11136,N_6015,N_6260);
nor U11137 (N_11137,N_6136,N_6011);
or U11138 (N_11138,N_7673,N_8781);
and U11139 (N_11139,N_6273,N_8118);
xor U11140 (N_11140,N_7513,N_7257);
or U11141 (N_11141,N_6337,N_8586);
or U11142 (N_11142,N_7504,N_7547);
nand U11143 (N_11143,N_6087,N_6814);
nor U11144 (N_11144,N_6329,N_7413);
nor U11145 (N_11145,N_8609,N_7137);
or U11146 (N_11146,N_7591,N_8348);
and U11147 (N_11147,N_6278,N_6820);
nor U11148 (N_11148,N_7804,N_8001);
nand U11149 (N_11149,N_8319,N_6761);
nand U11150 (N_11150,N_7079,N_7336);
nand U11151 (N_11151,N_8632,N_7509);
nand U11152 (N_11152,N_6678,N_6554);
and U11153 (N_11153,N_8614,N_8526);
nor U11154 (N_11154,N_8620,N_6762);
nor U11155 (N_11155,N_6888,N_8418);
xnor U11156 (N_11156,N_6110,N_8203);
nand U11157 (N_11157,N_7481,N_8484);
nor U11158 (N_11158,N_7751,N_6927);
or U11159 (N_11159,N_6490,N_8195);
or U11160 (N_11160,N_8152,N_6609);
or U11161 (N_11161,N_6192,N_6530);
or U11162 (N_11162,N_7013,N_7565);
and U11163 (N_11163,N_6774,N_6280);
nand U11164 (N_11164,N_6216,N_8942);
and U11165 (N_11165,N_7500,N_8939);
or U11166 (N_11166,N_6489,N_6970);
nand U11167 (N_11167,N_6358,N_8578);
and U11168 (N_11168,N_8474,N_7106);
or U11169 (N_11169,N_8482,N_8821);
xnor U11170 (N_11170,N_7210,N_6535);
and U11171 (N_11171,N_7272,N_7505);
nand U11172 (N_11172,N_8389,N_7951);
and U11173 (N_11173,N_8847,N_7956);
and U11174 (N_11174,N_8139,N_7307);
nor U11175 (N_11175,N_8958,N_7787);
nor U11176 (N_11176,N_7920,N_8468);
nand U11177 (N_11177,N_7085,N_6945);
and U11178 (N_11178,N_6379,N_6191);
and U11179 (N_11179,N_7815,N_6617);
nand U11180 (N_11180,N_6087,N_8417);
nand U11181 (N_11181,N_7703,N_6950);
nand U11182 (N_11182,N_8151,N_8392);
nand U11183 (N_11183,N_8083,N_6360);
nor U11184 (N_11184,N_8422,N_8880);
nand U11185 (N_11185,N_8486,N_8802);
and U11186 (N_11186,N_6262,N_7967);
nor U11187 (N_11187,N_6082,N_6854);
or U11188 (N_11188,N_7247,N_7966);
nor U11189 (N_11189,N_8485,N_6149);
and U11190 (N_11190,N_7628,N_8070);
nor U11191 (N_11191,N_6898,N_7468);
and U11192 (N_11192,N_7642,N_7280);
nand U11193 (N_11193,N_6825,N_7298);
or U11194 (N_11194,N_8273,N_7700);
nor U11195 (N_11195,N_8728,N_8824);
nand U11196 (N_11196,N_7849,N_6542);
nor U11197 (N_11197,N_7795,N_7266);
nand U11198 (N_11198,N_6438,N_8794);
or U11199 (N_11199,N_6565,N_6886);
or U11200 (N_11200,N_7878,N_6490);
or U11201 (N_11201,N_6098,N_7552);
nand U11202 (N_11202,N_8046,N_7046);
nor U11203 (N_11203,N_6667,N_8237);
nor U11204 (N_11204,N_7109,N_6109);
nand U11205 (N_11205,N_6602,N_6754);
or U11206 (N_11206,N_8385,N_7896);
and U11207 (N_11207,N_7009,N_8302);
nor U11208 (N_11208,N_6248,N_6433);
and U11209 (N_11209,N_8819,N_7411);
or U11210 (N_11210,N_7324,N_6713);
or U11211 (N_11211,N_8890,N_6109);
nand U11212 (N_11212,N_6028,N_7597);
and U11213 (N_11213,N_8062,N_8476);
and U11214 (N_11214,N_8523,N_7408);
and U11215 (N_11215,N_8754,N_7838);
or U11216 (N_11216,N_8935,N_7163);
or U11217 (N_11217,N_6643,N_6371);
and U11218 (N_11218,N_7892,N_8917);
nand U11219 (N_11219,N_6113,N_7440);
and U11220 (N_11220,N_7228,N_7748);
nand U11221 (N_11221,N_6311,N_6494);
nor U11222 (N_11222,N_8737,N_6414);
nor U11223 (N_11223,N_8943,N_6035);
and U11224 (N_11224,N_8245,N_7584);
or U11225 (N_11225,N_6093,N_6348);
or U11226 (N_11226,N_8482,N_7233);
nand U11227 (N_11227,N_8110,N_6000);
and U11228 (N_11228,N_7769,N_6208);
nand U11229 (N_11229,N_8464,N_6521);
or U11230 (N_11230,N_7437,N_8613);
nor U11231 (N_11231,N_6880,N_8540);
or U11232 (N_11232,N_8744,N_8331);
or U11233 (N_11233,N_8518,N_7830);
and U11234 (N_11234,N_6981,N_7292);
nor U11235 (N_11235,N_8968,N_8245);
or U11236 (N_11236,N_8828,N_7238);
or U11237 (N_11237,N_6158,N_6364);
or U11238 (N_11238,N_8247,N_7036);
nor U11239 (N_11239,N_6958,N_7730);
and U11240 (N_11240,N_7697,N_8268);
or U11241 (N_11241,N_7364,N_8615);
or U11242 (N_11242,N_8082,N_7237);
or U11243 (N_11243,N_7032,N_7707);
nor U11244 (N_11244,N_8733,N_8963);
and U11245 (N_11245,N_6364,N_8552);
or U11246 (N_11246,N_8505,N_6552);
nor U11247 (N_11247,N_6015,N_6713);
and U11248 (N_11248,N_6921,N_8283);
nand U11249 (N_11249,N_7300,N_8061);
and U11250 (N_11250,N_8027,N_6633);
and U11251 (N_11251,N_6126,N_6498);
nor U11252 (N_11252,N_7050,N_8721);
or U11253 (N_11253,N_6831,N_7345);
nand U11254 (N_11254,N_7456,N_7618);
nor U11255 (N_11255,N_7447,N_8187);
and U11256 (N_11256,N_6778,N_8844);
nor U11257 (N_11257,N_6926,N_7387);
or U11258 (N_11258,N_8656,N_7460);
nor U11259 (N_11259,N_7420,N_7941);
or U11260 (N_11260,N_6832,N_7342);
nand U11261 (N_11261,N_6572,N_6083);
and U11262 (N_11262,N_8074,N_8813);
nand U11263 (N_11263,N_6207,N_6334);
and U11264 (N_11264,N_8245,N_6250);
nand U11265 (N_11265,N_7399,N_6551);
nand U11266 (N_11266,N_8763,N_6990);
and U11267 (N_11267,N_8613,N_8977);
nand U11268 (N_11268,N_6854,N_8616);
nand U11269 (N_11269,N_8253,N_7130);
nor U11270 (N_11270,N_8716,N_8775);
or U11271 (N_11271,N_7339,N_6130);
or U11272 (N_11272,N_7112,N_7464);
or U11273 (N_11273,N_8689,N_7610);
and U11274 (N_11274,N_6757,N_7254);
nor U11275 (N_11275,N_8988,N_7751);
nor U11276 (N_11276,N_7682,N_7134);
and U11277 (N_11277,N_8560,N_7499);
nand U11278 (N_11278,N_6876,N_7199);
nor U11279 (N_11279,N_8021,N_7245);
and U11280 (N_11280,N_8493,N_7170);
and U11281 (N_11281,N_7198,N_8503);
nor U11282 (N_11282,N_8046,N_7980);
and U11283 (N_11283,N_8573,N_7114);
and U11284 (N_11284,N_6893,N_8729);
and U11285 (N_11285,N_7910,N_6430);
nor U11286 (N_11286,N_8362,N_7170);
and U11287 (N_11287,N_8526,N_8525);
nand U11288 (N_11288,N_8712,N_8884);
or U11289 (N_11289,N_6472,N_7208);
nand U11290 (N_11290,N_6147,N_8909);
or U11291 (N_11291,N_7115,N_7501);
and U11292 (N_11292,N_8353,N_7376);
nand U11293 (N_11293,N_7642,N_7630);
and U11294 (N_11294,N_8326,N_6880);
or U11295 (N_11295,N_7204,N_8265);
nor U11296 (N_11296,N_6904,N_7561);
and U11297 (N_11297,N_6733,N_8300);
and U11298 (N_11298,N_6928,N_7840);
or U11299 (N_11299,N_6114,N_7434);
and U11300 (N_11300,N_8562,N_7380);
nor U11301 (N_11301,N_7339,N_7763);
and U11302 (N_11302,N_8043,N_8724);
nor U11303 (N_11303,N_8836,N_6758);
and U11304 (N_11304,N_6503,N_8129);
nand U11305 (N_11305,N_6793,N_6795);
and U11306 (N_11306,N_8128,N_8057);
nand U11307 (N_11307,N_7747,N_6717);
nor U11308 (N_11308,N_8773,N_8448);
and U11309 (N_11309,N_6843,N_7542);
nor U11310 (N_11310,N_6946,N_7459);
nand U11311 (N_11311,N_7960,N_8118);
and U11312 (N_11312,N_6005,N_7593);
nand U11313 (N_11313,N_6740,N_8166);
or U11314 (N_11314,N_7977,N_6933);
or U11315 (N_11315,N_7259,N_6345);
or U11316 (N_11316,N_8835,N_7551);
nand U11317 (N_11317,N_8832,N_6213);
or U11318 (N_11318,N_6267,N_6633);
nor U11319 (N_11319,N_7281,N_8353);
and U11320 (N_11320,N_7179,N_8701);
and U11321 (N_11321,N_8149,N_8228);
nor U11322 (N_11322,N_6635,N_6754);
and U11323 (N_11323,N_7630,N_8131);
and U11324 (N_11324,N_6789,N_7907);
nand U11325 (N_11325,N_7418,N_6966);
and U11326 (N_11326,N_6148,N_6099);
or U11327 (N_11327,N_7698,N_6886);
nand U11328 (N_11328,N_7694,N_7065);
and U11329 (N_11329,N_6576,N_6675);
and U11330 (N_11330,N_7668,N_7623);
and U11331 (N_11331,N_8938,N_6879);
or U11332 (N_11332,N_8318,N_6225);
or U11333 (N_11333,N_8172,N_8134);
nand U11334 (N_11334,N_7289,N_8608);
or U11335 (N_11335,N_7162,N_6278);
nor U11336 (N_11336,N_6271,N_7946);
or U11337 (N_11337,N_8073,N_6251);
nor U11338 (N_11338,N_6552,N_7908);
and U11339 (N_11339,N_6337,N_7918);
nand U11340 (N_11340,N_6324,N_8062);
nand U11341 (N_11341,N_6542,N_6360);
and U11342 (N_11342,N_6375,N_7075);
nand U11343 (N_11343,N_8784,N_6059);
nor U11344 (N_11344,N_7386,N_8180);
and U11345 (N_11345,N_7280,N_7472);
nand U11346 (N_11346,N_8943,N_8064);
and U11347 (N_11347,N_8443,N_7014);
nor U11348 (N_11348,N_8700,N_7631);
or U11349 (N_11349,N_6191,N_6039);
and U11350 (N_11350,N_7932,N_7128);
nand U11351 (N_11351,N_6785,N_8765);
nand U11352 (N_11352,N_6241,N_7411);
nor U11353 (N_11353,N_6815,N_7834);
or U11354 (N_11354,N_7890,N_8556);
nor U11355 (N_11355,N_8587,N_6503);
or U11356 (N_11356,N_6258,N_8847);
or U11357 (N_11357,N_7220,N_7498);
and U11358 (N_11358,N_7936,N_7843);
and U11359 (N_11359,N_8201,N_6011);
and U11360 (N_11360,N_8301,N_8471);
and U11361 (N_11361,N_7207,N_7892);
or U11362 (N_11362,N_7219,N_7367);
nor U11363 (N_11363,N_8805,N_7937);
and U11364 (N_11364,N_6197,N_7455);
and U11365 (N_11365,N_8162,N_7472);
nand U11366 (N_11366,N_7848,N_6958);
nand U11367 (N_11367,N_7452,N_6076);
or U11368 (N_11368,N_7682,N_7745);
and U11369 (N_11369,N_6630,N_7581);
nor U11370 (N_11370,N_7884,N_8495);
or U11371 (N_11371,N_7925,N_6180);
nand U11372 (N_11372,N_8499,N_8757);
xor U11373 (N_11373,N_8001,N_8432);
and U11374 (N_11374,N_6935,N_8565);
and U11375 (N_11375,N_7290,N_7623);
and U11376 (N_11376,N_8844,N_7018);
or U11377 (N_11377,N_8937,N_8967);
nand U11378 (N_11378,N_7115,N_7894);
or U11379 (N_11379,N_8981,N_7429);
or U11380 (N_11380,N_6575,N_6993);
and U11381 (N_11381,N_8543,N_7864);
or U11382 (N_11382,N_7034,N_8915);
or U11383 (N_11383,N_7916,N_8434);
and U11384 (N_11384,N_6196,N_7330);
or U11385 (N_11385,N_8704,N_6672);
nor U11386 (N_11386,N_8137,N_8720);
or U11387 (N_11387,N_6021,N_8760);
nand U11388 (N_11388,N_6900,N_6651);
nand U11389 (N_11389,N_6065,N_7414);
nor U11390 (N_11390,N_7728,N_6972);
or U11391 (N_11391,N_7095,N_8925);
and U11392 (N_11392,N_8418,N_8050);
and U11393 (N_11393,N_7586,N_7724);
and U11394 (N_11394,N_8425,N_7544);
or U11395 (N_11395,N_8365,N_7349);
nand U11396 (N_11396,N_8686,N_6668);
and U11397 (N_11397,N_8994,N_7214);
and U11398 (N_11398,N_6603,N_8986);
and U11399 (N_11399,N_7101,N_6963);
nor U11400 (N_11400,N_7393,N_8935);
or U11401 (N_11401,N_7751,N_6555);
or U11402 (N_11402,N_6309,N_6931);
or U11403 (N_11403,N_7709,N_8193);
or U11404 (N_11404,N_7798,N_7582);
and U11405 (N_11405,N_6123,N_7171);
nor U11406 (N_11406,N_8610,N_6777);
nand U11407 (N_11407,N_8137,N_8949);
and U11408 (N_11408,N_8205,N_7450);
or U11409 (N_11409,N_8409,N_6770);
nor U11410 (N_11410,N_8648,N_8564);
nor U11411 (N_11411,N_8674,N_8169);
nand U11412 (N_11412,N_8311,N_8674);
or U11413 (N_11413,N_8347,N_6236);
and U11414 (N_11414,N_7598,N_7782);
and U11415 (N_11415,N_8186,N_7912);
nand U11416 (N_11416,N_7111,N_7064);
nand U11417 (N_11417,N_7833,N_8975);
and U11418 (N_11418,N_7738,N_7369);
nor U11419 (N_11419,N_6861,N_6291);
nor U11420 (N_11420,N_8380,N_8180);
and U11421 (N_11421,N_6645,N_8864);
nand U11422 (N_11422,N_8609,N_8930);
nor U11423 (N_11423,N_8241,N_7121);
and U11424 (N_11424,N_8402,N_8857);
nand U11425 (N_11425,N_7889,N_8166);
and U11426 (N_11426,N_7479,N_7302);
or U11427 (N_11427,N_6731,N_6235);
or U11428 (N_11428,N_7953,N_6404);
nor U11429 (N_11429,N_7922,N_8103);
nand U11430 (N_11430,N_6392,N_7968);
nor U11431 (N_11431,N_8578,N_8873);
or U11432 (N_11432,N_8289,N_8396);
nor U11433 (N_11433,N_8460,N_6971);
or U11434 (N_11434,N_7672,N_8620);
and U11435 (N_11435,N_6728,N_6117);
nand U11436 (N_11436,N_6978,N_8812);
nor U11437 (N_11437,N_6720,N_6692);
nand U11438 (N_11438,N_8374,N_6837);
or U11439 (N_11439,N_8914,N_6713);
nor U11440 (N_11440,N_8675,N_6390);
nand U11441 (N_11441,N_8801,N_6184);
nor U11442 (N_11442,N_8635,N_8098);
nand U11443 (N_11443,N_7315,N_6229);
nor U11444 (N_11444,N_7219,N_8664);
nor U11445 (N_11445,N_8883,N_6942);
and U11446 (N_11446,N_7616,N_6363);
xor U11447 (N_11447,N_6421,N_6931);
and U11448 (N_11448,N_7219,N_7669);
or U11449 (N_11449,N_6588,N_6919);
nand U11450 (N_11450,N_6193,N_8003);
nand U11451 (N_11451,N_7103,N_8559);
or U11452 (N_11452,N_6870,N_8226);
nand U11453 (N_11453,N_6498,N_8593);
and U11454 (N_11454,N_7156,N_7319);
nand U11455 (N_11455,N_8142,N_7778);
nor U11456 (N_11456,N_7303,N_8683);
nor U11457 (N_11457,N_7451,N_6562);
nor U11458 (N_11458,N_7317,N_7223);
nor U11459 (N_11459,N_7961,N_7484);
or U11460 (N_11460,N_6307,N_6722);
and U11461 (N_11461,N_7599,N_6294);
nor U11462 (N_11462,N_6064,N_7154);
and U11463 (N_11463,N_7234,N_8994);
and U11464 (N_11464,N_7478,N_8717);
or U11465 (N_11465,N_7671,N_7063);
or U11466 (N_11466,N_6213,N_8395);
and U11467 (N_11467,N_8337,N_6305);
nor U11468 (N_11468,N_6865,N_6644);
xnor U11469 (N_11469,N_8897,N_7511);
nor U11470 (N_11470,N_8772,N_7653);
or U11471 (N_11471,N_7200,N_8225);
and U11472 (N_11472,N_7531,N_7083);
nand U11473 (N_11473,N_6220,N_6165);
xor U11474 (N_11474,N_7969,N_6536);
nor U11475 (N_11475,N_6342,N_6209);
nor U11476 (N_11476,N_6454,N_7303);
nor U11477 (N_11477,N_8191,N_6879);
and U11478 (N_11478,N_8583,N_8003);
nand U11479 (N_11479,N_7774,N_8691);
nand U11480 (N_11480,N_8286,N_8250);
nor U11481 (N_11481,N_7397,N_8824);
and U11482 (N_11482,N_6153,N_8445);
and U11483 (N_11483,N_8837,N_6026);
nor U11484 (N_11484,N_7830,N_8730);
nand U11485 (N_11485,N_6143,N_7646);
nor U11486 (N_11486,N_7392,N_8318);
nor U11487 (N_11487,N_6983,N_7631);
nor U11488 (N_11488,N_6951,N_6788);
nor U11489 (N_11489,N_6459,N_7249);
and U11490 (N_11490,N_6869,N_7567);
or U11491 (N_11491,N_6431,N_8339);
nor U11492 (N_11492,N_7925,N_6689);
nand U11493 (N_11493,N_6929,N_6844);
nor U11494 (N_11494,N_7888,N_8629);
nor U11495 (N_11495,N_7853,N_7511);
nand U11496 (N_11496,N_7760,N_7615);
nor U11497 (N_11497,N_6678,N_7107);
and U11498 (N_11498,N_7978,N_7532);
nor U11499 (N_11499,N_6118,N_8189);
or U11500 (N_11500,N_7099,N_7986);
nand U11501 (N_11501,N_8873,N_8410);
and U11502 (N_11502,N_8863,N_8270);
or U11503 (N_11503,N_8073,N_7578);
nand U11504 (N_11504,N_7939,N_8155);
and U11505 (N_11505,N_8307,N_6270);
nor U11506 (N_11506,N_7550,N_8037);
nor U11507 (N_11507,N_8017,N_8165);
or U11508 (N_11508,N_8614,N_6780);
nor U11509 (N_11509,N_7104,N_6079);
nand U11510 (N_11510,N_8962,N_6431);
nand U11511 (N_11511,N_6510,N_8362);
or U11512 (N_11512,N_8364,N_7922);
or U11513 (N_11513,N_8715,N_6168);
and U11514 (N_11514,N_6201,N_6674);
and U11515 (N_11515,N_8896,N_7365);
and U11516 (N_11516,N_8503,N_8998);
nor U11517 (N_11517,N_8969,N_7766);
and U11518 (N_11518,N_7982,N_6271);
nor U11519 (N_11519,N_8978,N_7361);
nor U11520 (N_11520,N_8138,N_7491);
and U11521 (N_11521,N_6962,N_6895);
nand U11522 (N_11522,N_6365,N_7597);
and U11523 (N_11523,N_8921,N_7691);
and U11524 (N_11524,N_6153,N_8523);
and U11525 (N_11525,N_8768,N_6860);
nand U11526 (N_11526,N_7815,N_8192);
nor U11527 (N_11527,N_8377,N_7697);
or U11528 (N_11528,N_8194,N_8449);
nand U11529 (N_11529,N_8806,N_7649);
or U11530 (N_11530,N_7575,N_6685);
xnor U11531 (N_11531,N_6450,N_8336);
nor U11532 (N_11532,N_8574,N_7443);
or U11533 (N_11533,N_6752,N_6521);
or U11534 (N_11534,N_7797,N_8302);
nor U11535 (N_11535,N_8555,N_8774);
nand U11536 (N_11536,N_8249,N_8605);
nor U11537 (N_11537,N_6935,N_8913);
nand U11538 (N_11538,N_7460,N_7786);
nand U11539 (N_11539,N_8869,N_6577);
nand U11540 (N_11540,N_8042,N_6707);
nand U11541 (N_11541,N_6438,N_7699);
nor U11542 (N_11542,N_8557,N_8199);
nor U11543 (N_11543,N_8632,N_6404);
nor U11544 (N_11544,N_7572,N_8438);
nor U11545 (N_11545,N_6584,N_7360);
nor U11546 (N_11546,N_7023,N_6659);
nand U11547 (N_11547,N_6621,N_8059);
nand U11548 (N_11548,N_6778,N_8822);
or U11549 (N_11549,N_6191,N_8402);
xnor U11550 (N_11550,N_7634,N_6360);
nand U11551 (N_11551,N_7272,N_7338);
nand U11552 (N_11552,N_8696,N_6693);
and U11553 (N_11553,N_6108,N_6024);
nand U11554 (N_11554,N_7109,N_6636);
and U11555 (N_11555,N_7207,N_8769);
nor U11556 (N_11556,N_8029,N_8467);
nand U11557 (N_11557,N_8200,N_8413);
nor U11558 (N_11558,N_8922,N_8976);
and U11559 (N_11559,N_6650,N_8484);
and U11560 (N_11560,N_6869,N_6932);
nor U11561 (N_11561,N_7337,N_8823);
and U11562 (N_11562,N_6405,N_7896);
or U11563 (N_11563,N_8405,N_6628);
nand U11564 (N_11564,N_6963,N_6911);
or U11565 (N_11565,N_7015,N_6049);
nand U11566 (N_11566,N_7583,N_8387);
nor U11567 (N_11567,N_6698,N_6596);
nor U11568 (N_11568,N_6243,N_6354);
or U11569 (N_11569,N_7176,N_7027);
and U11570 (N_11570,N_8025,N_6181);
and U11571 (N_11571,N_6176,N_7708);
nand U11572 (N_11572,N_6647,N_7273);
nand U11573 (N_11573,N_8275,N_7086);
and U11574 (N_11574,N_7076,N_6921);
nor U11575 (N_11575,N_7313,N_6858);
nor U11576 (N_11576,N_7262,N_8712);
nand U11577 (N_11577,N_6108,N_7931);
or U11578 (N_11578,N_7646,N_8341);
or U11579 (N_11579,N_7292,N_8735);
and U11580 (N_11580,N_8857,N_7072);
and U11581 (N_11581,N_6899,N_8184);
nor U11582 (N_11582,N_6059,N_7904);
or U11583 (N_11583,N_8194,N_7175);
or U11584 (N_11584,N_6330,N_8858);
nand U11585 (N_11585,N_8473,N_6450);
or U11586 (N_11586,N_6286,N_7162);
or U11587 (N_11587,N_8605,N_6053);
nand U11588 (N_11588,N_7150,N_6485);
nor U11589 (N_11589,N_8183,N_6599);
and U11590 (N_11590,N_6467,N_8874);
nor U11591 (N_11591,N_8877,N_7181);
nand U11592 (N_11592,N_6378,N_8200);
or U11593 (N_11593,N_8285,N_7936);
and U11594 (N_11594,N_7144,N_8809);
or U11595 (N_11595,N_6291,N_6777);
nand U11596 (N_11596,N_6187,N_8663);
nor U11597 (N_11597,N_6851,N_8210);
nor U11598 (N_11598,N_8876,N_8804);
and U11599 (N_11599,N_8062,N_7937);
and U11600 (N_11600,N_8248,N_6028);
nand U11601 (N_11601,N_6673,N_6382);
nand U11602 (N_11602,N_8853,N_6714);
or U11603 (N_11603,N_6346,N_8954);
nor U11604 (N_11604,N_7538,N_8377);
nor U11605 (N_11605,N_7206,N_7389);
nand U11606 (N_11606,N_6287,N_7093);
or U11607 (N_11607,N_7638,N_8935);
nor U11608 (N_11608,N_8356,N_7320);
nand U11609 (N_11609,N_6632,N_8969);
nor U11610 (N_11610,N_7693,N_6832);
nor U11611 (N_11611,N_6200,N_7578);
and U11612 (N_11612,N_6437,N_6591);
or U11613 (N_11613,N_6623,N_6555);
and U11614 (N_11614,N_6009,N_6985);
or U11615 (N_11615,N_6504,N_8725);
nand U11616 (N_11616,N_8678,N_8028);
and U11617 (N_11617,N_7010,N_8957);
or U11618 (N_11618,N_8793,N_6783);
or U11619 (N_11619,N_6764,N_7533);
nand U11620 (N_11620,N_6042,N_7150);
xnor U11621 (N_11621,N_8568,N_6336);
nor U11622 (N_11622,N_7953,N_8749);
nand U11623 (N_11623,N_7404,N_6794);
or U11624 (N_11624,N_8618,N_7174);
or U11625 (N_11625,N_7947,N_7684);
and U11626 (N_11626,N_8215,N_8062);
or U11627 (N_11627,N_8856,N_6753);
and U11628 (N_11628,N_7829,N_6276);
or U11629 (N_11629,N_8540,N_7541);
and U11630 (N_11630,N_6080,N_6615);
nand U11631 (N_11631,N_7212,N_8276);
and U11632 (N_11632,N_7650,N_8751);
or U11633 (N_11633,N_8278,N_7525);
or U11634 (N_11634,N_8194,N_8250);
and U11635 (N_11635,N_8581,N_6965);
or U11636 (N_11636,N_8964,N_7381);
and U11637 (N_11637,N_6437,N_6115);
nor U11638 (N_11638,N_7752,N_8148);
nand U11639 (N_11639,N_7176,N_7262);
and U11640 (N_11640,N_6647,N_6337);
nor U11641 (N_11641,N_7616,N_8571);
nor U11642 (N_11642,N_8833,N_7445);
and U11643 (N_11643,N_8984,N_8777);
nor U11644 (N_11644,N_7971,N_6177);
nor U11645 (N_11645,N_7295,N_7262);
or U11646 (N_11646,N_7287,N_7820);
or U11647 (N_11647,N_6668,N_7048);
or U11648 (N_11648,N_7459,N_8318);
or U11649 (N_11649,N_8259,N_7947);
nand U11650 (N_11650,N_7384,N_7110);
and U11651 (N_11651,N_8085,N_7137);
nor U11652 (N_11652,N_6186,N_6342);
nor U11653 (N_11653,N_6187,N_8561);
and U11654 (N_11654,N_6556,N_6570);
or U11655 (N_11655,N_7619,N_7063);
nor U11656 (N_11656,N_8701,N_6153);
nand U11657 (N_11657,N_6148,N_6606);
nor U11658 (N_11658,N_8980,N_8521);
or U11659 (N_11659,N_7560,N_8700);
and U11660 (N_11660,N_7394,N_6066);
nor U11661 (N_11661,N_7566,N_7488);
or U11662 (N_11662,N_7472,N_6078);
and U11663 (N_11663,N_7776,N_7955);
or U11664 (N_11664,N_7961,N_7096);
nor U11665 (N_11665,N_6552,N_7046);
nor U11666 (N_11666,N_7383,N_7931);
nor U11667 (N_11667,N_6282,N_8454);
or U11668 (N_11668,N_8314,N_8513);
nor U11669 (N_11669,N_8468,N_7785);
nor U11670 (N_11670,N_6669,N_7600);
and U11671 (N_11671,N_6112,N_7502);
nand U11672 (N_11672,N_8528,N_7128);
or U11673 (N_11673,N_6962,N_8917);
or U11674 (N_11674,N_8429,N_8073);
and U11675 (N_11675,N_7466,N_7661);
nor U11676 (N_11676,N_8690,N_6094);
nand U11677 (N_11677,N_8401,N_8834);
nor U11678 (N_11678,N_6241,N_6836);
xor U11679 (N_11679,N_6135,N_6196);
and U11680 (N_11680,N_8082,N_6606);
nand U11681 (N_11681,N_7407,N_8854);
and U11682 (N_11682,N_8808,N_6443);
nor U11683 (N_11683,N_7389,N_7172);
nand U11684 (N_11684,N_6538,N_7548);
or U11685 (N_11685,N_8468,N_7764);
and U11686 (N_11686,N_7083,N_8886);
nand U11687 (N_11687,N_7807,N_8833);
and U11688 (N_11688,N_6329,N_6578);
or U11689 (N_11689,N_8824,N_6388);
xnor U11690 (N_11690,N_6621,N_6902);
and U11691 (N_11691,N_6415,N_8175);
nor U11692 (N_11692,N_6548,N_6505);
nor U11693 (N_11693,N_6256,N_8366);
nor U11694 (N_11694,N_8981,N_7507);
and U11695 (N_11695,N_6743,N_7389);
and U11696 (N_11696,N_6938,N_8318);
and U11697 (N_11697,N_6008,N_8331);
nor U11698 (N_11698,N_8953,N_8620);
and U11699 (N_11699,N_8194,N_7687);
or U11700 (N_11700,N_6891,N_7427);
and U11701 (N_11701,N_6298,N_7236);
and U11702 (N_11702,N_6395,N_6063);
nor U11703 (N_11703,N_8067,N_6327);
nand U11704 (N_11704,N_6075,N_7981);
nand U11705 (N_11705,N_7470,N_6344);
or U11706 (N_11706,N_6051,N_8201);
or U11707 (N_11707,N_7902,N_6241);
nor U11708 (N_11708,N_6967,N_6484);
nor U11709 (N_11709,N_8748,N_8353);
and U11710 (N_11710,N_8613,N_8965);
nand U11711 (N_11711,N_6894,N_7267);
nor U11712 (N_11712,N_7476,N_7485);
nand U11713 (N_11713,N_8875,N_7394);
and U11714 (N_11714,N_7065,N_6097);
nand U11715 (N_11715,N_7354,N_7252);
or U11716 (N_11716,N_8214,N_6618);
nand U11717 (N_11717,N_8792,N_6178);
nand U11718 (N_11718,N_8204,N_8631);
nand U11719 (N_11719,N_7140,N_6416);
nor U11720 (N_11720,N_7678,N_8830);
nand U11721 (N_11721,N_6341,N_8764);
nor U11722 (N_11722,N_8156,N_8579);
nand U11723 (N_11723,N_8545,N_8919);
nand U11724 (N_11724,N_7785,N_7658);
nand U11725 (N_11725,N_8593,N_8600);
or U11726 (N_11726,N_6675,N_6296);
and U11727 (N_11727,N_8759,N_7709);
or U11728 (N_11728,N_6781,N_8872);
nor U11729 (N_11729,N_8597,N_6935);
nand U11730 (N_11730,N_8686,N_6215);
nand U11731 (N_11731,N_8134,N_8589);
nor U11732 (N_11732,N_8407,N_8267);
nor U11733 (N_11733,N_6550,N_8197);
and U11734 (N_11734,N_6263,N_7701);
and U11735 (N_11735,N_8067,N_8956);
nor U11736 (N_11736,N_7190,N_8740);
nor U11737 (N_11737,N_6210,N_7658);
and U11738 (N_11738,N_8255,N_8780);
nand U11739 (N_11739,N_8818,N_8833);
nor U11740 (N_11740,N_6161,N_8254);
and U11741 (N_11741,N_7014,N_6818);
nor U11742 (N_11742,N_7487,N_8565);
nor U11743 (N_11743,N_8698,N_7840);
nand U11744 (N_11744,N_6285,N_6442);
or U11745 (N_11745,N_8300,N_6360);
or U11746 (N_11746,N_8627,N_8267);
or U11747 (N_11747,N_8197,N_7174);
or U11748 (N_11748,N_8142,N_7933);
and U11749 (N_11749,N_7777,N_6127);
or U11750 (N_11750,N_7614,N_7286);
or U11751 (N_11751,N_7887,N_8627);
or U11752 (N_11752,N_8435,N_6547);
or U11753 (N_11753,N_7728,N_8157);
and U11754 (N_11754,N_8291,N_7344);
and U11755 (N_11755,N_7933,N_6144);
or U11756 (N_11756,N_8649,N_6933);
nor U11757 (N_11757,N_6161,N_7156);
or U11758 (N_11758,N_8258,N_6555);
nor U11759 (N_11759,N_6651,N_6491);
or U11760 (N_11760,N_7366,N_7913);
and U11761 (N_11761,N_8125,N_7348);
nor U11762 (N_11762,N_6775,N_7043);
or U11763 (N_11763,N_8258,N_6557);
and U11764 (N_11764,N_6071,N_6385);
and U11765 (N_11765,N_6981,N_7606);
and U11766 (N_11766,N_6039,N_6973);
or U11767 (N_11767,N_6983,N_6907);
or U11768 (N_11768,N_6563,N_7948);
nand U11769 (N_11769,N_6166,N_7612);
nor U11770 (N_11770,N_8214,N_6649);
or U11771 (N_11771,N_7184,N_6516);
nor U11772 (N_11772,N_8911,N_8325);
and U11773 (N_11773,N_8456,N_8144);
nand U11774 (N_11774,N_6284,N_6954);
or U11775 (N_11775,N_8070,N_6960);
nor U11776 (N_11776,N_7586,N_7609);
nand U11777 (N_11777,N_7376,N_7622);
or U11778 (N_11778,N_8660,N_8056);
and U11779 (N_11779,N_6719,N_7551);
nor U11780 (N_11780,N_7973,N_8544);
nand U11781 (N_11781,N_6482,N_6579);
nor U11782 (N_11782,N_6830,N_8642);
and U11783 (N_11783,N_6960,N_8538);
or U11784 (N_11784,N_7170,N_6401);
nand U11785 (N_11785,N_6277,N_8443);
or U11786 (N_11786,N_6512,N_8044);
nor U11787 (N_11787,N_6453,N_6035);
nor U11788 (N_11788,N_7027,N_6239);
or U11789 (N_11789,N_6098,N_6791);
or U11790 (N_11790,N_6682,N_8205);
or U11791 (N_11791,N_8382,N_7786);
nand U11792 (N_11792,N_6603,N_8350);
nand U11793 (N_11793,N_7602,N_7060);
and U11794 (N_11794,N_6031,N_7999);
nor U11795 (N_11795,N_6318,N_8318);
or U11796 (N_11796,N_6024,N_7903);
and U11797 (N_11797,N_8469,N_8797);
or U11798 (N_11798,N_8807,N_6428);
nand U11799 (N_11799,N_6621,N_8092);
nor U11800 (N_11800,N_6984,N_8898);
nor U11801 (N_11801,N_7327,N_6741);
or U11802 (N_11802,N_7630,N_7613);
nor U11803 (N_11803,N_6875,N_8023);
nor U11804 (N_11804,N_7692,N_6059);
nand U11805 (N_11805,N_6419,N_7597);
or U11806 (N_11806,N_7043,N_6754);
or U11807 (N_11807,N_6860,N_7189);
nand U11808 (N_11808,N_7323,N_6998);
or U11809 (N_11809,N_8646,N_7569);
or U11810 (N_11810,N_7080,N_8701);
or U11811 (N_11811,N_8585,N_7127);
and U11812 (N_11812,N_6594,N_6909);
nand U11813 (N_11813,N_7114,N_6697);
nand U11814 (N_11814,N_7951,N_6185);
or U11815 (N_11815,N_7835,N_8215);
nor U11816 (N_11816,N_8553,N_7621);
or U11817 (N_11817,N_7364,N_7394);
nor U11818 (N_11818,N_7523,N_8839);
or U11819 (N_11819,N_8840,N_6042);
nand U11820 (N_11820,N_8216,N_6774);
or U11821 (N_11821,N_8101,N_7318);
nand U11822 (N_11822,N_6823,N_6231);
nand U11823 (N_11823,N_6501,N_7508);
and U11824 (N_11824,N_7051,N_7818);
or U11825 (N_11825,N_7131,N_7369);
and U11826 (N_11826,N_8287,N_8123);
and U11827 (N_11827,N_6088,N_7162);
nand U11828 (N_11828,N_7455,N_8321);
xnor U11829 (N_11829,N_8713,N_7531);
nand U11830 (N_11830,N_8505,N_6052);
and U11831 (N_11831,N_6415,N_8117);
and U11832 (N_11832,N_8322,N_7242);
nor U11833 (N_11833,N_6063,N_6066);
or U11834 (N_11834,N_8874,N_7949);
nor U11835 (N_11835,N_6074,N_8880);
and U11836 (N_11836,N_6319,N_8016);
and U11837 (N_11837,N_8619,N_7734);
nand U11838 (N_11838,N_7576,N_7704);
and U11839 (N_11839,N_8494,N_8814);
nand U11840 (N_11840,N_7957,N_8232);
nor U11841 (N_11841,N_8049,N_6697);
nor U11842 (N_11842,N_8918,N_6959);
or U11843 (N_11843,N_6547,N_6718);
or U11844 (N_11844,N_8109,N_7892);
nand U11845 (N_11845,N_7515,N_8919);
or U11846 (N_11846,N_6366,N_6522);
and U11847 (N_11847,N_8426,N_7939);
or U11848 (N_11848,N_7160,N_6945);
and U11849 (N_11849,N_8026,N_6370);
or U11850 (N_11850,N_7420,N_8779);
and U11851 (N_11851,N_8572,N_6342);
or U11852 (N_11852,N_6635,N_8579);
or U11853 (N_11853,N_7525,N_6056);
nor U11854 (N_11854,N_8996,N_6553);
nor U11855 (N_11855,N_6017,N_6394);
and U11856 (N_11856,N_6337,N_6201);
nor U11857 (N_11857,N_7591,N_7255);
nand U11858 (N_11858,N_8243,N_8175);
nor U11859 (N_11859,N_7261,N_6817);
nor U11860 (N_11860,N_8305,N_7525);
nor U11861 (N_11861,N_7711,N_8445);
nand U11862 (N_11862,N_8483,N_7275);
nand U11863 (N_11863,N_6689,N_8132);
and U11864 (N_11864,N_7800,N_7196);
and U11865 (N_11865,N_6114,N_7381);
nor U11866 (N_11866,N_8315,N_8391);
or U11867 (N_11867,N_6811,N_8799);
nand U11868 (N_11868,N_6393,N_8998);
nand U11869 (N_11869,N_6171,N_8257);
xor U11870 (N_11870,N_7590,N_8186);
nand U11871 (N_11871,N_7557,N_8712);
nand U11872 (N_11872,N_6913,N_8413);
and U11873 (N_11873,N_7475,N_7489);
nand U11874 (N_11874,N_7500,N_6047);
nor U11875 (N_11875,N_7855,N_6367);
nor U11876 (N_11876,N_6627,N_7277);
nor U11877 (N_11877,N_6646,N_6933);
and U11878 (N_11878,N_7447,N_7291);
or U11879 (N_11879,N_7095,N_8915);
or U11880 (N_11880,N_6670,N_8293);
nor U11881 (N_11881,N_7775,N_8482);
and U11882 (N_11882,N_8227,N_7627);
nor U11883 (N_11883,N_7754,N_8275);
nand U11884 (N_11884,N_6732,N_6722);
nand U11885 (N_11885,N_6270,N_7349);
nand U11886 (N_11886,N_6004,N_6399);
nand U11887 (N_11887,N_8781,N_7916);
or U11888 (N_11888,N_8418,N_8246);
nor U11889 (N_11889,N_6222,N_7571);
nor U11890 (N_11890,N_8361,N_7796);
or U11891 (N_11891,N_6127,N_8565);
or U11892 (N_11892,N_7446,N_6687);
nor U11893 (N_11893,N_8442,N_6843);
nor U11894 (N_11894,N_6398,N_7453);
nand U11895 (N_11895,N_7737,N_8630);
or U11896 (N_11896,N_6367,N_8919);
nand U11897 (N_11897,N_6086,N_8559);
and U11898 (N_11898,N_6500,N_8277);
nor U11899 (N_11899,N_8886,N_7546);
nand U11900 (N_11900,N_6001,N_6553);
or U11901 (N_11901,N_8957,N_6916);
nand U11902 (N_11902,N_8815,N_8402);
nor U11903 (N_11903,N_6693,N_8162);
or U11904 (N_11904,N_8325,N_7578);
or U11905 (N_11905,N_6024,N_7071);
or U11906 (N_11906,N_6442,N_6355);
nand U11907 (N_11907,N_8242,N_8429);
and U11908 (N_11908,N_7990,N_6905);
nor U11909 (N_11909,N_8160,N_7443);
or U11910 (N_11910,N_6167,N_6922);
nor U11911 (N_11911,N_8610,N_7847);
and U11912 (N_11912,N_7524,N_7779);
nand U11913 (N_11913,N_7931,N_8550);
or U11914 (N_11914,N_6153,N_7608);
or U11915 (N_11915,N_8412,N_7534);
nand U11916 (N_11916,N_6140,N_8834);
nand U11917 (N_11917,N_8969,N_8128);
and U11918 (N_11918,N_8056,N_8630);
and U11919 (N_11919,N_6672,N_6560);
and U11920 (N_11920,N_8041,N_6503);
or U11921 (N_11921,N_7750,N_7242);
and U11922 (N_11922,N_7262,N_8102);
nor U11923 (N_11923,N_6371,N_8445);
nand U11924 (N_11924,N_6838,N_8913);
or U11925 (N_11925,N_6356,N_6773);
and U11926 (N_11926,N_8592,N_7232);
nand U11927 (N_11927,N_6475,N_6450);
nand U11928 (N_11928,N_6771,N_6530);
and U11929 (N_11929,N_6282,N_6938);
or U11930 (N_11930,N_6677,N_6637);
or U11931 (N_11931,N_7127,N_6093);
nor U11932 (N_11932,N_7257,N_8630);
nor U11933 (N_11933,N_8098,N_8373);
and U11934 (N_11934,N_6038,N_6702);
nor U11935 (N_11935,N_7895,N_7482);
or U11936 (N_11936,N_8103,N_7386);
and U11937 (N_11937,N_6437,N_8664);
or U11938 (N_11938,N_6701,N_7492);
nand U11939 (N_11939,N_6632,N_6486);
or U11940 (N_11940,N_8163,N_6632);
and U11941 (N_11941,N_7152,N_6805);
or U11942 (N_11942,N_8436,N_8949);
nand U11943 (N_11943,N_6586,N_8731);
and U11944 (N_11944,N_6526,N_6426);
and U11945 (N_11945,N_8622,N_8154);
and U11946 (N_11946,N_8258,N_6404);
nand U11947 (N_11947,N_8025,N_7602);
or U11948 (N_11948,N_6999,N_7557);
nor U11949 (N_11949,N_8339,N_7748);
and U11950 (N_11950,N_8876,N_6410);
and U11951 (N_11951,N_7572,N_6723);
and U11952 (N_11952,N_6813,N_6257);
nor U11953 (N_11953,N_8482,N_7992);
nor U11954 (N_11954,N_6617,N_7816);
or U11955 (N_11955,N_7377,N_8121);
and U11956 (N_11956,N_6477,N_7013);
and U11957 (N_11957,N_8414,N_8479);
and U11958 (N_11958,N_7520,N_8069);
or U11959 (N_11959,N_6516,N_6762);
nor U11960 (N_11960,N_7823,N_7689);
nand U11961 (N_11961,N_6242,N_8001);
nor U11962 (N_11962,N_8926,N_7647);
nand U11963 (N_11963,N_7370,N_8725);
xor U11964 (N_11964,N_6432,N_7652);
or U11965 (N_11965,N_6942,N_6162);
nor U11966 (N_11966,N_7138,N_7167);
nand U11967 (N_11967,N_6870,N_8944);
nand U11968 (N_11968,N_8071,N_6888);
nor U11969 (N_11969,N_7684,N_8480);
or U11970 (N_11970,N_6213,N_6716);
nand U11971 (N_11971,N_7609,N_7200);
nand U11972 (N_11972,N_6601,N_8379);
or U11973 (N_11973,N_7865,N_6791);
nand U11974 (N_11974,N_8283,N_7109);
nand U11975 (N_11975,N_7445,N_8989);
or U11976 (N_11976,N_7804,N_8525);
and U11977 (N_11977,N_6844,N_6414);
and U11978 (N_11978,N_8764,N_7652);
nand U11979 (N_11979,N_6895,N_6769);
and U11980 (N_11980,N_8872,N_7103);
nor U11981 (N_11981,N_6021,N_6964);
or U11982 (N_11982,N_7498,N_7874);
and U11983 (N_11983,N_6900,N_7943);
nand U11984 (N_11984,N_6354,N_7036);
and U11985 (N_11985,N_8529,N_8695);
nor U11986 (N_11986,N_7288,N_7777);
nor U11987 (N_11987,N_6064,N_7332);
nand U11988 (N_11988,N_6634,N_7695);
nand U11989 (N_11989,N_7140,N_6205);
and U11990 (N_11990,N_6294,N_6051);
nand U11991 (N_11991,N_8547,N_8019);
and U11992 (N_11992,N_8962,N_8511);
nand U11993 (N_11993,N_7408,N_7895);
nand U11994 (N_11994,N_7302,N_7185);
nand U11995 (N_11995,N_8486,N_8675);
or U11996 (N_11996,N_7669,N_6055);
or U11997 (N_11997,N_8177,N_6719);
or U11998 (N_11998,N_6224,N_8914);
and U11999 (N_11999,N_6209,N_8176);
and U12000 (N_12000,N_9219,N_9190);
nor U12001 (N_12001,N_10325,N_9842);
nand U12002 (N_12002,N_10300,N_11690);
and U12003 (N_12003,N_9047,N_9350);
or U12004 (N_12004,N_11252,N_9306);
nand U12005 (N_12005,N_9073,N_11098);
nand U12006 (N_12006,N_9176,N_9434);
nor U12007 (N_12007,N_11930,N_11243);
nand U12008 (N_12008,N_9260,N_10823);
xnor U12009 (N_12009,N_10954,N_10492);
and U12010 (N_12010,N_9556,N_11912);
xnor U12011 (N_12011,N_10677,N_10500);
or U12012 (N_12012,N_10479,N_11414);
nor U12013 (N_12013,N_11706,N_10662);
nand U12014 (N_12014,N_9206,N_11457);
or U12015 (N_12015,N_10771,N_9756);
nor U12016 (N_12016,N_11322,N_11046);
nor U12017 (N_12017,N_10777,N_9252);
and U12018 (N_12018,N_10498,N_10312);
nor U12019 (N_12019,N_11184,N_11900);
nand U12020 (N_12020,N_11174,N_11927);
and U12021 (N_12021,N_11559,N_9711);
nor U12022 (N_12022,N_11526,N_9932);
nand U12023 (N_12023,N_10806,N_9214);
or U12024 (N_12024,N_11855,N_9765);
and U12025 (N_12025,N_11859,N_10458);
and U12026 (N_12026,N_10612,N_9376);
and U12027 (N_12027,N_10999,N_10485);
or U12028 (N_12028,N_9955,N_9486);
and U12029 (N_12029,N_9374,N_11581);
nand U12030 (N_12030,N_11281,N_11217);
or U12031 (N_12031,N_11135,N_9873);
and U12032 (N_12032,N_10246,N_9970);
or U12033 (N_12033,N_9263,N_10747);
nand U12034 (N_12034,N_9002,N_11911);
nand U12035 (N_12035,N_9622,N_9850);
or U12036 (N_12036,N_10045,N_10603);
and U12037 (N_12037,N_9428,N_9222);
nor U12038 (N_12038,N_10390,N_11817);
nand U12039 (N_12039,N_9918,N_9293);
and U12040 (N_12040,N_11109,N_9657);
or U12041 (N_12041,N_11774,N_11522);
nor U12042 (N_12042,N_9417,N_10124);
or U12043 (N_12043,N_9490,N_9150);
nand U12044 (N_12044,N_11040,N_9691);
nand U12045 (N_12045,N_11007,N_9045);
nand U12046 (N_12046,N_11049,N_9217);
or U12047 (N_12047,N_10464,N_9167);
or U12048 (N_12048,N_10765,N_10809);
nor U12049 (N_12049,N_10863,N_11171);
nand U12050 (N_12050,N_11875,N_9915);
or U12051 (N_12051,N_11851,N_9695);
nand U12052 (N_12052,N_11002,N_9975);
nor U12053 (N_12053,N_9478,N_10201);
or U12054 (N_12054,N_11975,N_9840);
nand U12055 (N_12055,N_10258,N_10210);
or U12056 (N_12056,N_11208,N_11833);
or U12057 (N_12057,N_9089,N_9141);
and U12058 (N_12058,N_10889,N_9626);
and U12059 (N_12059,N_9269,N_9198);
or U12060 (N_12060,N_10556,N_11988);
and U12061 (N_12061,N_10102,N_11654);
nor U12062 (N_12062,N_10003,N_9193);
nor U12063 (N_12063,N_9347,N_9759);
and U12064 (N_12064,N_9271,N_11982);
nand U12065 (N_12065,N_11257,N_9249);
and U12066 (N_12066,N_11455,N_11778);
nor U12067 (N_12067,N_11383,N_10964);
or U12068 (N_12068,N_11972,N_9580);
nor U12069 (N_12069,N_9629,N_11352);
or U12070 (N_12070,N_11715,N_9220);
and U12071 (N_12071,N_11905,N_11665);
and U12072 (N_12072,N_10017,N_11441);
nand U12073 (N_12073,N_11783,N_9609);
or U12074 (N_12074,N_10669,N_10558);
nand U12075 (N_12075,N_10749,N_10927);
and U12076 (N_12076,N_10647,N_9292);
nand U12077 (N_12077,N_9785,N_9940);
or U12078 (N_12078,N_9127,N_11807);
or U12079 (N_12079,N_9126,N_10590);
or U12080 (N_12080,N_9020,N_9123);
and U12081 (N_12081,N_11820,N_9606);
nor U12082 (N_12082,N_11646,N_10065);
or U12083 (N_12083,N_10750,N_9816);
nand U12084 (N_12084,N_9369,N_10744);
nand U12085 (N_12085,N_11513,N_10366);
or U12086 (N_12086,N_11018,N_9648);
nand U12087 (N_12087,N_9725,N_10900);
and U12088 (N_12088,N_9037,N_10281);
nand U12089 (N_12089,N_10851,N_11753);
or U12090 (N_12090,N_9329,N_9651);
and U12091 (N_12091,N_9281,N_11494);
nor U12092 (N_12092,N_9267,N_10444);
or U12093 (N_12093,N_11662,N_10235);
nand U12094 (N_12094,N_10256,N_9697);
nand U12095 (N_12095,N_9439,N_9088);
nor U12096 (N_12096,N_10338,N_9420);
or U12097 (N_12097,N_11205,N_10955);
or U12098 (N_12098,N_9851,N_11590);
nand U12099 (N_12099,N_10972,N_11255);
nand U12100 (N_12100,N_9853,N_9564);
and U12101 (N_12101,N_11587,N_9508);
nand U12102 (N_12102,N_10730,N_11499);
and U12103 (N_12103,N_9031,N_11969);
or U12104 (N_12104,N_10232,N_11287);
or U12105 (N_12105,N_11661,N_11775);
or U12106 (N_12106,N_9465,N_9750);
and U12107 (N_12107,N_10421,N_9603);
nand U12108 (N_12108,N_9114,N_11471);
or U12109 (N_12109,N_10410,N_10026);
or U12110 (N_12110,N_10654,N_10882);
nor U12111 (N_12111,N_11970,N_11449);
nor U12112 (N_12112,N_10845,N_9158);
or U12113 (N_12113,N_10212,N_11932);
nand U12114 (N_12114,N_9837,N_11923);
nor U12115 (N_12115,N_11563,N_9474);
or U12116 (N_12116,N_10249,N_9327);
and U12117 (N_12117,N_9264,N_10700);
nand U12118 (N_12118,N_9341,N_10143);
nand U12119 (N_12119,N_10101,N_11584);
nor U12120 (N_12120,N_11539,N_9589);
nor U12121 (N_12121,N_9442,N_11680);
or U12122 (N_12122,N_10920,N_11582);
or U12123 (N_12123,N_11592,N_10878);
nand U12124 (N_12124,N_11541,N_11645);
and U12125 (N_12125,N_9361,N_11472);
nor U12126 (N_12126,N_10119,N_10664);
and U12127 (N_12127,N_10394,N_11042);
nand U12128 (N_12128,N_9524,N_11360);
nand U12129 (N_12129,N_9243,N_10270);
and U12130 (N_12130,N_10541,N_10261);
nand U12131 (N_12131,N_11728,N_10908);
and U12132 (N_12132,N_11566,N_10014);
or U12133 (N_12133,N_9344,N_10893);
nand U12134 (N_12134,N_9944,N_9999);
nand U12135 (N_12135,N_9160,N_11218);
nor U12136 (N_12136,N_9381,N_10983);
nor U12137 (N_12137,N_10468,N_10666);
and U12138 (N_12138,N_10299,N_10551);
or U12139 (N_12139,N_9772,N_10623);
and U12140 (N_12140,N_11426,N_11015);
nand U12141 (N_12141,N_10775,N_9519);
or U12142 (N_12142,N_9734,N_11073);
or U12143 (N_12143,N_9803,N_9470);
xor U12144 (N_12144,N_11325,N_10455);
or U12145 (N_12145,N_11643,N_11967);
nor U12146 (N_12146,N_9515,N_11087);
nand U12147 (N_12147,N_10167,N_10808);
or U12148 (N_12148,N_9244,N_9030);
nand U12149 (N_12149,N_10204,N_11253);
and U12150 (N_12150,N_9109,N_9107);
nand U12151 (N_12151,N_9138,N_10611);
nor U12152 (N_12152,N_10745,N_9746);
nand U12153 (N_12153,N_10118,N_9684);
or U12154 (N_12154,N_10020,N_11622);
or U12155 (N_12155,N_10607,N_9122);
nor U12156 (N_12156,N_10287,N_9782);
or U12157 (N_12157,N_9038,N_9987);
nor U12158 (N_12158,N_10172,N_11258);
nand U12159 (N_12159,N_9188,N_11231);
and U12160 (N_12160,N_9621,N_9388);
nor U12161 (N_12161,N_11734,N_9120);
nor U12162 (N_12162,N_9427,N_9407);
and U12163 (N_12163,N_11843,N_10573);
nor U12164 (N_12164,N_10233,N_11300);
and U12165 (N_12165,N_10701,N_11892);
or U12166 (N_12166,N_11210,N_10027);
nand U12167 (N_12167,N_11175,N_9003);
nand U12168 (N_12168,N_10919,N_9674);
nor U12169 (N_12169,N_9592,N_9462);
or U12170 (N_12170,N_11798,N_11053);
and U12171 (N_12171,N_10778,N_11810);
nand U12172 (N_12172,N_9886,N_9957);
or U12173 (N_12173,N_9399,N_9348);
nand U12174 (N_12174,N_10594,N_11428);
nand U12175 (N_12175,N_11245,N_11291);
or U12176 (N_12176,N_11378,N_10083);
nand U12177 (N_12177,N_10052,N_9686);
or U12178 (N_12178,N_11038,N_9218);
nand U12179 (N_12179,N_11216,N_10398);
nand U12180 (N_12180,N_10169,N_10307);
and U12181 (N_12181,N_11437,N_11897);
nor U12182 (N_12182,N_10296,N_10079);
nor U12183 (N_12183,N_10819,N_9964);
or U12184 (N_12184,N_11844,N_10040);
nor U12185 (N_12185,N_9647,N_10591);
xor U12186 (N_12186,N_11395,N_11968);
or U12187 (N_12187,N_11211,N_11404);
nor U12188 (N_12188,N_9298,N_10066);
nand U12189 (N_12189,N_9831,N_11704);
and U12190 (N_12190,N_10129,N_11543);
nand U12191 (N_12191,N_9812,N_10311);
nand U12192 (N_12192,N_9480,N_10141);
nor U12193 (N_12193,N_11848,N_10397);
or U12194 (N_12194,N_10571,N_11066);
nand U12195 (N_12195,N_9018,N_11373);
and U12196 (N_12196,N_10567,N_9085);
or U12197 (N_12197,N_9937,N_11256);
xor U12198 (N_12198,N_10274,N_9009);
or U12199 (N_12199,N_9845,N_11037);
nand U12200 (N_12200,N_11168,N_11286);
nand U12201 (N_12201,N_9854,N_11146);
or U12202 (N_12202,N_9316,N_11830);
or U12203 (N_12203,N_9547,N_11185);
or U12204 (N_12204,N_11781,N_9332);
nor U12205 (N_12205,N_10377,N_9954);
and U12206 (N_12206,N_10980,N_10511);
and U12207 (N_12207,N_11978,N_11931);
and U12208 (N_12208,N_11574,N_10460);
and U12209 (N_12209,N_10953,N_9634);
nor U12210 (N_12210,N_10137,N_11689);
or U12211 (N_12211,N_10153,N_10095);
or U12212 (N_12212,N_10604,N_10523);
nor U12213 (N_12213,N_11531,N_10534);
nand U12214 (N_12214,N_10696,N_11172);
and U12215 (N_12215,N_11347,N_9340);
nand U12216 (N_12216,N_9755,N_9710);
nor U12217 (N_12217,N_10886,N_9542);
nor U12218 (N_12218,N_11752,N_10271);
nand U12219 (N_12219,N_9640,N_11572);
or U12220 (N_12220,N_10224,N_10984);
nand U12221 (N_12221,N_9092,N_10437);
and U12222 (N_12222,N_10076,N_9458);
nor U12223 (N_12223,N_9602,N_9393);
and U12224 (N_12224,N_10685,N_11886);
or U12225 (N_12225,N_10405,N_11248);
nand U12226 (N_12226,N_9041,N_10152);
or U12227 (N_12227,N_11074,N_11341);
or U12228 (N_12228,N_9501,N_9857);
nor U12229 (N_12229,N_11957,N_10525);
nor U12230 (N_12230,N_11307,N_10071);
nor U12231 (N_12231,N_10930,N_9270);
or U12232 (N_12232,N_11283,N_9367);
and U12233 (N_12233,N_11319,N_11655);
nor U12234 (N_12234,N_9923,N_9482);
and U12235 (N_12235,N_10636,N_10158);
xor U12236 (N_12236,N_10554,N_9163);
or U12237 (N_12237,N_9920,N_9087);
and U12238 (N_12238,N_10379,N_10108);
or U12239 (N_12239,N_9973,N_9929);
nand U12240 (N_12240,N_11213,N_10733);
and U12241 (N_12241,N_10514,N_11236);
nand U12242 (N_12242,N_11818,N_11435);
and U12243 (N_12243,N_9537,N_9021);
and U12244 (N_12244,N_11839,N_11928);
or U12245 (N_12245,N_9174,N_11101);
nand U12246 (N_12246,N_11115,N_11129);
nand U12247 (N_12247,N_11506,N_9694);
and U12248 (N_12248,N_9632,N_10347);
and U12249 (N_12249,N_11951,N_11889);
nand U12250 (N_12250,N_9950,N_11460);
or U12251 (N_12251,N_9299,N_10668);
or U12252 (N_12252,N_11890,N_11351);
or U12253 (N_12253,N_11310,N_9867);
nand U12254 (N_12254,N_10100,N_10349);
and U12255 (N_12255,N_10752,N_9246);
nor U12256 (N_12256,N_11759,N_10881);
nand U12257 (N_12257,N_10796,N_11529);
nand U12258 (N_12258,N_10504,N_11878);
or U12259 (N_12259,N_9377,N_9847);
and U12260 (N_12260,N_9716,N_10859);
or U12261 (N_12261,N_9383,N_11901);
or U12262 (N_12262,N_11197,N_9467);
nand U12263 (N_12263,N_11861,N_10853);
xnor U12264 (N_12264,N_9836,N_11024);
xnor U12265 (N_12265,N_11062,N_10635);
or U12266 (N_12266,N_9406,N_11051);
or U12267 (N_12267,N_10284,N_11362);
nand U12268 (N_12268,N_10030,N_11882);
nand U12269 (N_12269,N_11732,N_10401);
xnor U12270 (N_12270,N_10241,N_10907);
nor U12271 (N_12271,N_10621,N_9908);
or U12272 (N_12272,N_11102,N_10880);
or U12273 (N_12273,N_11749,N_9770);
nand U12274 (N_12274,N_9146,N_11834);
or U12275 (N_12275,N_10005,N_10113);
nand U12276 (N_12276,N_11589,N_10112);
nand U12277 (N_12277,N_11944,N_9389);
or U12278 (N_12278,N_11381,N_10157);
nand U12279 (N_12279,N_9289,N_11595);
or U12280 (N_12280,N_11239,N_9414);
nor U12281 (N_12281,N_10434,N_9693);
xnor U12282 (N_12282,N_9029,N_9051);
or U12283 (N_12283,N_9487,N_11560);
or U12284 (N_12284,N_11324,N_9305);
and U12285 (N_12285,N_10731,N_11880);
nand U12286 (N_12286,N_11459,N_10561);
nand U12287 (N_12287,N_9865,N_11993);
nor U12288 (N_12288,N_11617,N_11298);
or U12289 (N_12289,N_10002,N_9535);
and U12290 (N_12290,N_9313,N_10387);
or U12291 (N_12291,N_11666,N_9525);
and U12292 (N_12292,N_10988,N_10317);
nor U12293 (N_12293,N_9481,N_10675);
and U12294 (N_12294,N_10430,N_10507);
or U12295 (N_12295,N_10412,N_9492);
nand U12296 (N_12296,N_9712,N_11123);
or U12297 (N_12297,N_11108,N_11241);
nand U12298 (N_12298,N_11536,N_11685);
nor U12299 (N_12299,N_11361,N_10861);
or U12300 (N_12300,N_11675,N_9498);
or U12301 (N_12301,N_9262,N_11423);
or U12302 (N_12302,N_11357,N_11093);
nand U12303 (N_12303,N_10593,N_10251);
nand U12304 (N_12304,N_11162,N_9620);
or U12305 (N_12305,N_11676,N_10238);
nor U12306 (N_12306,N_11926,N_10588);
nand U12307 (N_12307,N_9904,N_10478);
nand U12308 (N_12308,N_10480,N_10419);
and U12309 (N_12309,N_10179,N_9721);
or U12310 (N_12310,N_9274,N_9485);
nand U12311 (N_12311,N_9397,N_11400);
and U12312 (N_12312,N_11346,N_9660);
nor U12313 (N_12313,N_11551,N_9581);
nand U12314 (N_12314,N_10579,N_9360);
nand U12315 (N_12315,N_9223,N_11027);
nand U12316 (N_12316,N_9074,N_11940);
and U12317 (N_12317,N_10392,N_10164);
or U12318 (N_12318,N_9363,N_11275);
or U12319 (N_12319,N_10252,N_11682);
nor U12320 (N_12320,N_11372,N_9878);
and U12321 (N_12321,N_9473,N_9096);
or U12322 (N_12322,N_9758,N_10773);
nand U12323 (N_12323,N_9717,N_9359);
nor U12324 (N_12324,N_10459,N_10860);
nand U12325 (N_12325,N_11660,N_10820);
nand U12326 (N_12326,N_11363,N_10342);
and U12327 (N_12327,N_9726,N_9512);
nor U12328 (N_12328,N_10209,N_9914);
nor U12329 (N_12329,N_10735,N_10265);
and U12330 (N_12330,N_9196,N_10957);
nand U12331 (N_12331,N_11165,N_9210);
nand U12332 (N_12332,N_11091,N_9131);
and U12333 (N_12333,N_10409,N_10807);
nor U12334 (N_12334,N_10963,N_9658);
nand U12335 (N_12335,N_9186,N_10520);
nor U12336 (N_12336,N_9022,N_11639);
nand U12337 (N_12337,N_11517,N_9189);
or U12338 (N_12338,N_9328,N_11534);
and U12339 (N_12339,N_11672,N_10839);
and U12340 (N_12340,N_10849,N_11816);
nand U12341 (N_12341,N_9215,N_10996);
nor U12342 (N_12342,N_11222,N_11910);
and U12343 (N_12343,N_10484,N_9538);
and U12344 (N_12344,N_9539,N_9978);
nand U12345 (N_12345,N_9216,N_9221);
nand U12346 (N_12346,N_10916,N_9991);
and U12347 (N_12347,N_10191,N_11720);
or U12348 (N_12348,N_9101,N_11260);
nor U12349 (N_12349,N_11994,N_11189);
and U12350 (N_12350,N_11048,N_9799);
nor U12351 (N_12351,N_11226,N_9148);
nor U12352 (N_12352,N_9333,N_10446);
nand U12353 (N_12353,N_10794,N_11155);
nand U12354 (N_12354,N_9204,N_9810);
nand U12355 (N_12355,N_11354,N_10146);
xnor U12356 (N_12356,N_10931,N_10121);
nand U12357 (N_12357,N_11393,N_10103);
or U12358 (N_12358,N_11983,N_11125);
and U12359 (N_12359,N_10902,N_9049);
nand U12360 (N_12360,N_10208,N_9476);
nand U12361 (N_12361,N_10117,N_9988);
nand U12362 (N_12362,N_10423,N_11621);
or U12363 (N_12363,N_9506,N_11057);
and U12364 (N_12364,N_11415,N_10407);
and U12365 (N_12365,N_9457,N_9690);
xnor U12366 (N_12366,N_10609,N_9549);
and U12367 (N_12367,N_9769,N_10308);
and U12368 (N_12368,N_10709,N_11332);
and U12369 (N_12369,N_9833,N_11960);
nand U12370 (N_12370,N_11398,N_9272);
and U12371 (N_12371,N_10189,N_11620);
and U12372 (N_12372,N_11605,N_9111);
and U12373 (N_12373,N_10531,N_9410);
nor U12374 (N_12374,N_9962,N_10802);
or U12375 (N_12375,N_10560,N_10742);
or U12376 (N_12376,N_9094,N_10574);
or U12377 (N_12377,N_9133,N_10063);
or U12378 (N_12378,N_11762,N_9390);
or U12379 (N_12379,N_11710,N_11036);
nor U12380 (N_12380,N_10337,N_11489);
nand U12381 (N_12381,N_9773,N_10294);
or U12382 (N_12382,N_9144,N_11773);
or U12383 (N_12383,N_11899,N_9208);
and U12384 (N_12384,N_11338,N_11937);
nor U12385 (N_12385,N_9172,N_9628);
nor U12386 (N_12386,N_10199,N_9555);
nand U12387 (N_12387,N_9752,N_9533);
nor U12388 (N_12388,N_10358,N_10470);
nor U12389 (N_12389,N_11219,N_10833);
and U12390 (N_12390,N_9766,N_9273);
and U12391 (N_12391,N_10537,N_9455);
nand U12392 (N_12392,N_11670,N_10530);
or U12393 (N_12393,N_9423,N_10564);
nand U12394 (N_12394,N_10938,N_9308);
nor U12395 (N_12395,N_9874,N_9916);
and U12396 (N_12396,N_11263,N_10216);
nand U12397 (N_12397,N_11823,N_11012);
nor U12398 (N_12398,N_9990,N_9735);
nor U12399 (N_12399,N_10789,N_10123);
xnor U12400 (N_12400,N_9813,N_11288);
nand U12401 (N_12401,N_9205,N_10368);
nor U12402 (N_12402,N_10687,N_9996);
nor U12403 (N_12403,N_11079,N_10724);
or U12404 (N_12404,N_11964,N_9044);
or U12405 (N_12405,N_10648,N_9830);
and U12406 (N_12406,N_9641,N_11741);
nand U12407 (N_12407,N_9529,N_9948);
or U12408 (N_12408,N_9043,N_9972);
or U12409 (N_12409,N_10457,N_9702);
and U12410 (N_12410,N_10671,N_10891);
nand U12411 (N_12411,N_10967,N_11344);
nor U12412 (N_12412,N_11694,N_10427);
and U12413 (N_12413,N_9013,N_9019);
or U12414 (N_12414,N_10280,N_11829);
nor U12415 (N_12415,N_11274,N_11456);
nor U12416 (N_12416,N_9510,N_10847);
nor U12417 (N_12417,N_11005,N_9719);
nor U12418 (N_12418,N_10761,N_11092);
and U12419 (N_12419,N_9164,N_11955);
and U12420 (N_12420,N_11597,N_10046);
nand U12421 (N_12421,N_9998,N_9741);
and U12422 (N_12422,N_10068,N_10417);
or U12423 (N_12423,N_11140,N_11081);
and U12424 (N_12424,N_11512,N_11105);
or U12425 (N_12425,N_9024,N_10254);
nor U12426 (N_12426,N_10139,N_10581);
nand U12427 (N_12427,N_10658,N_11417);
xnor U12428 (N_12428,N_9429,N_9681);
xor U12429 (N_12429,N_9334,N_10023);
or U12430 (N_12430,N_9953,N_9718);
and U12431 (N_12431,N_10592,N_10712);
and U12432 (N_12432,N_11232,N_9370);
and U12433 (N_12433,N_9067,N_10350);
nand U12434 (N_12434,N_9228,N_11262);
nand U12435 (N_12435,N_10070,N_9528);
and U12436 (N_12436,N_11616,N_10895);
and U12437 (N_12437,N_10160,N_11047);
or U12438 (N_12438,N_9097,N_9614);
nand U12439 (N_12439,N_10353,N_9154);
or U12440 (N_12440,N_11793,N_11995);
nand U12441 (N_12441,N_11945,N_10959);
and U12442 (N_12442,N_9568,N_11637);
nand U12443 (N_12443,N_10924,N_10862);
nor U12444 (N_12444,N_10008,N_11853);
or U12445 (N_12445,N_9665,N_9892);
xor U12446 (N_12446,N_10832,N_11863);
and U12447 (N_12447,N_11348,N_10998);
nor U12448 (N_12448,N_10683,N_10184);
and U12449 (N_12449,N_11424,N_11458);
and U12450 (N_12450,N_9559,N_11633);
nor U12451 (N_12451,N_11201,N_10577);
or U12452 (N_12452,N_9491,N_10653);
nor U12453 (N_12453,N_9426,N_10760);
or U12454 (N_12454,N_10659,N_9128);
or U12455 (N_12455,N_10111,N_10130);
nor U12456 (N_12456,N_11925,N_10132);
or U12457 (N_12457,N_11445,N_9859);
or U12458 (N_12458,N_10722,N_10243);
nand U12459 (N_12459,N_9590,N_10422);
and U12460 (N_12460,N_10306,N_9500);
and U12461 (N_12461,N_11285,N_10566);
nand U12462 (N_12462,N_11657,N_9662);
nor U12463 (N_12463,N_10227,N_9655);
and U12464 (N_12464,N_10180,N_11904);
and U12465 (N_12465,N_10741,N_11238);
or U12466 (N_12466,N_11755,N_10856);
and U12467 (N_12467,N_11118,N_9303);
nand U12468 (N_12468,N_11772,N_9604);
and U12469 (N_12469,N_11837,N_10483);
xor U12470 (N_12470,N_9282,N_9295);
nor U12471 (N_12471,N_10266,N_11705);
nor U12472 (N_12472,N_11402,N_9942);
or U12473 (N_12473,N_11693,N_11881);
and U12474 (N_12474,N_10059,N_10770);
or U12475 (N_12475,N_9180,N_11832);
or U12476 (N_12476,N_10034,N_9251);
and U12477 (N_12477,N_11663,N_10801);
and U12478 (N_12478,N_11464,N_9261);
or U12479 (N_12479,N_11750,N_11121);
or U12480 (N_12480,N_9336,N_10006);
and U12481 (N_12481,N_10791,N_9767);
or U12482 (N_12482,N_9532,N_10843);
nor U12483 (N_12483,N_9728,N_9440);
and U12484 (N_12484,N_11919,N_11561);
nand U12485 (N_12485,N_9117,N_10198);
nand U12486 (N_12486,N_9616,N_11822);
nor U12487 (N_12487,N_9939,N_9722);
nand U12488 (N_12488,N_10200,N_9461);
nor U12489 (N_12489,N_10425,N_9312);
or U12490 (N_12490,N_10453,N_9235);
or U12491 (N_12491,N_9472,N_10543);
or U12492 (N_12492,N_10055,N_11814);
nand U12493 (N_12493,N_11153,N_9183);
or U12494 (N_12494,N_11707,N_11467);
nor U12495 (N_12495,N_9540,N_11342);
nand U12496 (N_12496,N_9968,N_11870);
nor U12497 (N_12497,N_11127,N_9432);
nor U12498 (N_12498,N_10196,N_11549);
or U12499 (N_12499,N_9226,N_11902);
or U12500 (N_12500,N_10803,N_11915);
and U12501 (N_12501,N_11941,N_9584);
nor U12502 (N_12502,N_9250,N_9848);
nor U12503 (N_12503,N_9278,N_9777);
nor U12504 (N_12504,N_11343,N_10746);
nor U12505 (N_12505,N_10617,N_9330);
and U12506 (N_12506,N_11751,N_9187);
nor U12507 (N_12507,N_9119,N_10343);
and U12508 (N_12508,N_11273,N_11790);
or U12509 (N_12509,N_9835,N_9910);
and U12510 (N_12510,N_11929,N_10706);
xnor U12511 (N_12511,N_10821,N_9550);
nor U12512 (N_12512,N_9526,N_10759);
and U12513 (N_12513,N_11498,N_10756);
or U12514 (N_12514,N_10024,N_9522);
and U12515 (N_12515,N_11443,N_9801);
nand U12516 (N_12516,N_11913,N_10563);
and U12517 (N_12517,N_11161,N_10161);
and U12518 (N_12518,N_11292,N_10923);
nor U12519 (N_12519,N_11764,N_9424);
xor U12520 (N_12520,N_9827,N_10990);
nor U12521 (N_12521,N_10515,N_9372);
nor U12522 (N_12522,N_9631,N_10877);
and U12523 (N_12523,N_10356,N_11096);
or U12524 (N_12524,N_9520,N_9730);
or U12525 (N_12525,N_11917,N_11134);
nand U12526 (N_12526,N_10903,N_11154);
and U12527 (N_12527,N_9768,N_9656);
and U12528 (N_12528,N_9723,N_10522);
nor U12529 (N_12529,N_9700,N_9063);
nor U12530 (N_12530,N_9011,N_11599);
and U12531 (N_12531,N_10495,N_9479);
and U12532 (N_12532,N_11856,N_9477);
nand U12533 (N_12533,N_9259,N_10641);
and U12534 (N_12534,N_10585,N_9195);
nor U12535 (N_12535,N_9971,N_11011);
nand U12536 (N_12536,N_9325,N_11686);
and U12537 (N_12537,N_10982,N_9319);
or U12538 (N_12538,N_11629,N_10469);
nor U12539 (N_12539,N_10834,N_9653);
or U12540 (N_12540,N_11503,N_9385);
and U12541 (N_12541,N_9304,N_10084);
and U12542 (N_12542,N_9636,N_11841);
nor U12543 (N_12543,N_10451,N_11523);
and U12544 (N_12544,N_9574,N_9353);
or U12545 (N_12545,N_9471,N_10578);
and U12546 (N_12546,N_10672,N_9570);
and U12547 (N_12547,N_10725,N_10089);
nor U12548 (N_12548,N_9623,N_9201);
nand U12549 (N_12549,N_9380,N_9764);
or U12550 (N_12550,N_10267,N_9977);
nor U12551 (N_12551,N_10221,N_11518);
nand U12552 (N_12552,N_10769,N_9368);
or U12553 (N_12553,N_10192,N_10979);
nand U12554 (N_12554,N_10781,N_10064);
nor U12555 (N_12555,N_11234,N_10868);
and U12556 (N_12556,N_11564,N_11063);
nand U12557 (N_12557,N_10651,N_9576);
or U12558 (N_12558,N_10660,N_11004);
nand U12559 (N_12559,N_9342,N_10513);
nor U12560 (N_12560,N_9879,N_9899);
and U12561 (N_12561,N_11515,N_11606);
nand U12562 (N_12562,N_9197,N_9575);
and U12563 (N_12563,N_11006,N_9130);
nor U12564 (N_12564,N_11277,N_11521);
and U12565 (N_12565,N_9106,N_10714);
and U12566 (N_12566,N_10291,N_9014);
nor U12567 (N_12567,N_11683,N_11730);
nor U12568 (N_12568,N_9569,N_9822);
nand U12569 (N_12569,N_10428,N_10763);
nor U12570 (N_12570,N_10029,N_11187);
and U12571 (N_12571,N_11802,N_9371);
nor U12572 (N_12572,N_10690,N_10866);
or U12573 (N_12573,N_9513,N_10941);
nor U12574 (N_12574,N_11337,N_9976);
or U12575 (N_12575,N_9743,N_9704);
or U12576 (N_12576,N_9039,N_9444);
and U12577 (N_12577,N_11193,N_9175);
nand U12578 (N_12578,N_10374,N_9069);
or U12579 (N_12579,N_11405,N_11076);
nor U12580 (N_12580,N_9654,N_9137);
or U12581 (N_12581,N_11504,N_10614);
and U12582 (N_12582,N_11293,N_11309);
nor U12583 (N_12583,N_10831,N_10788);
or U12584 (N_12584,N_11267,N_10628);
or U12585 (N_12585,N_10193,N_11071);
or U12586 (N_12586,N_11664,N_10704);
and U12587 (N_12587,N_11579,N_10968);
nor U12588 (N_12588,N_9639,N_9234);
nand U12589 (N_12589,N_9016,N_9398);
nand U12590 (N_12590,N_9159,N_10155);
nor U12591 (N_12591,N_9185,N_11712);
nor U12592 (N_12592,N_11144,N_10348);
nand U12593 (N_12593,N_11028,N_11647);
and U12594 (N_12594,N_9379,N_10545);
nor U12595 (N_12595,N_11297,N_9757);
or U12596 (N_12596,N_11935,N_9871);
xnor U12597 (N_12597,N_10285,N_11401);
or U12598 (N_12598,N_9807,N_10440);
nand U12599 (N_12599,N_10400,N_9124);
and U12600 (N_12600,N_10663,N_10646);
nand U12601 (N_12601,N_11069,N_9345);
or U12602 (N_12602,N_10098,N_10595);
nand U12603 (N_12603,N_10044,N_11754);
nor U12604 (N_12604,N_9004,N_10632);
and U12605 (N_12605,N_10093,N_10077);
nor U12606 (N_12606,N_9326,N_9170);
and U12607 (N_12607,N_9762,N_10981);
and U12608 (N_12608,N_10830,N_10874);
and U12609 (N_12609,N_11056,N_9708);
nor U12610 (N_12610,N_10892,N_10844);
nand U12611 (N_12611,N_10411,N_9354);
and U12612 (N_12612,N_11711,N_9277);
nand U12613 (N_12613,N_10582,N_11812);
nor U12614 (N_12614,N_10767,N_11502);
and U12615 (N_12615,N_10335,N_11831);
and U12616 (N_12616,N_11461,N_10264);
and U12617 (N_12617,N_11626,N_11763);
and U12618 (N_12618,N_11421,N_10056);
or U12619 (N_12619,N_10471,N_10339);
nand U12620 (N_12620,N_9255,N_11868);
and U12621 (N_12621,N_11760,N_10288);
nand U12622 (N_12622,N_11032,N_9889);
nand U12623 (N_12623,N_10357,N_9742);
nand U12624 (N_12624,N_9203,N_11907);
nor U12625 (N_12625,N_11737,N_11023);
nor U12626 (N_12626,N_11525,N_10226);
nand U12627 (N_12627,N_10415,N_10380);
or U12628 (N_12628,N_9698,N_10864);
xnor U12629 (N_12629,N_10033,N_9211);
or U12630 (N_12630,N_9983,N_11547);
or U12631 (N_12631,N_9514,N_9599);
and U12632 (N_12632,N_10080,N_9033);
nor U12633 (N_12633,N_9994,N_9207);
and U12634 (N_12634,N_9285,N_10674);
and U12635 (N_12635,N_9666,N_11985);
nand U12636 (N_12636,N_10962,N_10734);
nor U12637 (N_12637,N_10010,N_9489);
and U12638 (N_12638,N_10512,N_9143);
or U12639 (N_12639,N_11510,N_11321);
and U12640 (N_12640,N_10073,N_9928);
nand U12641 (N_12641,N_9055,N_11516);
nand U12642 (N_12642,N_10110,N_10126);
or U12643 (N_12643,N_11791,N_11813);
nor U12644 (N_12644,N_10329,N_10042);
nor U12645 (N_12645,N_11656,N_10857);
nand U12646 (N_12646,N_10170,N_11736);
nand U12647 (N_12647,N_9729,N_11483);
and U12648 (N_12648,N_9943,N_11638);
and U12649 (N_12649,N_11583,N_11364);
or U12650 (N_12650,N_10482,N_9373);
or U12651 (N_12651,N_9010,N_10488);
or U12652 (N_12652,N_11151,N_10576);
nand U12653 (N_12653,N_11505,N_11149);
nor U12654 (N_12654,N_10784,N_11490);
and U12655 (N_12655,N_11537,N_9541);
or U12656 (N_12656,N_9321,N_11480);
nor U12657 (N_12657,N_11804,N_10075);
nand U12658 (N_12658,N_9392,N_9213);
or U12659 (N_12659,N_10727,N_11237);
and U12660 (N_12660,N_11299,N_10378);
and U12661 (N_12661,N_9995,N_10645);
and U12662 (N_12662,N_11961,N_11636);
and U12663 (N_12663,N_11203,N_10527);
or U12664 (N_12664,N_10336,N_9403);
nand U12665 (N_12665,N_10565,N_9375);
nand U12666 (N_12666,N_10116,N_9366);
and U12667 (N_12667,N_9026,N_11795);
nand U12668 (N_12668,N_9578,N_10846);
or U12669 (N_12669,N_11658,N_9934);
nand U12670 (N_12670,N_11722,N_11035);
nand U12671 (N_12671,N_11065,N_9256);
nand U12672 (N_12672,N_11713,N_10973);
nor U12673 (N_12673,N_11717,N_10105);
and U12674 (N_12674,N_10004,N_9946);
or U12675 (N_12675,N_9938,N_11888);
nor U12676 (N_12676,N_9760,N_11986);
or U12677 (N_12677,N_9035,N_11183);
nor U12678 (N_12678,N_10031,N_11785);
nand U12679 (N_12679,N_11148,N_11380);
or U12680 (N_12680,N_9763,N_9905);
nor U12681 (N_12681,N_9624,N_11268);
nor U12682 (N_12682,N_9435,N_11846);
nand U12683 (N_12683,N_10327,N_11214);
or U12684 (N_12684,N_9412,N_10465);
and U12685 (N_12685,N_9558,N_9965);
nand U12686 (N_12686,N_10007,N_11422);
nor U12687 (N_12687,N_10719,N_11301);
or U12688 (N_12688,N_10231,N_11132);
and U12689 (N_12689,N_11922,N_11269);
nand U12690 (N_12690,N_9488,N_11745);
nand U12691 (N_12691,N_9659,N_11411);
nand U12692 (N_12692,N_9893,N_10247);
nand U12693 (N_12693,N_10352,N_11077);
nand U12694 (N_12694,N_10188,N_11425);
nor U12695 (N_12695,N_9459,N_9960);
or U12696 (N_12696,N_9911,N_11588);
and U12697 (N_12697,N_11215,N_10393);
nand U12698 (N_12698,N_9933,N_11282);
or U12699 (N_12699,N_10435,N_9139);
nand U12700 (N_12700,N_9284,N_10797);
and U12701 (N_12701,N_10657,N_11585);
nor U12702 (N_12702,N_10140,N_9862);
or U12703 (N_12703,N_9713,N_11392);
and U12704 (N_12704,N_11466,N_10852);
nand U12705 (N_12705,N_9157,N_10145);
or U12706 (N_12706,N_11576,N_10689);
or U12707 (N_12707,N_9425,N_10148);
nand U12708 (N_12708,N_9881,N_9241);
or U12709 (N_12709,N_11223,N_11628);
nand U12710 (N_12710,N_10165,N_11089);
or U12711 (N_12711,N_10136,N_10313);
or U12712 (N_12712,N_10858,N_10429);
or U12713 (N_12713,N_11990,N_10958);
nor U12714 (N_12714,N_10214,N_9199);
or U12715 (N_12715,N_10785,N_10439);
and U12716 (N_12716,N_10009,N_9118);
and U12717 (N_12717,N_11723,N_10710);
nand U12718 (N_12718,N_11688,N_10320);
nor U12719 (N_12719,N_11799,N_10976);
xor U12720 (N_12720,N_10385,N_11864);
and U12721 (N_12721,N_11276,N_11142);
and U12722 (N_12722,N_10363,N_9433);
nand U12723 (N_12723,N_11469,N_9057);
and U12724 (N_12724,N_10828,N_9945);
nand U12725 (N_12725,N_9310,N_9132);
nand U12726 (N_12726,N_11192,N_10817);
nor U12727 (N_12727,N_10871,N_9103);
or U12728 (N_12728,N_10855,N_11681);
nand U12729 (N_12729,N_9872,N_10702);
and U12730 (N_12730,N_10481,N_9309);
nand U12731 (N_12731,N_10896,N_9050);
nor U12732 (N_12732,N_9900,N_9931);
or U12733 (N_12733,N_10950,N_11696);
or U12734 (N_12734,N_10738,N_10779);
and U12735 (N_12735,N_10737,N_11714);
nand U12736 (N_12736,N_9061,N_9917);
and U12737 (N_12737,N_10050,N_9240);
nor U12738 (N_12738,N_9644,N_9351);
nor U12739 (N_12739,N_11486,N_11308);
nand U12740 (N_12740,N_10039,N_9343);
nand U12741 (N_12741,N_9296,N_11113);
nand U12742 (N_12742,N_11382,N_11356);
nor U12743 (N_12743,N_9673,N_9890);
nand U12744 (N_12744,N_9430,N_9169);
nand U12745 (N_12745,N_11067,N_11088);
nand U12746 (N_12746,N_9571,N_10644);
nand U12747 (N_12747,N_11290,N_11692);
and U12748 (N_12748,N_11295,N_10197);
or U12749 (N_12749,N_10295,N_10202);
nor U12750 (N_12750,N_9924,N_9715);
or U12751 (N_12751,N_10207,N_9324);
or U12752 (N_12752,N_10438,N_11198);
or U12753 (N_12753,N_10879,N_10966);
nand U12754 (N_12754,N_10524,N_11478);
nand U12755 (N_12755,N_10835,N_10461);
nor U12756 (N_12756,N_11632,N_11164);
or U12757 (N_12757,N_10978,N_10032);
or U12758 (N_12758,N_10643,N_9083);
and U12759 (N_12759,N_11644,N_10230);
and U12760 (N_12760,N_11965,N_11186);
and U12761 (N_12761,N_9006,N_11463);
and U12762 (N_12762,N_11377,N_10099);
nand U12763 (N_12763,N_11329,N_11610);
and U12764 (N_12764,N_9669,N_10237);
nor U12765 (N_12765,N_9495,N_9104);
and U12766 (N_12766,N_9200,N_11305);
nand U12767 (N_12767,N_10681,N_9611);
or U12768 (N_12768,N_10911,N_11143);
nand U12769 (N_12769,N_11934,N_11573);
nand U12770 (N_12770,N_10486,N_11946);
or U12771 (N_12771,N_10125,N_10995);
or U12772 (N_12772,N_10867,N_10250);
and U12773 (N_12773,N_9171,N_10418);
or U12774 (N_12774,N_9179,N_11954);
and U12775 (N_12775,N_10331,N_11766);
or U12776 (N_12776,N_9952,N_11340);
nand U12777 (N_12777,N_9112,N_10597);
nor U12778 (N_12778,N_10718,N_9315);
nand U12779 (N_12779,N_11225,N_10454);
nor U12780 (N_12780,N_10178,N_9060);
nand U12781 (N_12781,N_10944,N_9888);
and U12782 (N_12782,N_11365,N_10876);
and U12783 (N_12783,N_9012,N_11496);
nand U12784 (N_12784,N_11366,N_9418);
nand U12785 (N_12785,N_11097,N_11788);
nor U12786 (N_12786,N_9706,N_10602);
and U12787 (N_12787,N_10107,N_9963);
nor U12788 (N_12788,N_11806,N_11567);
and U12789 (N_12789,N_11090,N_10473);
or U12790 (N_12790,N_10106,N_10236);
or U12791 (N_12791,N_10134,N_10945);
and U12792 (N_12792,N_11862,N_10836);
or U12793 (N_12793,N_11033,N_10386);
nor U12794 (N_12794,N_10260,N_11442);
nand U12795 (N_12795,N_9091,N_9266);
and U12796 (N_12796,N_11618,N_10278);
nand U12797 (N_12797,N_10219,N_9676);
nor U12798 (N_12798,N_10516,N_9294);
nor U12799 (N_12799,N_11086,N_10449);
or U12800 (N_12800,N_11075,N_9844);
and U12801 (N_12801,N_10816,N_10673);
nor U12802 (N_12802,N_11953,N_9705);
nor U12803 (N_12803,N_11334,N_11700);
nor U12804 (N_12804,N_9852,N_11009);
nand U12805 (N_12805,N_10811,N_9961);
nand U12806 (N_12806,N_9617,N_10694);
or U12807 (N_12807,N_11987,N_11488);
or U12808 (N_12808,N_11384,N_9894);
nor U12809 (N_12809,N_11908,N_9613);
nand U12810 (N_12810,N_9129,N_11630);
nand U12811 (N_12811,N_11072,N_9670);
nor U12812 (N_12812,N_9076,N_11296);
or U12813 (N_12813,N_10475,N_9992);
or U12814 (N_12814,N_10928,N_10721);
nor U12815 (N_12815,N_9451,N_10351);
nand U12816 (N_12816,N_11302,N_10205);
nand U12817 (N_12817,N_10088,N_11473);
or U12818 (N_12818,N_10986,N_11569);
nand U12819 (N_12819,N_11598,N_10273);
nor U12820 (N_12820,N_10934,N_10195);
nand U12821 (N_12821,N_9502,N_10905);
nand U12822 (N_12822,N_10447,N_11173);
or U12823 (N_12823,N_11611,N_9749);
nand U12824 (N_12824,N_9331,N_9956);
nand U12825 (N_12825,N_10650,N_11190);
or U12826 (N_12826,N_9823,N_10396);
and U12827 (N_12827,N_10837,N_9464);
and U12828 (N_12828,N_11733,N_9811);
nand U12829 (N_12829,N_10467,N_9731);
nor U12830 (N_12830,N_10012,N_11434);
or U12831 (N_12831,N_9582,N_9548);
or U12832 (N_12832,N_10371,N_9649);
nand U12833 (N_12833,N_10904,N_9786);
nor U12834 (N_12834,N_9596,N_11974);
nor U12835 (N_12835,N_9637,N_10997);
and U12836 (N_12836,N_10074,N_10072);
nand U12837 (N_12837,N_9591,N_10176);
and U12838 (N_12838,N_10899,N_10960);
and U12839 (N_12839,N_10242,N_11787);
nand U12840 (N_12840,N_9352,N_9102);
and U12841 (N_12841,N_9776,N_10764);
and U12842 (N_12842,N_10906,N_11265);
or U12843 (N_12843,N_11416,N_10456);
and U12844 (N_12844,N_9751,N_11229);
and U12845 (N_12845,N_11136,N_9588);
nor U12846 (N_12846,N_11350,N_9523);
or U12847 (N_12847,N_10932,N_11999);
and U12848 (N_12848,N_9709,N_10128);
and U12849 (N_12849,N_11080,N_9615);
and U12850 (N_12850,N_9720,N_11085);
nand U12851 (N_12851,N_9778,N_10354);
nand U12852 (N_12852,N_10804,N_9080);
or U12853 (N_12853,N_10547,N_10240);
and U12854 (N_12854,N_10652,N_9177);
and U12855 (N_12855,N_11948,N_11412);
nand U12856 (N_12856,N_10532,N_9919);
and U12857 (N_12857,N_11860,N_11179);
nor U12858 (N_12858,N_10424,N_9838);
nand U12859 (N_12859,N_9239,N_11436);
nor U12860 (N_12860,N_11725,N_11976);
and U12861 (N_12861,N_11914,N_11212);
xor U12862 (N_12862,N_11385,N_11858);
nand U12863 (N_12863,N_11550,N_9405);
nand U12864 (N_12864,N_9437,N_10910);
and U12865 (N_12865,N_10114,N_11991);
and U12866 (N_12866,N_9922,N_10255);
and U12867 (N_12867,N_9290,N_11973);
and U12868 (N_12868,N_9301,N_9084);
or U12869 (N_12869,N_10792,N_10463);
nor U12870 (N_12870,N_11147,N_11447);
or U12871 (N_12871,N_10897,N_9573);
nand U12872 (N_12872,N_9230,N_10783);
or U12873 (N_12873,N_11815,N_11394);
and U12874 (N_12874,N_11684,N_10496);
nor U12875 (N_12875,N_9149,N_10036);
or U12876 (N_12876,N_10360,N_10168);
nand U12877 (N_12877,N_11137,N_10466);
or U12878 (N_12878,N_10824,N_10909);
or U12879 (N_12879,N_9789,N_11003);
nand U12880 (N_12880,N_9311,N_11448);
or U12881 (N_12881,N_11789,N_9668);
or U12882 (N_12882,N_11021,N_10679);
and U12883 (N_12883,N_9738,N_9951);
nand U12884 (N_12884,N_10505,N_10223);
nand U12885 (N_12885,N_9788,N_11094);
or U12886 (N_12886,N_9958,N_9413);
nor U12887 (N_12887,N_10605,N_9116);
or U12888 (N_12888,N_11942,N_9567);
nor U12889 (N_12889,N_11204,N_9048);
and U12890 (N_12890,N_10290,N_9825);
nor U12891 (N_12891,N_11339,N_11418);
or U12892 (N_12892,N_11370,N_10399);
or U12893 (N_12893,N_11022,N_10257);
nand U12894 (N_12894,N_9868,N_9291);
and U12895 (N_12895,N_11731,N_9802);
nor U12896 (N_12896,N_9545,N_11271);
nand U12897 (N_12897,N_11962,N_9166);
nand U12898 (N_12898,N_10408,N_10217);
xor U12899 (N_12899,N_10813,N_9927);
and U12900 (N_12900,N_10365,N_11026);
nand U12901 (N_12901,N_9805,N_9001);
or U12902 (N_12902,N_10344,N_10587);
and U12903 (N_12903,N_11835,N_9140);
nor U12904 (N_12904,N_11122,N_11879);
nand U12905 (N_12905,N_10292,N_11568);
and U12906 (N_12906,N_11947,N_9780);
and U12907 (N_12907,N_10947,N_11228);
nor U12908 (N_12908,N_11794,N_9391);
or U12909 (N_12909,N_10314,N_11845);
or U12910 (N_12910,N_10568,N_9288);
nand U12911 (N_12911,N_11128,N_9819);
nand U12912 (N_12912,N_11333,N_9820);
and U12913 (N_12913,N_9685,N_11311);
and U12914 (N_12914,N_9225,N_10619);
or U12915 (N_12915,N_11495,N_10021);
nand U12916 (N_12916,N_11126,N_9798);
or U12917 (N_12917,N_10800,N_11061);
and U12918 (N_12918,N_9081,N_10890);
or U12919 (N_12919,N_10414,N_9563);
and U12920 (N_12920,N_11167,N_9895);
or U12921 (N_12921,N_10596,N_9966);
nand U12922 (N_12922,N_10420,N_10477);
or U12923 (N_12923,N_10228,N_9643);
nand U12924 (N_12924,N_9552,N_10047);
and U12925 (N_12925,N_11847,N_10665);
nor U12926 (N_12926,N_11396,N_11840);
nand U12927 (N_12927,N_9714,N_11050);
nor U12928 (N_12928,N_11602,N_9257);
nand U12929 (N_12929,N_9546,N_11410);
nand U12930 (N_12930,N_11545,N_9357);
and U12931 (N_12931,N_11368,N_10301);
and U12932 (N_12932,N_10600,N_11744);
nor U12933 (N_12933,N_9560,N_9680);
nand U12934 (N_12934,N_10638,N_11648);
and U12935 (N_12935,N_11254,N_10361);
and U12936 (N_12936,N_9843,N_11609);
or U12937 (N_12937,N_9882,N_9511);
nand U12938 (N_12938,N_10533,N_9401);
nor U12939 (N_12939,N_11084,N_11336);
or U12940 (N_12940,N_11701,N_10625);
nand U12941 (N_12941,N_10268,N_11519);
nor U12942 (N_12942,N_9017,N_9901);
and U12943 (N_12943,N_9527,N_10442);
or U12944 (N_12944,N_10181,N_10028);
nor U12945 (N_12945,N_11358,N_11010);
nand U12946 (N_12946,N_11718,N_10969);
nand U12947 (N_12947,N_9229,N_10043);
or U12948 (N_12948,N_11233,N_11462);
and U12949 (N_12949,N_11314,N_9860);
and U12950 (N_12950,N_10740,N_11565);
nor U12951 (N_12951,N_10799,N_9921);
nand U12952 (N_12952,N_10552,N_9042);
and U12953 (N_12953,N_11765,N_11429);
nor U12954 (N_12954,N_9238,N_9897);
nand U12955 (N_12955,N_11540,N_9600);
nor U12956 (N_12956,N_10163,N_9898);
or U12957 (N_12957,N_11433,N_9053);
nor U12958 (N_12958,N_10269,N_11854);
nor U12959 (N_12959,N_11106,N_11016);
nand U12960 (N_12960,N_11578,N_11909);
or U12961 (N_12961,N_10304,N_10283);
nand U12962 (N_12962,N_9775,N_10754);
nand U12963 (N_12963,N_11250,N_9121);
or U12964 (N_12964,N_11674,N_10518);
and U12965 (N_12965,N_9771,N_10913);
and U12966 (N_12966,N_10793,N_9028);
xor U12967 (N_12967,N_9075,N_10448);
or U12968 (N_12968,N_9997,N_9896);
nor U12969 (N_12969,N_9287,N_11866);
and U12970 (N_12970,N_10544,N_9268);
nand U12971 (N_12971,N_11586,N_11306);
and U12972 (N_12972,N_10898,N_10626);
and U12973 (N_12973,N_10922,N_9265);
and U12974 (N_12974,N_10062,N_11020);
nand U12975 (N_12975,N_9707,N_9984);
nand U12976 (N_12976,N_11107,N_9445);
and U12977 (N_12977,N_9740,N_9443);
and U12978 (N_12978,N_11041,N_10616);
nor U12979 (N_12979,N_11703,N_10870);
nand U12980 (N_12980,N_11552,N_11554);
nor U12981 (N_12981,N_10384,N_10359);
nand U12982 (N_12982,N_9605,N_9861);
nand U12983 (N_12983,N_9419,N_11138);
nand U12984 (N_12984,N_9824,N_9161);
nor U12985 (N_12985,N_10234,N_9496);
or U12986 (N_12986,N_11318,N_11872);
nand U12987 (N_12987,N_9416,N_9856);
nand U12988 (N_12988,N_11440,N_10936);
and U12989 (N_12989,N_11742,N_11532);
or U12990 (N_12990,N_10491,N_9536);
nand U12991 (N_12991,N_11971,N_11743);
nand U12992 (N_12992,N_10078,N_10974);
or U12993 (N_12993,N_11544,N_10757);
nand U12994 (N_12994,N_10389,N_10506);
and U12995 (N_12995,N_9056,N_11893);
nor U12996 (N_12996,N_11131,N_11811);
nand U12997 (N_12997,N_11180,N_10798);
or U12998 (N_12998,N_10884,N_11058);
or U12999 (N_12999,N_11117,N_11530);
or U13000 (N_13000,N_11943,N_11419);
and U13001 (N_13001,N_11603,N_11871);
nor U13002 (N_13002,N_9395,N_9068);
or U13003 (N_13003,N_10748,N_10048);
and U13004 (N_13004,N_9192,N_11757);
or U13005 (N_13005,N_11509,N_11673);
nand U13006 (N_13006,N_10720,N_9071);
and U13007 (N_13007,N_10751,N_10001);
nor U13008 (N_13008,N_10956,N_10245);
or U13009 (N_13009,N_11716,N_11898);
and U13010 (N_13010,N_11520,N_10569);
nor U13011 (N_13011,N_9394,N_9438);
nor U13012 (N_13012,N_10937,N_10994);
or U13013 (N_13013,N_9182,N_11939);
nand U13014 (N_13014,N_10615,N_10433);
and U13015 (N_13015,N_10728,N_11619);
and U13016 (N_13016,N_11272,N_10768);
nor U13017 (N_13017,N_10529,N_10815);
or U13018 (N_13018,N_9339,N_11176);
nand U13019 (N_13019,N_10322,N_11389);
nand U13020 (N_13020,N_10122,N_11593);
nand U13021 (N_13021,N_10822,N_10194);
nor U13022 (N_13022,N_9601,N_10309);
and U13023 (N_13023,N_11001,N_11452);
nor U13024 (N_13024,N_9212,N_9318);
nand U13025 (N_13025,N_11485,N_9517);
nand U13026 (N_13026,N_9493,N_11230);
nor U13027 (N_13027,N_9165,N_9745);
nor U13028 (N_13028,N_10131,N_11207);
xor U13029 (N_13029,N_10693,N_11933);
nor U13030 (N_13030,N_10144,N_9105);
and U13031 (N_13031,N_10323,N_10318);
nand U13032 (N_13032,N_11013,N_11388);
nand U13033 (N_13033,N_9447,N_9935);
nand U13034 (N_13034,N_10211,N_10987);
or U13035 (N_13035,N_9134,N_9349);
nand U13036 (N_13036,N_9507,N_10015);
and U13037 (N_13037,N_11527,N_11070);
nand U13038 (N_13038,N_11548,N_9320);
nand U13039 (N_13039,N_9302,N_10286);
nand U13040 (N_13040,N_9453,N_9543);
or U13041 (N_13041,N_11768,N_9701);
nor U13042 (N_13042,N_11294,N_9307);
or U13043 (N_13043,N_10049,N_11591);
nor U13044 (N_13044,N_10018,N_9744);
nor U13045 (N_13045,N_9441,N_11557);
nand U13046 (N_13046,N_11427,N_10977);
or U13047 (N_13047,N_10711,N_9499);
or U13048 (N_13048,N_11612,N_9276);
or U13049 (N_13049,N_10087,N_9504);
nor U13050 (N_13050,N_9732,N_9974);
and U13051 (N_13051,N_10753,N_10715);
and U13052 (N_13052,N_10150,N_10827);
and U13053 (N_13053,N_10787,N_11055);
nand U13054 (N_13054,N_10293,N_11992);
and U13055 (N_13055,N_9583,N_10925);
or U13056 (N_13056,N_10450,N_11729);
and U13057 (N_13057,N_9808,N_9337);
nor U13058 (N_13058,N_10869,N_9454);
nor U13059 (N_13059,N_10282,N_11615);
and U13060 (N_13060,N_10921,N_11019);
and U13061 (N_13061,N_10321,N_10935);
nand U13062 (N_13062,N_10550,N_10946);
nor U13063 (N_13063,N_9902,N_9703);
nand U13064 (N_13064,N_10502,N_10818);
and U13065 (N_13065,N_11949,N_9551);
nor U13066 (N_13066,N_11163,N_11479);
and U13067 (N_13067,N_11188,N_11501);
nand U13068 (N_13068,N_10225,N_10109);
or U13069 (N_13069,N_9093,N_11116);
nor U13070 (N_13070,N_10649,N_10149);
and U13071 (N_13071,N_11738,N_10961);
nor U13072 (N_13072,N_9065,N_9787);
xor U13073 (N_13073,N_9436,N_9156);
or U13074 (N_13074,N_9959,N_10688);
nand U13075 (N_13075,N_9779,N_10993);
and U13076 (N_13076,N_9985,N_10826);
nor U13077 (N_13077,N_11570,N_10914);
nor U13078 (N_13078,N_9082,N_10854);
or U13079 (N_13079,N_9781,N_11727);
and U13080 (N_13080,N_9926,N_10367);
nand U13081 (N_13081,N_11607,N_10490);
nand U13082 (N_13082,N_11514,N_11538);
nand U13083 (N_13083,N_11918,N_11825);
nor U13084 (N_13084,N_11746,N_10758);
and U13085 (N_13085,N_11852,N_11857);
nand U13086 (N_13086,N_9070,N_9627);
and U13087 (N_13087,N_11950,N_11779);
nand U13088 (N_13088,N_11326,N_11078);
and U13089 (N_13089,N_11726,N_10156);
or U13090 (N_13090,N_11769,N_11476);
or U13091 (N_13091,N_9452,N_11482);
or U13092 (N_13092,N_10676,N_9253);
nand U13093 (N_13093,N_9869,N_10388);
or U13094 (N_13094,N_10279,N_9652);
or U13095 (N_13095,N_10949,N_11653);
and U13096 (N_13096,N_9000,N_9135);
or U13097 (N_13097,N_10873,N_9585);
and U13098 (N_13098,N_9072,N_9936);
and U13099 (N_13099,N_10443,N_9364);
and U13100 (N_13100,N_9286,N_9227);
nand U13101 (N_13101,N_9699,N_10713);
or U13102 (N_13102,N_10708,N_9007);
nand U13103 (N_13103,N_9671,N_9323);
nor U13104 (N_13104,N_10489,N_11614);
or U13105 (N_13105,N_10684,N_10025);
nor U13106 (N_13106,N_9233,N_9079);
nor U13107 (N_13107,N_11952,N_10493);
nand U13108 (N_13108,N_10315,N_11896);
nor U13109 (N_13109,N_11328,N_11770);
and U13110 (N_13110,N_10519,N_10732);
and U13111 (N_13111,N_10310,N_10680);
or U13112 (N_13112,N_10402,N_11355);
nand U13113 (N_13113,N_10452,N_9753);
and U13114 (N_13114,N_9064,N_11353);
and U13115 (N_13115,N_9521,N_10772);
and U13116 (N_13116,N_9194,N_11777);
and U13117 (N_13117,N_11697,N_11399);
nor U13118 (N_13118,N_9724,N_10133);
and U13119 (N_13119,N_9100,N_10555);
or U13120 (N_13120,N_10362,N_9248);
and U13121 (N_13121,N_10917,N_11242);
nor U13122 (N_13122,N_9058,N_11511);
and U13123 (N_13123,N_11796,N_11487);
or U13124 (N_13124,N_10539,N_9783);
or U13125 (N_13125,N_11209,N_10326);
nand U13126 (N_13126,N_10166,N_11468);
and U13127 (N_13127,N_10186,N_11623);
nand U13128 (N_13128,N_11059,N_9059);
nand U13129 (N_13129,N_10332,N_10382);
and U13130 (N_13130,N_11391,N_11719);
nor U13131 (N_13131,N_11110,N_10376);
nor U13132 (N_13132,N_10661,N_9275);
nand U13133 (N_13133,N_9815,N_10776);
nor U13134 (N_13134,N_11786,N_10244);
or U13135 (N_13135,N_10215,N_10324);
or U13136 (N_13136,N_10640,N_10762);
or U13137 (N_13137,N_11824,N_10553);
nor U13138 (N_13138,N_11159,N_10622);
or U13139 (N_13139,N_10682,N_10220);
nor U13140 (N_13140,N_11821,N_11453);
nor U13141 (N_13141,N_10608,N_11406);
and U13142 (N_13142,N_11828,N_10369);
and U13143 (N_13143,N_10035,N_11206);
nand U13144 (N_13144,N_9566,N_11335);
nor U13145 (N_13145,N_10462,N_11784);
nor U13146 (N_13146,N_10305,N_9015);
nor U13147 (N_13147,N_9365,N_11439);
nand U13148 (N_13148,N_11507,N_11177);
and U13149 (N_13149,N_11330,N_11100);
or U13150 (N_13150,N_10686,N_10656);
or U13151 (N_13151,N_11052,N_9408);
nand U13152 (N_13152,N_10142,N_10272);
and U13153 (N_13153,N_10154,N_11408);
nor U13154 (N_13154,N_9095,N_9503);
or U13155 (N_13155,N_10177,N_9784);
nand U13156 (N_13156,N_10127,N_11601);
nor U13157 (N_13157,N_9925,N_10404);
nand U13158 (N_13158,N_9466,N_10948);
nand U13159 (N_13159,N_11709,N_11708);
or U13160 (N_13160,N_10883,N_11979);
nand U13161 (N_13161,N_9086,N_11403);
nand U13162 (N_13162,N_9415,N_11936);
nand U13163 (N_13163,N_10705,N_11894);
nand U13164 (N_13164,N_11195,N_11989);
nand U13165 (N_13165,N_10016,N_9866);
nand U13166 (N_13166,N_9237,N_11740);
and U13167 (N_13167,N_9245,N_10841);
and U13168 (N_13168,N_11025,N_10786);
nor U13169 (N_13169,N_9236,N_11104);
and U13170 (N_13170,N_10022,N_11524);
nor U13171 (N_13171,N_10151,N_11387);
nand U13172 (N_13172,N_11430,N_10276);
or U13173 (N_13173,N_10637,N_11317);
nand U13174 (N_13174,N_11451,N_9209);
nor U13175 (N_13175,N_11842,N_9880);
and U13176 (N_13176,N_10912,N_9317);
nand U13177 (N_13177,N_9832,N_10618);
nand U13178 (N_13178,N_11850,N_9032);
nand U13179 (N_13179,N_10559,N_10330);
nor U13180 (N_13180,N_11758,N_11407);
or U13181 (N_13181,N_10736,N_10445);
nor U13182 (N_13182,N_11631,N_9516);
and U13183 (N_13183,N_9152,N_11669);
and U13184 (N_13184,N_9993,N_10535);
or U13185 (N_13185,N_11043,N_9841);
nor U13186 (N_13186,N_11493,N_9554);
and U13187 (N_13187,N_11181,N_11546);
nand U13188 (N_13188,N_11082,N_10333);
nand U13189 (N_13189,N_11826,N_11279);
nor U13190 (N_13190,N_11721,N_9733);
and U13191 (N_13191,N_10038,N_9821);
nor U13192 (N_13192,N_11895,N_11803);
xor U13193 (N_13193,N_10277,N_9422);
nand U13194 (N_13194,N_9619,N_10316);
or U13195 (N_13195,N_10703,N_10943);
nand U13196 (N_13196,N_9191,N_11249);
nand U13197 (N_13197,N_9949,N_9969);
and U13198 (N_13198,N_9870,N_11484);
and U13199 (N_13199,N_10825,N_10510);
nor U13200 (N_13200,N_10933,N_10058);
nand U13201 (N_13201,N_9608,N_11141);
nor U13202 (N_13202,N_10951,N_9849);
or U13203 (N_13203,N_10391,N_11156);
nand U13204 (N_13204,N_9005,N_10375);
and U13205 (N_13205,N_9682,N_11367);
or U13206 (N_13206,N_11369,N_11320);
or U13207 (N_13207,N_9231,N_10162);
and U13208 (N_13208,N_9864,N_9650);
and U13209 (N_13209,N_10319,N_9448);
nand U13210 (N_13210,N_9679,N_11376);
and U13211 (N_13211,N_11413,N_9645);
nand U13212 (N_13212,N_9672,N_11885);
or U13213 (N_13213,N_11409,N_10624);
nand U13214 (N_13214,N_10985,N_10548);
nand U13215 (N_13215,N_9795,N_10298);
nor U13216 (N_13216,N_10970,N_9846);
nand U13217 (N_13217,N_11170,N_9625);
nand U13218 (N_13218,N_11877,N_11558);
or U13219 (N_13219,N_9579,N_10497);
or U13220 (N_13220,N_11491,N_10441);
nor U13221 (N_13221,N_9577,N_11613);
nor U13222 (N_13222,N_9675,N_11608);
or U13223 (N_13223,N_11996,N_9941);
or U13224 (N_13224,N_9046,N_11438);
nand U13225 (N_13225,N_9794,N_9283);
or U13226 (N_13226,N_10090,N_9110);
nand U13227 (N_13227,N_9737,N_10872);
nor U13228 (N_13228,N_10081,N_10729);
and U13229 (N_13229,N_9692,N_9505);
nor U13230 (N_13230,N_9386,N_10610);
nand U13231 (N_13231,N_11039,N_9663);
and U13232 (N_13232,N_9531,N_9460);
and U13233 (N_13233,N_10620,N_11374);
nor U13234 (N_13234,N_11202,N_10472);
nand U13235 (N_13235,N_10667,N_10885);
nand U13236 (N_13236,N_9155,N_11470);
nand U13237 (N_13237,N_10586,N_9450);
or U13238 (N_13238,N_11034,N_10082);
nand U13239 (N_13239,N_10810,N_11884);
and U13240 (N_13240,N_10206,N_11220);
nor U13241 (N_13241,N_10840,N_9378);
and U13242 (N_13242,N_11200,N_9884);
nor U13243 (N_13243,N_10838,N_10037);
nand U13244 (N_13244,N_11776,N_11535);
and U13245 (N_13245,N_11679,N_9387);
and U13246 (N_13246,N_11998,N_11221);
nand U13247 (N_13247,N_11916,N_9279);
nand U13248 (N_13248,N_10096,N_9677);
nor U13249 (N_13249,N_9797,N_10726);
and U13250 (N_13250,N_9818,N_11289);
and U13251 (N_13251,N_10051,N_10383);
or U13252 (N_13252,N_10517,N_9382);
or U13253 (N_13253,N_10894,N_11659);
nand U13254 (N_13254,N_11477,N_11624);
nor U13255 (N_13255,N_11191,N_10381);
nor U13256 (N_13256,N_9518,N_11805);
or U13257 (N_13257,N_11596,N_10723);
and U13258 (N_13258,N_11533,N_9903);
and U13259 (N_13259,N_11634,N_10598);
and U13260 (N_13260,N_10692,N_10992);
or U13261 (N_13261,N_9346,N_11771);
or U13262 (N_13262,N_10655,N_9098);
and U13263 (N_13263,N_11981,N_10707);
and U13264 (N_13264,N_10115,N_10812);
xor U13265 (N_13265,N_11508,N_9008);
and U13266 (N_13266,N_9696,N_10239);
nand U13267 (N_13267,N_11739,N_11465);
and U13268 (N_13268,N_11124,N_11869);
or U13269 (N_13269,N_10345,N_11008);
and U13270 (N_13270,N_9817,N_11819);
nor U13271 (N_13271,N_11312,N_9913);
nand U13272 (N_13272,N_10302,N_9113);
nand U13273 (N_13273,N_10474,N_10942);
and U13274 (N_13274,N_11112,N_10601);
and U13275 (N_13275,N_11836,N_11668);
nor U13276 (N_13276,N_9597,N_11157);
and U13277 (N_13277,N_11068,N_11054);
nor U13278 (N_13278,N_10678,N_10755);
or U13279 (N_13279,N_9553,N_9796);
nand U13280 (N_13280,N_9025,N_11103);
nand U13281 (N_13281,N_11640,N_9792);
nor U13282 (N_13282,N_10926,N_11284);
or U13283 (N_13283,N_11827,N_10546);
or U13284 (N_13284,N_10965,N_9912);
nand U13285 (N_13285,N_9610,N_11800);
nor U13286 (N_13286,N_10263,N_11045);
nor U13287 (N_13287,N_11327,N_9338);
and U13288 (N_13288,N_11120,N_9036);
or U13289 (N_13289,N_10253,N_10562);
nand U13290 (N_13290,N_11874,N_10570);
nand U13291 (N_13291,N_9855,N_11553);
xnor U13292 (N_13292,N_9804,N_10190);
nor U13293 (N_13293,N_9800,N_9586);
nand U13294 (N_13294,N_9828,N_9562);
or U13295 (N_13295,N_9027,N_10918);
nor U13296 (N_13296,N_10829,N_10634);
nor U13297 (N_13297,N_9630,N_11278);
nand U13298 (N_13298,N_9463,N_9232);
xnor U13299 (N_13299,N_11594,N_11492);
and U13300 (N_13300,N_9826,N_10991);
and U13301 (N_13301,N_9557,N_9054);
nand U13302 (N_13302,N_11580,N_10426);
nor U13303 (N_13303,N_11963,N_10373);
nor U13304 (N_13304,N_9989,N_9981);
and U13305 (N_13305,N_10865,N_11652);
or U13306 (N_13306,N_11303,N_9635);
nand U13307 (N_13307,N_9362,N_10940);
nor U13308 (N_13308,N_11160,N_9456);
nor U13309 (N_13309,N_11280,N_11761);
nor U13310 (N_13310,N_9814,N_11556);
nand U13311 (N_13311,N_11166,N_10549);
or U13312 (N_13312,N_11956,N_11152);
and U13313 (N_13313,N_10971,N_10355);
or U13314 (N_13314,N_11625,N_9834);
or U13315 (N_13315,N_10739,N_11997);
nand U13316 (N_13316,N_9618,N_11667);
or U13317 (N_13317,N_9280,N_11891);
nor U13318 (N_13318,N_10173,N_10630);
or U13319 (N_13319,N_9356,N_11865);
nand U13320 (N_13320,N_11235,N_10222);
nor U13321 (N_13321,N_9689,N_10185);
nor U13322 (N_13322,N_9883,N_11635);
and U13323 (N_13323,N_9806,N_10642);
nand U13324 (N_13324,N_11984,N_10695);
and U13325 (N_13325,N_10085,N_10364);
and U13326 (N_13326,N_11454,N_10097);
and U13327 (N_13327,N_9930,N_9322);
and U13328 (N_13328,N_10774,N_9402);
nor U13329 (N_13329,N_10717,N_9168);
nand U13330 (N_13330,N_10583,N_10262);
or U13331 (N_13331,N_11481,N_11227);
nand U13332 (N_13332,N_10416,N_11797);
nor U13333 (N_13333,N_11642,N_11270);
or U13334 (N_13334,N_11873,N_11130);
and U13335 (N_13335,N_9587,N_10203);
nor U13336 (N_13336,N_9561,N_11575);
or U13337 (N_13337,N_9761,N_10631);
and U13338 (N_13338,N_9829,N_10795);
and U13339 (N_13339,N_10494,N_11687);
or U13340 (N_13340,N_9396,N_10041);
nand U13341 (N_13341,N_10248,N_11345);
and U13342 (N_13342,N_11809,N_11747);
or U13343 (N_13343,N_9242,N_11650);
nand U13344 (N_13344,N_9876,N_9661);
nor U13345 (N_13345,N_11446,N_11390);
or U13346 (N_13346,N_10639,N_11867);
nand U13347 (N_13347,N_11627,N_11959);
xnor U13348 (N_13348,N_10086,N_9739);
nor U13349 (N_13349,N_10182,N_11649);
xor U13350 (N_13350,N_10053,N_9314);
xor U13351 (N_13351,N_10613,N_9891);
nand U13352 (N_13352,N_9678,N_10328);
nor U13353 (N_13353,N_11808,N_11386);
and U13354 (N_13354,N_11145,N_9688);
or U13355 (N_13355,N_11980,N_10526);
nor U13356 (N_13356,N_9774,N_10174);
nand U13357 (N_13357,N_11031,N_9593);
and U13358 (N_13358,N_11698,N_11158);
or U13359 (N_13359,N_11671,N_9885);
nor U13360 (N_13360,N_10334,N_9404);
or U13361 (N_13361,N_9598,N_9162);
or U13362 (N_13362,N_11571,N_10580);
and U13363 (N_13363,N_11029,N_11030);
nand U13364 (N_13364,N_11261,N_11095);
and U13365 (N_13365,N_11099,N_9142);
or U13366 (N_13366,N_10975,N_9947);
and U13367 (N_13367,N_10057,N_11555);
nor U13368 (N_13368,N_11315,N_10528);
nor U13369 (N_13369,N_9125,N_10436);
nand U13370 (N_13370,N_9254,N_9667);
or U13371 (N_13371,N_10503,N_11604);
or U13372 (N_13372,N_11756,N_9483);
and U13373 (N_13373,N_10536,N_9887);
or U13374 (N_13374,N_9224,N_11780);
or U13375 (N_13375,N_10627,N_11849);
and U13376 (N_13376,N_10589,N_11702);
nor U13377 (N_13377,N_9790,N_10476);
and U13378 (N_13378,N_9400,N_9475);
and U13379 (N_13379,N_10011,N_9909);
nor U13380 (N_13380,N_10218,N_10213);
or U13381 (N_13381,N_11359,N_9683);
nor U13382 (N_13382,N_9736,N_9099);
nor U13383 (N_13383,N_9446,N_9258);
nor U13384 (N_13384,N_9384,N_9646);
and U13385 (N_13385,N_11542,N_11938);
nand U13386 (N_13386,N_11883,N_10699);
and U13387 (N_13387,N_9875,N_10303);
nor U13388 (N_13388,N_9184,N_9727);
nor U13389 (N_13389,N_9642,N_11651);
nand U13390 (N_13390,N_11562,N_10104);
or U13391 (N_13391,N_10229,N_10782);
or U13392 (N_13392,N_9077,N_11349);
and U13393 (N_13393,N_11000,N_11792);
nand U13394 (N_13394,N_11906,N_9469);
nor U13395 (N_13395,N_10814,N_10540);
nand U13396 (N_13396,N_9421,N_10501);
nor U13397 (N_13397,N_10340,N_11017);
nand U13398 (N_13398,N_9509,N_9809);
nand U13399 (N_13399,N_11887,N_10915);
nand U13400 (N_13400,N_11724,N_11577);
nand U13401 (N_13401,N_9906,N_10138);
or U13402 (N_13402,N_9839,N_11600);
and U13403 (N_13403,N_11371,N_11782);
and U13404 (N_13404,N_9544,N_11474);
xor U13405 (N_13405,N_10508,N_10171);
or U13406 (N_13406,N_11247,N_10629);
or U13407 (N_13407,N_11251,N_9980);
nand U13408 (N_13408,N_9153,N_9633);
nor U13409 (N_13409,N_10698,N_10670);
or U13410 (N_13410,N_9967,N_11196);
and U13411 (N_13411,N_11641,N_11801);
nand U13412 (N_13412,N_11977,N_10289);
or U13413 (N_13413,N_9565,N_10013);
or U13414 (N_13414,N_11691,N_11431);
and U13415 (N_13415,N_9612,N_10716);
nor U13416 (N_13416,N_11244,N_10780);
and U13417 (N_13417,N_11304,N_10275);
and U13418 (N_13418,N_11735,N_11379);
and U13419 (N_13419,N_11266,N_11500);
or U13420 (N_13420,N_11240,N_9147);
nand U13421 (N_13421,N_10372,N_10697);
nor U13422 (N_13422,N_10499,N_11199);
nand U13423 (N_13423,N_9664,N_11150);
or U13424 (N_13424,N_11699,N_11224);
nand U13425 (N_13425,N_11450,N_11060);
nand U13426 (N_13426,N_9877,N_10901);
nand U13427 (N_13427,N_10370,N_10557);
or U13428 (N_13428,N_11264,N_9173);
nand U13429 (N_13429,N_11114,N_9754);
nand U13430 (N_13430,N_9595,N_9572);
nor U13431 (N_13431,N_11397,N_11903);
or U13432 (N_13432,N_11119,N_11313);
and U13433 (N_13433,N_9449,N_9078);
and U13434 (N_13434,N_10403,N_11169);
nand U13435 (N_13435,N_9858,N_9607);
nor U13436 (N_13436,N_11316,N_10061);
nor U13437 (N_13437,N_9982,N_10887);
nand U13438 (N_13438,N_11182,N_10542);
and U13439 (N_13439,N_10159,N_9023);
nand U13440 (N_13440,N_10431,N_11044);
nand U13441 (N_13441,N_10259,N_10691);
nor U13442 (N_13442,N_11323,N_9986);
and U13443 (N_13443,N_10000,N_10538);
nor U13444 (N_13444,N_10019,N_9090);
nor U13445 (N_13445,N_10875,N_9335);
nor U13446 (N_13446,N_11083,N_10395);
or U13447 (N_13447,N_10413,N_11375);
nor U13448 (N_13448,N_11958,N_11528);
and U13449 (N_13449,N_9530,N_10432);
nand U13450 (N_13450,N_9066,N_9793);
nand U13451 (N_13451,N_10341,N_10850);
or U13452 (N_13452,N_9040,N_11475);
and U13453 (N_13453,N_10939,N_9431);
nor U13454 (N_13454,N_11331,N_9300);
nor U13455 (N_13455,N_10092,N_11748);
nand U13456 (N_13456,N_9136,N_9979);
nor U13457 (N_13457,N_9791,N_9484);
nor U13458 (N_13458,N_9748,N_9863);
or U13459 (N_13459,N_10521,N_9494);
nor U13460 (N_13460,N_9151,N_9497);
and U13461 (N_13461,N_9534,N_10094);
or U13462 (N_13462,N_10069,N_11920);
nand U13463 (N_13463,N_10487,N_10888);
and U13464 (N_13464,N_11966,N_9247);
nor U13465 (N_13465,N_11695,N_9202);
nand U13466 (N_13466,N_11014,N_9687);
and U13467 (N_13467,N_9638,N_10346);
nand U13468 (N_13468,N_9115,N_11064);
nand U13469 (N_13469,N_11876,N_10766);
and U13470 (N_13470,N_10120,N_10054);
nand U13471 (N_13471,N_9411,N_11178);
nor U13472 (N_13472,N_9594,N_9034);
and U13473 (N_13473,N_11444,N_10175);
and U13474 (N_13474,N_9358,N_11497);
xnor U13475 (N_13475,N_10183,N_9181);
nand U13476 (N_13476,N_11924,N_11194);
and U13477 (N_13477,N_9108,N_10606);
nor U13478 (N_13478,N_9297,N_10187);
and U13479 (N_13479,N_9178,N_10929);
nand U13480 (N_13480,N_10633,N_10060);
and U13481 (N_13481,N_10147,N_10989);
nor U13482 (N_13482,N_11921,N_10572);
or U13483 (N_13483,N_9747,N_9062);
nand U13484 (N_13484,N_11133,N_10743);
nand U13485 (N_13485,N_9468,N_10842);
or U13486 (N_13486,N_10848,N_10575);
or U13487 (N_13487,N_11432,N_11678);
nand U13488 (N_13488,N_11111,N_10135);
xnor U13489 (N_13489,N_10584,N_11259);
nand U13490 (N_13490,N_10067,N_11420);
and U13491 (N_13491,N_9145,N_10599);
or U13492 (N_13492,N_11246,N_9052);
nand U13493 (N_13493,N_10406,N_10952);
and U13494 (N_13494,N_10091,N_11838);
nand U13495 (N_13495,N_11677,N_10297);
or U13496 (N_13496,N_9409,N_11139);
nor U13497 (N_13497,N_9355,N_10509);
and U13498 (N_13498,N_10805,N_9907);
nor U13499 (N_13499,N_10790,N_11767);
nand U13500 (N_13500,N_9985,N_11819);
nor U13501 (N_13501,N_9972,N_11212);
and U13502 (N_13502,N_11142,N_11392);
nor U13503 (N_13503,N_11683,N_10574);
or U13504 (N_13504,N_11839,N_9672);
nor U13505 (N_13505,N_11238,N_11923);
and U13506 (N_13506,N_10679,N_11122);
and U13507 (N_13507,N_10390,N_11767);
nor U13508 (N_13508,N_10475,N_9337);
or U13509 (N_13509,N_9862,N_9380);
nand U13510 (N_13510,N_9242,N_11425);
or U13511 (N_13511,N_10236,N_10145);
nor U13512 (N_13512,N_11224,N_9067);
and U13513 (N_13513,N_9077,N_11813);
and U13514 (N_13514,N_11042,N_11770);
nand U13515 (N_13515,N_10541,N_10384);
nand U13516 (N_13516,N_10055,N_11736);
and U13517 (N_13517,N_10893,N_10973);
nor U13518 (N_13518,N_9742,N_10850);
or U13519 (N_13519,N_11132,N_11926);
or U13520 (N_13520,N_10064,N_11667);
nand U13521 (N_13521,N_11737,N_11082);
and U13522 (N_13522,N_10515,N_10848);
nor U13523 (N_13523,N_9372,N_11818);
nor U13524 (N_13524,N_11033,N_10474);
nand U13525 (N_13525,N_10971,N_9233);
nand U13526 (N_13526,N_9401,N_9661);
and U13527 (N_13527,N_9720,N_9701);
and U13528 (N_13528,N_11792,N_11739);
or U13529 (N_13529,N_11654,N_11944);
or U13530 (N_13530,N_11529,N_11556);
nand U13531 (N_13531,N_11466,N_11373);
nand U13532 (N_13532,N_11964,N_11782);
nand U13533 (N_13533,N_10360,N_11856);
and U13534 (N_13534,N_9193,N_9969);
xor U13535 (N_13535,N_9271,N_11337);
or U13536 (N_13536,N_10578,N_11138);
and U13537 (N_13537,N_11789,N_10750);
and U13538 (N_13538,N_10256,N_10168);
nand U13539 (N_13539,N_9364,N_11291);
and U13540 (N_13540,N_9307,N_10843);
nor U13541 (N_13541,N_10563,N_10931);
nor U13542 (N_13542,N_9195,N_11365);
nor U13543 (N_13543,N_9145,N_10045);
nand U13544 (N_13544,N_10116,N_9373);
nor U13545 (N_13545,N_10111,N_11902);
nand U13546 (N_13546,N_9530,N_10428);
or U13547 (N_13547,N_10514,N_10291);
and U13548 (N_13548,N_9994,N_10641);
and U13549 (N_13549,N_9158,N_10208);
nand U13550 (N_13550,N_10604,N_11312);
or U13551 (N_13551,N_11226,N_11933);
or U13552 (N_13552,N_9441,N_11830);
or U13553 (N_13553,N_9656,N_10829);
and U13554 (N_13554,N_10513,N_9818);
nor U13555 (N_13555,N_10887,N_10205);
and U13556 (N_13556,N_11439,N_11119);
nor U13557 (N_13557,N_11033,N_11661);
or U13558 (N_13558,N_11436,N_11136);
and U13559 (N_13559,N_11556,N_10984);
nor U13560 (N_13560,N_9735,N_10423);
and U13561 (N_13561,N_11410,N_11328);
nor U13562 (N_13562,N_9292,N_9759);
or U13563 (N_13563,N_11013,N_11103);
and U13564 (N_13564,N_9877,N_10720);
and U13565 (N_13565,N_11419,N_11066);
nor U13566 (N_13566,N_11676,N_10437);
nand U13567 (N_13567,N_9938,N_10393);
nand U13568 (N_13568,N_11964,N_10619);
or U13569 (N_13569,N_10867,N_9847);
nor U13570 (N_13570,N_9906,N_9068);
nand U13571 (N_13571,N_11590,N_10856);
or U13572 (N_13572,N_11119,N_10644);
nor U13573 (N_13573,N_11437,N_9544);
and U13574 (N_13574,N_10588,N_11695);
nand U13575 (N_13575,N_11533,N_11528);
or U13576 (N_13576,N_9096,N_9192);
nor U13577 (N_13577,N_11408,N_10122);
nand U13578 (N_13578,N_9707,N_9036);
nor U13579 (N_13579,N_10979,N_10837);
xnor U13580 (N_13580,N_11329,N_9999);
nand U13581 (N_13581,N_11292,N_11906);
xor U13582 (N_13582,N_9201,N_9737);
nand U13583 (N_13583,N_10559,N_11891);
nand U13584 (N_13584,N_10543,N_10587);
and U13585 (N_13585,N_10528,N_11016);
or U13586 (N_13586,N_11077,N_10254);
nand U13587 (N_13587,N_9010,N_9534);
or U13588 (N_13588,N_10977,N_10396);
nand U13589 (N_13589,N_10605,N_10447);
and U13590 (N_13590,N_10051,N_10566);
and U13591 (N_13591,N_11012,N_11588);
and U13592 (N_13592,N_9948,N_9130);
or U13593 (N_13593,N_10032,N_9364);
nor U13594 (N_13594,N_10452,N_10211);
nand U13595 (N_13595,N_9583,N_11262);
or U13596 (N_13596,N_9678,N_11410);
or U13597 (N_13597,N_10482,N_9796);
nand U13598 (N_13598,N_11146,N_9242);
and U13599 (N_13599,N_11609,N_9249);
or U13600 (N_13600,N_11191,N_11467);
and U13601 (N_13601,N_10872,N_9958);
or U13602 (N_13602,N_10515,N_11037);
and U13603 (N_13603,N_10637,N_10896);
nand U13604 (N_13604,N_10693,N_9446);
and U13605 (N_13605,N_9096,N_10485);
nor U13606 (N_13606,N_10905,N_9431);
nor U13607 (N_13607,N_11007,N_11116);
nand U13608 (N_13608,N_9544,N_9748);
nand U13609 (N_13609,N_11705,N_11026);
or U13610 (N_13610,N_10837,N_9888);
nor U13611 (N_13611,N_11892,N_9001);
and U13612 (N_13612,N_9118,N_11396);
nand U13613 (N_13613,N_9909,N_9348);
and U13614 (N_13614,N_10602,N_11321);
nand U13615 (N_13615,N_9183,N_11869);
or U13616 (N_13616,N_9848,N_9229);
or U13617 (N_13617,N_9964,N_11714);
xor U13618 (N_13618,N_9843,N_9529);
or U13619 (N_13619,N_10524,N_11747);
nor U13620 (N_13620,N_11440,N_10348);
or U13621 (N_13621,N_11395,N_11651);
nand U13622 (N_13622,N_10022,N_11573);
or U13623 (N_13623,N_9185,N_9970);
or U13624 (N_13624,N_10646,N_10931);
and U13625 (N_13625,N_9188,N_9535);
and U13626 (N_13626,N_11996,N_10696);
or U13627 (N_13627,N_11654,N_11857);
nor U13628 (N_13628,N_9609,N_10719);
nand U13629 (N_13629,N_9482,N_9905);
and U13630 (N_13630,N_11843,N_9966);
nand U13631 (N_13631,N_10868,N_9747);
and U13632 (N_13632,N_11164,N_11703);
or U13633 (N_13633,N_11176,N_9130);
or U13634 (N_13634,N_10769,N_10958);
nand U13635 (N_13635,N_11841,N_9017);
and U13636 (N_13636,N_10661,N_10925);
or U13637 (N_13637,N_10733,N_11414);
and U13638 (N_13638,N_10542,N_11507);
nor U13639 (N_13639,N_9188,N_11353);
or U13640 (N_13640,N_11148,N_10937);
or U13641 (N_13641,N_11755,N_10910);
or U13642 (N_13642,N_10471,N_10054);
or U13643 (N_13643,N_11223,N_10341);
nand U13644 (N_13644,N_11904,N_9784);
and U13645 (N_13645,N_10448,N_10663);
and U13646 (N_13646,N_10663,N_11796);
and U13647 (N_13647,N_10167,N_10564);
nor U13648 (N_13648,N_10203,N_10470);
nand U13649 (N_13649,N_11908,N_11047);
nand U13650 (N_13650,N_11642,N_10908);
nor U13651 (N_13651,N_10906,N_11152);
and U13652 (N_13652,N_11949,N_11806);
or U13653 (N_13653,N_11206,N_10044);
nor U13654 (N_13654,N_9364,N_10947);
nor U13655 (N_13655,N_11451,N_9968);
nor U13656 (N_13656,N_9362,N_10162);
and U13657 (N_13657,N_10574,N_9506);
xnor U13658 (N_13658,N_9174,N_9804);
nand U13659 (N_13659,N_9443,N_10606);
and U13660 (N_13660,N_9002,N_11431);
nor U13661 (N_13661,N_11372,N_9037);
nor U13662 (N_13662,N_9068,N_9648);
nor U13663 (N_13663,N_11946,N_10034);
nand U13664 (N_13664,N_11636,N_9728);
and U13665 (N_13665,N_9468,N_9926);
and U13666 (N_13666,N_10388,N_9984);
or U13667 (N_13667,N_10163,N_10050);
nor U13668 (N_13668,N_9258,N_10699);
nand U13669 (N_13669,N_9707,N_11278);
nand U13670 (N_13670,N_10187,N_10776);
nand U13671 (N_13671,N_10614,N_9061);
or U13672 (N_13672,N_11375,N_9415);
nor U13673 (N_13673,N_11818,N_10734);
or U13674 (N_13674,N_11399,N_10990);
nor U13675 (N_13675,N_11567,N_9045);
or U13676 (N_13676,N_11766,N_10927);
nor U13677 (N_13677,N_10226,N_9383);
and U13678 (N_13678,N_11965,N_10141);
and U13679 (N_13679,N_11485,N_10613);
and U13680 (N_13680,N_9522,N_11537);
or U13681 (N_13681,N_9281,N_10989);
nand U13682 (N_13682,N_9341,N_11479);
nand U13683 (N_13683,N_10451,N_10857);
nor U13684 (N_13684,N_10451,N_9255);
and U13685 (N_13685,N_9307,N_10656);
or U13686 (N_13686,N_10738,N_11114);
nand U13687 (N_13687,N_9568,N_9032);
or U13688 (N_13688,N_11828,N_9527);
nand U13689 (N_13689,N_11299,N_9850);
nor U13690 (N_13690,N_10108,N_9074);
or U13691 (N_13691,N_11818,N_10296);
and U13692 (N_13692,N_11704,N_10414);
and U13693 (N_13693,N_9025,N_11851);
nand U13694 (N_13694,N_11893,N_11087);
xor U13695 (N_13695,N_11622,N_10800);
nand U13696 (N_13696,N_10046,N_10900);
and U13697 (N_13697,N_11677,N_11321);
and U13698 (N_13698,N_9921,N_10816);
or U13699 (N_13699,N_9171,N_10812);
nor U13700 (N_13700,N_11531,N_9045);
nor U13701 (N_13701,N_10897,N_10189);
nand U13702 (N_13702,N_9152,N_11928);
nor U13703 (N_13703,N_11639,N_9196);
or U13704 (N_13704,N_11753,N_9638);
or U13705 (N_13705,N_10269,N_10624);
nor U13706 (N_13706,N_10961,N_10968);
nor U13707 (N_13707,N_9834,N_11590);
nand U13708 (N_13708,N_11974,N_10317);
nand U13709 (N_13709,N_10149,N_9357);
nor U13710 (N_13710,N_11028,N_10095);
nor U13711 (N_13711,N_9496,N_11435);
or U13712 (N_13712,N_9711,N_10516);
nand U13713 (N_13713,N_11973,N_9421);
or U13714 (N_13714,N_11826,N_9326);
nor U13715 (N_13715,N_9383,N_10104);
nand U13716 (N_13716,N_10409,N_10888);
nor U13717 (N_13717,N_9765,N_10681);
or U13718 (N_13718,N_10422,N_10010);
nand U13719 (N_13719,N_11498,N_11988);
and U13720 (N_13720,N_9859,N_10052);
or U13721 (N_13721,N_10174,N_9766);
and U13722 (N_13722,N_9130,N_9003);
nor U13723 (N_13723,N_10594,N_11847);
and U13724 (N_13724,N_9969,N_10396);
nor U13725 (N_13725,N_11980,N_9339);
and U13726 (N_13726,N_9798,N_10913);
or U13727 (N_13727,N_9189,N_11814);
or U13728 (N_13728,N_9489,N_11309);
nor U13729 (N_13729,N_9052,N_9267);
nor U13730 (N_13730,N_9864,N_9562);
nor U13731 (N_13731,N_9677,N_10361);
or U13732 (N_13732,N_10538,N_9053);
nor U13733 (N_13733,N_10917,N_9851);
nand U13734 (N_13734,N_9993,N_11471);
nor U13735 (N_13735,N_9579,N_10482);
and U13736 (N_13736,N_9570,N_9440);
nand U13737 (N_13737,N_9158,N_9450);
nand U13738 (N_13738,N_9076,N_10410);
nand U13739 (N_13739,N_9080,N_9303);
nor U13740 (N_13740,N_9191,N_10044);
nand U13741 (N_13741,N_10240,N_11409);
or U13742 (N_13742,N_10631,N_11688);
and U13743 (N_13743,N_9476,N_9491);
nand U13744 (N_13744,N_10342,N_11001);
and U13745 (N_13745,N_9408,N_10574);
nand U13746 (N_13746,N_9575,N_10178);
nor U13747 (N_13747,N_11335,N_10245);
nor U13748 (N_13748,N_9552,N_10374);
nand U13749 (N_13749,N_10699,N_9771);
or U13750 (N_13750,N_11048,N_10099);
nand U13751 (N_13751,N_9820,N_10153);
or U13752 (N_13752,N_10435,N_10211);
nor U13753 (N_13753,N_10833,N_11768);
nand U13754 (N_13754,N_9445,N_11157);
nand U13755 (N_13755,N_10992,N_10370);
nor U13756 (N_13756,N_9153,N_11781);
or U13757 (N_13757,N_11716,N_9772);
nand U13758 (N_13758,N_9559,N_11699);
nand U13759 (N_13759,N_9946,N_10286);
and U13760 (N_13760,N_11983,N_10073);
or U13761 (N_13761,N_9005,N_11654);
and U13762 (N_13762,N_11482,N_10779);
or U13763 (N_13763,N_9466,N_10453);
or U13764 (N_13764,N_11637,N_10114);
and U13765 (N_13765,N_10994,N_9874);
or U13766 (N_13766,N_11634,N_11487);
nand U13767 (N_13767,N_11017,N_10344);
and U13768 (N_13768,N_9938,N_11483);
nand U13769 (N_13769,N_10593,N_9898);
or U13770 (N_13770,N_9659,N_11609);
nand U13771 (N_13771,N_10643,N_9372);
or U13772 (N_13772,N_9450,N_11186);
or U13773 (N_13773,N_10750,N_10704);
and U13774 (N_13774,N_11566,N_10307);
and U13775 (N_13775,N_10525,N_10702);
nor U13776 (N_13776,N_11668,N_10575);
nand U13777 (N_13777,N_11703,N_11857);
or U13778 (N_13778,N_11484,N_10305);
nor U13779 (N_13779,N_9123,N_10438);
nand U13780 (N_13780,N_10847,N_11554);
and U13781 (N_13781,N_11649,N_10834);
nor U13782 (N_13782,N_9491,N_10516);
and U13783 (N_13783,N_10723,N_10746);
and U13784 (N_13784,N_9292,N_10355);
nand U13785 (N_13785,N_9837,N_9842);
nor U13786 (N_13786,N_11493,N_10849);
and U13787 (N_13787,N_11133,N_11761);
nor U13788 (N_13788,N_10193,N_9004);
nand U13789 (N_13789,N_11789,N_11758);
nand U13790 (N_13790,N_10774,N_9178);
nand U13791 (N_13791,N_9144,N_9859);
nor U13792 (N_13792,N_9563,N_10554);
nor U13793 (N_13793,N_9685,N_9161);
nand U13794 (N_13794,N_10115,N_10693);
and U13795 (N_13795,N_10007,N_9966);
nand U13796 (N_13796,N_10275,N_11302);
nor U13797 (N_13797,N_10159,N_10619);
or U13798 (N_13798,N_10013,N_11105);
nand U13799 (N_13799,N_11024,N_10915);
and U13800 (N_13800,N_10233,N_10750);
and U13801 (N_13801,N_10004,N_9544);
and U13802 (N_13802,N_10760,N_10082);
and U13803 (N_13803,N_11278,N_10281);
or U13804 (N_13804,N_10987,N_11916);
xnor U13805 (N_13805,N_10554,N_11883);
and U13806 (N_13806,N_11440,N_10224);
nor U13807 (N_13807,N_9636,N_10083);
or U13808 (N_13808,N_11569,N_9181);
nand U13809 (N_13809,N_10856,N_10464);
or U13810 (N_13810,N_11163,N_9284);
nand U13811 (N_13811,N_9128,N_10591);
or U13812 (N_13812,N_10931,N_11319);
and U13813 (N_13813,N_9073,N_10384);
or U13814 (N_13814,N_10693,N_9419);
nand U13815 (N_13815,N_9874,N_10375);
and U13816 (N_13816,N_9410,N_9454);
nand U13817 (N_13817,N_9910,N_9035);
and U13818 (N_13818,N_10503,N_10828);
or U13819 (N_13819,N_11614,N_9376);
or U13820 (N_13820,N_9667,N_10119);
and U13821 (N_13821,N_11622,N_10439);
nor U13822 (N_13822,N_10096,N_11803);
and U13823 (N_13823,N_9541,N_11849);
and U13824 (N_13824,N_9321,N_10496);
or U13825 (N_13825,N_9609,N_11361);
nand U13826 (N_13826,N_10882,N_11219);
and U13827 (N_13827,N_10271,N_10086);
nor U13828 (N_13828,N_9117,N_10824);
and U13829 (N_13829,N_11582,N_10955);
nor U13830 (N_13830,N_9657,N_10250);
or U13831 (N_13831,N_10263,N_11356);
and U13832 (N_13832,N_10015,N_11504);
or U13833 (N_13833,N_9874,N_10220);
nor U13834 (N_13834,N_10327,N_9011);
and U13835 (N_13835,N_9260,N_10775);
nand U13836 (N_13836,N_10479,N_11955);
and U13837 (N_13837,N_10183,N_9361);
and U13838 (N_13838,N_9412,N_9103);
nor U13839 (N_13839,N_10578,N_10153);
nor U13840 (N_13840,N_9280,N_11697);
nor U13841 (N_13841,N_9060,N_11191);
nor U13842 (N_13842,N_11817,N_10987);
nor U13843 (N_13843,N_10868,N_11830);
nor U13844 (N_13844,N_9561,N_10685);
nor U13845 (N_13845,N_9021,N_10808);
nor U13846 (N_13846,N_9397,N_10697);
nor U13847 (N_13847,N_9943,N_9367);
and U13848 (N_13848,N_10313,N_11946);
and U13849 (N_13849,N_10803,N_9634);
or U13850 (N_13850,N_11153,N_11459);
or U13851 (N_13851,N_11925,N_10994);
or U13852 (N_13852,N_9489,N_11026);
and U13853 (N_13853,N_9852,N_11045);
and U13854 (N_13854,N_10711,N_11901);
nor U13855 (N_13855,N_11047,N_11724);
nor U13856 (N_13856,N_10651,N_9107);
or U13857 (N_13857,N_10999,N_9203);
nand U13858 (N_13858,N_10929,N_9737);
or U13859 (N_13859,N_10691,N_10107);
xor U13860 (N_13860,N_9300,N_10167);
nor U13861 (N_13861,N_11321,N_11728);
or U13862 (N_13862,N_9527,N_10942);
and U13863 (N_13863,N_11351,N_9156);
nand U13864 (N_13864,N_9621,N_10700);
and U13865 (N_13865,N_11184,N_11249);
nor U13866 (N_13866,N_11174,N_10658);
and U13867 (N_13867,N_9789,N_10896);
and U13868 (N_13868,N_11246,N_10531);
nand U13869 (N_13869,N_11902,N_10508);
or U13870 (N_13870,N_9469,N_9139);
and U13871 (N_13871,N_10452,N_10533);
or U13872 (N_13872,N_9294,N_11785);
or U13873 (N_13873,N_11122,N_11294);
nor U13874 (N_13874,N_11446,N_10061);
nand U13875 (N_13875,N_9301,N_11646);
or U13876 (N_13876,N_11860,N_11227);
or U13877 (N_13877,N_10331,N_11750);
nor U13878 (N_13878,N_11623,N_10636);
or U13879 (N_13879,N_11919,N_9279);
or U13880 (N_13880,N_11648,N_9992);
nor U13881 (N_13881,N_9654,N_10823);
nor U13882 (N_13882,N_10550,N_9850);
nor U13883 (N_13883,N_11307,N_11239);
nand U13884 (N_13884,N_10723,N_11321);
nor U13885 (N_13885,N_10627,N_9481);
and U13886 (N_13886,N_9731,N_11856);
and U13887 (N_13887,N_11367,N_9785);
nand U13888 (N_13888,N_9594,N_9919);
or U13889 (N_13889,N_10121,N_10640);
nand U13890 (N_13890,N_9202,N_11930);
and U13891 (N_13891,N_9121,N_9757);
and U13892 (N_13892,N_10297,N_10016);
nor U13893 (N_13893,N_9089,N_10348);
and U13894 (N_13894,N_9594,N_9998);
nand U13895 (N_13895,N_11238,N_11163);
or U13896 (N_13896,N_9789,N_9277);
and U13897 (N_13897,N_9573,N_11743);
nor U13898 (N_13898,N_11929,N_11569);
and U13899 (N_13899,N_9663,N_11917);
or U13900 (N_13900,N_11744,N_10947);
nor U13901 (N_13901,N_10219,N_9693);
nand U13902 (N_13902,N_11058,N_11109);
nand U13903 (N_13903,N_11404,N_10845);
and U13904 (N_13904,N_11857,N_10342);
xnor U13905 (N_13905,N_10591,N_9634);
nor U13906 (N_13906,N_10873,N_11510);
nor U13907 (N_13907,N_10646,N_10239);
and U13908 (N_13908,N_10272,N_10582);
or U13909 (N_13909,N_11018,N_10301);
or U13910 (N_13910,N_10562,N_9303);
nand U13911 (N_13911,N_10155,N_9287);
and U13912 (N_13912,N_10797,N_11630);
nand U13913 (N_13913,N_11585,N_10270);
and U13914 (N_13914,N_10095,N_11997);
nor U13915 (N_13915,N_9846,N_10422);
nand U13916 (N_13916,N_10357,N_11000);
nand U13917 (N_13917,N_9541,N_11452);
and U13918 (N_13918,N_10636,N_9331);
or U13919 (N_13919,N_9052,N_9823);
nor U13920 (N_13920,N_9145,N_10662);
nand U13921 (N_13921,N_11671,N_9138);
xor U13922 (N_13922,N_10174,N_10042);
nor U13923 (N_13923,N_11797,N_11101);
or U13924 (N_13924,N_9854,N_11031);
and U13925 (N_13925,N_9979,N_9075);
nor U13926 (N_13926,N_11287,N_10095);
nor U13927 (N_13927,N_10776,N_11671);
nor U13928 (N_13928,N_11585,N_11543);
and U13929 (N_13929,N_9678,N_10320);
nor U13930 (N_13930,N_10241,N_11443);
nor U13931 (N_13931,N_9159,N_9788);
nand U13932 (N_13932,N_10391,N_9639);
and U13933 (N_13933,N_11357,N_9398);
or U13934 (N_13934,N_10787,N_9042);
nor U13935 (N_13935,N_9217,N_10987);
and U13936 (N_13936,N_11543,N_9702);
and U13937 (N_13937,N_11232,N_9179);
nand U13938 (N_13938,N_9045,N_11664);
and U13939 (N_13939,N_10083,N_9083);
and U13940 (N_13940,N_10354,N_11108);
or U13941 (N_13941,N_9142,N_11553);
nor U13942 (N_13942,N_11038,N_9903);
and U13943 (N_13943,N_11069,N_11156);
nor U13944 (N_13944,N_11068,N_11200);
nand U13945 (N_13945,N_9590,N_9005);
nor U13946 (N_13946,N_11186,N_10725);
and U13947 (N_13947,N_11148,N_11942);
and U13948 (N_13948,N_10268,N_10330);
and U13949 (N_13949,N_10090,N_11423);
and U13950 (N_13950,N_9145,N_11845);
or U13951 (N_13951,N_10329,N_11149);
or U13952 (N_13952,N_11816,N_9110);
nand U13953 (N_13953,N_9049,N_11678);
or U13954 (N_13954,N_11098,N_11197);
or U13955 (N_13955,N_11425,N_11987);
and U13956 (N_13956,N_9967,N_10995);
xor U13957 (N_13957,N_9463,N_11216);
and U13958 (N_13958,N_10332,N_10865);
nor U13959 (N_13959,N_9174,N_9371);
and U13960 (N_13960,N_11562,N_10632);
and U13961 (N_13961,N_11358,N_10906);
nand U13962 (N_13962,N_10362,N_10718);
and U13963 (N_13963,N_9511,N_9941);
or U13964 (N_13964,N_9555,N_11184);
nand U13965 (N_13965,N_10991,N_10376);
or U13966 (N_13966,N_10935,N_10280);
or U13967 (N_13967,N_9908,N_9876);
or U13968 (N_13968,N_10029,N_10430);
nand U13969 (N_13969,N_10140,N_9714);
or U13970 (N_13970,N_10209,N_11481);
and U13971 (N_13971,N_11688,N_9751);
nor U13972 (N_13972,N_9753,N_11907);
and U13973 (N_13973,N_9767,N_9834);
nand U13974 (N_13974,N_10175,N_9513);
nand U13975 (N_13975,N_11803,N_10504);
nor U13976 (N_13976,N_9043,N_9896);
nor U13977 (N_13977,N_10063,N_10230);
nand U13978 (N_13978,N_11478,N_11447);
nand U13979 (N_13979,N_11584,N_11482);
nor U13980 (N_13980,N_9573,N_9095);
and U13981 (N_13981,N_9807,N_10596);
or U13982 (N_13982,N_11510,N_10881);
or U13983 (N_13983,N_11149,N_9219);
and U13984 (N_13984,N_11409,N_11964);
nand U13985 (N_13985,N_11646,N_11685);
nor U13986 (N_13986,N_9218,N_10180);
nor U13987 (N_13987,N_10879,N_11661);
and U13988 (N_13988,N_9493,N_10734);
nor U13989 (N_13989,N_10579,N_9810);
and U13990 (N_13990,N_9502,N_11551);
or U13991 (N_13991,N_9735,N_11388);
or U13992 (N_13992,N_10155,N_11168);
nor U13993 (N_13993,N_9543,N_10881);
or U13994 (N_13994,N_9136,N_11520);
nor U13995 (N_13995,N_11330,N_10422);
or U13996 (N_13996,N_11841,N_11471);
and U13997 (N_13997,N_10778,N_11360);
xnor U13998 (N_13998,N_11582,N_9851);
nor U13999 (N_13999,N_9674,N_11077);
nand U14000 (N_14000,N_9983,N_11935);
nand U14001 (N_14001,N_11702,N_10166);
nor U14002 (N_14002,N_11518,N_10011);
and U14003 (N_14003,N_11138,N_11653);
and U14004 (N_14004,N_10803,N_10123);
and U14005 (N_14005,N_11348,N_9808);
and U14006 (N_14006,N_10292,N_11959);
nand U14007 (N_14007,N_11671,N_9620);
and U14008 (N_14008,N_9041,N_9109);
or U14009 (N_14009,N_11920,N_10229);
and U14010 (N_14010,N_9216,N_10656);
and U14011 (N_14011,N_11459,N_11422);
or U14012 (N_14012,N_9295,N_9416);
nor U14013 (N_14013,N_9224,N_9450);
nand U14014 (N_14014,N_10335,N_10760);
nand U14015 (N_14015,N_9513,N_9329);
nor U14016 (N_14016,N_9683,N_9335);
or U14017 (N_14017,N_9766,N_10339);
or U14018 (N_14018,N_11466,N_9598);
and U14019 (N_14019,N_10317,N_11001);
nand U14020 (N_14020,N_11390,N_9240);
and U14021 (N_14021,N_9168,N_9540);
nor U14022 (N_14022,N_11265,N_9303);
or U14023 (N_14023,N_11958,N_9781);
nand U14024 (N_14024,N_11326,N_9625);
nor U14025 (N_14025,N_9792,N_10695);
nand U14026 (N_14026,N_9579,N_11256);
nand U14027 (N_14027,N_9816,N_9486);
nand U14028 (N_14028,N_9584,N_11864);
and U14029 (N_14029,N_9692,N_10187);
or U14030 (N_14030,N_10875,N_11654);
nand U14031 (N_14031,N_10902,N_9296);
nand U14032 (N_14032,N_11311,N_10941);
nor U14033 (N_14033,N_10380,N_11670);
nand U14034 (N_14034,N_11155,N_11208);
nand U14035 (N_14035,N_11821,N_10937);
nor U14036 (N_14036,N_9675,N_9106);
or U14037 (N_14037,N_9990,N_11895);
nand U14038 (N_14038,N_9635,N_9747);
nor U14039 (N_14039,N_11568,N_11344);
nor U14040 (N_14040,N_9533,N_10995);
or U14041 (N_14041,N_9616,N_9552);
nor U14042 (N_14042,N_9070,N_9275);
nor U14043 (N_14043,N_11648,N_10836);
nand U14044 (N_14044,N_9141,N_9247);
nand U14045 (N_14045,N_11013,N_11885);
and U14046 (N_14046,N_11170,N_9524);
and U14047 (N_14047,N_9507,N_9130);
and U14048 (N_14048,N_11865,N_11164);
nor U14049 (N_14049,N_10372,N_10127);
nand U14050 (N_14050,N_10337,N_11517);
nor U14051 (N_14051,N_9933,N_9802);
nor U14052 (N_14052,N_10169,N_11273);
nor U14053 (N_14053,N_10382,N_10803);
or U14054 (N_14054,N_10413,N_9443);
nand U14055 (N_14055,N_10391,N_10335);
or U14056 (N_14056,N_11868,N_10909);
or U14057 (N_14057,N_11319,N_10920);
nor U14058 (N_14058,N_9130,N_10766);
and U14059 (N_14059,N_10464,N_10022);
nand U14060 (N_14060,N_11021,N_9047);
nand U14061 (N_14061,N_11502,N_10310);
nand U14062 (N_14062,N_10591,N_10823);
or U14063 (N_14063,N_10675,N_10013);
nand U14064 (N_14064,N_11404,N_10689);
nand U14065 (N_14065,N_10259,N_11037);
nand U14066 (N_14066,N_10822,N_9938);
nor U14067 (N_14067,N_9970,N_9807);
and U14068 (N_14068,N_9873,N_10015);
or U14069 (N_14069,N_9934,N_9143);
nor U14070 (N_14070,N_11598,N_9305);
nand U14071 (N_14071,N_10752,N_11046);
nand U14072 (N_14072,N_9566,N_10573);
nor U14073 (N_14073,N_9634,N_10293);
and U14074 (N_14074,N_11557,N_10569);
nor U14075 (N_14075,N_11524,N_9193);
and U14076 (N_14076,N_9360,N_9775);
nor U14077 (N_14077,N_10412,N_10212);
nor U14078 (N_14078,N_10072,N_10508);
and U14079 (N_14079,N_11945,N_9800);
nand U14080 (N_14080,N_11783,N_10781);
nor U14081 (N_14081,N_10693,N_9107);
nand U14082 (N_14082,N_10022,N_9062);
and U14083 (N_14083,N_11225,N_10077);
and U14084 (N_14084,N_10845,N_10396);
nor U14085 (N_14085,N_10430,N_10899);
and U14086 (N_14086,N_9955,N_10219);
nand U14087 (N_14087,N_10206,N_10182);
or U14088 (N_14088,N_10884,N_9549);
nand U14089 (N_14089,N_10417,N_9931);
nor U14090 (N_14090,N_11374,N_9118);
nand U14091 (N_14091,N_11639,N_10806);
nor U14092 (N_14092,N_9104,N_9040);
and U14093 (N_14093,N_10908,N_10821);
nor U14094 (N_14094,N_9752,N_9935);
and U14095 (N_14095,N_9330,N_9362);
and U14096 (N_14096,N_9922,N_10468);
nor U14097 (N_14097,N_10326,N_11266);
nor U14098 (N_14098,N_11225,N_11621);
and U14099 (N_14099,N_9859,N_10905);
and U14100 (N_14100,N_9689,N_10463);
or U14101 (N_14101,N_9391,N_9675);
nor U14102 (N_14102,N_10854,N_10786);
and U14103 (N_14103,N_11089,N_9652);
or U14104 (N_14104,N_10443,N_10472);
nor U14105 (N_14105,N_9849,N_10984);
nor U14106 (N_14106,N_9099,N_11840);
nand U14107 (N_14107,N_11959,N_10033);
nor U14108 (N_14108,N_10438,N_9684);
nor U14109 (N_14109,N_10395,N_10335);
and U14110 (N_14110,N_9735,N_9749);
nand U14111 (N_14111,N_11659,N_11617);
nor U14112 (N_14112,N_10438,N_10020);
and U14113 (N_14113,N_11867,N_9356);
and U14114 (N_14114,N_11850,N_10440);
nor U14115 (N_14115,N_11330,N_11891);
or U14116 (N_14116,N_11433,N_10995);
nand U14117 (N_14117,N_9934,N_10740);
or U14118 (N_14118,N_11555,N_10741);
and U14119 (N_14119,N_9399,N_9435);
nor U14120 (N_14120,N_10841,N_10827);
or U14121 (N_14121,N_9662,N_10270);
and U14122 (N_14122,N_9006,N_10067);
or U14123 (N_14123,N_11765,N_9767);
and U14124 (N_14124,N_10776,N_11101);
nand U14125 (N_14125,N_10118,N_9601);
and U14126 (N_14126,N_9298,N_11207);
or U14127 (N_14127,N_11567,N_10854);
and U14128 (N_14128,N_9158,N_9921);
or U14129 (N_14129,N_11950,N_9876);
nand U14130 (N_14130,N_11730,N_9813);
nand U14131 (N_14131,N_10199,N_11047);
nand U14132 (N_14132,N_9000,N_11182);
and U14133 (N_14133,N_10017,N_10124);
and U14134 (N_14134,N_11484,N_11611);
nand U14135 (N_14135,N_10054,N_9082);
nand U14136 (N_14136,N_9270,N_9914);
nor U14137 (N_14137,N_9746,N_10572);
and U14138 (N_14138,N_10506,N_9405);
and U14139 (N_14139,N_10836,N_10997);
nand U14140 (N_14140,N_11823,N_10496);
nor U14141 (N_14141,N_11679,N_10218);
or U14142 (N_14142,N_10013,N_11226);
or U14143 (N_14143,N_10400,N_11836);
nand U14144 (N_14144,N_11124,N_10135);
nor U14145 (N_14145,N_10095,N_9097);
or U14146 (N_14146,N_10261,N_11940);
nor U14147 (N_14147,N_11061,N_11511);
or U14148 (N_14148,N_9202,N_9046);
nor U14149 (N_14149,N_10206,N_11135);
nor U14150 (N_14150,N_10079,N_9080);
nor U14151 (N_14151,N_9275,N_9089);
and U14152 (N_14152,N_9106,N_11925);
nor U14153 (N_14153,N_9226,N_9197);
or U14154 (N_14154,N_11045,N_10255);
and U14155 (N_14155,N_10078,N_10982);
nand U14156 (N_14156,N_11857,N_11153);
nand U14157 (N_14157,N_10679,N_11256);
nor U14158 (N_14158,N_9650,N_9041);
and U14159 (N_14159,N_11457,N_11323);
or U14160 (N_14160,N_10622,N_9614);
or U14161 (N_14161,N_10986,N_9055);
and U14162 (N_14162,N_9970,N_10721);
nor U14163 (N_14163,N_9786,N_9892);
nor U14164 (N_14164,N_10098,N_11618);
and U14165 (N_14165,N_9990,N_11922);
nor U14166 (N_14166,N_11856,N_11277);
nor U14167 (N_14167,N_9304,N_10367);
and U14168 (N_14168,N_9483,N_9390);
and U14169 (N_14169,N_9942,N_9620);
nand U14170 (N_14170,N_11225,N_9426);
and U14171 (N_14171,N_9463,N_10714);
nand U14172 (N_14172,N_9956,N_9479);
and U14173 (N_14173,N_9097,N_9106);
or U14174 (N_14174,N_10310,N_11470);
and U14175 (N_14175,N_11689,N_10875);
and U14176 (N_14176,N_9856,N_11593);
nand U14177 (N_14177,N_9998,N_10837);
xor U14178 (N_14178,N_10575,N_10014);
and U14179 (N_14179,N_11025,N_10991);
nor U14180 (N_14180,N_10162,N_10974);
or U14181 (N_14181,N_11817,N_10731);
or U14182 (N_14182,N_11125,N_10561);
nand U14183 (N_14183,N_9630,N_11495);
nor U14184 (N_14184,N_11385,N_11163);
nand U14185 (N_14185,N_11509,N_9586);
nor U14186 (N_14186,N_11874,N_10723);
nor U14187 (N_14187,N_11287,N_9757);
xnor U14188 (N_14188,N_9656,N_9251);
nand U14189 (N_14189,N_9358,N_9806);
nor U14190 (N_14190,N_11018,N_9122);
nand U14191 (N_14191,N_9662,N_10193);
nor U14192 (N_14192,N_10844,N_10430);
nor U14193 (N_14193,N_9076,N_9790);
nor U14194 (N_14194,N_11606,N_11835);
or U14195 (N_14195,N_10740,N_9008);
and U14196 (N_14196,N_9700,N_11632);
and U14197 (N_14197,N_11298,N_11667);
and U14198 (N_14198,N_11519,N_10436);
nand U14199 (N_14199,N_11113,N_10418);
nor U14200 (N_14200,N_11877,N_10250);
nand U14201 (N_14201,N_9516,N_9540);
nor U14202 (N_14202,N_10477,N_11236);
and U14203 (N_14203,N_11760,N_9792);
and U14204 (N_14204,N_9275,N_10954);
and U14205 (N_14205,N_11128,N_11078);
and U14206 (N_14206,N_9585,N_9508);
nor U14207 (N_14207,N_10528,N_11640);
nand U14208 (N_14208,N_11813,N_11488);
and U14209 (N_14209,N_9168,N_10157);
and U14210 (N_14210,N_11592,N_10996);
or U14211 (N_14211,N_10280,N_9619);
nor U14212 (N_14212,N_11694,N_11242);
nand U14213 (N_14213,N_10189,N_9791);
or U14214 (N_14214,N_9448,N_11658);
nor U14215 (N_14215,N_9408,N_11181);
and U14216 (N_14216,N_9619,N_9039);
nor U14217 (N_14217,N_10229,N_11704);
xor U14218 (N_14218,N_9585,N_10767);
and U14219 (N_14219,N_11580,N_9694);
or U14220 (N_14220,N_9608,N_9754);
nand U14221 (N_14221,N_9499,N_11243);
and U14222 (N_14222,N_9412,N_11441);
nand U14223 (N_14223,N_10509,N_9864);
xor U14224 (N_14224,N_9659,N_11818);
nor U14225 (N_14225,N_9428,N_10628);
and U14226 (N_14226,N_11309,N_9642);
or U14227 (N_14227,N_9059,N_11428);
nand U14228 (N_14228,N_9388,N_10174);
or U14229 (N_14229,N_10691,N_11951);
nor U14230 (N_14230,N_11959,N_10573);
or U14231 (N_14231,N_10510,N_11062);
nor U14232 (N_14232,N_11423,N_9786);
or U14233 (N_14233,N_9897,N_9059);
nand U14234 (N_14234,N_10319,N_10309);
nand U14235 (N_14235,N_11007,N_11740);
and U14236 (N_14236,N_10968,N_9759);
or U14237 (N_14237,N_9063,N_10796);
and U14238 (N_14238,N_11691,N_10501);
or U14239 (N_14239,N_10562,N_11554);
and U14240 (N_14240,N_10959,N_11811);
or U14241 (N_14241,N_11825,N_9587);
or U14242 (N_14242,N_11413,N_9059);
nand U14243 (N_14243,N_9845,N_9130);
and U14244 (N_14244,N_11069,N_11234);
nor U14245 (N_14245,N_11584,N_9135);
and U14246 (N_14246,N_10561,N_11030);
or U14247 (N_14247,N_11789,N_11615);
or U14248 (N_14248,N_10940,N_11457);
nand U14249 (N_14249,N_9324,N_9367);
and U14250 (N_14250,N_11697,N_10080);
nor U14251 (N_14251,N_9536,N_10874);
nand U14252 (N_14252,N_9233,N_10541);
nand U14253 (N_14253,N_10983,N_10288);
or U14254 (N_14254,N_9114,N_10779);
nand U14255 (N_14255,N_10529,N_10282);
or U14256 (N_14256,N_10372,N_11706);
nor U14257 (N_14257,N_11613,N_9308);
and U14258 (N_14258,N_11155,N_9506);
nor U14259 (N_14259,N_9190,N_10940);
nor U14260 (N_14260,N_10047,N_9999);
nand U14261 (N_14261,N_10934,N_9388);
or U14262 (N_14262,N_10425,N_11785);
and U14263 (N_14263,N_10809,N_11755);
and U14264 (N_14264,N_10258,N_10303);
nor U14265 (N_14265,N_9910,N_10700);
and U14266 (N_14266,N_11766,N_10041);
and U14267 (N_14267,N_11991,N_10871);
nor U14268 (N_14268,N_9875,N_9671);
and U14269 (N_14269,N_9999,N_9275);
and U14270 (N_14270,N_11587,N_10934);
nand U14271 (N_14271,N_11196,N_9311);
and U14272 (N_14272,N_10229,N_10379);
nor U14273 (N_14273,N_11762,N_9121);
nand U14274 (N_14274,N_10373,N_11292);
and U14275 (N_14275,N_9989,N_11360);
or U14276 (N_14276,N_9569,N_10593);
and U14277 (N_14277,N_11083,N_11214);
and U14278 (N_14278,N_10141,N_10208);
or U14279 (N_14279,N_11019,N_11046);
nor U14280 (N_14280,N_9240,N_11095);
or U14281 (N_14281,N_11853,N_11208);
or U14282 (N_14282,N_11281,N_9562);
nor U14283 (N_14283,N_11257,N_11796);
and U14284 (N_14284,N_9698,N_11482);
nor U14285 (N_14285,N_11107,N_11211);
nor U14286 (N_14286,N_9157,N_11570);
nand U14287 (N_14287,N_10262,N_9484);
and U14288 (N_14288,N_10654,N_10867);
or U14289 (N_14289,N_10719,N_11867);
nor U14290 (N_14290,N_10506,N_9613);
and U14291 (N_14291,N_10752,N_9605);
and U14292 (N_14292,N_11294,N_10449);
xnor U14293 (N_14293,N_9472,N_11685);
nor U14294 (N_14294,N_11077,N_11663);
nand U14295 (N_14295,N_10798,N_10469);
or U14296 (N_14296,N_9893,N_10168);
nor U14297 (N_14297,N_11826,N_11560);
and U14298 (N_14298,N_11223,N_10809);
or U14299 (N_14299,N_9375,N_9199);
nand U14300 (N_14300,N_11244,N_9305);
nand U14301 (N_14301,N_11863,N_9769);
or U14302 (N_14302,N_11725,N_9594);
and U14303 (N_14303,N_9247,N_11946);
or U14304 (N_14304,N_9936,N_11394);
and U14305 (N_14305,N_9786,N_9908);
and U14306 (N_14306,N_11929,N_9521);
or U14307 (N_14307,N_9906,N_10419);
and U14308 (N_14308,N_11385,N_11273);
nand U14309 (N_14309,N_10739,N_10262);
and U14310 (N_14310,N_10147,N_10764);
or U14311 (N_14311,N_9411,N_9282);
and U14312 (N_14312,N_9520,N_11781);
and U14313 (N_14313,N_9447,N_10443);
or U14314 (N_14314,N_10812,N_11523);
nor U14315 (N_14315,N_10936,N_10363);
nand U14316 (N_14316,N_9236,N_10318);
and U14317 (N_14317,N_9865,N_10068);
and U14318 (N_14318,N_9847,N_10065);
and U14319 (N_14319,N_9364,N_9878);
nor U14320 (N_14320,N_9553,N_10475);
nand U14321 (N_14321,N_10078,N_10129);
nand U14322 (N_14322,N_11090,N_11947);
or U14323 (N_14323,N_10679,N_10792);
and U14324 (N_14324,N_9085,N_10366);
and U14325 (N_14325,N_10326,N_10793);
nor U14326 (N_14326,N_10964,N_10554);
or U14327 (N_14327,N_11903,N_11537);
and U14328 (N_14328,N_11158,N_11353);
xnor U14329 (N_14329,N_9087,N_10966);
and U14330 (N_14330,N_9254,N_10592);
nand U14331 (N_14331,N_9514,N_11078);
nand U14332 (N_14332,N_10624,N_9346);
and U14333 (N_14333,N_11656,N_9451);
and U14334 (N_14334,N_11750,N_11712);
or U14335 (N_14335,N_11455,N_9566);
or U14336 (N_14336,N_11206,N_11259);
nor U14337 (N_14337,N_11448,N_9487);
nor U14338 (N_14338,N_9163,N_10836);
and U14339 (N_14339,N_10702,N_10610);
and U14340 (N_14340,N_10152,N_11129);
and U14341 (N_14341,N_9149,N_10808);
nor U14342 (N_14342,N_10855,N_9151);
nand U14343 (N_14343,N_10848,N_9363);
or U14344 (N_14344,N_9281,N_9882);
or U14345 (N_14345,N_9980,N_9990);
and U14346 (N_14346,N_10699,N_9116);
and U14347 (N_14347,N_9482,N_10562);
nor U14348 (N_14348,N_10520,N_11837);
and U14349 (N_14349,N_9268,N_11322);
or U14350 (N_14350,N_9535,N_11623);
or U14351 (N_14351,N_10076,N_11933);
nand U14352 (N_14352,N_11636,N_9509);
or U14353 (N_14353,N_11739,N_10747);
nor U14354 (N_14354,N_11852,N_10364);
nand U14355 (N_14355,N_11508,N_11130);
and U14356 (N_14356,N_11407,N_9628);
or U14357 (N_14357,N_10529,N_11962);
and U14358 (N_14358,N_9381,N_11235);
or U14359 (N_14359,N_10794,N_10963);
nand U14360 (N_14360,N_10858,N_9508);
nand U14361 (N_14361,N_11575,N_9153);
nand U14362 (N_14362,N_11079,N_9021);
nand U14363 (N_14363,N_10531,N_10433);
and U14364 (N_14364,N_10679,N_10113);
nand U14365 (N_14365,N_10183,N_11996);
and U14366 (N_14366,N_11734,N_11439);
and U14367 (N_14367,N_9716,N_9677);
and U14368 (N_14368,N_11860,N_11902);
nor U14369 (N_14369,N_11904,N_9347);
or U14370 (N_14370,N_10686,N_10156);
or U14371 (N_14371,N_10264,N_9808);
and U14372 (N_14372,N_11478,N_11917);
and U14373 (N_14373,N_9688,N_10602);
or U14374 (N_14374,N_10101,N_11080);
and U14375 (N_14375,N_10151,N_9332);
nor U14376 (N_14376,N_10404,N_9416);
nand U14377 (N_14377,N_10681,N_9348);
or U14378 (N_14378,N_10450,N_9379);
nor U14379 (N_14379,N_10787,N_9777);
nand U14380 (N_14380,N_11737,N_11214);
xnor U14381 (N_14381,N_10783,N_9333);
and U14382 (N_14382,N_11435,N_11976);
and U14383 (N_14383,N_9748,N_10232);
nand U14384 (N_14384,N_10229,N_10853);
nor U14385 (N_14385,N_10388,N_9597);
nor U14386 (N_14386,N_11944,N_10790);
and U14387 (N_14387,N_9857,N_11140);
nor U14388 (N_14388,N_11385,N_11444);
and U14389 (N_14389,N_9597,N_10981);
nand U14390 (N_14390,N_11760,N_11650);
and U14391 (N_14391,N_11992,N_11645);
nand U14392 (N_14392,N_11584,N_9940);
nand U14393 (N_14393,N_9629,N_9816);
nor U14394 (N_14394,N_9474,N_9301);
nand U14395 (N_14395,N_9905,N_9432);
and U14396 (N_14396,N_11603,N_9706);
and U14397 (N_14397,N_11548,N_10668);
and U14398 (N_14398,N_10691,N_9434);
nand U14399 (N_14399,N_9249,N_10404);
nand U14400 (N_14400,N_10289,N_10938);
or U14401 (N_14401,N_10216,N_10405);
and U14402 (N_14402,N_11977,N_11603);
and U14403 (N_14403,N_9993,N_11021);
nor U14404 (N_14404,N_11491,N_9515);
or U14405 (N_14405,N_9903,N_10588);
or U14406 (N_14406,N_10748,N_10409);
and U14407 (N_14407,N_9573,N_11300);
and U14408 (N_14408,N_10636,N_10558);
nand U14409 (N_14409,N_9933,N_9711);
nor U14410 (N_14410,N_9650,N_11629);
or U14411 (N_14411,N_11712,N_9559);
nor U14412 (N_14412,N_11371,N_11563);
and U14413 (N_14413,N_10320,N_10105);
or U14414 (N_14414,N_11540,N_9382);
and U14415 (N_14415,N_9423,N_11045);
and U14416 (N_14416,N_11749,N_9709);
and U14417 (N_14417,N_9528,N_11607);
nand U14418 (N_14418,N_11560,N_9979);
nand U14419 (N_14419,N_9812,N_11079);
nor U14420 (N_14420,N_9498,N_11549);
nand U14421 (N_14421,N_10156,N_10709);
and U14422 (N_14422,N_9033,N_10925);
and U14423 (N_14423,N_11941,N_11228);
and U14424 (N_14424,N_9332,N_10097);
nor U14425 (N_14425,N_10668,N_11329);
and U14426 (N_14426,N_10995,N_11967);
nor U14427 (N_14427,N_9804,N_11043);
nor U14428 (N_14428,N_11833,N_10684);
and U14429 (N_14429,N_10410,N_9289);
or U14430 (N_14430,N_9455,N_9532);
nand U14431 (N_14431,N_11752,N_11443);
or U14432 (N_14432,N_11890,N_11190);
or U14433 (N_14433,N_9673,N_11398);
or U14434 (N_14434,N_11478,N_9791);
or U14435 (N_14435,N_10009,N_11589);
or U14436 (N_14436,N_11644,N_10507);
nor U14437 (N_14437,N_10405,N_11146);
nor U14438 (N_14438,N_10672,N_9879);
nor U14439 (N_14439,N_10950,N_11240);
and U14440 (N_14440,N_10030,N_11328);
and U14441 (N_14441,N_10657,N_10887);
or U14442 (N_14442,N_10693,N_11280);
or U14443 (N_14443,N_10062,N_10778);
nand U14444 (N_14444,N_10152,N_10285);
or U14445 (N_14445,N_9989,N_11488);
nand U14446 (N_14446,N_11016,N_10084);
nor U14447 (N_14447,N_11519,N_10116);
nand U14448 (N_14448,N_11288,N_10317);
nor U14449 (N_14449,N_10051,N_10874);
nand U14450 (N_14450,N_11972,N_11178);
and U14451 (N_14451,N_9588,N_9359);
and U14452 (N_14452,N_9746,N_10015);
or U14453 (N_14453,N_9142,N_9285);
or U14454 (N_14454,N_10157,N_9977);
nand U14455 (N_14455,N_11317,N_10003);
or U14456 (N_14456,N_10209,N_9490);
xor U14457 (N_14457,N_10991,N_10208);
nand U14458 (N_14458,N_11353,N_10474);
nor U14459 (N_14459,N_9909,N_9658);
nand U14460 (N_14460,N_10988,N_11757);
or U14461 (N_14461,N_11870,N_11334);
nor U14462 (N_14462,N_10584,N_9941);
nor U14463 (N_14463,N_9498,N_9341);
nor U14464 (N_14464,N_10100,N_10309);
and U14465 (N_14465,N_11079,N_10140);
nand U14466 (N_14466,N_9809,N_10772);
or U14467 (N_14467,N_10044,N_10251);
nor U14468 (N_14468,N_9042,N_9133);
or U14469 (N_14469,N_10298,N_10527);
or U14470 (N_14470,N_10413,N_10939);
and U14471 (N_14471,N_11433,N_11163);
or U14472 (N_14472,N_10734,N_9890);
and U14473 (N_14473,N_11184,N_11012);
nor U14474 (N_14474,N_10309,N_10760);
nor U14475 (N_14475,N_10666,N_9795);
nor U14476 (N_14476,N_10662,N_11628);
nand U14477 (N_14477,N_11859,N_10306);
nand U14478 (N_14478,N_10221,N_9452);
nor U14479 (N_14479,N_10559,N_11173);
nand U14480 (N_14480,N_10186,N_9796);
nand U14481 (N_14481,N_10197,N_10603);
and U14482 (N_14482,N_10559,N_10328);
or U14483 (N_14483,N_10529,N_11393);
or U14484 (N_14484,N_10113,N_10901);
and U14485 (N_14485,N_11768,N_11596);
nand U14486 (N_14486,N_11777,N_11981);
or U14487 (N_14487,N_9396,N_9851);
or U14488 (N_14488,N_9169,N_9321);
and U14489 (N_14489,N_9008,N_10511);
nor U14490 (N_14490,N_9992,N_9737);
and U14491 (N_14491,N_9399,N_9518);
xnor U14492 (N_14492,N_11519,N_11871);
and U14493 (N_14493,N_9841,N_9524);
nor U14494 (N_14494,N_11770,N_10961);
and U14495 (N_14495,N_9608,N_9259);
and U14496 (N_14496,N_10371,N_11508);
nor U14497 (N_14497,N_11836,N_9799);
nand U14498 (N_14498,N_9356,N_10474);
nor U14499 (N_14499,N_11694,N_9488);
and U14500 (N_14500,N_10738,N_9879);
nor U14501 (N_14501,N_9069,N_10837);
and U14502 (N_14502,N_11545,N_9741);
and U14503 (N_14503,N_9646,N_10526);
and U14504 (N_14504,N_9977,N_10723);
nor U14505 (N_14505,N_11506,N_10009);
nor U14506 (N_14506,N_10782,N_9135);
nor U14507 (N_14507,N_9846,N_9454);
or U14508 (N_14508,N_11868,N_9847);
or U14509 (N_14509,N_9210,N_10303);
and U14510 (N_14510,N_9039,N_10380);
and U14511 (N_14511,N_9286,N_9598);
or U14512 (N_14512,N_10502,N_10568);
and U14513 (N_14513,N_9216,N_11111);
and U14514 (N_14514,N_10389,N_11721);
nand U14515 (N_14515,N_10825,N_11641);
nor U14516 (N_14516,N_9944,N_10479);
or U14517 (N_14517,N_11363,N_11789);
nor U14518 (N_14518,N_11511,N_9495);
or U14519 (N_14519,N_10096,N_10847);
or U14520 (N_14520,N_9510,N_10944);
or U14521 (N_14521,N_11756,N_11419);
or U14522 (N_14522,N_9348,N_10609);
nand U14523 (N_14523,N_11512,N_11483);
or U14524 (N_14524,N_11832,N_10270);
nor U14525 (N_14525,N_10095,N_10582);
or U14526 (N_14526,N_11196,N_11405);
nand U14527 (N_14527,N_9901,N_9555);
nand U14528 (N_14528,N_10160,N_9475);
and U14529 (N_14529,N_10810,N_10191);
nand U14530 (N_14530,N_10900,N_10937);
nor U14531 (N_14531,N_11629,N_11830);
and U14532 (N_14532,N_11254,N_11927);
or U14533 (N_14533,N_10765,N_10996);
nor U14534 (N_14534,N_11948,N_9137);
and U14535 (N_14535,N_9154,N_9361);
nor U14536 (N_14536,N_9576,N_11631);
nor U14537 (N_14537,N_9518,N_10659);
or U14538 (N_14538,N_9956,N_10519);
nor U14539 (N_14539,N_10873,N_11083);
nand U14540 (N_14540,N_9972,N_9704);
nor U14541 (N_14541,N_10871,N_10778);
and U14542 (N_14542,N_9287,N_10265);
nand U14543 (N_14543,N_11881,N_9882);
or U14544 (N_14544,N_9164,N_11343);
nor U14545 (N_14545,N_11704,N_11032);
nor U14546 (N_14546,N_9389,N_10924);
nand U14547 (N_14547,N_9165,N_10634);
nand U14548 (N_14548,N_9897,N_9337);
nand U14549 (N_14549,N_11152,N_9786);
nor U14550 (N_14550,N_10775,N_11941);
nand U14551 (N_14551,N_9641,N_11318);
or U14552 (N_14552,N_11641,N_9074);
nor U14553 (N_14553,N_11592,N_11537);
nand U14554 (N_14554,N_9590,N_11275);
or U14555 (N_14555,N_10481,N_9049);
nand U14556 (N_14556,N_11041,N_10106);
or U14557 (N_14557,N_11087,N_11806);
nand U14558 (N_14558,N_10907,N_10557);
or U14559 (N_14559,N_9821,N_11435);
nor U14560 (N_14560,N_10144,N_10680);
or U14561 (N_14561,N_9120,N_10335);
nand U14562 (N_14562,N_10596,N_11618);
and U14563 (N_14563,N_9333,N_11038);
or U14564 (N_14564,N_11553,N_9473);
nand U14565 (N_14565,N_11254,N_10796);
nand U14566 (N_14566,N_11912,N_10453);
nand U14567 (N_14567,N_11684,N_10479);
or U14568 (N_14568,N_10098,N_9972);
nor U14569 (N_14569,N_11572,N_11703);
nand U14570 (N_14570,N_9654,N_11192);
nand U14571 (N_14571,N_10021,N_11084);
and U14572 (N_14572,N_11004,N_11507);
nor U14573 (N_14573,N_11313,N_10591);
nand U14574 (N_14574,N_11015,N_9148);
and U14575 (N_14575,N_10591,N_9822);
nor U14576 (N_14576,N_10376,N_11754);
nor U14577 (N_14577,N_9803,N_9348);
and U14578 (N_14578,N_10522,N_9054);
and U14579 (N_14579,N_11153,N_10747);
and U14580 (N_14580,N_10983,N_9700);
nand U14581 (N_14581,N_9867,N_11743);
nor U14582 (N_14582,N_11825,N_10583);
nor U14583 (N_14583,N_9424,N_10520);
nor U14584 (N_14584,N_10012,N_11876);
nor U14585 (N_14585,N_10050,N_11765);
nor U14586 (N_14586,N_10222,N_9828);
nand U14587 (N_14587,N_9535,N_11272);
or U14588 (N_14588,N_9725,N_10725);
nand U14589 (N_14589,N_10154,N_10980);
nor U14590 (N_14590,N_10464,N_9406);
nand U14591 (N_14591,N_10827,N_11450);
nor U14592 (N_14592,N_11014,N_9263);
nand U14593 (N_14593,N_9439,N_9492);
or U14594 (N_14594,N_11166,N_10414);
and U14595 (N_14595,N_11688,N_9275);
and U14596 (N_14596,N_10196,N_10251);
nand U14597 (N_14597,N_9654,N_10851);
or U14598 (N_14598,N_10597,N_9330);
nand U14599 (N_14599,N_10898,N_11947);
or U14600 (N_14600,N_10670,N_11741);
or U14601 (N_14601,N_10629,N_10541);
or U14602 (N_14602,N_11074,N_10288);
nor U14603 (N_14603,N_11969,N_11366);
nor U14604 (N_14604,N_11778,N_9232);
nor U14605 (N_14605,N_10877,N_10087);
or U14606 (N_14606,N_9134,N_9446);
nor U14607 (N_14607,N_9881,N_9664);
and U14608 (N_14608,N_10018,N_9268);
or U14609 (N_14609,N_9678,N_11990);
or U14610 (N_14610,N_9929,N_9413);
and U14611 (N_14611,N_10268,N_11874);
nand U14612 (N_14612,N_10659,N_9384);
nand U14613 (N_14613,N_10554,N_9710);
and U14614 (N_14614,N_11311,N_11552);
nor U14615 (N_14615,N_10502,N_11844);
or U14616 (N_14616,N_10096,N_9237);
or U14617 (N_14617,N_11452,N_11678);
or U14618 (N_14618,N_10662,N_10713);
and U14619 (N_14619,N_11476,N_9689);
or U14620 (N_14620,N_10585,N_10094);
and U14621 (N_14621,N_9405,N_11390);
nand U14622 (N_14622,N_10274,N_10231);
or U14623 (N_14623,N_11292,N_10322);
and U14624 (N_14624,N_9426,N_11787);
nor U14625 (N_14625,N_9113,N_9072);
or U14626 (N_14626,N_9099,N_9885);
and U14627 (N_14627,N_9184,N_9699);
nand U14628 (N_14628,N_9754,N_9173);
or U14629 (N_14629,N_10925,N_11294);
nor U14630 (N_14630,N_11520,N_10725);
nor U14631 (N_14631,N_11677,N_10040);
or U14632 (N_14632,N_9685,N_10941);
nor U14633 (N_14633,N_11710,N_10491);
nand U14634 (N_14634,N_9117,N_11398);
nor U14635 (N_14635,N_11927,N_11306);
or U14636 (N_14636,N_10533,N_9828);
or U14637 (N_14637,N_9351,N_11899);
nand U14638 (N_14638,N_9854,N_10662);
nor U14639 (N_14639,N_10340,N_9767);
nand U14640 (N_14640,N_9305,N_11835);
and U14641 (N_14641,N_9027,N_11719);
and U14642 (N_14642,N_10381,N_9292);
nand U14643 (N_14643,N_9773,N_9262);
or U14644 (N_14644,N_9188,N_11805);
and U14645 (N_14645,N_11587,N_10984);
or U14646 (N_14646,N_10610,N_10401);
nor U14647 (N_14647,N_11551,N_9538);
or U14648 (N_14648,N_9417,N_10510);
and U14649 (N_14649,N_11212,N_11871);
and U14650 (N_14650,N_9897,N_11455);
and U14651 (N_14651,N_9212,N_11540);
nor U14652 (N_14652,N_9868,N_9752);
or U14653 (N_14653,N_9630,N_9935);
nor U14654 (N_14654,N_9459,N_9724);
nand U14655 (N_14655,N_10445,N_11426);
nand U14656 (N_14656,N_11937,N_9525);
nand U14657 (N_14657,N_10064,N_10140);
or U14658 (N_14658,N_9191,N_11153);
nand U14659 (N_14659,N_9985,N_10577);
nand U14660 (N_14660,N_11288,N_10934);
or U14661 (N_14661,N_9295,N_11783);
or U14662 (N_14662,N_10216,N_11469);
nand U14663 (N_14663,N_9244,N_9401);
or U14664 (N_14664,N_11227,N_9928);
or U14665 (N_14665,N_10396,N_10816);
nand U14666 (N_14666,N_9438,N_9306);
and U14667 (N_14667,N_11435,N_9725);
nor U14668 (N_14668,N_11412,N_9407);
and U14669 (N_14669,N_10307,N_10326);
nor U14670 (N_14670,N_9916,N_11308);
nand U14671 (N_14671,N_9149,N_10796);
or U14672 (N_14672,N_11319,N_10546);
and U14673 (N_14673,N_11025,N_10700);
nand U14674 (N_14674,N_10446,N_10835);
nor U14675 (N_14675,N_9704,N_9314);
and U14676 (N_14676,N_11763,N_11174);
nand U14677 (N_14677,N_11343,N_9796);
nand U14678 (N_14678,N_11156,N_11393);
or U14679 (N_14679,N_9146,N_10271);
nor U14680 (N_14680,N_9687,N_9554);
or U14681 (N_14681,N_9428,N_10655);
nand U14682 (N_14682,N_9530,N_10044);
nor U14683 (N_14683,N_9276,N_11911);
nand U14684 (N_14684,N_9040,N_10369);
or U14685 (N_14685,N_10190,N_10613);
and U14686 (N_14686,N_9285,N_9595);
nand U14687 (N_14687,N_11049,N_9000);
nor U14688 (N_14688,N_11638,N_10523);
nand U14689 (N_14689,N_10274,N_9539);
nor U14690 (N_14690,N_10775,N_9393);
nor U14691 (N_14691,N_10599,N_10150);
nor U14692 (N_14692,N_9070,N_10874);
or U14693 (N_14693,N_9344,N_9777);
nand U14694 (N_14694,N_10327,N_11352);
nand U14695 (N_14695,N_10896,N_11529);
nand U14696 (N_14696,N_10860,N_9623);
nand U14697 (N_14697,N_11280,N_9062);
and U14698 (N_14698,N_9420,N_9660);
and U14699 (N_14699,N_11109,N_10189);
or U14700 (N_14700,N_10881,N_11125);
nand U14701 (N_14701,N_11453,N_11612);
and U14702 (N_14702,N_9577,N_9578);
nand U14703 (N_14703,N_10005,N_11886);
nand U14704 (N_14704,N_9175,N_10566);
and U14705 (N_14705,N_11704,N_11387);
or U14706 (N_14706,N_10378,N_9880);
and U14707 (N_14707,N_10909,N_9651);
or U14708 (N_14708,N_9399,N_9279);
or U14709 (N_14709,N_9950,N_9123);
and U14710 (N_14710,N_9284,N_9469);
nand U14711 (N_14711,N_9138,N_9622);
nor U14712 (N_14712,N_10663,N_9171);
nand U14713 (N_14713,N_9584,N_10469);
and U14714 (N_14714,N_9972,N_9356);
or U14715 (N_14715,N_9242,N_9147);
or U14716 (N_14716,N_9133,N_9331);
nor U14717 (N_14717,N_11227,N_11777);
nor U14718 (N_14718,N_10035,N_11341);
nand U14719 (N_14719,N_9518,N_10452);
or U14720 (N_14720,N_10074,N_9253);
nor U14721 (N_14721,N_10156,N_11659);
or U14722 (N_14722,N_9778,N_9107);
or U14723 (N_14723,N_11408,N_9806);
nor U14724 (N_14724,N_11341,N_10812);
nand U14725 (N_14725,N_10873,N_11067);
and U14726 (N_14726,N_10213,N_10347);
xor U14727 (N_14727,N_11234,N_11885);
nand U14728 (N_14728,N_10536,N_10044);
and U14729 (N_14729,N_11468,N_10453);
and U14730 (N_14730,N_11357,N_10308);
or U14731 (N_14731,N_9120,N_11853);
or U14732 (N_14732,N_9981,N_11472);
nor U14733 (N_14733,N_11192,N_10999);
nor U14734 (N_14734,N_11377,N_10621);
and U14735 (N_14735,N_11991,N_10810);
nand U14736 (N_14736,N_11637,N_11260);
nand U14737 (N_14737,N_11934,N_9335);
and U14738 (N_14738,N_9490,N_10922);
nand U14739 (N_14739,N_11724,N_10633);
nor U14740 (N_14740,N_10732,N_9135);
and U14741 (N_14741,N_9198,N_10966);
and U14742 (N_14742,N_10717,N_10540);
nor U14743 (N_14743,N_11516,N_10279);
and U14744 (N_14744,N_9666,N_11164);
or U14745 (N_14745,N_9119,N_11706);
or U14746 (N_14746,N_9983,N_9135);
nand U14747 (N_14747,N_9084,N_11904);
nor U14748 (N_14748,N_11157,N_10741);
or U14749 (N_14749,N_11557,N_9932);
nand U14750 (N_14750,N_9620,N_9853);
or U14751 (N_14751,N_11890,N_9120);
nand U14752 (N_14752,N_11984,N_10460);
or U14753 (N_14753,N_10499,N_9188);
or U14754 (N_14754,N_10060,N_10558);
nor U14755 (N_14755,N_11633,N_11445);
or U14756 (N_14756,N_10601,N_10656);
nand U14757 (N_14757,N_10369,N_11895);
nor U14758 (N_14758,N_10572,N_11881);
and U14759 (N_14759,N_9304,N_11393);
and U14760 (N_14760,N_9746,N_11590);
and U14761 (N_14761,N_10066,N_9790);
nor U14762 (N_14762,N_11230,N_11515);
nor U14763 (N_14763,N_10414,N_11539);
or U14764 (N_14764,N_11093,N_11710);
or U14765 (N_14765,N_9631,N_11518);
nor U14766 (N_14766,N_11619,N_9253);
or U14767 (N_14767,N_9360,N_10427);
nor U14768 (N_14768,N_11923,N_9122);
or U14769 (N_14769,N_10586,N_11491);
or U14770 (N_14770,N_9450,N_11573);
and U14771 (N_14771,N_10845,N_11766);
and U14772 (N_14772,N_11972,N_9333);
and U14773 (N_14773,N_11216,N_11276);
and U14774 (N_14774,N_9886,N_10079);
or U14775 (N_14775,N_10936,N_9746);
and U14776 (N_14776,N_11113,N_10294);
or U14777 (N_14777,N_9797,N_10098);
nand U14778 (N_14778,N_9696,N_11056);
nor U14779 (N_14779,N_11744,N_10469);
nor U14780 (N_14780,N_10832,N_9929);
nand U14781 (N_14781,N_10992,N_10281);
nand U14782 (N_14782,N_9005,N_9290);
nand U14783 (N_14783,N_11989,N_9910);
nand U14784 (N_14784,N_10859,N_10808);
nor U14785 (N_14785,N_10992,N_11350);
nor U14786 (N_14786,N_10877,N_10875);
or U14787 (N_14787,N_10152,N_10965);
and U14788 (N_14788,N_10977,N_11367);
or U14789 (N_14789,N_9954,N_9384);
or U14790 (N_14790,N_10747,N_9958);
or U14791 (N_14791,N_11822,N_10199);
nand U14792 (N_14792,N_11224,N_9633);
nand U14793 (N_14793,N_11806,N_11290);
nor U14794 (N_14794,N_10047,N_10874);
and U14795 (N_14795,N_11860,N_11078);
and U14796 (N_14796,N_10184,N_11011);
nor U14797 (N_14797,N_11925,N_11721);
or U14798 (N_14798,N_9368,N_9006);
nor U14799 (N_14799,N_9369,N_9785);
nand U14800 (N_14800,N_9690,N_9828);
nand U14801 (N_14801,N_9316,N_11251);
nand U14802 (N_14802,N_9606,N_9847);
nand U14803 (N_14803,N_10612,N_10290);
or U14804 (N_14804,N_10440,N_10978);
nor U14805 (N_14805,N_10116,N_9102);
nand U14806 (N_14806,N_11874,N_11511);
or U14807 (N_14807,N_9991,N_9805);
nand U14808 (N_14808,N_11221,N_11161);
nand U14809 (N_14809,N_11555,N_10146);
and U14810 (N_14810,N_11816,N_10887);
nand U14811 (N_14811,N_11410,N_11926);
nor U14812 (N_14812,N_9300,N_9460);
nand U14813 (N_14813,N_10591,N_9375);
or U14814 (N_14814,N_9555,N_10958);
nor U14815 (N_14815,N_11208,N_9928);
nor U14816 (N_14816,N_10552,N_9689);
nor U14817 (N_14817,N_9587,N_10330);
nand U14818 (N_14818,N_9171,N_10401);
nor U14819 (N_14819,N_9633,N_11419);
nor U14820 (N_14820,N_11116,N_11497);
or U14821 (N_14821,N_10669,N_9020);
and U14822 (N_14822,N_9626,N_10586);
nor U14823 (N_14823,N_10786,N_10756);
nand U14824 (N_14824,N_9924,N_11759);
and U14825 (N_14825,N_9522,N_9447);
nand U14826 (N_14826,N_11525,N_11749);
nor U14827 (N_14827,N_9579,N_11037);
and U14828 (N_14828,N_9986,N_10980);
nand U14829 (N_14829,N_11014,N_11111);
or U14830 (N_14830,N_11319,N_9890);
nor U14831 (N_14831,N_10244,N_10500);
nand U14832 (N_14832,N_11049,N_9051);
nand U14833 (N_14833,N_10855,N_9743);
or U14834 (N_14834,N_9159,N_11799);
nor U14835 (N_14835,N_10544,N_11936);
nor U14836 (N_14836,N_9860,N_11841);
nor U14837 (N_14837,N_10521,N_9645);
nor U14838 (N_14838,N_10182,N_11917);
or U14839 (N_14839,N_11178,N_11927);
or U14840 (N_14840,N_9914,N_11855);
nor U14841 (N_14841,N_9589,N_9088);
and U14842 (N_14842,N_11849,N_11035);
nor U14843 (N_14843,N_9131,N_9688);
and U14844 (N_14844,N_9615,N_9812);
or U14845 (N_14845,N_11739,N_9094);
nand U14846 (N_14846,N_9189,N_9618);
and U14847 (N_14847,N_10137,N_9060);
or U14848 (N_14848,N_11529,N_9561);
nand U14849 (N_14849,N_10709,N_11186);
or U14850 (N_14850,N_11996,N_9730);
and U14851 (N_14851,N_10646,N_11583);
nand U14852 (N_14852,N_11239,N_11228);
nor U14853 (N_14853,N_10268,N_9273);
nand U14854 (N_14854,N_9764,N_11070);
and U14855 (N_14855,N_11893,N_9307);
nand U14856 (N_14856,N_9965,N_11382);
and U14857 (N_14857,N_11879,N_11951);
and U14858 (N_14858,N_9183,N_9957);
nor U14859 (N_14859,N_10691,N_10215);
or U14860 (N_14860,N_11072,N_11257);
nand U14861 (N_14861,N_10414,N_11798);
or U14862 (N_14862,N_11350,N_11844);
xnor U14863 (N_14863,N_11451,N_11019);
or U14864 (N_14864,N_10607,N_10609);
and U14865 (N_14865,N_9493,N_9020);
or U14866 (N_14866,N_10273,N_10783);
or U14867 (N_14867,N_11101,N_11684);
or U14868 (N_14868,N_10294,N_10783);
nor U14869 (N_14869,N_11397,N_11596);
nor U14870 (N_14870,N_9394,N_11102);
or U14871 (N_14871,N_11446,N_11953);
nand U14872 (N_14872,N_10100,N_11366);
or U14873 (N_14873,N_11884,N_10898);
nand U14874 (N_14874,N_9649,N_11998);
nand U14875 (N_14875,N_11614,N_11851);
or U14876 (N_14876,N_9071,N_10281);
and U14877 (N_14877,N_10175,N_11935);
nand U14878 (N_14878,N_9989,N_11437);
nand U14879 (N_14879,N_11927,N_10239);
nor U14880 (N_14880,N_11166,N_10007);
or U14881 (N_14881,N_9244,N_11832);
nor U14882 (N_14882,N_9448,N_11763);
or U14883 (N_14883,N_9105,N_9397);
nand U14884 (N_14884,N_10916,N_9364);
or U14885 (N_14885,N_10776,N_11342);
or U14886 (N_14886,N_10567,N_11851);
nand U14887 (N_14887,N_10896,N_11920);
nand U14888 (N_14888,N_9309,N_11110);
nor U14889 (N_14889,N_10121,N_10225);
and U14890 (N_14890,N_9771,N_10754);
and U14891 (N_14891,N_11935,N_9919);
nand U14892 (N_14892,N_11669,N_9195);
nor U14893 (N_14893,N_9482,N_10259);
nor U14894 (N_14894,N_9077,N_11845);
nor U14895 (N_14895,N_11682,N_9837);
nand U14896 (N_14896,N_11769,N_10859);
and U14897 (N_14897,N_11173,N_11881);
nand U14898 (N_14898,N_10687,N_11086);
or U14899 (N_14899,N_11100,N_9379);
and U14900 (N_14900,N_9184,N_10575);
or U14901 (N_14901,N_10290,N_9789);
nor U14902 (N_14902,N_11844,N_11518);
and U14903 (N_14903,N_9833,N_11778);
nand U14904 (N_14904,N_11558,N_9750);
and U14905 (N_14905,N_11521,N_9724);
and U14906 (N_14906,N_9283,N_11305);
and U14907 (N_14907,N_9236,N_10692);
and U14908 (N_14908,N_10728,N_11770);
nand U14909 (N_14909,N_11078,N_9357);
and U14910 (N_14910,N_9653,N_10938);
nand U14911 (N_14911,N_9768,N_9879);
and U14912 (N_14912,N_9182,N_11224);
nor U14913 (N_14913,N_9497,N_9817);
and U14914 (N_14914,N_11434,N_9304);
and U14915 (N_14915,N_11060,N_9419);
nor U14916 (N_14916,N_10077,N_9865);
xor U14917 (N_14917,N_10244,N_10465);
nor U14918 (N_14918,N_10409,N_11351);
or U14919 (N_14919,N_9206,N_10435);
nand U14920 (N_14920,N_9740,N_11058);
nand U14921 (N_14921,N_9206,N_10452);
or U14922 (N_14922,N_11559,N_11727);
nor U14923 (N_14923,N_11788,N_9509);
or U14924 (N_14924,N_10044,N_9927);
nor U14925 (N_14925,N_11625,N_11655);
nor U14926 (N_14926,N_10327,N_10771);
and U14927 (N_14927,N_9620,N_10505);
nor U14928 (N_14928,N_10623,N_9095);
or U14929 (N_14929,N_11880,N_11349);
and U14930 (N_14930,N_11091,N_11858);
or U14931 (N_14931,N_11004,N_9365);
or U14932 (N_14932,N_10703,N_10032);
nor U14933 (N_14933,N_10823,N_9933);
nor U14934 (N_14934,N_11961,N_11829);
and U14935 (N_14935,N_11089,N_10065);
nor U14936 (N_14936,N_10401,N_10061);
nand U14937 (N_14937,N_9738,N_10733);
nand U14938 (N_14938,N_9942,N_10761);
and U14939 (N_14939,N_11046,N_11517);
or U14940 (N_14940,N_9710,N_9938);
nor U14941 (N_14941,N_10903,N_10210);
nand U14942 (N_14942,N_9276,N_10519);
and U14943 (N_14943,N_10557,N_10318);
and U14944 (N_14944,N_11779,N_9703);
nand U14945 (N_14945,N_9273,N_10166);
nor U14946 (N_14946,N_10413,N_9000);
nand U14947 (N_14947,N_10132,N_9529);
nor U14948 (N_14948,N_9611,N_11979);
nand U14949 (N_14949,N_9655,N_11333);
nor U14950 (N_14950,N_9656,N_10841);
xor U14951 (N_14951,N_9092,N_9143);
or U14952 (N_14952,N_10676,N_11798);
and U14953 (N_14953,N_9722,N_9940);
or U14954 (N_14954,N_9498,N_10514);
or U14955 (N_14955,N_10439,N_11215);
nor U14956 (N_14956,N_10330,N_9288);
nand U14957 (N_14957,N_9732,N_11230);
or U14958 (N_14958,N_11224,N_10223);
and U14959 (N_14959,N_11547,N_11961);
or U14960 (N_14960,N_10191,N_10202);
or U14961 (N_14961,N_9894,N_9563);
or U14962 (N_14962,N_11510,N_10878);
nor U14963 (N_14963,N_11812,N_10965);
nor U14964 (N_14964,N_11295,N_9490);
nand U14965 (N_14965,N_9156,N_10483);
and U14966 (N_14966,N_10419,N_11485);
nand U14967 (N_14967,N_11124,N_10283);
nor U14968 (N_14968,N_10901,N_11440);
or U14969 (N_14969,N_9347,N_11256);
and U14970 (N_14970,N_9550,N_10507);
and U14971 (N_14971,N_10887,N_10809);
and U14972 (N_14972,N_9673,N_10964);
nand U14973 (N_14973,N_10397,N_11952);
and U14974 (N_14974,N_11092,N_9958);
and U14975 (N_14975,N_10116,N_11433);
nand U14976 (N_14976,N_11709,N_11786);
nand U14977 (N_14977,N_9401,N_10909);
and U14978 (N_14978,N_11531,N_11773);
nor U14979 (N_14979,N_11011,N_10967);
or U14980 (N_14980,N_11572,N_11584);
nand U14981 (N_14981,N_11131,N_11542);
or U14982 (N_14982,N_11570,N_10274);
nand U14983 (N_14983,N_9886,N_11714);
nand U14984 (N_14984,N_10945,N_9460);
or U14985 (N_14985,N_10797,N_10053);
and U14986 (N_14986,N_10003,N_9781);
nor U14987 (N_14987,N_11319,N_11052);
and U14988 (N_14988,N_10573,N_10381);
and U14989 (N_14989,N_11388,N_10224);
nor U14990 (N_14990,N_11660,N_9150);
and U14991 (N_14991,N_9040,N_9746);
and U14992 (N_14992,N_11900,N_9941);
nor U14993 (N_14993,N_11339,N_9997);
or U14994 (N_14994,N_11675,N_11370);
nor U14995 (N_14995,N_9141,N_11777);
or U14996 (N_14996,N_10161,N_11609);
or U14997 (N_14997,N_9125,N_11487);
or U14998 (N_14998,N_11289,N_11154);
nand U14999 (N_14999,N_9308,N_11863);
or UO_0 (O_0,N_13674,N_14943);
nand UO_1 (O_1,N_12491,N_14355);
or UO_2 (O_2,N_13506,N_12099);
or UO_3 (O_3,N_13352,N_12480);
and UO_4 (O_4,N_14541,N_13291);
nor UO_5 (O_5,N_13272,N_13246);
nand UO_6 (O_6,N_13009,N_13648);
nor UO_7 (O_7,N_12202,N_12544);
and UO_8 (O_8,N_12590,N_13657);
nand UO_9 (O_9,N_12335,N_14117);
and UO_10 (O_10,N_13961,N_12736);
or UO_11 (O_11,N_12145,N_14999);
nor UO_12 (O_12,N_12820,N_13090);
nand UO_13 (O_13,N_13614,N_12259);
nor UO_14 (O_14,N_13882,N_14214);
nand UO_15 (O_15,N_12541,N_13076);
and UO_16 (O_16,N_12756,N_14816);
or UO_17 (O_17,N_13640,N_12630);
nand UO_18 (O_18,N_14538,N_13954);
nand UO_19 (O_19,N_13692,N_13239);
nand UO_20 (O_20,N_14930,N_13575);
nand UO_21 (O_21,N_13566,N_13758);
nor UO_22 (O_22,N_14623,N_14162);
nand UO_23 (O_23,N_13974,N_14661);
nor UO_24 (O_24,N_14451,N_14577);
or UO_25 (O_25,N_14842,N_12050);
and UO_26 (O_26,N_14555,N_13788);
and UO_27 (O_27,N_13417,N_14205);
or UO_28 (O_28,N_14585,N_14487);
or UO_29 (O_29,N_13008,N_14685);
and UO_30 (O_30,N_13512,N_14649);
nand UO_31 (O_31,N_14225,N_13485);
xor UO_32 (O_32,N_12812,N_12941);
or UO_33 (O_33,N_13162,N_12871);
nand UO_34 (O_34,N_13848,N_12723);
nand UO_35 (O_35,N_14591,N_13341);
nor UO_36 (O_36,N_14892,N_12126);
and UO_37 (O_37,N_13313,N_12218);
and UO_38 (O_38,N_12320,N_13918);
and UO_39 (O_39,N_14228,N_14596);
or UO_40 (O_40,N_13333,N_14310);
and UO_41 (O_41,N_13311,N_14366);
or UO_42 (O_42,N_14875,N_13589);
and UO_43 (O_43,N_14396,N_12978);
or UO_44 (O_44,N_14951,N_13188);
or UO_45 (O_45,N_12311,N_14250);
or UO_46 (O_46,N_12584,N_14037);
nor UO_47 (O_47,N_12471,N_12787);
and UO_48 (O_48,N_12850,N_14804);
and UO_49 (O_49,N_14893,N_13693);
or UO_50 (O_50,N_14710,N_12483);
nor UO_51 (O_51,N_13550,N_12332);
or UO_52 (O_52,N_14747,N_12389);
or UO_53 (O_53,N_14391,N_12806);
and UO_54 (O_54,N_12344,N_14189);
nand UO_55 (O_55,N_14243,N_14144);
or UO_56 (O_56,N_14836,N_14786);
nor UO_57 (O_57,N_14473,N_13937);
and UO_58 (O_58,N_12498,N_13583);
or UO_59 (O_59,N_13347,N_12041);
nor UO_60 (O_60,N_12447,N_14696);
nor UO_61 (O_61,N_14978,N_12010);
nor UO_62 (O_62,N_13077,N_13426);
nor UO_63 (O_63,N_14177,N_13178);
or UO_64 (O_64,N_12229,N_13018);
and UO_65 (O_65,N_12959,N_14447);
nor UO_66 (O_66,N_14480,N_14894);
nand UO_67 (O_67,N_13653,N_12148);
and UO_68 (O_68,N_12310,N_14635);
nor UO_69 (O_69,N_12980,N_13325);
nand UO_70 (O_70,N_13254,N_13711);
nor UO_71 (O_71,N_12465,N_14304);
or UO_72 (O_72,N_13547,N_13398);
or UO_73 (O_73,N_13295,N_14515);
or UO_74 (O_74,N_14292,N_14476);
and UO_75 (O_75,N_12095,N_12932);
nor UO_76 (O_76,N_12230,N_14756);
xnor UO_77 (O_77,N_13897,N_13115);
nor UO_78 (O_78,N_12263,N_13414);
nand UO_79 (O_79,N_12937,N_12645);
nor UO_80 (O_80,N_13628,N_12221);
nor UO_81 (O_81,N_13348,N_14377);
nand UO_82 (O_82,N_13487,N_14899);
and UO_83 (O_83,N_12857,N_12494);
or UO_84 (O_84,N_12060,N_13292);
nand UO_85 (O_85,N_12464,N_13855);
nand UO_86 (O_86,N_14173,N_14539);
and UO_87 (O_87,N_13905,N_12690);
or UO_88 (O_88,N_12697,N_12324);
nor UO_89 (O_89,N_14149,N_13817);
nor UO_90 (O_90,N_14618,N_12983);
nor UO_91 (O_91,N_14622,N_13962);
nor UO_92 (O_92,N_14192,N_14021);
nand UO_93 (O_93,N_12552,N_13886);
nor UO_94 (O_94,N_14459,N_14524);
nand UO_95 (O_95,N_14518,N_12283);
nor UO_96 (O_96,N_13782,N_14468);
or UO_97 (O_97,N_14379,N_14837);
and UO_98 (O_98,N_13564,N_13059);
nor UO_99 (O_99,N_14323,N_14204);
or UO_100 (O_100,N_12132,N_13609);
nor UO_101 (O_101,N_14221,N_13312);
nand UO_102 (O_102,N_14264,N_13057);
nand UO_103 (O_103,N_14267,N_14877);
or UO_104 (O_104,N_14483,N_13943);
nand UO_105 (O_105,N_12245,N_12386);
nand UO_106 (O_106,N_14062,N_12652);
nand UO_107 (O_107,N_12185,N_13148);
nor UO_108 (O_108,N_13630,N_14334);
nand UO_109 (O_109,N_14599,N_12451);
nand UO_110 (O_110,N_14509,N_14651);
nor UO_111 (O_111,N_14983,N_14805);
and UO_112 (O_112,N_13119,N_12052);
and UO_113 (O_113,N_13919,N_12873);
or UO_114 (O_114,N_12056,N_12891);
and UO_115 (O_115,N_13761,N_12747);
or UO_116 (O_116,N_14911,N_14799);
nor UO_117 (O_117,N_12639,N_13404);
and UO_118 (O_118,N_13125,N_14779);
nand UO_119 (O_119,N_14519,N_14111);
or UO_120 (O_120,N_14248,N_13756);
nor UO_121 (O_121,N_12623,N_12591);
and UO_122 (O_122,N_13532,N_13324);
and UO_123 (O_123,N_12362,N_12199);
nand UO_124 (O_124,N_12121,N_12053);
or UO_125 (O_125,N_12281,N_13040);
nand UO_126 (O_126,N_13032,N_13314);
or UO_127 (O_127,N_13807,N_14640);
nor UO_128 (O_128,N_14421,N_13000);
nand UO_129 (O_129,N_12034,N_13196);
nand UO_130 (O_130,N_12187,N_13748);
and UO_131 (O_131,N_14941,N_13351);
nand UO_132 (O_132,N_13738,N_13278);
nor UO_133 (O_133,N_13770,N_13821);
nor UO_134 (O_134,N_14234,N_14147);
nor UO_135 (O_135,N_13864,N_12602);
nand UO_136 (O_136,N_14545,N_14878);
xor UO_137 (O_137,N_12843,N_14426);
or UO_138 (O_138,N_12910,N_13004);
and UO_139 (O_139,N_14005,N_12967);
nor UO_140 (O_140,N_13542,N_13481);
nand UO_141 (O_141,N_14505,N_13386);
or UO_142 (O_142,N_13934,N_14478);
nand UO_143 (O_143,N_14455,N_14571);
nand UO_144 (O_144,N_13830,N_12046);
nand UO_145 (O_145,N_13220,N_13422);
or UO_146 (O_146,N_13637,N_14565);
nand UO_147 (O_147,N_12385,N_14692);
nand UO_148 (O_148,N_13214,N_14226);
nor UO_149 (O_149,N_13752,N_14948);
nand UO_150 (O_150,N_13340,N_14689);
nand UO_151 (O_151,N_13277,N_13198);
and UO_152 (O_152,N_14868,N_13682);
nor UO_153 (O_153,N_12223,N_12742);
nor UO_154 (O_154,N_12558,N_12087);
nand UO_155 (O_155,N_13444,N_13973);
nand UO_156 (O_156,N_12249,N_13730);
or UO_157 (O_157,N_14262,N_13517);
or UO_158 (O_158,N_14360,N_14423);
nand UO_159 (O_159,N_12151,N_14265);
nand UO_160 (O_160,N_12650,N_12265);
or UO_161 (O_161,N_13755,N_12818);
and UO_162 (O_162,N_12592,N_12213);
and UO_163 (O_163,N_14070,N_12696);
nor UO_164 (O_164,N_13852,N_13020);
nand UO_165 (O_165,N_13661,N_14564);
or UO_166 (O_166,N_13559,N_12196);
nor UO_167 (O_167,N_14903,N_12674);
nor UO_168 (O_168,N_13979,N_13816);
and UO_169 (O_169,N_12603,N_12015);
nor UO_170 (O_170,N_14726,N_14767);
and UO_171 (O_171,N_14164,N_14354);
nand UO_172 (O_172,N_13228,N_13306);
xor UO_173 (O_173,N_13364,N_13010);
nand UO_174 (O_174,N_13229,N_13380);
and UO_175 (O_175,N_12952,N_14628);
or UO_176 (O_176,N_12047,N_12036);
or UO_177 (O_177,N_12627,N_12319);
or UO_178 (O_178,N_12641,N_14503);
and UO_179 (O_179,N_14722,N_12734);
and UO_180 (O_180,N_14974,N_12503);
nand UO_181 (O_181,N_12380,N_13871);
or UO_182 (O_182,N_13709,N_13649);
and UO_183 (O_183,N_14866,N_13528);
and UO_184 (O_184,N_13405,N_14751);
nand UO_185 (O_185,N_13971,N_13486);
nor UO_186 (O_186,N_12981,N_14074);
and UO_187 (O_187,N_14975,N_13579);
and UO_188 (O_188,N_14888,N_14938);
nand UO_189 (O_189,N_12653,N_12642);
and UO_190 (O_190,N_12505,N_12051);
nor UO_191 (O_191,N_13688,N_14873);
nand UO_192 (O_192,N_14363,N_14150);
nor UO_193 (O_193,N_14073,N_13136);
nor UO_194 (O_194,N_12574,N_12525);
nor UO_195 (O_195,N_12414,N_12453);
or UO_196 (O_196,N_12877,N_12326);
nand UO_197 (O_197,N_14067,N_14184);
and UO_198 (O_198,N_12330,N_12212);
xnor UO_199 (O_199,N_12150,N_13146);
nor UO_200 (O_200,N_12802,N_14011);
and UO_201 (O_201,N_13491,N_13420);
and UO_202 (O_202,N_13387,N_14869);
or UO_203 (O_203,N_12179,N_13636);
nand UO_204 (O_204,N_14122,N_13765);
or UO_205 (O_205,N_14012,N_12821);
nor UO_206 (O_206,N_14403,N_14382);
nand UO_207 (O_207,N_13014,N_14966);
or UO_208 (O_208,N_13379,N_13207);
nand UO_209 (O_209,N_13870,N_13923);
and UO_210 (O_210,N_14321,N_13015);
or UO_211 (O_211,N_13732,N_12387);
nand UO_212 (O_212,N_14950,N_12322);
or UO_213 (O_213,N_14100,N_13194);
and UO_214 (O_214,N_13247,N_12800);
nand UO_215 (O_215,N_14492,N_13642);
nor UO_216 (O_216,N_12501,N_12700);
nand UO_217 (O_217,N_12101,N_14093);
or UO_218 (O_218,N_13519,N_13192);
or UO_219 (O_219,N_12692,N_13052);
and UO_220 (O_220,N_12103,N_14064);
and UO_221 (O_221,N_14914,N_12296);
and UO_222 (O_222,N_12137,N_13223);
or UO_223 (O_223,N_14477,N_13986);
nor UO_224 (O_224,N_12106,N_12731);
and UO_225 (O_225,N_13633,N_12794);
and UO_226 (O_226,N_13382,N_13159);
nor UO_227 (O_227,N_12452,N_14879);
and UO_228 (O_228,N_14116,N_14984);
and UO_229 (O_229,N_12360,N_13660);
nand UO_230 (O_230,N_14004,N_14288);
and UO_231 (O_231,N_13970,N_14737);
and UO_232 (O_232,N_13153,N_13712);
and UO_233 (O_233,N_14048,N_12954);
and UO_234 (O_234,N_14527,N_13895);
or UO_235 (O_235,N_14934,N_14802);
or UO_236 (O_236,N_14757,N_14831);
or UO_237 (O_237,N_12805,N_12968);
nor UO_238 (O_238,N_13060,N_12303);
nand UO_239 (O_239,N_12032,N_13013);
or UO_240 (O_240,N_14569,N_14083);
nor UO_241 (O_241,N_12108,N_12394);
nor UO_242 (O_242,N_13687,N_14301);
nand UO_243 (O_243,N_14395,N_13110);
nand UO_244 (O_244,N_12404,N_12343);
and UO_245 (O_245,N_14128,N_14028);
nor UO_246 (O_246,N_13994,N_12169);
nand UO_247 (O_247,N_12001,N_12314);
and UO_248 (O_248,N_14674,N_13187);
or UO_249 (O_249,N_14715,N_14717);
nand UO_250 (O_250,N_12334,N_14929);
and UO_251 (O_251,N_14072,N_12781);
and UO_252 (O_252,N_13346,N_14643);
nand UO_253 (O_253,N_12699,N_13443);
or UO_254 (O_254,N_13476,N_12838);
nand UO_255 (O_255,N_13704,N_14650);
nor UO_256 (O_256,N_12206,N_12158);
xor UO_257 (O_257,N_13353,N_12091);
or UO_258 (O_258,N_13323,N_12811);
and UO_259 (O_259,N_13151,N_12716);
and UO_260 (O_260,N_14188,N_13588);
nand UO_261 (O_261,N_12675,N_14789);
or UO_262 (O_262,N_13473,N_14216);
and UO_263 (O_263,N_12258,N_14969);
and UO_264 (O_264,N_14792,N_12918);
or UO_265 (O_265,N_13553,N_14263);
nand UO_266 (O_266,N_12318,N_14820);
nor UO_267 (O_267,N_12765,N_13270);
nand UO_268 (O_268,N_14258,N_12061);
or UO_269 (O_269,N_12559,N_12301);
nand UO_270 (O_270,N_13315,N_12647);
and UO_271 (O_271,N_14326,N_14347);
nand UO_272 (O_272,N_12915,N_13061);
nand UO_273 (O_273,N_14876,N_12657);
nor UO_274 (O_274,N_13408,N_12356);
or UO_275 (O_275,N_12467,N_13879);
and UO_276 (O_276,N_14594,N_13964);
nor UO_277 (O_277,N_12474,N_14091);
nand UO_278 (O_278,N_13156,N_14573);
or UO_279 (O_279,N_12450,N_13740);
nor UO_280 (O_280,N_12615,N_13992);
and UO_281 (O_281,N_14972,N_12190);
or UO_282 (O_282,N_14719,N_13802);
nand UO_283 (O_283,N_14695,N_12928);
and UO_284 (O_284,N_13535,N_13812);
or UO_285 (O_285,N_13843,N_14931);
or UO_286 (O_286,N_12002,N_14271);
or UO_287 (O_287,N_13894,N_14810);
nor UO_288 (O_288,N_14644,N_14682);
or UO_289 (O_289,N_14819,N_14240);
or UO_290 (O_290,N_13577,N_12567);
and UO_291 (O_291,N_12998,N_12289);
nand UO_292 (O_292,N_14383,N_12807);
nor UO_293 (O_293,N_14551,N_12287);
or UO_294 (O_294,N_13349,N_12504);
nor UO_295 (O_295,N_12511,N_13784);
nand UO_296 (O_296,N_12867,N_12562);
or UO_297 (O_297,N_13624,N_12111);
nor UO_298 (O_298,N_14134,N_13217);
and UO_299 (O_299,N_14441,N_13157);
and UO_300 (O_300,N_13274,N_12291);
nor UO_301 (O_301,N_14801,N_12791);
nand UO_302 (O_302,N_13846,N_13936);
or UO_303 (O_303,N_13448,N_12810);
nand UO_304 (O_304,N_14336,N_13686);
nor UO_305 (O_305,N_13644,N_14154);
or UO_306 (O_306,N_12165,N_12507);
or UO_307 (O_307,N_13326,N_13212);
nor UO_308 (O_308,N_14203,N_14613);
nand UO_309 (O_309,N_14058,N_12996);
nand UO_310 (O_310,N_13470,N_12859);
and UO_311 (O_311,N_12814,N_12238);
nand UO_312 (O_312,N_14968,N_12144);
or UO_313 (O_313,N_14522,N_14198);
nand UO_314 (O_314,N_14105,N_14231);
nand UO_315 (O_315,N_14299,N_13521);
nor UO_316 (O_316,N_12823,N_13958);
nand UO_317 (O_317,N_12789,N_12671);
nor UO_318 (O_318,N_13534,N_12410);
nor UO_319 (O_319,N_12485,N_12921);
and UO_320 (O_320,N_12120,N_12746);
nand UO_321 (O_321,N_14475,N_12042);
and UO_322 (O_322,N_13423,N_13741);
and UO_323 (O_323,N_12920,N_13049);
or UO_324 (O_324,N_14716,N_13205);
or UO_325 (O_325,N_13318,N_12846);
and UO_326 (O_326,N_14328,N_12473);
or UO_327 (O_327,N_14595,N_13092);
nor UO_328 (O_328,N_13219,N_12232);
nand UO_329 (O_329,N_14699,N_13002);
and UO_330 (O_330,N_12225,N_13452);
and UO_331 (O_331,N_14735,N_13037);
nor UO_332 (O_332,N_14907,N_14706);
and UO_333 (O_333,N_14755,N_12149);
nor UO_334 (O_334,N_13445,N_12550);
or UO_335 (O_335,N_12929,N_13837);
or UO_336 (O_336,N_12182,N_13359);
xor UO_337 (O_337,N_14664,N_13541);
and UO_338 (O_338,N_12849,N_12134);
or UO_339 (O_339,N_13744,N_12673);
or UO_340 (O_340,N_12537,N_14843);
nand UO_341 (O_341,N_14976,N_13634);
nand UO_342 (O_342,N_14724,N_12497);
nor UO_343 (O_343,N_12569,N_13441);
and UO_344 (O_344,N_13289,N_13075);
nor UO_345 (O_345,N_12947,N_14761);
nand UO_346 (O_346,N_13823,N_14175);
and UO_347 (O_347,N_14940,N_14850);
or UO_348 (O_348,N_14729,N_13995);
nor UO_349 (O_349,N_14748,N_13027);
and UO_350 (O_350,N_13330,N_13658);
nor UO_351 (O_351,N_12622,N_14135);
and UO_352 (O_352,N_13902,N_12612);
and UO_353 (O_353,N_12830,N_12655);
or UO_354 (O_354,N_14927,N_14041);
nand UO_355 (O_355,N_13102,N_14762);
nor UO_356 (O_356,N_14163,N_12796);
or UO_357 (O_357,N_12531,N_13050);
or UO_358 (O_358,N_12896,N_14902);
nand UO_359 (O_359,N_13851,N_12914);
nor UO_360 (O_360,N_12009,N_14742);
and UO_361 (O_361,N_13952,N_13569);
nor UO_362 (O_362,N_13910,N_14935);
and UO_363 (O_363,N_12486,N_12455);
and UO_364 (O_364,N_13513,N_13045);
nor UO_365 (O_365,N_13753,N_14499);
and UO_366 (O_366,N_13388,N_13775);
nand UO_367 (O_367,N_14103,N_12012);
and UO_368 (O_368,N_12556,N_13610);
nor UO_369 (O_369,N_13173,N_13795);
or UO_370 (O_370,N_13561,N_12379);
and UO_371 (O_371,N_13597,N_14600);
nand UO_372 (O_372,N_13762,N_14647);
or UO_373 (O_373,N_14412,N_14331);
or UO_374 (O_374,N_14610,N_13727);
or UO_375 (O_375,N_12819,N_14732);
and UO_376 (O_376,N_14845,N_12676);
and UO_377 (O_377,N_12096,N_14559);
nor UO_378 (O_378,N_12092,N_13991);
nor UO_379 (O_379,N_14273,N_12934);
nand UO_380 (O_380,N_13337,N_14068);
nand UO_381 (O_381,N_12469,N_14152);
nand UO_382 (O_382,N_12155,N_14495);
nor UO_383 (O_383,N_14210,N_12542);
or UO_384 (O_384,N_14990,N_12248);
or UO_385 (O_385,N_12536,N_14882);
or UO_386 (O_386,N_12338,N_12286);
or UO_387 (O_387,N_14452,N_14227);
and UO_388 (O_388,N_13537,N_14094);
or UO_389 (O_389,N_12861,N_13258);
nor UO_390 (O_390,N_13455,N_14784);
or UO_391 (O_391,N_14708,N_14981);
nor UO_392 (O_392,N_12856,N_14809);
and UO_393 (O_393,N_14517,N_12191);
nor UO_394 (O_394,N_13477,N_14668);
nand UO_395 (O_395,N_14581,N_13708);
and UO_396 (O_396,N_12719,N_13342);
and UO_397 (O_397,N_13440,N_13372);
or UO_398 (O_398,N_14450,N_14329);
nor UO_399 (O_399,N_12840,N_12241);
or UO_400 (O_400,N_12817,N_13616);
xnor UO_401 (O_401,N_14392,N_12138);
nor UO_402 (O_402,N_12648,N_14218);
or UO_403 (O_403,N_13558,N_14686);
or UO_404 (O_404,N_12378,N_13665);
and UO_405 (O_405,N_12899,N_14159);
nand UO_406 (O_406,N_13336,N_13914);
or UO_407 (O_407,N_12424,N_12860);
and UO_408 (O_408,N_12757,N_13107);
nor UO_409 (O_409,N_13286,N_13948);
or UO_410 (O_410,N_13904,N_12917);
nor UO_411 (O_411,N_13276,N_14418);
nand UO_412 (O_412,N_13718,N_12304);
nor UO_413 (O_413,N_14707,N_12672);
nor UO_414 (O_414,N_14937,N_12236);
or UO_415 (O_415,N_13471,N_12837);
or UO_416 (O_416,N_13977,N_13063);
or UO_417 (O_417,N_12173,N_14180);
nand UO_418 (O_418,N_14349,N_14841);
or UO_419 (O_419,N_13393,N_13483);
nor UO_420 (O_420,N_12635,N_12530);
nand UO_421 (O_421,N_14324,N_12064);
and UO_422 (O_422,N_13983,N_12686);
or UO_423 (O_423,N_13800,N_13024);
nor UO_424 (O_424,N_12372,N_14241);
and UO_425 (O_425,N_12923,N_14325);
and UO_426 (O_426,N_13690,N_13585);
nand UO_427 (O_427,N_12195,N_13829);
or UO_428 (O_428,N_14659,N_14235);
or UO_429 (O_429,N_14992,N_14822);
nor UO_430 (O_430,N_12045,N_13316);
or UO_431 (O_431,N_12743,N_13850);
or UO_432 (O_432,N_12275,N_14358);
and UO_433 (O_433,N_14537,N_14018);
or UO_434 (O_434,N_12376,N_13881);
and UO_435 (O_435,N_13724,N_12116);
nand UO_436 (O_436,N_13472,N_14194);
or UO_437 (O_437,N_14985,N_12463);
and UO_438 (O_438,N_13960,N_14988);
nor UO_439 (O_439,N_14768,N_12509);
nor UO_440 (O_440,N_13493,N_13437);
nand UO_441 (O_441,N_12065,N_14007);
xnor UO_442 (O_442,N_13951,N_14445);
nand UO_443 (O_443,N_14634,N_14833);
nor UO_444 (O_444,N_13465,N_14115);
or UO_445 (O_445,N_13174,N_12626);
nor UO_446 (O_446,N_12377,N_12078);
nor UO_447 (O_447,N_12008,N_14533);
nand UO_448 (O_448,N_12684,N_14673);
nand UO_449 (O_449,N_12845,N_12433);
and UO_450 (O_450,N_12038,N_13363);
nand UO_451 (O_451,N_14467,N_12279);
or UO_452 (O_452,N_12862,N_13047);
nand UO_453 (O_453,N_12633,N_14614);
nand UO_454 (O_454,N_13384,N_14609);
nor UO_455 (O_455,N_13281,N_14220);
nor UO_456 (O_456,N_12588,N_14042);
and UO_457 (O_457,N_12661,N_12783);
nor UO_458 (O_458,N_14155,N_14080);
and UO_459 (O_459,N_12164,N_13236);
nand UO_460 (O_460,N_13912,N_13689);
or UO_461 (O_461,N_14142,N_12140);
nor UO_462 (O_462,N_14939,N_12637);
or UO_463 (O_463,N_12939,N_14570);
or UO_464 (O_464,N_12759,N_12348);
nand UO_465 (O_465,N_14964,N_14982);
or UO_466 (O_466,N_12839,N_12851);
nor UO_467 (O_467,N_14315,N_14587);
or UO_468 (O_468,N_13332,N_12381);
or UO_469 (O_469,N_14973,N_13197);
or UO_470 (O_470,N_13835,N_14044);
or UO_471 (O_471,N_12131,N_13831);
nor UO_472 (O_472,N_13164,N_13475);
or UO_473 (O_473,N_14705,N_14406);
nand UO_474 (O_474,N_13436,N_13053);
nor UO_475 (O_475,N_14463,N_14773);
nand UO_476 (O_476,N_13767,N_14031);
nor UO_477 (O_477,N_13834,N_12127);
nor UO_478 (O_478,N_12133,N_12461);
nor UO_479 (O_479,N_13369,N_12129);
and UO_480 (O_480,N_13591,N_14887);
nand UO_481 (O_481,N_12398,N_13048);
or UO_482 (O_482,N_14885,N_12014);
nand UO_483 (O_483,N_13376,N_13647);
and UO_484 (O_484,N_14608,N_14676);
and UO_485 (O_485,N_13154,N_14662);
nor UO_486 (O_486,N_12888,N_12748);
nor UO_487 (O_487,N_13457,N_14703);
and UO_488 (O_488,N_12429,N_13067);
and UO_489 (O_489,N_14631,N_12003);
and UO_490 (O_490,N_14464,N_13089);
or UO_491 (O_491,N_13428,N_14239);
or UO_492 (O_492,N_12539,N_12717);
nand UO_493 (O_493,N_14813,N_14840);
and UO_494 (O_494,N_14544,N_12880);
and UO_495 (O_495,N_14566,N_14925);
xnor UO_496 (O_496,N_12638,N_12048);
and UO_497 (O_497,N_12354,N_13916);
and UO_498 (O_498,N_13702,N_13651);
and UO_499 (O_499,N_14461,N_14909);
nand UO_500 (O_500,N_12395,N_14796);
nor UO_501 (O_501,N_12170,N_13251);
nand UO_502 (O_502,N_14855,N_13177);
nand UO_503 (O_503,N_14046,N_13509);
and UO_504 (O_504,N_13058,N_13294);
nor UO_505 (O_505,N_13006,N_14488);
nand UO_506 (O_506,N_13503,N_13134);
nand UO_507 (O_507,N_14772,N_13608);
and UO_508 (O_508,N_14167,N_13182);
or UO_509 (O_509,N_13999,N_13622);
nor UO_510 (O_510,N_14316,N_14484);
nor UO_511 (O_511,N_14723,N_14270);
and UO_512 (O_512,N_13580,N_14528);
nand UO_513 (O_513,N_13953,N_13287);
or UO_514 (O_514,N_13180,N_13238);
or UO_515 (O_515,N_13459,N_12262);
or UO_516 (O_516,N_13769,N_14327);
nor UO_517 (O_517,N_12079,N_14367);
nand UO_518 (O_518,N_14965,N_12244);
or UO_519 (O_519,N_12184,N_13105);
and UO_520 (O_520,N_13673,N_14874);
or UO_521 (O_521,N_14959,N_12271);
nand UO_522 (O_522,N_13005,N_13202);
nor UO_523 (O_523,N_12957,N_12487);
or UO_524 (O_524,N_12445,N_14771);
nor UO_525 (O_525,N_12411,N_13853);
nor UO_526 (O_526,N_13504,N_14118);
nand UO_527 (O_527,N_14320,N_14025);
and UO_528 (O_528,N_14385,N_13989);
nand UO_529 (O_529,N_14800,N_12436);
and UO_530 (O_530,N_14141,N_14407);
nor UO_531 (O_531,N_14257,N_13915);
and UO_532 (O_532,N_14602,N_14371);
and UO_533 (O_533,N_12586,N_12906);
and UO_534 (O_534,N_12720,N_12976);
nand UO_535 (O_535,N_14454,N_14979);
nor UO_536 (O_536,N_12142,N_12701);
and UO_537 (O_537,N_12895,N_12526);
nor UO_538 (O_538,N_14408,N_12161);
nor UO_539 (O_539,N_13355,N_14290);
or UO_540 (O_540,N_13362,N_13681);
nand UO_541 (O_541,N_14898,N_13584);
or UO_542 (O_542,N_12347,N_14224);
nand UO_543 (O_543,N_14991,N_12023);
and UO_544 (O_544,N_14886,N_12912);
nor UO_545 (O_545,N_14658,N_12118);
or UO_546 (O_546,N_14795,N_12868);
nor UO_547 (O_547,N_14905,N_12919);
and UO_548 (O_548,N_13898,N_14714);
nor UO_549 (O_549,N_12446,N_12522);
nand UO_550 (O_550,N_12025,N_12349);
or UO_551 (O_551,N_13293,N_14828);
nor UO_552 (O_552,N_14711,N_12936);
or UO_553 (O_553,N_12993,N_13344);
nor UO_554 (O_554,N_13026,N_13920);
and UO_555 (O_555,N_13723,N_14867);
nor UO_556 (O_556,N_13250,N_13170);
and UO_557 (O_557,N_12767,N_12970);
and UO_558 (O_558,N_12844,N_13121);
or UO_559 (O_559,N_14680,N_13563);
or UO_560 (O_560,N_12237,N_12991);
nor UO_561 (O_561,N_12962,N_14924);
nand UO_562 (O_562,N_13189,N_14063);
or UO_563 (O_563,N_14607,N_12235);
nand UO_564 (O_564,N_13595,N_14169);
nand UO_565 (O_565,N_14009,N_12521);
and UO_566 (O_566,N_14656,N_12188);
and UO_567 (O_567,N_14921,N_12403);
nand UO_568 (O_568,N_13328,N_13001);
nor UO_569 (O_569,N_13370,N_14056);
and UO_570 (O_570,N_13145,N_14944);
and UO_571 (O_571,N_13734,N_13596);
and UO_572 (O_572,N_14540,N_14364);
nor UO_573 (O_573,N_12878,N_13749);
nand UO_574 (O_574,N_14549,N_13839);
or UO_575 (O_575,N_12135,N_14849);
nor UO_576 (O_576,N_12246,N_12081);
or UO_577 (O_577,N_13797,N_14276);
or UO_578 (O_578,N_13460,N_12088);
and UO_579 (O_579,N_12295,N_12508);
nand UO_580 (O_580,N_13976,N_12337);
and UO_581 (O_581,N_13210,N_13556);
and UO_582 (O_582,N_13413,N_14008);
nand UO_583 (O_583,N_14212,N_14444);
and UO_584 (O_584,N_14101,N_13260);
nor UO_585 (O_585,N_12328,N_12997);
and UO_586 (O_586,N_13516,N_14791);
nand UO_587 (O_587,N_13867,N_13906);
or UO_588 (O_588,N_14803,N_12217);
and UO_589 (O_589,N_12679,N_14342);
or UO_590 (O_590,N_12680,N_14770);
or UO_591 (O_591,N_14314,N_13434);
and UO_592 (O_592,N_14049,N_12327);
or UO_593 (O_593,N_12769,N_13482);
and UO_594 (O_594,N_13116,N_14397);
or UO_595 (O_595,N_12226,N_14201);
or UO_596 (O_596,N_13023,N_12890);
and UO_597 (O_597,N_12325,N_13334);
nand UO_598 (O_598,N_14351,N_12421);
nor UO_599 (O_599,N_12768,N_12512);
nand UO_600 (O_600,N_14808,N_13186);
and UO_601 (O_601,N_13451,N_13548);
and UO_602 (O_602,N_13683,N_12456);
nand UO_603 (O_603,N_14486,N_14287);
and UO_604 (O_604,N_12711,N_13827);
or UO_605 (O_605,N_13288,N_13957);
or UO_606 (O_606,N_13033,N_14330);
and UO_607 (O_607,N_13185,N_14994);
or UO_608 (O_608,N_14750,N_12829);
and UO_609 (O_609,N_12027,N_14121);
nand UO_610 (O_610,N_12488,N_14127);
or UO_611 (O_611,N_13523,N_14260);
nor UO_612 (O_612,N_14311,N_13456);
or UO_613 (O_613,N_14043,N_14576);
nor UO_614 (O_614,N_13367,N_14870);
or UO_615 (O_615,N_13847,N_12076);
xnor UO_616 (O_616,N_14977,N_14861);
or UO_617 (O_617,N_13621,N_13450);
nand UO_618 (O_618,N_14859,N_12028);
nand UO_619 (O_619,N_13766,N_14665);
nor UO_620 (O_620,N_13191,N_12267);
and UO_621 (O_621,N_13401,N_13003);
nand UO_622 (O_622,N_12585,N_12606);
and UO_623 (O_623,N_12822,N_12393);
nand UO_624 (O_624,N_14920,N_14466);
or UO_625 (O_625,N_12608,N_14589);
and UO_626 (O_626,N_12841,N_13932);
and UO_627 (O_627,N_12573,N_12677);
and UO_628 (O_628,N_12415,N_12468);
or UO_629 (O_629,N_13522,N_14047);
nand UO_630 (O_630,N_13038,N_12707);
and UO_631 (O_631,N_12181,N_13392);
nor UO_632 (O_632,N_13887,N_12798);
nand UO_633 (O_633,N_14436,N_13735);
or UO_634 (O_634,N_13086,N_12775);
and UO_635 (O_635,N_14642,N_12710);
nand UO_636 (O_636,N_14388,N_14233);
nand UO_637 (O_637,N_13298,N_14079);
nor UO_638 (O_638,N_14252,N_13375);
nand UO_639 (O_639,N_14333,N_13560);
nand UO_640 (O_640,N_13305,N_13271);
nor UO_641 (O_641,N_12884,N_14821);
or UO_642 (O_642,N_13412,N_14754);
nand UO_643 (O_643,N_14474,N_14278);
nor UO_644 (O_644,N_13232,N_12801);
nand UO_645 (O_645,N_14458,N_13252);
and UO_646 (O_646,N_14448,N_14120);
nor UO_647 (O_647,N_14023,N_13203);
nor UO_648 (O_648,N_13861,N_14738);
nor UO_649 (O_649,N_14123,N_14512);
nand UO_650 (O_650,N_14213,N_12624);
and UO_651 (O_651,N_13402,N_14880);
and UO_652 (O_652,N_12666,N_13435);
and UO_653 (O_653,N_14060,N_13750);
or UO_654 (O_654,N_14275,N_12578);
nand UO_655 (O_655,N_13468,N_12054);
or UO_656 (O_656,N_12546,N_12272);
nand UO_657 (O_657,N_14433,N_12909);
or UO_658 (O_658,N_14818,N_14255);
and UO_659 (O_659,N_14621,N_12345);
or UO_660 (O_660,N_14052,N_13317);
nor UO_661 (O_661,N_14730,N_12058);
or UO_662 (O_662,N_12203,N_12607);
nor UO_663 (O_663,N_13993,N_14432);
and UO_664 (O_664,N_12478,N_12724);
or UO_665 (O_665,N_14956,N_13743);
nand UO_666 (O_666,N_14394,N_12070);
nor UO_667 (O_667,N_13321,N_14462);
nor UO_668 (O_668,N_12373,N_14997);
nand UO_669 (O_669,N_13300,N_13619);
nand UO_670 (O_670,N_12869,N_14787);
nor UO_671 (O_671,N_13810,N_14743);
and UO_672 (O_672,N_12874,N_13803);
or UO_673 (O_673,N_12166,N_13171);
nor UO_674 (O_674,N_14908,N_12517);
nand UO_675 (O_675,N_14912,N_13406);
nand UO_676 (O_676,N_13731,N_13046);
nor UO_677 (O_677,N_13857,N_14918);
and UO_678 (O_678,N_13868,N_13464);
and UO_679 (O_679,N_14416,N_13892);
nand UO_680 (O_680,N_14217,N_14718);
nor UO_681 (O_681,N_12815,N_12293);
nand UO_682 (O_682,N_13618,N_13035);
nand UO_683 (O_683,N_12443,N_12006);
nor UO_684 (O_684,N_14497,N_12893);
and UO_685 (O_685,N_13011,N_14236);
or UO_686 (O_686,N_14017,N_14196);
and UO_687 (O_687,N_13433,N_13601);
and UO_688 (O_688,N_13890,N_13427);
and UO_689 (O_689,N_14185,N_13598);
and UO_690 (O_690,N_13818,N_14069);
nand UO_691 (O_691,N_12568,N_13396);
and UO_692 (O_692,N_12346,N_14574);
nor UO_693 (O_693,N_12198,N_14759);
nor UO_694 (O_694,N_13978,N_13790);
or UO_695 (O_695,N_14075,N_12282);
nor UO_696 (O_696,N_14971,N_12605);
nand UO_697 (O_697,N_14138,N_13950);
or UO_698 (O_698,N_13620,N_12457);
nand UO_699 (O_699,N_13409,N_13764);
or UO_700 (O_700,N_12305,N_14174);
nor UO_701 (O_701,N_13168,N_13411);
nor UO_702 (O_702,N_13431,N_13684);
xnor UO_703 (O_703,N_14844,N_13172);
nand UO_704 (O_704,N_13120,N_12611);
nand UO_705 (O_705,N_14249,N_13418);
nor UO_706 (O_706,N_13554,N_13629);
and UO_707 (O_707,N_13458,N_12019);
and UO_708 (O_708,N_13094,N_12037);
or UO_709 (O_709,N_13143,N_13876);
nand UO_710 (O_710,N_14110,N_13733);
nor UO_711 (O_711,N_12189,N_13056);
nor UO_712 (O_712,N_12987,N_13668);
and UO_713 (O_713,N_13502,N_12490);
or UO_714 (O_714,N_14698,N_12889);
nand UO_715 (O_715,N_14521,N_13538);
nor UO_716 (O_716,N_14823,N_14350);
or UO_717 (O_717,N_12664,N_12147);
or UO_718 (O_718,N_13833,N_12007);
nor UO_719 (O_719,N_12960,N_14345);
or UO_720 (O_720,N_13140,N_14215);
and UO_721 (O_721,N_13224,N_13540);
or UO_722 (O_722,N_14137,N_12984);
nor UO_723 (O_723,N_13065,N_14469);
nand UO_724 (O_724,N_13496,N_12907);
and UO_725 (O_725,N_14106,N_12031);
or UO_726 (O_726,N_12458,N_13605);
or UO_727 (O_727,N_14140,N_12515);
or UO_728 (O_728,N_12706,N_14453);
or UO_729 (O_729,N_12750,N_13525);
and UO_730 (O_730,N_14504,N_12520);
or UO_731 (O_731,N_13613,N_14378);
or UO_732 (O_732,N_14126,N_12533);
or UO_733 (O_733,N_13500,N_12073);
and UO_734 (O_734,N_13126,N_12990);
or UO_735 (O_735,N_14798,N_13093);
nor UO_736 (O_736,N_12595,N_14390);
and UO_737 (O_737,N_13365,N_14854);
nor UO_738 (O_738,N_14376,N_13926);
or UO_739 (O_739,N_12297,N_13339);
nor UO_740 (O_740,N_13719,N_12745);
or UO_741 (O_741,N_13149,N_12298);
nor UO_742 (O_742,N_12940,N_13826);
nand UO_743 (O_743,N_14054,N_12609);
and UO_744 (O_744,N_12130,N_14281);
nand UO_745 (O_745,N_12146,N_14641);
nand UO_746 (O_746,N_13856,N_13670);
nor UO_747 (O_747,N_12192,N_13526);
and UO_748 (O_748,N_14156,N_13555);
and UO_749 (O_749,N_12454,N_12315);
nor UO_750 (O_750,N_13578,N_13956);
or UO_751 (O_751,N_14434,N_13371);
nor UO_752 (O_752,N_12109,N_12514);
nor UO_753 (O_753,N_12152,N_12938);
or UO_754 (O_754,N_12477,N_13395);
nor UO_755 (O_755,N_13938,N_13266);
nand UO_756 (O_756,N_14506,N_13664);
nand UO_757 (O_757,N_13356,N_13051);
or UO_758 (O_758,N_13552,N_13759);
and UO_759 (O_759,N_14604,N_13319);
and UO_760 (O_760,N_12689,N_12513);
nand UO_761 (O_761,N_14030,N_14245);
nand UO_762 (O_762,N_12178,N_14033);
nand UO_763 (O_763,N_14113,N_12694);
or UO_764 (O_764,N_12000,N_14143);
nor UO_765 (O_765,N_12177,N_13269);
nor UO_766 (O_766,N_13840,N_13290);
nor UO_767 (O_767,N_14133,N_14529);
and UO_768 (O_768,N_12240,N_14932);
nor UO_769 (O_769,N_12561,N_12979);
and UO_770 (O_770,N_12824,N_12124);
nor UO_771 (O_771,N_14646,N_12506);
and UO_772 (O_772,N_13227,N_12773);
and UO_773 (O_773,N_12614,N_13399);
nand UO_774 (O_774,N_13137,N_14003);
or UO_775 (O_775,N_12519,N_13248);
or UO_776 (O_776,N_14526,N_13524);
nor UO_777 (O_777,N_12646,N_12277);
and UO_778 (O_778,N_12834,N_12254);
and UO_779 (O_779,N_14442,N_14575);
or UO_780 (O_780,N_12887,N_14684);
or UO_781 (O_781,N_14422,N_13794);
or UO_782 (O_782,N_12816,N_12842);
and UO_783 (O_783,N_12528,N_12094);
or UO_784 (O_784,N_12966,N_12176);
nor UO_785 (O_785,N_14510,N_14420);
nand UO_786 (O_786,N_14753,N_14222);
nand UO_787 (O_787,N_12702,N_13691);
and UO_788 (O_788,N_13343,N_14556);
and UO_789 (O_789,N_13462,N_14195);
and UO_790 (O_790,N_14963,N_12662);
nor UO_791 (O_791,N_12163,N_12062);
or UO_792 (O_792,N_13710,N_12122);
nor UO_793 (O_793,N_13863,N_13081);
nand UO_794 (O_794,N_12879,N_13017);
nand UO_795 (O_795,N_14308,N_12269);
nand UO_796 (O_796,N_13421,N_12551);
nand UO_797 (O_797,N_14624,N_12420);
nand UO_798 (O_798,N_14922,N_12375);
or UO_799 (O_799,N_13494,N_12667);
nor UO_800 (O_800,N_13720,N_12833);
nand UO_801 (O_801,N_12741,N_12350);
nor UO_802 (O_802,N_12442,N_13184);
nand UO_803 (O_803,N_13742,N_13139);
and UO_804 (O_804,N_13679,N_12601);
nor UO_805 (O_805,N_13869,N_12294);
nor UO_806 (O_806,N_12625,N_14095);
or UO_807 (O_807,N_14731,N_13087);
or UO_808 (O_808,N_13685,N_14207);
or UO_809 (O_809,N_13499,N_14082);
nand UO_810 (O_810,N_13896,N_13357);
and UO_811 (O_811,N_12399,N_13242);
nand UO_812 (O_812,N_13213,N_13095);
nor UO_813 (O_813,N_12582,N_13786);
and UO_814 (O_814,N_12357,N_13099);
nand UO_815 (O_815,N_13571,N_13069);
nand UO_816 (O_816,N_14513,N_14542);
nor UO_817 (O_817,N_14954,N_12329);
or UO_818 (O_818,N_12613,N_14401);
or UO_819 (O_819,N_13705,N_14588);
and UO_820 (O_820,N_13331,N_13080);
or UO_821 (O_821,N_13279,N_12405);
and UO_822 (O_822,N_14958,N_13109);
nand UO_823 (O_823,N_14362,N_12950);
xnor UO_824 (O_824,N_12935,N_13701);
or UO_825 (O_825,N_14055,N_13028);
nand UO_826 (O_826,N_13832,N_14181);
or UO_827 (O_827,N_14470,N_13814);
nor UO_828 (O_828,N_14814,N_12437);
and UO_829 (O_829,N_14343,N_12644);
nand UO_830 (O_830,N_12251,N_14061);
and UO_831 (O_831,N_12738,N_12201);
nand UO_832 (O_832,N_13747,N_14353);
nor UO_833 (O_833,N_14019,N_14901);
and UO_834 (O_834,N_13106,N_14780);
and UO_835 (O_835,N_12777,N_12575);
and UO_836 (O_836,N_12368,N_14783);
nand UO_837 (O_837,N_14165,N_14605);
and UO_838 (O_838,N_12872,N_14508);
or UO_839 (O_839,N_13796,N_12302);
or UO_840 (O_840,N_12678,N_14050);
nor UO_841 (O_841,N_14558,N_12753);
nand UO_842 (O_842,N_12825,N_14620);
nand UO_843 (O_843,N_12214,N_14523);
nor UO_844 (O_844,N_14863,N_13780);
nor UO_845 (O_845,N_13998,N_13461);
nand UO_846 (O_846,N_13302,N_12434);
nor UO_847 (O_847,N_14373,N_12097);
nor UO_848 (O_848,N_12721,N_13249);
or UO_849 (O_849,N_12848,N_14014);
and UO_850 (O_850,N_12897,N_13098);
or UO_851 (O_851,N_14479,N_13889);
or UO_852 (O_852,N_14520,N_13858);
or UO_853 (O_853,N_12243,N_13570);
or UO_854 (O_854,N_14197,N_13360);
nand UO_855 (O_855,N_14546,N_13245);
or UO_856 (O_856,N_13124,N_14145);
nand UO_857 (O_857,N_12013,N_12353);
nor UO_858 (O_858,N_12208,N_13678);
or UO_859 (O_859,N_13152,N_13787);
and UO_860 (O_860,N_12341,N_12875);
and UO_861 (O_861,N_13072,N_14132);
or UO_862 (O_862,N_12112,N_14884);
or UO_863 (O_863,N_13783,N_14679);
nor UO_864 (O_864,N_12029,N_14501);
or UO_865 (O_865,N_14387,N_12117);
nor UO_866 (O_866,N_14051,N_12604);
nor UO_867 (O_867,N_12119,N_13030);
nor UO_868 (O_868,N_14161,N_13308);
nor UO_869 (O_869,N_14655,N_14794);
or UO_870 (O_870,N_13221,N_14637);
nand UO_871 (O_871,N_14059,N_14437);
nand UO_872 (O_872,N_14593,N_13262);
nand UO_873 (O_873,N_14949,N_14071);
nand UO_874 (O_874,N_14375,N_12285);
nor UO_875 (O_875,N_13225,N_14740);
and UO_876 (O_876,N_13706,N_13280);
and UO_877 (O_877,N_13945,N_14417);
and UO_878 (O_878,N_13531,N_14457);
or UO_879 (O_879,N_14638,N_13514);
nand UO_880 (O_880,N_13799,N_13721);
nand UO_881 (O_881,N_13726,N_14856);
nand UO_882 (O_882,N_12300,N_14193);
or UO_883 (O_883,N_12044,N_14472);
nor UO_884 (O_884,N_13022,N_12174);
or UO_885 (O_885,N_12462,N_14563);
and UO_886 (O_886,N_14962,N_14957);
or UO_887 (O_887,N_14400,N_12722);
nand UO_888 (O_888,N_14615,N_13204);
and UO_889 (O_889,N_13969,N_14084);
nor UO_890 (O_890,N_13997,N_14414);
nor UO_891 (O_891,N_14578,N_13849);
and UO_892 (O_892,N_12364,N_13592);
or UO_893 (O_893,N_13510,N_13135);
and UO_894 (O_894,N_12977,N_12972);
and UO_895 (O_895,N_12407,N_14319);
nor UO_896 (O_896,N_13263,N_14701);
and UO_897 (O_897,N_12292,N_12323);
nor UO_898 (O_898,N_13036,N_13083);
and UO_899 (O_899,N_12945,N_12804);
nor UO_900 (O_900,N_13760,N_13424);
and UO_901 (O_901,N_13338,N_14986);
and UO_902 (O_902,N_12577,N_13808);
nor UO_903 (O_903,N_12139,N_12422);
or UO_904 (O_904,N_14303,N_12416);
and UO_905 (O_905,N_12072,N_13931);
and UO_906 (O_906,N_13209,N_13781);
and UO_907 (O_907,N_14365,N_14590);
nand UO_908 (O_908,N_13155,N_12994);
or UO_909 (O_909,N_12370,N_12527);
or UO_910 (O_910,N_12186,N_12589);
and UO_911 (O_911,N_14776,N_12782);
nand UO_912 (O_912,N_12417,N_12989);
and UO_913 (O_913,N_14871,N_13141);
xnor UO_914 (O_914,N_14405,N_13449);
nor UO_915 (O_915,N_14380,N_14081);
or UO_916 (O_916,N_12175,N_13985);
or UO_917 (O_917,N_14811,N_12059);
nor UO_918 (O_918,N_12074,N_14430);
and UO_919 (O_919,N_12242,N_14339);
nor UO_920 (O_920,N_13264,N_13034);
or UO_921 (O_921,N_14238,N_12894);
and UO_922 (O_922,N_14782,N_12597);
xnor UO_923 (O_923,N_13128,N_12992);
or UO_924 (O_924,N_14900,N_13133);
or UO_925 (O_925,N_13466,N_14065);
or UO_926 (O_926,N_14987,N_12355);
or UO_927 (O_927,N_14277,N_14076);
nand UO_928 (O_928,N_14774,N_12949);
nand UO_929 (O_929,N_12247,N_12913);
and UO_930 (O_930,N_14024,N_14148);
or UO_931 (O_931,N_12549,N_13062);
and UO_932 (O_932,N_13567,N_12157);
and UO_933 (O_933,N_14562,N_13074);
or UO_934 (O_934,N_13557,N_12256);
nor UO_935 (O_935,N_14725,N_14254);
and UO_936 (O_936,N_13959,N_12670);
nor UO_937 (O_937,N_14384,N_14040);
and UO_938 (O_938,N_14834,N_12391);
nand UO_939 (O_939,N_13825,N_12563);
nor UO_940 (O_940,N_13806,N_13694);
or UO_941 (O_941,N_14361,N_12444);
nor UO_942 (O_942,N_12854,N_13677);
nand UO_943 (O_943,N_13900,N_14108);
nor UO_944 (O_944,N_12799,N_12788);
nand UO_945 (O_945,N_12017,N_12090);
and UO_946 (O_946,N_12594,N_13676);
and UO_947 (O_947,N_13283,N_12828);
and UO_948 (O_948,N_12576,N_12718);
nor UO_949 (O_949,N_14998,N_13963);
nor UO_950 (O_950,N_13070,N_14683);
and UO_951 (O_951,N_12274,N_13617);
or UO_952 (O_952,N_13114,N_13111);
and UO_953 (O_953,N_13085,N_12714);
or UO_954 (O_954,N_14677,N_13593);
nor UO_955 (O_955,N_13573,N_13361);
or UO_956 (O_956,N_14332,N_12557);
nor UO_957 (O_957,N_12089,N_14817);
nor UO_958 (O_958,N_13841,N_14424);
or UO_959 (O_959,N_14633,N_13179);
nor UO_960 (O_960,N_13498,N_14318);
or UO_961 (O_961,N_14611,N_13663);
or UO_962 (O_962,N_13778,N_13805);
or UO_963 (O_963,N_14053,N_13530);
or UO_964 (O_964,N_13562,N_14229);
nand UO_965 (O_965,N_14919,N_12384);
nand UO_966 (O_966,N_14970,N_14681);
and UO_967 (O_967,N_13941,N_14913);
or UO_968 (O_968,N_12599,N_14211);
or UO_969 (O_969,N_13480,N_14777);
or UO_970 (O_970,N_12016,N_14853);
nor UO_971 (O_971,N_12853,N_13824);
or UO_972 (O_972,N_12374,N_14087);
and UO_973 (O_973,N_14955,N_12035);
nor UO_974 (O_974,N_13166,N_13599);
nand UO_975 (O_975,N_13144,N_12371);
nand UO_976 (O_976,N_12460,N_12313);
nand UO_977 (O_977,N_12901,N_12156);
nor UO_978 (O_978,N_14136,N_12749);
xnor UO_979 (O_979,N_12852,N_14657);
nor UO_980 (O_980,N_13285,N_13643);
or UO_981 (O_981,N_14671,N_13565);
and UO_982 (O_982,N_14346,N_12268);
nor UO_983 (O_983,N_12755,N_13345);
or UO_984 (O_984,N_13602,N_13632);
or UO_985 (O_985,N_13307,N_13377);
xor UO_986 (O_986,N_14089,N_14435);
nor UO_987 (O_987,N_12423,N_13190);
or UO_988 (O_988,N_14157,N_12299);
nor UO_989 (O_989,N_14482,N_12725);
nand UO_990 (O_990,N_12669,N_12995);
or UO_991 (O_991,N_13474,N_14393);
nand UO_992 (O_992,N_13697,N_14297);
and UO_993 (O_993,N_13862,N_13484);
nor UO_994 (O_994,N_14341,N_12581);
and UO_995 (O_995,N_14440,N_13021);
or UO_996 (O_996,N_14617,N_13327);
and UO_997 (O_997,N_14348,N_12598);
or UO_998 (O_998,N_12250,N_12693);
nor UO_999 (O_999,N_13982,N_13875);
and UO_1000 (O_1000,N_14917,N_14936);
or UO_1001 (O_1001,N_12205,N_13322);
nor UO_1002 (O_1002,N_13793,N_13243);
and UO_1003 (O_1003,N_14313,N_12632);
and UO_1004 (O_1004,N_12476,N_14151);
or UO_1005 (O_1005,N_12636,N_12649);
nand UO_1006 (O_1006,N_13949,N_13768);
nand UO_1007 (O_1007,N_13079,N_13801);
nor UO_1008 (O_1008,N_13600,N_12093);
nor UO_1009 (O_1009,N_12228,N_13419);
or UO_1010 (O_1010,N_14739,N_12534);
or UO_1011 (O_1011,N_13255,N_12771);
nand UO_1012 (O_1012,N_13091,N_12784);
and UO_1013 (O_1013,N_14764,N_13215);
or UO_1014 (O_1014,N_14552,N_13320);
nor UO_1015 (O_1015,N_14335,N_12688);
and UO_1016 (O_1016,N_12210,N_13544);
nand UO_1017 (O_1017,N_14648,N_13158);
nor UO_1018 (O_1018,N_12985,N_13656);
or UO_1019 (O_1019,N_14298,N_14601);
nand UO_1020 (O_1020,N_12583,N_13966);
and UO_1021 (O_1021,N_14872,N_13646);
nor UO_1022 (O_1022,N_14493,N_12779);
or UO_1023 (O_1023,N_12728,N_13432);
xor UO_1024 (O_1024,N_13625,N_12104);
or UO_1025 (O_1025,N_14630,N_13268);
nor UO_1026 (O_1026,N_12510,N_13865);
or UO_1027 (O_1027,N_14022,N_14826);
or UO_1028 (O_1028,N_13240,N_13981);
and UO_1029 (O_1029,N_13275,N_12439);
nor UO_1030 (O_1030,N_12321,N_12004);
and UO_1031 (O_1031,N_14952,N_13572);
and UO_1032 (O_1032,N_13903,N_12951);
xnor UO_1033 (O_1033,N_12640,N_14439);
or UO_1034 (O_1034,N_12580,N_13201);
or UO_1035 (O_1035,N_12933,N_12288);
nor UO_1036 (O_1036,N_14744,N_14419);
nand UO_1037 (O_1037,N_13866,N_12441);
nand UO_1038 (O_1038,N_12239,N_13842);
nand UO_1039 (O_1039,N_14839,N_12125);
nor UO_1040 (O_1040,N_13054,N_13438);
nor UO_1041 (O_1041,N_13507,N_13568);
or UO_1042 (O_1042,N_12154,N_13947);
and UO_1043 (O_1043,N_13713,N_13680);
or UO_1044 (O_1044,N_12266,N_14490);
or UO_1045 (O_1045,N_14746,N_13400);
or UO_1046 (O_1046,N_13161,N_13859);
or UO_1047 (O_1047,N_12730,N_14209);
and UO_1048 (O_1048,N_13594,N_12105);
nor UO_1049 (O_1049,N_13237,N_14282);
and UO_1050 (O_1050,N_14029,N_14317);
or UO_1051 (O_1051,N_13844,N_13604);
nand UO_1052 (O_1052,N_13955,N_12207);
or UO_1053 (O_1053,N_13888,N_14733);
nand UO_1054 (O_1054,N_12359,N_14443);
nand UO_1055 (O_1055,N_12786,N_14261);
nand UO_1056 (O_1056,N_13103,N_13160);
nand UO_1057 (O_1057,N_13430,N_14389);
nand UO_1058 (O_1058,N_12654,N_13672);
or UO_1059 (O_1059,N_13988,N_13127);
or UO_1060 (O_1060,N_13909,N_14131);
nor UO_1061 (O_1061,N_13809,N_13066);
nor UO_1062 (O_1062,N_12075,N_12926);
and UO_1063 (O_1063,N_13335,N_14865);
and UO_1064 (O_1064,N_12660,N_14896);
nand UO_1065 (O_1065,N_12881,N_14827);
nand UO_1066 (O_1066,N_14187,N_14077);
nor UO_1067 (O_1067,N_12827,N_14386);
and UO_1068 (O_1068,N_14806,N_14429);
nand UO_1069 (O_1069,N_13725,N_12426);
nor UO_1070 (O_1070,N_12617,N_13208);
nor UO_1071 (O_1071,N_14431,N_12529);
and UO_1072 (O_1072,N_12956,N_14438);
nand UO_1073 (O_1073,N_12427,N_14728);
nor UO_1074 (O_1074,N_13296,N_14597);
nand UO_1075 (O_1075,N_12712,N_12942);
nand UO_1076 (O_1076,N_12866,N_13980);
and UO_1077 (O_1077,N_13699,N_13836);
nand UO_1078 (O_1078,N_13329,N_14612);
or UO_1079 (O_1079,N_13968,N_14208);
nand UO_1080 (O_1080,N_14129,N_13908);
nor UO_1081 (O_1081,N_12739,N_12876);
nor UO_1082 (O_1082,N_12312,N_13655);
nor UO_1083 (O_1083,N_14247,N_14183);
or UO_1084 (O_1084,N_14202,N_14200);
or UO_1085 (O_1085,N_13310,N_14995);
and UO_1086 (O_1086,N_14688,N_13100);
nand UO_1087 (O_1087,N_12600,N_14766);
or UO_1088 (O_1088,N_14496,N_13921);
nor UO_1089 (O_1089,N_13746,N_13469);
nor UO_1090 (O_1090,N_14825,N_13901);
and UO_1091 (O_1091,N_14864,N_14026);
or UO_1092 (O_1092,N_13791,N_12628);
nand UO_1093 (O_1093,N_12744,N_13574);
and UO_1094 (O_1094,N_14883,N_14456);
and UO_1095 (O_1095,N_12365,N_12572);
nor UO_1096 (O_1096,N_12516,N_12587);
nor UO_1097 (O_1097,N_12270,N_12540);
and UO_1098 (O_1098,N_13671,N_13389);
nand UO_1099 (O_1099,N_14675,N_14654);
or UO_1100 (O_1100,N_13773,N_12924);
or UO_1101 (O_1101,N_14704,N_12284);
or UO_1102 (O_1102,N_12555,N_12925);
nand UO_1103 (O_1103,N_14099,N_13390);
nor UO_1104 (O_1104,N_13884,N_12020);
or UO_1105 (O_1105,N_13231,N_13536);
nand UO_1106 (O_1106,N_14697,N_13104);
nor UO_1107 (O_1107,N_12264,N_13811);
or UO_1108 (O_1108,N_13350,N_12971);
nand UO_1109 (O_1109,N_13029,N_14305);
and UO_1110 (O_1110,N_13415,N_12351);
nand UO_1111 (O_1111,N_14775,N_12703);
or UO_1112 (O_1112,N_12082,N_12479);
nor UO_1113 (O_1113,N_13259,N_13576);
or UO_1114 (O_1114,N_14670,N_12579);
nand UO_1115 (O_1115,N_14253,N_12493);
nand UO_1116 (O_1116,N_12683,N_13928);
and UO_1117 (O_1117,N_14721,N_14191);
or UO_1118 (O_1118,N_12057,N_12278);
nand UO_1119 (O_1119,N_14027,N_12946);
nand UO_1120 (O_1120,N_12499,N_13891);
or UO_1121 (O_1121,N_13819,N_14295);
nand UO_1122 (O_1122,N_12030,N_12183);
and UO_1123 (O_1123,N_12419,N_14230);
nor UO_1124 (O_1124,N_12361,N_13815);
nor UO_1125 (O_1125,N_12049,N_14337);
and UO_1126 (O_1126,N_14583,N_13097);
or UO_1127 (O_1127,N_14107,N_14765);
or UO_1128 (O_1128,N_12682,N_12772);
nor UO_1129 (O_1129,N_14923,N_13366);
nand UO_1130 (O_1130,N_13972,N_14812);
nand UO_1131 (O_1131,N_13529,N_13383);
or UO_1132 (O_1132,N_13930,N_14889);
or UO_1133 (O_1133,N_12704,N_14835);
and UO_1134 (O_1134,N_14485,N_14712);
nand UO_1135 (O_1135,N_12255,N_14895);
and UO_1136 (O_1136,N_12792,N_14862);
nor UO_1137 (O_1137,N_12705,N_12400);
nor UO_1138 (O_1138,N_14629,N_13257);
nor UO_1139 (O_1139,N_12656,N_14752);
nor UO_1140 (O_1140,N_13129,N_13495);
or UO_1141 (O_1141,N_14502,N_14915);
and UO_1142 (O_1142,N_13551,N_14190);
nand UO_1143 (O_1143,N_14481,N_12865);
nand UO_1144 (O_1144,N_12110,N_13508);
or UO_1145 (O_1145,N_14283,N_14797);
or UO_1146 (O_1146,N_12797,N_12159);
or UO_1147 (O_1147,N_13925,N_14168);
nor UO_1148 (O_1148,N_12969,N_14112);
or UO_1149 (O_1149,N_13084,N_13639);
nand UO_1150 (O_1150,N_12219,N_12982);
nor UO_1151 (O_1151,N_14606,N_13244);
nand UO_1152 (O_1152,N_12406,N_13019);
nand UO_1153 (O_1153,N_13990,N_14989);
and UO_1154 (O_1154,N_12432,N_12762);
or UO_1155 (O_1155,N_12366,N_13607);
and UO_1156 (O_1156,N_12382,N_14356);
nor UO_1157 (O_1157,N_13199,N_13880);
or UO_1158 (O_1158,N_12141,N_14666);
nor UO_1159 (O_1159,N_14465,N_14598);
or UO_1160 (O_1160,N_13893,N_14807);
nor UO_1161 (O_1161,N_14713,N_12892);
or UO_1162 (O_1162,N_14158,N_14166);
nor UO_1163 (O_1163,N_14272,N_14543);
nor UO_1164 (O_1164,N_14352,N_13378);
and UO_1165 (O_1165,N_12758,N_12774);
or UO_1166 (O_1166,N_12564,N_14130);
nor UO_1167 (O_1167,N_14760,N_12390);
or UO_1168 (O_1168,N_13416,N_12709);
nor UO_1169 (O_1169,N_12863,N_14498);
nor UO_1170 (O_1170,N_12418,N_14720);
nand UO_1171 (O_1171,N_12629,N_13234);
or UO_1172 (O_1172,N_13454,N_12440);
or UO_1173 (O_1173,N_14357,N_13381);
nand UO_1174 (O_1174,N_14104,N_12695);
and UO_1175 (O_1175,N_14626,N_14256);
nor UO_1176 (O_1176,N_12948,N_13488);
or UO_1177 (O_1177,N_12222,N_14603);
nor UO_1178 (O_1178,N_12864,N_14993);
and UO_1179 (O_1179,N_13645,N_14172);
nand UO_1180 (O_1180,N_14736,N_13716);
nand UO_1181 (O_1181,N_13581,N_12903);
or UO_1182 (O_1182,N_14548,N_12732);
and UO_1183 (O_1183,N_12435,N_14269);
nor UO_1184 (O_1184,N_13587,N_14399);
and UO_1185 (O_1185,N_13700,N_14057);
nand UO_1186 (O_1186,N_14851,N_14500);
or UO_1187 (O_1187,N_14700,N_14090);
or UO_1188 (O_1188,N_12402,N_12780);
and UO_1189 (O_1189,N_13669,N_12770);
nand UO_1190 (O_1190,N_14098,N_13226);
xor UO_1191 (O_1191,N_14206,N_13772);
or UO_1192 (O_1192,N_13729,N_13518);
nand UO_1193 (O_1193,N_13877,N_12593);
and UO_1194 (O_1194,N_14182,N_14114);
nand UO_1195 (O_1195,N_12847,N_13429);
or UO_1196 (O_1196,N_13261,N_12882);
or UO_1197 (O_1197,N_13545,N_13527);
nor UO_1198 (O_1198,N_14409,N_14001);
and UO_1199 (O_1199,N_13118,N_13407);
nand UO_1200 (O_1200,N_12518,N_14415);
xnor UO_1201 (O_1201,N_13838,N_14369);
nand UO_1202 (O_1202,N_13546,N_12571);
nand UO_1203 (O_1203,N_13175,N_14404);
nor UO_1204 (O_1204,N_13299,N_12068);
and UO_1205 (O_1205,N_13828,N_12026);
xor UO_1206 (O_1206,N_14691,N_13654);
nor UO_1207 (O_1207,N_14890,N_14933);
nand UO_1208 (O_1208,N_12974,N_12215);
and UO_1209 (O_1209,N_13241,N_14312);
nand UO_1210 (O_1210,N_12115,N_13650);
nor UO_1211 (O_1211,N_14381,N_14916);
nand UO_1212 (O_1212,N_13410,N_12153);
and UO_1213 (O_1213,N_13068,N_12916);
or UO_1214 (O_1214,N_14286,N_12227);
nand UO_1215 (O_1215,N_14178,N_14306);
nor UO_1216 (O_1216,N_12425,N_12691);
and UO_1217 (O_1217,N_13233,N_13927);
nand UO_1218 (O_1218,N_13933,N_12466);
nor UO_1219 (O_1219,N_12098,N_14781);
and UO_1220 (O_1220,N_13942,N_13123);
nor UO_1221 (O_1221,N_13216,N_12535);
nand UO_1222 (O_1222,N_13044,N_14858);
or UO_1223 (O_1223,N_12136,N_13549);
nor UO_1224 (O_1224,N_14015,N_14242);
xor UO_1225 (O_1225,N_12102,N_12986);
nor UO_1226 (O_1226,N_13698,N_13917);
or UO_1227 (O_1227,N_12397,N_12475);
or UO_1228 (O_1228,N_14446,N_12168);
or UO_1229 (O_1229,N_13163,N_14829);
and UO_1230 (O_1230,N_13944,N_13358);
and UO_1231 (O_1231,N_12931,N_13611);
or UO_1232 (O_1232,N_12886,N_12339);
nand UO_1233 (O_1233,N_14259,N_13872);
nor UO_1234 (O_1234,N_12621,N_14694);
nor UO_1235 (O_1235,N_13626,N_12532);
or UO_1236 (O_1236,N_14002,N_13965);
nand UO_1237 (O_1237,N_12063,N_12651);
and UO_1238 (O_1238,N_14000,N_12316);
nand UO_1239 (O_1239,N_14125,N_14667);
nor UO_1240 (O_1240,N_13230,N_14153);
nand UO_1241 (O_1241,N_14785,N_13403);
or UO_1242 (O_1242,N_14411,N_12171);
nand UO_1243 (O_1243,N_14170,N_13489);
nand UO_1244 (O_1244,N_13309,N_12128);
and UO_1245 (O_1245,N_12953,N_12813);
or UO_1246 (O_1246,N_14370,N_13924);
or UO_1247 (O_1247,N_12113,N_14579);
xor UO_1248 (O_1248,N_12681,N_13967);
xor UO_1249 (O_1249,N_12538,N_14410);
or UO_1250 (O_1250,N_14530,N_14428);
nand UO_1251 (O_1251,N_13253,N_13078);
nor UO_1252 (O_1252,N_12668,N_14550);
or UO_1253 (O_1253,N_12643,N_14289);
nor UO_1254 (O_1254,N_12778,N_13511);
or UO_1255 (O_1255,N_14425,N_12358);
nand UO_1256 (O_1256,N_12066,N_13025);
nor UO_1257 (O_1257,N_12200,N_14741);
nor UO_1258 (O_1258,N_12964,N_12388);
and UO_1259 (O_1259,N_13055,N_13391);
or UO_1260 (O_1260,N_13113,N_14066);
nand UO_1261 (O_1261,N_14947,N_12018);
and UO_1262 (O_1262,N_14946,N_12502);
nand UO_1263 (O_1263,N_12413,N_12160);
and UO_1264 (O_1264,N_13218,N_12194);
nor UO_1265 (O_1265,N_13284,N_14251);
nand UO_1266 (O_1266,N_12553,N_12687);
nor UO_1267 (O_1267,N_14285,N_12760);
nor UO_1268 (O_1268,N_13297,N_14036);
or UO_1269 (O_1269,N_14338,N_14307);
nor UO_1270 (O_1270,N_12905,N_14727);
and UO_1271 (O_1271,N_13354,N_14669);
nor UO_1272 (O_1272,N_13206,N_12610);
or UO_1273 (O_1273,N_12482,N_13131);
or UO_1274 (O_1274,N_12252,N_12071);
or UO_1275 (O_1275,N_14016,N_14547);
nand UO_1276 (O_1276,N_13101,N_12708);
nand UO_1277 (O_1277,N_14413,N_14645);
or UO_1278 (O_1278,N_13873,N_14176);
nand UO_1279 (O_1279,N_13490,N_12084);
or UO_1280 (O_1280,N_13845,N_13112);
nand UO_1281 (O_1281,N_13539,N_12224);
nand UO_1282 (O_1282,N_12858,N_14536);
nand UO_1283 (O_1283,N_12965,N_13108);
nor UO_1284 (O_1284,N_14359,N_12204);
or UO_1285 (O_1285,N_14340,N_14769);
nand UO_1286 (O_1286,N_12958,N_13132);
nor UO_1287 (O_1287,N_12114,N_13582);
nor UO_1288 (O_1288,N_13368,N_12005);
and UO_1289 (O_1289,N_12412,N_12180);
and UO_1290 (O_1290,N_12383,N_14146);
or UO_1291 (O_1291,N_14309,N_13031);
and UO_1292 (O_1292,N_13929,N_13183);
and UO_1293 (O_1293,N_12369,N_12431);
nand UO_1294 (O_1294,N_13016,N_12481);
or UO_1295 (O_1295,N_13181,N_14847);
and UO_1296 (O_1296,N_12698,N_12634);
nor UO_1297 (O_1297,N_13273,N_13874);
and UO_1298 (O_1298,N_13096,N_12543);
or UO_1299 (O_1299,N_12069,N_14702);
and UO_1300 (O_1300,N_13041,N_12663);
nand UO_1301 (O_1301,N_14838,N_14860);
and UO_1302 (O_1302,N_14300,N_12080);
and UO_1303 (O_1303,N_14639,N_12548);
or UO_1304 (O_1304,N_12220,N_12342);
nor UO_1305 (O_1305,N_12726,N_13211);
nand UO_1306 (O_1306,N_14232,N_14627);
or UO_1307 (O_1307,N_13975,N_13142);
or UO_1308 (O_1308,N_13467,N_13256);
and UO_1309 (O_1309,N_13659,N_13722);
or UO_1310 (O_1310,N_13627,N_13007);
and UO_1311 (O_1311,N_14848,N_12902);
and UO_1312 (O_1312,N_13453,N_14897);
nand UO_1313 (O_1313,N_12616,N_12401);
nor UO_1314 (O_1314,N_14582,N_14179);
nand UO_1315 (O_1315,N_13043,N_14034);
nand UO_1316 (O_1316,N_13071,N_12043);
or UO_1317 (O_1317,N_14690,N_13666);
and UO_1318 (O_1318,N_14449,N_14010);
nor UO_1319 (O_1319,N_12231,N_14815);
nand UO_1320 (O_1320,N_12911,N_14266);
nand UO_1321 (O_1321,N_14246,N_14832);
nor UO_1322 (O_1322,N_12408,N_14186);
or UO_1323 (O_1323,N_12472,N_12735);
or UO_1324 (O_1324,N_12484,N_12040);
and UO_1325 (O_1325,N_13612,N_14078);
nand UO_1326 (O_1326,N_14553,N_13736);
or UO_1327 (O_1327,N_12930,N_13631);
and UO_1328 (O_1328,N_12085,N_14160);
nor UO_1329 (O_1329,N_13739,N_14199);
nand UO_1330 (O_1330,N_14824,N_13394);
nor UO_1331 (O_1331,N_13714,N_12021);
nand UO_1332 (O_1332,N_14749,N_12908);
or UO_1333 (O_1333,N_12898,N_13492);
or UO_1334 (O_1334,N_13447,N_14494);
and UO_1335 (O_1335,N_14678,N_12733);
or UO_1336 (O_1336,N_12308,N_12448);
and UO_1337 (O_1337,N_14139,N_13543);
nand UO_1338 (O_1338,N_14402,N_12290);
and UO_1339 (O_1339,N_13039,N_13798);
or UO_1340 (O_1340,N_14852,N_14368);
and UO_1341 (O_1341,N_12554,N_12943);
nor UO_1342 (O_1342,N_13397,N_12197);
nor UO_1343 (O_1343,N_14793,N_12162);
nand UO_1344 (O_1344,N_12665,N_13984);
or UO_1345 (O_1345,N_13777,N_14237);
nand UO_1346 (O_1346,N_14535,N_13130);
nor UO_1347 (O_1347,N_12713,N_13301);
nand UO_1348 (O_1348,N_12409,N_13235);
or UO_1349 (O_1349,N_14516,N_12961);
nand UO_1350 (O_1350,N_12740,N_14653);
nor UO_1351 (O_1351,N_14788,N_12340);
and UO_1352 (O_1352,N_14891,N_14790);
nand UO_1353 (O_1353,N_13771,N_14085);
and UO_1354 (O_1354,N_14560,N_13122);
or UO_1355 (O_1355,N_13792,N_13907);
or UO_1356 (O_1356,N_14119,N_13662);
nand UO_1357 (O_1357,N_14322,N_13745);
or UO_1358 (O_1358,N_13860,N_14534);
nor UO_1359 (O_1359,N_13603,N_12618);
nor UO_1360 (O_1360,N_13922,N_12336);
and UO_1361 (O_1361,N_14734,N_12785);
or UO_1362 (O_1362,N_14096,N_13505);
or UO_1363 (O_1363,N_14507,N_12392);
or UO_1364 (O_1364,N_12547,N_12307);
nor UO_1365 (O_1365,N_14532,N_13728);
and UO_1366 (O_1366,N_13695,N_13707);
and UO_1367 (O_1367,N_14102,N_12751);
and UO_1368 (O_1368,N_13854,N_14554);
nand UO_1369 (O_1369,N_14846,N_12470);
and UO_1370 (O_1370,N_13304,N_12492);
or UO_1371 (O_1371,N_12209,N_14032);
or UO_1372 (O_1372,N_14592,N_12193);
nand UO_1373 (O_1373,N_12489,N_13804);
and UO_1374 (O_1374,N_14660,N_12795);
and UO_1375 (O_1375,N_12430,N_13703);
xor UO_1376 (O_1376,N_12276,N_12803);
nor UO_1377 (O_1377,N_12067,N_14567);
xnor UO_1378 (O_1378,N_14038,N_13590);
and UO_1379 (O_1379,N_13533,N_12100);
or UO_1380 (O_1380,N_13478,N_13463);
and UO_1381 (O_1381,N_12280,N_14268);
or UO_1382 (O_1382,N_13913,N_12944);
nor UO_1383 (O_1383,N_14881,N_14942);
nand UO_1384 (O_1384,N_14687,N_12560);
nand UO_1385 (O_1385,N_12211,N_14219);
nor UO_1386 (O_1386,N_14045,N_14745);
and UO_1387 (O_1387,N_12790,N_12870);
nand UO_1388 (O_1388,N_12596,N_13641);
nor UO_1389 (O_1389,N_12352,N_13813);
and UO_1390 (O_1390,N_14961,N_12086);
nor UO_1391 (O_1391,N_12835,N_14244);
nand UO_1392 (O_1392,N_13282,N_13586);
nand UO_1393 (O_1393,N_14910,N_12831);
or UO_1394 (O_1394,N_12631,N_13885);
and UO_1395 (O_1395,N_13064,N_13899);
and UO_1396 (O_1396,N_12619,N_14284);
and UO_1397 (O_1397,N_14223,N_13088);
and UO_1398 (O_1398,N_14398,N_13940);
nand UO_1399 (O_1399,N_14857,N_12523);
and UO_1400 (O_1400,N_13267,N_14491);
and UO_1401 (O_1401,N_13501,N_14996);
nand UO_1402 (O_1402,N_14013,N_14980);
or UO_1403 (O_1403,N_12438,N_12253);
or UO_1404 (O_1404,N_12331,N_13996);
or UO_1405 (O_1405,N_12234,N_14039);
nor UO_1406 (O_1406,N_12764,N_12955);
or UO_1407 (O_1407,N_12077,N_14035);
nand UO_1408 (O_1408,N_13195,N_12500);
nand UO_1409 (O_1409,N_13520,N_12999);
nor UO_1410 (O_1410,N_14374,N_14460);
or UO_1411 (O_1411,N_12011,N_13439);
and UO_1412 (O_1412,N_12832,N_12658);
nand UO_1413 (O_1413,N_12317,N_12922);
nor UO_1414 (O_1414,N_13946,N_13715);
nand UO_1415 (O_1415,N_12729,N_13442);
and UO_1416 (O_1416,N_14344,N_13167);
nand UO_1417 (O_1417,N_12776,N_14511);
or UO_1418 (O_1418,N_13176,N_13763);
and UO_1419 (O_1419,N_13138,N_12495);
or UO_1420 (O_1420,N_14619,N_12900);
and UO_1421 (O_1421,N_14086,N_14109);
nor UO_1422 (O_1422,N_13754,N_12123);
nand UO_1423 (O_1423,N_12033,N_13939);
nor UO_1424 (O_1424,N_14302,N_14274);
nand UO_1425 (O_1425,N_12233,N_12260);
nor UO_1426 (O_1426,N_14020,N_14489);
nand UO_1427 (O_1427,N_14294,N_12836);
nor UO_1428 (O_1428,N_13200,N_12808);
nand UO_1429 (O_1429,N_12715,N_14006);
and UO_1430 (O_1430,N_12167,N_14625);
or UO_1431 (O_1431,N_13623,N_12975);
nand UO_1432 (O_1432,N_12761,N_12620);
nand UO_1433 (O_1433,N_14928,N_12565);
and UO_1434 (O_1434,N_14778,N_14514);
and UO_1435 (O_1435,N_13373,N_12763);
nand UO_1436 (O_1436,N_14830,N_12363);
nor UO_1437 (O_1437,N_14471,N_14568);
nor UO_1438 (O_1438,N_12396,N_12754);
nand UO_1439 (O_1439,N_12727,N_13117);
and UO_1440 (O_1440,N_12988,N_13374);
nor UO_1441 (O_1441,N_13638,N_13785);
or UO_1442 (O_1442,N_12083,N_14663);
nand UO_1443 (O_1443,N_13774,N_14758);
nand UO_1444 (O_1444,N_13717,N_14279);
nor UO_1445 (O_1445,N_13822,N_14926);
or UO_1446 (O_1446,N_14616,N_12428);
nand UO_1447 (O_1447,N_13737,N_13757);
or UO_1448 (O_1448,N_13776,N_14586);
nand UO_1449 (O_1449,N_14291,N_13303);
and UO_1450 (O_1450,N_13042,N_13606);
or UO_1451 (O_1451,N_14092,N_12566);
and UO_1452 (O_1452,N_13779,N_12449);
or UO_1453 (O_1453,N_13878,N_14088);
and UO_1454 (O_1454,N_14904,N_13150);
nand UO_1455 (O_1455,N_14124,N_13515);
nand UO_1456 (O_1456,N_13789,N_12333);
nor UO_1457 (O_1457,N_13425,N_12055);
nand UO_1458 (O_1458,N_12973,N_13446);
or UO_1459 (O_1459,N_12883,N_12524);
or UO_1460 (O_1460,N_12216,N_12367);
or UO_1461 (O_1461,N_12766,N_13265);
nor UO_1462 (O_1462,N_14693,N_12039);
and UO_1463 (O_1463,N_12273,N_14960);
and UO_1464 (O_1464,N_14427,N_13073);
nand UO_1465 (O_1465,N_14636,N_12022);
and UO_1466 (O_1466,N_12855,N_14580);
and UO_1467 (O_1467,N_13667,N_12737);
and UO_1468 (O_1468,N_12306,N_12545);
or UO_1469 (O_1469,N_14953,N_13385);
nor UO_1470 (O_1470,N_12261,N_12570);
nand UO_1471 (O_1471,N_13147,N_13615);
and UO_1472 (O_1472,N_14906,N_13635);
or UO_1473 (O_1473,N_13820,N_12024);
nand UO_1474 (O_1474,N_13497,N_14672);
or UO_1475 (O_1475,N_14584,N_14632);
nand UO_1476 (O_1476,N_12257,N_12107);
and UO_1477 (O_1477,N_12143,N_13222);
and UO_1478 (O_1478,N_14561,N_12496);
nor UO_1479 (O_1479,N_14945,N_13012);
nand UO_1480 (O_1480,N_13082,N_14967);
or UO_1481 (O_1481,N_14709,N_14097);
nand UO_1482 (O_1482,N_13169,N_13751);
nor UO_1483 (O_1483,N_13675,N_14557);
and UO_1484 (O_1484,N_13987,N_14763);
and UO_1485 (O_1485,N_14572,N_14280);
and UO_1486 (O_1486,N_12752,N_13883);
and UO_1487 (O_1487,N_12963,N_12459);
nand UO_1488 (O_1488,N_12927,N_12826);
or UO_1489 (O_1489,N_12685,N_14296);
nor UO_1490 (O_1490,N_13935,N_13652);
or UO_1491 (O_1491,N_14171,N_14652);
and UO_1492 (O_1492,N_13165,N_13696);
nand UO_1493 (O_1493,N_14293,N_12172);
nor UO_1494 (O_1494,N_12659,N_12809);
nor UO_1495 (O_1495,N_13911,N_13193);
or UO_1496 (O_1496,N_14531,N_12309);
nor UO_1497 (O_1497,N_12793,N_14525);
nor UO_1498 (O_1498,N_12885,N_13479);
nor UO_1499 (O_1499,N_14372,N_12904);
and UO_1500 (O_1500,N_12937,N_14925);
or UO_1501 (O_1501,N_12639,N_14260);
nand UO_1502 (O_1502,N_14930,N_12546);
or UO_1503 (O_1503,N_12505,N_13340);
nor UO_1504 (O_1504,N_14442,N_12257);
nor UO_1505 (O_1505,N_14040,N_14965);
nand UO_1506 (O_1506,N_12646,N_13509);
and UO_1507 (O_1507,N_12021,N_12793);
nand UO_1508 (O_1508,N_12340,N_13696);
nor UO_1509 (O_1509,N_14082,N_14446);
or UO_1510 (O_1510,N_12654,N_12710);
and UO_1511 (O_1511,N_14811,N_14788);
nand UO_1512 (O_1512,N_12152,N_12795);
nand UO_1513 (O_1513,N_14253,N_14276);
nand UO_1514 (O_1514,N_12853,N_13853);
nor UO_1515 (O_1515,N_14605,N_12795);
nor UO_1516 (O_1516,N_12602,N_13984);
nor UO_1517 (O_1517,N_13447,N_14784);
nand UO_1518 (O_1518,N_12539,N_14071);
or UO_1519 (O_1519,N_14003,N_13468);
or UO_1520 (O_1520,N_14035,N_12172);
and UO_1521 (O_1521,N_13223,N_12175);
nand UO_1522 (O_1522,N_12989,N_12601);
nor UO_1523 (O_1523,N_13610,N_13882);
and UO_1524 (O_1524,N_13961,N_14514);
nor UO_1525 (O_1525,N_12430,N_14369);
and UO_1526 (O_1526,N_12304,N_13880);
nor UO_1527 (O_1527,N_14652,N_12969);
and UO_1528 (O_1528,N_12033,N_14064);
nor UO_1529 (O_1529,N_14361,N_12852);
nand UO_1530 (O_1530,N_13228,N_13849);
and UO_1531 (O_1531,N_14058,N_12683);
nand UO_1532 (O_1532,N_12425,N_14619);
or UO_1533 (O_1533,N_14671,N_14780);
nor UO_1534 (O_1534,N_13007,N_12722);
nor UO_1535 (O_1535,N_14633,N_13290);
nor UO_1536 (O_1536,N_12940,N_13672);
and UO_1537 (O_1537,N_14654,N_14772);
xor UO_1538 (O_1538,N_12572,N_13198);
nor UO_1539 (O_1539,N_12245,N_12581);
nor UO_1540 (O_1540,N_12336,N_13150);
and UO_1541 (O_1541,N_14794,N_14350);
nand UO_1542 (O_1542,N_14307,N_13839);
nor UO_1543 (O_1543,N_13858,N_12825);
nor UO_1544 (O_1544,N_12249,N_13326);
nand UO_1545 (O_1545,N_12273,N_13134);
or UO_1546 (O_1546,N_13959,N_12394);
or UO_1547 (O_1547,N_12709,N_14963);
and UO_1548 (O_1548,N_13557,N_14501);
nor UO_1549 (O_1549,N_13395,N_12078);
and UO_1550 (O_1550,N_14063,N_13860);
or UO_1551 (O_1551,N_13973,N_13646);
and UO_1552 (O_1552,N_14058,N_14481);
nor UO_1553 (O_1553,N_13720,N_13656);
nor UO_1554 (O_1554,N_13618,N_14331);
nand UO_1555 (O_1555,N_12240,N_14125);
and UO_1556 (O_1556,N_13854,N_14341);
nor UO_1557 (O_1557,N_14839,N_12475);
nand UO_1558 (O_1558,N_12468,N_14418);
or UO_1559 (O_1559,N_13089,N_12206);
or UO_1560 (O_1560,N_13099,N_13383);
and UO_1561 (O_1561,N_13680,N_12708);
or UO_1562 (O_1562,N_13219,N_12334);
and UO_1563 (O_1563,N_14035,N_14325);
nor UO_1564 (O_1564,N_12429,N_12249);
or UO_1565 (O_1565,N_13106,N_12594);
and UO_1566 (O_1566,N_13170,N_13611);
and UO_1567 (O_1567,N_12525,N_14787);
or UO_1568 (O_1568,N_13687,N_14352);
and UO_1569 (O_1569,N_12780,N_13143);
and UO_1570 (O_1570,N_13699,N_14830);
nor UO_1571 (O_1571,N_12739,N_12139);
nor UO_1572 (O_1572,N_14153,N_14166);
nor UO_1573 (O_1573,N_12813,N_13403);
nor UO_1574 (O_1574,N_12962,N_13764);
nor UO_1575 (O_1575,N_12393,N_12467);
nor UO_1576 (O_1576,N_13211,N_13703);
nand UO_1577 (O_1577,N_12914,N_12243);
nand UO_1578 (O_1578,N_12423,N_12665);
nor UO_1579 (O_1579,N_12836,N_12235);
nor UO_1580 (O_1580,N_12200,N_12126);
nor UO_1581 (O_1581,N_14637,N_14882);
nand UO_1582 (O_1582,N_14951,N_14601);
and UO_1583 (O_1583,N_12276,N_13907);
or UO_1584 (O_1584,N_14600,N_14990);
nand UO_1585 (O_1585,N_12770,N_13331);
xor UO_1586 (O_1586,N_13251,N_14742);
and UO_1587 (O_1587,N_13478,N_12378);
and UO_1588 (O_1588,N_12960,N_12151);
or UO_1589 (O_1589,N_14167,N_13183);
or UO_1590 (O_1590,N_14919,N_12729);
or UO_1591 (O_1591,N_12021,N_12474);
or UO_1592 (O_1592,N_12894,N_14673);
or UO_1593 (O_1593,N_13049,N_13442);
nor UO_1594 (O_1594,N_12372,N_12554);
nand UO_1595 (O_1595,N_12384,N_13103);
or UO_1596 (O_1596,N_12491,N_13161);
or UO_1597 (O_1597,N_13930,N_12907);
nand UO_1598 (O_1598,N_14861,N_13154);
nand UO_1599 (O_1599,N_13055,N_13409);
and UO_1600 (O_1600,N_14514,N_13933);
nand UO_1601 (O_1601,N_12075,N_14636);
nand UO_1602 (O_1602,N_14107,N_14420);
nor UO_1603 (O_1603,N_12066,N_12153);
nand UO_1604 (O_1604,N_12241,N_12769);
nor UO_1605 (O_1605,N_12869,N_12712);
nand UO_1606 (O_1606,N_13170,N_12298);
nor UO_1607 (O_1607,N_14866,N_13820);
nand UO_1608 (O_1608,N_12999,N_13652);
nor UO_1609 (O_1609,N_12581,N_14637);
or UO_1610 (O_1610,N_14932,N_13117);
and UO_1611 (O_1611,N_14225,N_12242);
and UO_1612 (O_1612,N_13868,N_14627);
or UO_1613 (O_1613,N_13434,N_12465);
nand UO_1614 (O_1614,N_13081,N_13916);
and UO_1615 (O_1615,N_13941,N_12422);
and UO_1616 (O_1616,N_12422,N_13802);
or UO_1617 (O_1617,N_14724,N_14042);
nand UO_1618 (O_1618,N_12130,N_12984);
nor UO_1619 (O_1619,N_13236,N_13786);
nor UO_1620 (O_1620,N_13823,N_13688);
or UO_1621 (O_1621,N_14595,N_12001);
or UO_1622 (O_1622,N_13196,N_13705);
and UO_1623 (O_1623,N_14395,N_12824);
or UO_1624 (O_1624,N_14356,N_14641);
and UO_1625 (O_1625,N_14852,N_14272);
and UO_1626 (O_1626,N_12223,N_14645);
nand UO_1627 (O_1627,N_14653,N_12471);
and UO_1628 (O_1628,N_13493,N_12632);
nand UO_1629 (O_1629,N_13962,N_14130);
nand UO_1630 (O_1630,N_13763,N_12174);
nor UO_1631 (O_1631,N_13967,N_13801);
nand UO_1632 (O_1632,N_13714,N_12809);
nand UO_1633 (O_1633,N_14501,N_13698);
and UO_1634 (O_1634,N_14603,N_12984);
or UO_1635 (O_1635,N_14330,N_14172);
and UO_1636 (O_1636,N_12738,N_13585);
nand UO_1637 (O_1637,N_13233,N_14637);
or UO_1638 (O_1638,N_14341,N_12561);
or UO_1639 (O_1639,N_12558,N_12894);
nor UO_1640 (O_1640,N_14836,N_14571);
nand UO_1641 (O_1641,N_12963,N_13508);
nor UO_1642 (O_1642,N_12699,N_14156);
nor UO_1643 (O_1643,N_14658,N_14310);
nand UO_1644 (O_1644,N_14025,N_14614);
or UO_1645 (O_1645,N_14232,N_12759);
nor UO_1646 (O_1646,N_12622,N_13305);
and UO_1647 (O_1647,N_14480,N_14815);
or UO_1648 (O_1648,N_13886,N_12926);
nand UO_1649 (O_1649,N_12144,N_12763);
nand UO_1650 (O_1650,N_13023,N_13291);
and UO_1651 (O_1651,N_14342,N_13414);
nor UO_1652 (O_1652,N_13736,N_13001);
and UO_1653 (O_1653,N_13179,N_12421);
and UO_1654 (O_1654,N_13168,N_14208);
and UO_1655 (O_1655,N_12819,N_12457);
or UO_1656 (O_1656,N_12608,N_14318);
nand UO_1657 (O_1657,N_12688,N_12931);
nor UO_1658 (O_1658,N_14932,N_12672);
nand UO_1659 (O_1659,N_12980,N_12921);
or UO_1660 (O_1660,N_12340,N_12746);
nor UO_1661 (O_1661,N_13385,N_12578);
nor UO_1662 (O_1662,N_12243,N_13953);
nand UO_1663 (O_1663,N_12710,N_12260);
and UO_1664 (O_1664,N_13692,N_14802);
nor UO_1665 (O_1665,N_13738,N_14609);
nor UO_1666 (O_1666,N_14876,N_14059);
or UO_1667 (O_1667,N_13248,N_12552);
and UO_1668 (O_1668,N_13299,N_14788);
nand UO_1669 (O_1669,N_14977,N_12712);
nand UO_1670 (O_1670,N_12393,N_14388);
and UO_1671 (O_1671,N_13866,N_14409);
and UO_1672 (O_1672,N_13161,N_14280);
or UO_1673 (O_1673,N_12526,N_12062);
and UO_1674 (O_1674,N_12641,N_14652);
and UO_1675 (O_1675,N_13158,N_13120);
nand UO_1676 (O_1676,N_14871,N_14329);
and UO_1677 (O_1677,N_12767,N_13081);
nand UO_1678 (O_1678,N_14363,N_14984);
and UO_1679 (O_1679,N_14897,N_13085);
nand UO_1680 (O_1680,N_14175,N_12638);
nand UO_1681 (O_1681,N_13063,N_14648);
and UO_1682 (O_1682,N_14089,N_14418);
nand UO_1683 (O_1683,N_13763,N_13046);
nand UO_1684 (O_1684,N_14507,N_12265);
nor UO_1685 (O_1685,N_14448,N_14522);
nand UO_1686 (O_1686,N_12799,N_12078);
or UO_1687 (O_1687,N_14667,N_12270);
nand UO_1688 (O_1688,N_14571,N_12726);
or UO_1689 (O_1689,N_14777,N_14627);
nor UO_1690 (O_1690,N_12881,N_12203);
and UO_1691 (O_1691,N_14944,N_13275);
and UO_1692 (O_1692,N_14162,N_14736);
and UO_1693 (O_1693,N_13693,N_14713);
nor UO_1694 (O_1694,N_12155,N_14190);
nor UO_1695 (O_1695,N_13452,N_12478);
and UO_1696 (O_1696,N_12745,N_12502);
nor UO_1697 (O_1697,N_12530,N_13167);
nand UO_1698 (O_1698,N_12483,N_14619);
nor UO_1699 (O_1699,N_13239,N_12952);
nor UO_1700 (O_1700,N_13499,N_12864);
nor UO_1701 (O_1701,N_12302,N_12890);
and UO_1702 (O_1702,N_13090,N_13245);
nor UO_1703 (O_1703,N_13186,N_12719);
and UO_1704 (O_1704,N_13270,N_12107);
or UO_1705 (O_1705,N_14788,N_14626);
nand UO_1706 (O_1706,N_13368,N_13695);
nor UO_1707 (O_1707,N_12015,N_12160);
nand UO_1708 (O_1708,N_12861,N_13342);
and UO_1709 (O_1709,N_14765,N_13587);
nand UO_1710 (O_1710,N_12892,N_13296);
or UO_1711 (O_1711,N_12118,N_14302);
nor UO_1712 (O_1712,N_13014,N_12022);
nor UO_1713 (O_1713,N_12680,N_12543);
or UO_1714 (O_1714,N_12460,N_14094);
nand UO_1715 (O_1715,N_14767,N_13137);
and UO_1716 (O_1716,N_13052,N_14983);
nand UO_1717 (O_1717,N_13970,N_13971);
nand UO_1718 (O_1718,N_13698,N_14065);
nor UO_1719 (O_1719,N_13821,N_12194);
xor UO_1720 (O_1720,N_13477,N_12207);
nor UO_1721 (O_1721,N_12227,N_14934);
nand UO_1722 (O_1722,N_14676,N_13257);
and UO_1723 (O_1723,N_12375,N_14765);
and UO_1724 (O_1724,N_13072,N_14616);
and UO_1725 (O_1725,N_14400,N_13035);
xor UO_1726 (O_1726,N_12356,N_13238);
and UO_1727 (O_1727,N_12816,N_14089);
nor UO_1728 (O_1728,N_13411,N_14667);
nand UO_1729 (O_1729,N_14134,N_13155);
nand UO_1730 (O_1730,N_14838,N_12379);
nand UO_1731 (O_1731,N_13074,N_14634);
nand UO_1732 (O_1732,N_14557,N_13236);
and UO_1733 (O_1733,N_14786,N_12370);
or UO_1734 (O_1734,N_14865,N_12859);
and UO_1735 (O_1735,N_13554,N_13135);
and UO_1736 (O_1736,N_14780,N_12617);
nor UO_1737 (O_1737,N_14416,N_13521);
nor UO_1738 (O_1738,N_13789,N_14524);
and UO_1739 (O_1739,N_13774,N_14574);
nor UO_1740 (O_1740,N_12465,N_12399);
and UO_1741 (O_1741,N_13084,N_13296);
and UO_1742 (O_1742,N_13974,N_12970);
nor UO_1743 (O_1743,N_13046,N_12109);
and UO_1744 (O_1744,N_12717,N_13828);
or UO_1745 (O_1745,N_13573,N_12590);
or UO_1746 (O_1746,N_13991,N_13007);
or UO_1747 (O_1747,N_14633,N_12617);
nor UO_1748 (O_1748,N_14150,N_12054);
or UO_1749 (O_1749,N_14609,N_14285);
nand UO_1750 (O_1750,N_13053,N_12830);
nor UO_1751 (O_1751,N_14738,N_13863);
or UO_1752 (O_1752,N_14723,N_13708);
nand UO_1753 (O_1753,N_13969,N_12824);
and UO_1754 (O_1754,N_13409,N_14054);
and UO_1755 (O_1755,N_14512,N_13545);
nand UO_1756 (O_1756,N_13690,N_12624);
or UO_1757 (O_1757,N_14995,N_14749);
nand UO_1758 (O_1758,N_14143,N_13978);
xor UO_1759 (O_1759,N_12198,N_12124);
nand UO_1760 (O_1760,N_12530,N_13372);
or UO_1761 (O_1761,N_14904,N_14833);
nand UO_1762 (O_1762,N_14400,N_14517);
nand UO_1763 (O_1763,N_12130,N_13179);
and UO_1764 (O_1764,N_13458,N_12832);
nor UO_1765 (O_1765,N_14469,N_12770);
or UO_1766 (O_1766,N_14681,N_13656);
and UO_1767 (O_1767,N_12649,N_14734);
or UO_1768 (O_1768,N_12194,N_14765);
and UO_1769 (O_1769,N_12627,N_13406);
and UO_1770 (O_1770,N_12722,N_12358);
nor UO_1771 (O_1771,N_13418,N_13097);
and UO_1772 (O_1772,N_14193,N_14952);
nand UO_1773 (O_1773,N_12679,N_12212);
or UO_1774 (O_1774,N_12836,N_13129);
and UO_1775 (O_1775,N_14362,N_14351);
nand UO_1776 (O_1776,N_14799,N_13946);
or UO_1777 (O_1777,N_13125,N_12632);
and UO_1778 (O_1778,N_12764,N_14971);
and UO_1779 (O_1779,N_12568,N_14348);
nand UO_1780 (O_1780,N_12827,N_13814);
nand UO_1781 (O_1781,N_14094,N_13502);
nor UO_1782 (O_1782,N_14265,N_14612);
nand UO_1783 (O_1783,N_13428,N_14524);
and UO_1784 (O_1784,N_12298,N_13884);
or UO_1785 (O_1785,N_14755,N_13722);
and UO_1786 (O_1786,N_13194,N_12185);
nand UO_1787 (O_1787,N_12808,N_14622);
and UO_1788 (O_1788,N_14859,N_14121);
and UO_1789 (O_1789,N_13374,N_12235);
nor UO_1790 (O_1790,N_13140,N_12153);
nand UO_1791 (O_1791,N_14935,N_14639);
nor UO_1792 (O_1792,N_12243,N_13235);
nand UO_1793 (O_1793,N_14282,N_14091);
and UO_1794 (O_1794,N_12174,N_13786);
nor UO_1795 (O_1795,N_12399,N_12957);
or UO_1796 (O_1796,N_14333,N_14303);
or UO_1797 (O_1797,N_13058,N_14888);
or UO_1798 (O_1798,N_14375,N_12793);
or UO_1799 (O_1799,N_13688,N_12055);
and UO_1800 (O_1800,N_14260,N_14573);
and UO_1801 (O_1801,N_12079,N_12679);
and UO_1802 (O_1802,N_12461,N_12724);
and UO_1803 (O_1803,N_13059,N_13583);
or UO_1804 (O_1804,N_12436,N_13710);
and UO_1805 (O_1805,N_13829,N_14241);
nand UO_1806 (O_1806,N_12874,N_14185);
and UO_1807 (O_1807,N_14416,N_14696);
or UO_1808 (O_1808,N_14129,N_14119);
nor UO_1809 (O_1809,N_13868,N_12352);
or UO_1810 (O_1810,N_12456,N_13122);
and UO_1811 (O_1811,N_14319,N_14958);
nand UO_1812 (O_1812,N_12561,N_14772);
or UO_1813 (O_1813,N_13536,N_12814);
nand UO_1814 (O_1814,N_14228,N_13264);
or UO_1815 (O_1815,N_12008,N_14017);
nor UO_1816 (O_1816,N_14925,N_14099);
nand UO_1817 (O_1817,N_12361,N_12234);
nand UO_1818 (O_1818,N_14491,N_13470);
nand UO_1819 (O_1819,N_12679,N_14733);
and UO_1820 (O_1820,N_14161,N_12943);
and UO_1821 (O_1821,N_13067,N_13886);
nand UO_1822 (O_1822,N_13066,N_12853);
or UO_1823 (O_1823,N_13784,N_13598);
and UO_1824 (O_1824,N_14868,N_14087);
and UO_1825 (O_1825,N_14749,N_13962);
nand UO_1826 (O_1826,N_14981,N_12236);
or UO_1827 (O_1827,N_12045,N_13994);
nor UO_1828 (O_1828,N_13791,N_13375);
nand UO_1829 (O_1829,N_13097,N_14483);
nand UO_1830 (O_1830,N_12121,N_12970);
and UO_1831 (O_1831,N_12033,N_13205);
or UO_1832 (O_1832,N_14686,N_14792);
nor UO_1833 (O_1833,N_13632,N_14589);
and UO_1834 (O_1834,N_14937,N_13284);
or UO_1835 (O_1835,N_13261,N_12382);
nand UO_1836 (O_1836,N_14100,N_13297);
nand UO_1837 (O_1837,N_13861,N_12624);
or UO_1838 (O_1838,N_13546,N_12021);
or UO_1839 (O_1839,N_12658,N_13187);
and UO_1840 (O_1840,N_12927,N_12204);
or UO_1841 (O_1841,N_13660,N_13756);
or UO_1842 (O_1842,N_14229,N_12682);
nor UO_1843 (O_1843,N_12361,N_13205);
or UO_1844 (O_1844,N_14679,N_14923);
or UO_1845 (O_1845,N_13247,N_12470);
nor UO_1846 (O_1846,N_13026,N_12926);
nor UO_1847 (O_1847,N_13815,N_12240);
or UO_1848 (O_1848,N_14890,N_12932);
nand UO_1849 (O_1849,N_13483,N_13762);
nand UO_1850 (O_1850,N_14990,N_14212);
nand UO_1851 (O_1851,N_12693,N_12422);
or UO_1852 (O_1852,N_12770,N_12580);
nor UO_1853 (O_1853,N_14282,N_13820);
nor UO_1854 (O_1854,N_13922,N_13694);
nand UO_1855 (O_1855,N_12517,N_14493);
and UO_1856 (O_1856,N_14004,N_12898);
and UO_1857 (O_1857,N_14350,N_12190);
and UO_1858 (O_1858,N_14007,N_13992);
nand UO_1859 (O_1859,N_14097,N_14943);
and UO_1860 (O_1860,N_13004,N_14885);
nand UO_1861 (O_1861,N_12317,N_14981);
and UO_1862 (O_1862,N_12875,N_13925);
and UO_1863 (O_1863,N_12659,N_14626);
and UO_1864 (O_1864,N_12095,N_12870);
or UO_1865 (O_1865,N_13031,N_12297);
and UO_1866 (O_1866,N_14172,N_13006);
and UO_1867 (O_1867,N_13228,N_13406);
and UO_1868 (O_1868,N_13212,N_13840);
nand UO_1869 (O_1869,N_12387,N_13501);
nor UO_1870 (O_1870,N_12445,N_13562);
xnor UO_1871 (O_1871,N_13451,N_12953);
or UO_1872 (O_1872,N_12350,N_12625);
nor UO_1873 (O_1873,N_14889,N_12066);
and UO_1874 (O_1874,N_12649,N_14387);
and UO_1875 (O_1875,N_14761,N_12927);
nand UO_1876 (O_1876,N_12442,N_14178);
or UO_1877 (O_1877,N_14165,N_12602);
or UO_1878 (O_1878,N_14158,N_12414);
and UO_1879 (O_1879,N_12740,N_14334);
nor UO_1880 (O_1880,N_12530,N_14703);
nand UO_1881 (O_1881,N_13603,N_14959);
and UO_1882 (O_1882,N_13588,N_12762);
nand UO_1883 (O_1883,N_14685,N_14317);
nor UO_1884 (O_1884,N_13838,N_13964);
nand UO_1885 (O_1885,N_13723,N_14939);
nor UO_1886 (O_1886,N_12153,N_13825);
nor UO_1887 (O_1887,N_13697,N_14828);
nand UO_1888 (O_1888,N_14687,N_12657);
nor UO_1889 (O_1889,N_14513,N_14680);
or UO_1890 (O_1890,N_13901,N_13181);
nand UO_1891 (O_1891,N_12956,N_13207);
and UO_1892 (O_1892,N_13045,N_14629);
or UO_1893 (O_1893,N_12330,N_13601);
or UO_1894 (O_1894,N_14960,N_14921);
nand UO_1895 (O_1895,N_14397,N_13045);
and UO_1896 (O_1896,N_12692,N_13852);
nand UO_1897 (O_1897,N_13852,N_12059);
or UO_1898 (O_1898,N_13711,N_13443);
and UO_1899 (O_1899,N_12641,N_13100);
nand UO_1900 (O_1900,N_12759,N_13374);
xor UO_1901 (O_1901,N_12514,N_14851);
nor UO_1902 (O_1902,N_12940,N_13634);
and UO_1903 (O_1903,N_13915,N_12281);
nor UO_1904 (O_1904,N_14725,N_14013);
or UO_1905 (O_1905,N_14725,N_12790);
nand UO_1906 (O_1906,N_12645,N_13434);
nor UO_1907 (O_1907,N_14417,N_13169);
nand UO_1908 (O_1908,N_13369,N_14990);
nor UO_1909 (O_1909,N_12789,N_12289);
nor UO_1910 (O_1910,N_13130,N_13355);
nand UO_1911 (O_1911,N_12557,N_14769);
and UO_1912 (O_1912,N_14621,N_12834);
or UO_1913 (O_1913,N_13722,N_14518);
and UO_1914 (O_1914,N_13739,N_14757);
and UO_1915 (O_1915,N_13496,N_13874);
and UO_1916 (O_1916,N_12517,N_13652);
nand UO_1917 (O_1917,N_12826,N_14891);
or UO_1918 (O_1918,N_12726,N_12028);
nand UO_1919 (O_1919,N_14215,N_12902);
and UO_1920 (O_1920,N_13547,N_12118);
nand UO_1921 (O_1921,N_12462,N_12654);
and UO_1922 (O_1922,N_13873,N_13735);
nor UO_1923 (O_1923,N_14482,N_13652);
or UO_1924 (O_1924,N_14795,N_12431);
or UO_1925 (O_1925,N_13211,N_13073);
xor UO_1926 (O_1926,N_12833,N_13433);
nand UO_1927 (O_1927,N_13686,N_14157);
nand UO_1928 (O_1928,N_14681,N_12253);
or UO_1929 (O_1929,N_12766,N_13896);
nand UO_1930 (O_1930,N_13456,N_13363);
nand UO_1931 (O_1931,N_13247,N_13890);
nor UO_1932 (O_1932,N_13625,N_13476);
and UO_1933 (O_1933,N_12571,N_12091);
nor UO_1934 (O_1934,N_13644,N_13567);
and UO_1935 (O_1935,N_13293,N_12417);
nor UO_1936 (O_1936,N_13035,N_13640);
nor UO_1937 (O_1937,N_12294,N_12624);
nor UO_1938 (O_1938,N_13844,N_12279);
nand UO_1939 (O_1939,N_13273,N_13301);
nor UO_1940 (O_1940,N_13627,N_12665);
or UO_1941 (O_1941,N_13117,N_12768);
nor UO_1942 (O_1942,N_14124,N_14245);
nand UO_1943 (O_1943,N_13774,N_12259);
nor UO_1944 (O_1944,N_13222,N_12502);
nand UO_1945 (O_1945,N_13135,N_14256);
nor UO_1946 (O_1946,N_12369,N_12078);
or UO_1947 (O_1947,N_12566,N_12965);
and UO_1948 (O_1948,N_12785,N_13963);
or UO_1949 (O_1949,N_14410,N_14666);
xor UO_1950 (O_1950,N_14753,N_12151);
nand UO_1951 (O_1951,N_12345,N_12883);
or UO_1952 (O_1952,N_14681,N_13919);
or UO_1953 (O_1953,N_13066,N_12289);
nand UO_1954 (O_1954,N_12145,N_13045);
nand UO_1955 (O_1955,N_13179,N_12304);
nor UO_1956 (O_1956,N_12416,N_13119);
nand UO_1957 (O_1957,N_14485,N_14548);
and UO_1958 (O_1958,N_14694,N_14710);
or UO_1959 (O_1959,N_12562,N_13100);
and UO_1960 (O_1960,N_14974,N_13613);
or UO_1961 (O_1961,N_14141,N_14355);
or UO_1962 (O_1962,N_12528,N_13789);
nand UO_1963 (O_1963,N_12094,N_14320);
nand UO_1964 (O_1964,N_14366,N_13027);
and UO_1965 (O_1965,N_14966,N_12703);
or UO_1966 (O_1966,N_12232,N_14273);
or UO_1967 (O_1967,N_13938,N_13607);
nor UO_1968 (O_1968,N_12696,N_13879);
and UO_1969 (O_1969,N_13345,N_13593);
or UO_1970 (O_1970,N_12145,N_12124);
or UO_1971 (O_1971,N_12270,N_12698);
and UO_1972 (O_1972,N_14979,N_14233);
or UO_1973 (O_1973,N_13958,N_13267);
nand UO_1974 (O_1974,N_14642,N_14101);
and UO_1975 (O_1975,N_13079,N_13095);
nand UO_1976 (O_1976,N_12425,N_12809);
nand UO_1977 (O_1977,N_12623,N_12465);
or UO_1978 (O_1978,N_14239,N_12548);
nor UO_1979 (O_1979,N_13005,N_13889);
nand UO_1980 (O_1980,N_14980,N_12131);
or UO_1981 (O_1981,N_14875,N_14009);
or UO_1982 (O_1982,N_13725,N_13123);
or UO_1983 (O_1983,N_14771,N_14044);
and UO_1984 (O_1984,N_14828,N_14171);
nor UO_1985 (O_1985,N_13860,N_14617);
nand UO_1986 (O_1986,N_12065,N_12448);
and UO_1987 (O_1987,N_14715,N_14314);
xnor UO_1988 (O_1988,N_12071,N_13052);
and UO_1989 (O_1989,N_13085,N_14061);
nand UO_1990 (O_1990,N_12469,N_12069);
nand UO_1991 (O_1991,N_12638,N_12611);
nor UO_1992 (O_1992,N_13331,N_14929);
and UO_1993 (O_1993,N_13148,N_12943);
nor UO_1994 (O_1994,N_14331,N_12320);
or UO_1995 (O_1995,N_14379,N_13477);
and UO_1996 (O_1996,N_14896,N_14805);
or UO_1997 (O_1997,N_12755,N_12450);
nand UO_1998 (O_1998,N_12026,N_14749);
nand UO_1999 (O_1999,N_14038,N_12829);
endmodule